`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
GEfvXn+CYJWnRpahCRd6lGW2ZOPGm+FvVePMj0wm98TtxkexpqjKimyYHP3tDAXfLzzZxks9U4G0
VEr/MFT2fQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oYvnUGXz/ynKVacP65M/XJqOmbIsKVnpEWci3of0oRPZ8FIAu8fomjmAPl1jbMstZtZ1dVpNyW/Q
9SNzooLfc/eiU0VbxthuRR1VdtTNKiMhfR+pJ4ynS0vbh8JUynCj3fW4+NvFnC0pVaI/BmRiggNX
Wwx4OTANjlKG0g4vvqs=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
UajxnPAMvL9P66D+gvtZtOWSWQosuM22jDUJow37J9t3wEl/qpKxMIm1oYL76aKKPcyM1hkouVPV
R4bVz92cs3STyEmW6AQaFyPbutUJKQ1DI5IbxzDP5QsxYPlS1726brZjmVOPHLhqSHftfV1+yW8j
9cISe2a7AIpiJw2gHWU=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kkWKcNfeQRsnys921mm7wDIkarrnlnOR5BOd2CHwJ+0MOeaI6NDXAlNUD0il0RWAPltNXC8cu0tw
jYePAHWicDk6CGzMlQ59CxFKMd/ygzMUiOhHJCJgYjuxQ/YHylF/bBrVR8ALGL94k784C5pXEC0Y
/HYJ3Le4qQbBGe9bOZG5X1FyVqZ5PaLrUwVD0ppRfhiVe0Nd6wOn/8Qba3PIksAaN9U9uthJUHnL
fYxbTEaNjBJ8KO0WN6ZXlLMgXFVJABum2V2hq131C3Hig5ebSbUnH74FAMTUoyyWERWs302lOYXp
IF6bi7NJ13vZo8Ya5thIzJcIMvvLr6McCwM/0w==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Wjiw4qdfvbJLOPknf/5meBgqJxV3tV3yfLBiYrXnouh3dDe0ClSR9LCu3a2cOK24iS0ivP1XnPQv
PLtZuoNfB/8ohGKtz2wdNLS6mAWGT4piCe7tFh7IoPq94zR31KPKOg5LiDP1o2JOkrvZzfEEoYij
jfumJf3qONCPzIQijSWh2kl6FWX/AF/xokanwRLCy51gLSKAXZiK6wDuXgWK9cMxlw1ZPdWrjLiA
pr5w5o1bOGWBUXlrb+z6QYU2sHPZ9LzhS5lS1CuQtsEdO2muUgYbzKn5aGMeeFnTgDG00IxufWf4
0rhSdVMcY/Q09EPMJd/AHEoqlx2GvcdbY3jxxA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
reFJr7mSlypn/enU7H5TZvAI/ZyTp9+kctgFsmumqE7GOBxqSUowG6MGAaQYIE1hOE4uT3VBFWJw
iQsxWtnwhq9VwskR7NbSyN5SPFzDEVDI0NAwcjLNEP8WcGxI4mtuwNaIDEKTKZM76+MTJ4N6FkWJ
ngmihXto3VLJs0AE9DrVsluixT/LsxkGIzuVG0wNsUsx1UoBoUOqyhKp2a2TITKIAUuONBlvWYPm
PSR3aSnsCKnaU8ongyZz0K2Okj0Sv2V3jEK0eRsg49lcZyCHBuZOYWvaFZN+EgYasLjS64yuj9eb
ucldGP6eUfbVRTANgpxKv3RolOBABC7o7hSngA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135936)
`pragma protect data_block
BnAR5YpZ8O0NjodbyjsOzg7Dq7Y2Ud+fn4ebewNNqxPk/okNCmPCwG5sot0e8bM9l/1rBhLN4Shy
JDYN8Yf9NmRs76TshyHCmwQO/E/CxijOX/s2srzJw6rw4QYclzbWsYVMIa60wk8AEMGUtRgI3GZo
VF5Tauj/fHYx7Q+eVGVsAae/PRUfh1jseGHIbzBbg67ugz8hFwZwpgMepA5JLuRZJbpxu9TjbJl/
4B+P+NVohiSNZVFWMjLa/RnB6NuktnNxxqhcWymIHcYPOOdFuyj3iPZH7tBdWWr89ybeJaePUdle
Dha1IXBC3A50lZLU6JL464gLWcxk/6KNAkd9nEC+QfhIcUmruHxzfY7RwxZk7ZWWGQmvya8IS0Qy
w705ZjMgx+Knw6g3geQgT1Hfa8MlfG4VmitGTqwUGhlu4LXqH+OLPiPpDP3OsHgkgXbI6C2kXGC6
XHfpabyaEyHfprJkTVfT/6+OTEBoaJJgZ4WyDsoJWw3G9OA3SrlidfwZoNWwCkqcTbDT6oHsg8bw
VGQnebwCr+HCWbLFgFYgwBFJ1B4sw8rz16fB8z2vy2AZT956x1a2dewVxC0mWPtCRE1Y6OC4JPqV
4r7IT3G582FV3Z0Jzgju1Qn4/nqA9ctJYBWNaTxuG5WqqWkna3cX2eZ7VQZra9CMdjG1c8tB/eaY
aL+OhyftQXpS1v16yaoeFMoIRj5Uoy7P2v2LyVhd+N9GfgoU+8iS1JDQ5N1H4nrX5B51byvKlqvN
JvPV0FGtW56vEcIOV7Rf0GtJkD8B/78UYC104Q1m49jCKkNufnCTylcoJaYjnj/EXqhJhrZ8Vd5o
lQOE2kCTyKvqjOyMJN+xqVOCU30iDfVityI4Xw1DWc1nbILXCWIx+QSTc3oGlNzbbvBkgJpDEdpF
8B/NfpeWM4SQTyZtIKfCyJ9D/jcsZoo1mtOT5coYB0Mz0M2fdahi7rXGcxiuTqpvAup0gQs29+Iw
MjG/yqH6Sp1ySRk7uCik65Dvnh40p1m55O9W0KyxpU242zRW0f1KttFUcJSXr8fjpa4qTUjf4QCh
euCx+Qew/GGI2eHbhI5mhfqeAxuadP6hggKq6EaBY1FfHFv6Wbwf8cFSBKmToaY7j8aNgs4mBnen
uHUj7qA6IkvzSV8xjCPsYQ97x3+yPrdi0U5DXKLX31Hl08lYkYx1RJ1k/xIPaK1zA7QZMUCpqMEK
DcB1G5lQzPIWMw0MUcRTad7WrcOzNRmyXxBYcAWx5n+aMOkMqZxX43VkvkYssWgSp5SwDqHrCbzl
M7EZI7bNy7lfXQJ6SN7hwEgEoPDB6va9EQ3XkPez00mRvYLvOcI9t2zUgiumHhajVJkZ+2fnZTv+
21XhboBMqx+k+Kpcs9TyMUnnjYi3m3AxgfNs4KRk9m82dGooDltlGBXscxdkaLzra+BRWdV48yCz
QmTVQGPrk6Ns2v4LEnWrcla+ZW+j1c8XXU64UJ2DaQbV27Zz+i333jV1MZFKs/SiBZ8URe3N1NTd
BELHVAtU9uPUkYTfPQl9ET7rE1aiglbz1wccUb2GVL6PEz3cYNj1pK9eVZIZ0fUPWEVe/9D2qLUj
HIPs39aY2/j5KL6Og19HYizknLOHB/zyUsXDp/50RLOEYuQRsaNwSy0EIisfY1806VJWbhCc1XTA
ScSvFccvk2lwt+1mhuN1skPrtZxoJXLKJWnvhCnq8O6dXRljJLEkNvmT0G71yQ7uUw4zEuPbORHN
YoP8Mgyv3CNbvxN3LtlFJ7cnxYnIaM7emJvT9BqD3LlQAsZsIIJvG5j7eCdV2EPaII5v0NAeQXCN
DSvVQOIBisU/ktoeGpgMSUbOpti7WgT0oc2US10BcWf6+AmLeeeiYlfLcf0UXeaUUkY9z8FJTjos
yRY1qJFLNrgf1JIuGCUYh7RpeQHT8gvF7SO8dw7Ig0cEfDEAXg0dSQkp1CetOMWR4fycSwdxCToC
o3+NIQJahhXn+c7T5rLOQs60q0E71p9BfQ6hqP/dMVHKzEt/zOxIukOyc6h8OgTJNuyW3oJ7sM1W
zEW147R0fQUZyMe4iNstCHENu9lixPkD8BJ0D8fiVNDpl31x49XwolQ12A+STFlHVGwRziEq6Oz3
SXVLUT5+OJV7aPuDaOnm50M4ksXpa5MPPHmrYL+FxA0xCz7wT540693PMpvGGcBaQlUt5ITcaukq
lKQepwGjnnmRIZqNtFqLKahjyObUoyg35F2+PX1qJTu7zZ0d6gMgHq3qR6FshTBBvbwZOfazJqrZ
CNIkx+4jxAu/FSJ0OfWjNkyvd96TFroFxz+Sana/TRK/jbr22Qwjm7IAnlCF+5+i47bgGFPlitBm
yl3l/x5da14aObo6CLrZRuchw22HSDULaCixOrartFjAxlsPccXMc5yoGZazxjqoqBGR43BrC6vZ
X2mi2R0THBiD/zg3ZXK00DywfS0gF8/mLeOc5ihDSVjVCiw9voaSdRhB91N9t5kbskJMqX3gu72L
agjWIL4k80atA2KDe/ARaAbQA0gkNuO8azbcROUtg5lF0AdvuR+i9o9OIYkBs4+Ot3JFjFyNoyWQ
0CJ4imJW+weObA9TBc8h65pGgVQjLgSRpVKqsuVQYt7jGMNj3g4yTpYOakqqk1b6p2GKAVoAVoSZ
VAFgfs7gMt2aEzCOb3L/4LRmPW+2nq9RaqGL5a59HgdE96KKAJpeMA8Os90R3UQxm19u/HeTwTfV
TCN4JJANo4PQEF9dWAh3ldqmKkUyJT44mlqFe7R2mLcY6uZWfEVixlAUXubIK8LFE+DXvCeocGdr
B3EWkGyrWfx6i5jhnxdJSNAM7G7KUGhtXRYEdqpsmuNN+XrsZg2HgvH6DQmvGa66O4YGAe+DA9pT
x/Mln4A7Zb34JNxBo8VgrNokPbmh4Jry0r2RkZKNjgR994aFLDm3boJt7MRus2i7Z1WxpgkNmEId
3Bjfy48/VERatI3IP2syLEne4Cc/hcyjWcw9Zga5VVvLMJTdSn26Dq3uAcSY5Vsdpbg2tYcgocGE
67qIw/Bp+UDw+031u+yWTd+4sPj4tWn/vRtFA5S+UGeU4DUHHiuQ7n1w79sh8GSirRJmpWUvDzUv
jjAkHfPLkiEnjKHhRdDnB44Ws936Q+P8k1IbqXVTMrxyAfKmkhPLqW0YafEzv92MPt2CVWdCy3Ve
PH++0ES8x1yVpkPWQ91sjZ0yyoSHcn6PucwIAz//+OkxUrGPHfeCSNxkLdERrhLtZPuPT/sHuYE4
p2BjcGPcPlisxUWad0LAGe/KuTstAbL2AbwqT8KaJ0Cu701pVoLOMeuwiylNsWYuZJ6mNUR26X3x
RgvWwFuLTS09FTQExCrHz2E3OBygBRX3P9y7/osdXqFS+SsE65WCqVmI+ifiZHol7Z/WfVrcaPjh
go6dBGNzURQY0uTS4SxmLZH+leZKwo8amG1zoKfGydxXWqFyUmz8NrYUdn+pQ9h8NCmzcDUYW1c3
F9bCXvKl98SHmjQPgQvCaM/tZOt/75A/masA2TGhdC8RkZw7jvBqoEB43A+3+tjjRGH5D66Ncm08
MPsut91Xe4fFc5OE2sdf2Ya0Bloi16UrgzoBs47nV74WIzcm5++g4sU6TvmC0Lfo+hVnAzOuuYS9
PgAE8LCa9nf7qL3PafDJhRucV1K/LcB3NfB0Cfsrs+2FXd8mV2KFdU/LyklFjKtna9SwelkDYMIi
y+nupuODwRbOBtAuBExZY0HFZVLFegof9TeTEgQ+KUWR3nFIyA48htW89MWs5iewag+9E/5tyS16
MyPrllj+tzYJSxM8FBPP5UW1ODVNvxivbRPbHiKMqryzNBw8sM7dZEuf0vqNLGSyJJfC8hh/X0+t
K4b5qBL/YJMfaDcBDrHEzXnnvym+C9ti/9zIjJdH6P2bHX9BCMY0TPV4Wg2jrZJ+4O4NSdIT9kuO
bz/fFHb9bdgZrsFf9Z/qyWn6cFVWvcIEsgDHfwFoma8ENSYaGcivEP23SUA2JK2a+eZjfg5Rmx75
sVxF1Zz4aVXIbXFZcgguX7FjW8gqgoTPMzo+GUCK+/MxGERVDqhpUU5A+ON0zJls3P6K6Ta2RO1G
Cof2GBQYPBsxbL0KoSR6aYMxtcBZnllROkFrAOkBOmuSm++KHZHR15qdelLBdyoBj5MwrtIMEUbK
XXlrNad8chMFR1n3dvyhFi2qrDl8yt+698960pnw6rhaRKrHHW78iBd9vuBLC8FT1Urv3vp+O7Of
FNiNdSv3dpQMWSCZ+yQacIOTCmUFVuIUd9LaJEGwZGTMsr+4GlTRySAnyqfnu4zP3Cd6sll5+zLE
/9x+KsknGbOt6pXgLj6BpNFTheANBsoMmpdtXFeiGXxeOMy3CzwPk7ZkjSLSDPn+qpvwKv3+BSrR
ZJK/jtuaYeHxShWiRdp3EybZ7YXSSADruCZiMB5TD5pl0WP5KC6K78VlgmfRQRn04LPX8zuftN1E
PzKL1qhMWaQqOTLxzoZXupmGo1CC73H/kUuC5v47LxPFNrywUee46wczVuXgeIGjXT/oTtTIlEYU
DOsaRDMalnUB6idmZLaYmu2jxZ78An9Pa4UYRa3ublnIe82+CIbAsfuIpD676a9VKMoAj1H4Fnyz
Y4+v1raCXYaozeSh6VoNVoCgn5ZUEBMv4baBLXQyaBAytkwhE2oMuvt26L4cU2Tab8FdGxoBNy2A
OhU65JajfHaFH6dl9XMW30TCmFD6zE0PQNBpGFf0CnBewo5yyQ4iARTgn9lbp/bAnWZaSS+931Uz
I7gYx2DA6ulOwjF9jVNnUTB0ZZZiTpdqE0sLiF54Em0yaqrmag3JztTyYg9G8Hin/BIdKL+rOwb1
GD4lIQTFFHEL0hfKwnS9hWY7zwmkngFpfR7fRKRodrvb8xoL1vz58qFhvM94pYMEAxFoK4l1RCTZ
8/gxmJmYXYh4xzaMyaK+92+/iKuwYpxsFiMwcuI8/utrOYsLWpaYXIJrnqNhc7shV/+MgPvhIrGa
29TrSgvqC3HWCqnshWPkIAooIaR8AwuUTzJRDY2e6uLweoK+fEM14TlQHjpDUeWMZ0CBEmT6Wt3C
ifQOdzDsJgbnrWedzGFj+u4RDe9nmc0ePJ0MTrv02GsuMnrhaoObiFscor2KADlCdmVYnA7R4s8H
qwMJAxBwhu9w19Fae0acoPqljR8iacfuAPussdMWCVoSp43F6oRreLP1Ncm8PyfFU/tvP8JpiwqS
MaHF1YpTvv2at4Wx6r5XGEs9pSKI6HjryZ6FHTPwlwVCIt3SIS8dBdeRhHlbuiUhAR3ZDol8X27G
GemcdWS/W8CbtWJlKG0eAGxAkHJNvQLNc2utMhA/6q/99ttNfmg+oP6j9dNV5hZwQHNhJYtxNwDR
9++lF2X/tI7ws2ik/a8LhxuX1jLfzz/Ji/apfEAH/YQU3eYA+f7Rctjj+uBr82Ms8y1uqt2KMY7q
TJgMEofNPqNdhkJSIDFrVITcCRVDlDAynfp3ho0kEB7va/AfWeUzLBHUGSRbSXxTbDHLsuHgBRKd
op6o3Ypmc1C3C8bk0JyL58ylScw3NRFgiaH1nH4EPleWVNVsAw5VITIsIC1Cz8944K99QkVMMb8O
S3e2jrMliVq1zjH01+dWpjwtdLDrn+4apXGUkQZhChXhbK8nK/IrYXGR7rQFmOd2Bpjwdh6h30PJ
P9mw7Icqq6txUPEC1PBVZt6wZRW+L2WSzloK1wcymh8iZaz7fFHOFloU+NNML6ol9fGyW/P+ueNH
JyeYDXOyDOVc7N3YZNnyYdvk4lihmCpmRsz5v0g8WRXwczbvCxgXXhAk78PadbxmdfhKvzPYqJB+
/7RJaV1seAbbS+TgAICLsoBPjt0ehzoCl5RPhVb+EoUl6HO3BB6wVIgaQnkikh2H3ZdEHHoOhOM2
Qfbu+yujzBbc4UCXPGKpWBEhRh9CbtpJsJ8/bV8R+N9hlZnf4UYVqTjOzNvYAt7lalgub8hXCUJk
fk2KesKxfhShKwMGUTg5tZes8Tni12Ng6sKrRywBApTT7+aL6UrsnAVYkLD5dSdEdKbJksk38tkt
voNUVdHxTfh8Une5rZ9kv3BWNiS5DGNgQLSye8HcWtnwZPW5SvddivpimSxCPmvXKnbRjiof6kx4
shxn5AEJ6HPAn1sJpomHtbxkDSW18YH6r93khk+PwCLq70sxChON5qamdQ5dUez3oHLs8rOYpl+9
GUPRJGEs+Bet3MtD1pyMOVDklOBpCCyfbIXbwlwCRsKkRwqxk8iuv1nTuuA27yfZoGUQcvThoHQn
7Zq2UOE0a0hi15ofmtq8ODfYTV7lJdASiIbXhK2hShn1Nrhk4cX54006h3QYYXuxcSWTvBfHAPjS
13TFtqRJqS4sgmrXHO5nthjPY145RVYSWMPlqKjiRCFGXCGJwPtk2J92SqfoxOp7efl+lhGznE/W
sRKUCCVJuH1vU8vngZQ+f+Gylbsb8b/8LK8R85npdozQFaVL5J7FtwGMQO53sBPPr4gB1rORvMyU
xYrm0ntexoEZ6hOV1p3MX6Up+I28eslJuEPc9bumHHnbI2TWEFx1jUbHlBXSrwcv9hHPlpcaoChf
6cRsHAzE7s/TUiZWfQCbSLuroHGJ7LepInum/Xyvo0rsrW4pg4jBXSelTF269MAMN4jQCn1C6Qvo
FNTL9GFK1MMUQvkCrgYoi+MUmQmSAla6snTTDG6YjVUIJYJOnP/EMV3tWZxHPiwfWBtwj/pXRsr3
C54L41Jotd2EFK7N/v5ag8zQFxv4AnJs7FxhnyDmDSvymPaTw/xhMp2GjjBDRN38FTbat3R0ZbnA
moZcCkwR1cMiUUi6BCSNqli3NjbOKMiV3tTi9fyoEvEchDgfhGUYdR0b3imYqIiyAOerDEvzDRqI
TNyNBYE0fqXM5bzw+UzOt/FNU8V2nPhDNbczcoevPLu3hXZfRxvKYZDeHu06zVOVWMzTNkee6Kp6
meeto6YN34JnRFQ2s10CVSSEWOjmk6uctkxnka6e7PfFJjmqlykXx9MlkwZ0msfFuGwlX3G42IDC
viJGvrWSuG5IvNtpWqqaWPvMsx8lgjK3xpcjonlrGeZv+3bKoTqHhtkwQLWhx66TN4xJ30chv3Tq
2Sry+hlwVvWZdo45AUKBpNn5/MoM/tzq/Jg8akBa2S6UfB0lZ7G0erzPINn2NeAxuKpKvGs0pCHG
71kyinhRRo/ePpChSoFWWoUytWTsErQBU79QmdF9coco7YflgL05CV0uaQcpvw4oP2kJYcHTRkqu
oNmPd7M2qBSuQPofP1wg/GVwav2iFrNcZz/DDmEluC4dyhh2bs04FdfJOlQJtvGmm7xa2TQTnVWl
Wor9YMcwtC8+TsLZdZofYW9jHCp52SiGJs26WEGJsZKBJnytl0Wi1f/wFvsIKQdg2dmcdUgjAsnE
MiJAm/T8Qr2s3jpSsLq+S+XE5f6esuZHccjdwja73hVeQUbb2tB+jFeO7TCnoCUjepDEGqV3Tein
Oop82qibvES7hOe0buDO/d+xDHI2N2g/hgUlj2rssE7kCjE3UfSE4xAjyH2sAgdzF8R8PSvT3xHG
cb0fTHsWkkshvnVSRXMpfzstP6qiyexFO+aDoiOEImDI9U+m6yIMjA9Nsz9ejhcGHnq+yuR7SXNO
93BaeexUhBBx7ex8yubyCnTd4N0Rq8G70uADlMg2XQXbflOUDUUUOixM6CO8+utLut58TmWz1iTe
7hNO0TVnXgQ7xXtC0YH5qAPZ3PJvS3h3see1ajAP898t8ZK3SMNmZ+e4PgcY88JOzjahWXPNyO0V
mubNgH694sQHdL470UGmo6znraF48yFsH9QWNRgVhMD+DMIB9yP9U+3y/+YaMeBrTr51zR63v7cs
6N0nuBMJo4UaXWppZnMdwVI/iDyvWzh1+1lrOUBOLwYPM6r4ofM5MvQm8/DfUMZq7RyHxE4YjpN2
MTeCiBC0zwei8eoCzEpVkFTgvP9IIvOqQcqjFxykY+UtSFWQzD+wih8nZ379faoRzjeAGDY6b8wh
wyv2R02GJ+Xfsmq43lJOzCuemaHwcr0nwv4451SixjyjJpd8PO93hmMfcJ2qyOb/JlSGaWXANZLA
PhQwsjUJw4sJWE8/Jp1Xe0nMrh6xPPyX3s+CEVIRD4ZW1oX7UsqJJiI+1dY1D/XfaqCYdNeH3kPl
c+39HvT1XgO2VxQiJodhL5lN9FTp3B+6YteckNED2glYneoRJpz37RvV0/qGK/ygMj+l8W4661EA
oONkzIASLeU52HcKAN6MD0eFczHlzsntj0z6lUpu37RCFmVw9C0h6QJN4e8ilu/rI/WxybX5iAWR
M1QKTstjWrYI5pVHp5ciDk4jsoRxOfdZaOEOCgZ3khEegvMOQzts8XkvFPfInNCL0UErf1EToUqG
qppOnjCPQuxykkxQmokRBKby7JfRef0o2GpARG6M0yjMUO94f4h98xnX/8Aa77u0pcOnNt2WSyXl
yHtHEsepZYPbzxCvjYB0Q6IN0ukOwgr6vQTgSr/a1hgMBb2mWFNTbnN0YPD3mPc95HG5C5g3FKQ1
ajAVGL5XfCM0xXZVEr48P9nDrw1R0SrcuDwIrSMFP9Q96eut9ISWu/V/7b/Py4Cdg94oe5EtaeUk
DJUUVKMvO4QIGyUmS+UYrkWNWtfQ6+/jFSQpCPycZNGDWaETCZN+krCVe0ubH27RmEZM1ZAmaYrd
2x5MuYrCUIeXd4EfaE//EZGCkbPMijGfdyDzG8FidviNcKnzrg5zQ4mhHyTjEoCgyf9q9r2M+ffc
YvlEG8Hn15lgWFWux5VMSAm4gpLP8eJX5UEkCCG5+rkJvsNdTqwlNKp1cy73ORI8L3DkS9PxLIMe
yMt7gebTEhSLZPehv/UAG5vMC5s8TfdRn8OTiGCpZQg3bLUjxVqOgjacyKASwImS5qKHEXsRrQ2R
1nag3Vw2lh7T1V/Aq7Paojv9VwWBVsh9znLeXArM4Sk05AARnPaX91225oqtk5opioC/YfVWNyeL
V+SVB0iWRWzTY8ir73diu+zHdSdpdHH5/8jr7Oxs58RsM4OJCi3RVZj8SmHwEfLi0Rruk21e8u6s
gLWMcuUSkxWjqAbeomJ8vGk8JPS7lr3cDqpkYjZ3mylyan1kx+DV5rw3RG2zGOJooBewFAWIv+V/
hkkS+0a2LpjiwI0FQgYFX/lo7VsPZS6fwVwk8HjQhWEPfQD1lEgen1+t+QWAjuF7WcxhSGQG94Aa
Phvhj1O45vDxTdTk+pvf0BESLFMOHKwaJ2lYU5s9a682BbmDgyyjHHIz2iy2+VCMtV59UsgYsFb1
eGw7fwg7hCa7oqdd0Ae5+XLv9kquUd1JiySXxlLgVujSFAXuCmc5AW4lEkhS0S3HoQLPEFKNXEX8
T9GE9NFy72Kf7RvXayFF2OamX5soDWz8hju/CgtnuVq3dRAuo+VSo8QWaxuqWjldDCwEcgpJLrD3
NM5shyGoZ1FcCw0DOs8rHn9Y3SWLq3GiZr7ddKhw/I9QYpZUCu4pxHjEqW4y498Q+wLUgR3MIJyP
kwyZ1Z/dfFMDytRGM3rWJEx8gTnX/kqzMeg6gPSavWvZGNTPDOvpfiIWIk3S5aL2oYWLlT0hsbJQ
lpmLNMSMfnho8W2sf0a+SqKM968UyqxlDvovODeXja525oLlZhqZKiXN70QkGhlj/klwjGgtkPoJ
5GmhwmuVqSr7+54rTQrknKkzzJtKNZC7JtPPotF/c+o+SZc3MSWq4+UD4GK1qjrDfKNrH1C/vycc
HnHQX2U2OsCiNDvxYJ7TTt56kvWPKEW0XUEzJ6jFgHczuAv8TjZnPNed4JNUJ8r6gKCZu17dFoPv
oxg4odtmEAAH8gcHm7HTYE4J8rfMtBaCVFoeu+gT03YpuJtwIemrezLZk6fU+DsQx4sSIb/wEM2E
SNFAu6WCvUIrWR/jEsTnHCu9uZN4pfxu+0pdAie7OmYowydxeYacnmeeP1UPhwro/whC/HvLgPR2
Xac3gtbUHxX0FcnzcRYFfVkt7D1IvIrdk4ch+CivUvG/lE0Y6+V7Ifsldq/N3+ANivF7GXRoTgIy
Il02mH7nplcSed63wPiUzKX+dskqT3pSwKHq1e1s/VmjXY5Fd8FN2vmA0xp+CLE+2QsDUheptCMv
QDFl9V/Hl3sC/3C/7YDoXl1snP+Lb1MkYsZp1uVRSSUjwfa+i21LmaiJ75WSHCPQCL8y5eONU9/h
8I5CFwLgkThPYgCs2VqWuJ5CJOdg8aYfTvWrEaWsHwB29tXBJ8aIigKtj+H54hqNmb/f8ftABaDT
EfXx/5n27ZrHH8HAHNH2CIcHkdIyCWlueLxmhQ8i2L6q5FlIS3jtPw5sfljLkW9eD1Lb1SVzwiTN
2LPjMUgWTUFnJq+jLPlXb2l3jB6E3dizFVkBDIuGtp5dqnyZZxNjHnX6qM8PH/V57qrmrAZBdgyr
I36r/mSgab+poiHzAHc9yeiLs5v8WmomlPzu7tfNT6JO7Tc70Qrd+qV32H1QI8mhK7huJg2UuwWD
p0/TexKMfEW3TaQ6yHbKrKzLTtp93uGHKP2MKaaxovSLTwIowsmvwWm1/O+ZmKBEmaiWY5Bunfbq
DgJj8eeD7MnFBZjiWKOVNCK7rs2jih4NzvbVnFSQ4Kps0MlinHhvPPq7TYTLEe07uL9Lw4w9Wk0r
B62AC3MnOyqaQJ2mV/IzgkylFRBwfMi6C2C6rdCfAJJWUJz9w6W0BkhwBOu44iY02h1CigDFq0KC
gNuBZZ/pZ5gkpPICt3NxwSbOxXeL/mVZ6C7kLOYpVIKJXqwD3SlEUkL9QqKgosjseoXnfxDss5KZ
JdbDHTnQqWsbyETaLNPTi/k9/UyvJIr4F/aJGr1zxAqk5VqpftJl37aAZsYwg0LlMcv8FF1eI+J6
EbA8hMI9Cmfa6bti5clSo1+J8KDHPUtM8oylBAVz0fOubpJEkVCpPRo8sfxqTAN7pt78wkFGY7PX
cy4/0T6ocPGIwkGDgw9XHHTUCdSowqPKq73Agirq2A5UR+0cLdG+PuEoxfaF2agQ6K3hSpFzvFaC
8/LawxPs8RkUbtS2CRp2DP1LzJQtpPWTGb2io8LKQ6tvToFI2eiUoePAtDNBikYgvn26QCjgaE7u
Bzvji/uYUKnHiUH9AhiAW4jAEey1dYdJqvzLT4PE1O5eXuuNdWL+p3X/yOql7aWdguzjM79Aj6No
99bkNPNwcqGRkmI4pSma8RshxR86nFisO0F0kkfHCCGDf42h8qW7B+xxVfNZ401zriv1IywdVz5r
pQFRF1S3/9vDs9/taKUy47P14wZon9tdLzRN4qOUMQ/1AsPbwzRMZ8YdwgVs+0MroMhmrsRfvBeF
QllAWpXeb0csJCdvb2nL6y1nGavcjqQ0Q+Q8Dw8tSd8Wx03qDyjspw3PttQmLvwpweVujMTnxi/P
iH7ploQ1gZU4wfo+CHWp1IRXTSjPxmFDhCi4dMvhwpGbVAdGkam1AlVhAmBDOgrYuLdUm8dMkHeC
VgYZS3irJ0ZdxcStPg4j5Tq/gZWdwYM0Bul7UsDff82Nv5Hs4gXnWfrNaIvX6L4diDotNHEIZq46
y3OPYeAendtJNkcBRCiuWabGv1NQOXkq97RzF+2M4Fa+w07R5JNRU9qn8nYFXy+O1XxfrxGq6Qaj
rfTwOZ/faLNg1+ifHmx+BmcRHinKtiofzZ23x1bBr0uCZssJ5Zdg5rm3xE09dzX3OmWWyI1ABbHD
6/xRNcA8F84Dxc65WUQM7mNiNVP8eIh7Ey6yZN4eMNLXxXwBGhwFuUdQSF8YVB07h/Zpt3WUB/e/
bAZRmnYKx9QoIBmB5afyfFUk+Hd5Io7aA2EJbdjm3kjcTPhu6iiZJhQUmNywLNYGncJ7GjTu69BP
HJ7bnxIC44BSQgc7/7lFL1w9SU3omLEu93v6einYEv4V0fMrAM83L2tBRKLYPa2h3W/yxY4whH7m
pHl1cOlyudQytKMTayp7VU8A6ldO6TpR8R2J8rabRG9YjYwnOCmOKs4eBrN5vwA4M75yuoAnfmQ8
FVUSpQ0Nme1FSvilGM64duH6gk9gmemkMMuQWbS65SAPxhKyMKM9rORr0hPwdSZGLgJCZegvt6XF
LG3xlsmlZ/Dtx73zmL+hc7LeEAthRDmD0s6dY8HGCYGcxCqpDhVKK5yl/cZgzqIy4gmryvoXWGSj
c+n6cyTYrTb2Fskb1yN+96aT3hjzwGrA/c3w6aJ8uV/Uk8yhiJS5ng0dpDESPMsRjAeadBbqFmeC
WVhwre757Ew6DnC5ljMdgAJKa+rAhJkr8leRZ3ai2wMa34hWYrlYZ7w1lyy0dojri1HAvUcBPJo/
CfbReeHVJmonRJhfMF7zhjyrk/i2j1cAg486QQ4BvmQGu4VoS9As/rd1+TObS83Ji759aq0sCtVv
rEBGS7F22IjImlxwMADGEDlKs9LoSEJzpLkehNuHQZqgTOPSpeM0P2x9p1DkBzdCdKeo50GGCwz7
6t1xsIuUMTfQlobOsVdhw+Q9++jZkLBMHMp3dKWEmZ9VxTYtxhN45Ol422TMdIZQpD3DKCrpYeNp
56ZbqZ57Og+bdQCuDc7ktFOVXpSlPynO/kGy1u0lk2Lz2MKb5wIh3p5Hf3eeeSNIp+nTOiRRIWFH
ELn1T1CSCfExiT5UWGCRiLA1Wwm055Zrk305BfUYbyBazS5rTh3rcvLVU6Ryn/wDW0X1yBbFmGlX
xt6k6lZDDYT3GVud1t+fEIZHlklgHah+mi/yJL9C7uC4HZ30p34DimLnL0bPvWVkfFiCxRjZeD0a
kP7YnO+sZYz1vr5F024v5wUMTtRlVuvWJYpwJnB1TEEZN+j5p8SytTIh6S731MN73T0guBDlZKxx
DLM56uLbh4w9fVh8icKuOfOH3nNkowJZmcaM12s1jo3ybFqEHt929o8TS0k069CLsX2YPaVH+Zq2
8gJaNOErYQeUbopJglOk96h8dosHMW/O9qnbNo2TTpGFz+6ieKC/r+sqKKXkDP/b/xmB4WDZfe2b
KU8UfJPWJ2hf69iwWa4brzV3mHjnPxqq8LufOikZJ/zXm8fh55DtweL0mib4LGcDH7xJSUIOwQnb
Y3VaicLIl/EuA9WjeRXoC7oltz88xxv/1Rc2dQB4MX+9f/QqMtctLrB0pZlvc9QA73NjTo4ob9Mo
8AyNCBpmIsZS90+d8lsrJ10Srgzo/O/6a1LUrWge7GQC8ul20zPHgd7Rey/JQ38ofApe/pjmam2J
7dS+KcRrmO0Jpz/3ShVSit+ueyofvFwWbEqqDJeSL+AU9HzSm5N20BSz8OlkUYkueCHo9f3msppL
9op7Ej4EQrJC3nEPKs2I/qcKkG/iockRRAKc+kT+fetOZfo4Zw8k9wdj1fMAYunBY149U1CaZ2Ss
/W+sZyt/UDAwKAOW6jLV6ODYt0C+u0MVVvmklSrBk1mwX8CWS+0JrdYFdLnFO//XvQBC77o/JX5P
a8xGhrbcgFOpsYvhkbtD/ksMyGX+uwKinUn7Ohp7+3uqQcqaQmYH9Ikd9K+qDYZOFixSWf0Z/Pw4
zvX6pMpYMb4/WvIX7IwKGRKSw/VbCDzStKV8Hcq35iWtPuaOaTYBEk9w/FP4rimHKs4vZ1+ouPFo
GYrHUaYqHHzEovg7ZBwkIkbtveXQ2bB/Mao6CGOCbMaWCdenIWxYxt1KNlqFC2qpWCpgeyUn4MhM
DNJBTI9vM2rIpReBVp0kpSvc4F6lFD1k9LNOSnKo4kqnp8E6AlnT1DmSMxOumU2EDeAKfUQsnQq0
JT3iqv4UQFJzSGpArzY1dQnJWRHtNW9+nQePK7OqUbrrZCO+H0M6H+VIf9iv3ipVQaSshe6O5VjC
pW7IlFfHozKvJ/hfglGh95sPolAXRb4/o5MZcmAamoVFrBVJzO2ZN3AY7rdB87+nYSPX5dZ0Eu2X
Si/AHbxovexrz9T3hXXI28HArYerziVV7XDjN9aTJPNvD4wlfmMKqDxYfjhgieNTI0XlCjlXcknn
jqiPRb0SoIiUvfCPs7YJYJIBhTwe0388hgHQPDuBYEfozzcN9O0Jbf/xxryuhW38E6k44Lb1D1lx
2pZKQYMjJAduuaor0+bXRkUbynllb9lB+lGHD1Q5FPMvN3ZIJ0pmVQ0q4HF8Ihx2V6nz+WhiB4h5
2gWvQtonRGC1Jqbjj9r4U0+zg6u3VuFQNvHCrHxwsmoPdj4wfNU3OebwcV5x1quTpx+ZTRBYYLej
YywJmDcvjq6xRiK9AKs650C7+PWooojUOtuQI12idWcRngnjEnDYaNf1BqVn3CdYogZo/FWo+UzF
m8bEbscbMgTRz7f04SRMQYvFb851dUaWN+s98cILLSROtVrd295qi5NcfaDZkmM+qky7ZoCOawvk
slwGeXB6aKRptO8qbjVQ51vl+qkwcIYS8kEAvwPYfVg5Sf4APoNQB0uXknF2LQxTUJlvmVDpE/IC
wFoIc69RWMM3k4T5Dh6sjNhTGvV1cTNtIByh6ESHD/toPcwypG1dBzyAl7D0OJ3iLPWKgAxYF8Hp
2A+rWtWztQ2nGcbHpfMD1e5MihcPHIvl4V/pn0sdZl7+YIbuX4nuWHj0FkWn8K/FlIx/e2t9tpVd
mvQr8T6ZMe5vzuPQFhwkrAHQN9VSnoDpXPj9OSGCy5r6ysu/OoofKNgKjiaWDCVTRYkkYNlM7fiO
J7Ebrjas8SkR7BaE76Xh8Z9Dj/Fprbkl4vj6KYO1Wy/H55+DI3ZzgLdn9UBa9DlxrkrCMBNnLZHx
TlsfWLtuhuFfKvbCDJHkxZhlfOESqMplIJH2cTs13KYCTi/gW0q98W6YiY96OKnf6+rpuaW2bLST
iXBk3+bVhlEyBa6zuXXWHos2MmLD4QZw4t/ThQjclDNiV8cHjzc21LSmdw3qX+ntHEaqEeOXd/WF
E2BEGaPYYIOkeDgGlopMAPNXmts+N1QsxKrwyac9SnoJSWBJFXVAHO9t8lN3Rze8nlXmBSgw8T/7
8U5SlgqdHIrjVZL38/C39EKwJLgjB3rY6dbWqLWzkMGBgFDY9BF5A0W33q6YgB5oOQPbXO4iSst6
EeyHqFOm5wkIZM8YRc+GspMeuWkwmDLLOmXZX8yKe3YQFU4tM5nFxZlabxVQc3KtgQ0iPS28YVJZ
NSl8aBXIOS3MW63c7vfrZcI5z7X+6dgatHvOyzOzjae6jnNBj6vPsJrvpHdC1A4SOFJYjh4N716l
OYN3L3FYadJpAWvj9oCpzsTRZZfNEK2P4/1eI/nQ+glXMgJZ4KMKSQwMizvpJaYWjI1WiA0Wovbg
ycbGGoOmtVkIIS5BH1+czbZq/xXxsKd5U4UCpg6FoOjBGeMNmJ+oag+Pu4s3vamZ4Jpx6ogk4YaF
gOam+nIVOKpumTsDZBIiVf2tXAuA9XIfRvG5kPfeUejj4RlwvuWoaiksajHv/o9DFAiDW+mN6Rhi
4110Bj3Peq81crAlKZS/dPmK/NgWhA6kbtPfGq0ZCiYkKTKEbHOv0+MfRSP5KlV/y2llbzkt6sgW
X1pt/jmPnqdEMaoq+m8xmyqOJgW++9ABghoQnPhfeuCrEhguw3AIXvsqLctFdlwPuR6bkJI/tcbi
0TFUFTCkbd3Gf3aH/b4O9KfegdDnieKyulSdudEEnsxD+o14T8NOzgtUjrYl32T5FR8f2D0w2Dme
wIA1MzI1P1SIujYxwZ3eepscZTx7a9eNufLyLSCo31ZbTCrg6S6bHIPLbrY95VFVd3B+DNCAATqB
1/uCuGPjICtu+ujs/xeadk4AfjYETkD2EFA2VPQpa9JA7OoQ/9Bms+n1lPc3bozozA57gfgfI/IK
YB7usaqLIzxR8SUGNulZn2diP9As9sqjKXw66pJOG2sFANK/D7yaixeKNTMaTQtNbYaozH/q7rHx
htLldN3cHjKr4KGjNebW997nMfNnsfwAkmnyct2jUTcxfdNuiiWzUBuoDK4GAU2PKduqhBS5+IY7
rKlkEfPkltnlkekyvxA2ECRAba7/bszwXinG92m2FtnLoSqAIvTwaXhwvDtVHx57Sf4Myxb60C07
KfKCAlUz4xujzDXNdaAoUofJNWcaOv/m3M0u/rmNt3pmB4Uv4ENvIEFQ76SSgPxFwfNoNMBpvOqw
KJql/jm/ypYIEbz8PCPP6ZZ4mWijLli0bbX33qbFGiRyRlSU/Cxn+owEo2zxNx2mxzT5BlXo+uFL
xZ4Ptyfjt1zhwf7+wwuM/Gzs4AZXEYlKc5bm0ifQsyMF8BhKWzhjE933OWzyl78cc6DkDftBJLsa
F7IFVFy8OfguwAachMUDiZwzCgxopRyw7Vn2toWtpEPxNB09E9/Ek40mp7BUCqSfLdD7hSkV1sc4
vZA/e2r7T1Ur1jpmzflyBETlozRo/u9bnZe6TcSGvzuXdhqfJTubc+PCRti9ddwlbMpKoxdUPDra
qyt6yEUFk8HDm7ba1NJasARDJXHuMzOpamMVAkAHi1ySgzkUK801iyfEkNGNcon3hZUMiKUKu5fv
EJ03wneOCAjs934//DAGihF9hVCZ6lMnvw78T2Ao/oWKvGC6u/GWXAvvnh1TZ2vWWkx82iiH5cK8
9lLf2tUySCr9/J1TrlaxC+cVtsd6/jXEdvpmOh0I0okAQFBd4QUNjhnsmi3JLF1FWjTSYFifo49t
QozS2zcCgNdXYZTQZ1nhGJwJOMRCActgTTNHaGEVHE7qxJReE2wWvP0rlTuAMp89nPm8Qn0vL7gX
ZeYTNS6U+zyNUoc+2xOQoNV47X+IrjZ824D28PkuKN6H/WwGdnlQ5CwRX5mfJ81SJTxD7x3PPWXe
h5vjoas53gzKdeE58Cl2kSVqFF0y3Wt3m9Ab2eJ0LMVPVzBIeQ/pDoy5RR/YMzlSJ/sAe+l0YcNq
39vWbD9GrN89Tl/1LiABEcJW/ktLPaDDl/XQFc0F69U+DLR4vtPb7CoxhNtgPK7aHRroZTTHfaFd
jcowLl8tRQNrUhRQsSt48PUsBC6euEXDmvvwuMR+4zwDNV0/gVjCXUuAyg4Qp+lr1au2vKeEFeOH
ORJqS4Ix2J7sxn0hzAVN+gH/0FUxdy80jh2mAjlNCCiySnX59QO2VVILNIMaM0ISAF9kK6s18Vsv
PcsYi9D/CgbjcRtjfcXYlGcLSNtVY4+y2qWEjo4baIqZmnVK57EsTU/UJnpW/npd2q2hF1hGcOE4
qu/GFC7351MxQyB+WZ8N/Y0c8ENFDhY7+J5mKpKNZ9XmVOOY9UrnODFSEkmBWGSa2PLXcGL/czWt
RZawK/FpcGNYdyDYqKXdzS74x0JGPAeKeF84UGwxuclf3DtaWtThbS/yPeXVUZvWZ5GVm242SuQP
E+9KSS+7mv4sxoaaDIPeEYcQUFRcLnkUHlRLHx4aMml7RIASdUto7+914RIU5a5/XsTAjLSvoeyZ
mjwEiQZhhGFNH99BdJiu3LySAexs3PlA7qFdpwKd4TLNV7IhwMGRITxn6pQY98O2zFq/THYXNjF9
uS4ME5C/yBWcxnUaTVJ6FPZH47/HFh/pDwa25+mH6h57IpJQbfFw6ZDK/HgJaV0yc5eUFcd5/R0l
mkzmOqphyh9U0+wymF056rGWbZSde7KrJLWzcnmGAx1X3xFSbjgXVLi3eoiMy8SAtcT+ja3c5lxg
BXijlSsLVgaLJwYTpDaFN8NcrdpbcQVlPrkOINtls4fLSlSn82APhSAbo0hKD99RRYVGnE28Ezz1
OwTAB33/Pz38hax7txiq2OomiJEIBOipMDFqEw/3amhT9fHb1dXo5//q8iH6JP5DHoTZXw5YvjBN
9ooObti0OHz1hDOw1lqTsV0NlCzG9px2ufIvqnnltu/BKm9H/RpmRMLD4CgspAHYf1/a/ecFwhOB
FHIL8UC4vM9NDDEzATCL68nNqcTB+aCNbTXtZJgsCnN1FqAPNXUNdmSL1hhYLx2+Nhq7rbMn9NfS
KmbWtcJbWSRLeM9EM28N5Jt1LJj6o2oPRi0ZRrptyIG3Vrl50XPmKFcEGlzcKsDGnj64J2X/vBCb
bglginQj9tlaTaulY6celieH7mp4FI+KSjUHxU+b4E2MpmodLG0cWwLpAQ2wYSbAxN6pUnrlTWXm
ZlHHYrKmo2PZDIbOCEcw20c7NFKEq5xzBKBmoaesg+p/f3JjtereDU6hzeJb7ACvgIefQltnpQIB
f1oojOlTZPqaL1NVnTb1cqFP5N5BBMJH1Bj9wzotuLFqzG0Np5aX5luMmEyRujKqi0uqLq4DVv5m
axwpV/weEwMJrFqwWeStUV+JwqS5oSMkC/cPjS9wL27dcH+f6yLbErnqqJS2W3+xIzetdM6BReLU
SrDpRzOdreMsbRHqLbmVL3zvHQGracXPI7vNloalLfgUrdZUNFSa+1yB2Vjv7BWGjpyJzkoMMZ9k
T31sEwgVOxRgJHhRBntkoz1IqA9U2bbRDTAxI0EbrYaFA2Uv6kxQNsnUFYvSWVlt5gj6fK5IXlUo
T5uAvebUBiPdzrNNJn/weI3K42VxpTwWb5BA3ur2mWapwHKnX9m6ep7F3x6ZCmvI0r28jh3M3zYw
WL6wOdlqL90BAPb1Si1wsPGJra6v69VaucLIhCc3pPzZt8oaBvVE4h3Yd8s1UUjmsrsIEvW0hOil
JtIHjPNQTNWyvsdXdjpF9ekWCSce4WJOrcyFYgA5RvddlBcPIuLewKGyjRjerHX6blUSmFIpRTKD
GRpSEmfWvlqv0/jo4PW23+dVdGLl0m/AKobz3VPibH2Ji8ynnav/17Rkuo8Cqgd88CoC2dTnpJA3
EmzEm2qyG/ypyYsY0wdKuFdJljvzCQzYt8DjhfAuZ/epBYbhx7R8kijITry+oERhSGqeYpG+AdQb
dTvDY1o3AVeQbi2qUdnC0SHxZdt+cXJ0Jj8Ob75ffhCZdGC++8yaJdbgkiENoK7Tv45VmHd13eSA
Xg0qKki4/rDrtoy+ppb8tOQaqjTB7iqHAXcGah2LHLvyEwmFhqC7Ih11umAbLTkCvRYKrEo1CjkW
Wke2M7GZZkYqmp+vqEpVG0Kc1C4UXacx0fSYA2VXu50duyEML7rZ2gpV1KG5tgENXIUZeiY5DXSI
+gQqm8jZA5Hv4GRHvkrMAMsjhT+0PpWu3zxEfY6Zt4BqbfrDOoOqZK/8Tx8OI87Lv53PuoLo2E/e
rK8X0F2XVYGnB6ZECnQWggQ0UwnT4cnpNnbZ8f0+ynQizluo3X6N3BNAVCReAKwGiMqa2Y4/9FK5
hrz+nZfKvJBCqnfrduKtD8/1qLzWuHhRG8oTgOxgQFdUufy9NFm1lT69IAmKsfMXs2h+HX7hqMU/
GAqPD2wjgQnKvw/JuTKVQ3GguqDZ531MFW5k/8I8u8OswpVnmPP+ftKc7lPbw1pkfLtN0h4nm5fd
TwX3aSFSax0XW0Tkz9NKBcDwrkpxT3QruPlJDl5BYRutvxfAn/q/iY/9uARu4thDR81Tf7MWy6sl
Qi5Esu6YRC0Vb6IHApdIR4M7Gz/HodLdN/7ssb3bC/yfR3G1X7vekySUguPYkS1EQP3NDq8L3qDz
ORPOYWBjx3I8arK/4F59aLoAf+6JGQP9h2HS5CbvmbgMpjhN0RFI/jA5cFRGxKiwOt2CV4urx6Jx
+JZlbFn1qLM2wdR/MAuGYYvT6l1Cb1xIERfJFxFNWr13nlmv18b1tMKrFSQGewPOZSf9Fgozlnay
ncD6s/kBJJOxafZN1VMix9D1UyrXPxxFpdGeFioZsveyklGvYkeJyAyhyekvbpP2OGREte3c27HR
aekiseRfDXrzBc0Hia+8/6Rj8NLL/Y1U27FquVla90HbZa7VTHPrbjkPOejXGWao8woGQg0iHWsR
ku4B+YaKnmQA8ElKSjZO0PZFvPdQDEcTWx8Ig53pfVK4mn0v0S54c+TlMYU6KmNrfIA2dpcruyyM
dMJshetOSiqYpgb1w/o6yeytxazHdC54qvkHI8j4ASWt/zOxbnAujCFQ2MeqFhPXtdc3s1CMczFU
jPwSq04jz3BcZr2vAdjcNCXutVxLlaAqPaf4UN1VwfgkHHN+YbTlmUn03+zDR+vh8OexUcxaveHE
zma6ARwl2e22dEEX2m1V4s9T9TKjQMV24Gt5879k4zO4b6cyndzt3LTlGtVJhlZopfnrG4N6hf3t
NvCaacbRea01EOTW38qebQMClNzezuKQ2hb3T/ynCkhTk8vyQA4fYrTcf0BDWgZUiBp6MvBv2AeD
WnPhQCNMIw7r0+sXpmX7CzUeIJNbqT5YuiA7YiHB2lTFIoR/YlzdK59O8mMRE9Dy6j1o/zX8kxko
PqpnHhOeVymYRono5nBvi4erl3Ai6O1Z0UdwRSw2FPrqcKTf9lfTzRu2SXyxqa9d09VhtT0rFF8q
jimS4j6OZfU+nk1Dj1kSgdvPWR55OOIjmQZuQkSfEAPLaFE+gyEQOFjB3IQtJ9d8GqLItbgXX0dW
TDOcnINSeFdSFWFLYWlw8PA7zN4gqj+pe9Akyjralv9m7kPWxd3Oy+rhQ6sE6Fy4Rc5OXU0Tkwyr
RVDySq+63A3pks/3e7H3yV+KwBEHsQlv5kj1ppdWx9jSps1rnFU7dAqTeLRK6ZM0SuRLd7/X1lp3
ztcyYuVuE/IiOBMiWI/JZ7GOkOnOc8bEOQQT4tdbDBqjlSv20l/mmMIC7VCw3udT1sZEnKQxNDZ2
jm52yh9DCTK0BhrTmyuh4v0Yq/cz/2aYGhxmTMz04nhFrBeIPg2wxS5DuXvNnwLwDyg3iupZbRB7
b1h/uccw6kUf7I0HUaGftWF2IgetcGZunnhZylLFhE1wBZcqwumJD/6mm6iJjdDNV6YHwm12AvRL
S+cD5K3j6siYAwt3wHDF3PNymrN2lpNgc4lnuwYH0kufQKDbRtW4bxQCqo0QTHUNZiRhphHmG3p2
ETVQsmG1Dq7p24VpeesCcgfwLblXyXNach/dFQKAB8OmlTifuo+wGvuBt+CqVTLvV+3JUeI8HXlC
3A/dlR3HkAPVcEJ1JE9Yqxg0xXD+vNRFhV7VpM8TLzrJtbzw0hTQ55rxmJwexhD4yyvS/BJQaAab
vLm7h/U6VBQOXQcJbyWMf6+q4HsyFjo/ovOa3ZqUqUPRowUhxS+MM/xp/ZRLF73vk2ggpjgXf0iE
GgxNAtz7lfkTrPOC5piclfVSmae8uVl933xlkklO3wRcdxGREd4O4nXjgU88Acn+6I8fNvveRrtk
APoCyVQrzuookpT7IeP/a5xImC1SI7DJx/9Wq2Xi6Cwm3MsWfVaVdko86ezLTQ2L1glTW9D6OWfW
hfnQuF+LEIEhpbwlGJTimmiN1J9ej+z5GRVQ1Zs49s5o8SZ+iIaqkS71wg8+UZ86YN9ubwPk1rbN
wiK08uYTauBUvvNZ1zivdole8PRH8JMsbiKITGOOBfvAGoI+TBN5CDVAo/rZKwmU10cbF3Ysa/DT
qPZPPFgUt+xE9y3GjpmAL8fKiAI5rHqM6Ep75oT1EMIi1GV27DT90MR/2qXZMhrWF6AVA6nmbMg8
cKJEUFWvhqyPQ8icKQv85BJWVDAlvn5LlqvnkhYo4ya9grce09mOsCSzBKNXkLNephhVqBidG3BI
yPN4vvr1Dw3ZN9+0tLkJ2QU9WGF7a9DnRodD6LDUblqOuWMPFRDHEag2Sb0ktriXXnZ/aI18+1DK
WVRXwvgBsZeGyOYTddw+CFV+fxM8T2PQTgN8QZAX0ot1/AgOmbVRlKVDpQN+pJy5qi0JC8mzNZvQ
euWPavl320HS3fiUTYuuxBxwShATDotg0vLcYGFPZ9jyuBxegMkLiFkWGGSpep0uu/wRe1ZTA7Do
6nVgs3VrtYe7/bBRKI46gS1atgS7+HndTbG8p8pq6GOwnOX2CxSpCTCwxxL3eNwPEgNPrcW6zCCp
ANV+nvNEdy4tY6te7v3qYS5DDr8YJ5rT6DnXAVRXtUFmCoJ2Ar+XrCiEoQ5C76AYNogOuHxZZg6y
t3nSeQdbvmHKTsP/gRmlhXU+h1+nCApiH8KqtdhPliswCLubwgJx2hdtnEOJQZaHUHNU0ANGT/LA
CMx5n9PxZLTDQBAvg1jW3Mo7YcOEaS/ZtKHqj+JDpj06T5FaAruKBZpvVCG81X50ncmaCTBe0Bgu
ta2PGjDdBlz5ADGsGKY72nK+UzfhmFzyZejP1HtCobQb0wb/7V5MSoctwJ6EWzb0uIAxjT8Ic6Ld
5pGOqeJ/Mxp7j5dLg2zYBHifAST1nNSMkdG3kUsLFgfaikELaCWzigOp6RKDN9qBbPlSlNQW3IB+
fmJDVAWmgLdG9ppFF917RQN4vKAQicr/bmkiOubqJVNKVNvqN20Le7+C/Cn2DHTW14+M6noeM5p2
/z3GH8NvRN7biFbeK6Z6x2gYzuc5iUvaD//MS8IkhAvYjxvPxOm6P+NNRKef0GIgdGHPoCzGc2gM
ZWGDlCw5ArL6dnZwc8A0f9JZ7FoutoJL/WgBWpxUmdO+Mz8FUcS3ojErj7kokI+iSrvLjQeto7FL
jbCspngxl2mAkDtvu4lqE+orxPp6D4lGZcd0TRKt8xb7q5WR25FER0uBUIOnEnd1/n/gJKURYoBb
hO9NX6nM6ynVEft5LaXYHioQbquhky4iDz856xgbP3Zu9WqykR1KANef3nqjasrF6ZF9Frqeyjc0
uctjCXn7MJt2Hn6+9gStPKF0h+6BC1JGlvV1oLMG3ozQs9LgkuRNyRZuMkdbtm6BeeA2fxJzkyDy
KSEVekTHaXF3SLHh7AI7pPo5niGxmKIOdzdBUq+DMb5GO/hyG1iKr1JLXDsFlxpUqT/sb38hssry
n8F9e5eJB6pEqZdFPWU2e3oDHQJ5UbiYS13cPZGeLaPkxGbeW+Gbl4TXUarX5n9Z6/QqjkoPT3/n
QeFHv+qOopDfJBkf0KKatnG0/uIsKuDryzb2EvzWu+vP8rKSpKMIcCJj7XxbrJXueLt29uhcdqP6
gc/Pwhoc6/zP8Bc0dCgJXEZ+JDlTTKNOPTkYKgPhU6wZo4cEOVBPqOEuIoHpquhBY4Nlqq2htVEA
il13EermOcUM+PCbqeoT0qTvUlrB9a13sHsT4zGk8Y6KT8F87qtdyYMZuD1fJbluHGl44Yf8jXTP
rAwHhJPiZ25aq9SJhMacBEOSlDs1vN7hQQ2yOuVA/ddOv8znTf6PYXgCqEy2mm32g7EX+yJTS1lX
/zAsfLbvFq7gZw24A/mXclvrxvrPahD9h/QX4Sikz0HcGZL4VqUiRt899i6QVLM3v1B9zWqmrZkk
65J6Or72EhS/jBdYgwvDSI+h1NYzoIhZBZXkO8NSUpZPIy5D9y21r807664yjZVQf9fYO2aZ7oPO
xCEjyekwizkj4G7LR4CjLvnSjC6rY9xILwDp82oMwsJ8g/hzOaWhHTFySXQZy1KZtnOqCJ/FM6F+
dzeElOaFYLXtZN7ooyKJZ7nUYG/xGq0TdrSSmNkEZApAIBwHfz1LJBvUomiO8fhOUb9U1cld9KsY
PORKlcsqKRw+aQm1DnI7w2ZJWXOqNOcN7VODN9t/yJAQcsUCocDyQ1XPT+vBpsqIE3Nbw5FU5FTz
sqjTsPy7MGMyLL6hiwwMn1a8il/Sh3YhDV/qBoAZ/R9Y9BShVrHZH6PLs5eFjoR4VFmLdyXvHIt6
rKjfg0BPJzbXlrJaUlHgDZZ1+m3dJMpZkRLiJpVKtHTn9Oh8nKIK/eNPMoSQRdlS+q+6saI5owB/
LB3zRxaP76KzUqi495rMvczZ9j7hDRuWn0pcchZsvQFRAWvjTCiYshj46i4B9en8zU/SyXN/sjBV
hitFbfLKuPeVi6v6j2wn6h3RagvdmPqM4teM3fhhCOGqrYfYs86P+6kW7KYathcIv1RcB9D7monm
d3TfEASfPMiDC59StMODRylFB0aBcY0qLzF0/sXOHhp/h7qNjpHzl0jGBHf1qWfdcy7qBPwVUCLZ
jmKs8zKgSo/g7HR6PXa5jVTFCnTNW1EgSm+K7hPYmICj5VyQdSy8SAUH0NCik7kKK6HCyGWgQv0z
2I3nprTNRfl3Z0Tdwxqg7dFYHJAATnWFH8Vlsbs8K8+oMaB9xcgBaq8J/Hcjxxs7zrqEl1w3seXF
uRRNkFB2al8k/QX+0guSPUv3d2cMBNu+R2HEUXPNvRyb+u5H89L86YPcolLsQT/Ep8aINCYcXqWF
W/WH4O7BhqvnFX9Lsm3z/uq6g2NtzH94DhyjYcBAZHAZfeqnCPdfBN4y4EAtgLRI0ZIp19hGOiK2
IY3i+86xPfFOFAvff7ed9cMEU7He6DcNz+UMLiY7F6tct5AILLDUE1A+uNvfCIM436ZoEDDHO8nb
Q9JUeU0j3FS9b5tvaKeqBOvxY6PG7gGBmeP9dwAfkgsBPbwwbGHpSVfEyjssoirj2LF90uuqRDTK
1TOBaeOWflSxCeUUWjuPJElrCeqAgUgKECotF/pyxH+tQdbMmTL+kHhDpGu16eqCceznmk01PH8l
T5/n5IBYpU1je2hDGLNxfs5/3WDNmb8sAbrX/BT2ecYP+7tKM6xkU6R7xKZWHLCu78OyeBDReEZ5
OOpLUDpXtB1BBTBTOj9Qgi/DaUMgQFEbY4qenEskMMRdrkPBR3Akp4lkczClu7s1etNLlJOL93wG
8UqmaFO/xF7frbW2yuRYqfApg9Alq2g3UfWv8cCkrR2OaRmNVcy1/HnsS8MukhFYasnVK8VgbZ5s
R5oYDSYwMVDKGoFU5U/9bUHPAFw7Oto3E0C0olSucbv4JaMSgV7G2OqneIMiW7U9b9ZDVny/6x8U
UKDCbCOFXao4QJMtha3tNGdSVP1ejYq5/FgsjXP42inNxWmJw9smsiWhE6EBaMmgxTDzL4TBwxIf
hHY98UoMJTazrCdbptNhqA2qKhnrN10cCU9djvmzIgoy02ZuXQv6PXKV+1CFkdCvWtAJ8AMZ1M65
XjeWTjPZ5CZ3TojrW2eivAbe4Ak2kpZUiQEabiAbEKFDAMJJz3Ci+HIEitRIi9rc2JZ7js0T1DUI
nOlqekzPs08GoLiuUwLYyFqGvc36rZiMOoAWrkmweS6dvND9vH2qFcS+KXsYQV/IMAHtHgG7g5S9
WefJImtHP8zEzSx4KAXf19JWymDjkDnwOhJpZi505EKMkTkO3HPzu0161rkBHMKLMfPBSug4LFq2
rktcWouDRCbNqQBtFL1o77MjWuB37cGO6BWGI7DjDyFR/ySxYx+Easu5JkPx1ldWc59bK/V+rdB0
pUk7Xu8SrrQYAzFcsJ0TqFvI+zl7GjB4uY14fnHoJx8/Q8ukneTblJeuIMvi+aH8OY4MAL9nRSfa
Pyx1klmVb9uICl8HkLOFPQOulPKke8PfD8USv6tYMLYewN4orPTTmWSriWlkptL3zjLhZ9LBiN+l
xiamdsgkDBIJZERl/6GpPwMKlLnYBhqBkQ7rel6d4AZUjN5PLHeNFqnNgARvUXOGQ4bTYtwW+aez
Fi7cePfyY7BjcPPscNFI+NZvXNrgArPHE9K2oE7gr/uHHI7xmvCuzqtbaZedIrIDBRBuGJQh5is/
EdD4p0fT4p1Caq2vGoAOtH3GKx4Zgqy+QFLC2KCZTvXAX8mg/vKUkPS4kuG7preo/eh6Z/GO+k7s
WUccUa7/SrvjAVzwBt349/On6Ek80EwHX/7t/uWTmcx7gETxhCufLSaqV4Fto9xk9GkCuNXDEp5w
LcjLG22snC5GyEjJ3lWxB+HuqxRj6S3UcvoL2dVQTjwbu2TliKLhLCs+Rpnre8HdXbamDcn3Vg2J
qisoygRJ1h8dUfL+TCCS8b3fFHKI/4sPu77tT2R+hktyRsndVGMD6oV+g4isXZYnFrGKgKGgoPyf
c5OaShiY5AbSsIexr4B9Yb2pSpPkJCMJO2WlIZxtVYznAL1007oLuDeOEWOWOR90vlCQHsEFkB30
XPcD9ZeDd3ECJgUMCHEF0AeFMX/vcjk74HR5bvur2PT4ht1g6nxCcRunfsEBCxUL92CvYQoIHreA
Z9lmCatwtzmMY5E1lWq1dasVDFKJksT4m3P34ssP1SCg/KRZow671pKPCghmRebxzVyhwl2rQUYv
HtImUKXNxtC+8+Kg1cZjo7I2AWqNawTeHYtOWR7RR8zB5kyY6xmQMx0C/jJutuGalUFDas65Hk+4
Q+lIBkPa0CGw2NPEqHtvdk1g7JM/oTBwduCTgEnYKxQGmAsH1lNQX34k1JC8t/WtQ6uFunYI87KD
2ev5bZYT66I7Sqxcrf+yav5+g6vyzZ2vUFVwLW7bViMcazaSeN++a3VlQv+jgp6030lDoJKPy28a
h6qS652RrlvcTGLL1/oP6zuMzEvqGOCVXZI0964nht9j4VxofihLKYyLsq8zekOVyLKzP9HXbMnR
e42Hx4033SBXRAN62nUqibrngEsTvQjpeRt049/Bi7trLludWVAfoMyaa/kLah3xC0G6pftBserj
aISU6xa3adz50AtoCZIF+kIE6oJ40xSQ7329BG0kEMDzADBYZ4xWiUk4YeoPvqebK8OdJ6JKQoz0
/0lKOkeGRHzi0V8kv4HLToYvh5ySL7J61iaP2ajipaJDS5RbPEwwK+6Aj0yo2l7h8lLYgmS6SEWj
AQCHfhDMGymcbb92l8uHt2DK/oPmwubGU19YAf7OPDWSrTAKplURZDCt52dE188QsFlJEpP9Ff+i
rb709MjL1ETsmRgWv2lZ/BOhrzzWEUfaKN3bMbFKL5hrP+Yy1cVEFMG6A9x6vp3ISU5GC1Pu14Dz
X7w+EqT3rmAxmQ4Vr/LItwebUTRu7GzW85lDuIo28XvjeoVV53SOls/JpcrB00nt+OGAolGuY4XS
bUJ5S1cvLwTbHKhz+/ZHHawqtRhJ3vNsaxiNCixXf5S5a7oTgoNC42UpGJIarUyftlws8udAcI5n
VJcZay7cKJbXAX5s8dfmAQ4eH+DBTvZVsjzrYym+Xhy4LLClZo5Ip/IweBG72tm84Ak2Ikaizrop
qiF/PlXYU6yj9yT7xx24CIraJOVK8ZRzZoyqF8Mrh+gfBQTdv6zetVh0W26IIM/GBlokYfRjMTGT
EvX8h8fpZW+HEm7kazdUxEU7c9vDU4ZpHHw1cQYfoAxpvLfnlen+ureYbfU2Ga6OnRKi0JmYEKvI
Ab/ghyrV83/M7HdIbGEdWOYW5e1p7mZmGKjPZ2MmCeYabKvUbnU1C77UWM8C++QyNi0FJdY4eVba
CSQwAAI3FEq1mxD6GPidxSvf309c0KskRo9mudjxD7RYVkr6dy6Y06+0oNSwNpkGawB3mIQCxcfi
7/ZjHsnfoF1o8a29NQ2fcakAsa03h58/qKGXS6tKgbaRv6w48ZIkLIHngzh8LvzHiCkRCehVT5PG
B7PLPDfgV4WcOTDcqStamlT0g+XH0o/dJz/Qi0jhcgX+uUWHmrF2r4dLc5/LFA8P3DX+1sb5nmWX
wkR319FNVik9M/smPZD2Z/rPJwfanjsEdyLbUILtpBqqLuW3J6YVMZJ0MOgDHY3tXAEq9sOEkd+H
V6QpQVXTvz9nZt1h72Y1jnELFtCR0mkEV2iXdKVwF4LP1LLxOz5LovJFblxyJPkxWqx7FLQKpbDA
f+G0Oo3q1ZamwrKxIpxKKpoYlPw5DV3bg6A9l6Y0zRcmUg18XlLRxA25T+nwS5h3Dn1pyHRqys2F
cG/fQEBmCijgNCQnWnnUYh8QOMVqAZltHxWZhvnROE2XDok32wVMSrTxkf4LCSXwPyWhtReioNCY
jY0AFKjBuLKvDJSadI1+DcvpqEbNfJ0CyBK+3/3jRo4JC1XgfsqY3ok+QV9VKZkUxgx0wosU4RfG
02R1/sQLMFBQcF3wTuPQJR3nlSTkSlW/98/VYa5tGu+MBHAqz7IwEJQ+/2VdVZh2/9eqW8+hoOUV
1BJcplB45c00gBGpiJdbsg4Ht/JET+vcY4zs1XWf7HprA2cN3zk1KICwQIHYFWt6kNiFVl3TSb6F
Q4vJ9v30humI5TNxO2t6tC0DV3HSp+HR+goHZfxoQ9SGD1ha5h+6gz0wSRxnz7L1eejSScPu0FGt
J+rqVYf9kx6d+CdqwEKNGBSqcQ1ClPi/Rxla8DzX7z3nhXe1g/teKhn1zyW+LxhnTa/Zdl0UgIpt
jTKka6Cg5np6SGxeOezt4pthFr6PSKIxPnZ811MxqJANtkeoDCrnrKvogFgzETh2alYlYkrlOfQZ
UHEoR+Nf3AuoQAsPLZOzHFJiK0HmcSIJ7bD+Nw15vy01ssk/Ul7XSPXtAxzumNemmaGVtcbcwMww
vPAIDOoWqbqvEYQkRKHOBgVmE5N4is8zsBLuHepcMNOnlSXZfCr3bgx3xmq2mQEh+n1PFY5fMQth
P2hXmc37bTArKccgmGDdPBmtyTMYkdPGNxz4pnzxTnmtHydJmdpSEoiCA0c4/XhDToBsJoZZenYM
64sfsVLgmtwKQj3A9msGd4QeH/bqjBvFNdAxbo8CpMq8NZGv6ujmU8I4r2LH6LGFWDnocG3l0Bge
ewfnW0kANgGke61SzrlsEgnzIi33+Sk588vaicc4yXPL0nvCAatOvkBWgzBwptz8sl2Lqj/sFATK
JpaVSokPBgGgI+jSDjWU3D7HtAxf5WsHyBzoREWuYKbUoeSkb9V95LNKPl5wgD6XJqe9n8G+1zBd
PbPMtezgttVYqh/yEpyUtZjVbHMY5zKduBD6wDAGPTkCncz8FYGMvhm6cStlsSIU85e6qeZIHE9W
FmWfyZ5qx0FZZOfRHPLMn5NZL42rh3yyab2aohMW12438SiW3uUgKinOiYteWaX4LGYzG5tXw/QW
6gQHn+sv2rPNdKNYcxgiAvY3Y2eUBjSwtro64j0BHWinoMQ46sLTqOg5klD7Bo/l7I20jUc2Mrux
7gmAKo3RphXox0U01gF8g6Nu3johB/k9i6xx7r8SNjqAKst3540dr/03yZ1MNxXpX2i9mzwj2kpu
yMMCb6/skvb15nRDYTKLv8P4LUERS6Yn1yZcwWFggnB1yYX8G+O+xP2wNlj84q2K2nccVWf1cKz1
CCIBub1AWX5LQ5jIEu0vXTjzTVR+TSpzQDvfJMKuHmJRxUE/tpspBFsZVLvHpP0GgIY6sDhp7iSs
/2p1gSo2RfuJmLjmYGNiaMvxLR9E0BJliwBSEJgCo2/tkIzab8gK2H5WF9WFTQ1gSoQaIACA+mKA
C0Y50iSvQBVkDmRo0um+HpWsFf6Crol4SJWA4fUOM3zS9b4Uq62NfUycA7PYEnyhmCw+gKmGy/EO
iRbiAU5esbnXmAN1CwJZSbkiGYMK1eM8s7fMGjffDWSU8si8JHBNnngo01FZDiziQaWapIni7k/8
FH/FiZjCcRdRYJK9mKKP2P2k1D44AK0pjXHAkwIuA73h06QntlHAA60aBVli03E0PXp9pwDqDlUD
n6rmLnfBKguvaWtxtPfOyBaj2jHeL7qAohD+mBPCa2xnl+weGyXHiY/ZtN6w8Lrnsmpfp87llcQV
b8xMni6uFUmoVyU5k7QjwXrVa5DZ4mog3/auhthzy3w4IFbjv+1xZFIat0qa+a/pKUq3QW5njiBK
1yaC5pMBgWh/AoB1qcJ2138eU0ZmFgjLKK9TZh1Hjj6p8ITG8P3QIlqQ4Pj5SzXt/4Tba64GFMAz
pxlzkZZHg4KKy0L45YZ9H8XhMQ2e+qX2WZPZ3od9mYtduIReCjc5EYReeoQNgFinVK6bmugWhI+o
ZeRy4DAQuTy3JiEnHZUFvEfQq9MHzTiiOv6KssoESDmPkdc5QTB2vRrqYMCTAeGZCczEVtJzfKee
q8lZHypRmURpdMCI80K1GHNlil/iS1J32MaN8ab2w27t2hRWGu5rn4Wu8ewbdQqxgOdMcqt4VMZQ
IFrL/ofEgLB03rqULOJ5qrP/JYCnJG9LAaZsLlwOycz6qsK8URn14dQyExC4p/fvZTUYZP1pc2Mr
TPZ7f7dYpzoet2Sqq7DmH1mNM7o7wdvdMo582kAic2P6HhkRTiYJ1C2M+RM1QUj1jtkeVFLHgDM9
eAksapj0XCkO4cEyu3/Sd8iPCWvQq9Wjiksrwr7mHfXuJrrKFFwQ49mXJgQqia/CEbHMomOnUUNn
FpW+y23AmDsAIgiR9x3oDd/xcb+dCrM2mPYXWW6jBaWMW8M5XArmdFkAXj3byJ9X95wcSncMbhil
AdkCFlsFeAfgmmirIsNUR0MNMkVqnzwWRWl575iGSUt44rCcpqLshxllP50kL2MKFH4C3GWhjVGr
klG4VXzFbtSv45BApjxV+S41cICFXXF9XsezMEUHvQCZjBBLFF08+R+cjmwdhsiWQqmudnVCNFf3
/TRnHayiSM4pH6MA4o6yO6KphVjbpUoW/qUxbTwkUfkpLZ0sGQRoarfc7rWreOCDsOIQd0cfBTnj
7LKFp1pMhx1KBhNe2vyiyE2dgbUPo10GCDY5IY2ZYL0GwgovNWrd9bjeKBVPdPQuz1cfgonqadjk
/WnmK72gnidjnQ1pmPXkhH+tdGPbizZaPqog+2aMy1JOKCn7bwlxnFaiTiNUitQulbtLR/Zed4Su
7LddBbRimiWwq8eawQomCz5LAu+Xy7WKVZ8dujwLV6fWPptzB2vd8YK/jnm5sUXbZTsU8wLH9knG
YpOudd25ay44OA6GNaF2/QWSaJLKvUz7w7VhKRtbhF1yl7Ddg1OB2kKZBPDerVdRRzw5tC2EL7BW
77LTBuad+4vVM54NK2zPPPxoAZUSmG3yA//PEhHSv+fLlVxj53buK8WDdyBV0rGS572efTfzpQa4
QHYxyi+U9PNmJaxQEyFYLLOS944HVExEtEkF+CSKXtPZXXCmcNvM9kkTwrDJOmrvloDDw4u4vnbs
J0PkNzY6xmJRvVVutYmJCzPRrNTmgEdItrv7SpZ99Wu14OJwls2zZTOoTpxHbEst8ZgE/HTZ/1ie
+Vb/Xr1VoEgoH5/QuMYbz/gAB6x0A6LayM/5D2ROeFa1t62I4kiuuAiv4T+of/0hIaAO666CkAFo
Az5LRsZlocAOgq7VBEuZsGGFb3jQSf7Z6uHh3XukFYEEQDfjiMXi6fVhX5XqFcD5XfR0yQ9rQULx
hWLgY039HHI4h1CHuax7sURcfabKQr/Tf7QWVvu7pqb11tB8vYP7xnJI7vU3XFuOUDlQwbUvNMcb
mYZqJEMZaNdjUecAzqBxEcP+K0/yDmogKzB8GkqHNKVle2+XHIzKvY3awj+75ZH/rn10BtlZyREc
Yd9KFr4FnrSLFqXguiw7GVWeyrME82lZMJGuWzpwG/sUJQrYQw/syXfpurQNATbYxT/u8o3BzTrv
3qNDaV2ZBoqMRmvm0CTAg9KWj4yR+X6Br0pLvigYtWdYWxnJ16GeU9qvKWWiP/3ZtJncdgf1NrhD
MKh4g/MtelCLxRhU0Nf4fAj2uSqDWqWHeUoqD8UbH6b1esdx2yB28CSf5GsXlFp9jNh/L8KfoMGy
UXA1/64OiVIa4ns7Wsh0zgHUFzdyMIfuJiGAusF3QIzfJC9aTEgQIUBjOgWnnwNf53v/0s3DHKHZ
O0HZZw5ObYqPxwUcU+8wN9JFa6oEfJGCdkRCPwCfJBzBfhix/78fV2S9FLGrPGtf248AI8yImo4y
kIspBw1cgTbFSO0P+K7/aFhFEAitjRS0hHZAhgMWGQdLG7FWwVnX2BGGlXyDnApmxvj+/h+kDteI
z/HS4FiKqPefUkS/eZlBb3eacOSVo1Z6RuixvIhpJv09hVzmjLKfG2niP1oxGaFinxOck2aMJ1DJ
kFQm8pGe9vkaOQWq9yWFBFzeiEsFjWnSHekdW3nr66VoWArHW29bO4HrocZB2ZtFCU7VKW6CYXk2
1owrz94Zhkh4olJ56Zcgk/4xxH6JO7ApvOZwnYF4O3LBnUeNo6O7GW7WmToH2zTmTsDuGBsE9uxx
rHkVA1M6WyREGEUA9r/V+rLyi9JpK7J1GV9B3WedzV6mYbt36qYlf+VcjDxHsgsc9WlUu2aD1wgd
X6CNk9X7vTC7JbZb0SsL9E7kg0fIvAhMu1/0HoWYSzfXYS4+J6GDZULNTa++btYNGoI97D0lbFKq
Q62vUgAv+IyElydMVTVR2Q5oGPMM32aUcGEEb0NdaCYjt4rICC5VU5ZlqJlbKMbuvNNxCtW6TiVX
ZxvWIs+243AJy3q9zIJOO88rSJuOkyNomBbH1vsChOEhSPDnR+EfzVMlzAkNamqj25IKAf4yAoht
A013TeROgW/o+DIfl+wzIPBlJWvxU0bZinl6kelYT+18CdHVQxD4elPkON9OfNYiJK0NSrDT62MR
tgHivOTq52knN7NWgp+zm8NOXvqyQLrIMSU9TKcgC8gI/WXvWc0BF/a5SHCCqz+u6EDbAWTNRzHp
rEKLcXLDL9w7gWCXWry2ncQGS4FMAfB45tEqXpHVhV4k++e6utqqI+5gSvdKolK+wPNZsYPEkpxG
iNsiVZVsSu78EmqaaC13xrttdR5SONGP/oaj0q4ydy2J3PWu8v2/pHH4j/B0nnoqvxE0bTdfd5ZV
WKrQxe0DxikBnsNkKehNrv7uhU8JIBufYG9BQ2WQ+s5ceEG9npZu0meC9BGC7X+28aT68/CWCnrU
b2B8v7wyQ7M1gehHVz1i9zmWutbfZULFc/lOFpMfMod8fN6hF2rxaR4DiiTZm6xu9dVKlU+2lwwY
6AoOaElp3RGTdEHG750t8dWZrEEB6evwLHzWjhENjlVyH43nSJKEiP6+juyhLA/ApNXFG3AbPq0b
evXuJWrzQRPwfx9XK41+AExWFwQ4OQXEmBZvz2bluSfpCQchZYL1b4o9HzOM0YQ48uuzAEFpQ43K
elTPbsg1+NHBW5d+DuazkBbkhWppp2zldjYaGdhAm0nlQg9X+ihF6n6xJCvIM/nbku8GGW125qT4
scCJ67aml0L/5fWAWrskhSP25vdlUyXPZ8CNmLmLVCJ+YmPsiXEA5uVRxP4u+4YkUzg9C6QFZUw1
Q47etR5QvD++2mBspRvUlYLS/i4eXnqBTtOnSc4Yn5VKEudyoo1lVXYwS5rJnKH9n5iw3akrKSL1
LTnPm2x2PNTz4RdhJHFK/lkbuder131aTqH1AlqNt3MbMBEfqHFSuGyJvN6vN+dBrCpZGNuAWiWJ
+QrzcUsm1ClTjgdotzYUQnMnb5JT6g9cFdzWGUP44G1KR4aRiE8qahr72H/TSRhs4Zdvc3NFX0MP
3A6DBJm65lVlgi7qS18FOpuFvk250xDuM3oa/fcBrPSVHautS6UZA1Dd/yg4Ugit01zrAMKe/kHC
k93poXGSCAsyKD73JfKF/82Hsu0pg+iHosAA+8Wv6S1lS4jeRI265uMkQ9h4ylzFqe/H5/XxB9Xy
5WUnxem2GHpeLUFzZONPFJFtF0aixaUJpaGg0yB9zQ5vQPdABnlkUuCC2ksKwYhx3ufRH4X1p8TL
NcFloc4u2FsVJJtm6HpFCw8SRJVYFo0EZD/YE1u908ZY+XJxMZGhxhpcFzv8EEeYsisByQPaHI/q
fTje+lpPj/lNnt9EQl0604DUNvAshvkzB1rF7kaHgf/9vZd8hY4yUahBaraGAMoEl5AqqZu61n8u
YP7nT4wUgifoNOYhB3lF/DYDZOMdV6CNjIfHbkia+7HImJL4r+M39GfgPmoxW7Ph17Mk6MeseGg0
pZQ+cUvaRd8gjyr2rEhniNkXGuHgSuj2bH9pMN+GHG7rX/mOYsPzKePyn6y275OPdp83Y9mdQrtC
qchrGoUxpug9P7NV70mPXH1ay9hNlcgg9gdK/LlH2FP/9DJCzs9mpjHGvoshf+9B6nOyjPznOvsJ
zMVUWskiohXWlIK3AE85MSiRTgIQ5zRVl0GayBVSoOt+R1hw4yLsUQCQcg55KLD3995q43Uoe19C
2G7F6B7FSoLeMjiu7VbKDbrO2BYr0iVcjajZZPJBxMxucygXutB/J1V6jc3IK/pwwnvWtEkn/67Y
IJPj8VoET1RU0hmpGSoKf55qIP4ASj3BYWSqRZE76cOdwuZKRiXdHF5oMtddZYSVHe1QN4VPr8M6
end5Aplz1WOto3VMA0NakCJAGoPhDPg8PWjQ36oRp9uNa5lgGK1SfmRqZYt6hmL9E2lY+yNA87O7
c0GYXUj3ogNsbx2gVGAtYOVLzvhCrcj2mDoZlEVcIyPrSOd8W7VD9uIoGKm3WP6hje95Sj8N1VT9
zc24Qm7igHJV3pkLTePlD9BryxGoxredTRi3u1d3ObwdCtQeX12eaU0/jTgHoJ12Fsr4vTgueaqk
Y62GcYw+CDUC3YlfEGjK3XNBqCq5yV3yIDYECLf9EBTqPBlu4U5R2bi7N0ECldL3kMZmZlrB9XNQ
uzje/skXirYdm2BE4gc1J82q1gu2nN9S17mZdiFVXU8DCHZwS+h6qUWIRUllLN/h5j2bb7oWFLQz
YzsM+jBeu/9i2eLrkw1Gbvw1e6lp9SJPi7aW1Ofwa8i//jzmTtHrIlOoQJaxZUf1Lo1/CU07lQ+8
1FMjtvRsadX6Ek6RnoyDCTszLjYOqUCqkPnVwmN59k2bbFq789JaaPTZcVYAIVGsXFFsT9Vck+k1
ldqSEFYASxwqSd22VSubM6B4YAFVpGjKVUctTXzfHfjsmKMoOjCCCSN7Vucpo3t+5ZRFctSDUOOo
/qlETd+PvabcW9yzurnW1dmIrWl1kSBTEUWNkf8q04WozDb+G5A0qa3iQUDmnjheMhfMdBu+SBlh
5j2luVft2DB3oZAowOqvL8j7IFdk13a5S4PGnC1T8Ww3Hhn0eVfl1Zdds8AAwpFXyw/5l4/T6AAg
mfQRNKFjiCLs6AuMLhQ1VwtkUhFM2Dk9t0UxZF4IGGqgxq1t+DksYfQK80SLCVo/nQl0sGtBDz3C
FZ6usrg+z7lQHye9ycu/G0giML4dbT7NV9CCanKUZvXF3bdRAcc7uUDibY+2lC7HbofrgL0gm3BG
D5k30dqwMfP6FY5iUlbZbloo2JEPHiQgFI7SsZsOlpv0f4o8DWN8rTulxYrOP6d1oSxoL35l5a1n
OfhJhGtcSzhFXUzh3MyRAXbBFON8EKQw3NxzxL7uZQJVGdL6C3WbgbjO7pzsZI4BgUscmynuB0gS
uMdGzUJy6/iZym86f8VRPNDews67b5nUEG/ufN8FcPlddkNpq74CzwlxODaiu3z3XptLm0NoB2Up
2zoRtGm4mPAYco+bhKrj2X4oWI/PWZOhhlCnW2Y5he/yA8b6mnsXl+2Q22i8+t5HvZFxeO2iCfts
1ZfCQe8KeKczm3CHpXYRFw96WpCsTS80GVk4zsH1Q1mrvC/QqcVwXXTKAFGjZdsF+bLMysNN9GEn
2M//rUGSA4pDrp293AkK0Ty7mc5nvyU+brG7mJddny+WaySfqEU8v28vwTvNZ4JPdQdPEPO8g+g4
X/XM7bS+HCSzVFUhL7MSnEzE1ndhnk7uOlFSe39xRSKYAMW26raUxxQir1uRzDOdMJbkljmc6ZI+
nplCfW1jGtl/BkuaxQxyj6pK3arEyN0SeSt9uzgyV20r+jOcv6nSCZ42Gd6VIC1wkU6xMGLs255g
aj+nkndlHnSYHF/vFb+XuKgQ1T2lNyC02XjWEz2MR/J57woZRI3o4PazhaQzCBx+NSd+4epM1e7K
4B4zVmQksq2XzY08RPpqhV1StgWxWFJNeOYXnF8wQF3OZvCw1MvSl7b7xFC29Io/twHixFdpqq2f
bauZeeSDZjSH2zknDTCJzbt1YoTLqpLJaG/eDMSEAThZbS7xo4NpC3HdXrN8Bt5SqDKHz9RZbSu+
T0D43yYVjiGMhOfh2C9S2olqJok/Vy2RjvQeQg7cM25QAUys822TrYPzActeMJONePcmUmt1FdKO
hKkJDpjmTTPg86JhZ2FxzoqNcfjDPt7YDyOdRhRQwUTsFqIzkfKBsXHQPfSh+Ex8A5Z346ayNsUO
8VDoKXzGtV0U/aakj0+a8aQcz3cGNe+QE+7pWzEC3KHgewGoWJd418ZbPhNohkOUkZili+JIKG+0
i5CRXSInziPZS9FIQfmuoQO2hEEA573oeh6+agLYgR35oeYvNyYiqQiAm+mQXUTQ/HQmYIX7HfOU
6DKbE0SuQhMZlg0yTYmU6dH9VTH1Xl2P24hjZoWfQqbYpjtF0swsJpZShlpXZkpSql32pHHVBTZi
C4KfcedzXS1br2vjHwAAAWWVJ+TvYFio/sdRYeyjhjsC6bDlvYHJkc1mxo6rxPHMqjlFtOSEi+FN
auKVCLWHvNTmIdhrfx2CSM16LXXtLx88rdpIPFLGgDKqnXRIHagPZMg7R0N9CeoLpRRwXmgND75J
xXLDLB8oAVLYX8cVFOQ46oPHHNqo1LOq1MITtA1rzU9TgMU+sAMYYBOttPRUmb58QwWwTeg5kyHZ
a4j1pVYm/bapvF8SJGNEWOvYdrhIWLsVMnj9wI9Cj/OI+xesJuea0fgbRDz0PToITtrnGChLjhJI
68zmK4RuGAnzqLVCNgeHgXh9Nny5aBmWrXB0an0HDjE+KSjaSCaaM9S9DjsXcRVXYLRuTaF2pbv3
BGe0megfRSemEaIXfVGgtbhxb/oEv0c28uncKVkWDlqT1tkczLGQAarE8TlM1IZMrKETmeofpMn1
8eC/s1GFXRNkJ1ooVIEx2ARAaPLzugkPfkwX/BRpzmt47WQFNGnEncjS0d/CSNH+RM9YL2mX4lHY
IjmcmGVSBBJSvOwRMMrNg36dyxDc9qG9OahCnpUgHVPLB4RI0X5eKW43TZ054gAVb5pqzIhx/QNa
l/MQkreOjrwEPAdvc5jFmZBhyNbPjNJbNAIqGYcCp9FtW50t0RfYJxbAolzoZNZxG3MczlTAkBai
Qp7jGuSF9PKcZkMTxdUMW9bC6ddLi5gxroaC2kqpIjXUI892WbWweRr1pMdeDaztDTh+0RWMZHeS
Bq2kDuUNrJ1h3YA5IctrHbfNY49+mUvZ8KPviYnxBar9SWfD1bkQ7pEpBwxUK3+n54XuyuEk/B83
DcYV4Oy/4fLWPuNGyESCXn5KI6A+lUoLBcYC0CF87MZ8JVGm5i9MX2EWiUNUsMyUu45d+xM6Y+E1
Bw+unmAHM3oJtf2huUaIwhcewgmyij+J/xgBG9z5HHx4FKl30pAin23T4mXxvETb5Drl7pc9ey8L
oDOfJtQqRqf00w4F+ZWV3mAep54fO/7T2O35E/Qg70/r17H+T6Gj7oFpdH9+28P+QYuga5f+3JJE
+hvA9slyIL1gz9vzKNLk/NMYSrsvSwp04dj+1TXCRxEqY+e2F8/yzDdTRhJ/eM2be/DgMLSBgADL
wxjV91CqfEGYQsiffncYcZyMk5tq9E7njhF0aYET2EV9hnPhWMF+acPEk3K9yS10Sp5qlljKAEuE
VjIpzqQtblDeWqUP0l1mFfA759UuO6BFVCZ9tz5kkmYs8M4O0XkzcWHtCEkc+XLNM0Kp89/RyKOy
L/YGuzABUwY81kTbDE9ACchQBuudRIo/bgicC3T0QoDjd9JNvRb0t1DPUsyWMhcg1fv6usPAOUVq
z4HRrEhVNkS9kaoyrDNM5VpuhPgJYJWudSRDnktthhHgz6uSB8zptJR8ekvMvtK4qbqlCkJ5DqdY
2EMd4y0/9Wp2nAbq2afVRHcyeFG9/mkOZ29GAdFReNGkOJgMJW6Otn7BDAjVOoxoZF7Xr6SDOIRy
FvnslFNXqTGBO4pWsUgIS+FODauKqQXeKDBJQsZXFaV6GGKsxgs1MSYmfGRzKcHY592i+y5dpYRp
8VFqbHzv1HnraDgtYTz8HDkjqjrrRRmvrgxjDfgDLODHerN8mXYuY9SArARQerBel2DXYIely3z9
bLrnUef+aJPC5GZJheK4efqwekWu+60Q6LOO6gOrPZ1pPvPMQbWwxWz+2K8mULhiCnMMZ3Izq0RS
XPhg38jvb72vZOl3exhSpT7lRdC3/xuDEezObCDefxzpfnmz6Qs/MXQTHZQeNvDnNAafoCV3IHyH
5Rzoj5DzcoGpj9enFlFeDXEUjbdrUVCrNm3HClU0c6Aa3Mz6vBXWlZavmNucsQxGnEY82X4e/3Np
rrERDrNPwEhz5EfN4W+MI23yM0NMaHB2tfXIcap1Kzf6frDpLUWcReq3o/RIaz6W/yIYHJd1nuXC
Hc2hcm2rpj+V/+jJt3LYap0uf1jjJM7ONaCJH+f809asBaNGwDv/z1ZZxN+ju7y4iv1aHVGD7BFe
GQ/5b1t5PzAXmomeqcZBvx9zqGtnKiLAjAU9LtUR0wNvtkSRu/HijqGpuG+mHYaM29JYhJ+DERa5
TtHb+bRRFwY3YYUBtnCIA5/0FpFJD1wbtxCgTNlIxmg2Wnp6yBynE6EWtJADxEtUQHtorUWEuqms
s1c9ynjj/jHpNiQ7aUbg8BcQyxVWBgM7Sb2lWs5m5bcAPVpFEdZDAC2PRidKZscvyETSlLnAxgSX
xW/4fd+vkSPAKg6ZjYYni09d5gm1Iwr30565MGveIWVIdZJBrjHV9MKZEn+qEcAOg8XrcJSJHATa
sIBk4CCakk78K5QDGctIUZCCywBElTrTirGzNwZ1EUXIKExDSYBDgp56nRxs2th3yTxDJwoRc+1R
O/ZOeVYxJOXrByznwSHX0NbUwS8HqLpX9YFkHd+H8YeWOWNNeCMAD4ytukdlweuskJAfL2duza/F
t4/X5fUF0+RMFfdBykZ/Q472Ey0YsCt0usEuCe+u9dHSAI87RA/yRIegDHbG6pFjeeH17yXOWe/q
XXL60lURmlVwkL8HbhHeaAfSRil0hPuC3hpv/GN+NF7RviUmXz4ZCj2o/JY3wAYfYcwfprcL4L18
+mEH/AnDY6cvmT6SfA3YRDA+wVsaa1pqRDlcbNFHqoii5Y1GebwJJtE4os5PT+OJxSZxgAUnab6X
C6iqkTbigqDy0j/KaNtFSVNlPsjxAVCplTUlJS4ObCovbq6zqQPxFN7XGw8Lk6d3/rZnefAURWa6
XedQ+kC7T6ozjdOv5hUD5FIQpdUhRjL44sEkZiVsSdfP6641lLWvJ+fGy8viN6FihoEfJDw2uJJL
U1OHFrsQqMKt2/KpZ0LkXhW+mXuogvWHUp0YRImdey+MC+IzACItzbCz6WkQ95NDYWjoY/X7aXg1
ml69ubFaE69qdedSNhuaSFvOSmgIA4Cs1k06K3KbPrk/MrMhIBOMWxB+t94PvyGG//Ta8mNiV5F/
jMLulXoKgH2XLc2Kc298enF/LF23S0Chc5qCAPTRgoIcVDmus0UQvNvxVb3bIi4o6IUNKenX56pO
ElqahojZW4SVGx711vKw+YzAt6lEIzBnNzqB6jOmgOdyS+SNNj3qfowl79f/MQ1t+nsOqtmPCRtZ
1bqvAJGBJcbu9tzvMQZ+vxamyJgIgZQnNPLz2w4FO+58sYqEv8Fk2/AvJFiPXNuzF77R7XTCdr/2
dc0RPK3foq84NgVSVOtKU0UZAK/AbRTfNJoKlej4qGVMs3sWkKIC+sYn3yRqbgwPADFepgH8Vz2T
Mju1kW3KJ+Y+nHjfulyl91phb5W38knwv4V+yR0eXchwXXYwUSaEIOinFR5zPEOq8uIiCJ8NmydR
R4eR9AZ2K8I7RZqEMj2a7rL42pHlZ3VLsg/8D5v8fdO9gPRWS1Ms2hLWawstIu+Jg7Sdm5bVF7SU
o4mLyDr1DxE58dP8x76qDVbsCGC/X4CqOLW2QQqsm/rxzjUkXh79uVsKmlCmyauHukcvMpzaMZNh
hoy3nfDdc9YFMTjTtf959395yD6XrXLetr257h92HusZJiqI63lnbDmvuDHikqPEtrfQS8ooU4EU
78+KfcC2ggYOntuUH6llLyDEJ0sLNZ7/BXFlADQi2Tv8+xohAq3v+0XDrwsHgW+PsQmcxt7E1r38
q80CvBWTr6fiNY1zjFnu9wZcbwPlNE10CNy4h3QBc9akgCLuAGysYvlm5mkwPzv9Ko5r/toTOsgk
5SUuLUrXPLMxW74H7xrOLg1P6lPcROVhfs1Rpg/TYbvWRXNgWZ720AMdS0NjpZn9izzyamajnrSs
Ewi/A+n0DBCzUIgrM1bdaVSpVDe6ZVR7AYEVD4pUkmpEpNqxcj5K2DWCw97hYrvUnm6EGBgatAQE
XzAKC+O1gDSUQSNzou0dSHf6cIDWbmtgr2BJnP447usimzYf0BFn2bwqQ4i3LMLBsoTt1Dxv3Ysh
/hkqXm9veiXDPtZEmKIQ2f8wQj5HHRyyFlrTHrG2cJLrvm4Kug3hnV7NFkBJuyv8aISJ0CBHnAA4
RkRB/dGyKkwzR9akKEWOIR98/5qWZyAtYESz1b650OGO+JVCLqlOk6cfekWJ/oIG2WIaMCeeDfQo
ilF+mma6KoYD8CnV1E/k8FRySDo6EIwsOL7Oqe6azzVz12umO5yTi3ed1TeiSg8/yC523o+w5tqM
8i/fylinkXuD5+CzwTUJ3s0EI0rDkOMS4Jr3LbVH8SvTdJgLgsKAW8LoZ97XVnhquxtpSJdFpiDb
9TYl8SAxI8rjZ19hO0MV0w8HJgM6EgTcqlZdMyV/k5dykr81U/nzPqm7aS8KMBCFIHKOdAmvRXZo
hs3JJcuAqnxYwBfMaiXJzgteAPoUMPFEu7g0hmE+fwk28SEyrdfFLiu42O+Xcwzz0B2r3lZws9b4
15jVvgvRkot2iCqW7s6IRpWGoAmWYQGNc37RLFZtamCEFyCibTKpIDAmhliNb9SqBR8qdh93e0jM
wSL0ngN2/bJfD2OS9auD/3QZvyv1HKKSCymNVjTw3RQ2perIDP3DOi8O+Jh76b10dKaSSEm8/N7K
y0nWrEUEpgodO1kbl99NpsJvNwBHUdFvMfmD+aDtKmDCJwUnbQ4KhUhzKmTobwi5xy+ighH3NGJT
4ep9/I7+WxOi2InCQlxamPQ3CBytZ+ou6E2w4XkbyLac3os1tAikwO8sAYsVFb6uUkozyx9NIIis
1btawSB+C9B2eacr4RtbAvlR2w+tYT5ntwTqOeJOocF5YiP1Gjha8qwINsESvu8E+CCRO8LimYdX
f0PI1aB42a9A0DWyeWDstwRmCWju918nMJb7S5VoaMAu/zeO/TflRP6j9g7d205dsmgNrOVNewI8
9MS3Qb6yYST0GHuNBmreUe5aLKAIHaM9H3mDCmC7tRHiyt4msBgSH5AzsVnRu9BmRJJrWAXsDmW8
aDMF9XO3BTIj3Ry+XLDLQdDH8jSURbQ7WjptjnA5o+rZLf623TR4l4JDQoQyMtbwnWLuCaFctToa
BpTq9ecGp8NJfsDODgCfF457s8SvXLxkauYhfwMd8uGlr72SLRav7kUiPyqUnn3iEKe/6t3Phy3T
EopJhVsDOIDa7SSvJ36mpCpQhvzwSFjgTSyQT1S4ePtzy9v0/v4pJhBIQ7J2TXPow0jChgTqix2E
mvlbEZDRXhCY5aLJSgG7q04PxfoEI4o+mfCAJqKPtPaMjbfQo05ivPi9M+o593efa3t1F3K8Sgll
i4QwFv+hnAgRtSMH/KJy+sTjHiA6nISemCxJ+mZ5+slefCaSfNHlDpwK76wkvu2e+Ixmb6c7zL2L
0EGpq5lIEo/fi5ALHkw12PT5u12h/MisUxUKTbqWANr+AsRzV4RLLiOuulxIv1OnbzWgb4692ddZ
/ol7APVyRT0cNywBMHDkeogNsPg+/NrqNIMHh48okcxlZoLKZtQTFS2QLh/FR7+WifhhYO/6Wpjt
pDEtsrD3AJ4JvNQhYkYqupnUaXZYQy973i1vYYaYZbS+yo55zl44CDUo1ay3x8tIIO0BciUVs+rC
a0AI0MILTly19sEi2KZ8XWa9hXLn1rNFt6Km0ulSaJXCRnoiW/Xr+ThqH/ypPBE2L/4UcPNm4Wdx
3BoVMPLHLX2Bk7HgRMcWrspqG/kiYB1RqGb6W7HzKJ5MDjTehCmi8TIj/YJUPM0bkQJqw27Xg3WS
Xv7X7yuui5Fmx89WYy3GHZJxPalbyvBZRvUOX3Z3D1AaQn/f3/ia5cGOzH8fZyLaNEihqcAcw/EZ
UsjhUTIeC7cDDw3bQwuc02+LsxYA0NvbghY/KSF7JEkBrLzObyyLg9XQo9N2wEgJVC5s9UVH8VsK
Z9LFsNTEgLwA9JFCs7PT5XoT5jj6bZYN1PpgPZosjWSMFs3xC4BB1Zq3C1YAk4Ud+7OgO7sKhYyi
Bzb9ZY6KaTXaIelfoXhwgK6UB+grfhx8kw1+1q494uF/Wo51Mz88PXaDGYmJlRs0zgU1JuvLyBTE
5dPqVE0ow3q2gb4r7Znu1ZeDMC9AOdU/yMcob5TXlYbj/fEGbvkgIlPzSNW3WGGpG6kuJMtiiWMW
g9Jag8ukpDUbjSHSuYd4CWYsI9FTSK1WGfa0XXOxgWyTvX3m2KCU5Z25b7HfulIocvwo/yR3S6i1
lxnOIebHodw2bVRFonVqJJgXnWgDZXnlkpdDvkrvk8ZF/Zy9/fsLT3zV2G3n75/v6erGsjigIY50
PxG37ubBDMIcacWbrMAxRPMKjZtoZ7uHj9Hiho3JK6Acp11+SJpI1nqoVEj/R6VRshGBCf7nmXCA
n07Y7T/Hgf1uhjyMXhgsV7x1WTvy2cnxbq6aR70SnfJGu91pxHCreWByrDRCN7Yodh6MHZpUgfyw
1OX9LNon7/DrCyxgqZrye4h9drhDhjfLKjN94WiTW2MDH9296eUUUKIt/rcDJqoCO7y0Zw3R0JX2
COvU/wC5fxwhlZMjb3iZKHoFOYMBsaavDx/YsqBxTEOcKXOUsod2OhdmQm0m6IAJQ7LFDU6Iqykh
Zg3VJCybIHvLfrEyr8fG3fYMAB0pM9f1KzfpyLaZy0uc2bs9nwO2cgrBCgUS60cDUwmnuWPWpM7j
rT+stYb42CBGAU68IxQUO+eKmXICHb5AYoayaHUz+pkIKxqzL7N2fStcg3CizWhH4fby1BTYYO3b
pK1ZwmulNHrYpq5WdmExjek1NyuDbxWqYp672F7jmsF7AdHMAJxEiY5qQVqRWW/eR+3HeFjTWjOx
w2kOldfHAKgIQAm2bf3+oXvlPprxhCEfgcdvVRTJVMeqxr6pamrIDbvkGv/xRXkeUBm2udFHkdrC
o5Ok5fysbjyY7kHZZ19KeZi8Pc+xdbAf75+h9kg/8nPbuq2Fg4RA1fcFl1KzVniVDr6dgsq+j5cj
o+b7YabEfVeSqq499nFUTAfxqCBnN4H+7xJShYFIogx6mVLguxIs5an6udGBTLzQMJ6OwRMYvJEM
5/4plOQU8eU/6jZWkVf41MaqcXU2PsEebakEM8z1xW+T+YTguXVkA/T1beGBXHYPhcmfxzLjB0vW
R+ZyhLkviISzr+7hAn3zyhsMWnPRZ3vfdqn/KvcU0m4Fl8vbewzYLCrfI9obzi8XntBS88UR6kGA
yhPWenz1+WrNlg+w0WObflPRRXvtd8QXvgYwYt54nhFgD12CW6dTdohVuNu47B/udFyhNRrbKQNa
eazOtB876eRG2E9PpM+YUz8T8uJUlnL32K/oq7KpDPOBrDIwmAMpDXEONVLWHYVPhrijYfKic1IG
IBUzIruhEOH+rEJzld2TUTCxi5ovF24Qn16MCBX56eBwRLi2fUwTEWr9fjUp82dhzwzOSPOinNIe
/J/+k5h65+xlNRnGiP7q3KSr3jGr6VKj8Jtp0vPZrZJAXQCoE/QAp8AMGy388iN02VSjbyvGdzh+
mfhyVxhCe/c2MqARBJSgDnYbJqLZcLepzGtisPVNObWR53W79EDJBOVnDnRoShIlG3optCGsfPQj
tbpdrQyOd6slQF3LaiWWHaLtx/8iQnw4nTinOgTVHPfXN0AGb1MERGI3RdHdL5BOCdqGJjQ/JA0l
w3WW9WQTJro68nbr2JwMNbLSvYgIb/K8j7qB2xnvc1OYR/MUNOORBvdT58G+9wF/QbnK/3m35+Y6
8uPecGCylcfapVIxsxxo3OLUOIlNzHaIFCm3mPhgxMBcYVcyu3hTuyGxyTYYGIo1zCr40D0loAKv
gKldKDq8NuhWtWT7D6cc36gsUJMjTOUEi06Y/6S5f+lLUyzDsH4bihu2zb67GfISsurSrZ2mPj6G
OiXkHzmOF4KrvT3iFheqI4BdwZrdJwjFjUl4eg12/k7rQhQkVIqqFaEjQWJc0/2qP/7BcrR3UJBT
qSUlhNTO4ELl1moRP50KOhJ6kn52omQ4vA5JCH/zUOkitvTptDXm//DFgRAI+LhSeHhBi4oermCb
vIjCMTd3kMmULi5zkPnAq84+a+j/wTui9dPYP2hp531CifcKJGQdBLJd8jIhdQSYW9zCxY/gEarH
CWUQ/80fARogD7DQwxJmpNSw4s2QfRMJVIT3R0o7cnHQNLrx50bQaj3ELXGiUIsI0MXNPrg75wau
wTizfJfLQ92bu/GdRQDsZm/YIVo2rLM1atcumaa2cMyZ57qC43iGJ8+mVeKX+3Iu/QBp1UVnbtRG
4u9OVAEkIvEZ1bYlbj8yFkBUiUEXw0lS8JQntxRuKmEuWT8FpJYv+7JW8jKk4Gcvyt0YRo7/W8a4
m05S1Sx4JIZqoSVO90o2sBZAbmphWAejtcevftKUrwoIDGhfWdLwGPLaSPEQfh5peUzxMJqbhFQO
OsQkAfNxizgsucFp9kjx8CPg4EU8K7WKA6+9SeqWwPyZIBrIeOqnbvYFVm2lGGUMJFRPHO4GBiF0
4XokxpznDlhk+ejBYkLgJcnXsMkQLyXLDa1pNXldeLFYO+IyrGwM0+aBRX89vMRJ30q7JZHXLqiT
G/CRWY+8bzZQdy5O/+f9A+ne+U74qfgAzO/IntAToPl/nJ5QLH8oUfG1RmLdWfyMl7RWGFCRph7Q
nbUi25tdWP6j7gi1gw9ZUpL7SqgmXCBKGOJFE0v+/vMJhgYKPQbBTbCqErMCrwnTQmWQuAOX0ZSC
NkRK7WT3Dw4S0QT0bBEfVqpQdQ3bM5a5PKFK2ca8rPj1gwYezzE2Bwwg2bM5YD0mF02Zbu9ly4Og
0jhvOSEIPFtaCSvirS82ZY5LfgvNefKjHQZm6NqvFS1FDy45tnjToHtJxRR0kwwoj10Narjib+PK
bejFPb294vf7Ob2LeEKE+zcSS5c3cKAbSfTKfxd6tvfhJ79PLyHJq6+Pjnf/KYO8Q8iJf8ajt9Fq
5rpOdfb2stLR5WW41FAoqGJYbjvXNoeDi7QOQXnUOq696rROj6FjvfEoALpC3xz6xQ448I2iUKQS
7xJrslA6OzqAqnxnqbmuNIeXGksm0v62cyGgE1VFgZMi0TaB8uJ3IrOX+s9JK8dBAcDllAuJC+j6
9cHy6yU58h4y/Xgd1Nd6JVxzLrdzeZrWkesu7qyQj/wH2kQMc0xslYdhzjacShvk1jy8/tBN09sw
Pt93E7gX19HnW1DV+3D+KRk3+ZIY7A/3cDM+g+qWrce1z3QBn2xOPwVK7YAPJGgYLdduoZItYiSD
ItPUiSvPQ/+XmakooofEyUReApo/nU47MZxphZFaVzrSZjwiQMqAv/0bgwZ+8zWF+6eDV6VT2eFB
Y8xmhOkke6vMbbcGoI38A+6wjA7sbs6MIM0VyVQM7L1nALuXJtxp1aGLCfn9EUDfhbAc+9QUj6YF
UGzPPRYpNrGVH91OfG187qf5t6mTHLluSwORiRQnaMFSznq/SAeri5ZZVRdi9GRR66S5zKGxtzZL
QN3P+WB5n7HNYG4IZntbT5rKhBzhWoHd6Sn/UHzHIJmecWc0ZC5legGt0Df/RrJ4AA8SRmRrdrXH
DS+l3ckCxbSEuAnj3cgDEKCxPm4/iF46Z/PWa8k0c/cyeTvDFG7SGtf5+C0yDFp6jY4cneaFxYAT
uD27pAonLx6+FxPWXk6b1M5z0xBlIM/ova8IsRT5UAKnf8MgewxER3rolBBZY1mrEWJW+XaNIIbm
5xFk+a3YCULTqjhrTNaleEQz2zIHyX7eXmovvPbx+kHaw9NJH7/xTxqgFMeSfv5F7DzqioYzG4VU
OiNV44EyCV0AwqNTCnLdqApLiglpzFw6NJTSKa5/AoGQseBHGY/ADWOxFKk50H24tcBW9oc8SE1R
gL5Hsk+9yGiN0733mXBmIyNJgb18UTYGHcl0Lqoc7ptWBWEkBUlhaSzmewmcn6jzEesNQSm5HeCT
ivbYuUbv6xOHKC7xqpEjDWBSTx+wDS3bp5cbrL0HuD5Q7Ckwnyck4wOKHFCGmWp4tyf1LzcSakIK
j3M7WR09KB9ielRQgtWyDY4QnGiUtqfpC2yOIIf1zf4XfU38L5RO4bEqtooepXtFD/oi5prEhoLt
M1VzApzlsWSjYUdLcCGnNGNm0vwiALpvdJZgiF/sjegg50fKBJSY4YgeyfwcfQXjKbaUrvzeghqF
Pe/DMlCNk0izsTFOV6X1x2ckh0GtI8o32hvcm0MAWK4nXP0HGlWdbAEiPSUChwZMKltCrcRMpYcZ
FPQ05cO8TYoJGXV6PTWAxP9IZi76UAR4kVOP3S7OQhJXE0zoUoH+SslPKi1ehNKIplccsOXFUjUL
hGamT/KYAlHgzNPWyoY+IN/iwBKlDsYzUCw38xTTIsGE86vDnyMYZ+YhvuER9aCb2rIhg3uJb+Jg
DaQEJIaFgtyGKYTpF7wAXbF4s97gEzHDV1aDg67aFoncn8dYQCESbImqKBSOu0DBZlcLRLkIRiau
plocL82qmV17sYDPYczlzk6ghCKtDVllmbeLNwTdvIMOxESaANKkTe1vpUR5jDPv0cl9I8Ne9k+v
LGrJGIuuTv0OksLGLfJ0AEg7wjglP51n7txedJOIn0M2NZS1emDcuRQuGQifmVmpn7B/cisxHSRE
DR/0hwWZQciDOiX5mnyoYPpGjD8QcThwBqDp8rnzWC8LloHFk5XOirNybYb7kpLhcz5QkX8UPwhY
vx6+OLxltUltE3GIGIFXuKpndD9GR+e3tcb+csSovl4589RquO4WsUfU1CG87jehUrE3F9Hyel2l
uQ4yF5+7dbVKHTGiYUWJesCfjDUH0wdo6+223Q4Xot+nQSXTIKgvC/kPPS81Mfl8UOuThVuuZZEo
4N0aQhdYnV/2uYlZW+8HDyaKyyPHwxcnK4DKKIfq8o57FS84DfKVMqYnGN2SFNp4fUhTAAaNp2HI
wzSY3O00GGoILp5rkcnYyTClMzzH+3v5NBJlJssTbMnJdkNJ9QWqV1ow86ClCi5m62WX0m/w5HXq
C+QPe6h+XwFBhJJyuSXmzoxV0gjLIFh0FDZwc4yju6pOq12pGWY0psHLmVnfLhPv6VYertrJdLVw
tJAK7OkGabm7mk/JRZBuHf81e2eXQ9z3MTCNoxadMDh/ONlhq/0vflVqGdfgesXRkCM4btxRkuOF
6YYaWoqHeyNPr3FrLHIaxREIXTmpKb3N6V50hGUWLTlqglgJwbL2fnz8Kt684mYy8tOzHKvNInH5
CFY2SBxmuo2sdfupPSsV6ttxRBq9i7TLlJJMDVBlqTf/xLmH+XFZMgkrVoeP7yfi47UFUTlrAVFA
3C3fPnR+i3BazA9g6pKBbbQAqArt3wG5QmzoaeTZztl/EPcX4yMxP/0zVfxbWguL1L5vC9Ph20Bp
TibtgIBCfeoTxjmjTzlUAYAsSqWhztxWYiknmvRKD7boRBTcyF5Yl2YoM77POmbK2Cx6lo4KjrYj
eTfKNw0Taez0Z+Y8IWkhQ181dwgkMeHs5aW1x4LEVNSIKfjScOJ+ckdN8etyflKL4kcTEVfqfSDK
mvDchJhLp2bpUFFnBSkS1DgY/YNJDyF8tsD2AW6j23WIxOzkxgJp5dq7HkyoieB09yNTJ/38y1mh
oubyGiob2pgdCW5Ma2usImpViKpA9D7cF+928le8sWeZJ990navCPSS+jDa6b3IN9+fQyJYJxZs4
o/bf0BtQPkNS/5x7dkSPXsdEoe+UY90kgQHC57hdVXwwwA8NB4Kh61neF2vO5Q3wmmiIPdmsb1Au
fG1AYxNtqshzXa33yYKuKxp4GaMwPD8V/qxBcdJVMXG0B0E6hog+0pSfX+pXIdSJ7jvVxhEmVju/
UaoRO7dVRpYDXqpA9lYB+5GvZAfakZ6/YC0t8ljjtngHFpXHkiScp3/l1L71pe+7LsuBYIvL49is
+Int9/cMKdLBATV0THcmtBBXvqCsGs8xd4/6Bb+hbhh7MqnJibZGMne0PvG8SzU9l+WKvV/1kcDB
guvRAR6w4/jkQ4AKX7bOA11g9T7MwpDvcAXX0pNt7ZN0qSfufBHtuAwNQryrmNqXheeGDAbuSkWV
sh3GJOKEdkALeFz4CIkmwE55YXaLl33vWEYfa2c8EmTiGuP+d1SxbZMGd6aMy3pg+EfLiG+kHMCR
rdEhyqDBxLtAzPxaeu0cWAlwZk/jMitx2FitpMX4PvAkAzo/sQKJQnMBmLfZkFbF3+4rci2/QG4O
Yh316lq8ng3Dkw4qHz5F2Mx9rKbg/RbVudxGvQ980AKrWifH1NxZK12aBhzhquSc5LcqtdAyrUiO
uPo1LM9+PpfJIWlOEfqHa1ZoMetG7xyi7nN3n3micEA9iCJyAO9dUSf0uaObugtIvr9ZRzm2d3sD
yY5qujkDjOZ54A0uRPCqsPRSI8WnOa5VQFhrIoJcmypU76vU8yGjAOrjCV50hS8zazq6wr6C6Eb8
fIc5yYU5kzuSJzY+Fykt1ZtxaERcFWQ477YGkj9/RVF5j14xRVSY71a+/RrgMbqT/Vw5R9NURU+X
gO6FP5sdCTqf+zRSmou3vM7uv70wYyMecOCCwidpw6KYV8x2Chx2QktIY7OGKMrsDgJCggnIBRNe
oKep634ZuRhPcZoOatFvOH+mCLfqfLs/IcH0MEtEtP9NJIhiYkEvcdOGRPzOtTjBuytdV42tBBCv
zElnecUJgD2wagEbtq3gQVFZFR6kk+FpW1hjoLcBjNVaYYWsxcfLuQDMvb2olXORu6NEFRNNel0E
CLlWuj6oJAFANDKlItcfZQl3Da1qP2W9lIKUeS3iCKFfSi1yYdtZAdLt+stFhkUzfFCG4K48secF
ebBmD7bKYoT8i9zOps1V7ryAojhZgLJKUq8yCoRReGc8ZzA1lDVXm92JpXqd7peL0x997f7APWIQ
006/EZcaWCn6dribRE/nDSgJ4e65LJX8yU+PYHHf8JvOzBu/JxlCVYMykFyHRcaECBnPoLpWem42
Qu27ynr93Kfu3aeCjcvY2r+UJtTCZ4X93Ek4b8di3Z4IsD2Cc7vPAdmmSH1fvg5nYJSSzOZ3braJ
wyWu+k+WjjiTOlpBCYzkcNfPdtFCzRbE9UcIS7qPVoMgWcuG9N7dLQOnCsOP3ovbKAVhPaNEvDrS
ACdrygUNz+GfYEsaVzF+Zj1Lme4XgUiNIQYREwhbDhh3lQtydZzghxnYSiL/S9Hg0o5jksl/uyA+
HWqu3LJZdiqryoOxqx/2gYg55mgsJB18NCRipf6eed91Az7D0lEHGQLSHKaY+BWuXGk1vAh2EPo7
V2bn9rNRZjsvPJLy0xbn1AUAo+Vp6Jek//WI6SkjSlZwh6/RY8/x8owl2lOTvO3/tgUalZE1Dm6K
GSYj41StzxELDgbJpjgT4uAm9wcxCCW0lwGoI8HpR7IrOFur6uIhKs2k6kLGxIHfLFIBgv3Qy+X/
dE46YycqzT8vf66mk0UtzHDHPoJ3SsnRPREb+LWiB9EzzQJ81ZUR3pQAtxGaU9sJDHbsxY6RW34v
omeWydNDp0/EIeanhVIZusYhLOnT8mBeVp3L11qrJYqCmNVAyRsnMCAYsSDmUNzCvewi5rCHICy8
Ozm+DcILkX6H3M14NrJJAxjGejHIrpeFCIGu+RGmb7tChxwqnsU3yFcRGDLN13pNxATiO81c9pkV
M6vXmAE53RhkbMq2A6eNzbEzYLTQCXtSM8AC42emzgcbt0wA6Jynv7TiuBOOlcuThEZIqFfBO+eO
esIYGc9gGcBN8ZmnCn+NKinRSFpRBCRl7pRAjCfB2I3HjI+O4AOLmjF/+0yTBcZcRIoiCgI18ZWO
qz1ISaT/IANHEHM07ZtXAEbU2x5rAD4uI8hPY/u1tSkdVbGvZ+D5utpWaVcutlbIQ3HkfU3qgMoL
ef6yAO0s16/k+j/ip+LWv2gi2Btp2Kd5+E+qCpD8Pd9EJ6kSSUgS/u3U/Lb+cv6A3JhJSeQjTqOr
zEqmOZsnWcpDgu5IGjbIcImv+lHeHOm9wwYxSiMYhjW9R3P9VeKjHMRSJd2v0QEG3/4I9baenLf/
ashzs9vtizPdWx2fTKC3Wze/JcECqSkc75tvQsE7tMbMK5hvRyXbvdDa4jRiHAEQPornDzGgxlLZ
K6MMgw3mmTxAitzevnQRy7h/bbhFj8wK0NOqZsv0BENg7vVp59N6zcU7Z1+gRmMxSNhOsMZ4V+BW
YrnpnWQFxh9lYXNtt93rb3tahlbd5xfEXBmaTPpHp5RFEwWkkWPmw8HX4lWKdV27DBXPO7pTxZu0
qXXxb0swJrzDDH4OcNjfnOxhtqw+i5Uh9/dHlbosa0jhJI1/Kx9BflxtgZsaLm7ARN3E9jrwusSU
tvBR14IyHr9P7oICb4YOS2ivv7x2uszLj0cKzOMx774syATDhdbJ8FpcF/slsj54j+FtyzstKav6
1VM3mCEFoXHnR7orJqYJrODy7GJs9KMiwXCgPr/Ig2fyuSYAK25RDZCkmLwkSqCmhy8B+ricVlVd
S0RBGY3GLu7soAEHFoEAW15hS4ESjGFXAu573Q6oMMjYNqIa3zCvW6zZtknwm5SPLBhiuX1m/0MS
j8a2gyGIbvzpxUmZS5wSrRUQ8RtQlOBYQ6b3YnQI4xGg6FHxt+VQDhpbUjzFDRDj5YjGGqGDsiLx
hUIFK18r52cBGYo+HpnwdY4ql1aOmjMg82CEdfdrBuZA0xqoAm6V1aU4MHPS9oUn1MiYzbT4tuHl
bfINZNGcmchX5AbJ9CUn0e0ga32Fuj/9261aBkTkG4jUmFlVU5ltbhaLqEvsYLaGRUrVAwwXjBKZ
f5rKwjwU1hI/fRsZNnUd0hmlmDK9a3gfjBm5NdvqWDb3sBOb+KbedeFNQjZ6hc6NbMpCZpmd4aEw
KwN1A64CeMkACyM5TJ7fag2cqWus7tUumE6XtpQe0SsJf0uRz2nuvrIFeR2pasQJtKkkEZ2R85rH
2lNJfG3j1KeRUdKf7a1ZebxOkpFql56yVdgPMpo2M/62pg/n+TxZ1hcNe68npYJ1pg+adiwMOB16
AnJ2sqkrBJEdlElmMFOfn0pdwkiUx+KZlSZHOIUpWBCHPTYNplRgw5OJrRHQeVOAqFMxxFFtsWaY
HzNa55qGYSaRb9oA8Y7mad38nE7WKhUi/5F1iDeoVK0gC+9VdPIWhvkO0WrFlRZiMmJ2E9lKLS3g
3/WuSMvRKpKat49O7taCdnrYAaTpKu2wDrRs2whuuzoXrSOERna4ykxIcxNZneJo/vT6D++O4cQk
AZokHCIXtuLZ0CRHK3qeufMY4Q3gYJFERnmkBSpf9dNuvYXnwwo+FoCi3dva1/RcqUXYS1UvK5vu
pFxWeSW/KLN5hbaYr8gc1BAslSHuoqbPzIjpLrBN4EUZi+qppLYCdX3UgvBF7mLnL3Kl6MUOCqWN
HAEe3Lk0Xo/LT3Hq7aleq+W3Dp/tpJ7iVhSx76pQRzfawC0Mqc8sV0rYJuSLN3LUNlLppFcHZck0
lCkN2P/ZBJTy7NQoVgBDc9c/w79lQycCYR0PeV+y+B9UCjKlzd/ZzMT94gcAMoBrWBgFmVBc8DFY
DiEVYW1ANoydRjMKgF39wVfRNjQ3TjTxJSLmH8ozN699JE6gvTum9LCTK4Uo9k/m399LsvQ+u4pj
lgMFKxIiFRZMz96K2N+u2n4vqTGOxuojBOATFFA5Nhto3hVZnPEsgXotubkJLlPdlIP0pzp5DM9C
M7+x3vrkw4wTvCaabexMI1XsXYyVaSjiazeObV/LM3b8tWN4mmA04IGIkr7/HNr01DHrFNKKFPtl
2L3onfxXydJWd3zgcqDs1myXadehXW/PyzcZkuCYoa8DGD6FFuWcqQ1AYCu93hH8w8dvBpSCpzPD
TXFg/gRyHqdIedsgOouRN7roQwVtm9AaO26gEHpEa3b1zUchR9ANX3fAz9w8pgKC5iCxD81Qg+1Q
xyZhVme4S+KGlw0oCZ6DMQVQygN03GjWpysNcL6Rax/Nav75tiKxh5kpmhSIOiUvBKaZwzgixN+Y
uKA9Uwz7a0UcIxGVVQSRA4pjVnzgb6YiM87m4yZsx8koZuVs++Oc4ooDoUc1slj9dJzzSv1G08Kw
bMgv6PtRHybq98Xobu4InvlDxWjQhzIcaTFTkIMQKilPE9TDiVwJEo679snB9lF/f79mFOl8iOmR
QgtWdSSPJM7SrO4szxtuJQGm89HhQl9nOJ16n31kcKXmNDxqpgwAu7K4XNLtNUsH1wm9iX1tVgIM
5y6S6n7lC1HtJkh7WB5sbXeWNf+gSBukYO0TX9xHsruW5CtS0uaMRyUFrzixMsh9ZKyELO7Ut0zs
HG6rx6sNg8hBC6hETO39uYnIOTExEGBz3Z4Rq28AXXNfk9olNCozix03PvIg8pWFPEfsJ3hi8Tdz
JMl/6UIDd8+4pC3tQO/bNxhcEcJP69JyreEvghfau84Om5CIKgT0WIaUXjCNz/spLQLkKRvB6fvS
bLE1mFsJVWpHwyKLoKNE/YDOos8DxZHyn5D7hzSdiVRVlpfoiAvht2lh10pjU33nISUuM7HDNQK2
GFV5BUWuiamRAs1042+G5mtMnw9EDlv5C1FqfFDaeDfjN73Of8IC2t6zZvoIE6OZCVmnhISJLhEy
5hnM8ST0GkvI6EGIxeG0m+dslmtdUMw1UGn9wA5P1ba3nTe6/1F2JoY99w6QhIVdLY0gb6pp5TBz
vkA73yvQCJ+pgVL+V0fC0D+l1rpjEE3Z5TFgyQjhjDpFEM9FzhGRRcsrThZm8VFdLnrchw+Db8AA
jBWyW8my+uFARj4jiHZHKfXJbPt8vunxsLpbKQGF9w4LzF2oi86lcJe6nwSGBxx4BdOxGAsC7AHl
peKbGfQC4Kp8gn/5o72eGENsQ7T7bswV29GSmN2cd8RAn2g+NX3V3FV4MvcunwpM2NTv7UNGCGfH
pqtNzHYyrnDCzC5zORZ7EAmdMe7i8JlViGw7H9iaJsmp5xmXlBbwRFHbg+JrhmzkqYMpFR6V2yRB
tsyaCxsAPYv2RAsuJapbB1bZaOBOMsPDZmDCLN9vNgDBmlWg40uY4kJLXSXdip1VDxG1bX0uCTi+
UjjffH210ARIxwQx4YPJukM4fuwSKi+us5cW4c/jEbr/Td16HYnmO0YYs3QO+cNMxlQn1e9O/5eo
zqSkgcyIHvFqXk99JIt84aXQMVV4ldYjWqRfyiVcPVuwwYMh1y3zL2qiqXKCgs+zT6JAW5OYaz1w
nDHWsqRAHvJZccz6/eBazvLX1vy43ndEJRdEcOg41WhZ21nXiRikO74rae52P+r3nZcbLQxfSlKM
rkO8+ykDjoAPvQ6dIETQ5jcjLt9toaKTCR20SyYVH/3ROWIhpaXv2GgEhACS/FhubpdxWjHDnAIj
xbvDJskek8p5xJkNsqTGqVnxZrAChLXU5pyddkmvGz5Ibe+zgLV6DB7gi/5OoSDjgyBbLtxlQN/b
k6hR7TM5RlvGzeLzO34/tquEFUHBhwJ8NYGBWRaBkKo8KSaAlRdidyt45WhkP+o1QBcL1d5C3lSp
PVpvzvkgo1mJhUAOINcQZJmCHzApMVEufrKLPZMAvvYfDxshP54SCIO9yV33CXHXQmpP3Cy12scr
P7L7drs8Pyx8hFl1vFl8sTRAxJ6Zm8HyU8Tfq2dMURR9Q+sEaI866BQGbyp60y7UponHH8kCsaHy
sIPzRJCZgkk1dhcLPye1JMbGPmTwxGDc/JEoBptT7BAr0PA2ogPmrcy8GomubOciEiyAK7mgbver
G0OSg8id8UH6BDk6D3AvOjIoHUE7iyUC1u6OKjJ7zH367SMgeQyYAnP0HCMpx3pqkBZkzFd+U00j
G81XQVOKQ8tzmQ05iZ59ejBJ/AaHORrVhH/wS1DN78XTEqZax36c0Az4z5iLmpdTWjyC+GNwJC8w
WoKCZDk9l9Yh6qDcR6AE7tFXuHbjvEkCfb8Luvuw0+eygn3IhKsaX6TI40rWXN0ssNKSd/VWJ1l7
H3QbGZXCbSsbOZJX4kjQ7236fA63yiY3AO4Dtxt7fCfwSp3ao1WFyPauhSI2RKqjaIUVk5nSHfSR
02zOJ95d/Kv7CWP95aZSrbInCL4Ou0JrOzrMSPMW+3KRD6Yu6Kec18vCpEJ4L68xqFcK04rU83fl
s6HwW0uCtsNqUCednEG1lWtcTHlMCXQjNOhQz4mL0zRdR9JTaEPH7hBJ24kD0L48MMZPVVXNgOjY
sZ4Xo2RqAze8FFs8chVr7zFBtKkOM6g+IzkJl9RFbSa7snY8Pe5h0hOqzZyQBKZNtH0iRH3AOVUX
S1mvOkdDzjKhpwDl5i1oov0OLCx8i4dHPfWbi3kPMx36cV9s4zhrIgMyXDMZ6YBJv2THZ25vJO0/
a2ypeclatxl8LD2gcRi6LixZqS9gTVlXB5OBWGVbMtdvx2HcEEHrxvWUllPpuZMz95tPFKyTV+n0
n5VGcEfN99xiXSNhLCNoo9g8z9YEI1wGYuWWuZqNTtx9tHAmK2qMIk2otot6LHPxxQYaZ37M/pmr
1vO7sXoPIVL909j7j71fYbKpqVDKMr27Z/60eaeWmHw4wDKUiN9vAQx9D6AXC3KXg8M3RHy+b2Jz
nc62EnnoKsJTB+g3S7Mqtd4XUHoHuWDTx9ntUKiO3o93XHPlhnT14ExWTdrNVF+Nc6quaIMU+1Vw
YPMJ/Jm7kzhJDLVDOMit8HGYUj1qGwFlqlX2T9SBHkCfdfD3kyWoHjLdbduVGdbI35w8bue7DuFE
D4BGGKp3gExVmgZDa809XIl+XOnNlTnm8fDQtRXspfTs/JMG5wd7BNvwYzsjXXbNzHM6dl4BCPCc
FrrpsmwZCVYDiu06r4dLD0jXAjQ7xr69smry+9V8DhBzfN7Squ17kocQ9SbFHeaU70w7j9KuCz3i
xEm7Z7+5UxYOCRIUP9d+kE8llEOJaakC8+efUpwX48cxPRPojb8RfJzBM1oyTPX0Pxuw/k7TDeQk
Qbi0jGBMvxTS8OvVOidq/IOxDPmJmKVwh5DdlzWAq7B/jEicZm5U7V+3DSc8RM3zxnqCg6ixhmyw
ADdUrtXha573zHY5T95BZPbuBH9n4pmNGVcXV4b5rETwY+6Im57GpC5fA39uzb2eziE5/9cVld6p
WpeqrxlneWVEk9ezNRzhnKZLaf2nZIyWhRu+R3g/Gjo9NjTXFJ8NiVMYDaktNpvremaxFtmo2Yvx
Clh5RCdP8tN6bHGoDvZQEmojCYmUGp367LnhnYDoPnUAIwuP00pH03/pIQrS6Ex/C2Jo0nho0Fgh
BR5nGJ2129w/izCyK7clWVI8xZL3+zvZbKSLjSoBz1rIG4xAIux7EiIn4ImwMJQRQcgWA6QYhUx4
byw7nIGuytX+MlYyPGVgW4alkqBZvMA1DjQpe8j0sVJfvjULbHGleKs61CRZmgKe/Tvvh1q7dWny
qPJ0FQB80mZ4S+XK+nMA0JzP1WruQJwvL00aXipuH9na/QA2ceKpjvDNKLJZSIepUsFDzqLpxN9Y
RFP+/WIF3/YV6RVt1VrcnrO6b6REA1kQimyd2dKbvy/5uTRBH12zasB/oDgW/qOerkWm7OCbkuQR
FMT+akE0RaBZkIqURfvWdR4gdMvoEZajyo9BFoCA5GqkWRmnwsX27MX6LV22LTk8KyrUivMBYEuE
oARtm0Qg0YmpZRqGcX+QbzZqUUyseBIFw3vv45T54ea4VkealQvnxH1iSyBDbJEijOhdMrZ7Jo8b
uT+nsrOOpddzvoBnRA9EJBWdfNYqQb39YBIElOd2UxlItEnNC4enin7/2TF8muOu8tYSebGBJ3Cb
U1HpA0KfMpcMEykQVmliooRyh3zZHnA0VjN9i7tKdj/FshzQco5Yoh5UI2zRT4Hi7Xpj4dTDszo1
r7CTtIQMsUImwQdZOjzpqMikNz9KpFMFGmkLOwaHph+/dEJyByqkcybJ/NrVB4+E4RxvCONoWLjE
3w/IREdXwa9PlK6UAe6L8xSSeMws0fmouE7xKxd3wgJ3ON70QxMY33xNTg48lc+qj6cCXJ3weQgK
DumEYieBxDIbzDPumSgaLJev2xyuPLwy9O4ci4eRJo6HY9mZxhyWVHIE4uCLpBEdPejqkdVzXukR
unvEYHUXkl3ZsumEsVUqqPjxsP2zIuYUEhtAMRYf6KLsv62yKqjLqKUz/bHNaDEi5x2Z0cCc+c09
h5i1wHv/svP92fkr6RLJL+yY4n5W1cCp7FDC04/Z/54WjtdreixPu1+uPWqdtOKwxwXoDQjLvMUZ
2BoDYBGbWSOsqCQyM805Pc08AUxx81ILMUlZ+8ZO5VDXkw5LT3nlJcdBJ4lBYXURfR3I2aqNu8ys
PIQTRi1kVP2scQHZt7IgBA9bthcU0SavPZCk1snqaKIkp9lg/CjPhFezLZYVFhHMQ5yyuDa/DfX9
0yv6EYxUZFpTMpcWg3/UOfkujyVEoVmvQtGBr02rlrW8rO3j9AH8qHqnPIKJiZascRdylSS2iryJ
4AAUTTi3ohI1J4NsQ0mZN6/mAxO5pkBso3/uVadHNT+NFLb0yvMSQSHatfggr2PrRfDYt99S22H1
/BIEu6u2T8eT3GdsnYP8fV2wElKMvzXYLKq+DxtApc84QvycDKQKb+iZQQJ9bvNbX0K6IpPvETPM
vd32SRIKy+o3tcxqdcunAdADy48ysIJxU4axzhs5Lvf4xZjw2xuzWD8XDq7DtFX4LhHnlN992gCv
Vr7hWEDFEnaQkzeLoEtwDuEe1AFhk8Mikxhx3WdCQ5V4aRSr7QbymzjcebkCR6uBxL3WkC/69TBZ
8f5nJY61dLa7c0fhkqamGw/GoSw8YWpKK1Z3JxaoOPtrdPUtp+kN+qzq8dCzooYb6hXL4iJvGrS6
wqc/RokcVhGTN2BflbW4G0JMg0MkJxaB9TH2LeCHkS4HQ///p4tRS0KybciplMHM6lcNVLuqWTn5
ZkgCfU9G7/eSpke8HM5fQCtEQGo+tKb8PBw1NlHUJ2KW3jnwBIR2aqg0QJJE7wCAENTQJzrgDk+x
ZuS8S3izLsr5kncY8l26wuIcDl9e7U/eiXARQYZXauRRvW+LZ+sALxI9LIp3/VIafGqK5/d68sa/
aewoQRiVGceP+M2TPgx0JmNSF6j6cNZxHQ38hFdBtVm//42aK/jr8SQdTI7sVay9IBJUfkPbD3QH
aGJ+7Pr8/k79k555TTh9Dh7GOu0vgfuNTPMxcdu6k9mgzrDBXIMzx6IquUMk7EhOdm1hQCWufPiG
Er20bn5dWE9qJog4rPxIsqOM8ww2zZqEsYU2rY4bx4NeFavjr2gSvD98IVDTQDhJirrhZ6kjfKS0
YJwytfxCQ+sYHubC3EJM78SJ1xhIPsuQa85b4qbGCYiI5o0w3jT9lNVNXUQMzAwD3Azd5XDLUaJt
OK7MeUBpB1a2B5hnDm4sFhR1IXB3Z/kg/kmFm9iP6N6VKzbs5gUdRFaBGB/9VtEpgQSsLzhPWtZI
2Q6W7m33PSyut4GP9sWlqHoEq2m4qWiMUFo8hLagFyfljKv2JvmyNstJ61Vjsb5e1eyOUMmKhdCd
nr08mbTehh81NFgLLf/e3IJJk63UNiNO5mntP69JX7FLi049RcBH5nB3wToYU3nHyaADlgnbupJU
kUQTqBU+8hFux2rrBRcubeLAlaIlMclDqTQur7evCr+iD0GxCo9EFm/jDS8xC6GAVVROGlzXLZXW
vclBXuAg8YF+kv1yFcbdCLOG+HX3dvg9vnF5AMAp+/1PM8Ai8eW8Bt6VgYXPLBgEEqH7cEJEZkmt
91LmxbVIMARgqhuwj4ErL8LNJZ9QAxK8KdsxrqxEh+RTxHMkladUYrl1ojMFO8EARZWMk8xG6Re2
SMbgCvNb+/4Cxo12oLJiytsmAa+d5pxcvaqKfaZWS2NBY3dbRF17wxCrTDSSKICaIUPmba2MMuTm
X5VwfVOChpPyfK8Uj6aQRDBOEdIFrd+9msLjfVrEBS9xj7cdeQyMoZQVYWOPL8+e9eWUNzCcQF+6
R1Z97eSqAlmJY9d4Addq9FAUS5kN5eiZNnwrI4MccexaEuOe2gq1jUGYRpRfYYyFauYlnET7F2Q2
WUxluGu+8zP8mOjEeXxg3GWiGX9jE0gMIYtRLzpnml10vLWUdlit3HRm9RtIglo//0JIEq23YiyP
MZ/u4RejoagCqgsBM9ktzEOhKdJe39ELC2LZF522stmtS3GFFRlDXaD/lgmYYxGcsSTeRhGS6Q6L
8Y6scJJlWil2MLQX1QaiTu5R7CyIQz77871deg1daD3f1cuRSydHs/YDawwCzGVW8m83Eu2kT9wL
DcuVvPVWpFVjmUAVVJZhwvpYk2tmGJ2vGJIAHYcuGojVjHs26tREwJBXAVhdr28xdASQ+SISdZ7O
UhUZCjys7Cnh3NiiFFY5iJ2OKltk7XuOMiPXZjBXtEIyBb+aP6ZCdMetn4QQowvcrfzFgOSyWk/+
x8CaHDH1Jbvj6Ib4vYIaogZTYssDI6iTLpm7fnFFO6YB98gzwv+S5XerhK/XMtP67zBaS5UcNlk0
/D/o6JSQMR1QXR4s7911ata0M2ohT1iOqa9mKfIDCzxhFKzEcfLPz8nns5S+axR7jHzI1yCApc1b
tDNMUL0jvcLm7+THQKi/Gdg5Ii8WvbhgImmqSd1Riwv/2WRmTA8Mitj8kluO4sITylwtZjMwj0jQ
QXQYImMi+KHQauHu/WSC8f7p4jjVgelJf4Z4B6v82Q2TB1/T3C3f46z7vPLoLW+EipTKhyYMAw0N
MuMFtIGbyDV42rYDU9HcLjRgapXlcLh9M7k4ZeZAhI8a46/MxjhSBrMwBXheJ56uPNJODO5mYC0p
JFpdIdb/B0Hz5qCJxm1V1Vk8602uciCya7KiWx4fnx8zrmEd8su7mkCxya9CqQbnibRSoiq3x5+K
TAspqrXxY5xXI0nG4zK01D5BtRMHFGEwfIIZD8oi4HuO2Y+XQ1/N0wSrSkvpLVSfqbvhPSZn333b
C4HO3mv59Ob6No0qgvAByDL8yiK6cOmIDTd9n7Zmz3oacz5ucykyCzM0WAbmnH9HyIrhnOZyECOV
KXpi/Jkv9z8muBe/QysNNsVcF/yYOPPyCWHPaFpRjcBwOQTTsi+81/9XF9TE/NqvNxBZkMN01spq
Z853UK4RI/z6orRYfPBwtalUbL5f7wle9eT+M7m7a1OsIkdPzhlmkP4WooP+qm5yR51irG9unGJc
OxKAsJgCSS/gFleN0Yyq/4yUMXNkr9fI9Q28AUvqcKEIgIqQgyA1W5nIpvmruuzLKuVkPF8FYC1L
Wdq5xxh7eZCtOoGmKZBdHYSxNfIvYykjppGgvfP3drcN7ECdJz95+dkrDINzhibgE6sQJURWkRLL
FFGqPrUx1wR3eMVRAPeeqhGgZ6feTxIsQENQPtv+fRnmnEbBDbk49JpfPRJvW8OZtfWDv0hYjeeu
I1VBuWYJ2c0+1m5zu5kiOMo9+ZIeN4I6bGLCvQoY7YSOHWMAUcb+ubOrUwAdT8prA3vTADO0BAop
K9tJTcXltfVUkhke6a8bz6a80i3eGbCgtBerW8cn40bcJ0qAMCm7LznwmCuTdK338EGTxTTXDf8r
G7PSJSI+/1WZHdUBeN3U3CBRoym17g0MLQrHRf94iirFxFSQPLsoD3+e5qLSnFFNgrc9okpER/QK
De9ABiOYihSIq6K3Ru7QfKHvc+fxCQIGPLhp1bPm5x4jbjlsbPv/gJjUh63fht1si6w9/ncgf6eR
3bHWzqK7HZt8Gkajo7tx87rl2s+g0U1zUyVKp5POhcZm5UAVGbauZtC3REbar965zrdz51va+Z4R
TcKRQcbn/bm4Grom8bjm42d6y3aAVvYs+QHa1mwLJK8s4hddCykA1WbLXtL5T4o8K6dMYfSHv5cv
Gn9mUac/J2G2XzwTiGarUbkCykTosDPQSoaRl672CFRnHZe+sEDQNfp6RG3iQtP6G5HEwtT2cyu0
AxAOdIFDVlmULZrVxk0FgrbSiVzEm1xK26Pe4SbGpPx9myxzdXxu0yNrFZqFz5teW5sTgJG6RyWM
eKAem7pUKEFQOfZ0ujLHWu8D/75p7l2kRsJwZdoP4wlINeYL0r7Abb3e3of4wA6feG7NO1/JhWp5
xTU9V5sd5XRR3hb6dRUQ4qrhmPwXAyWEW1EF44Upx1KDEEjLE6NVJBEV72U/LBHL/Wk8/2QAIKZl
KgT7V9blDXX0d/p68e5UEgH+FmAM5p6GqwHii1NQkJj9FCNddOw0pKasO/U9Si3hoIgTo1XuPooA
/B1jo41uEZgNNyPrWxWUMKGcRmyyWOwf6BGlJ6fQmvC6lDJQ0zvPjFWxTKb/YsGlYmdz068+4oKt
P13RZwaX08XlHxguZpnLS/ig0dKHLeD6dkTs0hvAig4tzdlnXK/zZJRLS12AxMRLPrjV6nCS9lWs
5LqEPcnWgywrGCIpM4V/eaavP9tN40JrWgII/7rwhNlPQrusUx765CRVk6e2elCKz/DFAZRwvFVb
qYQUtuPswS6qu8swt6T1vujLcpFmRWdaAtjeM04YPf6lAG6u+4zXGT09PTWjQd8ATEAmbjdRdqcm
NZS08XcLVAV+vN2NbQeqTpvEO3SoY4UTYkoB9/vT3kNeQ6FQAHqjcHtSob7x7FBf+A7o57SyUbLd
dZrM6zPg+zjZxDcvXAOpxJVYi7f8oCE0nWgpFDZ/ApvVJBYX1cljhzP2MW4I+DVhQuMk/cAYPVBF
r4LBQMbLZaLUYxfBPZwO7khZi0rCJ+FzyQHQOK7rMaLM+DxaFifT94oq8J4MExd/OMYmPftMQJ8Z
GVzBfVofNs746vRwQBdZaZBefFKsI0v8s+50fjqys8tOg1/0wQRPiwLkDirD1bTgl3uvcTGrRr/G
3jAoAmPCRBmcfMNOkQmTdXuTsxfHp7sTNWG/hOYpDqkPTkQknxXXYbSlkWn4+1E/rc3Eqj2mozXk
kTjT92bYMoMrsPpOKIPGhcrpjG/POe4hpQ6vQKXzcT7hAte7b1GZU3zRxt7q7pAxxZMron7Ve3ob
7ixQiaf+D5lSBaZP2s9s3z/CCVJHhr8lh8CM+cBKvMJkvi9nDIdi+YbPz2w3SOrLBTu0JTgBamu5
TM4n5qw9SkFoRT9n/RUmlOGQMV/5gJZFqt1MURFNnRQXmvWXO5VA3fneqvzz/tKR56kzlTXQyMpv
C7dhv00RlN9miQaYMr0PkD49P8hrM1htUQh3bn7HW7GwS7AksqIbv7vWfGUIVQJMGEyJ8/iDcYPS
cqa+P2dQLjCvVsqH8s/ytlC1GtlQGR0wt90iBv0vDxF7Pnk5Hq6gtRW6ERzVyMw/McDxPfNDziIg
FKXixA4cdEXn+Q6N8qT8AARniyMSMEDPK1jqhSmeGIyA+OQyWtaataOxYlNEC0pp1eGTrdiLszsm
seIdOnNFOR7hIXIIyQyp+DXOhNiH6PEPVwJGh8+HmPC3Nb3aaiFLpCtMTlyIDNS9O+JcjqC/riuP
Prr8zZelvK/SRktHMFaazx3wlYZ097hnaOdRXA19+RsFsgIPG/NcV+5OAdu/YK5P/VeI18RMygcy
t9XXlXABv8BedfQY3tfKUpm3XtPRFAazm4qwiMBiHyrL5+okTdoDzZMNg98Nvk29HAnwscBwSZXf
fP+r4t3HSRdMQEJeAZCDZCqoA1Gkc4ECOITTl6rVnd9AmIOi+UC+9jMdVkLzo+IOK85QJ9QRmR2n
iPvm7VBnsrmZ4gFKsEPH7xPEePOjpmfbxDF04weXqZga8nFx1GhIzzuOQmUcyXJzfYv9ozDKstfX
Hoxk1J/fOAwDq5zNvW/Sa7/54HFASjTXQqKXXnPlDDo+CTSUFgAoZumqbtL6WZmvqhKOaPTnl/dB
Bm9e3byocoWEQw0unErHjv1rF7VrWIbqV3EtkcKCoahGE0CEOzOz9YHYhota4dPfMMbMoystpdte
ayi4HwzMOy/GFV2iH89We9a09IPt0vL+2MYXCJoJ6KHAdEXRgCAp6STTk0DuoGJZpkEh+8EOo2Gf
aMXSsrPd2i4zxgWwd3qhpEb4osXKAfxY2jdWOJBrii8Di4Z5BjMSfCU9CkNWRpAWRdWOhUxE5/qa
oSxBNvGASy+eQJtBZDLOidRG0K+16oBpC+9v+xz2pMMGozMilWn2RT4+MnogXi7tGGBa9A2VqF3f
L5u7ZdzHp3bbvYKOMW2oCVpcVadngk4hi3H93e4mYZVtYB3hAZsPf5rUZhlrfv3Oae9TnIUSZ/wO
zvDn6IZu3G+RIx2Bpo3WS54Co7scmkWqBdJEe01MHOYZv4bifZ2OggkrgINmI/56gyIpTfUHt//j
/R2rvF1Cngz8fQVQN/pv984+jwR/X28VcoC6KYJlSP+Ise1N0Yn8UwcQxZs5rOCWDXX1E/X+ejtF
QPciVUzHoRDccVteqdDGzmSUycmG3Ho10cAii3CiPmzbGyBp/cylPl8dUlnbry4bjGc5ttLm3d3Q
6yOR+pKVer7Xtp+fLxonKUV1dde/aYJPBt1oloCqVOdrtvfk9XiWrx95H86YJW6CRI3b117CLxUe
H3f3sOZrsy5dXqnY3a0ZDZ6BrG8dgnLEW7EC194kS3kOpDpL77FOUxEdEvgsNQnnA6wbHEpzqEDR
Yu4EMCV+QIQggNB8GGtujDsr1cSvhHmjdC9yl393Qi68oqf+T0nZM5MfxgtlXOjaWVPL/eYPQTAo
WLl3INRvGCdeVnzIzuG3067nLLE/Rp6CHaQRqfcWNoEh/5ZwKRqGMca6g7lhFtXUF14EQSaJrSDn
e9BIXtFat3QPs69GXA+ctTBYjED3DvH2efRmj341lO/pfz9/eX4x1qg2oQTidf7c5FSvXMlEmlmb
fbNGR9hKB0UycjiCsSEVX/RU2Keo1kF2HfQP42hgGASGI0tJ8SLE9IfjJ2t1cYJKSlh4zwh6z8Hm
G2NtW5Gvz3P/6Cw0QUFXYk95zHi5Xgu9DseJDkSlNCF1mqUOn3FbFjT4BcOvQfHn6weLr6cap3rW
FVhl/oqK+SkP8VY/vYFBZM1RgpUQRu8ulJeNl6eTROCrtaiKydOVjpatXtd6nYZjqrJ0Cs3k6LLF
fUDgXgmsjnMS07ZSsdUZulOAVotD136kLMDP3g3UVrtYYIHH8q3ZPotDkt4BF3COsajxkxW6ecgH
DEJr3kLhJm6bGgazNJFKXuf9SweN4YXGSxSse1j5n9I+BnFR2MidK9gEFGXNem+moxDDY+tGfeVE
Y1c1mVBDTrZQJJchOWIe+RMq4sVP6kkoaUK9MS1Bk8tAwbSIlyspSr7sMQSNuvuFWEf9ER4a6AJK
qMSf3S8sl2qx9U8uVzmaoKVbcVR8m50mtNGEMtW7fXfgSwleCnc0OcvA0pvDJ6ur+peMAS82/avh
O0sY/DUJkRaPVTtuK3Hv5hElDzM5lIDTtNjexCo4ciCTvoXy/Ekj9Wsp8Vi+Amwg80Y3QtVpPQUY
nyWeCGpWuoW0hX4JYG/RPF3WU0WVwHU7cPOgnh/KqwTPWbUHwx7+jkCIVmQieaa4HEpD+oheGbL3
G4KUYX30QrMY+WhZFy+SUSB8C+QQYYYfFvRkGNF8ouHvjpxkKWTBh61tHKI/wmHHAjquH0FUr7Ag
gDt4aMmJGtYbUkt67LygTMnMs7fuOvuB5WIdEf2g5DpaPtnCM3P2V1dc0k/O4HdZZsV8pYXqrMQ2
6F3xxdsNx8T4dD8zf4V7GPjYsJstXtfr0x+Pu8yPWTNd3nZpr6APwD5TSVLRqbt9ZopUYljxzAfa
8UdymY+fTl6N0w2U2LZO7hZjEkv67cFSEudGAeSyLOL63C6naGyoMur807QGOsxZvPE//FuaMl7t
6AOcwfVlBd9RpHqZEv21W9T8G8/XipcdIUFAtcuPv2Ob0T9XOhgXrO15jGOOzEKjdSEQHavR/RLL
qXzotaVL9hewk8ChyrP56EySCxOLT6dEDfBAFu2zhpnoi9wU/CpIk5m3C+UwnqHppepjh+YkJ5Mu
oEd6W+pDsfU0dGIin6/wSMheu2364XErbt2jExh6vseR6q8Ju/LLQsYQrCSFitvZJ48cq0RhOK5F
6GJbIGsuiaDqRrl0KBRVmOLbGE0Xtc+JfZCHbLBIZ+Am5mFHjAaZEbU/ncUjfFXtExJoSQPWwoir
3KKKH1xdw5oILfQ3G9NDxt/dXFwNqvlJICk+Eir97uIxiu/7K19NHTYv1RVU8ZSWVhk8J3og55s+
/NsZ42e6RmSaxJF8sPsCI6b2BkUuP8vKPKx4Y6HtYwHpjLNxgX1BDQ/cIpY8MjM9V/1E39guw/n2
n2ZPUYtS4CtTf4DGtswGllXjun8N0rzwG832MLq3ajNv+P0yWD/RAKbv2oufgidJVjDDq/1rj31f
YHRCxJRjctpo+EqIXWDG/XghQhkQ4B61IaSI0tiP+9aDAOcqx2y1H0gx/+SbSXvdi0QLujW7oM8o
nYxXib8p27UQIx6ocLd/aei2oB+jLdNyeHhmwwh1joX39lTd7Y4wSiPZAVz8/L0HwPsI+ceQsLSR
o16isAxCcjT0PwvMnBa2FwtJNiHREFF+aUpC6yfNye5/sx7NTEyCNSfJ10uk8MDkPqGBbHS7XddT
Da2s++Lo9GJKFIUOQg6vQQoGIYDZeQE+ZEcrzafTPAqUE8uk2TnZE0TosVzJeDMSo6IFMdBVeV1n
eVeHp1/P31Ap3mmohAp1OlaEFNYwEn5ZUO3UzZshBAHSFIHCaDlnDuBYJLDHGK7rU9Uv33/Fy/bo
BFwQ6yGKVO61pod1BqgeG7PYILKqHi81Zmk1gMUuNd4ZaSvQN/4iMWkYMp0l4utlbepvC5cvqNu2
bzINcKDHMwFnHl3KPJe5m5QvJJDqKqm4ZwEbTEJNo022I9nRV/qwz5Ulgw1KC+FOLY82p8Oyd0We
QI/Gr4Az4rGXVffyRjcYA09d+g8AkT7sc4aPyGe9JI99DfI8dwAOnlpAS6HK2FO6i/8/sKA1V17n
EICauQK0ca4RYS2eL5g1iTohHUo3wfrIZzDADzXJsF4tlbgYvGQMqixJpcaSaXZyyPlrvaNIbgqN
klvcYqooe8ZORW+X40D7gvheIcS9KGBrUWYF/cbBWBhwtKUnRrxF/bi8kOsiynDU+lFK+7sXfPxU
GtK0LIPcT1zC7X4pN7gur7C0WipiKJJehLiIpgvvhtyDq+9ITYOggogTSu2e4B9rTkJpFhY72BUb
1pblI6JQlEU5HodgE/fxXhDqTBWmJfm0m06uwTujJY/+sMfG9RUpDiEjghbIou5zJtNZhI0Rnir2
Llwk3moz5tF3qVjH7xi6V4vkELavfJSTbgvboIH7WjaLf5Bj+8bk+o1bwrlI4AzHPDAbOHkwPz1w
V4DBCO5i+s9j1LQI03d4R8ywvR5E9KuqnvaLjInQChD29aZ/1neZFaWQmH3cojf5mlMUMMMEKznw
+jueMwq2lU8XrncysPWC4LpQK5XvUdo3Ws+UV9mh3B2vFJyYdZk1hUzrHPpcc4NQ81CfjacZK6s9
CgNQCW/K9VFAVLhet9CSCHMj9cVklH3qUIjEg3BEshRMFvonBHqh9mt0eYznVGEkQceWgwTAG3PG
wlQAAvBrzuXdgXgCKStHobf1Z0z5IwLnRmv15Kgt65tDF6QoIFvG0QObSqqQu2h72F+Yf8f/wVIN
W+nGCOsJ5LpyAx3OwQ3Ae7LtaCtDlyi0KkzM89Yojq/Sjvfjgw1qpeKmrB99IUaVxB5moQ3HCb9g
VLGLoDG1PkvZIT1GE8T/oWHGLl32qAHzBIBo5ZwrWl/EuPWciN3Arr/9/CKgUrRb77s5juxukx45
rZSPvAiqfYIOS0HXZjHRsujhXsXEuJhMHngAIHfK3wpdQYOaD/1rS0oeum4AMwsVKu5xwleXHnoe
g+eDLpyJXHus28Kukbmm8OXE8Z0Nm3am2JEpCDbILGIBKYvQII4YacvG6tC7fqmCPOV5Vs3sIqPo
PkIR/ta6Gk7ZpndT94VpDrKb+/ZWzgcEMaSgHnJyC8ZBa9sr4TdDjIjE08q9u5d33ae4R2RXctEi
cCAUwTj13+v+vTGLCztibTTc6/p3IyHC1pW6lorQm0ybLfkewabEOOFEjwTYqEZkcUvQqSCuSKYa
D9knOHbf5c8BLJ5iZ1NrTiXXVoigiDVjMTtrnyDJXWdORW4KVi3ksqFrZQKNnqtIpWag9gh5ibQU
XmY3wo1/VXLzTd93w0RU6pYgpueA4NtvKfNpqkyGIvLihI726bzl0e0OJs1WltX6TzUoaDxzM5Fa
SV9m6336M8shk/A1YuhQpSM1gaMKoGa71ZKB7Fl2agIWGWK1Q3kMT6q1pkOCtx9xfLQJS6/i2xvd
0ZQkH02wLJ4nbgusKKwdQ3IgBMgE5hnHYBCdtmys/XDm7yhO9WkK2yDjhgDTdCr1NAv4gl6qC7FY
wYejHmPs1i8fSZ19qiOlZ48QYRAfGz/p+2po/x45dQXeeAW/WboNE/nUkhh3p/3RrM+O5s6Ps4bA
9m1ObTWBy8HfUSaendlP9N9jXfpFIBzF1qLSSGSo/nsUnKsg4Ujm49ee1Gdz+5WGIJ9opb6CClae
pA/YweDWnp4rN6SJV1VDYyyOjvWBaB6s5TBaxK8KAsvMk83lEm+eB0d/QKKqJOACfQwe2V+J1WpU
SuiCZvtDoiqoEgU4csVpS7Kk1w0Bo71r4a9/874jIKrgXJbmCnQ9c3m4ReYHt2mrPz+MfMQjozyL
kziIk1DBTP2RSwWOwc0A0umXTO/eCRlmhW3MHwmyKpcAbzCPs/mlDRoy1B2NS7p1f80/qJypx3Wx
2YEgggJid5RLQ2w3KepYy1FIoWApiWMLH7zuFY2kKxeVaNodjQU1mfbeKxrNzs0mJUIMpJwZDRC9
aVNbS2cMBLql+LSkb/4tf03/U7qJquWw/tsgJf5Fdn5d145JhtxbFbccad2cl6DH8jbXahH21NUx
00k+lCVxDXWBdf3Hc8O2wYsAPjHaQs6aQ46pDZbEtoMtzgFdnhCtLRpIu3iZnIV4lqpAuJEmjeqT
G4ZigEIjPbDFsysm3+a5O5YvOfxbWpJCUkESwzMvkDKSv0wsP7cGhxsiFHrF665i25lcFP28+6zn
0rDtkqHTqqbX/iyHFYl2VAXDgR4BPPMu3WU2v0LRTsY/sqyTdk1YLcTpg0XjS4OvgPksmFBjylC5
Eq/x9BD9GjaAvXbSTZUE8LbtMmSPlktMLjTUNaZdBPWgEUCVfED8Ojf81IGz5OXCT20t1m/a3Iis
YZEdYXo+LIS/B4vp/FMPejhOmY63V2Pq1YyTKe9/rwalM/uzibDYUN+uJhSw4pYN6UKjmc0xy17q
+f98D8FTLDXIS5wXt9PCPQAdOACyl3D8JVa3gzJvDK7tTRfNy/3lc9IEgD8bur2dTLR9BBeKvSwS
wZqqCTgJhqZ/9e9P6usnHFiJux4+0Pqjcm2Nz0ibFHKJe5j+leS1ZS4Xcm8yg+A8gh9OIQrcHEvU
GowqCycyGLK2DcRhV8ovC5VX5AmlzEsJOfEAQi7nftiOiMETeseudPq2QtDGqhRBmXxBWScXaDOs
zCOyjGo/eON1jCSTRQHuToiF1ePKtHyB1QgOjjuQPe1dOsbJHVH/mxEciq/NwyfKH+Vk4nxm6fxE
yXDKGvXKqva4jKi3GrDl5kEryqTsB1Szy7+/fCC79DPbfq44qXubw01/PDqGONGoZaMn13wjfzZp
Mmdpvg1BkQ2RSNWdOBSgwkz2a2D+UOUQYxXgEWJzsSUubDAvd0pmz5qG2HtUcSpiuc4pbMo4qIDW
T6Ma59oGDomsOEuZ/K24wshM8EjKwRsWfJFw44Itqxoku5j+jh7FW/etWBqTcQop3+vkgOMNXbVj
VsJiaZv1FcFTC53psCMPwmJ9NWg4MnekPLrPr/E4fUZ4H8q4emEMN3PgU4zITRq5+wCEkTuuJZF0
DhXqZpxcOX4zK0+hLPNRr3/dCs2yLowBxZb1tyUd/ieQ9V203OwU6lBksOP9aK4Xrg1eAdrw9JJ2
/fd8nw5R/wWMlnX8xTh4IPPe7azF16fY/HMM4AkaDj/EQb75P/5Yi3W1dsPwpxnBd6b+pakZfIi5
BwtN1S8zt5W0CJk3yXwYUtXpVHNpsLZbFG0Ok4oPUG+Ra0rf7KwNKCnFN08JqM1XqA8rLuN1xDy9
Huo1Q4L0CQGM8P6R1CMibVwJ2TPnxEJH2TXkDlNUDeRDGLpngcdfNI5f9nbBR3+hVPsADOB5i70Y
KEdDHXayTdmYiBSXlswlXmowsXVeiAwNUK3GDjHCJIFBQYgplUYyDDJ0Y5B3ZumcEB2sAjJ9Ppmz
7kPueICvmtTdBMDEM4f1NHIhBmYF28Ih86zc28JF6iIdTTSBVwrX1Ipm8Yq8974RkKVtPjM0XXis
/67PBRj41q1U0BWoxXIKQuVI17QgVeq4pp30MQsW0tlQd23wqjU1PBt5vE9tZPNnu0EPrvXLHSna
omfnWjis31N69ANNvCzUuuX52KQxg36WUsSwAigqaEUozHVqbd0n1TEa4W9vrw3MpErLgIVTLcQo
DAXPMcEDj3rXO7+ldcWG1jfK2NwtF8boYXhExx/QW9L8NIxeJJoDbxFSCtwu1kA+HnKwuj5qIsKe
BHhPXSzE2YNIlwHhdZIAJEZKszsplhGv8Tisy/AcRQVluRl5I9jNyWpHMv08Rlhno8/9fMOcY7Ii
ny1RRQxZulaYJiw7p8z0g6RMJKnoDc9g/Ux32PXytRj1QQGj5a4b6HOIb3Sxg7Md3AB22sjCc1wH
5MlB4W1piFR6OVm5fNv3RgSUvUiIcL3kI9sOC0xkx90vK5E8nhFE6h1OYJeTZ7TNy3rsvlk5SWkC
Xs6LKXESJNlsTI0PgejjqVx+FBUB9co0CON+qQZwoJp5PcurrZz2APl5VjeWiHbY5Sf/s0ZsiQ8w
mCJPFpYyxW8RXf2WMSkDxjCVTGJM54XSjbpoBRv5CAotVv8UHnOeqMdMujl6TQN6a2s1xbo3qQA7
+8iFIv3mMT+FgI9+u5eRMm3qX/5MgkoAoq1CPa9ze1kgTgc3WV5ORANpdOFJCokyNiJVXQWwP5cj
qZc6ngFjvDUMRO8x0+DS/NPh0z2RBYgVlvquSEV/LkcXv+MWCMDZPeEqXRRwRVZpMU/qBCkW+3bi
04uJUhuHUVI9u7r7QGCe0aCUosmeGxhcTRKF7lnQIe3EZhBp5boqsDXrjtmhj3nr3nPirxv8wPBs
EX2Lz5phmSMGf9SzhbcpMGGmJ/yxDmodx5jIKgmuZdIIoOIEcruoFr5wAcQNPJ6pWLAaPRhc5Eq0
X4oOiqIY8+6TAR2pJGiWX83W6f6VpK3ZwYHEEi5f+IPecntFbHRmVCKvDyy/jX3GW0+Qoa3BlDlF
rFu3yIKNPWuXRk7ax9rCjHd9IC46lcP83xTPGHaWNb4Q7Mr5isLDg9GyHAGqH+n55ppNUFnVphZF
Mz/5Zq4/4ef6eiQHyODbTKOuIozU9gb6gmEbapnzdPdNGn6+5bka3FdAl0cP/H869AUuoHbfKEdY
Gl4QSuUYV3f5ERS96jIPJNafs/LVJWsMM41+KFnNRNK0BfEBXeeMwAWO+o8UoTxwt4eKN28dJVpo
u105KyKOdDY4DmjJP7yNlRnOu90HhevmZqdK9bTAS/kNdHlV+44NR7XImv7+CJRj99CcMboAO2aZ
bgD4ihzIZS1JS2aBm0zUyUHqi22a2/LDIsKjVi4kiwhjlAFa/E6X4sqLhgc8jXseZqMR3C6uGQ1o
RuQMsSWUuFd/IVOtxvHx7M703gEH3bbVbb7GKBdmQh0CmFBCqZNkDtkLL/qzM2oluJv8emuqqImg
yYSg/Bjo1wvGA8+WQIymWHt9dktXrBkQDe6daPzoZf7TfCnyu+H7C8TORjhPwS/CYF1hBfBm5adY
HFqouxGLFkmZ6zXTYY0QKgpovUKB91e3bfXYvYX1WfUa/ISsndyTNqaT67DvmzAcWd30W/Gc0inq
vjc2zzPyJ4ljvTKPmplMt954OjnE3ES4+sRCRSe/gQRwaG5+iBqbMRv5Wbz44F8KOhUdgoFlqL/D
pfemvd10JphIL0Oe5Z6trTuUGF81bYwBuldNg81rqsPxgKLORtvCp+5WfMJkgyfQK/xOr6LgD5RB
a/IkmIecZ4qA0TMLa1EQHNasXuXhDR6bq2ho6ZJAy/PV9txthGyKME/AsHDNep0xnm2suuJ9gBcy
qYEGdUkINNQ/W41zX6SZJMlFEtZSvTaqMlvb/jkPCFZwXrE7LMRTiSDPq7WFZhQ3tXJezAPkwZ6M
kXBrugvQAkE39ItieEU3uFuo4DY+OXgveNBah6dOlfeDn3uldA0ddMkdJfTISJiEWTgPYKjiGNfJ
PJyXvwsXbJOpQ6//QoJpd+MqQcQz5VwTpMshObt9a872MqHAvjiSj9Cwg2JiWnm2WtkhbsB07clU
lNGCpi7smUyG6YJvZ5g43wyAXiSe3dJ28G7cMPeEF+yux8JLdkCv2Kjr088XcGPyA8GdryGMpzmX
lMnaXGOxYBITIGA7GUNFZjRYXxCaOVaa5sR4P2gkmxNTQeovZ6noj5sP0rBXm/SEXE7dcKdwpujA
BWAk6Y+r8WZmZTkVRMk3p+EnzNiKkFddWUoIXO+nQqh1sdAiADMTRVP0hwVMz38kz9nVhjXnbdle
ify0ct0VRXtgA2oMeMtzHrm54R0u9jUE378+Y1DfK+Inl/Zz3pJLygzIWN4o3foA1x/lfgWIzvKU
bdP+RcuT9dgS8/ZF6PdHZCIbnGYe7MV+G4GS1ZmBwiqrqpjnKUmy4tVvv4BuGDl9RSqerxMMkSRo
rLu2AnZfFWkyHHEhZPB2gxZDWImGxsGe8R+gIzG4X0tycqZbmBeGrtrDOFvsNXHVZ4tJ0SHdgm3c
dB4BdG2wnpmdmresuk1I+l7G46l5acoYMYN21H9MJlHmqfMY0rT93E02QvneCplLCHD2n59WHE9K
zzPn116gUZ5mWXfthALO0jFbRhUhsswOk7UplZsALBi7DH1vSNw+NnKgeh4IZOGRmGX/JQQK7izo
2HD97183gZwabJ1p9OrlLAXzv+089JoHfmXZaMjDA+Z7KzXdcOOpH9dhdwtIHh5ESV22ESbtn0lR
miA+dryzKLBOieayHl2Gvpmxyrm7aG31zSX55QQp8KgzxntedgCVJSdbgV/6M8H2QCjXyA6B/WVJ
iTvv8CaEOt8d597Sh7ntp63IEvSI35liJHS8W7c35sTgea80qEP65qK7hOSxwWm3TyJZ1m8TiZ8t
o+rMijrsp+4pYpvXaeBPL8VnGU/dZCyGqyN48o58VGJPMwvM2cc0Mt4CfQWENw2oslL1BBSkzmMz
B1d4idJv5R25G97u2nDkVxl/Q133GktUG4jZvmJrQ2n7cXTRdpLnEoOrznbERXtg7zJXoFwiKgso
EbsSZ0I2CKoh0pvlvtxmcpnroI5a4uTIhe7PY21jBTZKEJU406yt894UOBhA2oq+5g/WtyNQHeUw
cUcK0YEr99DR3cakXeSvvhmZrj7RuKsNiS140549CCeb6iozJC8wAAL5JnklWwJmHa/HZfW5326x
YdSasFgA1jjyiD+5l25MoKKzUryeE6oGVNAavMZ9RMhG93lkS36Jn6W54wLARp2tU3oDG5cTDTnR
uQJVe44KNThd7oNBWQIuUXWf/e8oZT6UJ5Wa/wi7iAmz2Ge8Zoe/m/+x+OinLvOG1++Ni6AYF0wN
9QBapP3PZnP6MNBf0XqzHiRQEu20Fp+9kL9vsBXQfsaeYiNYjTQdIEiDI6ywwrtpLFn45OFN4PpQ
e51VNPHRexO6NbLLOM9KC3tHtjT+5RND40sWXcIVeRC/rQZufSHayOr0hoQw+33xoKyJQKiHey0l
tJWj/dZRC0WYDDI5ho+EoIa3/Gtuhx3YY3f+0465ACUHt+VGfUnbpvHGgdPgFPBwIrzpxlamNy05
/bDxN3DEBQAjIhCVCSKXotB0vwWa3QdQoX4gXFxSZ+u54mX+Ejij83YJTDx4wUbK8JgkY0eIFz9m
aibDGfQimONx/+i+PszWwAX7O88HYDhHBHnDoqt2w5gxXB5pjP0DUI7TLJ7/yI4c5m/r32HTgP1e
GrOfzpMMqbFuZamS6AQMRkyCrkjeewSI386N8i5W5O9t4Lc67K2JBcHFFXZDibCbDuNTIT/BuXB5
8CdWBjE5F1ltXGkP0tZAUN4e2dH78uBReGCR6FjCgVq/3B8IEFGUoUT8Ratr48TPPrQdAQ9MQMoi
2Vz9Dd2iO4aS8cSmMSEoR8/drxQ+Gn/hLFLiIM/0S+KZCGD5BYPv4LYSNl3/9WuaJEWXJaoRn06c
yrPo6BkSmAeK9a1SAVIrPQPGioVkIi/3y/hZCIAgZ2DHecqB3V60buc2t/uALUAqriJEIhSAWqmU
bgNSY7aBXeSj5Jsb4K7DrVM/PA/LyFYS/QX+XuJImo6Ni75LziePOMN7i6u6Zov4zEgLDXvrZeCt
g6KbYkN0fC9U38cGbXI6VP6H2OD4DkVUApioA7ZlvHT0Nv02GdFuOVq/NPAxLCL72Vm+p79T27xu
7ZIKRK1iY0bI2UyWi7mNR547gDMHyQvs+v2UBs92xq3hYuL7hVNbMxxkcm0MYVJZvjJcPfDGtZmJ
Y9Q8cd/g3rlx+czhFRzyB7zB4E0vPe/fiU6Ulwob3QLD+0QOqf0HCxz1WqTnLsOzmQZp5jq2rqqX
9gxH5aSUHrvmb2q/w7Yj0WUoeDEhU1+lyFySkgKTrSQJf8zRuGWrA02d4SgSk7OiDAkWwTFfVCxH
6zB9C+XKn1q30HmThzy9+yg2bC1wndYl5KwnMnDeAjlPj62NxReijNkuRcqpB+6d4i2cZ6wP+vR/
SlFNh82ejvE5EWCNJD6bYLZMkopkRpbnojsqxArAzX/lHKtaypU2P7pbJH50pSZ+xBiXyI3H/DMs
nSIZqOWUij8ePGUmb8n8rhkyXu10kiprwvFGGFXGKcuqL7p0EJ5QsLqUKAY2MFN1S34D6k0TDS74
9VDNq+1cWezRxrUvtD38N6XUOECRlu1WmGxFxn2ZAsBeg78nMN1et4MezTU6pgwcLbh6hvr3qoJ9
jFkg0VXFd8G/NLEEwvVIYZnzhFIE0ULtgrfhZQz2wlrc3R7qD6CT3HmhBqpdhnstHIWktLmjkBE1
q3XIiSTVgJU4PEfvR5xNlVUFN+Ajc05a0bcIUP4ECrpBEFtj2tWBHpCH+CbQMousOFJzNHVOnwEH
7JNkWciifBIgq8A+iscspndwuU0fCHFVOPUb6bNhaqx9C/O/VvZdTIuAoVSntM7k+dSZ2kgS+Olw
QlvocKUs59BGRKvAyaNONC6YnH1g23UGGk/txzQPdze4CFUfFR8chb9Lc8S+gozaQhDpBrLeFWox
rjydP/9IENWmeQUWjcrxAdTVl1IZbzbl53s8T+zIMIDUdX18lWBaVe854tl1k12r9YW4LXSvkuw2
nw7+JMM0PZLRG24pZFLCZuGClNDPik2C8aZflonfX/MU7zRkKLyQuWGIPhsP330vr18XFfm1J5OV
Sg4JV9YOkk3EPbYLPyHHX7oOOf6TPwY+t15UFGMKmnVwlJUAv4JdUd7YLfuBw5c4tXcWLSNjLddO
0XqKH2he7f6yVm5BnjpKUsV0HUfwUxYYVHL96stI43MGGla3Xs5Fvim5QHN/2Vh1e+FXNTi2CFhe
JHnO4I9O9cyfR7A0UXuJkCp+Ll44Lj5LeCKQAGh/AXClxbHX/kAs70c2yt2VwXk33nSxLYwawx3K
9P0TSOJ9NUfqRedV+TrQjmh/4pu2zK560QOkr3ULe3iT0C2HmDxiuHH3YqktCg59fpx2PxD5vld4
d9aPUKXhr3/vQiRJ/uH3kddL4Bz5qROnp1AZ+dMx0qOO06BpB9S2cq6cDID5vOAGy+RZ4S321m5X
ORVJdFKb+Y9P7rcY0x3pAABahMqN+WxJC409wDPUVWklCeyTYo1voRbRYbMEiQ/eQYmfZgsVsOBM
8Z8HPtuBD3i0ZQyDV7oU1VIV/I0xVz0dwR5X8Bgspyxu+ppnEc2a4xyOiA4lNhBHifM8/Iv0h0w8
bUvtbJasNmU1Vi0veN6lKAxFz2pUkPVhgjw/WMgEEun/UQVDYhi3abWn3NZbBPdGXCsUG6OKUjL0
KNEMYIewcPPB/WGjTncMOrcDwCuHh3QJhpmIX5wRxhkk8+OV3zGJv3yfRDgf/45MJpX2+s3uUjTK
+bYZnwIRXGnXyBxkde8AcssvR6yF1fIw42wsIcF99octz4tTqv4byg6h4SnUxzhptV03nZ1CYSnj
imjBsK3pVykhSOgemynt1AI+TeMY1ol28EBJttRslvpSzeFvnoGF5TxznFQbdvFfjo0QgVjPgS7f
O9OsMz7mY2jMZpipKz3cIubuSWcCrTjXkpXCJcFx1A8PqI6PODfK0q1QWC2gKv8UpEo6xqgcm1jr
oYcdLCw84xnT3oIfJFz+C+y9vHrQjUq+zAG9lkWjgNrLqtsIaowppPmcg1kuUYKqfrq8LpdnVZ25
X/Jiv2JNh+7KKaq0ZyBVQpOWjdmxYsNwTeMqNzoeR8aMcsQbfLA6jSWsL1Rrpv7l+rCw/W0VNybu
oYqoWKcesByWHCEVGkkweMOTbZhy1542VwPfzSu37PN50kD0c5FWWjiWb9pxRuRk3+XL1YRHmcSH
1QgVaEGl6gWeJcStihe5Refanv83YRe9V8OBjGKeV2bE0IZfW6TERI1RSg64Gbt0VeEyGO1/wXEC
qwcYsD5/VtU7dgL/u8gUSP1m6cRA5Jj7lbeNrCDW0kZFPJ3nJ+GUiS+GDS9sxGL939fNPF4CBchu
V+ZVnOo7aPSEYUbpTIZdx0UQyTYj1UrO/So032yDymE8Sf8+LAkdTxCJ0W3rw4WTkOJmF0ihJVAE
8WhG7dv0T0kfanmBWk48SWlBG6ZFKJxDzx/93Itsknub816dqXVwqTfGA5QG8UDF6Xdk9AyMNwUC
L2xLXyFhj4UJt2ZAGgvjMAmDkqd9RoHF5tocIqKeFFilikShinVu+5W9XiDSUh8248eCKt3gfuwa
QvUmVWw/i3oRNbpM9E+1XdIsnl+iW0VWvdVTEE+KOaAemHNPmk82Vnz0HT2r0qWt7P0T50+EE9jo
TMir88Q8+SW9KpL/JQzhfJUorJw9PzynGwZqPEY1r94Flpx7PQsosLVQmQPbrsf1val9q84hClwh
ilRiwMn26HVvl/akNiw3OxP/zwLjYllBjUD0rWSiET4xqlh0EjSL1tlRUm3ULk984JyMZPFPbTIG
mu+bsYU9hdtq2xcp4TPQqIaBaeOR8K9NB4IEv5Ir0yiLBQRIGowBkCLoB+iSUkuajdJwU9kwBva7
l6lm1mOfSRRpGuUtPe0QdY6a8i/bXo36xXvlgpqtxrMTd7JhDtaVAvbGfREfB0UvoSgpOjLMC0Mo
K15IjkAbV7fsBfsP0WmPb9dsSoqed+QCh4JKOmkyl4SBp0dxzVAuRx0rc+HLboylKlScU2u4zSQu
0V6ApnBRJasHeRq/D1EfBWTw7i6x1SkL+SZ0OEoGni/FYLj8xARoo/+qrnWSBb6LE2D+9TmqSf+O
FdaG7CcScU09BOPfCC8rslTYNUX+j/l8icSzKfCYxpsm/Nz+q6JNNaJiOiKu/2X2a/NhpTsaLwav
EHWRKX8xi12miRiqgke6u3P86xwbj/tYjrg4Lug2cNFY26ShtEqhsjrapXzc8C7CaZBtgbO5NUby
rzTVSte25rVieRS6/mfLDJTOMIGrBVk/LR/L55vdM+gAKZ6VYnDtphT+KJFr80tId97zYbh2lBXD
6oIMsi13h2l86pE484kad02dJl7DjpekMoOdwjDy7utgPeZ4O7k4ZjsUxBzIzgMwyLhyCPK73Pzr
CNWFeH/0MAg0PPlRjIhFsNI4P29GTbq/rSDS3J7tYCFLFroJ62YQrQi+fcyBHKU26UkmjZ3mbAnT
5BCkh8hS/Vre7dNjjTUhta8I3RXRGBj2/q0PzFKSxuaPMnkx4rCyJ58L5oYS4id6gprHh+zCmlVR
5SkVnD8j7XbW6S3gw1/HhQNyQxQGeh3dAZiAvS1re067iufomQNMemv2VN6d/IqQIKz1WJbKC4La
OpMaTugLNMkowkFvo8dn7N4iteyodRBOn93bLR+HU2pSRRa9pWUN8acVYGgYxRsZS0yg+rgM5cqX
74CO5jZkj2HyegbNDujLFFTz5ZnAReApEYBJwq7NkpzhcvuIGQQ2zCRP4WwjfuX34dB7N7q2GX9K
xUdL/G53gZv/Tqn7P/BuO/zim2zN/xYheRu/IPkXmpl6ubHMO9sBfcyW0wwBwEeadEb/5uJXLRJN
+NNZEE4QdOVReGjMk0uYAK+kaKAHGSKhE8pcbLBEHQFuN3L47qOKwkS8OVlEuWqT0Segiqos1vug
DgMTgLpWqvvVFI9HBOXtm8kf8U80wTnEpxb7LMhdPVfRmDlt6QM1cI2uV/gjPVxWpRduXqaWsI2E
0/EJqPQ91HWH0o/DEa3jCs+8YSdfrufBjYf9oGEA5sj3lnlwdjoAbgbhklCpR09vicqdiEMiKZMK
WvHE6luvgtG3+uSF9lclwhy6HJ8lkUDXE1854+oHiU8c++vkmJXA7BzBmvVls+k4Nf/R/ZcJM06w
onbY6v505Qwvy4yt88kEsuBMBf+Qv9YUSCgivQYHOj+AtkljFftBgEXQcovQZuaFl79BzVkjOL3B
s+25EHY7FwPbZ5aU0fKv8Dzsks1+hWRUzqAz47x3AG5z/adL60fskrYze7OURl4owq0PRXYx5H9I
UU33wgwDke5bD8YG+W0gAQDNHMkA2AMMSDoZlbCxerfoCrL2c+gP0vpAO+bRCPBZK4TKdi0VvzKq
iuPS9p7duizvksy/yEpm5199YykextkD6l99zNJn/QS7anSajF4VJbfb9pCpdTljZuQg6condiwR
zJ1fpt5NPtnjBUaMIU3hy/zJ8Bvv64NNi6DNG/vu8CtDy2rQCoTtUqg7TVQmSNR3MRWPIhbDuCzk
IgcOfzo89y3ldJMbi1/+vRPifojQ5i6Lanr/2KKIT9n6V7TuwPh0L9U9Y6qwC9v22xLY1Rli23pe
jZeSC5GrMNuVhpOIUPChtgN2uCcnBuntTMohxL+acliIgGwjFtkOgg3bBQKuP/OXrP2jfJq5ZLSn
WWnOZJC3X5Uae7DjehIt9QS1GRsfhMMMYZ1KpFhqLg2e909WblWO2G0bTiH5ZCxZ6ALUpzD6y5GF
+3sN2NAqR15em2tn3inIB7UWS5umgoID40O3jpy+rBlqPWva9VhD1BbOOyn1AhumipvjCYvyoXPn
fjahWL2xqKVCtiP50jtFVIQvpBXMFYdm3m54ER20LhTYlne521TuKrXxK/siDMt79bE9sLehFqkm
imhBlngqbVpya3Tqldi0laPgf2rm+CEddK9y7qyaiUo/pe27zeppacpl8DL8SHuZmcEtX7Y6xbrQ
vtBT6xCsxhYW2GH7j1YsO52Pq4QUaA/r0QTlAeW+BI2+NEhQMes6C2cfb8StAbHXiQ3zNlQWmtI0
0KRTMqEvnd0kEhsqQTSHl23aogj92iWEu4hpzwM1VksYTVb2HX6BAJU511PDfO7a6XYxATNn2weW
Ulba3jVHENa7Vce2fHljuDx6HLJeq3YVWBrjanbQGyKBlZ99acODKc7S3AmZ3vWM0q0lwJ4nOdN5
bCSgSyOwFIPqi59jZ7TPpc+WL7pn0jLstxZB2ZTVR9zQ+CqC+V+L5+DGwrrXcih4nnP7t8l2CH56
ATrytO/i1FrZReOEol87lnT2WsBURoCAaqk70Jh1kgmC8VAGUP8x+TPQpTXSIhetBxFMXt290cU/
G66NWHha4PXplh2LT+bmZ1cZB08qXejLdAtvlOLkXdrcQgvsxcR3/r3njimE83w0ylXLR9phxGSO
+gLdOHzfoBdYd6vtr2hCPKWJT3qJGbieCQwwmHnrnJogxUKcdUU44YL5PhYv09q0MPP9rJcjRhG5
y3E42cmiW0PaiL+BVzLLIGQE8TxcKCo32UD7OekdALgx6M/NJR2XXp7bZP0tvx3lcD0nGrYLYUhj
XrXOP3p0zx4GMLgDObyWbLj73pekkQwFNLL7vPFcWryOwTuNmJDAdkGayGniBckA1KfVNNUjXW9b
16F32BB18jwkKicqbaCIry8LwzHLKmOlgFv9e1DndXuPOvf+O1lY4xY8dGRPO8/Ep1jEllELUBd2
EqYZI3DjqOEFl9ShscO3eceZ7TmrlzRIQFW1MrSAH2KStvHV2Vqm5lbJlcOjsqC5UbMWt4xS9bES
PvIuZ8uWa+YWNKtJZOGSfvU0riOGiPM+8LNNThnFltifYT7+D5+4ekENj+bcawiNDvDh9vW5Xzf8
BCwK4ObhjfUANgk+8kEjqRjv2ODHdubK00OdLNbrFAqXVCjr/+rhqWEYAh9M9T63AodnTba5ayqJ
dIxHkqMNBgWa/mGO5eq9IaTvsve0dzW09yKY0hUddzpUMphz9aWGVBkLfsw7VNf7CRj//LO9nr0u
soqPImJ6j3lJFp+y/m8X9B/5mBBF1bPtK79gwyOuswy8WqxjUwXBpjisM2fNQgM9JnxZR6tdahSr
vSEx3jCpwPQgoUhtqkFNhUAWAhlOt4AzdHcgCey8hbw61BhLcOawT6iB1DgZIxMUz2vXGHckHE4f
Pk46ifUA/Ltm+OOlaa3ZbkyT55tG4aXZBeARKy0/HfIjn9mVfKb9ji6wExZQyl1fwffJX4GYrcuc
1qrUUzVH1SN5NuTyroh97+GVOQ8mRb+607RLQd/TqzK/7T18XYFGHGixy97xOQA1AFWE9/nhyZ9l
grf14poE9yfTJvlp7q9ue+4a3SaeS3+pYByCb76C7VTLgLAVVYa6EJLbQV8LL9gW/FHGo5IX0kqp
c49rDN6SBXcH4T2pc+a3MnQ81Xik81A5hOJZvz3w98clpkMdlnJvtyFYkUGswffRpkJPZQmkqhNF
fCgzdc6RW2s79185BQ3+AT/vVtRMMc9npt73i5ElbHbzEmanKlvr8msUAEuBFXsDEfcqwJ1ljPWF
39IotAWmGeKiZSY20HCHLip/B5XuDIwFQmvzWyqf/aIi1Tfb6HabZCrHTsO499cMAc23LR8+UyO9
B10vwo1aEpo637kuSpo1oU+cXxDglxZ2rOVRKKcE8taajiz6/klN0Jgh2iFIvk70S0i0N5y0ZnSM
af8rWWIAm970OZss1Twkcc5T3/J3KJqXNdBMBMQ8a+/+xS2KPwTgfrXlNsiG/tk5PzMJc8xwMjn+
sbcVBwnpDxE9O+Rt9n3xSMTFfatwN6tf+UKr4h2M4SI6UP29PNWzHHxXVtPgV6VjSF9r1/lYf6Hm
crDw1AsTB51YTI/iBcAnSDRnlupY+D4A9k1OJ9unS7O2A3yFEmvnNLOfK3on7H960E3xTTu2mXxx
SeJXYK/P/0aTaP3guV7LATKIEkHgomSVKc93e8OH9GfSd/Mk36rUa4ckqw4drsTPYiXvuJIszcur
Q76p0X10wU7cjxT4u+3ij2+wld9kEnMCMV7Wy6hpH72+4/L/GA4PaYvrYiwfHdNVCNsKfLpFoI+F
3R/ZcdtOWoF7XMqnQ/XDyirfdlWnkCR73w6exEjTofRbCEUKS3sLtTizEy2Z8W4ZXubhbYSXqGrE
hzZ43OzVI7JiH9EfP/aOfRiCE+LXXNJzBTqCKooHO1JOpCC1CEb9zNPHZVQRhlZMKk8DdWgR1xPq
XrdTfnP5eEUAgPuG3BeGHcwYO/hajeh3QW9drXv+H2I/I8wGA6zauBpRQRaZz3B8NoIqA6QIRu13
3DxiHCAw4QHNn3kBE3d9w7d7dPJvGOlV/NvOhx0YJ3WDTsvWl+EAFFWznmhMHMRNiLKRnXbtE+3G
WAOUtdxzxNIGjVWmXq2UKywMEN8rxwj8rZw3kqSIgU8HWs85V2NLdFA58itTIJIk1S43wKGjt4t5
5BfDDa9m/gXYIE1nxHjb/faYT9G2yxeITZpiqWws7cskKR3F0uQ3gAJdssUraR0ko2xcwSBoVHv+
oa9qJLbH9TtS18z2AuffhDEoPGHhzKwfT8VkGUGkVmUt82Nq+33OEl++358spRFZNqlQIbawbjvV
43eMF4hJrrDSbQXewaQ3bb2TgXA6R2KttZ7x53x5JauYhy5jpvJt54UmJDt141f45Qun/3f1/Fbp
XN9evEat4T1f2CYEgshHBZmPKt0hQkjZLTCdmF/thD0XqnehncGkRudYoYnkqvSFNAOXu4zaxOK6
X6T3j20XpfFxbSD7zVETEKpnsPe1G/55Hu6lskRQGMydxQPdZTY99NIt2PdsMV8rYKAgVq6vD82y
jim4oLAgq5OhOyY7CgPpeBaBk19z0nt2Q2GzUEyLMVm5VPU0hysffsYz49aTcx+LQv2MMNo0l5sv
4L4P4oojG3+QRgYFi6NGSVJzHHokmA4wn/7PMio1ZsbO6KffyuVRFMR7rHFMMBph2ufiB7V/cWcK
V+EQFWeOiVVKWXqQP6D4GoGXWvjU895yyjcSrqbtqzwtFjpq2fEO9iibPbPtpm9JEN/NeXIwhjy+
sa/Kn2G/+pnBpS+M37rIhy/YHPHQSzJBxPXIoB82tYc0Js8HzGXUKNGphabCU18H94Ypx37mHJLz
tf2wV4q+5I7rKwI9om2DQexkGkOgIScIMMea7RXAlJKvGgXX3W28Kiv93xNLyNhsN/BS8k0GuRXM
y9TZB9t9YJnY0eABlA8JonU4bnaXu4yvY+mzT3Gvaz7RVUmO0qpeNR9vj/fAw1RtdLLxagFJsFin
XrVEK+PtiSVf2Aaki2VAWQnLEkse0ZOKEsxXGO5O743/qRRDhv1QXIXZQOH/MB0qiNnrr4MFvtfu
j1+IZo7FlFIXSlmv7ISH1atIy0PS3q4HpLJ5+fG/p+mNiOc4lI4w1v01QE1jxMtksY8g8bcyni9r
pdyTKV7TYKKcvToKLLhH1w54v3BS2eFAzFl6HtEH+ujeaK6TSyGGsU+el4P2E65Pa/gYNedC13/6
8/52c6mF6t8NZHMqQ1hgIV1qQD1aBR9NSwcLu/3DMjXyuxrZ0oOkhrpv/uNyiHZbHTwLj2EbzEXc
EmqGuPt943HYOxJ0JySRWEsV25kYMHjzeMJZ2vLvU+kuhK0OhfBk3LjSc22eIT4BXTZi7Jto9Jj5
bgEZxiS48lossiG6DRTGWQmICCruCX+JzzpKfKuZh9+kqfHWFSS8XrEZx9zmkAAi6Jhk1cNUGscX
86vLPF0Ywo7/RvcFlUAi8a602D0XlQkp/g2Q9QjDbsO+ZpmuZPLW8RalxyTJjAzavvbslQtRdhsu
YcM8O7CfWqypCu4teC9PUhOki+J1DGRsca3LnKwcjqwu4CET8gy15aUo8874gQvOEIkau7FmwDfm
CH72PBlhGubmWG/NxYQBWevcegTD6MIRCEGiZTvL3aJG4Dor2dao4pIz6ejBqLZD+iqTAxp/apkz
1/dPLsVJWCySUJ/33yC1pGEx2sXvkvOAcdGge9K9n0bMxPE2wg+tvkTrzANrPPCnccuvvaXjltz/
o1EG9BfZi/MmdcWR7beCHTc5dlVfDmiECkLWgo9D0O2f/WQifvvzpmcZVTigO29oqYi2eSCefP0S
/9TBwK3kdL8M3GUVpLLgUwxQWooR4TtpTPuv12kgtR+VYe1nYLZgoC+B5PDi+OnWamZpsStl0KKi
uZ7jMOXJLfORv9mg1pouzanIf7pQB5pKNjxb+xSIwm+MweJKmEDA33QGIKcnrvnvY/OmO0JT7bSo
iMyTP3tXgg/Dl8AcRkBZMwK8HSCNZ105bLwnaSQmeEv+nxmvEpD9UOl3ueXKPr26PopChwg4TWzu
8hcD/cVK3cWvRDI+8XADuaaYdR2dDha94NfSoaHFwtLseRrv/P8uvoAjfXuc85d1pdLLGWLd/x0E
r6DfKSvEsj+zQWqSuWb2hQ8JpVFpAszo4pH/m5zdo6HisTcQOSqOh+1Yb1a+6raQSYszHfIuM4wI
9e63EtkkH6zlCynyP0mt4MqTOwWB96rZC1iYJ3H1Bm3envHpUe+o244yVJJS7b7djOj7wpyXFDrF
QXfJiEHPf6Ek5yC7DxfupArAYtEE+/k93XgiwsOcb/GbhBsOJvkyI1JNQqxrMFAOgwaJBjtfL07V
GNHj7pZNAzIhuUge70JVxwTFLstB65fjtQNw4BlDuCVlYuQpg32kRsppjGI47cgNW8YL4RGru/T0
PTYDk1u09NX4X/TfyOee78l3JJ9VQ3gGW6lH2Zh0tlJ6MN+HDoJhBOHXvKfiWSDsqxBhlI8Ma7a0
fHYMK/+K6SpFdxlLUQ7oDqrA9tMX5Yqbg4fO78L/53Uzk6jgxxMaQ7Eo6vgirHtsYrKNo+6vd2MB
xKerbTaBD1zcOcCE8aqn50kcOGVZxHZDo4dEGs8JvFQuftXOSjp/s4lZZSu36ZkOmLLK8+Lok3qL
rr27p7Ke3xrorLwygSNqQvemp3M3jyMukClHQpWPSciG9IZLJmO7gldWz8fcwexpHgrPHzEC3u7H
KepGhQLpICeblvEXSGE0knNL2DxfrujQ+AdUlAcF5HyneG38tDKxWuHlYp6BkKGmzGaMaR3qmisa
BhHRMYrwzhiJpXVt53njl74jwD24UIDaiP4B6KnY8ug6gIC8o1yMTk2qkyj3+goGohAe0wwX5pDQ
KWza3EndIvJxdeRvwnbYaZhM9uYMrkXPc9WVQL9Kt1sx49F1PC2SLw3XdY/U0ET9uMoXx7E6RB3a
zEbUSqNV+6W5VBSHhW0iQnA6rslpwTbyzc0S862urJh7t6ovxOcOjQAM8U/NbQ7MPIFfzdW37r1/
11pTLhcCq3+0pgXUbndzToZEVe4uwGUWFyzYZ2ZVZxJuas2++zfm+9NF2DBKdDc1AtzEgceiPtvU
H2yF7CfGBU3FGf1nYA2O6goEvDSQhDrH+f8Ob4FGlSZ3PI0bkmwsJ4rP59fLfb0JyS6E9oJmN4k7
o22AFb8WQzQZB08h7Or9cZokM1x0y0iG0Gl9Kpcy2DeAu4kosri7RLGtO/clENDEBgTE9zyn61XQ
gDsF3uS0bswPL2stfq6aTN7Y/I7APpzMiOzPXdqc2awxKUpg3ZjhY3rc28RGhzzORNmMfa3yU0RF
cSvxMM1S/x1SYGD5mjRCgQjZtIcyNVQQh1IGgsQPoFQqTWZfOljYHYp0OLrZcln3zf1gHrDOEEYx
XaI4Nw0KKFf7JaDMo1l/fKlwfBAgG8fYRWizqFRAZpYGvrQd0CTPn4OsjORpGFghEvCZB9Ez/rG3
RFAf0XMJumque8imeREX3s6QuMvvSlF5jDOd/zWUdkJppAMqEzCYGN7BgS1TDdtoVTteR0LyTP9i
E0GXzKhUD81APAn+66RJ3XRKBLacHkiF6CuNybIBqkwb+vBBhFtiYjI80gmrxaKPDZaHHC9jI0OF
l1gX7HExjzvS5NKDJeoP2ryIM68jreEdliSXt2nLp+kAJboxfqOdZx+Fna7MBgafuE/rK0OHxNcA
zwQoHAOr3S5efL3i7XhlaIOGdr78KYKqWXLBKmEd50m9VpfmoWvJG888yoQP1Wgt1nZVVhcrs85w
LHtPI5/TkK5GqE+0HVjKu3Y90VBxL6lJHS1XsNwAQJ0ASS0dO5YYqKNiSEpbYw1ecQBhzlMwFF+P
3VHbgIdJq9N6Xgnn/0I1uwGXlDFKlRX7702SbDItJxJ1zo8EsF8/hO9ycnmdsiss/jQSXPylosrl
92nwKQSK8HfYOwh4FeD6wwUpz24fzdRtDP1e/KZl6lS+VeNox4DF7iKgfs/hQlX64AAJ9RE8Iw/U
r3jqCx6YrcYwJNQ+2ebSoLxm//N8gPclVIWoPDGAgzbcIrW5i1/yIfP1rUvKCLGq+vlTw8nZsJvk
tpVsZAZNs9YTWyvZatpnxr2UVm4N7f7m2SJBDRDxVyDwuAuPAg02/oS6Thbn+WmDQxcirYUy2Op2
l3EWOn6sOzI1csbQ1Pjvtoe8wy6FgRLPF5e+MrbqtbAVRzrlfQ92PaJAbT7PMutAsTjdlPLou5pZ
MZMNIYfw/AzWi6NaORobcn2groZKNtYmOHgQXhVru7O8NDkY3IifSozYO/PN2gJvJqHprnHcmIG+
f7UcueckKwK+FNHqqc6K77AXLX+tuES+T1tx+y4+JOl56si6gUzfWAQx8sYDqVo8N/m52AAHpVW7
h7YnulHnXoM/xU2fhVstCKX0oxbII/dalfuFuzwpfBlwAGk2pUPa8MXIMwXJhHuwvF+CjaJCc0R4
B7MBUCqKLZl1djaFOLSGf+fN+xP2S0aEIhnGy32/XogWpM7vTkLvVCQ2TELcYss1a4pXepRPmPP5
g7HNd0QYDxTwbhRISDPxeDigHWLNa3QiPSQQUeLhdK4+irkUv28FoK4NUcLimb6+H+bv7ycUoWsh
u2/B4b7DtAPaKzsfKFFwMFvjAKQU00bCujAmpvmdGeApQHLZLK4w5Tkkt1CBAfh8UZ6djsbVByUE
GpSfPi/E2BIwtaV4z8Ogj42WXVxAsjNI/NFEWcFt7aoNHUlZIjV/JtNa9HKX5+NU2fkrDt2u9Bpj
A1fFCKh3MwfJt0KRmwDxGegB85fjQthza9Wm7DjsKF+6O9ii6+b+OEoXxbfykud6pHF5vF4pB00r
1LWyKtRAMmkVuC9oZjzxDLGZ3VukatHaRZfl51fXAp9AqxY6+QMG5MC/PNok4b2ikxs839rR/OU0
0s9al3xSkG31b4XinWSs50qWeLULeofoTGLPZeLKC2mP8W4qLWvIWoPX4Q6mE92j7/Hbwhjgt6xi
lTBjZBQpEvcSdCczghJfrAQTGfvuLfXyw0VN/V6evcSqhq74mBV4sfb16C3miTxQXopipiwndrPY
go02/UuZuveQ5h6AU2dpprn4tGi5XbL4Q3wikgtITUJTJLGQJk4DAYDohAWiz3C16JdIS24HvfdJ
NnNzlowLFP8fnMI9J5JzBGpMw/el3+sMm4Oouv9ZyegIt+XwDNRmtnjYaDXibFCQIMoL/IlrZZwL
UNDILA+w9PUihPeRSSuDWoK/9ThbbvKh+nWZaARxpPKd6iNAqHBwTwURG1oAjal/5YS38X2kNXzN
59wUkBW+P7dPMd+GH3BunDou32YQa+E59oWGyScmwphu1Y4esMUktqTXAyAQo6x8bZ9CXlHJbnTf
NWOIrfdmyii3GL4RPYkQ/mK9nzy2ffWSJWtkymvotmc36sQ4oAP+K4UxWj+qMH6F0KpGOj55Sw+w
/fLjRbFxWGg9+US/Ks2sBJPvKVacqPiqZBqYr63vgqG9xdYwDNEF+eFOMN3M5/375hXeCl47MvlC
Ixgi/DRaq0kCyI1wAbgHH1wR+3W/wQqOQQV1WILcC+wV+x8xmVmK558rqhHKejRyEvVSI15bvIv/
RvyGtTJa3PqylaWLIPnlYKxNSqNnXv1VTt0aBZyWdpkvhHWYL2RA/i4EmvgvIbjUDeydQAovbiZm
QJRgPsOLBk3gEwJALadGs5jmjo77TOwj0ka4drUv8r6T6Z7hVRsJOMcfmA7hLRDFduouTRkLTmfK
Z1kLhNynXxBsIzOcme2NsOcemL8Fjymgs4dP0NNAFC1K29m+v5EnuOoxKLdRiRZc8XR4z/muKtLq
AeLBUHncZx88pf/E3lTfRQEyJpSFMHRo4n5bnBB3TIadp2+yhHH+FwZ81UOlhssZ3j6HSg9/FbjN
QJ7u5b4JIdKrzRBtcwfl5NwUZ72GFCobXuyFGZMmYQIUh2s8gXsaJiR8pOg87JmFrMl8/2NWMxDV
qod0PUb79J8bCgFI9aqljBfpnAIjboSSluv7t4Tzio5flYlqzZwMvrztpUiGyDfWIHPggoelz/rt
9wL89jbz1bXdC+btt35mWO2O4oyIXqu44tzi7Nij+we1HXsWoW56D3UBZbEYL6bLJzjR6olIoO9K
iTU0BER9+Md4apATtN+/+qfGwSuS4E5TxsbpVhqxOAFK/lAsHK7cxIWSCdXCD4Jvdfm7f7ZKhWum
s+2s3faFzxfBGiRPpoGqI1W01FY620yV3bo8y0rL7zBo7TyrGQgiAk6uJa6Dlc8nsYpa9QEzbHC/
zrrzX7XfkV/V9QcbYTqeVHOtXhbaqoVxhb9Umvu5bjFBRHDG/88HdSZGu4Emd62lpfCH7Fw8tFxQ
9KnVfZo9TfUJH1csoVpOqxWGG+K2H6CE4fRMaTCXG/sGO8SfET5HCOGlsjvABSqI9Y0vcXyPrxMf
hJUzQmYUoeZhsabFUtncOqENooVcMvVFEo9lXwE4USFDm8NnQXNyqwr+SJlUhG3CbgmSs23ioqu3
e/Fmt5fmvCR6XiIXZ99dmQBf5EbvOgfHldejYuKHPORiQkQd7rm579vdOAicGaxieuB1RuECkhYM
8ReyF0Izxvp4vkpc0jiCvLGlEMM7tsFVh4l46rtaxk0tDHgoe4Qb5oqqcZRUzhCfOjhOZnGP2mer
KOzhAiLxRLdGn1GCiReQA7o8db51bioRmrFVCtv9GtfPrw0F4HZqdkuwwf4ofXi8uVpxNxPctQIV
0mrJ5E8Satc4+RLbU3fsi8bS/Z2fSDP3xBOcm9QJBPQD4yvqcTXoxgnRn9YEucXSIlWQx0PsMnHp
TnF9WWdqhgaRd+txrJwqccDt3fXIAOT21QfMr/oO4zibK4ZwZUvHDrDsLzbs3EhoGuPrLiJuU+g9
a++MpRZc+rlCYhlM6vZEIdQno/y+I5I2WxUSJP5pWFaspf8wD8MvNd6TYi4s4Gi/2s+ZZj7p2h7e
urExT/tot77d/pf1az2h73d3o8/vYvpEfWEGMis9g3TpQUQKd8hxnd5JDSiulTlUaR98KW79Wwsr
QCaOUSTMGnFpPnsVs0ZkbLYsjZpyMOnfjB/uz7WvslIEIZMfKBTeMqX3gJ+HM8w3EpqZaGz80SNO
XjZMP+B+LTN2CBUzthJvLsgPfVWGQ5D7oNDZIXIMV33fPHS538f6qU25qeBcUrKvoNIBKPmKA5+B
Pq2WMjbsJL9Os+YiAR1vpNQeWaQuxko+RGkB92xGOtg9y7eeNKKZKDPVfXLJvByeOtALLA/ySnWx
spXygvQ1xIoATPRC5ya/mItqU4KuiBgX78eT0ouU7LiPrj9wvfTmjMfgZ09c+20mz8zO11j0DiDr
Iemk9U5DGaQTEQm3snC9l9CSZRIuGJVELxK/ITl+obckzIMW8Xxpp/1xjYtd9NxJjH+23L+XgwO8
vfyhZ6yBET/WQM+sHUSiLFIcZPcf4ch84V3SMXpWG84wS9pJDy0AjHo9W9bjWR25amvECxag37gl
BdDmsrVbCeKrKP6xv4OCaUXXnqi+Gl7Vm/SvDs4Wq9ubUDptGLjoNYDFCRfdhTRiSWed+OLuAHwN
uPM6JCd5jR3j1GeNPCLyUbt8LVh3lFU8z5b9DnFSP8Br1Akf+e1xSzcfp38TRVfx0z4ZtDV9pC0F
FdkkALu5WfoK8HyzRYdl5Stv/QGmdEOoCSRphgDTN1UB4MC1YEfLhFAosUtPH8bxplG7hVbTYY2+
0defgc0lufz3O860lUJMPwtkB4cHzZuTLbiwKZwYy1m483ym2R137FOixUCisvxgLfTIBD4pOIB7
t8si2nePBZinm5n8V0xnlo8F4fOEfuU29yPDS2y7+9DOy2Anc6Rpo/Qp8O2ps7Y6o3TYiNxTKwiU
2JCgtitDi2wrblwyqbo8rWBD0udZYjCJM8K6e4ToUtaOYEl7pmJR0Uv1kAuKupukUh5EisHEsnpw
/KxsJ4zptF6JKPlf/juwlN5pdpdMU5T+P2cmVgoPevJz17kymFMmb3DlGAsF67EwuyJbyOdqE/71
+rpOk6UxupEsDwzOmddnGDub2gB8qakLmYN8i7QGZBRMXtp3eTuTUKerSkVKpyIdywMv6S6nAzW8
PprwsmAdoWJ3aGKYnWE8gDqmWEBIlHA0z7C2qKxUuxHLtgwrbNN5ZjzpyoB4N9MqlyKLOg/iSaZQ
K9w1ZQnvQEtSNvzJlAynmwnETMGVhitKRW100Dnxy2WYJA8XmrXvNeJqVWjcgvhDihbGYGwKyJ3Y
qPEgjXPChh4+rwQOar6BB8PK1DO5TCXb5B/76UhOkY0h4uY60PlVnwcB4HebeRfOib0gnOZOQut1
14Sg5jmhDAoIZ/weihmebgZTNngi0+eIG+OVZHbekkEpwLXuL5MKKUxiEPaEFMv3prpMEp0vyqSs
3v7uLsLypLX87GfXTNTSK4QN7S4ey6nQVQcjRYnzPQzBNLOVGNI5Fo4Qy/6z7POTf/1yvqemYtlz
d+j5mfT7glSxwb6ZPk2vhPm+Hv2kkEXIapn/38EHQIQGg2LeShauV3mEemmY6XgcYuzgJPlE+i4n
KM3YRtoAgObRf5sYbt+MrxvgKZ7XtgL3pxdhduyq648APSKQDLsbHAuNyTYhpUKP+MHGyBq4HYTt
mHWoTRTRVe64ouXrhGwBBRmarv9eFzl+cyN0GuFKcvuD7o9xaUtAmNW6/WU2VH4kL9L96Wr0o2+A
tvAXrnRG3otxMzksLRpLbjj9pb6VWesZ/8XKcgD1e3BayIUjSGG/VAepjGeeWLefeXXofsRwFGCr
UUnSNxE8/KRTHGlllogiNCImTG3Ss+S3ZXCCgGRkX92a8Sq1/rdbsNLcOUVGckqZs9H9Wi8ptNK9
V/nNWFb3YVoCXdxK5vAkScqm0TJzV/iunqeDXi6CA64WVriyxa0/ZTZbZv9c+QjzCeBp2+4rO2wL
/U0MvmetMqbQ4vNa6bDrEO7tKCPpqi+NwS7A28LQIwFF44dqJWqjY2bCjgy9v1i6EB3h6amo27Nq
X1SycYzdRIvm9lcmg2ugQXyGgPMpbEn0Tbsxr2D01d3OwdkJQEejocLWjVNjy2zqbL72sEZT4UpR
ntAXMHgW+VaT9EqOueeRTAZU7IbCnbqW2Ojl8AiQM4bVDL2SKPdmI8k4227c2REVYQJgbduAGxx0
YDa5paNMmQ05IgWSimrHA1iiG5IVLm1NUa47ZLBbWiKBrjRajysxwrAyjaSinAs4bwpnGxc+v/c0
z1u0IB0BwMDEaYH3yTjfQfK1gYCU5OCEdlQwwq1Qm55Ui8RX5PUpHPyj3Cosl5oW6+Xj8BYJrPbL
BuT+eQQSUi+gyg7ickmyhwOJY7Xp2C47ECTKALKzTmluL/k/Y1Q7zkqzr3WI//p/Ua/HdLb6suIg
N0MQ9u57uQgqnCFxKBtqN9k09QPyrEc4qFpVWS7uYRd4GSS7Sj+iM2M0K0IW4Qnm9xsQaTni8ehp
uIlLADGBKfTfU6j/kWRt4O2+30n9WQTx1mtpmp4hdqQQVkWCh+H/MrpuuR451ggIMOlf9ZvIkJa/
uvT7TMKJY5jtAgGOC6a2dOftVMErGqSU34DwTs7QC1JZ1mBXCGUI9XquyYgsH7QiL8YLHOD0JeHq
2EGxZDxqqwSVIkqrJNtkk/iFotFo6BhVZfW2zePLnIFaWIuVQy2RUMCgG9PWvOXMq6mXGPP2/WAz
GXTKqPHj8/ozlWT0qlgnuBd+DFC+n3LzRlWsj08vF1P9/7Ctro4cTYHu8XZYFNNSH8y1m0QbJN4H
ZFYAWUXew58Excq29d+hfP/AxvrQ94dyrjFaYHZHEeq3+StD1YlI83ygH9T1sBD1q6En9jEd6ySr
9JiTLsLtHXKGsoukcEJETyiT9WWN+Xy0ZNSzf4mpfZk8W9xD6bzZLrR/AkX2sKfmMGioEYrXrKP8
AqTRqoJ2sXxFmRwDeYYUepabckz1sQod9OaTurde1L2y1aZXGXq/Q1bk+gGmrIZmwfdcGlC3y3mM
fjVJ01vvGqbvIOXI7jWLAi429yVgXb/rNuircIKjmxgK1Xz62ZDq6RS6nj1taExh3JqzpczVUTA0
BCwk6os2SOn3cik+Ovozf0OHwwbUBGruzq4M1IeN1Guz4GyUGHw6QMnkWRXuMPJ6pCTk9krlrTwh
Dgf59NREI4BIFPg9TPo1Pjw6iYmqzcgpoEcuDiO+OverLCvINXuQ0WS5y7UjQXOgtsJ5kIwEjBTL
XaBxozAOdxvOYvZrywCU8/BWU2Fw2G28Insf+HABjH6PXsszXOkJvzmXwd/4sN6U+QxP56NZ1Iwb
O9HbqllqrkqMyxm2nneO4IwXZCgzj/On6P4nhCVpCivinxZrf8Ye0gqlg1Y6i7TFMvOWwLn/noo8
cPong0Qn9CLeKr3h26OwBqFc97nLMK2qBlBhkkZ9+B9+kkdBU2gcj8S5KqSzWyVOnqXX3GonVlAf
1BVPyZxg2HdOYj4Se+r2jBsKb0Kc3E1K1HNUL6rQD2AFGvhvl1xeUCsATKTsV/tMI+LDfe9CBm1r
aT9rFxVpUkLEJSJfvkqrlaVF3K87sWN3AijEu15cHlv/Zldb5/1kNRyfwu7vdJ9o9hb9VmjUYDAr
GX8znmJ46aLGZoaRWMCWGn6/4x3kEn8NP8evAeppx/Wf64RHmEO+F75zQ9bnUUJE6+k79TXNcVl7
kw5aJozmmSmIF3+NIcqBfA9OJCydSRHf4q5UqbSwBLhVeO1EObkEKNsIONvcUuuoK+YkSv09NSrm
qiWvLgEn+riNmfvwNbSZO6Md67HUN9YyA6A97sL0VRHjveh4dp7xDDDWJ48gVcdEF+EWzBUBBkY1
fmH2QzfrdIchRnUOjRuwTzyGtiHX+XjCsPy2bx6d9flprLFaD/y3KeoPHQyfyZVZbwK8q0u4LtPF
DOZx/l6Nj+mJTjrBZyFrR6VbhbgF92T57FBgL2i6HZPWpDaW9+Wu6kGsRWZgqRBBSxoljgYs9EF/
rxmrIUP6E52C4p1oh9VJcrJmugo9OPZ81/3YGOKWgq03rZsI4KyuOOU3MSTcmEP+c1bhRfDpU+cJ
YnfnDKFt3DAUxEANYNkkrFwF7B2jOZxr3fZqCQJKYT3ZlGRqAZNbm2fxbwVgVVUpLt3NFvr9Seo3
pyY6PLiVZnhnoeUDZ1UxwC4gCpzeKvZDylo/CP8ZalnJ0QkglWIEokWn1dxzroRjMhxmo0JFuriQ
MPADqGmudWVDV4IZtJRkG/gPZ3ywdxZiwSO40uMmQ6JZpIJt5j1DnC6Sc5wLZovkxQ0HSBXGZwal
lPbBgRE93hw13SFip28MePaq7pQt/irsH8nxAM551Y1fc+Qg6awTYZKZgVYFD1lAlIIGHKoZhAj5
j+xXqIAFIxGQcyQ8/GXlxJWYpoiZenhlyoASn6S7GhlQlzHtDd9gX9kEVfzygCPPwId4xa4pM1Wc
LDWsvhb04KBD7catJBluWnMEwdEAeBb1+pR0YttGV4SPrjsy/UynaQsWgOffOSZgLP5/G+hO6Uz2
Uwi7E/uUqDnKY7d45Hv/I0qqMWUXBtZlfIe9voMMB8LRiim00SG+MbnMD2y3SufgLP/EcCNxDTPU
du/iERrfvzjlq1omEZmeCcjfaDUSfm3bK11t4zRkejzdU93K7lGa83Z5byl0/jAj5wndfn9PsxeH
K8Op26crNfDcKnAG9uoFu6mwxWmtAMPcJx1uE0haYDJzVtmfBbxiRGP+oDk6iOKhqhSZHKLhy1p1
+RgRzQaRTO+e52untpZtAOMEsWyaM6Pzg0F1iGa1RYunKNpqdymxJNyEf4jcYgdJv5WCddQe28/4
zaJjcvTvFxNLSB2Zp8tuSnfRy2sPdtxdGvk/TK5pL3hG8ZPrbE2z7Qj7OdGOIxFJTAj/vYN8zYnu
Rezr4nebiw8Js6txmiIy2p7mpfYDnfKYLxs0+GbWBVqVIBWCFrRZbpFyU5zhA5JLCCx54LEwXZNZ
DufuHiE9Jq03WpVV1vzMUucpPhxPv/4lBez1HE9RfMT/BH3EkKq2lOkSLvaQr+1FVSykOgJVThU7
6/HJalXHQokVihiTovBTVFzsHyXe89oGoSuZRqiuQ9r47/eIv6O6x1iEQR2mLtNM/mbg5XqcJFCo
/QrJA6n48sDQvleyFSAJZ3Ppvl38f28InjKaMZGsoeY0DWVeYtdd3/Ce6oAZau8TReRipAAQ3vff
77YqJ2pqeDojlwlZ22fkcVgLXmwLAfzeCpsoSPkBKuOqARdRjuk3250VZz3LqV2+Zxqg38WXp7Yf
C6qw+1Dav4hLuhX+8lUfKK0pFaGytn9TtZGw758UWY3lIk8dOADCwGVwpMmNJvYrGOjRLrKM2/35
0UaJoFs6DXcwHdSzLk/bsYK9Oyw2fLahRt9DEb6lthyJEcttjNejeggzLwhJW5asWFVAboUVwBMR
mu0TmiKFQXn2VNSCYwYCOqgaXT23GgdFt39hBw3DhpKAyiIB8NtMB283NvHOjFnF5OgRyqnNOlUN
RMHun1TmPSc5Mtc0ZS3/F6XCJUteMCLbXRyY0JjfseJYyq2WynzgbKe+vzmnC7Hc3BcHHl+0RO3n
29pfoVQfF6yUbSp8qY1XAWUCEk3ppqwC8B+fWIvUFXzZJjjvhW5nLO8SAoVCYZ1LbwSzqAPI5P0B
ggZIEXOBRoRbaUiVf21a4e1yusyjEIUJOUj8OCpwPYe/znp74i3qPs1h82Da90zWqLS6b1D9TEAf
YZj4p/MaXUH7Rp5H9/tW4mR8sQiqR5AKrhV2oMFd9/JToucZKj6mLW7wLdPsJNut/uKGzMJRnALc
wd6hXtuxd97zf3fVVECDlahA1hyFSCPxkXm4wwGyodqquA5lq5tc4YVLLxNF+nsDQ1vYU8ZZBwAX
HfprgkVh3foTcf9a3MiBtFp/SU05WrTzwkU9qVlhtZhJr0TL+u4U/wCyMHw9IgAL4+4JLWb2yyfP
zbKAXSjEw9FIGeXRml6ctf/67GuTzNZT11/JIwEcUJU9Nb2p7fBwgCUMbzZW68ntOvZiSKJmb+pU
751XXaZBZa9MTCCu0mQHptvqB/QEcRxCooHHzhwkz5EgoBfpl1Km+i6KTbcNqb50fFLPVXo9uBLw
b6AiDDGrVgU2dAMv4t8K71aQELtuocIWcy8kzeESzLPzR3TrUWW2oJw+8YM3eiyb05XCPQLLGIMH
thgRQiBd+JAae4CH8d20wgp31WWMf6IW3TrNNHpLVyCNW8Be4iNoRhlpsKH7I06TDRTjDRW3icEn
+OhOaIu/dasCyCxIkEMbTwxPKFB5uDE6oNqBuX5zHesxjebRH5hmK8cd4duzWu7gegKxotktNN/2
WYmUU91PtYDdsK86AOvnyUeyI+k37hJEWeMWYT4OUYVH2Cv9TX9cho9OEHsCxMMRqca4trDpNybF
YdrDAB7Hv/dPRaoTwEtG7GDk/Ndt3cVRLGrkbHIiTP4D6hyAY5zToW5KRNXSoF++I9KYn9p1Rht1
I1NajySaUQXr9F/4bW4KDmV9SMYLJ53fGgLJd1dsgNqlr7SdXVhBtu1zqxy6waFNtk3OY5CBsPaj
jxNnAT7VwvauB9VqYLpgfAa+ktw1y3qbMWPrYw9BHtHD6c+Lh2jNwByl+aWUtpXI81sCnAo/h6NF
83RtIJAa8sNVsM8ugtQLIJBWFQ36SZpdZR4DpH4sfnRWHc7ZokpuaXYRo2TcJylwYEjDd90JmLyI
PdwE7ODGinD96Vep7/ibAlpcm2gL5bLKAKfmezzctsP4/n8IZvJYFaygd+Mlo/61hPvCk9ZkkXQs
8ACCXhY3NwcE9aCMQ1aRmZhYLtMlmTeRbd9KkhVR+fKXjcN070YHFlsPCR2Y7qHH30QITDikLkiI
Q+C72brNe0kgSgQwfM9Mm/PNR5PVXyNh4TF9/lXaSuDEDNVNDrENs0hiDm+4LJy7UBRk+B/OnolB
tqJ4dtLeQAscifs6IwNwpYOSKKThBBJrCto2PIQBOuLjFa5EUrDljk+cXp1QnJ1+txRW5nsX3U9a
Uf4n6bGcqEYoTjv6aR3E/mJN9ADmTvCIDLqqc6dEUbIEUbeiyxdmVMGaxPRjSj4G8FtBYMySvX8N
3HvpL9jpxXzgYna/MLompxPpYI2dzUb7KssqUXt3T8KeFyqdAWGf4d6AAbziz/K2BCtJpnZ61KBB
jM2GDn9TBNo77RTyF1blGjafDvWDAeE1X1jO7VzgeJEzbVS0XtlTw8XSuwW9BJhtxmaMrdNzlMDl
EwnWpNnfC3S7j6Xw4VV2D7xqvSU4zK2JrsQq+nNSqW033JN4Tt89Xy7RaOZWQkGonOW/XTNgCQPN
JEevCWAqBgVQDoM82QqBYNR+tpT5fKKVkB6Xec1i1qujG1zBiegLryPtHBuVsPv5+/NKvTnJ9HYj
O05T6mHHFT5z6TAIjbmTzDtEzWkgie3BlzERb1bBp3XM11j7ykOU52NCxj2z6G2w0rMPoXH7AmGx
Z559Fx8mJiQbcFvV+CNdE95q8TxUAl44HumT5qKtgJ7EettGjMUdk4XUY3rSM7SuaAYS3++r3BEe
51Z29nJ+96KA9/WAUaCeGegheQjkKjya65OGzaHxJ7dX+Zst1jyW23/73vc6DoIRi09nQEZXqkrh
EvRKghiUwHWw0lQSu7QsrjvvN6AiK6YGD61V8zvvZFJTfy6X8NOJPwb8oqpznSQeGKSDjoRxLUrw
U33uGJNZhxk8CJODges1CMxhgUnKUSJ/3TEFcrWI8VmXGB/qViJFKqGKUfvWYmvytn7gDT/K5Zy7
wmBAkBLQsss15sxC2y1hP1F6tU/+eSLAkvk/y06nSH84ddDNt1c+WodjCf1c0Kstbyd2CLuLZhOV
Bgzq5rlftfzGSOWA8GanX3qd0xIVYyFkmGDbV+NwaPGLHMhJWViKQlxs7JLK53PWzRNp+c5D8h6f
y+vxyjhI58SJR//FRWnJF3X4Bc8OGx9CWiYj3t8lrTXlMTq7uoeiRLamRkllOsAwybc3hnZpitPT
i6IIzAZUe/Ii36jKaVPjFZONqzRulImkTA3ClyrBJhiFQ76uNNPvVyJIvoCl/l0b++G4K1wObaqW
BHXGru5xqzkWVWq40Fcl91lwoiOBW0La7FkICCEO8lgtKl63UCWUhjzep2bP3Nst1RcL4/laH1ET
RYWdhAviUwmBwtLwJlBy5wVLJLIkalXBinLWpBGXmMOkagh9RoJom9wYFe6nNW9s8QxjUR+NGFEz
bLkJdzIw0eU+1aQ31WQrF9AQwjGtIv83JBVCtN8ki+XWBM9wxH2gomKA8MJbZpmYBc+9H3Wb+VmB
VJSjl05YBYA9RyzmGSYWIvGl78v+ebEfQIjbv7b70oaT9RzVwkic1Ody6hdF+D43xFa1XgcdaQlI
/pM0r2JbR6zBahygTMaLk9YgokSTwcaAtkts3vgaQAOp+7Qvs3vbMBpYs9F8Eem3oa6auwCxFdHu
wuZ3DDi5qAQJWdQxcfu0EUCwZfpdkK3orMK7ly0M0Q8ctvzXzN4gtqyehwVo44oUamvfDJcTteni
Y0jm5vf4sVp7RAD2ozJ1rG+Ucm0C70oicbJZSb993FTFbqHg/6VcHJqnoaRaY1GVxCU/jZs0cwyX
r9No2UboB59cqmq5CGtkz0ACvzG6uTHB2G7zCndJldy6M1awBhChIRAoqqimtD3aGgBwGNKH7CWL
A8zdge1VQ9t4ohIwdWZNt/MIGvDO/jEHn2dTUtmT5VXi1wcPIZPpo7d+8mBThNKItEXK5DXZj/9B
6O9FyoVssrEf25vh66fGVyJJZ574zUIl67vtZNa8hlJ/cRvwpRk4Np0owV6kJa6Qiv2HVvw2EO7a
y97uwJcW5gnh58dBb3zYOdBVAb2j3BNUou7Nk9f6/nwtZUvhAvrIWZ3b/rNuUpdzSE78NZqa1yCN
GActPxeLcNiGFCobDB0ioyI2kj4aS4TPvMXpFkU1mUTWkr6UrQCnJwv17lrdvfbbCVKWXYEMdUd4
RXDY/B9Io/Q63EtM7tB8aWLEzMnOCFWh6IQrvtwkxwYF9fJzUsO97c08Mczip5jwgM2T2zw0Z14t
L3jJiYOCpoNeNRpdkyPyAa23iKGmgoFkeXKGUvS5zHipU+lyKRYaeGKjIDicleSL9MUsniD9zbyG
Uf6aJm2iziHlEyq/RV9i09WBkoDquJimd+4vyKVU4zcDoha+ANNgA5ROgUrorJ6jj2Z1Tv5ILRgs
WmZcjcrc6eLP/nDCnvgszYDVbrRp0E4wj5d8T1ROWnpX9qLryh8o6Zsa2z/8JWefWnik2g48U9Wl
yS8E89h1J5FQvLDrEWoPi6aa4/s8Q9fSv+kRdcEET/VV1R59SGiuue/zmQRiigx9Zfqca7+IBIx0
dFd2KO2nRC4/XpDdN6LkNwR1C2/e8nn/uZyMgZA/KUM4qXTlnd1EOHqZoqSRscziA4+5wk+q1b+Y
2cM+6aldGon41YCuzMNxSl3EPFq30ZB4phIFExQimsxyVZc82y81oi3/d+SGwvtSoMeINOjE2sp1
JTQol6rDhfeL3PT2X1asNCbWZF3XalCMCoz8Rcv37tFIFVlClp7O0CtpPVDANAGeOTFMaRazrYMN
wYTiYqQyKcKcyJBM1y+5Pt1yQp+NphmpYTeZrWfOtjCAt6x1CINfHaj0ThmZUBqMDTmm0EQo1BcU
v5HDPypDKOeNVbq9+ugRQ0GCXt1gpaOAL0FDGX5EeaDsenoPhBoR2Byf7f6e9RdCzZ4HrfWdwc9N
vVz3z1jnwiutDfZgLExx53+LbyjO+qGk2JZV1hb4kZqxaxaOJcGqikZG3QOMzL0y80xrs17+QLtm
EkGZOt4jBIyStKQfiRfe4p8i8gYRjolJXJtQ6KAEvjk7ouOYu83Sxa16WvM+SmsnMV0FsUs254kZ
0RHQCeHBVZiNxXDZcZde8eCf3N42/cZzN8oslAi3eeXL8hIAw06yxlX2QZmExucpprA/mrxFEzEE
nhNs7zagpSxAUgCx/KiIzGURzd2Y7IweVqBGo1L7kOeOCb4ppgsI+IFFGADTYXyKfHQ6sjx3glmj
0dQTjUCUXfWHNpw/Agmho4DQEMREo43bcWgXWGLglMGnnLyoSutjpZkviyE9cUCGWQ0hnHskOhuJ
I5FGPAN70S7iNj+lQq0usB2wkIgvq+ATxJlqHI6EfxBTirxbkuKPz2SACCTT/edzQY0p/AYRIVBf
52te/fvSk1E1l1RdxdxOZt5PbwWN14pUUSjJTr6EYuUmJbBvMiPuK3TBQ6cw7gx9Z/WTBwVercS7
CcouROPnHvvxkjb5d6OnG8xl+yucFlZcpxVehfZQ3DBAGlV5WckScrH8nlzERuzFJeELRnU+fKy8
vIR1hF9dwJZ8L1kRFuOBSCjCFeBoCbi89DDmmlpFuNzTfmmxJH9xzr8oh0XdtoaPtRIAwMYozOB9
/KoMSHMdFJNUQIdr8h6nVuYiF9NETes+Vw9ayRhAfiUXGgJ5l6taYtsjXHvkoBT4OAdJi/j4L8zC
acNSCJsdbEHFzYi0DhDLrpiPV+c5Q04MUHOgz0KHh4+l9+BeclMcUA8LEfAZ0XqYAlbOvY8xr9uq
zSGH84GHRZej5omLCwKeowR8LMY1mTBI4KelWa2CziiU+cVyopOzJzfoRa4ETReh8yLbGO+XA0DB
4EnLzR7jbfUIsywZAE5BHIb8cE+frI/RkpY6dlmz1VQmDWxuQn+MnKqctF8e/5K5XGubZR3zU5o6
Uc644I5AN+2OpoVEh2pEY5LCygQAA7wjxepk55BGyblnPFRboMBayezCZvQdQWlt0ulWrda1AOZP
ltDnfxt3aGRu/5EuGLsbpc3SILrm2M78tb6Ecmw3u3czv+Q0qGeJwBxTbF2X8mjq/I5QZ7+wKF+g
hNr+fOOx+JMRTnMxyHJgn+LK3tnolAeHQvmJAiG93sj1pPUwCprgf48wPYwGJVo68l8Ay7goe2O+
aPbHtgr6afqjTNbwdrr5yIHJbMYcbzMSVt/CJN5UnDzGt92bKYrs3Y2UbLSEyezYmi2HjZjmTg9/
mAJCxCOrJNWBRk8N/LADjGXy2p2dmWkv6y92H0GE+5lKwOy3gacxobsh+nNY3sc5PLNMgAIuhlkM
RrAdHzG/hePUpSY4aOC2zTX/cYDbenlyn2FqtTIaFNy3oK/nHbzZ5Mt6h/Ea9eOaH/HNy9b8i8fu
/Ui5KCd8Mk4hfVrIoJYKFxNS8kfDZiR+MXvp9nOljIVmYcNj+gHVfO/Js1K4cUVcX5juMei2XWpW
ohjoxw8Heg2ngBzZugNvuSLR2drhl9GYRRf304ns+p4AVQKVbPur0TxYh4VFFL1xJz0dXd+Rc3+s
dOksJYBe+AI2D0TuVoYVP3XKLMv7fu2qRRAxhzBLAWaREEnBKz25Wj8gpFyjtyEE8vkH1Z42W32x
eMsQnJK78l/021s0P2cOS6NAvc02JuFPU6Ptt9d0oMjT5dtrxVnf3USsrxSKgL5IjotXukA0ht/+
vMRUkVGcDIKFFp/q5/60+gwKRKAuWRamDU+ATE0CoYfynBq1VAFTS0eotjMc56ps0Xjk+xuGbRGm
rus6fE/SQVf8TcbCAkfmGuygYFU51LxsTAVkVg2D2cysAAjeXAfZLbOvtWo1+uqgDO7T06gQJcTF
gfhQjYN6Gw7j90Z8RM9Hf4qf+2vmiVL3HpCJQen9utQduvgeezUQyHvexK0p2T2wAbkkvzVKVFtE
0H3UF6XZKE3k+/NUDjPh9XEs2CBTP3D30F2q9dCkDOdhEYXDAIKb5oIp0Q65F0lmUP8OJ5l6npEX
y6jF/qkmbm6hyXoGOUVR6BKpa9NejFNi79FsSsaLqsFpD0U/QOAAM3tIrS3EMkcfTMKZLZ7cQotz
IHNkxYbAGDMdOZ34a/TX+KBR/jT33Vb6XCU9W3eOoTU912LxAR0Nf/awh06+BBOBK71tDH0w8OTH
O48fDIf0Rmr27Z0tNLTDJKmYQvr7RcRwV9ewIdyIbXiPAXasXkZfFhFMuPSCB5Cur9KCWCNGxu0z
D/fa+51IQ1yiJa8kPbV/mjRXx6IgComy2bN2t7yZVs7sUgIWX2E70p55d/g9I8bO4CfKZ+9lhvt0
mruTNMzrFxu9PKlSrLLLP/xbyMzjhM6mz5Wkm4G88bztC3LpPmYgnTu5SA6I0nhoY+BESq2SQTCi
Nq0KUcEy0TqGa7aA0+taU2U+v6thVZa8L/xOzoRRT3mVJh6M19V24WEVY/xARpfvxyrLk5dxUfSB
1weMpogKw5/TsaqCMpV3ggWDeFTvSRv/5EhXgh0XZKVOVs1KtEsqEfOhwxvWkj08a8C8qxDe01P1
YBp5jog5WGQFTdq+xc6vaWOWmu6ux+iE8DcHpwYZGINNZKLWP668v2PSYNltBWO5cHl+ODzzMlMG
fRHxn1eo/qQ0xVnrOHovch8n31WADFtdKDmVPzEQM/WfO37QcD8TZyiQ6oVZ18vWtnfdKyi2/z+g
Nyqmmtq0TRG9Z7DwJxUmOkIWEDWp0mr0kMxhmJDLZc++UDRwI3DP7x7dhkDwt0NECXzOx3s8nlWQ
mvcEbiiwOyBWr3XvzN2tc7xcd7s5YhpDSgVBfvEV89CuneCRrsAA06ay5gMlc2Zr0+qwLPjqhX21
eYM7TZm9D9ZQ6S1HRmgSO4n/zFJFFp89iNvwkrH37wZdpjXV50av70Umrzxxkx7ljUyzGnPFs5Ks
C5EkGrDipAB0wApghO4j5QViiJr0dJrq4LQAvVu1VbE9zox9mBV99+wioFTujb4pWj48EuaCGYmP
2+6IXwTHkJ0ycyQ+2O8Xv7rIwIgJaJzlCI2tAAIHzfNb34iCHVDSkrHWz3QZOyGYkHpvVZ+Id4E1
iE9hXUIcT4Or0JAavbl6/8KN1S3hvXmnLwTex9OapS+ytsK1gTF615eLOIOjr7s0klS71qSqzeIL
RJoTRJV8357+V/17JkPaJyB6Nb3lHjlaV8bbhn2qqsBtQylP8Ar2yYE4i8ThiYsmyPV+xAALy9ss
HHyGmYXctcf4+zW5H41eXmGI827d+o4XBmhTpaEYjqrpuOQ7tBcyZsbpg4PTLrpdsJV8k73R7juR
wOJN5sXGUvPa4hEY74bP2H6GJxgg45+kgJxvBB8M623P5xOvl38BjayNoEcMHGLr7Kk+emTjlkOC
hJdfjf8CVx4NWFpMCHxNvPD1I7HvlSLbsaIcIew4KZMWLm9O4PSqj9CREXdmy1cIwD9jfp19euGi
fEIXkphPwqyaNcqJ3ctZZX/qzwcDivvrkYkWlBXPfGTrZ/GOoJu+b3TgDIRyRt+k6fNczey2TSKG
mRYo420m+TXoK9zve6d+UC5ROjzrBjz4pCtInjlMG8Yc3AFKmwooTkdYfUO3iPkG7y/Sakq2colV
784ZmKx7tNNLOM5dJLwqsXOrbtSrTUIFHd/Y09qMuTkHG/0NNbO7fOmF+3hVkK9KtQqbt1EihSY/
JxWYUMEGn9y8yzbDdc5tBCACMklFCE5aPzblymS7nFFo0T66BSfR7PS0xzk6l99NiOOH/MQxUfdC
Qp2BKLK2+U2tIByoLz6Bl0vlcfkcgtAr7HWEXZU6r7lqJm+keU8K+ghQ0T+1oay4Mwz2PJstO1q/
SE/GYzAAzAmghyJDmI18mv7jI9urLQs6jtItXg3uv5DSEepkgU8AxS570ObKveJ+RiH7JYQe+eDp
ZmdXuGGVud/lyEiZJgsaQsz3MRsNQN+M1YlRdFKyb8RxO5SMeontNN7E6UqS5vMvK74WAevhxE98
EMMoxpA58Ci8ur6TvQ8tAnTVoFRKQn9UNI5ZKxc+XVZZUC8wg9MfNo8V1vzhdGsZTVdD6GYoWElW
OXPBYpr2sqX0KYWk71ZH7XgTrHARzvM+h6s9DQnhD4ySbBKMqKxKwXRCePMAxJE6uxSYTaOIPdVe
vJmKc7EhXykMibvhJD9L4BfyzVeeNxT+P9hHvb4rHjA0EXn0JMYdKSDaF19eSCR948YecszO6fYq
L3UV7hB/f/w47fy9rhwfgn2yKasKVwkTONTn69ys1hGILq7z/dSsckMLWErfuRJSTM3Nop5jw57S
03huGjPMbqZWNMMJrvwWanNpe2Ns54fNU6Hyg0kUdbnxkS3fRioDQ3KVPLwZpG17+Aum+dGEi3ws
v9AAnb+qrQaCVtRSMCBtCkxLQrq2XUHJho/I7Ug38+S8fMZ4LwlhF8bkTvj64qhObqDQNpA3LZ9r
WyWhskhONZc3noKtOG33TWMskbogiomW0ukojVgig+6tS+y5aWXol9tF2PLt76zJixs/brTqVfyD
LzbNrECWuVOC/ASdrBSTIYeL8n6Qa6ccyt+Ro9uYud9y79P95o4UitUxZkb90ypuByhBk+rZ1GI3
qOAdXV1Wp//u3C5mPFZhpKtNGZZ1mxL+SbGMhjEJvJTz6Gl+sRXyoxpSvH/Q4uXZmESP4UOp9m4L
feYIyWWORJS9G/lsw/NPE9+I1U57/JbjmQYuswtQSs0QiYQg3wMcRRtdLHIjlEEMPa7AD53yLJzC
5K5MDhFCPZgarvesHkG3oknz1EOqltrz31M0yMwcReZJ7VBpodEwkwA06TwekeCTtOfIuFrm0RX7
STFeuB6nenwT72ChO+Sw9mF9ctSsrsdCVs7RW+5Z6FWhlmcSGDWkycJhit2hi6Ni6VBcK8Fu+yAw
CGZIhjMAJhj6tI6QtWHejNeLa2KNL/ctuRmajVCpmOd9ktqGpQGDSDDlhzDN6Rz2QKtaLtJ9LM8B
xPenpxWMwgenwemGwd+r3bXR6tRgfz0XgTGFv+OF4HimF7A9dctMciehphsDONqGrkRh1IuvLdpW
tVMJjp1yLjviXW67MOOZX71aohRXS02GrfhRX6WQB7rVMurr4x3a2/+Ynw90fQSQ/SzhiU0onE5y
0xyl28+Vp0QlFWfkjb7OpcmzKglbSgWlJBWYLMjaKZazPDUoLBkiyUgRPs5KrYkI3+9O9qPSTAhn
cKdgxwA6osrtsfo1xmhDMIAZpa9SW1pJJto1MvokxvU9Lf1QQJ5Zv/gwXBX8Svk9USZrG6LMfwa5
wJDExtl2qeha2X4+Fi8BdE/ebM02n8GLDIWpNulmVGeSrsDManY5Fwr2NbLYPuKxVCmNvieV7Tu5
ciHEOvU5H6zOYKWWlFyI/K56DtrvzrrxXVahuJxzhCy65+q969HNbAfAwQ0OFWUhT8tLEN1p3Kza
bekySz6KjhFwDQEdezILil3HqA3mKdJL9/VkhJTUcfDs2KV7yoKJYd++FQiKbnj4oxSORpVN+IRb
VaHDczmlfWBvQ940YfjitfVSPaC/Lyl+tTWMLewFYHTZRjHSYI7cw0qNNJGq2JT4mOYpIigSuXw7
7ztREMl17WK0GAr2c9Oa9OIJl7EmK+hJOOPsz3MhrtjecA1PX4o7TF9U5fGMsl25UZSW/O2vGsiI
0O0Nj8IgehbB35iFy0me3pd5YrlsnjOsNG7dcz7iBzhN+ajK3c2f6prbvQTVjn6yIsXyQlQDpwZ9
PMpw+Gk8SFZexTJSkXbrIn+B8vu4Q/1xH0bOtiBCswfwB9CS+ShV3GWZ+hUMVnBS2NIz22z+umF2
hQaJqE5NIaxPj7JGu3BHG/RR379mB98U9cuBMkP63EFmqPDYGYniJBv34pxzbe3KKWIZmtocgMFS
P7n4yWFBaqzBVHuyTkfAPhBgvYht087ls/70UFLRd3JjzySTq0/RXnz3DBSvIQ/fn2DutaxS/6X9
pwlJ2pauY5j04bcwZxT58yDG8M9N6gOlHWE3D0+wU2k+vnqycBEvXS97UE3STsDWCABcNhBTPp3t
mzmj26dWxdTnwNdPLoj3p5mkF6Pd2D3PTkxJw0LTBJQGm8bcM6NPvbvV0RZnQQfAOJYQLhe1Tbe7
Wsl+P5SZ0uuN1NhMc7JoX6KCRJgKcZ8XQlDtp3B/mTbf/5o448J6jkpj8vAKH+tzpikVUQvYDrDd
YEs3hpmuAzuLNgyXIjqLjlUAVvb1bLJbKfGZuzgT+uOPPF3A6lU4sKB1Cu4Fw50Zv6L8W0AQg3rd
L4q4Kk9Kqom1MkopF5uRnqAI6I5KYTGrWtKXpG8xcaq2fwGxMLvq5IVKOp24rUruOLaHI0Ij3Zij
jEUIg8aEimlLv79imX7235rziDRiZbJ8l5EftlM5whp4EZkL6V1iFMd5p5t8AN93aKwD3ZaAaOfb
OYNXWO+skenI7Xzr5MxJD5MoRfqrFfJZQHUerAxzPBgtZeum97V7RQd465GstI+/jUJF20/e2e7F
K6UID92aUiwgOq5gXboaC8ajVfDGtRvzdy1TlEP6lW4XLaPrXbm1rg0gXOWdBOWczkHr866ldhWM
DRpOIpJ/ScKSZN0/lfzxAdhaygMXOtnh7QlyJ+M5lc+fGVViRkOOhPrkem6fvqFWjojANfcecCSz
Dt367Fa5Z5uFd5X1NpGme2b2ln/ZJfhLKpD4UUqzCZiBvZ4o6+owxUX7Z9Wne+gV6SqQVgqqolQt
WteCfYVi0DpPc3TAVXKDEx5jj2W/ZADb4Up55fS1+OcW43HhmWRWzvkKthKJJcj4uiJbIMw9Kyaz
dhLvIlOcDnqV4c2a/vLUdywPrpR42aUDNZ/C5e9ZuWIH/4VyCVlhdpzazD7f9Wje6qQhiz4rdl7b
mpX/2h6HdUxvaBgj7FgVmkE+T1atYU2Fo36ACozetOhTxmdmFnvH/sfgUGoSzxffd5IUEiJuWio4
uAT8LCxfuFLgG0w6MPgVpxAUTWAXlGkKWY9JiRLTxfzEMAfP3jjrzrb3yRJ9Brl1JmUbKwZgi3qx
8XpZSegajxVsBHjqQyOD1GFZx8wsB5ucdrK0kUtv/3XW3UzwmVPIde6Vpb0nBdhcc0SZCz/p26xS
SBTwO1UWMRTDcg39oG7wLDXG8sARBGJ5bOlxux6Dd0TZJOgWKDvKkdivRp5W9Varj7iWBbHtDl0/
9tTb4PeRLX6PXAu073HCmQAU7yQmhNU/9PH6Qfr6/kxl/ovY3UGD5x+228Cv61Gla1NM1qTvqbZ/
E2gAC3EYtjpGCv45MPPj7T8k4Uask5Fbum8qwjQyBuFCr5iSYiWhByTfaUm6qR6lIqxx3DnVc7Gr
V1Je7f9oeCdefhmFrPnYfLLBTj9I0yHiZs774PxBqfeSo5Xkr3UyIjqDBMYa70eQIWFaTNsyB2lA
Wd4V6Ryj3oQTmRzz8wB28ELRCQh8nCBxj3dZemU9yKELU6rPr6V69Y2uPmoCR4Bv3VsgIs8ZV2Uk
1rCW5Y0sCcufLwEU3dXOxFQbOXmg3/qo3GD3IlEf4nsy/0zHmCZaqSt4hLZ80+AcBRUgcXT4aFye
6E/JSBaB4iFYMUjfqWgQqNxKcx+PJm0SsJgNGSc3Zrfa+0XyYxEzY000g71AJ7a3DMuq3le1e+k0
+mhmK4vyOhKkonFrtRdxKDRDt0T7f4qEjwZcotPC+BFPBqZQQ8b51myNvZmrjK4kw9JfE3tiCw02
Dl32ElLBg1O3DJmmU+Emyvk/eGnRsl9kau6RdBul4cy4TUsEG4kH09TgnfKuaftAcbwgHm954xnv
PEZjfl953sJrcD0dbAI9VXcMqJfCMgl4K4WjeRthKPweTBN/+7FXezvhtAIcu1GjmCtHzBiF5vw7
9w8RWceR8oRrPF6Xb7nRDGPdIZmPLJPB3qes3y9zftWl3SUXsFMyfhMdQEDGNqbgmLFTZs2iJ/Qg
nuRoNii5Ouiqkq6T27fTbONkFRrZqGEWjMtQbx92febXbxq7QDHtGyikOou7J7+GDK+/ra4qqw6B
Sq6rM/Uv0UqwBTebRu/Qs30pcnMLIAeniOeAUaHQwjSprOBLOzZN6z7CB9HktfdsEIK2cHwWsk3o
JfV6tGiLK8JQGYxDTP9AIN7Pu088Oc8guXf5Cqu4ZBjM0U0jc5PnlS4QwZKK+VQIxiBrm3tNcBUG
PkeM4rVWuyJIGemHkKVqFj1LKZgwYi8Qqsab8GoWhat1auUwBd76YqD8nR75MciUEOVieflKq5IZ
AQ3pxA/qeIL3odwJUHAqJOMlK2hmVn+IJ9MGXpWLanp61ibrq8eKgyUPN0slRp+w6ezxmsOqB+bX
0C+69zmN98Nh8utby5CYpLyc8XiDM5lBzgdhjEVDjJBR8lTbhfJN0oMjdH+XrdiRQqwzVTV0zaxJ
/ak/wWze2ZpdJVYzZqHr3Tcu3EHFUg/1sVmBfhzfodcs+bHCzF+Q2yi/dnuvMJU/x7uhTF08tPo/
/qjsbILWYclJw01GabRTE+FIiafpRX1kbvaQSB8NvaOh0I2/A3mMDTz5zstI7RtxeQ7J62qx0rXr
IBOgA+qaCjMuMX056g2MeKqJldffHP2lWgTiwLwBqSbckJ3qJ1sor/3K2jSzVTIbHN6YXoxWpoDh
LWutdtL3ywXKnS3G+sh/STD3hNOK9AKKC1qMt0XiiJPOPMzll+wkA2BaxcVGbYb51aimMJVATzWq
Y77OWhy2mYkdwW8GbItAxgoajyHLBqRnrYQrr0IVuiulbDxSMoa9SwwbV8x7WF6o+Iil71QWR0qL
2lS5TuoG7z1dpqeQMQ4tuH8C8pv3x0OHKlMEP9Xe1q5Y3Viv8dpmrv7y0iIbz+RCENoLv8oMGVeM
SD4DoVVrahv6eArzC7kdO/Ad9dVnNhGaZ019REnieXTr7dKcgAlZ8+hFF/CHzPB3wNxMrXga2qhg
S2OO88Etw+5xM4+sRP8R4te0hL3D5Y6ORdzOANxC6Ho1VSKGAPF5eYr1qoSHYIHUJjzYl25kDIMf
w1ybj7WuTPkrf3tG7YjgAukqAjB0msVBq5OKgQtqvztBb34NSoPyZuevX9pYBJaTg/7eQWp5w6EA
f6DEk7V4ZYEGp9H/QBkxj2BvJ8csbiGYKhNnL0Kcb7es6Kwz2t5dxD0N0B20U1TTWZ7e4Uw96pPk
21kBN9v1KOleaseKPtlkw6fW82JECTM9F69/gmD3C9hjhq86fyLyksd+B8hEV4UpzQ8WSj1GGAVs
d6kGdIqFAQJNVGY27L8YLuC18y3wHM7yg+PcKCOoOboC9K3ODfJd3ttuTj7EdbpxnU5wkbGBG8ke
cOHM/jvcE7lRWZFpXv882RKFcE54TUoRuXW3dYcCWEaso7C7W9bV9ere9OCu1AaIf+QJvhrxGc0U
66sKEE+YFJcial+YCvd1GIyLFguntHLT46i2zoFvte4UC/1IQghn9Ezd+4BXMdpGNWt8l15fdFmd
AL0GHlxgKwMs/765294CAHrX/6VmeynkMpjW/itDIi5VM13/uD5L5A2GULOmppBssDYaM8q7lC+f
4/Iko3glOwz8DETOhu655wzfZXtx+rhnf4WEP6sZPs5AxtErhYEpgay2bQ64ijcjUgdKkVeA2dvV
8krAgMx2iDq2ks1iSMvchtxspHBCxQXbMWnrVI8ki162Cu6YnIl/RJntLxtZF4S9tgH9WdW2dQyG
dQAcPnSAIkPuyECQg0LPjy4x9MukQ/6FspKx6HEjgRHhuM9QDdM6HLz9Q2SFJCYRTRBfVAZZMaTf
92g4qwP7hMeOXrQkEc1v7D3TDsQu65S7pT/DODvOjUYQmv5sS1K0eoe69NHKDSoBn03Do81NmTb1
pcLy1+bNhCjWH2Okvu69mmSktRU+uiP9wdy5ri1iEjMclddE25uBEJ2OV0fllNU+sXB5zaJX7Bb1
lsenm7ydG1Lyv/iQ5EEb1P9ln45NgXuYYJBsTnTggRXcdOfQ5i3UwXdkpvdnsAsG0OcrDwu1tUxN
e1BKUuzn1UNkkgPiVjr1sBQpNuGEnPGEaBLfbEE9ACJNad1XVLvS76tONkcDtrh9IJcYH2LXHmKh
OYxPh61ZuFieaen1pBu1hABn+C6qpj0tdUZ10iRqtdXJc6xQiNDD9y4WY509lixzThQEBbL4rQrU
5sKuUuPbdb5ALiNktwdH9LxO9TQ5VoXt4s8kYlsVOf/LIkv4ftBElCxxUBjxYQAUq41/yFjIdV4s
ogFqWTNYLCV1BtOGe9Zb1GBCYUK8N6omVRQFKgd4S5vkkpjTgxU7Hw8gdmf8jH88ZX/6kLRZk1Pq
Yk4BZlispmnT/Dr2i5zf4qKZ0whaWFIs/TJKWO4knYZhrntcMipgutsipGqSMHEa+/31bC++GYcV
pRyP/fLL2oLppm4RvioxQ+tXTazT9Vhe5ba+PxeRkueTburzeXaVxHd6J1p+HivKk8X1mE268o7f
SkC0PzY1H+tJHrR4hoSo33wq8/qKZwR/45dC559/qclsP64PjjQ5AE5vsC+jhRfCWGid3z9U7YyH
zrQ9izrIVvu/olafa/lCDwlwYSXYVoOK8bqiQmR+kZ23L5fV7IoJExdHI2mGy53hVZmQet2aN4DE
Z3t2qRb09kHeBhb42akVvGRNf2Pj0sDM8gcfyHCxxK09e++2FX0oIWxPU51Bmcy8X5hpfxBYZLwy
3UQL2Nj6uYTk0sS3lAI8gBG3KOPol8p7GSjVUqwrWurYnEbjv0BhtkUurwcVTpgKY4DUfhuU+GiP
Xl5RPMDVKXYLZJ5y9w+vOah+9Orh1ZnRkuJAtCiUDNt6cCJ9oIBDLFz645515+Us4OtLuXV76Z9C
8gh4lhlz93BYun7q/GrUgpcWMRwAMt5fKTlcby57tRycBG405E3XxjwS3DMtlTx6EUa3OgYp4kWB
oxqKgYalEwJ4yd94xCkUJ4j1la5/acjHOUs3JtnCguHcbudpwplFbAhI9gnRlNaUD7GBThSr8gbT
lfivayXfka0c6b7STjcO5RtoW4uE16y97Cd/wxWhXNPaBuf8gdBu7QmvgWTcpk+XXM7pn204y6xi
Xnm+cKFgB/8KF8vyD4/y6lJnwXKKRcJQhBVZ6XAWY0Sx0tqUXPO0LRn/UXE7O4Us0M7yrmwc7z81
uabXPZH9Bx7g7vgRRfAD305JSsF+eVMeZ2lLKzU3mrwCkI7yvirXdXt2DRnYjfzZ/mJyp3iJrXTF
fWuBhC/oBoaTQRtJo3U9Vv1qfZG1MhoO/UfmJooIz+VO7jcffvieOHMQf3VkwdYPWGIF8YK0FwTi
T1HaFKHFKBsoZX0rBV7IDWDjTlJOYKX2mo+Oh5gI7SpWZLepa63Eps/LD5hEBZZyL0fK4yjhHkBV
LiRXbRk0gkeMh+s+s/OdInhyCm9DyLhNq+M4lbeorRBTDcr+wCKnc9yidHorb4XEOKKKFdNnFK/A
O4s5XIF/s5AyXbV08yacJHedPsK+J6JkozXnw4KmA0cnDc4UdEB/VUFiCiKJ3jRz6IC3x+icx1EH
qyc6TZSpMGwEdLHM+faAQ1q/yLN9BQMyabb1PTejx7fvdzJpCk3I61b4WI095trpHuQw29aXjdhw
lW2o/EY8fd8Reu/UiR06cpWxZJ6eqapUKUq+b63FvNSC0qKewL2uUNpSUf0Naos+y09tLrOlzQRh
Z1BBAz5GSGzLiMkyNS3tx7S/Jvw+Y0IBM1TFMbNmk2Tr8cAD5M9FS8xYZAuNPcSxNwldOitqT8CL
FGnHRiqX/lB4U43Zhmbq3AmbZxWbjjeRQzH6G50RQWKMBd3bwaOBJ6rBCCBMuvV93Xy46sTTM8ge
3CcslT70yM6nP1SW8VfDOt+xTGxabrgQZ9eraLVB+XIy4E5g1D+DWWCtvzFLQLSOb77QVJm4qi8s
7ZlyGO4tRO3ISUqWLpnvrDDkwRYNgHcB/RTYSo+MeAADvCBFY/vdNlYVTcukFUD53IiW7PddzGbK
YEHQdNFtCcOQhtpt7THHZ4zKasXIVeHC8bspBs6CIPtOw+qHyG7DImzw8FtOV1CPDY2+mIRNcqR0
qP/EBizb3UoeEVrYVKOCyiAvm3/JE7fwZhHH33wj3JIDQtfENOWnn/xp53xznqwSaXfy1DMmswiL
OojZBP7r7sFEu6XAYsORVInIW/iuxKM2j66DtJSqS0eBc3ZkwX7M+RKlnGtEoDnp3uICB5CWULfN
efLxjHkmHO6aHMN0EBkYJPsRZeywWqD5KgU9vHK04am0y2g/Y06hBpAVtRD7xjj6Igrmd33zJTrH
SgdvI/G8+XA9pU99556zUt/MgdMHgwh+Yw3K076Vbxg2PYu4zsKnXzAfWUuRO+uvSFrT1kbnM2fg
N8oKy4fQNzf1xa2lCyoD0oHHr8LhE9m/jq3f4I8WlMGtgA65gzFfDpTBSd4BLj9oEyT9MYsNEkYZ
CeBv/4sLHmaoXK2KavrGCvuv1evAkzm7DtxUzn788LTxPvsCS8iMLlbXBeLN05AuZofR1pmctv7I
JOWNuG+Eno17RQSPOrrSNYt2CpU5/wuGAoKq34Sb79qUbsIYGcWhrUzYKsrAxgkFTa+5oCcQuMyy
ueG6tdFCWNTDmCF5zgoF2YfLJJrVNJ1lFQ3eiDDO0OWOgYG7LT4KGxXz6NmcvsCwv/eE1/jNumtW
k1ex8nqGB4sz7HoL6FvWWm1s2vEscNR5k47Y3DspDsQMQWuBRxu4Ee+WkaJxXdcvzI5wxTNv3SPY
tw/ncCVzEDTqB+Eq+o3qXbVvegwx4OLj6XnKmBfcyKsMSbanSbALRCjQ0mjKW13okKzUmP7l0Wq8
T8+Lpsx3TEAtjscSrUQOkXIQETDs2dAprGVE0IttxXhBFHNKau0YKMOSpp8dBVHEl5+5VdRKcisR
FpPNtmqR6UlVt1rxbzCW0ozkGD27gH3u+xT6WpE1aNXwy9fLmRJbLobNo1hr3rXa+K4IpkD0qa71
cF/TLHekMxd7vKmrhF720ULka8oErbxBHxEB52or8mRRnjv9PTH5vmz5AuwJnT+mxmQctSAsVO/A
Ap3HizBVgStG1m87AlSUeD5u7/cO85yjGXRB2Odndk5wUHqUjVEW3+G2/36l3W4Y+WJ836udj0/3
HDJXd8n8TAPMB5QU4epo/HHhHFwgQ0KayidfE5o1uz3xH+cVY630rhtYkziEBPxGTDbxeMKHfxOx
kLKjaV5oB10cy1mAX8BVAge53zoJGi6CYo48pE9uoy+Jh6IYAGDyPBO+rOWWUbPTUtZ0OzRpOAjM
BPJv0lsZb9Haij6wBdh+v/riQvg9BRZtA7fgDualKkwOCB1zwHhxx+2QP12CAnEo/eUV21Q/wZb4
5sOS/53cJM6YrqdzwEivUKaJvsk6XmQ4CXE/CXVNc0Kt9e54/xisRDGPl9DGHPjoOWDdxpMkD9a0
5cuukkEYblIFEJPlNG4tXUp9XrujWFdlHTztTFwXDpSdtmbEZpe4N9zq+72BYMVYxtqpvf6qnrJy
xIxoP7mWcb0mDar7f/J74LI6vsCl1uML1DPJi+AnfGHCGRP66Rct85bDIWr6ROtZ+Pz0trLTQ/2F
+BAZBALk9bxh5FQeb2rmRBQKK8e8b4hB5o4rJpo4NLr8jk7+Dh9mRos0sWAA9hHfdURQ4RlG+/qT
/jpXfnNaArYe7jBOY1OW4E7VMEjGwpmv2VnR8JRffz6n1z/cYK47mvKGEzC0m9kqLLH51azF3K+/
TW4SoZJxFDipufGo9ozHO9V3xc8JfyxPg0n4Y8yueSuVYF6k///cVBz55LXTbz4tWt3AP4ZUhXPk
b95Y5ZGXmVK9AP0Dp/9/9wFtiJxUgqhKzNWXLImxih2iMp2vQAU5B88hEgv/k7gQcLrrPzpNzqqW
EAIMdaWiUmVazaLIZCMNdgSmg9ZA1+lsRaYxfrdUyqfVkq9bghyB+JBcZ2wwe1r/zjMeAN2ChDlc
C/mN8sw/dsd76lDza0buIPmLjKPobI4s8K1WXYk4qbLO9A6n94fbXMP3bcsbQe7AN27pyd4PEM++
z3hFkZ0WBmuhDnZltFPylfrbTpBCV7dJ9wFNL0dDctb80R+7TdrecZHhaKgcqMiSN5uoJu7tz9wR
osTfk6/ngKSlGQA29tcAtFPyKztaOgdtww7ORy2vuenQrS9j9X17ABW6SRKed4wCjKZ4MO69W4p4
6zZG2q8roqMdHAZH6+gCSY1PuPgKWQesB0Czwj0lBEHazrUhJs1KSwpLFVbIyj6kR2rADvPlPIuM
qziQm2FD7mt54R3FLv6wkq6dPnHXo/HPjiqNR8dxIpU3qVSjJJ8ybcEw4qOMVdttkZZsxfPVkhZf
D/l9wm2cDoqh9xqZkXKcHyzXgOCi69sQHKm3yLBjcMTPQAMzhEyAlDeBcJ5ZE4IJBt3Jrd3QfqBq
tuZP9THe8Z8CVfPzYP9Iuu+aXiK2hjPBzvyIiUVe1GUROYIE+JGeLaoiPVJw7AlGE/0LKsAoaQln
ziVec8ObkU7FzX+3QwSzkhhxQjC92JGIkaA4LLX3iEG4DxGo5BQNAsoHwkeslJ+KUlHfy1aol24/
x2izdEPDP80PLYKl8CRZq/ngHXC5F3j7CEFGC5DL6j/OsQIJRovp7sKDrw1wO0W0CRvrD8HK0Per
9EeeKv9P4BOJbbdMds1GAsu/pwpZ1ECrTtGeuj80HGKed1e4Bz8Yz0X9kPMXAHN+D9/RIBdiIHJL
f4VHyzITqMiXZmwb2U3vLyhzQ2qqRIwvSDb3hTJ6AOdFEnCm/LvhIx20/Df3bINR7aM/Kq6rl2vr
OZ7RfV8F8CNmSLv+sijU+jIY8LOztvQEhmWjG4I3LNMQCL2RYPmewisP709H4PAPaStv+JcJo67O
bfHcg/HWC9eogTOkKXLM0IYJhyZjymBDB0pirCqs/HWuX+lKUWMpMQYyn1WBuVwP6yKFnDEwNdr/
v1NoMm7zsI0sLOSHQP6emtPc5cRA1fFBMoMIWGWOzE27agYxbCpVfS5F3w9m99NVbHNj+ll4dn4N
VZ/rMssKx9UqHzrkxcIJY/yrse7G/q2iQkO+/fZUsYPuBrh3KnNa6skiKxWxBrkXvu664Bcs0dKa
FnX8evbGnBdrhybCsQ13/26HMmiewexmiu69npxwNVFrXv1G3DBl+hOzgl9fb6h4baKm5eG/0Zki
+cPvxtfqE4FP/PaCRCpPQlKX/mCfJXzRlo3V/Ivf9B/jy4zXkSmkvBFgCseaQYwowzR3sVu23cli
FU/ekHimELDsk0/b5GOyW1ngfGML6Q6Uy4tfz80pTOU1mcdJWHsjT/ZY1Mjq8Df+cCmGMKxc12w2
yYLzVF5IU/NIPG98QvmjM9lq8AUjBU5CFCQY1a73W7AB8c/awJdz9P0udbPiimOiUfZFeXFIf6T4
DuK273Kb2wKmKhgsnxltpGPcCjK7oOu6es/Y7welzmtzMTxVUVI9bnIOh91/4UQkq/Vwmq644k6j
sqLaYkpz5Lx/rrbwJ2zUID4CW8m5AC7Gypwh1XGm0uo2ZlGzzeC3wgHh7hsSJYUb4HbgYmukLusw
QsCrAn7Mt341qhGqwqZScK5CqMVqN+8OVsEdWkPlFHNcnGU6GOaEuFj5aOcuomCeAWcS3dbGxVrp
5g3KqkFPczvxEtFtoZ7h5yL6A0L1DeiOl7c2BfXGn/tv+fUz4x1/vSkC1PVRzI8j57GZpH32Xty6
phyRYnSUSiNk4BEJWgvublCA+LkW9eAiYx3koFTrTVXtQvCvnaRgjR5UUu2gDNMpHgARUhtGDSiA
1Zfrkaz+oEaUWbOXOmNOEf6seWu/BKQHtLt5ngcL28sP0ovJnhzMoco9vmVYiKi0tdEYzheNySLq
Q0TDUCGAxOStyOIHh3B7TRNo/wvJeVMXPFhhvBl+2kx8h+dxnjwzTMSgY+jlNMsDb50YyKySOSlK
BEcLagMBB63kdd2oFBpxJnEruSH1yv/qBWpyDvV8+eIKKMG+HupP08tTFOkHF6VgWkMiXe6bsSFC
Y8mj1t/HwU36hLlNmlCCWJeE0zM9gvnpcIOE9qLiHWn5LMg/rtQTN/Dzl7FiJ+QfwrSCTmhXB3qx
WxU4dpWsczj2SbnWGOO75Z8o2n9tDDdAJrKt84iudqJ3p2iNV0dE95PjKwLnhdMDIWxu7UkrXdZj
R06T2iMpQqWojVgRjuCVsiKCwDVSOkfL7BmFmrcAaMfHIENIAzA+CkpZmr5Tcxi0g8IJ2KZ4Y5H0
5nA/+tYuSQWN+c/UZ0QeElme49no1P4T2w5Oho2g0cvUu6XlHFii+/UsQRd+2aouUs8zRYtRvMi8
91rhXT7SheOybdZhzGc0rm+YM4ANccAU90tP9U1cfm4ho4wuO+ArNk/+H6B7tOvc6tl/JHNyBaLb
lMIfqbM1/O8pw0L4XoKPM79cmDxXuYb3mNS6C/qCUKolwywR8uLznBR9c7qgBR2zLbqLyJj1hsXf
MCGuTgpedC7GPxHurtYkzD5JtvDU1gzvlasmVfx/FJZg0TCbOzZJ4O/SrCbTxh5DZBalWvDV2VQV
6e7VWyu8SvTpE4GPZ+5hZ5e25MFSjHEelwM46INhfBDaQAh8jsQxKoMlWKWYHFLtVYE52woW0FZM
SbyYnC2pIzUu+1o35m10JTdSnzLbFuLOOhloshclRK6CTb6Ls4irTwHIcQnUgUU9e2LZxzovBaBi
UuoIGY2w5ze6B2oRbymvnL/FMe0mOYKBhLEiiAHSljqmkzLtfzXL/OObcBLSpB2poGymxNQBC7UZ
t5+1JFBFQjYVy253yUv8bqZUwFJ6lzPpvumNm5OdtuUVY79K0p66NJeIHHi2Oa80LhP8ZXuARmwq
+wvWyIqFB8EHUYLN8/zhLeH4LG7kyPerzpq0O64eGGcT7Xy0fnUSCVWg04aXcs3NvT1cKaffYZpg
E6s/qJ57Dm+cyLQZDiS21FGQ7s81l9GrAxQnusn5tYR7HiXlTxuBYfjml0LGd907p0+eEgSnp4/+
/GSt1y6Cl11a3eLbFOVkqtWftZ2/hatHjQyCF1Zamp/Fy5EyZBcNgW5gJ10XDe+BNx9FUlmuaRgV
t56V0NrzWXTaet+fXOkqzwfgDZO0rms93sl5zlvQf58ExwijZg6PFve7BpCJwUVxqPmBM5wbh+8s
QIFtpQzx+18DuKQHrx3aW4+/0dqPUquerSqVu7OnrscsaBgnBzRj9kdPLiUkWJmGETpexOjm3BSU
ayV87/iDKBTUmcM5QRfZCj7/H+GPYzRSo/CLySe0EgiDM2fIV7kS/vlUbULHz4GBMzADfqf4/4dS
bETgS1+hYE41zhg8JdAWYeqNrGAeH67chIJ8qC0wEe60ZxVZerm5DhumLZYnwL0gCLaBEd40IsDD
BWqauJxjh5OiZpRl6x1T+cTSfch0C2Gx/w4hZPHRE4SAifnIViRF30YOl+RHn2VwL5C5tZZDN15o
dnJgso9uKYtmLtyUjiObegzJcRGHp7bMdDpD7YXkHIeTKzAB+3iSAhfnFEqHJmHbKdtaWqkz/Ytu
PxOZ7nVyi6kMwmlSjE01Y5CzEexSeY5SehWen7zCGPakPJ4qNltkt8mNKkvDkZRlFPnFPUQhPzwP
4UXS0FLfTSbSw2xclTWjoc4Qi4NboOK++tIqcgywSAXejbikV7JeUfrqmv3UpjpxKEGTb/UvNpJq
QtvR1z3LS4RynXwd+sffUbNmY+AVlUk5nV3Zm0azPUba/4oEV9JWF83j/JB06inQGg/x2crUDGjo
iKFTe56pgRZI3PJ3/4pglfx6977DqeOwUj8hsQUCIEyMKS3DgtdQUdXSQBAnRxxGZQ/4sgg2jvSe
t+cW67IcrTAGagk9oCTrFwoEvmquAaqVsQiJ71n0CZOT7Tlz+7FDHd9ut5B3gqkJ3Tk7jjKZiRHe
KQeHZEvXgQfzETiuAZKZIzLSF6G6wejnhmzJDDTTRSxqB3WbnlvULA3ZlBiVM0yn7PiP4ZDeR1ey
9OD/LblGTa0iFARWdv6lkxmJMfowKqB4DD8NZVdpJkczR9y7jd0QxgUcG5LGOtzJ5ffuxTsAtyL1
eAjg0ZvWegv0FOY5rPV0BdD+VwCfLUdvTe3UnZblKnE67BFz1cLzD9H9qkBzpPyxPrSIMRY1rvJB
tRKrGtLp2JZuNQQaYO/1zdU0GvpJND1dbctHNYq2CQ+E8+wDGqlP9Qsu3gpuMlvFZHpsqXpsic9b
fvd+Fnlw3n34V4V3p/jRjTFPGSgf/563tFcW1yG+1nNg0QYFTgdt8U6ndzGMRoydqsCNGsRTbvT+
ajHWe1ObxdC7mJpyZmGjK277Afp2FzeOV61BPAhwBKO8cZyERsgicQpKz+bw6NJHxepqzQK6af4x
TG1sMKWHtjp3ZjLVSA1r4lhSiuRVE+nZ71fwRhY5x0irp9aN/NZOjtuXtKb2Hl6NQQUaXsEvaahT
o+Qp9HBl970GsalKxbEeFlnE6b7lQcxN3yVE72eh3hgfdkPP9Kpd45JhdPqaH5zCNCT2uMSjdiLI
pRkYHkeMHkQ94fVruqiWWSF1r73aX2bg5p3zQqg1DcQvFwrlJep9dxz5N7kRFFn1KmOEJ/NHbb4M
2aFAcsNq9psD9sqY7yiorjp6xsyFXyLHWGioAJHw8G1ilHY+yJPVFPQICu0mWKJs1ekrVB8zwH7O
lJ6EHzdPtVIH23CZRYR96Ddc+tnUg4sZ474wWYfUkrdp/hXiUUDbwbneMeTRH6Gbx2dNkYXrLfDc
AX8hQSSjMotHKCiNMaHdKmAl/3CCLC7cMtfCif6HPWtjZHR0ymPsob42j++vfepuF3m+McmLhwYy
P3UH7RhG0FAUDVEhBNX1oYrH7lbUSPN0CPEDiFk/O7vs7xZAk681WtFvXGz1OM4z3fCHVQHRCfDs
KPwN1twACtKwpw+ftp3G27o7E4N3Fxob3enmfyX7Rxwsx/bugrBouWTWE54pwPaM7Xs0UpT/E/QH
0uwBW6+WUglqkj7OvtCximdtl35KJYpErbPf0Z71vuGdJBsmlCVcYdUD5cDMKps7DNk9xUzmz3zv
iNMgTFrlcgoqxcs0Xw+uxb3fgZWnzaCJk5RW2jHgEDeulX+h8ZkDAPh0PNnFNKi7UfdJisVuUoVe
vxLBzfkNBg7ri+/AbkuZk1FSOQAfO/fxl6DGs4V5zawqhURb+BHruridx+ledgREFAMNRpM7kE7n
E0C3ugVV1AzxrRzeF9sPaUUrZflmekTSsNy/Tc8Lx/bxNQ6s3+lFXtFQEZ06Ykz6aznynQRYhAYM
rcjXdvXo6TxV5C1MSy5nxIJdxlqPdi0xN3iAAnThFH/bYzVCWdjPadBMM7uDxIKbcuZeCyH6ulgf
MDVQjSv7n7vyq2gHo1RUqlonHa343Uj57KRYrmUFX1M78tU9zu0BwDz4RormgjNxUqCyL3G6yAel
GUoMWc5j9bRXFnwgRit8QYawQAeG/CUnVm33ZdfDlaib7dBR3GcLgoUfwAJzGNvHHUm6bKXhgGjI
d/umkzlHfsXtBB9LgHaCM4e2AtyfVeqHARn9wsnYgVFy8dPex0GcdcH5qisF7DnJ1l7GDWRIV8Ak
L3WSEvjFNguVoXaH7z68tM5oWYnVozpN+oIkw87MoD55gxqwBdCieP7xSs2pltH1t+GjvC87YIA0
fKMOJ+EWPH/MQHFqo0WUBcfqaaTr7yMR43DgPU5mJOmaYsxm2lI6pJG+PVbMcWWRZ6GLiCXQJ12m
W56n2v6HYZjuiv5bfWfhQIYRyOIzpV3tQQY7l/UJ1olTDF0mHfWCnmQ6NcxSRndHw/mbzD6ySOm7
fY1aww20wDaFsulml5X8UtjW9PTyFEfESYyrSkkW3qQ2gAqveOlRS01JA6D0oaVb3c3lTTHLYrrx
w3l9vb28t8eRWk3vuEcR8jzgvTLjq8IQzr5uSop3GsP9FDSYgsgSdxAivmykWA2bM9l6PrtUB/tN
lO9dGihOM1GthO6GYq8/tpOLFBPawfm3DaZZbfij3f1le2B1YZWvu0H4PZ18WRliKXIIpRqoitf+
1cXJ406WosFE25maKaOGGeYb0kY3AVCrCYacH466UYIU+whOELKbElpyiA4nRLGcD+905vzqUmBg
iUbv7TNy1SBpaRnJVi6QpUX9gpoHliikUFfHZmoI7W+tL1+uG3yUU7yU1CU5Xge3o4gZbpk0hk+H
Z7dZEQBMDyJjaObn2AVgn0LGUfcfyISid8/fqxQwBLBg5NwGHTno3liPVYNmmpFbltkHxPBU6+sz
w73pffg1zYe1Ps/r1c6euClFef8xw/3wyoYhjkdISmsMC7EmdVgKamDbZ9F6Zm4vCVu/jVk41PPA
66RJgcEv/mqIdam7Tq9eU7QeY7Go6nN19JcjpRNLFrRqjrx+Bv0uM8TPKWfcK/Ngodv7HWHhS3pf
M0fANIhO2CTDeEcTQb3AE21+Cd6wTVhj/1Wwa/J9EPNzN89yM2r9KIoYzSTTwkl7zLO+w7POZK8C
YL55E9/GTMerUOZ09ZwTflDwgz17j6az6Afe/TjArtoBF6+KhExvgRen2NcSFLvM5yUr9CDCLdwO
+czlZ0k6viIHu4Hs6He5bjVW8Mm5uUgRZ0nWH9/wKNI2GodKyqZ+dPrT/ujCMpOEHndYdmfoZZIO
77lHif2PnXGxDVwRYl+deXwPno3mBZwL4dcPibr//C2nTatUZmYvXjMiiSqotW0xYUkYUzQfAYxh
GrSa00LYD2LUS/vte6ak4Im2v6vzchOIShHDNc/PJxYWGBy35cutNzFu65Boy4s40BzspGpRrdny
e6lnr7Mav5NYY+hc7BGSqJT8fqF4yXZlg/AntXCT1vj5hlVluJ+6qFqabMWLo0mnNnbMUF3jPCzu
7N0NI8r20aCUBoWiPW4AauE5zNgyZAmobWy9J/YRDEcg+/88vHQxk/hhel4VnVBGAwgAS3G7f7dt
T7YSFRSQXYJXC20Ym6rvf2hist1huU8SEg/a5EI1XGkzfDqpDaslZAJDlWp9aaqgq0kgwaf207hz
yNF2sAFC3Z8YMlfv0eYkHJ16nIZMXET8bx0Hl4KOkUU1J8QwjMa1C+djGLYzjHj0TfjxkVeCiFgf
7cMcsfwa85RB1gpfzeWviBtZU0+tZSUr7NFAReSN+qk9xXmul2Bn0GfipB56Ophfj1yRMvqiLAwX
mwy5zZXr0XenVzRuc1vjRDnrm2e9g4zkic+p8GOvU5kDqAIlMr25RQYsubUI8LrgtGwUuX9AZnU1
MGi73F7hgMbN0LqV2RlJmku1y5XR7zShsWG6gHxMXXnCy2vpEmDGZYlHJS37jqpmhQQUQfZa54mL
2Yv12SkTlZk88o9dG10I3XiH0hEAV1fLXSFeYoVur5p+GVTImCV+zXOfjh7o5wjYFt/t6XuB+pBp
/s40nuFTkuyNXFn3553tbM6Jyo9fOy7+4skOipHAb7rcstv5hoN6hemMvZq61L9sRQhPsbDlmwJs
noEFP/BJoLWLQwi5IhtjCU94naboMGJCGj+lEgBKDBEljvCuQPPpxlTonCU9AvJE6QtO/xgevm5A
R+sf39sSv3x+BmfRW6d/V8XqsHaK9q3nDPZ2k9IVyMXLMf6gnsYMIOwY6ZVuBCSavZwpbf3rtV1l
1hXC/r8FXpZKf7IZhSiOTrX5LM07Dl+op37t1m2DsN0cgS+C2+DIFB2o1st6p6361le2F3kYNbFE
uKviUHzmQm304QrUtdDAmxfnNOIbC+b06fjaJtO3qABPHz5nYlVPi1La3999W1ngie0M/4eJKZY3
NFQzy3C06X+ZFaQ1RH5SXu6l08TmjJYo2D9tQ9WKqfup34Rv+D6id4MH1gAx/JO1QOSPG7Nrkgbh
jQgMVq+kXulcKFe0EkgOtx2g3baOphx5VS7dul9Icml9fvjpBfRUVfogQvZ/NjEoCqm8K8yl2sFj
wLmcVdP4aIMJe8m2AA2uBisSS7VvK4ak9+Spn5iMAfw1/ev3jZgxWxHNxpyRbP9xoMiBCvWoX0Vw
bp2YsskOgxOn24mFQgw63OyIXFQQ8ZNJwXBzY5e5+IEIUtFT+oa+cMQi9b8dbilhRwcfM2h4cQMV
xZkWA2bRloGzKqvFAEc0nIqdztFeP5Il03Wd6mPiPR8K/s1QBCafQw09H39jg9++jqpgJFhW7NMh
/AmpdyypQJ/JurSdtmWdFA7B0Lq8xLmBSIMCjukmU2d7QCnOPBogpy9pz/1bE13ymKKc0ulPkg8G
grm26cYIR9ytblTCY41dhBG6jrVgG0se2dZ25gZ4+IbTdkXXREtlFro1VZMfCLJVahBN5RrrH/pm
/d1JbPrbsE7lJvGMj1lCdszWPl3cI+xsw3Am/q20dc/jFvQpiQHeBa3HeCd6CNFZaHkrmlpup2Nt
gv/e4Os8bGTy2+yGXk3NVxB7KqvO7JHteuTLtO+G4GdiTEH9XAXwoEAAspOD+8RaWRxWejyNoBNC
1VJAwVwkPgaoFts7R6gE64BQX3JcfdSpi3TcoLaRaY3JfXsfWaKP1h16wnUgAqg2TZOaVBaO7pvF
J3cAIIDMHTmBsxlBVIHKt2ZWh22taw+Mw5V92CTurXHlP/8PlCn3mUwpG0wS1jxlzRqyQh7Q2+7z
/03WpSsBdogbjhMS56qE37UUqGt9Erz1rMTWXpGfSKYN4mDYrgi12xMKRK9p1B5TGWINsqEzGlrs
B9G+ZnUxWpYdC3dqWKA5vb70EgI3eMx71gSl7BtXvrOtJMnFUo0FB/qzjvMGGshah86MlJhTkIed
2BSzQjHgYT98swVN2FvYErnYZFN5tFEDmxZai5uDz1dZ8r86GHUNFSX+MWNvFPritV242tif5ACK
ObdaolsdAWL4FoRslQ22EASURmyAsjhKzBt4nPmgcSI2pV8LQAdBZM5lJEdyMVlBTmOk0UrIjIf/
TqY1DCJx2EVTzSaB9LeEcWhqqxTkl6JJMM47trETCjAr//zheUigaJM3R4+ylI3ThiKNTkaTzpdU
/W3XBxkiHh3qj6PzqqNxL5vNOL/y/obQa7NVebW8wQ2cFM+DygpbmYWZsXUyJDspfu5fRATesmr5
Al4NPKLAO4i9v9Bj5UBrsnMy/jGsaQ2cTAp/gq8cAHQDmZ7Nv7f9/G2y0WuLHCSPGv1nk63KxUTX
0EXXMw78Gh7WjygNIyQfb75STKg/jCO/g6atsUnK4xq1KBYbm5MKLD0JV5XY+GxmTuJYRU8FxvfK
Czn2+SLMrjI1i+f4vSY1VFPsRX0pif1fFK6FMfllMzawgYPioJD9TnoK2m5gIG34Qg/eL/xPDMEJ
tp+8eio6l1Xt9Wg0Xex5siOmzEKB05Ds7kGAcIJvVrR5xNM1FAqVICsz/e+vG54pd1PNeaQusNIg
+UxcC0GoMB4vtusKSjGxjCBwC6v/E1WzrunV2AJegQwg4moh//z553CkQcrXcMu02nViZwutvxdH
X7uj4QNBCZzZVFq3s3YCfLvYulDGwjlmogwYfyWuPX9fWy2ms6nX/nvD5ewqOA892x5ytxKZ5R9U
75U9x13hsKsVJzdkp4p6Ig33HOqRCPSNJ/k1RgBmRFTApFmKIgfjgkISN95rlkEY0RxsarbJhnY7
qDp1ozAm79bD87wJhlgLbnmDQ5ruSTno7q5idqtvP6+6R/Tqdn6vsRuC+oc7EInrUfVXlTV01Io/
OFqwoMWGC7pIW+tsPKZxV54qHravx6kSHXboifXe3bd9B6nZPBejs2nkvhmLMx0YUWc1epmS/QX3
/PzuhHllBf0M/rX/EBwKW5iwd6r73HdeSz4cbu3hg/SI35bFhwQQhd4nm5IK/RNSk/m4K7z+Fldb
6iFQIccNbByWx8KEKC3h9tZYiHnHhK5ymRB6Pd4OEtuZ7GKPyu4SA+ckKp3R6S+oiWGSYMtufAY8
oMb2xcJseNDdkhEBdALXEAmlIXFCC3sB9d6prETiFuM7U0wNvU5gjjhUjJ2E5jmz05h7zyNdy+S5
Lc07Pg3Zr5hLYDnA2bI5LVNVfbhuwNDKc9Y63yZSEXGMsVh+ILkgxAoMaLV6gLxEE78WhcFrRlyz
ozEWYkGg5O5gTB32tD7YrJHoA1lvEwXtcNz8uqRZbPw947lJ8aFSDnFac+SaeEi+oRR1+klt+3XJ
ab//WrF+XaaevLVdFMiuwQJsDPPqzOEtdN2im5LzYfeU5R98gsW8zKZAcXOWzafK/38K+0nQwh1h
QWoR3m1+nCw6z0vToQSizH/FHFRJ6L5JDpgI2LVgcgfjaddgKZEOeuDi5L7c7xCeMFWwBiXgiC9/
hoySoZUeaI1upqh3o9pssinObkg44ZvAav2Lc0yG8KaNmYh4WAXzazyTkFn90z38/Eqytg78+gcJ
eVQjIQzyZ5MZ2Ow2iee9ZEMoxNzy7HbIfD2bmwy7jTdlMJPiAmwRECiZcfOZulTJ8MWrt8mq/OUK
P0yurWq9sLl07+yjSmsIRNftNPSoD79znp7aGCR1km70VWNdyZcL3KaNqCp7J1MeJslesz4siB6j
A2mqca9UTK6dsFVuKVx4BEw2AOkK6/sUlpJdDoTOcONnRJMKOkHl8BItHgn1nOw6W+e2Hq2Jwz02
4ogEWfYjVA5IdyOy6etHlUDOKMPRvrfn13mbP5gJ/msSUHQZYr1qM7HHVTeSXMR39xtbI0qESkwh
gGO8/Ee9svS5eCRJvFAWZoE3jjCQ2GxEmo2aJLFh590augrvEfy/2sViO0qpvp5YnN/zN06Q/0JN
E7KXVvMgVvZSlfuQbWUTu2pmmsE+eerXwiFl4+XpogqMHIa1OPO8wZupcqQY2e8hzzPX2hXcVpX2
hdOq6yPjTEwQS1U0NTSpg5m/X6HS36bRWa7j0zHZ104Mkpihm14Aye+u632Uwe1XG0iVIFqyAOTi
mi8F8jvUuT2+pMmrS1/RZRv0mmKobdbuNG/87pbt7kwcig6VkHh3VK1MNH+zF3Y8nwROoZ8S+5lC
LW76wpGi5dEDIcGYIhFIGo5ULCkHh+K+jzQq4+EM1u6PT1DvKdVhp84ESCjBp9DmRkgukLPwWvzJ
EwZv9slXBE1Dx9QMQ8GQzC72AuS++3bSnpkeYgTPHAx5h9muf7XJBQlxtIGKS37+uylfdxhhJD1b
n3r4mqDsnIqIPhRFCbXxzoPy+pVqtlsf2GlnTkYek7UkRYIHdBUhkbsWfpgJosq6+tlyk+ueuAe6
N/B7s5B9eyyw+Ejr+C7guZ96wPcDeRTbdpLdSl+9cYv3x9WUXBuPaZHQtOVS1e61KP8RPj4jKinG
Tdgh1vKCbjLRFJ4tM7j80lz3VFkWQI90petJ3kep5LIJvcnwxHJazFPcvBQpBQ5VhZQsDvaavVVi
Hu78sShNjLqziCsrSHIsCNH2jg2WsEhySOyl60s7P74HD9CbKWYeGReIqQJeRcOVsIGipWhFbU1o
swNLh3cavQY7o7l48tmjNwBAgOPvooI0bYjE3k79Z83bO/X102NILJEJR87ikMiJJg87AbBEAMp8
kG+mGrdhPRNtNqfhasz1SrwAFU3g6B+nQ8haGF6cvz1AQ2UE9TjBxLO4Z6F1JJrYYRJs0xU/TlN0
mNJ1FdD5eF5qPkl+MQu4FAgeTZG7jj5OBAgzzQ9uilLB7XD1STVQyNFjAzWGDLvV0GbkXHc1uqYb
LHQjNWr9qrI0X4s5gYNIVR2M+hjC83fIGNqMS3tZLup1zOtJPc55KwNg5qG6mh/SVDKsMPHJd98N
4Yui9/1IVpBlM4+Hk7O7Gyh/173Vv4/Se1cluQQl8SOZRlWlkvPjjY3maU+Mabyl7fht+u7P/wsI
C9h/MDQ+fJBKEq/FL9QxSmEWohSyZ8lKEUd9F9sPWoyVl++128qKZ1zBTJ8f4PfInXq+yZCoQM3s
OklllmiBLT/EtUKnkiM+w/IllFKFaPg4o7aJShpa3NS56EAJAHINnEchx+BRskdCcOGYyDuDFj7C
k9rBcpnsvGWqnGjXHj/pMWngn7DnYS1yRFIevipaIc8ga9XVO+MeJIF1rxfvDLmWW4XUUv1mUwe4
I6z4rGPYKQRnozmFlozSaLvufQglCiPoUQ7tNLJZLMHX3gILa6dPoBxz779hnZ2qsz0hGE6k1CMK
XHbVranw/hhLuJAN/eZkfTr1c99P0cAGiz1/Q7OQpCaHd3nUzZ5ynA7voKuFajxSuI5zyOXqPdEG
/oLTlGEAHnecm+0CbhbIpW/wrvFT83nReIH0S+2Lv2okWafTDR93X5D8yjY5/s8SBAXBNqSVMfxL
ZODW74LYXUlIEQruOErYHy2Lmpo9ij+vN8ogJs+WHMoHVqZ+0bujRm/O9XiMexEFaV/RpnX1w5rD
3Mnfs3Fojb514G5ICU30Fx3ilBbXhddw+QLW76wWP5z/wDMpvjqmxND7h7qRIQd9c2f2J6g/lf9g
66VKQAD4FJTm/2QAqd3UNrYoyjMz6BaXRQ9YzY8p5db/v2OlwRy8NHE+KlZ+HPT9b++xJAlz5Zc0
4RgSWuLxP8vBXXuGYuD2hAIc+x8GutPS5f9Y6t+Rds9Icnx3M1ldVbIj0d9iTd9caVaFE/VoRDkc
iL/AuFSzK/xLxH0FJPeUQVK+Fb5HazevG1f7+u8YE0CHVfdOmdpwgZBBWewcNk0C6UvmmkIAfZhy
kF3lMG40n0Z1QGU2zNyerWyhY+DgMm8K+Dxh8cf1WRirJsi9nQU48Vh/mBymsAiAREpkE90FPEIW
GdXjhdyyj9QbwDLrPYt7iyzf2rSF/4+HSNr6CGDMjEvcA7IEqA/W3ZP7h9oye0GMGFznq8WExiGL
UuXx1/xmhOAM9ZvvJW1x96SA88uOR/bUKtJo3KNRu+/giXCM7/zQ1gaB55AnD1LNctC7uhCFKMq0
VznOah6LhICrP+oLOM6vYZVLyDNCVKEjWpqEzlPWAwaXtNGKQ/xJzvpQPbi4hM8XGXEI9up15ee0
a4fU8QIbKGzRYoY3yUDcM1bwwfUA9p9YYKoWPw6g1GdzRSQzQ8datakVNHs1D9SUMO+8lKtf6Yth
x4CHLeI0Fv+5jmQEhtY4oIAqGMrkwYpQjX2TS+SF5M5Pkd8tDGHrEGj0OBT96k4QYdqc/WvqGmSN
GdKkjWzuSYX7/yOtlP/isQvQDcWyqINVX32yD1tUhguVfbXyzwiNUDyjlKLI0Kk475GWvN+xKaRX
35D2go2yfgsWLsPt55YeyrKQJhWuZp0ypazohSpEjhe7suI4mM4wyb7sinxGE3eSE1Ysb+i/HXjW
mHfQqt0MEx8XdwxEFhld/sIJl84icQfA/XARCi5rgi6M9NA//fkFVL89r2vfN+AUJWJSTonNtGSc
jaudWhGMb+R3wHMrgEKdq8yV6j9AYQ1Dcw2VUfon47NsYVLpVECbAl/gIn/EeizorjJRmH/2hKeD
4kPzGgK9EN+eqVCKJJL9jf4JSxIcYR7rYULszG0JCy/0VSStN3bd057TGYQrMN2LA42t92HhusEn
y/SUv0O505Np8Kmty4nGG/HS+kcVEv+B1HhZipRMHnlvXQ7RkbiBvgo9zqZIynUgvY2Gp1lvYxUP
WiKnXYrw+x2iLhqmhvsYQc+j/Y/JTuFYMxbO+U1NC1ie8TDzYfyLXRVu1oLYQZHyp22A4NzUWsN5
H4m/8ffAgUbYI/St8cocPfq5K6YDgx0VuddIDQXuol3qIeq36ODjq2LKhHqvDDMjpuZxEorygQL8
0gnNp4VtaK4aE2XXtSFX63UGJ6bx2h4yhL+hG2aY5d9vyD0RdivejlhplF4vl+EGsF0HaKhpnbhh
hfFM0In6xVL+bsZNl74kIwgcp5c5yCBLIjtJUhKbKLOpzi9yhss2y8dPA+mivnvA14RF4BL4wVwe
aQdWvRw0a9ODEINfiDmVlrUNC5ghz1AupHeN9MLZbE4J/VqpF1Os55zBHQWhBcJ+8QXinW0ptM2f
CQyA9xdAzp/MG/UQsErdSlZwX8Sw0N2c/aczYEaLju35WLeTaizq6m8QPrzyV0v0fRUfmyd3Ize8
hKftjBImxGfBjWK8S24zRu4ycxobNwJ7tfvllhavFMbgDVjNJ3lLVNgYgZvAce78V1wKqQNdnLvF
TjB1A0nRHWv99pvAO70V+VyMuhEM7XozPdCEnqD6aJGXGdoOKetLPj7O+/8jNQGN+id6TScJAsRu
tnyty7Xtl0tyyfnZbTe4L6Ngs62CMoeHfe/sNyeWQAVUPaSs3Iu6jOavNgIIS2P999cpYwLJXiDF
zofVts2J6cCQ2QwBaq2CnUhtLvnsYdZlrUKswMxyyYnfrvbGnB3ooFpcPW4F5o8qtAU6IVdlTPgw
jHZ+n227oet5cempA0c6a3OevnNuNdMBeBDhE8IBFB8pYI4iPJo0dhvCVC+u/u8HjMGbdWeEXhi5
NadjUT2ZYSPcUa8m3Feyg/9Xwp+vQnPSaE+FyWCJsDoWpcGHn1OusCzhRSGbCKQIA2jA6EV/nKgp
+OffxZlLhfftv2KFwn2jRtMqI2pn4u7e30t25DwN8I7PskThQb6K/cULqipsd+y610i3OGKbCE3g
Bc7hqQXltW9NVnLn/nRgjS7Lc1j0bcO1dKb0uV/4ALQYVgk7hVizLwQ72uSzUMrn8QePtrsV/Bb4
y+3h1tL+rhMNCJ0z3njNImgtrKlFQSkjLey/a9Gw5rQVgyCt2v3qHTz1ndWsbkfBLq9sZP+pMgxd
tNMdCKPYfFmfiQeZa3Yg7Nes0RyngVkPxuxqwY2sdJwaCAllvuxsm7lNKe826021jimrt/Z4Gu1c
QeWHVT9MWg7Jvh2bD6Ubq1yFx27e7+YZCBkuAqPIr/Ll7UsGLxVe20eR+aUZhu0KJ5tURn+XnxGu
CiJqEPmL4XlwPixeshwkybXDnUJ8+AtjLK4HxhdWTN7pimAOX2bfhV1tZnJ4DxYONi4Lge51kb1X
TYYIB91m0BokJNH15IgxTZwQBJW3NTJFkJQOk/ULbJXotSSYM1wuQ2RVO2scA/0ABICImSqH4Pyp
NmeqCZQZqpehbvCotXqPR6Y+kVuolqxltsMRae/aXnBbWwSSY+X+8nkIjPJ/hLKXL9M78XIANM8s
d4x3W73XVaft2A6tRsajx0FBoREE5TDePCZd+qoJRwRcNLxNc7muj/JJpcKX7qbQcnFaOo0KSUSx
XNkrPZF1pWhyYPK3CzGrOo8d0qaIGnlPDyyiIDhZntFoBrQbE9CVNf5tURJxFTyKZcvL1waHOi1g
8wXh8MJrOyN30Df89qslUd/OFpEbVpLoKSJhfgMjQ7P6zrIfAjZmEXKn15WjTr6KejVXvUqLjGOE
tWUMnJ81VcrwbjXpdeh1Frl9lInJB/BP9aHmTVrq6HP6dauEV/ky33XqxFulLWeO6Es+SbcGWEOD
amPkoU65DtDJ0PS+y1S8IH0yx/+BhwWKz25dh/FNXhixh95ddqc0hK6mAFOQV+XyCHw8viX0u2Wy
LZxG3Laa8gkA+gJiKImDj1gQp2hDGZCPeWA7vMCPoM+Y06UXfZwGvfwVlunDN5tkNsPUyxfOFeti
QdNB8CrZBCF/ApzoYF6OclozWbHN2+0/8Hiw9Oma9AmCdLyJiS0ZIMyFTjfvmyNOPjp2u+cL1oMg
rhq15u3CY9kL3Z26Rk9phAMszmOoLY93zp4Jy0pR4FC9yw5zJOcEYBSw+kz34c2M64NoT+wkmVjj
aW9YfKfZJfPyy1H/YMfwabcyB57g3HPpoTqragN01K1zgytqipFboNj+TV3z1j9/FQqHCtWT3vBh
wrePB+F3MGBEF7yB2BKjsD2KzhwBLDNP8zNR4pDj3+qwDRUlUWx7iMmshANODqNuJS/V86zsmR0n
UCQF+kRrARN5gTq/jjMG6v9cxvNnlsRF5gH+XlwvTKD43BcAKhbF1L8UdzUFUNGStJSYNPUnnc2f
5V76wGnvkXSozQcpJo7NZFD5o4rJ51CCBvqmkKU+hpjjkccAXXBC5ykt52TQHSNOmoPIwwEVliPC
5HfDYtSltnHuyXgXXT2T0+e7urcoYUVnbFYV+2pj+J1toijUZTtAJV8aVRl2c9iDCcl7msfpj8jS
CH0Q2MF+M2PrwhzA6YnaPiHY9CpAa/VE6/eOmb1frqhmZdpKitolc7YZUkaLghb3K5cTz+FF858R
h6AnnbZcJFVXxrLNcmBQh5xGL4TqvOJkKw9PuCHR7+Ov55kHETdEj7Ga7GejDvZHT0vvFYQNq7A2
FYa+2Fsixgdc6eu6VUbDVO6zhxLbi9J4QaclzHfmdqCk1arlteb/LfSUKDR/9irvgpfkL7i4EHeK
Kag0OC3GiEfWZfk3uEx9vxjgWhB6Uz7ZAbC2NAfTcge1YS9//Pr+xoUd0UNGsJ8m+NAVKM6xL9Q4
S42GkjCZEDWRm+h8q03ZdrDu+YU+Jxa+L1mA+mEPqLndM+c7AshAeXA2TaFEiJ4+5oaR8CS5OT/x
ew89iFq6obDCPm8m/wNQr9Qjzme0wPQhp0taO8Oxsi/lqoNpmPXqwzrnw4RCGmq8kUdQYc4mXUSe
pMq2xOjzKL/0DldFngKTMhfEGlZaDbeNaLdaLKjIgGp8vxJsjSGEE3ocHsclwVwyY+hYgI97+612
oP5DyT0PbWWdcrJm02Zbks0e0iFWQrkAYLbKRBRgWKufWlQ0Sgy/+B8HDbBJDmyWkd6qgXJqYLS/
aWlfYaRAbCmaAhbMtngJnQpusHc3RUdTVXB3LXcWGLp91BFVpKI/cGDY9FTSvsrTs/M0rqWFB8oA
di/H46Q4qS9CUPLBMwSesIV0mO4OF3MvFUzBAkiYx8wxVNBfdOElFF172MUtZsN5eDCC2EEl1jiX
PVK3rZmRIgz/AvdEkxY4ozJJ7VFkr4Nt0O4XgkaTpWosr976ueRe/PMfX/KLLEbYNPCuo6+kWdxB
dGGv+tvPj80YzjkGRRWq5iID1PhThsp/fiAIM8LGdqdahlwPdx7SrbvMIlMH+CAaCUO7BxHcoFw8
6jAiSkxfei2QzH3b5WVjvxaESwwtP7Rb7H07QUI+qDpEmSLCShtz6nYuohwoXAvJXBISwORCp/un
gLOVxKy4AmDMiJBk0WBDXqHezFjDbUY8gE+LQqHJ2DXH4QgHx/6Je8pCrcz6qrMRLqUmx3tdxfot
FFfprcYvhyl899YY49R5IF1Sh6LXF3q+J6MIlUFYKMHheSv2rLRiONquMVGxaW3v/9L1fBeRBuhe
y8yjMGcbcQqAoub+okTpN6/sIBWSXSx7K7y+06LFGLiETGib9r4+W+S3V3brNxzEx2HRr2G5DBEp
5Rz1eX4X74M9R564UeEZh/h8//FHlH9gWAnAQYP0J5LFYZ0sSPNDY1U0DAcBwayF1tMSMDX38ebM
Pf0aOmqRyHo2CqlN8HKE7vATzPaFUaM4hKwxLh0V3Y/WKJCUEZGgceRemOojWx8ekEaEyLZSrt58
UTW1B8NdUGe+lX07VKtUjdc40n/JiCa75wpLovWCfCZiTFY0MU3M+gxaRwxhaiJQ13MNEd7na10T
ii4gh1KQ+C8WHs07MyyHyaLpJIPdPBgGhznY9YdTB+d6MuFLND7c0Xmn16riqMV7UJ0prAGA1M4v
oWXaO+8pMYSQT35WCpVSWY/Xqq26rY1g++HHIZJ3XIJ8aAxSQ8nkTDUBznXxmCPfZgQ0eAHMxrvE
LzfaF+ueSIW3dTxJ7Z7CK17AZ8tghRjaJES6IiikJDLBPEoi8hVxg3fRPaImEOjFXDjlhEz1rWEH
D1QKFsNoLbfK4lEDSMLLQf8H47g7/ZTymZFAciX/t3NdS0BOBoLNQGy53zuTI4qOmlp102zKNsb1
FgGF7xFIQ1UDAtBRsPKmU6p4lsQubiND14dZLt9kbdbVokYzBxGSm7zmYckMZnQGrAxdqgeomoJd
DQiq7Qq/pnSJcWrFdlyY/aEIxEqjksJbFMSbO7gs9TqSl5RNOQV+KQ69hwmchdrhGZBcf84FJU7e
pnZHhTruE0QPZaoW3DF9aqGUeTd5jKi4/NK50nPBW9sS+zb+bycf3z2TlGHYHzLPSLRpf3A+MdMb
ttKZiRJUjIg6rXAl1XIef0ZAfLtNkmM7cqmWyQ5KJrBOoGT1L45NE9p1/G7OoimFZIu3nQI6se+j
K4fGHTad6ksKvZLIQlnKi3JvEWLQqByQORcUZHt9/A6un7mDvXDS8B7vAU6599MANmE5u03uXDD2
dV0wQo9jfjrG3ReHWpUAPghsmzneW4F8ekL6JHES/nDFcqIR1+WVeBvCgik64E3pKtBmfS4ZMMJp
PVfcXXe2XM3g2p1U1sgagOntRC/DFPZG//+oF57w5g72IdY6YT3h3riBN0Ifup9M7iiiE08RKlNW
SYwmTfsRJOdsw4pr5jLzfZKCsiz4OiEAMhB9Ym4irzh84vlt8RUfXnv8A9BrfUdeyhmP9N67xozs
H05UyCn8k5Iiqyq/9aLbQdF2Z8CGoSiuowCRCt/+kj5ecTVzphNfZGDpkTyRHpI0OYLHx7r6NGUj
UgtdwsYuN+1WVWtU3QpboAP1w1hXil2X5kG+bhS/IgGqu2esdrv8bbzxpatq0ROKntaGgQYxKz8+
zWjc8VtJ7aeu4VZgDKef/wSccP1xZ1VwDl/PVcIv7GenQC2Wed9k0ZGQjsE4JHe1BrsSZzGWjR1L
pWSNXJx+VGfz6XIigl6luarN5Mr5EK5ZKbRZrETZ7lT2XNaqTJ5AcVWMsMKn7Hr5yZv8QQtTZpra
UOCt70r/U/h2Eb4P7p7LxtjdJHNb5vFOwdTs+bM9doZFpICceVHKnyBPO2mPjUZt/q2uLiptc8fR
kCm7KHMIlZ+lnGaFTQSUo/be8AGXOYeirFG4xAnyNOOZyQ383pwgHFFH281YwaRRa03Nrg3bZnUf
QEbZp8WbadSML4gqLOTQ83zc4vzq6a5T9ystc5UTiiZJShr3dphtgzgCGh5B3WAMt7x4xOGGeFvb
vtszfSYpqMBqx2dEmf9bDGzlMy49qP6NST5be5lyHSVga1R9BkIltwzVt3e6AatsF4KlkiqH9zDy
hyjuZJQL+/2HTAYcHIHctZ4f7GNZAfgm5mIUjxJnw0B49bnqVUUwEWvQ1d0+SPzMAApr9ObV1Z0T
NlYqf/55BDyTMW76+krufG9aKwLr5bwa5dCRMeQoYFaoMIkUXEUm7B/dVp+umGJ6xAvoZmpprZpb
dPow55K8fhbfTCsMPKYIzX0lr14QiHEuoxXlSi7wEtG5xev6azG5d6suh2v35eLI90feDRUvkb/i
JAc9oodT/L+wNkLkMHzPmE9YNXrHY4yHenfUPryiI1hssSuDRJF5RhE2uAcIhDrQ35vkZ5lB3cx2
hLF8dMfIheW+Ib4v2njnCHSZIruwO60JBw9wfJ4XJRuyLmSbZ9DKz0b3cHQoEutNOfZRP1Q3HVvs
/vUV6yURuCV/XaqgGrOqFofhJfze7uUsQ0bWAnfSWThVGCcOIQptSMgj8BL9K4alZf/HS+tm4qPE
U3pggbWSrnevbHPiaMmZD1vcg/kn9xA+PtcY4tNY2C6xtdtKQSNd1nktJYLtVwza/oHWDHKC5W7n
VhdmeUcFA068HoIeLc4rZXRqYYS4DGOZC+IG3Wx5IVN+r1VgOmM15ZcrTJFBcaJxmwIhX/BdUP1F
uG4gxXY01AeAGjNd6uRWi9TzBQgB1GYqSv3aLORurbTK87n2NhNbECiXdc5IuY5DZvHqrouHLN0A
fphQZ9tv3GatUuvr5Txba5+yZw/eiXQYkMmmX+t2QGY6YOMSLbdWVp2a7s9C+2HK6eUneRzv2jCM
ESzBbmfM9puOS+Io+DoePVcTJyvtc040gFM8MrA/uyuaeIhib0DsrEvp8lBheV3S3yySbMp0yays
uk9skSp9vDB29K+8Lkef2UYHxyHUmKZSJpeCa7RrfY8xPtiwlK1KumqspFaHAwYUPBZKwqLbdXrz
efpSaG7UWD0uMWBpRwPShf3+/AUVSOuz4yecKCMHgmLBmEHzu4efxfrEV3dqp+Kq5pBMtCbRZmjQ
EPlJGcoAOAGOSVks512BVCg+ZJTCG34BPz/DYOt3LUQPH6uq59BQsoh/Rtm4XDBIbWrYGat1mSzH
QQew9mPIBGFlJ76z+DTeXwdMBXToDNnxIVAa4QFoUDFk4kttDHoq7Xm1cy0tvoE6h7uUthKmgULS
KNRYtukGHCDnj7kJYR/oZnGx5VVyrMRZtNdeN32X8bWIbZxYZDEyQENvgEjtI6AVePWURf8lHwfl
lhUWbP3N37eqTSaos9DcLeOdnXzbTD8QMdVlBxnPxpfx3wN6wDvKQCII9+CGQ0HKEBQ10COCSO8z
8EmmNOBR2y7CKCtGfja3SzjLww//v4IyaqU1A6c6yBpKCwvk7tLzHhWfIsQsMqEncticcmSqnMex
eJ8/SNCXd8d6qm2yt7cjQloMdHvw5pMoJZoXjsn10RuqrrN+b5g0IJPf52J4Tc0nLgy3KYaWsrJj
nTF0G5etpWbdw7fsFxg1aPgn2TRcU+pAT6Shyj6hUCPyrAWOZUH+V903whWQsI0tk/WoQiCuOHec
JUfFjW92XyLWrkbA23Yi539Eeph6e/jNCmE0ttBjHvhSi9vncWeSxqdT3dX29AZwD0wcnP9SrGrS
wE528ck4TRUJP+3kyLaAYmAFC/66M8h1lJy6MnzpUcrWLbOT3Tdsjh+fozNcLkahkcL3hsoKtHQ/
Vi/Eo87Xc/fb1shCMhufXLGxUShydcnBrtBRQl4IaGimJ0Vb1dBLUj7ITiOOhmJf/kERU09/B/RA
QhY2QU1iXVfKmvJeQ8liHfe/H/unAiZChLw5YdugzJiKYs/MiMwHBW9jA073EeaeNWVRdM0VKKIJ
HWvLU1pk8JK+PIwmVB7xw8Kb0il+8KTMKLG3R7CoCl0QkUaItATe7Yj7mBZUrKbfGfJXTvVKZ1t2
52dGnLq5HVKiM4UfBKaFWpOeuH1wDbxcBBBetCKrPqLlTM9mcRmziml2BQY7x9teQjHgMN+A1HmF
KFR2hS9yxe4C5tY5nG3uysarBcSNs+kbPj/XPbsk2QDUPAaXvH21wsRv4cE3W53dTXGjuYQ7sHvO
5Pngkvc7fJrZZyjK461CbBazzHTUeE3z2I2wuLLDnFr1TgqtQk298pj3wVWU25G6uO+dy3cwviXY
Xxvs1JkqooqnAuf6tnDxoZ+Kikzm4HKZd0CUym2YyTh0A83BXCH6Z/Gaon+9/S8XjqQziG4tDa2D
hcV7iYO2gtnQANGPNGMMCs2tc1xKwZDyPX0DeN3o/ElxN65P9n0AID23POuH0elmNKCpy6YYumZd
mBEV5qDbNj290AYKdgPnP9OTalbaqgEEU8Io813pK3mdyQyLpVvk/0SR5eq8T7HAb3PQjAuAcLj7
Cbqe79T3nFx07jB+IGcweQsxJi5JPc45ZnBQpkkGK1BXTzEOgXIWlyHcWJpei/sXFz8FKuQF7qkJ
PqB732YuCUxTZJ02W8yojAJM/C8qB4bY1SNxPZQZutwIlquru3+7VLYBOmoSL50dspEAoiGOnpR4
nBo/ytlg6zMMFzrfdVpCgBi4mo8vwIsKtd/3yor+G7tySs4yUK1fP3bCBJJa72ZINkvhtE8Bkuyz
URyAES9lAfHDIky3mV2DFiqt8t9mRHCim7X1fWwYPPLAUYTNwnMGAwC/KdCQNXxOnhpNFlRWIXHe
kwDNz5dZ5YzsAh+CJvi/lrVS0otTdCYu8FrjcigokX+GXN340hzrNE0xkDTqUZzt8X3pI6lL6Cug
w1L3b/6u5jO0vgm0/WHUd1ylxUke2bRUyYL5hxOn7lmPK789AjfOR3CxPZ7h9fYHDULWtWV/qBTH
z3gBStsWOhCmuyPMYHP4LdawtlgT1RPfLQWoH81+hgev+YCYbq0pzj/pg7n7BeqY/K1jeyefzcIo
po8mylIKxh8fJZm2x18gY63/aH3gBkMQh4aIIJNh5qhCALHdNXFsk3eLio6Xx6BqbCLc3uIszI+7
dcwVfbHn4a9/VF7YNTTxHbir1GZN0odb8J5Up811aC8ZKRvstTqAUV/mJS//ikVU/9sjZzqlkktb
evH9cUX1Yboy/xo7ue0P7fytGcyeDSdwpoz0YLIfDHEzel7gKnhsDn0L3eJzl7ZHOty7lQd9nEyW
fcOaM7AwGwG934PS2yjrhujizAEM28JbXYvswuGh73w4zkyOkW7q6OPqIs34kmpkfVpyh291sreB
4iXd767cR0R5L2M6IeVV2lDNHAVQ4JZ8cf64f2HF2WQskPmrYWxxAkwZemftnnIQV6dQB+s9gAfj
I1/W/I6He4dvjFTVDrLk0MYh/USfHRB6GpzubqUpcHY1eZKsyPIli/eqm5H5WOAz55Nwwxvgat4j
IPmf+sEvIg9EXxcxH7dp9cPMbpQgyojxnHr9OA2p8gFoOZ5CHDUfxIiOZq1/5PYeYXmtbTf2jJNb
TnLn04tZFN8b8Py9rnfJCtdHt3HrDLmyYt53kQ/HfsbtlJxkdDsw35OM942Revfz/RIhdbNGO/k6
naW9hXIcXt6sViNOD2BeymssjLuJPnMVPUbPgVo5BVD6cTLVsVAowSnGtuksj0wjdbTo9MufcJUD
o8HpbV95+aMRVlUmCnTB21WzE4B2MUXnMIy0iF3KvU7pJX6kd5ZXwI5nD7dADAhA45wjZsNINsvH
WsUutdIXUQHpUOlIqzDm8is3VwPIqjAYPgky9JW2l095WB/SjxW9QBj7tL2ZGD8ZUfTnosnZJJ4C
MalcIyk+dmyInzVOeopHc3guFDEV16cV5YXm6nKkvsSlWSVOMtTng3rWREUXZxkhnQ6WyB9psXbN
eTZn/Rm+4UQI2hDoXjrbVqvE4xp2pMC0qpCxopm+sbd7DyeBKXOLbZ8j6eBZU6lWLmjz6PpxnAgc
gRf6+m8gzc0FGzdQy0++p1gtu2Oyg77Hk8oyUNRGII0CA3/1KDjvNdTfkEuEwYIf+G84uNQurMH9
/gPyDJ9AiZz3UicQKejeyekxOlENYoJYppzRJXo6wusvRHocXLmGVNRqDWbiISYmEfxhQWiXoNVY
KjIYwL9vd7hS7LM49UPCmXBRPGoGB4Sbi1UmllmpNSCbJWmkn9nA7Gyfyjt4qI+29WoFjbDJfn8B
bSShQkm0zsNDPPcb0cRpgvq9IY8TIZ7la73hrmXasq1yA7/SXlhRUCXeh1PiXT6gNzNJGs9h6zcw
3gEaxehPV56Wh76nbsw9mA7c6d14CUPZh9gjfwsf/wY3XqhodoMQsaKfuynizSuSHK32tmKnds8r
eCdtDbAe+Lg5kK4q0hY3lJyJx9C3sWrwX+a2U+krtwK9tA1YusVagq9+9z3hdHznDsjwMa9ULIM4
5+byllCq3VnT9yAAgbIiORFzib1ZBWtpmh5Z0VNOg++u5LKc9UNYTIuZW+1b2K1S7Xoiakp7miZz
olgqkDxsv1VoJvao68q+/hY6ers/jpGx3i/qA6JygRgRIJS6CBpcWszUXcvJC8pIxkQmVOP/zuES
76DsHb3j4X6syknTD68jcvRW+paYddVyl4QgygW8bCTa+z6zcfCKdYp0MgI2i/fVh7oSRn0gEUCk
rFWWa5c6qID7ZF+7C5nj7fum7nUS/6lQzXGlwod5kuK9S/z5EhNXSycVW4zSQ55rUAXlEONmubW+
vnVVu32/o+N8CiTTvHZ9fJRVxvrQx2zvFrJBkN+1mhFAch91CdAWChimTssTCt1P5QnrbuNvKu4u
hPs9fi4O1UPtPAdJlAzZyY9SUhAJ2Y+OOQRojNu7ORqpf2yc8/iT5oshPjL4kdryMcHmFVaxi6lS
CLcAItkOYgCWHVqh7MJ2mrfyCXysWnwCTZPFYgZjZ3ysVIgLB4ufHX7XwUCyKPbR/vLyRSQKMIBP
gxlDJ4SHIEBSSiAXnNZdWvi6SDvX+icZhUl/VmUyncVakrTGpJpbmZBnKdy/YkgZFWhJQNOkeLSL
3ACQw9X2nk6yjlFlBGAd1gEAWPBhtwFuom+g6KW6G0fbNSN8hHtCfP/9mhO+XMqRj5R+KYleth/j
CGJdlmkEUhikHi5y2K6kGhk9cj3+4bP0JQqY9oqIrUu+SPNCSpIHuHfzU3M6H8UidBDgJloebAYP
HTyr/XZ89o9aVHSIQTpJQwqST06te7eMlWNDL+n0e2XwaHpo1HLjl2ZH/4HqOl94gAc07tmsxfxt
JXRq/vzR1kJxs/tnIdYsSZUMRYkf4U4CtkffDnH5geg9GLGP6iow/g/lwBk8b5HlF+rMWDCW03kR
CZYKU79E0Zvmym368S7fobbrPQioNhEn0sP9vaQCf1nyovSk+kXaFYbPprCRhjlt3EkYxuVeMpG1
Fj3JaA0pP18WXNP2DgdsjkJyYqCm5rXWigJo6rzhA8jzdmnXbIQcC9n/arL3mSdv5u4c0UtkrPZe
zXuH5P6mvxb0i80Spb5aQj7fcxrezUBZZ4Fz/lj2CBuxFv7MYOTfR5zoOjyiUcW9tvwMFn9Ljtaw
38rxLwYjKER4erade2ULuFoxhrnbNAXJUr0BcL2pkip2/W8WqUyLUO+zAq7e6YGysoBJuk0d+H2R
TCYE0wObCSvRHUiSaQQfTev74SGymjIQrcIlNNVCu4jUle1MJnPguyEL47aWhp01hMUeLd9LGNha
jebX2K0Lmvnswu2ugL2ke/e5iCIjzmZZlvCpPHWUD0Cc9vIHSlboqWh6ufabt60oKYJg/daBJThL
oWPvz15/1HkpEJ0b9+SSTpoDMAjclrsJakyYB+sTtfmRtLUQA7f46h4OvkCeXWkNd3pKzRhOs5Rl
5DWyGHXzvCmmbODAVtioS440VnuEUF10qs0de3Dy2vj257PlLDcd8uQzWlIoa96M4X4gkAMr/0mY
wB4dMa02d9UM+ygb1qtmRS7JQgEjM+9cFkxAJIYJO/R5d6kBuLj/wzun/REavyZRp8HxO2qdimrb
2Si1xfrRK8h9aPDJb5Z8By7lK8nmgvJLCMNPWIvfIC6x2WYGtSyIlWrBQaB5YwipzDot5DI5oWkc
3wU0TzEzRt9+AsGANL44b0dKeNInxWPwbuaJeWp3SwKJVP0aPYkJCf3esvc2cBPHxwEQc+Jzjpm1
vIzo00jBy1ogcDnO3Un7+J7ceKVPjUgvfexb6teuLC48e1zDpjD0PMb2F8KLFVakmbg63U7682Kz
GU8qoGcX8eGE+DKYN6XrCF7epS2q12KhgZk3cQ6C/psZ2r6QNTMNhEm/467llcxHmvAF3NRFnVZM
ov1UBlhl4Kf77qmYRQBvQTRnBgeNtkHj/pNpQ4+aRwj7dWiIjaG9h4+z+6Oh+zY/uSNoRIclqlGI
fD1cd5v/x/bEGER4wcn7XBiYUrSJywp2nxouaEEoe3URBIwxyLnJ8y1O4kfNNiCg+rR3KU4u295H
6PKeOtIOeQ0OwrFkSlFSetfZ+s4d4A9nSeX40g6zdGMFD4hurfi8WcMtZV9hc5cUyirj51LaRSqA
iC8lHegt2Q7SMira7OKskg9wRasRkSlgImzi3gRqQkyygPXpeevHbFcyHKhnHmN4asMCp9UzD49J
ifZh2bZmyuotb2ANqgL0DGdkEdbiDwbf2Ph2b6KgnUdWxiC9C3Ocxmbr+56bkmemCRX5fr3OGj1p
fdap+UaiDxYh0NlTh82ShUOEr23aKwBw8PcZhrEhOtu4R70/PuIqonuKsOIJkDNyjrBZFrqiKdNJ
u2YZHJ2mOmMLOzcTe9QvZ9z3bOE3DC/QS0Zk495hmTQdTKAMDNIYct1zw+rLAZnlR8nlYCmK9A0b
cmqIhMCPpczD11/mDp4DRZ0z2hcAV6ZOyz4F+w5n57+GSRDciZAk2lP0W/oP2s5BsjOKZk4zf6Y9
QoNtR7+/377BRhmac4OpnOWblWRWjZRoLzyXXWzs3vtbgMW77EsUdtatv+xCMSe0DAsoMythL5wT
4WFhGmG8BgZgFW57vOP2xdK29Gdh9oCWlnp01mwNY7hWiOgYooTwIsHa1kLIHuNCLQFlwlDYKLF8
3hiiK8SDIubPRujCFvd2OyFgqCvhqUSadTCfVNuPb9Wg1l55kEVsQzoNSRzbxo26I9uztckj4hj+
JGwKL237WJDboIEo4/csRvWqBn5hQhuHkWHXY319TDmvusBFV/l4Kn9J8cAjaes8MRbiJWstc8Bp
kCf2cFbfUYonQqwFLk6GzGNwiTs5wsUE0cnmsGzeAjqUuNR8WGMYuSTodqaAFT4Jfr5OSM1XcVPF
w9oks8b8v6+c6ZUNcQjPh6Muw0qhPp58qiC4hlYmPh6LW9n8lyZCFa3p2qiNfp9doCJf9vVSwKM/
p5UziNs0AqCXyGxoyfyI7AfhAxoj/ZdrjcYthMwmpQkeF+bOEriJHJJdd1miqUNtHR+I9ht6eiDU
9VliyuB2fdTYkreC86SsNixIIrsVEKgbEVcP1oyPIsAlOqVYQIorAjyM0bcuUd6f7N+kbvWcIcM6
hy1R3PW6Khezws0PA3Q1z0Le/RdS4Sor/NE8MdyW+ov9eV8CR1ZtcanFKY8lQpn2Mj1QV28ZidIl
pCcu/MwvbUWaiboOdZOo4GRZP1iKshXUrgbflgWMCs5DEIT1XcS7UMhJIN3++otRnu3c7rfeS/L2
p27neiJ8dEwrpDwZardKynJmjdc/iRYi08I3jl7hkMTdJHlsv1YKLeLFrzBS3NYsQdCmRQL0qVLj
izmZQiOw5+nMRAhzJWI4f4soDUG2mSMRotPVaDOxaiWjh0bOQTdccg38gK5bzxcPRt9qeh8VQrW+
nLZiI9HOBal10CqDLvwLgq/e4GLmUT+lgdahzHncNi3f2gJa3EtmHrLZBe+pgF/oSd3QLbgmCz2Y
J43oKanHobbIJ1uObeprWZGfgVBvmgedxE5HkXFat9q3Sag/HXR0ZF9ZxPy/wm/ojR3nhG2HFxQj
bmU3aaimfjX3v7ewZx2T89jg5+tD9NPzDCyf3B0bKtW6D3oF62gv8TTzr8dV5Lq0QLzvDwbZOMLi
cMNnAGcHJrLMvX6QOCSoZ0BqS3GfBW13vJC1aiy3y671eeAjFIPls+DQqdhbqU3xr/xwyHaP7eB+
++WTNCkTUOJ2jyUjajmbe4g7xZmKPRC4ebhMKUNvXAVd2DMr6iDDgLJhy3ZFFnvF40L93Bj9jtDg
SXI7GVnJ7E4mYLjSJlGIy1DxLQFsqPX3PQOd9E/7ZXrynVSsIe+HMEG/HOPsozcYtLFcNMrAEpTd
aRFNYKY2GQuQFR8HpPpQC9LapMzwEmTkfVJd/9TgIVT4zg+g9uG1OCxtjN0xrxE/qffnvckhMzgX
G9ivJD1bBgFHLRvSOPHWixkQ4dA4UdJrPwbgrql2/iHr2xGxpSFrwJy2td/q8ZCfro5dDQoTCsoX
XO0PpC0ky78Ic1DsiNWJ/zsykwnWVq9to4RocHC3I9DusUA3KWKya/aJgBLC8s2LsOgDojrG5PYw
zfF21umVKzm4UFkLl0LtDFL7hjmB5Xbv5EicLxzwo2QRnzuRF24F5TP9PWOjGG7gto4csPZVbb6s
Zgg9by7Cz6dbllb8V5hrJ6zFD1j7SocuRaSh9fGaNTd5EegvazILDedC1vWXYZSDRTxCUwSM0RR0
OjgJ8QYLH0sJUPu7ObMXJrG67qwvhV907wFHnTxCI8zi7UzHLrPoXZBXASKGgRKsnsoH/IweXxql
YeCLPM4KYMTeaj9m0eJXpfAz4OrJQDcS/4IVYsdnU4pzAJjtZmcWP9q9KFQOb1hEov+7/uHv4u/B
ZY5VRmLb0yKmu5LqjNuq2gF/fmy54UF07KlT7TW22yo7yaaMNwdpu4uI+GmVxuUkiwmBAQh38QxR
YyFIM6KT30L6PU1MhChrOonlPXsqkfUqKurwSEIsDe80cM24ahA+u9SpvuOovo/rq/b9AtkmV5wI
28IqG6ZOQ34B5ira6+ibQwoqYsCTGINGdO24Q+v/WnxP594pLk+QpRn9QifOQJ2Tl0tTvRP0NPay
DOgqyGcRlydQ517bGigvGev+X7pdRIVcwSTiUMPIvySenUno8JaVJbWju1gLisaiXPVjhOLawyqC
e7YI5p3v8tcq7dR+dJ6sKUNlXQaBj8rYfEoHKWHi4iAgVYwuBf8kRyzuFFka6MJYZK3p22ZO4/Js
tX6xO3sPzwqZ+A4UN9b9D3BEe8W74lLYp7/pjx864UfDA9+bKYUOcna4FDrTX6UrykJuCA2U19ab
B58EYYfSRkAqJWCDFYedQMjPBat7nkTXH/dEKrEtAz/eNnia3TX/pU9lTuSXnEPx8fT1rurMqCOS
kqlJTZ8pIOVBOzKE0olycvYGvJvW7TfUkUIMbotryCg9W4f7VmwbEjAl5X3B5Bytv2mjRrTwjQXB
EiSodxlVXkZHrGHzzAGpCtg5z2k4b34/sx5j92pqt9R3aa9f98l6aDaIYR+y317dy9TnsO1elxIS
siBoQD90x1Q+JWvf6O8GzZJFCRz1jpkDwZ++p0F97Ouvwdl2zp6TOhSRyrSHGM411IhntAzEef+4
AH/tJF8h1CnPUI24EagFw+FPeoHZ+NBIWNs+RcMDEQKWREqcC7CP6Cbf/SQGzs0c1Ou+cRJAv4bX
Jtc1j0slsLYesiHqRVFyw6r1nep+pYHHfzbp9w5Gb5Vn7s3wLtcACig/rUI34wwNFDS3rqRv63eE
1u02Fjdpmuy9I5d2+JoqFDGrvv5kFesfjCo+ZPuD3EP5AFQ/1VVxTgE4yoyOtiIzgAl4ztp+OYdc
Iq5N+/AUqjZAqoxQLmNUgLVGgxjf9MHaFjx7oUaXvErlPi/YvlI7qNhlgSmNHXDHaULLKs8Blahm
jAQvEwYfPA9UJBIRpEsbgimTcaZIc+ir6b50x2YoraZPzHGdwH+0KOW03YrhaC9XbuWjBBV0BX7e
wG7qdqFm7O8QHFRAu6vQc3447KLkVvN71zNhKbF3NWfOZ7RM6zhvx1lcauCtOjTajIYGdGX/qFRe
Rw4BXunbuNNia6FpZvlqMurIK/wu+bzH2UBL1cPPR9MNtHLdUnW4J+xWSl0jJosilTk5hbb2ev+p
0Mqcl7kt0kAfFhLKbMcbB5bpTgypg2bwJKwtIg6KREmWhKtkxUQdcntQ9yNe4NeO/wMbR+x3/xaB
VSME77jW9bbivhzfsYbbiI4aRRhieu1YKPSBNnf37X7sJCu5p5Q6S9HGgIM1VrUPw1kud4ztNewz
zEMZx0A+Gb4crNl9Kkd9yAkYHedLw7YCAgLbe6Z9LcXOtxiQit6UV1INJYE1Hxune1ntv4y6VuXT
Rrgs0dozmViO32iUw1QZwo/hh2fC81t1pY6QMeBPs4S0OoFQRBvZoiaiSAUqJEFaEPaqs21YIQqi
67MAl6oWdcZ5skvxjrIal2snl9Km50mcn1T3Ll3Yja0afAN5A4ilbnCPv06x87cGeg8DGCra+8HJ
qX6Z7eLaXL0PRTqh3m4xXjaTT7z91HOib7JIqzowwhaR5WwZJg8YZlV2sCMdefhv4H4PCllTikoW
boyF0x1AchsdXgZRnma9LMhYx5xV3pRf8DCkSafyBSgtWIlPal9EVsR2S2OgGs2z7D54pX9cKVJD
ZTsKV2A3/O+fXcYd3BbcwB9uast7PJAsRqw+y4BWBO48gqpBwOVpP7XBwhONvSLzH/6VzXPQBWGh
nIqGSb9ZFFJy5UJapLCv8YGNOh6dzNjXVhAjxg37Pexr7/gArZKGsT+1Qts4DMBTgYMWUWRUQNhy
XJuMBm8MZDdzpkCtTw/TTG6MTRLVxKxw4SrdADllh7BijU53aiDu/Mfbl4g2ngUivJwoXtppxCXZ
DfTK3m0DWnfUmcNuHaBM5KcexECP0NhHEWv0mnVaZRLsxCyJovPisbV1OkBSZDdL6fZ8U2TZ+Sof
CLm0rMMjXrN+pqtLMtn/dt7AC9oHEfrs0hsoptpDuhEk/qk+Cbuz6HvCoZCz7+W4tFMTF1YDauT7
xTnu/4eWJWnTVGhDWMrXniPUjHNKwIiQ5IhlY2s5rhinkioiMas8UBBazeiXrjhhzjQcDea1z4z6
eQUNIiFC69J7moT3D7PehIokuy39kNcPbzIkpJKkw9ccsh3CXctlsSisSog1fCVO/VfiGu905OtU
LeVBsrE/zYYrgsKjK+gcZC0lTv+Q0ZDmMay0tYtxxyVAKr2wd1snVejk/sElugpzxC6kfYbDL53m
LNMpH2FnBvXdGM5q6LDBPSyn8s/vUYic54z+jgILjYsKGu4ujecar+LYmhIGjGU9IOfy9czhjMUU
hy2WS/MrXapCdcfXYzXzdNikrTT7s9t0SjVuBmDY6cDwF3rSa30U887ElGWUGZABU6wVhXDLVPwu
pkTl/IxEYAz50b3H+SD039dSUu5rNh5/H22mGFDD/5Ja0PmCYvMrnrlOLRsy+GP+mwsEZ76yZ51k
gCtPptciW4cl4hjjfm3c+FtIzFiCVP19Y/mOl4LltGwm9YWe96/6gzACQ9eOnX5DOIc0+9MwDobT
wpwDqQispUfOvcAWrQAnYFymajjmsoJ0ocBxmSm97na5jYpDn//FW5HP5ffxouuNzAJgbPUfxAPq
76b8rX8vvkUzgbt66SfMsOVQfUdoE1eGpWSDpPxgqM+7zzz1JBmorN23LECdORWnIvfe0+Z6DaXI
dfup8/T5S6Z96F16Hd+8g4SzUwftiVN0Af4HxyJWYy7ceLhbrwrEYtJVMKW+zeDdSRZ8hId8Prgu
cOnzVpUx21RFywBxlYFlOlwCp1zOGdveaprppF8gpZmgqCDqmHKDyNbTfZIORcbffDldGCgJiEg8
KCdllThz78sPYtto6udT6ao5O5ci8RJn/0VkcvPgGCuW0spov6SUwGq0cfypSIURp6fSTagm9ggo
2CEiCfsKZwB4UEO8Pr+LTpnORXUGpJzBbnsNp6tguxtiIQ5lvOmqZisodyRvQsJTif+wsp7g4PQN
GB3nRhvS+RTSdmX/oPjG81XloXfVynDG1qiQXx6ArCSqOjtrrb+vOPALxJ5KLo69nKbVMGec7jbE
1ZE0pkvrBsuzlT2tcGx/N55jTfFO5PGIJ3h51bYX1Av59pdeYlFzxpwCDjEOXSulgFRQHfAvs0sP
LyhpmnQRNWqbGy3THwyNR7kbxXx+JY2NjNGc29vUDptBcLnj+5szSfNu/1jfQA9AAB9DfX43i9tE
mghlTR1xGIacSySmYBVdxOp6Xw0DRAwO3WKREwSe4XjclyNapG2Np+fOklRnIdIuswfXSaaUfPFa
egSzW/XDKiM/mH29ffvvLBsJbpFikrkH/MARuP/tViP/K/xPyCwLHD+/Gqw+H0h2tQ1G7unl56Ln
FBWOP9q7I952Qa9yFLZsA0osxJUhl1rl0kdC+eIu7YPL5eSdUYBLys8kxNbsv+ybWZlTaTNcxNUz
4DMxVTVuQI06Ny1FgZxvH/12spHyyy51A4W9x5rHVcxPOPy9XGO4R8ni2GxGF1GiaOF6o0/RSbXz
tAOpRtjOn0AbVRy64TxuA9D2LyqjsD5N25z4DvFcx9EJIj7/iDJKo6pGgH9hmil437sgtfsD1qAU
klbJLXcHdb5Tl7e6LqvqLSjQqOAvUdn+NFBByxQjXcQ2+0/5jIqUurin9lL22JiiY1UQlOHEdjhW
VmHdRrE4Cdnv1HmpKi2VnMACGB/k3Mi1LBDN4sqg+vEoumxx0RdT0GyjAWm8eFTY49K9vTeLBZcI
b8ZfwTQ5N2heCuE4NUPHeIG5z+Ath3alrjCkBWePzddIWf1kajqzY6n5Z9Wx3ET/xJxtdC+iPWXb
Q1kVqJIp0WlGFivG2s+4igd4aJl/f78jhy5d03NAK8+Awf3TL5nYzPcxZYKQLWO3Hstn4U+9+VM9
rXWcoZt8O6u5Zw3TKoyHBr5L0i6b+O7exIQj07MGynAYjcB4EktySSRmA1yc4Z5K+oaQaU2HwHlF
ICh9BeZ6WhKQhmT9Wxi26jx1Qp1Aub6IMu7SX+6AuzOxP1zzIta5zmCc980a58hCsXA+PnbZjDq4
R51aJJWvDmAhmsT7yta/K6ptZADWVtJrS6rIw8H5qQv2LuCefnP0vxUkx8NAPjPOcYH1Fecw7lHM
dGdtIqLFtHesf6tkqK/jxP5CeFHKu9cog2/3s+bmLbIwAjtXk9nggK3EXmRXItEaQjulssOg3TFT
AhA+rUftDQckGaE1Cz9sRuAmvVB3MtR7PvW8hbO7yaupyRpqy0qCeKNPQ0eOT8qmQv7M6+xbP7e1
CfJ6CyIdrPEejOCN+Rsh9VjZ6ZTQpIH4TNLUk4EedAWzYFqHRRIpZDAzjdLuKIGIXhdT8+TCPl3k
65j7yhnDMWn/DpgeTWIat/RTDT2fzlbIWi+wQkc0qaRG8Br7ZmGYdRFGYWijNdsEIl4ZLPVmZPd0
QyEXsnrkgLMcgNJQsEe8jpjg2ZXqsExHWV2sWXeKdf2ieZLSIqoiiUbFZgxinLMdzc5f7DYcyaBN
Y4S+JEEnthl1lf4SB5j1qcNl81T5Cblb92oK5bG70Pt2TpEVucaW294tU+yS6F3iOq1e0bWdNixg
QlJHlD6SRPw+5hBQcHrzdbXg7hXM2eHhKRVJhRLfTXn2aclI7GHtzF7nj+O+9ErK1XS0y8PijAQ3
J9Y4JJzi/0lflhcYaRnlcu+H/f20L5zPwC3l2bqwPOA4eobhRluTlkyZrZpE8X96+PmNqJe18PJu
pEFSFBiZca5hs8OA47SWotJTbzUf4AN/KdK19YN2KeG2ZEpnTsQwFFjQE6iaswz1gxicyQk+XqhQ
u7qCC+PBhQGMyEPfcWBPWChL2KAhFHrtXyV5RalTMdaF9c+v0YIO16/pnyuSUB1dwJSrm9LFMfA0
x+fhXD+jteSn3B1QV8+q0Un7j2h7AsI52zZRvqpFS2IGEx8rQcTmP3ikkW2O/UIi9oLegd9ZM4FO
J9nzJt1wdtTle/4KTzywMcfUf2aV71pWj6L80KYHkFo00b/XS3TPNqWerG//3XzJ6PKa7RqgXtgr
DqbjhAr2UYwNzcgbV40Q4neBUMwzScWODMxecznnl5KMloPya/lErUfyTiv5rUELsuz7FJgkx8G9
8XqA63crije+uw3JstYgUpmQ6WvZYWAefl+joD8f36bSgmfFAAyHQAZMCXuX53hn2oC9vuh3PcWu
DqVJE5uFh5QKONzd+YcK6lrZhAgE2l+TpdnFTZzdYA8X112WvRNWjJfDL11h4clZVOaMTUTcATWI
kq3txBm4H0sgF/c1g+CJJcIG8FqZZqFgNWz1EV0gc9uZbogM0vxcPL3rYg9t43ggNRwghHCRVrsE
OotafJ/+rvyLiz2Wb1p7SctcuCFWivQJuz0fIgZt83O5mOuDgSA7kcLn5keciBe/71bRZNBtkPLB
SFmRgmnz3Unf/yWI19c4LaAmwG1zWqhbaPFaeNFxFoDYhdSQXqNcJkjBlPGs3y6P4kSKNr2DYbqB
8rmtKO4iU7I5AOvwV8PEr03cji70ed+ltwXYOJkVWkfWowIW7ISjAmRhRmyIrZ+fp9UH4vAs4MCk
ZHrwjXIDAcHdPQAnrdNjPRmZym9IAc63QdwnWUcCSt1cEPqx2vEvtlMt3HjovhRZlfsvXngNzMg7
wvnfHRYEegFDAzIVA1w/aRLZ1NR6233noT4PX/QdWplPCgl6hDAGarjLCXdO5n9g+Yj8iJX72VYp
PxJ5tVzuPOcu5bGCwjIAEERgpmYfEv6/I081WMTiHzSvdACXE7ohCBOzRySaT8nXDaeJf1hP47BF
W6i2D7oFSYzBoSd1SDM4C4oxD13Mpn4PPcoIbXdljHkG64jcRF+6QZI2I+kOrflxTL8gR7i5aEq5
Te8CQnQ1CnXiUG35PGcPc08jsW7eyUZh7I5wfILC1j9puWLGBD7Sw5YuvEX7GgoBi5E0CTzVQ2JD
D3MRTgqDrAlBfjnCEmoNwPTbI6de5LZDmiwjE/mJ/jvzeIJJyxXwtiTIPa1Mqh1/0a7jiV2BqqO0
2mxMf/fZ0TEhVlmtUEJCVnU3vY/EpfWZ+RPhsaFkhSM2MqrYJcaBJ+/u51ozdYVNZGtxG3kD++I+
UCSJEV3IH9yXvkLn521VzqL/7MbV5jRjpOeSjN3R52/masVJ8mWjfkTiiJicASZWNpAhfwivLNrJ
iZiaN2LkoC6AUKphAbIL178yYWdRyNLGDbJgZ4/DpCQW2sfTYXzzxd4ReRz+b14KFekRAb5YSKfk
DxeBFdcolcIwfCK0A2O090j9bE0Qf9JJHGgHLfWXf/tkwDROw8a3DjA0WpJ9uVdHPWocd3TnUxZx
QF/1b2yJhsyVEUiFh3CN8kW/d0IhsLquiDeRV2Z6F92h23elz7A29RsbtD3A638n7QcqJwSMnuFk
Wcp0MwrNf0bpJWG5cRcZWZWKXhLibU/bd2pHEMCxzRN4izeU1KfiY/Th3hvXSV0kUy4lxrZZH8rI
gcvfe4YI40mBaUFqaQMWEmiK6JSpIwmQvIvgMec9TPAzA+XInV8NECiUoifZRVVJixqa37oxiSwq
kt1seyXT4ghOpD+TmSTHdS8pdNDorfanzntQS2hkqy2FLlHcsaLNMZ5sZM1brjyMPJNUI7N1K1Xq
vfTBdXcS7BcMCTWHtWBfuBgLBBbIHr5Q1o4uAiZ/2si/RrOKzljTOvKj6e4EX/Rp3uHdCY0kYrBN
eo+dK1kNM1DiaU7DyuuF79K5LNP6A7SBy0GRBvR6DEEsFhTUj1th49/eSX47b7emKRaVIuQdyXG/
VY1JHFEMrTow1jAE9iDMqpBCem2T6qk4H8fvIU/wARlRBU60rT5KBhCo7Ov6uY2NdHnPz7qdpaqx
Cqe+XsJfAESDo+8JffALcBH0mR/Ub/uBADh/MIBD8MS4HgHybai19z2TQi+0dLVWUMuh8X0vhO3Y
xwFhEwiw75w6xcHVVmIBw9W1wE+oJhZ670yGRiJGx/KpfgI0zyHSI5YbdSu/4OXCz9eXUy0yoBTE
xDzLT4o3IvDQLQOMUql9guDlT83i6FDlbmtm0COKRfjB1nsvTso3KulStZBCkqQZWLlbRyUe9xfE
DuK271j+0Kb9Lhppiw0gPweWfouLL0D1ZhjazqHzjlTWVDzAQIrimZ567tDLjW2UiGLcWJ5zkC+j
9kFYUnaC5VH18I2TAMi7cLd3mWD3e4xBsoDii2og8YXPe66TW7OYhyyhhsmwJRdXzHaTmlVnOzDH
SjyGKnI6qc4kWbtdpSshTQbKbzDFTx9l//cWrjOjGzG60aMSJAEc0f9PDjNP/ZCwrcS4D8SvWbEa
YUOBDuQSU3WfbJ8hKk820EaFQ0p4OuXYazaLvRJ8HqaxMLygQjnoou19xFlPnb5Hxu6Qz4Ohx19B
ed6RWHvyXTH8ZIg8giaWL1+mhY4uLemTGl91XnAT55TuUH2G0kYCrE6jU6VrcCXk4+PWbihEXkgC
adEk2mU2PjiceCVdXdv0+WNy4xdbf7pWiVPxsNE/QY1C20sjPHeBfiX6ZAQKR+bjsH4MnIq0wKHZ
yTF9110RvLmX8791RWkOC6ux+XKx01jFwv8cZbXJFFilIX00r88s7C4CMsj2n6iVVtnQR4wGLjze
yheh577SNCftY5hWIlNIrrzr/+ss2poEu/fPTDVGcIyK64fQ5XJ4IX3EDdk8Nd6T1sc324uTqylm
RHOKrAr2rVdlAeiDfngQilOoY3VXeMIZ5V/1cUK7jzGCQbvcFUd/wVdUN7gO8NEd2aYqjn7Cq2wP
qPyDPa/RrIfbeSnqiNTMqe1pGBvsrAR4i1dANJ3cSuZP3aizfSnQzMY+vQo1c1KIzRZsEZBTBKPq
MtyRUe1zBOzoqYcjZwqkN90Jr7Hv9VQF45ACKPwkZNAJokaRNgLqSOLivZE721NkhciL92Vi3951
muhXyN5kmdqEnL13w5hBuI6n9/F1iu4GWsdEL03xJI0sCMHOULCZdd+XxIA4pPZNc01FER9I+aCw
DdkT6NStImcZuNEgDgiK7tNXe+UylMFhI7fFRSTLghT9ha4lUEYWo80KK+9riCUu8fvIkfyKakE8
8nRdKcHFLHm54CBcLd9b2u9VGzpDlB8L8BJB6xvUsOXXVRKKSbWUYNGdU93ZtRjiSQWHOUiz9foQ
B7fJVJ73SwLqHum8CzE2s9w9AtSsUeKkHhPVV0U/C0dkAr4kccTTiR1A28o7b8S4jWd5Vs2T0l0u
hkt/FHInFJpZ3BP5WTMwudLRpcqFLzqYG0+pGxF8Iu1kCrlK7hkC2NA7v7813CUyYv13CDtYIZIT
PiD2Ny8osmh2IyAH8PEecJ/fJuTHuDLZK8AZbXoiOqDWgVV/2PWNVsHbgxC6ZQcdx+BhZirMSjIA
doEGsxzlRusWYPoH3rKh9jJt8quesL3Btm2I/7zAPZmh0i/h/f1zlfKsr17AawnAO+MKZC6+gF3T
DZLgPXWxhAfkSNWDxPv8J3o9caHtVXxigjle4g0RkmMKLM3qjN70XWn87GPMy4q8x0N8GZh1Znfm
1lXtJgBDOJxat8aCnI8u7D6wBHJbkPYMk737JlqhcqS2VFmLpecrmIEihNPiwgX1Y2M0R1xZ9fc7
0uKcw4bFpL6BbdI50tUZSMf+51PeEd5ngy9wI81GkayMbRqu/UgHHQCq339iDAmPnyPMZUkjiYkD
72X7h1Q9crI7eAwCuummcQ5K/Q9TdJIpLSn9rqSjefQdroacZjlUu5yMnpL1ehjHG5oLTVNqe0oP
kWWcR+HoXE/iBsjhVzZd6vtJyk6eHegVY/XtHU8H9PkBjSR0Pg1uk/5nEt8by8ntzW4AxRKLpG6P
+/ZNpV1vgA9QmV+RfnaoF0WcZfQVRICbPuAi7RNu2MMcbsta80zhRZAUPY+kwG3MctAVDdkoDnCk
Pne14ntwqUegSlc9banR0lK6vlhsvKsLttIHjuPofVjs9jiLmcqeDegRSIoivrqKwL59hAsvKcDl
b+IwpL8LUbetZEs9CPnJ9FOvA8z2aObnt2lNIBWvCf63EnqwS1OPQPvWd4duR9Ca3NxdgFcuXrMT
Jt6oAVzu9LVVh2eIVx/9eXQF7AbwEblUkuhgyg5mNWkbl3Fm+91AJNijwCQIn5U6lPmP9mzgZ0o8
YbMqfR5YY9tlWMYILPVpQzEh8QE+JDBtkWPDboAM7u2+ssrmDRlMjlphxTlGma2hfpuhPbE5d4/b
uu+UmFn8vP61dksQFVcQEfZLuuCPS364WU3SLq6q9B7CQp4GIBiLL8pHeIqvoIzkgp5AlxjM7OQT
ug7YOw0mbLqU53OvAeoP9UE7Xr7s+Du3MJGxuJP3HKLwBWbJTxn4TUaG3yBwoAZJKYayIBHWKij1
mGyTzvMeDUB1D769BmBa+zWr0SxAM+OKD1RDC2n2lfpVnKDUDLEqnIBd/j1KT/1LkWO8tBBnPcpc
H+iuV3NVl4I2EdIGWKQrK+w1Blv1jqGNrMHNEosPCYvPVLrKFLaGAsSf3RS6ytBkd3RgNy+8sGzZ
ZyhNzTZEJ2r6GHtXtyOT27PoyXjbPS5yVrGQXZ40EslnJIXrfFgNkATKvhlTd7zBRgUnYorPYk+V
Qv3dtJXwdAdAVcrHDNGrmbCvNh5KHVCGlMxeHjiPz0tnhezyCzPQ93HY3i/3M/GVdI9Kypkqm4mj
uJsfToVBWsqiesSTkwLreKBc+iIArtCGzGgQjRNb1L8N2E+9ebohP/5E6m3k/rKkVqvNzz/5t+sJ
LD+rz8Otkxo4LAZGSZoAWTa+DMyf6xTG2SQiwABhY2rOo1MQAk7nneanw8w4uwb43+tUowbvwXbu
4RnFLElZbMk+Gw8RZqVTNQfrDO92WkBKAWa9r4fuvEZJlWNXlpL7GnZmKMXG2tMLolBXLdxGshD5
OkMq11CVGr4gLkCPlvPDapw2cFlO4GXwFIW/r1VFUuqOZOeeJoKRnCa3bguIphi0aiorfgFPRlUb
/cnDn8Fekola1/WRxA8SIP8ULaV9wvca5ckYdAZBGX+glZEvpx6I8B4DgZeQ61X6jVm/IfdzdpOF
VeofPutVPL+x3HPELX5fP7AYbt0OMKeAjZL8nRZV97uiqxyqlpkTG8/5EUp9N2fsEkiQzZ3q1X5t
UgmmdolbJfZA/NqNb+vrC+C89z6i0mo3IP6aHbUQutteEoIbg2HXY9xKOeIDHPqRi4/0Sc/EG1Lm
lLtadzDmziinecOfDh7Q49gGGEMCkCcI0HGx6SSzgufp7WHpqCnYR2P/kRdOvm2YSfIc9WrYSs9O
VmwOe0pKsNf9xQph1y3PKjtvRb1HJYgUWNoeprkn93sywyPsnS/FLS6FkQ4rH2S33GMvLTIOg8N5
fUJDBATsn2IoiAkc3mh3H5uHZTQCPts5LJtmY4XJ95RtcY258aj3CebuTsl3H9wWcWQ3ufEHHaNz
QK0owDwejtXSGwcBXHPUYktZyFCc3fEukoaLRxQmcXBL7DH4KBHhUlfN7x/gXOxhZICTv+q5CSKw
LsHDyhzmPj9Jzdg0G08BDYQT1I+xZ1Q9uUMOqSPr33nGDVvIq6jXDGGnPo5nwnFJsToMvgjR6Xrt
oM6FIi86DDhNKXahcx8uIQg5L2OCKhx0P0Pg778mNO+yfDDf2v61voPaHy1Wq377fkkQEUJzpa7v
7qgryGq3SZ2+tnMe+V9Nwhy3/1mHJTca2oivY9uwzdnote3OwmHuCsozMUbc6BNWjBQHBvrzEH1o
8uB0l1Omhs+49YJkMHpYuMCSa+LNSOK6mtkXT5eawCqAqKEzUU20SC22JiozUDV5x/Kbdu0xIAhg
vZGlhHwtfogXkxOR3NRiIfl2PFwAHY4OqeUVaiNyEQNpIVYgbSkLr3lFvp43PxrKaNgA9+kFxZCf
8qQJMH7USPKGtt6vxIyIygtfNz1tc0ISd2TWX0yZBMYbkr0+aP8DllfI5iNM4Jl5Ph8HafdYQOJP
9QiFtoyphuDKBKlzu438Zs2pjZMT4z0CybbNCnU6tUv+LQgkR+A9PHHLUuljJ7Nn3J5Y6c0fXyUG
MGYU4zHBrwhKihjs0VJ0j5C7/txhCS50U4J6ms6nJ5Kv3HIjNoSXy1lxMjkv1/8wl/SI8jxn/imy
V65Wg4ANV3m7x2ZhVJDC9AfPQ6Ja48KwajXFYJS2q3Ces2fWUjYtMwrcc5JA5pysVXU+j/S+goul
uFQCaMt5O47qUwEMRiak5akhxQWBwSNMR2RR+AScq/4OSq5y2QLpdDtb/WMnltP0sN1xpuSHXFBg
w0TZ3c4OdD8qvRm0VKjHluwTcqmz1ninmPlLKoCtSiiR7OuDmOjalVb3nnimp36cIWKLBfMSBFnP
nw4K6CUos4q/R6sMNQ6ZvsRk+oQ5mcAEeRc4HNQGdh4vOXl2GDRc9COQgWeK0jjm9vuqkhGRPPqc
ZbI1/512lV91+9tPBFnLI30HFOAkIvUgGG0lkSPeMJXv6zgn+hh7JhBKN1LKCjrqQHqn92UHIYmj
gEhP9xAkqEh49K3iad5geItGLu1f7CMfvbg45Ckrc6H7X1lkwayAUG/l1kUwLtPCQWOrNHnN6Oj3
2rmaiWqRkLiVELZftVtQd95/gGqmGvr5q1pKjjL6UaaokSd2rXw0kD2S/lwLSp3VGuF3Jdr5pFdW
Rd5B7+THYIuzR3uYm9NQYYiJyGZTUfKpYBO9ax9h+sBaQG2lWT0vdXR5606e0E4Pv5PXKqQbpv5k
Yc5OB4v6sh7TVCW2wcyoQYf8VmRLgAK5tRM3B8Mylsu0QlkNCt7jslbP20P60cCYs/JG63WqykNU
bE9Kd4jiPY2SfzjaKrRt8Pt3UOkXeetDWjUg7k6OKmexfhhFGEwlW4Lv1Qet/B8objAzmH58krUA
0BjOdPgiBWoA4l+MTCueSm19oI/TShLERpwwHOKHzlwNZ59EWVzEmVMiteaftqsD7E0J2pzov+UG
ZX9gTyGZxOms/5fHWH+l0DjeedZdgYByzek8UBzvoZtT1tDKJuS+t2wcgsQbHFyQWRMTNinfsOu3
w1QA6+6kG84VLb4OB79y2lMbKK1GfaMq9doLASAcBymmG+H5DpMJCWQibFKe8/+sZUYknBOkSVNn
+0I0dKYg/1HQa2W5nBAQh0UEeAztosIXgmQ8TpwTfEQPrl1DKfx+yUGyH2KlfPGf2yJ97HqkwdxZ
gLMBsKhzo0xbq5Pd34ZZ7VrhWs7gE+UtMhNH2+YobvKAInfkl8tOh1ES+jpFWhah+53fN/cddd/M
J9T32ZICwKaTyKv7vuqXqYMgkGPxqpvmXdKk1gwdUzhhsxxcN03OhaKTpGSbEVm+5xF8y1JDA/BC
Kd370gcCOqL7v5asvBMhsUsogFlQTlK0XKo2BLzCejPoIQl+KJ/5Ap8QXmY2WiK7zOnZg0NuwPQj
678FxsfIbtYDy6lEsnnWGh5TjpwJn2qNlVKnk2soH/78FyWECcuos8Rlx0U2O0smaZB7b4IqziE4
3LIJALw3AYjO0P76JCyp3am8HpoDyyioXZ3OqB4Csp9HJy2CXbGfCp6idWNDpvEqwqhwDxxVZzbH
pOLnidb0zudSwbKePy7PdQnp4di3iKBPGTu4KVxpP7lJjHSFT1aEuTiBca9n6Xh2axKiUlfSvRSZ
RK5cbv+uqXACUyXUkMUDq2OM2ax5ChVUnIgbCPAkYTZstKYY6ViQzJNQv+mOR82C/2riReTXOCyT
E+SexEdSgXe0e11YW6nVFZcWU7fdCwhcGEvAwsnCYrwW8qIDRJnjs996tBQah+cyphIcNIEg8w3y
BssLZR447p6egxoQWHaMpqid+4dbB+GDVu1A2cM4SiB+CFomAR04uk/Vg+pR++2z7NLgnuRxfd2X
Wn6YEjBBwmmUQGxTQCQLY4je81vXWUr8e04DInrpxu4qAIsUrIP6x+2ynCplQTF0EFZ5+S3qkKGU
os0K2xV3BwnEZoONgNPWpixqeMyBqyk8wC4hPAss0P2rbcuab/lTIJIga/dszLQs7+3DjLiQhHiA
YbBGJZAu9oy7m/VkGHik7Wf0+iXfrIN7NU8KG4ovnAj+b2NxbFRw2+NMjXga2fQ7ujHXAKkooqd3
OfInKnrVIb9wQV0Xd2qkdwSpVqFZgThYsZvTAuvKvjdwkg6cI5jNwbTYbS14guJzgCdy7W53RWzh
qlgAly8d8X1/jnT4DmjTV4C6d0X/fiyyFBPxJ4Z30JLQVXLXeMd4IMOWuiWE8MexgG8ETi0iH0hy
rmHXwbJK2yMx/q4Wuh/o0WDzXOO/ymXePMdEi3TNNcb9RQeIRY86sxmgCl/4ksQhR+BsrAPJNhw2
8gz4oGHNe5k5DHTFk0nxLtriOzo/br3rWLHUd8uI544WR5c0usH8F7G1JkDLVacKemZqYImWzcXx
nr/KLfj/iYZj02HL/BW1R4KKgPBbfDTHL6xUAeYyBev4I5JVR3VuRQPvUtlZxFtzfkN4YKLvaZTI
PbtJ1AA/bjCwnLuIpnHueSjkR00hy3PFHzRfUkVzFRWVwCU9wZdMm1NckXQOk77MtYf4fHEZEXn7
1Qhfuk9++/dOe+adNq5goheqHNu7iJ5omOsRxrit6pG1lYjW/o1I8BGW65MSjRVTAHgkSBVQwNJi
hsFGNv9aH/4cUIKvZ9XLrMvOlylm0tuDPthriEXneOn3GSFyDTJtfX7YYF/nRw2P7IUiDzhdauL2
T7kguDn3gcDHRpfMb3aHb4K6DK0/ot+qo2JQO1WiCjM1RV+AWJ2UoIy9WExBVOpLxjbV4zdROXxS
6zMz7LfLmfbyKYRCheiz60TpuWm2Z3KurY1qg3nn4Pg5rCxfs5GSYPbuQ0Wi2vvmkt2yYjYf4JEv
kEUMrR4s2XRJ1FHuUXfMzDPZhZrG6GgdjyzSate9w3BfgYJ5H3CR5nuzG4qr1gs0QljixHSHK9Zl
f9GDSzmHQzKScmr6SQvncaJefRqUp/4m4gEtFLppN6hSTJbJ8rLDAfaAoyIFCyXnjYoTLmOkyIBu
l5saAfxTmt3q5msCu97kMEgvi8AzKXE27Vd5JdwCndrUBgt1OMVX/V2K/aELAr49toUBBviN1bHC
Rt1w5zWgyB7qeJksqgWAYPYALWvsQYJ9rgZp2XazaUwJQeeEpZisqWEOiNar1ybhJwGefcXwWfsW
FLAxVUV3sDM8gXTyTZEwMZKx77UgEbHEThe9U0Q3+CTUWDPyY0BXZyLFf5Ln1YPMCpKcZOqxxp/1
MvzQrKAt5cAeGwdoKYWc3vYtgDgTwOar5rheYVzkyob104auAXqNOjq+VoNsySLf/R26hU1CpEqc
vHTmd2yAu7wlaA0z7BjbAYvoSSw21JimlEaAZEVb+ENO4T9y/B1d4zVkcE6U1NABZtdHSwEs30YP
VotZyr4fgAsw5xbFu0Bzup4KCNIgwdlapejeVX5cElqKML6X/i2fqsItdTiQPuJu8JXzra7DY08x
1e+26aISj/IWRRjDF9Kc4AkWs4SSqjPz/8vRpNUvXXnkQRzn2Dy75cbxydritNfhB3z75z9nVt/i
YB+hwX/4CB8rht3up+rdAN9/8xUlU7UWFH75FdKACJf4FdJXx9pyZf21uFdbgLLh4+KZz0oBg5ix
v9HuyCJ7gJlsjOmHfqQwzrlvUuXHM4vTNrU4z4pzwCczURy9lcn8RyZbWsPe+Tm9Lixtn7ccw8eh
2nvWrd0wkQexszJjTaFes/uMGbLo5/AqiMPlYf/BA23lTk82p4m0dpFkwV4+14bKRGAj73HlO0U3
SljXretxGWIGe8Rh7ZP27QJdhdt8CdDhSMusEcZaE+rUTeZ8deTwxVgpzur2FTWqGlhfl16quXRk
Hy/38UV8ll6h8xUTO679+hspX8leWNC71COfqdmeMcbDmVSTw0ome9r4Mm5TQcD+Yaw8pE4rCJfU
Xh8FaiI2kO12Bb5+vf19PqoUhz/E2Y2AnNfA2q3ejU5uYClCtIVVvy4DKysltCE/VMG21TS0ZKVl
Ix0i43i8QeqhK/ohsqUaB32DppXFA67w4VaxggGs0kZYGOLR5G1ogKnOIzV0AJADtq5qZMInGBkZ
QZmFOen1LDuVy9q7jNlTDFICno6y3zQgHglft+xfr6/fAztWJWNCw3c1wsD+n/PsBCtbgf/Qbrb8
YQat7XQ8nhUAkSwD0IX7zcbR/+vKZe4rT/MwZ7h7xX1bE6LW/u5/mUygcBr5u/rTTfMr7Ogus3Dw
zDfhFo313ytEOuaZ7VBXsBkLo+ZoWubsJ4EmUQHnYESc8uk1PMypGeon0AmjlEofGL6jU244IB8o
GrdtPsW06m380hXTU/CMmBrQ8qcqnwuSmjsEhlhGbET/CXsw4ATJqcMLXpsEKCfLN+frCw+LDfTQ
4nxhNxlCs52WeBpQ61Kh5FxaI5IsmnC89K+nJhpflLWv7SDUKDguHUsKmjf9BoMt/jQ9KDFmnUVs
U7hvdoF8+bL+JoBVMrKS0o1CGaxz4qRDoEDHD+vHxXfBygA4Pk7WhWQtPajhWSfF9xznFPZtvAhw
KP/pRDoivvPNp2EIvHoo/SCMjAWOuzr8/vXP7UXucnDfsslPPflNE95HfAgC0c0z0GvhWCMppJ7e
CUZSy49CS+1bkct7P3QQa5l0Kk//xoICG+4OhbqUCvWgSWv5OEcsc7sHZGbsEk7c0w5i4HZBRz+o
/My0gJt6SmDtSXY6OWv6kXBzYuXrTZE2ixr7LxLRwkpVTgeM+n7kIEEMwsIUSrxXHHxHpeyewE8u
uYvo1T1EE0mOuFiU1zOlWmLktJTayvQYAYjWn1rV7d9IJYpNHZsIp6T399LmIoGnlS77vn6yj8oE
4SNOT2GNcBHqZpLW+jhT3xIlbcfF/MkMGysQ6bY8OZ9FXUljfxV2IaH2QKKNJTT5LfNGXCFJhO/O
byO/BlhSNSQAgrJB5Jdd7ctyjEsXlTnDt2hy5DenT9dCO6VQFH3CI2cA/IS+54UIHdSUAaYxnOxV
FLLUNALUwn11WVd+7WPXCPkGSRfJ7ite7okymIrhRBAGEMzZrO1ucBViLxg2AU05WPoRM1LFUjW9
Ywm+YiyN08XJrFCjltXTkYMtmGEAfwoe2dijx6+ZbfKfkPFzWivH6kiF/CfZsN5iednAUv1rvFdT
hemMo7wSXuJL7boyyiSvI1thBJKKqSQaIXSI9Jh9OfPCdOciOFYZM/2ZXlb2ge1BjjpQKQ+h5//8
jtg3JSt45nJawCoHk8utR/WTkW2fYDqERRJLKUdyEzRDQT+ClFsMzarx0cKf3fT+Oq5CdGXzUQcn
4B2/i6SrtHrHa8Jkig+CqhPgGJOWoK4TNrEF5dXkXMS//+OmdZIh6TP5GZAqxeiEAEw08KmtjIR4
8pA4Vh5j4X3F9qw7NDPyiKNeqdCBuN/Y1rp9qgnu+4lRrgLqPP+BCtnvEFrwSxVtFGPr62xiYW7J
rCNAutCJ7k0LJPpyspLm9Hh02FYJ50c9vRjhjqR9u7gLZPS6meC3Yu6Gcyb8RQyWQyend6nMX13Z
RP3NN58pqfjs1uR/uJrJg5NNghZsvszjQKWJx1lmhJJWLGbz3zJiTs/BLza1AdvFb0JBhMFz42xG
rmjO7Jl6HIk+9sz6WckgP3odHEY2QwHDVbj73iza01G/ctKfTQJGUwykqLk5uEhAEA2ubhBQuSrV
rM7rmQ4Vnklxi/gTCDfLG36UACr1ws9dHZKVRR/5qKMgPsJB0dd5nJbDntXt+ll4j5k0I4bGB0kv
wk75DzPxZTTp0Sz6D7YPl9TgjqHyR550122jvxxUVcz1HKc9I6BW+eb+NN7uIXnXJOKNPJtAW8w+
h92lmMSvgAzntAyPEF6rVFd1jyRfPrcjaM4ZEk5P8n9oxvQu9lHbjOg7R71UpLpVG2NsOR/1DPut
KFTIK0AXA8Gm3z7wXN3dvbtawhqlzLvAHSPxAtlsWzIZdcwcLZgFQpkr21YnE9cgj4eUGguV0dlH
fhizYNi4ZIbgL8imrz0XIYRWFOu0MQ/TUEgpfucy5LfjoiY/pEQJ3s+y+yulHvO6Ncw9SJQifJyz
wc7RsAVCZ8mHfbQ/7MREmtaeHCHURlsKV8agnAdc1ruu3uGFsO+QvgO6gg3Vq1lLW4SCiwjTLlJJ
2CfO6W77T5K/i0y22xTOurkyUVTVpG7fN3RlDNcq9RuRvJ+yQvrutGdogHdD8XkRr8Gla4AkHE0L
HiPoLsl+vlZ3oldfykdqNsaoHMDmrixk59SK8rbA3a6fv6xh+Ao76IcTI4b/wI4psl1G59959RTZ
5WDJtkD4GwALapSRjkhglWzWc9GrhYGTwrpadSCSYLj1wjsw09HdJ6Wzaxi0OB05xTATm2z8rHU0
3vctEyHZ8Xt8Q4+fR/HOR9cX0UbVW3Z8hXeZKbRMCErksnfQESyLZ9dOjmVuoFeaw1FVrXu0th4Y
3k21zHKH/VssZvsUGFIZwoiJsM/fscbuY7Qpq+7YSvK17Lzh1ls62kM02zjPODKWja8babduo7Dt
R57DAFqejxx16kybbuCcZR2/Us7WEcUnhsRXebc+HXLXz20LINw3ICWnM5YCl2LLA7S2Kf/XQqLz
nQxWI7p0i5UOzwIMOAvt+4XKQzFWN3mfxN5ZGrWDnd+7IAAvST250DrgqFmCudvgD7u7mBJuyCSO
y8f42whuSklauXNoXjhROeoYu3liRDX7yViEhvsurHbYDLXXpD/PyND/P3YZ+GkqglQSjKwSk4Pv
3Ggx1/aOCRa2UfyfZfsjnppZgxv8n+VcwpZvdh2/0yCZLnnHOGepCWEn9BH0SnS7ehHqyd+AE0pG
dj/+ZM+/OJIqpxNLTAogUZeh232mHp7Ypy4GGkGF9dhNBu1oe5i/3ppiJAoQf91kN6Z9Wby1aRo8
aP26eeBfHoh5T6LyZsqdExra3oFKvAPBHEZ9a96u9Si3GhPrlscoVJWZNj33uiVl0eKsPq0J3PKT
BK6CCmvZL6hMUpWsTYyaaC57BqkOI4Gvj7EQwSfMZIzBefKt2NmZ+km3Uy9hVLogpYUXDRl3g4Il
Ri7EJK+h1XwTo7oxT08EHlVg2QzpXwkRiVRVAfVCxKePXG2Xc2rE59LV0GnNtocpcLkbNJN4p5IY
GiKaxlNB89dkp5C/V9UgNn2ytlqG/1JQka0fJxdGDgZlTtwe8sybXUvr8uvGm8/ivVC3aMaI4Uiv
MiJ/bn7cKyQ6W7QY1dwGjeJazFLtVKptT8+bbJtc+ZVvD/ktutlPHllNQvjZA3lqO2o/pF2kaeS8
gHkQKt9RFetXi1VKene00Wu1wpuVyqzjIExpwhZnXaNdtBTfMuuiWcCOn+BrN5OKPbDxeHRj8Qm+
YT8P/ckaHE0b0Zt7HfDr9oKJuIbuiA1KcTAw8El0EAqukcdXhTQbWIYaPSU2QjVrxCV1DVGZEX9K
w9qn6E7ff1giPjt1+RRQrJVw92UTq23NF5Hj8OsAOSK83dfqIej6rL7Lby0yDImpkNn+/njVaBBZ
xQ1+0k97335ASF2p+ONWCM6wCAzHTVbjupPw92KhqpO0WBsNil35CXrlbQQbwaJXTUtVB0NpAxIH
Bj7DAf7rEYwNNXGFQQetlD7fwLXAxE/F4WYbH1IdwymKnDWosvvAgWE7CWg1m9LeNFoHJ4TgMm61
AUEuLOUPXmqiTX/PTgk/cBlqOTnXhBi0HKCUj2V2uoJlmyP083NTYMcAa317pQowa9HqYj9ZuYAB
YHh6DZuaoswM6AAg9mVkJfF+Sl+9rx0VXeSPyCDLYL7L1SwJp7nWAwPviXmZEQSUmCi0NDhOeysW
0zriKGEi1p4hQrTzl3VS7iAZ7tBwPIkB2ojwCDnDFu8HYxLeOA1afMntdmQr3ww9x7NNWvepctDh
BhksG/ZMfHitj90o0+b9Rrv67/AjlYsHvXxcd2vUu/EWbxAnOoCXMrciLL4yj8sqNpt2SnF+I4GR
FskjxbVOMN2SdqfBDVjTi8H5lXsn0cwNtVEiXsTx+BiaR86Ipkm1l7TywJ8C4gotz9CV/TyECndp
/YP7IQbQ+yhMtRtn2E1Q/pPwrIyiBCCbhohRXwN1hdiiPn4AaqNFT6BoxvEEKBGz4MNJokHwhAte
1zEFladuQPwgV2MQ/rst17G45G7ejolQklgnsGVPzqNwRGxt+B0OExBQnMZyQ0UxaLtM+sqMGdN9
bIWAw8+bCPBItqbAhR+amwQYBPwcMwflT1H7kdBxX9EJvIE5PQaUU6IIFuCqMYDQLAINsAaDZhQC
df3P8bWYDTRaDIflF4+mJut06235MuocaE9LFD3Gy64LnByzswdRC7FC/1Lg9yCcsJnGAwM89Mzz
yVnSQ3zT2QMWay9zWTJDSCRlrazeddSWxjsHpyXnWEfIDHbD9Tp0E6LROrhIbIGrYp9hw0oj1C4w
joN3suIOx1hJ1olmw+oqxFuHWChczUfgAXJWidlzBAigoIom+NEUPZm7Q0YXbZJ4F7PzC3Sh3V1v
6Wn1yZBewJ7KVcXgdaWi5b5wuGGTJJgwjo7/nICbc8un61lJJK00rqs2QH2fVCJwB4I3Imny/J6v
T6OQtajGW3zNiAyl4oFJwprXW9/jY1xZxlkvKuf1UPuyiokrVa1S+56H+n77i4sIzfnX2sCLLpj1
2FHlwPr9vDyissVUDxh7FzhMEy+zMRyKKV+Srun4pGAGCL+3NCo7BoGKno6cngle9VhxyAligsPw
1mXwuQQ1GC8YvHMnz6X79NA8HgjHkGel75KJjoMM46RfWZe2oAHJsrwbE3Kou9mdoGTwCJ1zpZ6Q
HKVuu1qhwZkslsbxRhYKH/GxWSw6UPc6g0LEajy40HnCp1607Brv9D1EdXNSRD74OSAz/rLxp3Ss
mvGtSx6LaTMaWet0xepxmdTPWtEOXIL9BRNChe45cUxwWhvJJKcH7hNsvnkUeoVQb8b9R70ukcxj
vNT2Fu99o24jwMrDsntqVFjIMa4AMKc5tix9M0PEOQZrLvsJBwxo+UDUae6lFlNe73X80eruO9iY
kHZFanoWGYbC00whwURgwVK2evFfsDpCzTKCSSN4dCGMAUcOQ0JIZFWHrezCww1Msee2NMc0QAEx
xs8oJNLF/OqMPRmTUxJB4jvzwGUSYKOxlbfvCSFRyxr8tu2J7Elo8QbiZKkWL759G1sjv8C4lwk4
cZ8KxJffLvyx5ehkCAvUJVkVhQWysRr/Z+tiziH0HyEUsUBsl3HB/duipYjogq3tDupiaxGjjVsB
kWMJ7LDAJ+QMPZHYdwl05eiFGv/+hkFf7llaLtGaXn1BMOE939G9yfvK+WzWoB5EIfZfUwHKx1AH
FBka+Qdn/pj0TVlpo6v5yHK3bBT49FQTNwqTbWDk5cY4M85Add+Tg9a0QkJNr1k9b5R0XZq2oRlx
zYfRNVsFBDXtIBWp37exPQ5/c8T9fHBcActo1C90NxPxhZjh/IfKZNHJVvJi7arbX4Le/Kiph8YQ
6yZ7/hs5zr5aD2wqyneoBhPsLhzBb3Hq5LL/JW/SI51/HUyXKblGnGOQOjtvpil63uRaNbVP5qpT
qmCI88lY7XVpug1AOTZSRBVXWvjOCL+9Ln0Jjd9CNyBq4gYa3FUlmaulxVZaMcF08zJzpADgF3Iw
LePA9sNMwssvlvpyEWCRLdWWcbyhhkYGxNTArSR0WcrEolIqwUfrRmjz+9LKA0p5nJuuFsZ7WZ+x
uhHZ1l7Em8f8myFzjRwmj5YCa6ppZ7mTiIj4N1hEsX/l7d5CUYLeWA4RFhr4Ijrrr/kDZPt81xUR
iICybOOKRiNfNZkTiIF8Uhm10GN6ERKYrmKjUDNYR/lmSwGx9aIhS4UX5XSyyL0jH2NVSxo2O7Pk
VldmyGSbSrwowckY9N+LVcpeS7wDhhWyDyPMGvfE/icBK17YUZFolvh9+NsetVP3ZeiZKZ3/OeOu
L6kNS6IvNna8wj70H4pqU2pa3SqgaIAdspCDJ/rrru1IzyVMZoTBBrT9y3sHJUf5wPg0+edbhf/a
353k3jM38fxe0iUS4LvQdSu+VQmir+mRWhcWP/xfVAHEgzC95mUSe8wVgx1XKmLQebdFp69fuOxC
bRTyKl4nZTTcx76rpcYDpJA7i2GUxqIyrrLy0IcppPqGBUH5TycM14eUVDyz+Zid9l2ZOB6toK18
vjF35a5QyPCh/KXqeB2f3H44ywTQ+3VaeafVwq3JKJw66Axpk99m4z/s+wfPMNwvopdDaNG+2Wmd
G3aU+2ruE0h2NrX7R/9K82tUgGgp4kWkXC/EYEblrIAVy3d6Nt/QYuYBob1/9lYLq8eqG/uKTp5A
R8bmcDpLPDBtqYUY1gq4+3LsrMxkEpdrJ3amSzzBD5YZbu1RYUlK4/Q7v6RLajmj7zlPt3IkEP8X
wIISsJ9HgWloDvHan5dOp6qLhxxWx4JjmNwzVOT2LbWG0JdvHpk8BBpyRtjcnRPyAwuGxbU95XV4
tfIOHN/6fR4WF2y27EoQT+EnbwkkiqLXdMp0CZacyjxRkWf5xa2qp6Q/O/yvwylrTrjZ73i4nLV1
znrDYPaxf9b0F0kubhMIfTrt5+NxajYf7fQFlSQbMHCMCaIZiuJu8/nbb1SL+VMDtPLoBoZXsVuK
4eUnFqvezAyriXqDvnRFycN0dA6Mqb5duTcqUc/vNoTs9bqdjnzRLg9TbrAIOFEHK4gE2yy9JcsZ
Img95i5zHIp8ecZzEz0w0dyqkZls42WbctwgwvHJSbj/88BKjdEPePqwsKq4kIsZltwPiKJxvOpr
KXqOzd5cOPD4LcWm2lu/JipbP5S/qKmR3sTH6aJjEKYAWexIK7mkYO5i3f7rncx/YQgs3S0RiTru
FlN4VR/fr9iU9O9rZEq11XnmVvGykGZbbnJYOeLOq1rVyEwXsetB2F89PaycUT7iHX8ztH+iOxOn
GgI4WcaMm9EOba/JEJgjfy6p8pK1dFOHzMYIp56mDc1ifBClJQeA/rboL0BIAvDU6U7hs2oMPVHD
6sD1eHDQ+laTTRYt09Yu6uWJgLIQp/ggiEElZ+SzQXNKGU9c6ELVX3JbPQ+A3wItvrf9t4XP8gkq
1OdM6LC/kDjUiiUEgQaGoWUQ2qvRq46KnT3n9Asj06D5xIfb0GQXk38Wu99UVR0Od25vThh8cWY2
pplldISC3s1MVt/xYy8knZwP9TJ5meEhU10aUO344VnztSDcTukezsfchmNM3k4BD/LP3zxQhF8D
13WzlU2HrevqxdM0s2TR/qW1/YRf26KOYGfbxezCwSYXkenIGTnrHAxKcKwJQfifujwCZ6kAUNry
cgZ/bkSJPHFY1u7Es/6iR+iMqC1Ex33Wx73ZOP/9RIgSZs1EWbYE/FB981s3VNUNEYzw23FbBalz
lRWGucohbNqKbqlGkkc21TFR9TfLsNMA33uUqZAL+bozCvUwm+rc/33gfkXQAGNfBMZ2hIh0TPou
iZUVNRtt/75iFXCQwjF+GYjbKnECyCGLK7zvetp210Huh0wi/FGbDPEY8M7XSnba3yHDAUGPl1p+
VZMNPRR+/Cj9j4PzOvMeo8ZIj7L0zFHooQxmb3D97xiUbJx+LwPFgxL+izOQwE6WHphmAB3AI2dq
jo2epfhG0um/d32IwS0WFBTF4461qtp9yZjvnObE99NGTtm0B4zjt9JSHGzjuohoEmLe3l6Q1Ogx
uXCe+9lRFzEVJbFL5U7PnbQOoPejtfP47cwE/+SYkZwWLsAp4xT7X7DRdkm/VKl0zZHODO5WdOp+
6IK8OVnmxpmO5KmOhFLO5eMj5u4uGJ2iJy3djvXQmO8Y1Swm0NJTvR07BTSOm4f5neR0bjH5hLGh
JKv2Djs0XuPZJ7mMH42WWUgGK5K6spNv11Q5NKTQt8MUXNU5DwL/04V7ZJRxCCrG6FJW9y0p/oOJ
PI1xdg8Igw++l1pPironfXvrYwZAKXMY/QaWwl048/aOIGKvSIh8emIFbCClmdQ89O//r50JzL12
20mTa9N4jeFseaYBDNAAICMrGbqPLe5SXw8GnE/IPZ5LU4PgIUopO/MLpaovGDdIK+zGJj//jEQO
9oYrtVmosBGwJd/t5WH9mt1LFS/cHfzTPqJnz6DQTHSL+C+0HXXY/vHwtGyTKmvkaECp85R/Sl39
+9UgaW5ywb63ZgvLA7nqrbOogT5e2dCf4bnWbQDtSkH0nC8/zvGraOkzqAITkQQaCE2xg7I7frt6
JksZVEDqdgcbCrBc8/IMAVcFX0QM3UyFrbVnB1Imdvsdtv611Vk2Ltj4r7ygT1pIRuEYa4O/sfdo
ltSyEaS2WG/qt3OBRwSjHz8MO0mC4RWeJdTMFNcVDIwAjFegVWwuiZtIsitdgaNGxF5MRjQq1JaI
gztBWS4d2uCJ2M0cuVIE1xNS0F7LZiwbAZ38Gy/IjwJpB12Xp9NM36A5BqWmUjV3UE7XfOaiV9gN
MXgapEyRYgsQnIgsMvrg6Fcvg5ixAR250SsOfgw/EZ+cVDMlKkVgzxmVBz3DwDTTY7ZyWUGOXDwn
ByeLs97lZi7ihHsBUHggKG1Oj6seHDv5aVmLzwqdd9N2r5x9nLBj+bwl46fJaYGaql7LNERcVU7N
IeduMHzsL23PgsGeIaV/WTuYDcqg4G3j2NjtLDonbrsEWGSw0/oCU+aSrCCxuiQexx7NWfdT6ilU
txGJSFdY/xkLXnZ+E+2ge996yHbw2ytLzlzSDsKduLsg+T29+JyPj7fty7hSn372swJ2ywDpogqU
qyxv8gQQIvW5E1U/XUzzTWn2YBqEGrHxcnc/rZAjTCE6hj18z8sqpMXqaGJKkJK78Fx7y6FOcEN9
MwYJobrXi9JFZpVfU2o9JN5aLrXaIuKhvnprdyETLM5wRBP5haWPCZA20OqhFZwZwyh2xxBgtsXc
fmrw/NK7AyZoMkqJmziel6YVzCzHC2BxmVfeC8fg1q/3Sgj/mbxYTKDc+i/h0pZTb4byM0l8ED3M
/WQfeIcKUxstFHwm84cXv0ClEBCuhzu2zy2i+U3r57i5/V2E/N01/tUfomRv469s3gdfP1bP1Fxx
Mm+BnEBd19ZZZ2i9Yf16Bm+E3w9g8s50rg27uUsfz+fBytNjcnCr3FTFXJJM9DUTuR3K35b9rdyV
bejZtjqhVeSGzJKFAAY3LemvHgyMbfnZEorB2eMgn0pdVrwHyAQrsYptycdyLzay1yXnpTWq0Ju1
uWanD5ElNV3sUL+NZs1sCPHc5GVwVWsJYk4xt4reAUHQ1YCghv6L09dvy1jDE/oLOtoXvFjDwSqm
sDx6uc7W7R4zvhuptIpRUiOCj61KEPJ8CPm6BtE1PHMI/wQHVN3/g/0r4GUJheC9M5ADhDG5qQtc
Yepl/ENXNLFbnodl0g6M9h0mdJvk+8cveKou1gVast8j/liKwjaF3WLfogbF/29DYLN+I+7Mzn3B
xsL7UD39xiUnf3tBKuR91FPisUCMr7lMHwFq5C7+g1wekWJMeUArL1DZK3fcz2SbSP+xkAW7ICem
hMOkfCDksP9C9g0fKjBqFndoYQXTHzZsuxzqzlEr4P6lcy6nw4X9yanUGQJMgvuw0Mflc6zx+6vM
PDB8wbRBmNF6Rv1K/jgLRJhx2s56XvfhXJBnh2soutv3F4LKOgAlxRDYU93kXMBrANdNUi6Iiqby
EDjOyXG5538+hpGVRq0B4cNHNQK8dpxt0D+aW3MzQN1bjRg63SmZMva8Lug36HNkCcY8o0Vl7GA4
nDlVnbqGyFC/mHHy7/+zveNaNyl/tlvUFq/VJLIBDHGW+W4PkK8TCd0J0HibR4o7gS+PJBHbM4AK
t9NCODXfVa9CjEJvJ+2tgX2rN5kUrERaG5rGKcvsUnPySNrIlOOIzgYmjcwWLwOY3W+aZVmjwxBP
kd+wGATkn09OYAK8sVpFx4UliqXOOaKrtNe6lwj3LfphVwulXxq580p4hexcqnYzB3bq40drl/ED
cktQBdp/r8hU0y5g0uHwB92Ase9OOkBl/XfgOHI83XIr+DZtoEcqDK0QK/uJQHg+Rn0vq28YLYIR
eWWXOn939JWnV7Wds3EgTzxf7Fvtv07iFOFUlzIbjSbpdNppAUrOYGPJOeDSejwcG62s+FeNDLSc
FXusgZ6jxV1KoPRLcoIJ/DTPfX++zJ6zOjoITuIz2ihT/MlCTbTaPWGoHYNHyrAeMR9HcdbIb3Gv
/l4MDizrK9Y0mulknFDmzLAq10XXrWbWAxplQLWCPNc+FKAJ/TqcLPOmGdmsOfvP5fVaX0OHXGiP
J6IBC2oMzV/l9UWZp1g3PNpK+Am/+AEa6ruvjuvs0lZJszCgJqpKN8HCxr61dI45YZA2gHLJrU24
17Ci6HBUlD/XKdujun0CkJP4+8D28Cr8piZHxQ3dDlCOA0Xibco04GnQYQVt0fDRlS4t+mGjkjmD
TZW4S8heDe+Smk/MYCmeOvcwpkYrTU/3F5WExYJsOteCgk9s8K/qd6h0RkYceYMN+j0IQ1VyggHW
tt+JRQmcPdjI92HsPb1EUHDxZsK0sEnhCr+YFrO6geT50ecILI3ZV1lG/08NrJEoCkicwRySrTOs
wlp8MqQtccNATxdT33RpgGzzzcAMGkcvcfJAYK0MVSchpNCPgMVYJmT5gaQ8D26GObEtyekZY45q
Gm3/t6m5truiH6sBJmpt6sGczDdp9CD8zVDlDAkbKNcQz6iF5TsQMxZtGf1U/kUuQhuWvoTr6lkc
v5xt5o+YUaDGnt7e/E3bBkuO22oLo+RH33YVo76tNHk8ddEn+nEKxEPbZEFzqnCRbujdcqwNsU8k
LResC/ISfpsAcj+YfnyQzwliuOY1CkhJenvECe0ZdAifGIkaXyma2BaEsHUkIP2O1WnE0B5ayTwp
abzWcjKMBB9tVc2+EcomirZUp0GgukQD/cBdrdEB7iPFuS6F25PpdbLkSSmHkAeX9vxWYbr2sDae
DD6AwjPWE+ImiCK6P6J5GzqGShzTdstAByIraRUefZtlbI1cE1uLnzwGe4yvPtqjweLXgetot+We
Qzr4oce8skir0dxG4SqGv81dtdoyvnpzcqTYZ/6qi3zjiQM0BoTsY0C0oO+l0olfUeIBhNmB74T8
+1+oe0uINI5KdwUgjKYmIW69EOIpf2/QbC/DLO9MljQZgd9DMS7+qPclPEmHuIN3AkRNn/uWWZra
qZtUTdAggQQtkPBwB2jidQ41T4M4/bKBAY3KX7u2kyrv9IFcnk0PB1e7XSdMNAo2Qpz2bdTaNo26
dqsEvrY70cxNhypK+GsjUK55sTNyaMHiNraJfOkuRKFifQtjzgNALEPWWxV7ibs+i/OGHnBTG6jg
OdVdH6wre/PkusHpS3WRnp8RvkKyG8Jogy8LZ2/MabRfZvk/EPwjLrfG10amlFr6Gq6bFOgOjHJB
DmwmuI/hrw8kSMztW59Bj6wX9K9KfH2QD/7MrVrPunBIFAT19cYv+TRYVVUddTtBsfQwWOWkqpKq
qSLkQTukVifnmqCP1tUt6JGWftdXYXx8kLkZoYDc/2LEAc6dPEgZ61J9HIGxFDQRS+zZC8LhHSFb
KmaaUX2c131mAbhL086y/Mc9pEs2ADK91qj/l3E9P0sf92LvxboJOOPklMOGyMcFRcU/1UXH1Va6
dw86Y00b6OP/XeCeClz0EeCRVUGqxuO/oGyMq2w5rmfXpP1RVOpMUO0Jk2yn+Y4tTfDOUGx0OMBL
5GZaSRx5Dv6/8GuA36BRHArDEGjisBl+d/GBG9APMW5Zx4KxJ0ErCDq1oj10fAsukrHO7InvO3s3
qB+vo+qPhE4szPdDPloN4zZnG1jJaiTQcd5Wo1dN6WxhyVb1BZfQjUJ0+bUUKxeMsZdI0KisnyaQ
+O4sKL5BKKGcRUdYnSoUpm41Miu3ELV7Q3d6y1o3mFGXCRHh4NLT3MWLOwIdgJU34QWYLqszfmHx
j6ZNmu5I9s5LGJO6TsPNJC8naoIoa5tTSptD4oFHAjlYTh1VwGkmLVod/cGEs9stiJEwFatUvpRQ
KAxtxbGTSSGFevT0N5SKzmaanGyKRSLdNYheZEr+cFaCDlNmacAbHGjg5GElxVyuEVCDkADGpsze
ofk9cfp9n6Js+6ncPEcayjrJiRI3JoDeuCYRM0LUNF/8dmaCoPinZQzO8KjvbaUfb2ZcQ7bT70YA
9VL5aX9GKOUSZXFBLC0y/wYAOrifqV+okmVSZ2VFXzmbDninVHtbPUqg1Ogniq9qipM1I4pqr9eY
/dRZuMkLxTEAAAgHuFPB+CilXgpBuHSHS419YbPyYm2WdJDsePXuKbnr0QPLItC9TsE1whGp/ra/
iqKf+1haI7u5Ycl6T/im/YkFHwO5aQG557Gfj55zyMoI6BLow48CRxpkg6s+M4hmVgn1qnqXyIhJ
a0MOLxqD8Sjq7Ve2uwssD1gt5NkqzpxYICICz87mRWAGZp3cfJv2hcoNucoa+cpsXoGbdmmAvLPt
Mx2M7BDFrPAWDkssG9hAKtP1TB45JAPNJ5cXzgBDEsx9VPKeR/53XrXmLL2XfWjm+muiPBPehOqz
ifhrDnDKhS81c6dOO49LcEKvKN+Epfht8imycgpFbefOQFttzKRaBfdHBKdTww7HRi84iThx04Rq
q2x7X7bZCpReQsNm/WfgtIUyLSRadmNPMxZvtrzKVGjnkkwWKKK0Er7dsvWu9qVAo3KD/uAX2f0W
Yr+AD5vdMsSHIRiGZxDuPFHBJAruysEo0ZuNG1aRHLcGZiGytMsGyhG9ysuGSv3phD5j/usEHvl/
MXBkXAWe0kIVyKBctxpcWf5h8oESNvHPzgFM8dZgjkFpy1EDsQdBwGBJxY7TPTFD3nq4wBEOZbn8
OHRDi3Z4vu0akxnhzyxUnX1ghcYXrwAvKAJBClHJ3L3itXNucYHLW0kod8e86/44jeDduHU0qdTL
hQPFqWNfHQ9j53zMq3Hyv6Z6BuoG1d20vXAkQqc9SJ9C3z6D+/sglymYsEs8r++M/gHcoGIG3ibi
8CWef8eaqs7BOEzoISkHJNyambz8Bgxz0g3AcI+phZwGiZjqYkAi4I2wVYgKL3nVjJVHLCw0Xbw7
fE5axaQi2/p1bln7HReO+HJD61W+CEnXmWH1qpxZqvSY/2dpewCL73uIMP+KLdxUzVTQ55bO8BlK
17CrkYrwbWoTBKtKJEUf6mYzKz0sAYAYWdmziNwhZPXI5pgBekvYL/E6Xd1yvMD3KI0u34laRZGP
YVB/kCfMd0mGLjiKT+mLhEe0ycE2/RYncxvNCq5Lsg5ePGqkTqNcwNI0y2jSTDf+TOQD5stO6b3w
FFsfQZlPl/T2xw/YQ3OLXxL9LztYVSo3tcmDCuVO3mGoqgQn7Haz6y0zHkwbIBiIdYSLQkSE1kpx
uUu9aPso8fdgKOSzeJ9EI+2gmzuSJyvFfQGyjRhtoLUnjPqkIXuEIvBsr5Zj9BAUsb0pcG+bWVYN
DzbIZs8UVYFRz1x/VzQGIvKP2HMq+3mcsHDP50w1c0OJMCiNdqG5wjxGOx8V8bvup9onztKROvDa
62FaV25nb3QpG6in8Arom+2EBp/cE6aIjzB+vVGiBjeasmxmZQoovdtT+HNhMA+kChtxz3BqfZq+
LsfekOfkZJZ9XSxsdDaZE475K4vxBMiGsChGn8nC8RGgGlmcmpjDV2p+J7+V2D4vZ1zaydrmqYcJ
zmWrwIWPYyOs4P7Y1KhmrIeYbT45XS/ahAZeO1Myjx92O/e9mBhoiDFYqrF//06CjmwXSorg/446
9j/DwCFk2qwbk5wrLuFtF1ijpddVl7g/DfF3ZQYtw8brdHIxfqr4Fpm38qCeKNwCYpa+ljYdWP9f
kXvadhub2X8vguQk5xB29AYDL7JHDp6SELMkrJoxbcbzdYnoK7U0FcK2hpNmQ/0KZUshh4lTwQkW
LmhCvtuuCoo/kBdcz5lAYMujQ9Uf3ZunBgl/FqYYFyehhmCTFq/D82W/QaxvWp1qEoNnbWXF0v7h
PLo24Of0TGUR/STF/fCpIOk8D1pt4rpg5zIwEJ4GEsM7JN5rivLSyPBi3viWxqsDaoXJs2xDiQjT
m+18Af63hNERxVnoBtncyHruaxNIG89LP+Wye8g8oBzrJR41nPn8/eOq5OYpkc0F0rLCqdllVj0a
i2eAjIDheMr9JokbDlT8jCUTV7ojkjdhQJKN4m7aXJE9v0EH+alXSjxpy6mX9HfQdab6Du3OcdKs
PW4NEfFgTde3lNkC3vB7sO5GzgDR1pAgKslX0IeNIhZ6XWd+EwKv2CSXcy7tnFeG83zUcxY0Nvly
dQFp6i9t5zelTuKNu8Uu1Gv8dnJpLG/S+J68buyR0R2qd+dAsDbhCCs7HQKwgatfM3pTepjKtBVT
gPvmJYqg+7EHRu+xQY4Uq+1t2eCY9ObWLpeJfyIgPKKurMC5xB+oMR3WsLNSnoVLS5WAmPFL1O3n
NFck5Oim/l88BM+mpmcfbHxU7oVfQVek9SV9xjdMHtxwfBaPCwLyTAVTd7ralW6GPfpV4bDnpo2h
a/WjGSBoh8zoxJdYhTeCO5trPksDTIFS12L0rDd51uqpwkYiKdkort04eC/DFZ2dEJifklKhth6T
IAvcm0p6Okss5XoDTAfGq2rsQwS94rh3C6siDM8YdmJ6bdMTjjBLfAHbI3f0eDR9go9hn0MrDrjQ
B57hh/gQHi2/bktvJsuerysoe4gtVinbsig57lOcoSGBqv03AFek64/Zo3TXBO5vgiGD8BgqL9X1
PfpweMoXVFYvALZV/C1eO9Z5LzuuuJgGlVMtYvlpmatA+l3Y5ijHtSU5jmvgsGHvMo+9mMY8J2cT
9cwkdpC3lH3ZX2q49NWEJbpa23t4icteARu2c9RjG30v4Q8wwpdjpjRtb61oddmL/owz6sMGvytT
r/e9oOxM+bbY0jdi2MM5Vi8aBijGoi3e99m9bH8at+WsvpeTAvXlhkVnxbuu52nAPBSd31MQOtGx
P2bjl1Iy3hB2Y3JNOZcZMlXRQgfAVJDm9V43GaqCj9wFGbVECSLcE3zDK+bBLeUqkPmkfPeLl27z
XKbRfimSO3RgQPhauRG/wmc0P0239hPlFhVdZu7unYovZipTGbsHH56GJVInmpym1C1xbSLUVbSO
v+HCCzL0XgbSK5t1XdehH6riAaRmfGVeVR50ML8iYGn8xjrELZNH+gFNMJ8ZVs6QLuOxXp3nI7RX
2fnKVvRcnbHw2OulOqZ02Xlqs7mcqXiSzMrLyGnmGUqHBM+7Rz+T3rMtgrqpZmba+xXsXzcafQTf
Ul7CtBurKrrAgkwYYRjcRGo0qbW34r72Pdks8f3l/1ZoKPHJkmi8xPvKbh+cR0gLF82aemZZSad6
HwQ95Bd+9rOjLt9NtKVH62rfvGuHs/H7gkf8PcFlKdDDWLP89/OXOjrG6S27/rdhn0ebAk0AQR11
0rWmPayG6ysO5NofFQE7tK59yEO4e3KG8y0PUUgQyUXZrggHEvFBmIpriiuotNhHvPRpol50ZQiW
rcBJJjPN9zANkTIAQtfXYqsXhW9TfQU2utVPdU3OAxsyeGqzWRRkEtyJ8HVrICXD1swWfHO08eI0
5OrVtiJLMo7PGbc0Nv9RMZT9XhrXH769Gig4QW3TYwZG/zdVOHz6LhMhKFKNMtCilS4b039MZDeO
nnjiu+PamQTgdLWHHINWoQN8MH+Ec22XzrIBl5abADowsCHIWidjEGofDbrRnM0qphXMA7jQIQDZ
RzkGcanbVcfMnOorj0dOivw3ujUR+h+i2p45oBaP4vWGlySpdnArWqVNQRu6rIJwOE1w92JMtDYu
FQioFWebFK+Vl/IikzUMO+XHjXFvg+LEXywursoGK8SMTbyTG9imI+2io4fO+fcI424ozyoPYfWU
D8TjpPxE5PSdtxuSWqjPNgjbuX8phKY7daSaDOyQ3D1lnopZLXDEsT/cNN3VkxGcPY5CR5hoXAWV
hkpx+42y/JpBFXP35D77MoiKmbHYNUrBwKtRfNCDml6ZACNEexZtl/G9MWsWhWiROIRjqtryNZ+C
fcWsS+5j/hNYcSLqCfyI5loURaADzAS6N41hoR2NCn/8vKbqVV15Ar6oqpVWu6JSe03cbxkJdwJb
plWxCW1qRjQGStw46+Hr2PICPVdsxAKTGJZQxOyN7gMraPskaFBS+JGU4jOYJtYG5z4jTqwFQqJL
3aBBxtwyOinkGpL6rWYHwHs3fEi/CW1uptI1LNV4E2dysckPKCt3Lu2mzB3D0rJweWX5D6ANGWSq
5YR94Q7B5gj3RGde1DYi61JOWVFSj9TC8DPlv6jDKIoKqj/hyjRGV/uWfoyoJxkn4Ilcdh+s0OgD
RBrjRq/cczlqZMU3N6SiPTIdd4hImCskTuoDXkRUhknJchagaWlQwXkvR+YOf5YKdbxYV384IZw5
yBfNIerb6TqgH4XBqAJlnX6qLwPgqTPgnFPbHYdtNRmXPAxcwCaE3F38QHOA8Gun7bmaTZyaQkCK
CGeRvad+c9AF6xnbE74GnugT0SOD7zWMXJ1QLNZAlvX4gp5Wqnq+ylir1PAY/H17L5oHsDvJxEzr
deRiSyUDu1+l47T/rTUe8t09jEeGIF+RJy0z+TCPXUadhchcHcM/5+RjszAQtP1Cmw9dko92T93i
zIF+QAp/X9n/7CPv4Hjw/xL2sCGTOvQsWwyDxM8TsYoX1oTrKLKHHaOCXgcbgDCM3W4CDW9c+ntT
5eDomfdK1LiRhvTGC7nvQP6hxB/2lQfxv7SK6aNe3caH8Lqsref8QBecJMoKzHGNzBfWZpZAjARj
2Un4sLNZV8wGvhM3iJQBV4Fcz+0579hhFL34YxvR4/r0Vqpx7cMeCiNOvMZ+GpWsk3UlPXFt5xT9
ZBPj/QcuIxB/Rpnyc/KnBTY1iq0k6JgPi3W6HmxBg9+BDXsoGle1IwGREXh1K23xSlsLKCePDQlm
jdPNYbUVO5KtFnGIMOws5zYDIvQ/qtYh6oiEX7BS6kCWGpuAbGpgNv0s8B5OIqWFTpEqrtkoR5tn
7IfHAcWsx1+A2NgjSpQScHI/G5df/eeWeJqiGUtQF7aaUjmad46r6EaJK0dshsP72uqrLgICmfwK
Rmjp7D+d3Wp11UBb/ZZNkuJXvrKW+UGk/eDBuC3/89ZHa+tkJaoDQXDVzwVl0e92HTtaLSDSyXYF
2tiNvlQAM0Smi7p/bbPHJDKQw424M8JKfunvYSepQnVA7UToKHHKJrunLafsNoT5TW2hHOf6sbmH
o9opd6AnKAeVNZMkUOVw/ZwXfeasdYHRgk3ZtFr7RY1O5sKPsJpALRUDpv/Cij2Ysq0ZvUjBZqDG
9X4HJhrd4oMsABxNTWoXkNeDiZq+KpFUaIOOykwix2nkFYob79KP499qo5tPOMAtNZ2Rh2u11ecV
AGSI20ASecU2cihe39lPQLHycz2C5mY7hqbjAH1Br5Qr7FBWzo0vktoWPT5fIWAkATTmpLleXe2j
bsRHVoiBGvIBXoqWUhtOVb2c4wIR2cddMSwDBs1eVHC/TzGBcBLIRBy+7jONBFKKVh+bkvs0LYcG
oPrg+hFm0dBQzZDblzSIo/Ij6MrCbIT6Y/dLFkbMFuTJZOj/XCUpSCMfdQjhC3STiB5VEPRebqaq
OmcgtnCJpohz0LTkqH+7HSzSvB3i9TafTghxjpc5RugfDxlHa/VVN681tGzwa331QWL92CNx5EbG
pEPpMnKDeDPZuqO2+XAVy6PiS0dD275Eyoqi+pa6938+yifdwCtf/3jfsyysHL1hCDRdzkNnZQEU
7eAYrlsmbwgHFIAoU1YWeVOdDI31DGTslVVPVwCJZ/HKiNgqV6fOwk/ej7rrRtmA3v+UlTPXw9/w
cNmEgwwXuzQWGURvLHMGfnUG+JFfc6VoLAb0OZsyZPquYAPN/KQqLeGACLkFKr40zs/ZlrafRYSB
I+ICD6W0DMYwP6qg/AsmhlV+0BsdrbwkJYk6/c+3wm1khLjhMjRJxoSkTaSo+qDqurayypNVSl0M
MEsUm3YNXDQtKpO12fvWI1THmRamy5NxjmEFGzKte8XYfuVfbFCpln0udSfIlCuAdmzSKFr0i6iv
IWOeF5Gdtm7PIAuL9D/lTlxibpgD+/ZHf/VoVZB3lj7+ITojmOvf/6o2ZfVU/bA0OO52mWSqY4XP
PAG78Gdm7/kcGkJPLhbT59oZedThVhzXocetNihPzRSRf++i3Vq1g1HGR0y6JXu9Bx4X5oiKo0Jf
Xyg2+hyablrIpFK/Af62KtcHlMX9jM9vjLON2H4XKRc9kl038esA8uhsC5cQSMfwD3d93Np9yedV
u2sntlIru+KjndjkUXsT2LxAoaRViBPCk/HgkGjPNd55WOYveDn1Q7PSsq5VOIj7DOMhauk71rDH
Ec8yZlTve/esD2X4K4UKEnl0B/JkYTk2c1FOxAkSfBje8p+IPTvMyBCsDixY4Ch4pQlihq5x9FsS
va6mXqTD5Z8vwtREDQegJv7F34Vj+5DP4+uS/vwNepzN5j8SU0UhvoKCsZhZSiQq36eDIAlNe5qx
miHOK2bOhPhRsO4vB8QSrurm7ku+CO6ySf2NkRi7zmrFprOB/3Lx9hynQDS0FOVyueRj3zoqsdUp
uFq6MkS0ZApYFgmJ8gzJb/jbLM5LZlPAojJrAt46KAWMsJKqocFuWTIoqK8msegVOtD8pF07gjNr
pW1WmPZxXqTXTK4Jg0IK+awSF0gLt8F9BD4R+B8BWRauN1jbUrax+IHr+Z0Gu4SnFuweoT9VjN/F
S04jSo4tZqwubk2iATMkEv8wu4iVc/NwlK0PuGZMOxJFbfzpozK0pV2o5tjWdSEWcJkarei6+l+T
sW9SqHAyNm6tLh0RaZYx488kf23/G/QK3t7zhHOcVQ+eqEd1j76VYuu2inQAPQqRUb1dAMHkN19R
vxSoI/YeDDrcrGVpY2qcOavEZgNZgjSHK0zXW55eKKP5mgfgSLo4xT8Rwxr+4hyl3/HghTMkoXis
RQStCe9TQdVFCn+j7Ppub109mEN5ROyTAsKZPTQMDpvHu24T39/YO8KmNFiM7Eh9Imu+G6JfTQ44
tqTbHMEyyMBW3QfTR1ja8qN85DQutPMYSp1/SRPuusoh9mX7FNYGWOIYAgACUeYBfCCuXMpCqptT
yQfPADLPsNRAJn8y1JxGRj6kk013/fcSt78kIJiDZ4uSUz5tMeVl+c7fMUqMoDK60rd2Dlkd2hd7
Q/xTITm7JEOI5Lo5n0FggQvshvVH2+XVfMRiLGYNnY90kgMD2dOar9cP96FjlZc4Joi3e9buInlG
KVVYlHkyvbx9kSm8c7fscq+Jx7Duy7hDS68gt1iMoyra2xSEXOyGF/UJ4NFT3ynMuB+jPJ0VmNX7
l3cmYc20vi0fn+KXcbkGuSjeIRlBZDHd3LlB3ldbfCh41kxnKRrY5JMgMlv/PqUrlR9GLW/S5Yl8
tfYeabJ+OLE0bYKBjZynrOyX5jVV78AvLLem+yQmmjxU79hD3rLwmbkinTjj+XHpK6oE3OxE18d2
BB7MrzaSDUG8zftM1j9NE2zc7htqpsziNjSqDaddC3XNeNmcRDbvhgs7bdbLKv014fJAbsQrhsBv
kWA0RsBqrNYZe6l8OBIT0dQIU5bFssQT0sN6QX70RXP5Rm83ta5y9lqJ8+r9SgQyZxVbi8Jricsb
T/ODUTHWFxgR27FNZb6Vc0dZKktE2w/jWhS+el4TpBe85UQE01OdkPyBJYB1WpbsmaB7wAERWtv7
u8w7YiksgkodcMkUIUmL8muMQGet1OdFD+2qeM4e1Ev2fQHsQNRNWgXvTgvriOlQGL7rEatS9bjC
RLGWLG2J88y5cToCUdwse5GwHICJEe2hxWLuL3eJkIJefEY/yMjb+kJYwUU3J1ksTyF8ig2QfH4J
msOUbwjGkMTgo5QCFq6z86z/VnIW5DZv2RS9+kloaM8hvYJ6Ld3x1hhtKJgq1bTL4wDGtkG7WTVC
LFuH7nRFNh1ET5+Iu1bYhrdOAa5gqrR5OUraRUgQUD/hPMzpvyAxKI1LyDfLreNRNwCqzAuJcX4k
jVlIYQuSnIq47VR6yVmXO++CpHsvzjQNAT2ylRjtLMywaMiYxV9+IeK/LU6vzy3lMRCMF8f4XWDw
68EDBoQHXlri2VK7Mvq7KRkFojFgKGGe/wXqvnil7sfEOFmciJyu+w+EBpimxP7LtraE+toJKBgR
dsoG0A6PWKPVp3lIPtP/NjSlLKVlRGmgT1mvhJwLM7elb/zD0DGcU4NFxmGas/oKGqDxRYshp6Tp
tIWQHU0ms9DuHxlfc10MgvocSiGoNPFiizHzOlrZwy63WwTmopJihlWfrxRsNzKQGkc9VFBnHGLW
YQULEYX/3ItTnloho04I/L7YiReXtvIijmN0n6SR+Okr48RE2kfSkkraQ0xqwHAptv795WP0AyT4
xc2xGvHd7DnJOGe6XlnZTUr8UzRoyS2R0oz8+rgRuWC/dedBuMQJomBzDnaavdP/wx5vblJ9eAvD
pmXe9+wRP50atFPDZOF4iM8M11StzASCwTZX4mybapfE4WkZOpw4nWg+h7tlCQOxWAwdXDIr6nk+
0VpAQHzqqDxGMiMoTymp/LZe5R7sMTMfRpLI5bFaJ6koj+nk+Yw1NE1atT2AMA2fARyCUNs0Cyhh
qxPlISSaJBYIwqSbmED7tAOOC0BYCGtqqo/s3Fpj+dgdCyR8VsAPPvmm/b9CShA9eUK6zolrMdGt
s3wxv/9Mv190Nx6CCA9+5iaMlXaCqPILuypQM8rXoduWzw6wrMNws92AucrDms15fjNNBFF8KXkH
J45SV9P59jSRvBYL6xgUGkXg5SXSTaTf+cnG4p7nWt82s67dlgMwnU2+JfbPxe3MjuJZ/wgXQKE9
RyF7DOIu/Iq1GfI+iaVwEWM6LeUxA7cMOgsG6msJrbPQdPv67uxWJjxx5S0rPlQABGtgBUFL0Ec4
DEEgq04en2DcLsDaYTT8JnAf6xBIYoa2MpcNQnIWcRUjNS+NcM33S+HIzHBbGLkYxTHxmyHi3I13
BR8jwbCPS8hJ3+FvstsRS2RRcB31LtyO+YnlZLakDr1ECAsiAWbyHJrhjtfM/GNBRVUmGWJoADuO
xA722zwrt3c755bXUiQVj8CM4yYi/Y9VHoiQHsExZYtB96Gyh9sNKaHvTHSSkcq/Lo2ryNsuFnMc
uEnWSVowrWggZVSdz2ZxvNWpoOj8mRS753AZq52dYQHQsRGVgW5PUmfx5FYPXeKSQXV/lYABuEXe
T0NFfCB01G0ZmapdsLcLn/r/4XzWR180qyBPHClChdEHuJHLmxi7q9KJlU62e1K31fDXaVNxG9UU
wUhFMa4TcPCMF8pSSxDsdttFlUfykPjD8lIKpn8LVidc2+7dtpf3XnWyy7nSR2TGPaQiF/5Vg5mh
gsOBZg3x/jFH6iX3/VXBVc6bd0WC9mIsXokESJ8ttacqMw8/XrbGlfKWfs8pe7+ZH1pmVCUcJjlf
ALi/1iWxQgVT+glrNpA8J1U2u58rf/dlCe5dE/ykdMEAwdi8oGDXP6qktDxGN07ll/vwi34plkfe
gc65kumenhLoj8hmcN3Bl5RK/Bss8CTs1A9zS0LtX05+GbReAaU40lBJvqoychEs8wh3eI0y79+c
Gz12bkIfLkNg261tYMwKzVGmEy9buuFn6/GtJgVQAbSnoH0Wwr1IJ6AT88Vd2AS19LX7Utrlav2c
nLNpUZmAqhoMXLufR6bdHTo8oxx/m54ZpVkXbm+kd8dKXEQcv2Sj7Ku4Cz/lgAZunDhzUIm+MSXA
G2FITJo4WyHmtMff5+Sb6bZPmvEUzDxzp+or5vJ+5O2yY6yMlbVdfwNr70JrWxopGaNLsoXMTEFZ
6UIGdeLrzB35ACOpb2xmuVlH1Tt5+RQg93e8AE+gJh/xL02v0PG8/aNgiSO0XQQuxkmlC43kITpd
33hvOTtcGhsNFbZz6rpLCps/Z36OSulTljKDLxMPfz81k0HH4wmprIH5KhQzewISgT99w+xEZE7R
S702JVOGbQTRhGivEHsWnN7pzQppym+jwognPLzbbjODRlsTqGSUFN0g4DIVBfF0gAHsJ+Abz6Z9
BEndEIzjDPeuTvYAwKNrBgtHCMe/FWI21vlL/XggnCC4LXR5sBK7in7T62214fA/cEy3KMd4UMEn
n/ivevIHJAksbDJ75HgVqP4bRwoKpxQ2dEdXfRjQpIepoUVTnMQWLSuSUGYv8FtW010fqxln6mqr
MPq/Y6+/bOnjXnjxf19J8Qq3boiBYdbckWBuCr2aLP9CsLBzJF68ugMi40dNal7hDO/O6x93Z5Az
Z9hcfHDh4bV/Q5QaztZmc25NVheIMNNL4d/ODFehnPvk7aOt4vK1uKEefvf3/oBzT4lxVAiKO/pQ
Bu8PsCsVKTG7vI9sWgus5vtGeLvEAU5TDmMDmBHYf1FQ2YFs6ah0pmZgPoBlhOojsNLsLx9RPVfp
knERxXwsX0EWdIZtWLUUu83iEAxehIUb6XqA13hQEUd2eZEkn4Kd0zeZdtoTs0p7jMbuz9G+1F5d
mBry/lJ/7WUx1rME8WIrxpOJ9hHe3Mr+AWmhzrpugODsSADuj/gXwCTetvswHJt2pkTJ9NtVvfX+
kkm+xrhXRcY2KUvuht/i3Djmx+S3Il3rt8Jmz375oYIS7Z3Ne1J6yjpHUFW5JZSV8PgsKMD+ZpQq
BchZsY3ytB3jRzvhVlGHMTlMBNXrY/EhLAqCL3uQponPG2Zm86ahtdfYRU6/1OcdIeXzKEbu5trx
LLkH/Lfv4eKGYFnMyFBYDxlWy84Yxp45lVlRfbNHyxt7rR+ytkI5i+nKiq7MZKCDi9KO4R8u/ZLr
t0z0QSL7uMjcJahPfgAKG0uj4QGPxxYhN/1Lf8CdWEs1LPGQ38bJA/f3qljQhpPylj6NhvJk/x4Q
JCa0iQsyvQfLhXHSC4runkXn/HSSwNft+kbwxtcTMPogqWaL6VvGYxv1heVJpSiK8EtApDs0iGSP
tKkbpM4XFrje+j7trTwpwoyt+ocIT968b6f9pVb1Cn+kTK03ndbnygP5LKWHNbkhwM2VMOVRt7Ra
O6EKD//F+mCPM2ZaeQPwFX5DNtK6QyvnmUX+SUiG+ADXQwhw6OmeBOB5iuVlhvw6U4rNnHzdxXul
VoWJ82+ObuGiPteOioW1jgoqe7FH03DOOI6gk/e0WLrOm8kw1oVJYLY+6NKBVoywMei02AygX5kj
dIlBnF0HdTqtI6Q3XAH8PWtIQsPJBeCi9q5Wq2YD2TEu8/MWLmseHnXl8jbRrqJJ7vNIHEHbFdwE
kZu1yXfYBi47Rn9PEgYp/Au8BjgNUy1Lcic8Br8tXfPCtoHKr9FZf906GL7J1Wd0jxgUCI+SHt1r
tIDMv4YbJ7K2f6S1d5qJpWgEj2Iqhsod6/OPVKYykmeGxlBX94sVeie9c4RmXQSetMnbVbXhBnlY
k1u9U/GFkkLyqmWiae2i+QJ0N2fi60eNEEgs9hLU7NblaT8Oqhny0LlIugUzb0zxe4ZBTi/QaRkM
BZKq3UDLoMm0Yk3ctT18ZPtHXGP8At8NgZK6P+BODGkwAy0XMvkbUlupAlalI4Dua3TI3hBFCf1x
f7MXkxPcczc/NXIXLMLiGiIgkmeKAiPLsy4NEoLmfUgSOH2vb713TI79g3EHfdioTNuHxV0BMiFT
sb7UGWVTQAm7C+h1GJRmIxOEXPMYQ6Zt6uVgVXTzCuyLx/WzcSDttVYde+3ZGuX+6jKeb2nvZArV
o/99J1baxmiTV2BH3pkmnM+HdOMO9DRVSvsiRgCYYKKZ6jCH5z05AerGUMh+ltgWlze+arhtsD5O
5LsPbvgxya63XZW16BfDST0WYtPdNY0geZDK+Qt7Q0CTTuaR3xJYdDbV3rolv+dRjRP3fQWN47v1
DSlfB/oisaBG6OCcmIx4W4HtkVNd6EMbZCxtuqUvH2tfdnBv9HTopmiKVJnien8Je0bjqHm1L/sq
bRjiJiDiRH6zzXpU57uLBmIUPS6SSFJ0cmbNdqTAjFkwEdR8Jn1yQ9kvJeUUgQTuvZAMWHw4zQAG
XOvIaMXJHzHJwLzk6JW5TOkpJ92GmlPiM4nzdpYEjphSHjwVSQcyZ4Q925QSl3S46LynrlrhMMbl
UfJqO4wbNw5Ejmo0jFHtMe5j0B2fKFJSigCqf+eVkoDN47eHP+ZPwGKp6rg3hegdg1PpD7e8CaLf
/xLVsdTUAiHEkKA5elHb7Mae93tbBdKon7lw94KPjNcjQGf6SDHxlYRc3KUE+FIXea6ESp2NgwOf
NMEzKgrdDw+vP1lilwfIwj9jP1tbWPVKa5bEdYx8Mf6S4LZtLfI0RA8lyTfQEBgHymN/OpsLFGFZ
pccTG8UZOwcIaC9yQU5M0fMqavyx9mLzgldKmDJ3XXFUPVxH7GONpw8J60LOOyDQ/ow8aGZBWATw
3oTqd54VnGR/rcRaiSF8qEnHCZ82bIpxZVy3cDJLqCcJDt+OMe3tJOheiERSVP2+k2jo6lkdXz7k
Sr32Eg3djcZueKOo2ySDQkprhFr1VKBRtfJPndINrl6+0JFu1PfjeO9E2/MoYsaoeHi2rDbCk0Sl
RwCXDEXfnUd05cdRFnrlTlQmrEs+wWtu/sLj3kSo0WOHmvMgKCJDBT0HbX6Vq74YTJ3M82NnwPuD
uVv9Uzy/o0VHHqguk3L58xnoMkXkMqGreTJPCrLMMZRjcQYOfS3eg581ntu2c/OuvA99cNNYSJFO
P6rmpqtjAC4CXy5zS8DAA1P+waLj07k7DDK7GlqIwlwUV7kucabyoUHV8vc3I+1Br8WY22xbCTSY
lnr2B7hzZZ75J8IkhV85f2oBnn00RK2rF2VhFnSbGJzutPfguRGjFFszGRHyK659FdHjvrLHTdGl
/m09Q82n5edfZe5c0k3NQoDgWqDI22D/MHqQcTkXtrsTOIQK9oh2+8f/hBlEf9VkuWQGu9dh53id
rzO4d1fAfY636NXsnBQVadiRhD6A3cRR3BRdd5E4ZiTo0aHiZ9/r++m+kg8xweznPPh5NM75REgO
rgRrD2FmqvjDY4zQiOBKLRYEehvBqYXcThHAaHUefqW+lQGA0PVTrhZLmCz+OOe0QolkAqZzS1ix
j89julpjrdqZagGOhbHYFEVRKDK7OjyppF5gdnFNDMuFbVBZPVYt+Y4IEL2GYcKyLfuamKqpneWZ
/v3UF6im6kHe7/iUR12sQ3wClOtqKaTmSWeBBXolhvr1rgbV++BAx4jchD7YZdpI/UgjX60BD8RK
MWPoQvxmrA+F1SFqQBABN9f3n63kbY2kvRbawVuiB1Tyh8rD/bkCNFWZTmaAxGMfVaZEcTMFP/Fn
AznfX4Pp3513Kinc6EjnAsd8mr776WhVNSSrqdIJfcvwhMeUzhPQ4pT81sI0M0IbyIh5xeQKBV8R
a8c9z8IQFEh5WJbLeEIQDwkle97tYV0AG1Vv5P0Gg6NLSMy/aHYdb0MOQwIhsoBfUyKG07HJPeji
mhS/IOGSPnw7r0RBsD66mUGCSF1+N6ItSH0hO4J7qkzaQE5mrqfi+E3x9wmKy8az2lhhc9dVpKm6
V7BB6cE4Ozt/1TA8JLyo1wAQ928kzchvSZ3coKCPhm7wNqSt58tAqgy352bn+X8Q10CTFok0Vwda
qYcUdjT7iy7LhT7ZXmuz8dTvUpSNWYKgJfhs1lbuqjJE6pfGNxSUr5Xs6qtxtL4/cZvAWqUu7lyL
GfZJanMyaKsNrkBzQ9PuBpEb7z/NByhhBH5nom1iyRTdBHtLsLAw1+MVmbovynTBHogidIIpG7fM
a/A/GIkR5pS+e/knwr/5RD+FMYCL4u8jElA5NeXnuEKJJLxLrPXIT8ESBeVOL32bYQm4BUKXVECH
WUp1XcskSX6syiiV2imfOKo8vDt1G4vj/Rny8sIGXoZM+GOaxVerijGn9Fuhog8nvljQR9lF2Iod
tZ7y5YQxxqoophEplXzfWwUz0an9Vevqe9Kn5dYNhfS4nbJuxQnccdTfQhC/rtLHp0E6Wiw+GDEi
6uhOTgbgmPskJHpwkrznVgkm60QC5f7nlkH7bzIl7Qi5xS68VV5mOfH3ZJQTHWxFEqVHY06PT0Oy
nBJofNtj22I5578N9QQNBT3GjfoYrObrqHModtasrYzkd35uWwtRwF/nn+DwR7WFqZa+PqE4JAoj
Bh89VxOqetqWblSipXOWyXFGxgSt/DdrgoMmoMPq2VnKR/Ohh/PGAq+rCH+yIR7swzXaKndpdcQg
U4w9oO6RnOTtrMVeEfN3GbgefZirQV5XL1jiXS290N1Y8WCJiXfW0TApK06AEPXi7OsBrRkwN7Rf
vIPbAZ7BY5leLOB+TqcZOvP0c6n4zOHRi1JPFNuljbYwS9e90Pd8k9UWyDOjM78+eOhl0RVGjiyr
APXayrIn0Jo954vInO5NJzK7jbl5njGVnyyLu9UCfiA0lI4pRvTI4c6nNmaqQjNkM1vd3eZVverv
rS3k0y42t/ZdOr4RMNkRQj5nf5r2NsSROISbh5iL6gjExIqosOmDiytVu89b1BrJ5QH/nObG2g48
ZBIZ6m0W+Y9ZdiG0cme2fhnDt629hjr1VNSKZS20a3NXw5jxlkbkjqXgRDedtN0P6NztoKb5zDyV
2L0r2an/Enh5K0zDeOVABt8+WOF8vG8vXJhiIuqY9Qm6GuhJcnWqChqBNZq32swISo0j4+jV4zCT
yhhW4hk9uX2f+P0xtVSHWYJ4qZ9saaT1RkzJzpJm+idDx3MgpnER1NbA+m0ku+L9/VY7M59HV/mb
hQvlyKwOrdyRdN3QU3OUAV/x+jvm1uaXOOU6hl+ykMTVH+ut/M1BxsHZyjxPpbnzzSEqCxPOp9Ut
Hholwck8Lx4j/fzHQ5G/T8lwAtyM5ygNRGr/L4z0qZHCR580M1/8WPKAogIGFJSN/GsUAEhjG+eU
+ZSdVHZQ2j22wkTtAf4WOQ3s30XQ/CkLYtfOu9c7LANxeHgD+mc4dR47E3CeuSp+ya4O+WZX+l6o
+xxH6vSppAkrenvnbM/FuP+SetrRtdp/Qbea5ZyhodR4khnWdyELzzAT2ciIpQx1RXj+SjkKgSwE
gtW3m+c2p4nn+c1lSdJTimMLDueocRe6F/bwkii4OODdiexWjmd8DNTXmgw9lp6vsw/VYqwhv2Vc
W8W28JC4MUFhlNzPgs150Op8eFYC0Vs9lp7BMQ24xrRQb9bVzHfyGZT8EDiazebX
`pragma protect end_protected
