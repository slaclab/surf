-------------------------------------------------------------------------------
-- Title      : PGPv4: https://confluence.slac.stanford.edu/x/1dzgEQ
-------------------------------------------------------------------------------
-- Company    : SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------
-- Description: PGPv4 GTY Ultrascale+ Core Module
-------------------------------------------------------------------------------
-- This file is part of 'SLAC Firmware Standard Library'.
-- It is subject to the license terms in the LICENSE.txt file found in the
-- top-level directory of this distribution and at:
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html.
-- No part of 'SLAC Firmware Standard Library', including this file,
-- may be copied, modified, propagated, or distributed except according to
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library surf;
use surf.StdRtlPkg.all;
use surf.AxiStreamPkg.all;
use surf.AxiLitePkg.all;
use surf.Pgp4Pkg.all;

library unisim;
use unisim.vcomponents.all;

entity Pgp4GtyUs is
   generic (
      TPD_G                       : time                  := 1 ns;
      RATE_G                      : string                := "10.3125Gbps";  -- or "6.25Gbps" or "3.125Gbps"
      SYNTH_MODE_G                : string                := "inferred";
      ----------------------------------------------------------------------------------------------
      -- PGP Settings
      ----------------------------------------------------------------------------------------------
      PGP_FEC_ENABLE_G            : boolean               := false;
      PGP_RX_ENABLE_G             : boolean               := true;
      RX_ALIGN_SLIP_WAIT_G        : integer               := 32;
      PGP_TX_ENABLE_G             : boolean               := true;
      NUM_VC_G                    : integer range 1 to 16 := 4;
      TX_CELL_WORDS_MAX_G         : integer               := PGP4_DEFAULT_TX_CELL_WORDS_MAX_C;  -- Number of 64-bit words per cell
      TX_MUX_MODE_G               : string                := "INDEXED";  -- Or "ROUTED"
      TX_MUX_TDEST_ROUTES_G       : Slv8Array             := (0      => "--------");  -- Only used in ROUTED mode
      TX_MUX_TDEST_LOW_G          : integer range 0 to 7  := 0;
      TX_MUX_ILEAVE_EN_G          : boolean               := true;
      TX_MUX_ILEAVE_ON_NOTVALID_G : boolean               := true;
      EN_DRP_G                    : boolean               := false;
      EN_PGP_MON_G                : boolean               := false;
      WRITE_EN_G                  : boolean               := true;  -- Set to false when on remote end of a link
      TX_POLARITY_G               : sl                    := '0';
      RX_POLARITY_G               : sl                    := '0';
      STATUS_CNT_WIDTH_G          : natural range 1 to 32 := 16;
      ERROR_CNT_WIDTH_G           : natural range 1 to 32 := 8;
      AXIL_BASE_ADDR_G            : slv(31 downto 0)      := (others => '0');
      AXIL_CLK_FREQ_G             : real                  := 125.0E+6);
   port (
      -- Stable Clock and Reset
      stableClk    : in  sl;            -- GT needs a stable clock to "boot up"
      stableRst    : in  sl;
      -- QPLL Interface
      qpllLock     : in  slv(1 downto 0);
      qpllclk      : in  slv(1 downto 0);
      qpllrefclk   : in  slv(1 downto 0);
      qpllRst      : out slv(1 downto 0);
      -- Gt Serial IO
      pgpGtTxP     : out sl;
      pgpGtTxN     : out sl;
      pgpGtRxP     : in  sl;
      pgpGtRxN     : in  sl;
      -- Clocking
      pgpClk       : out sl;
      pgpClkRst    : out sl;
      -- Non VC Rx Signals
      pgpRxIn      : in  Pgp4RxInType;
      pgpRxOut     : out Pgp4RxOutType;
      -- Non VC Tx Signals
      pgpTxIn      : in  Pgp4TxInType;
      pgpTxOut     : out Pgp4TxOutType;
      -- Frame Transmit Interface
      pgpTxMasters : in  AxiStreamMasterArray(NUM_VC_G-1 downto 0);
      pgpTxSlaves  : out AxiStreamSlaveArray(NUM_VC_G-1 downto 0);
      -- Frame Receive Interface
      pgpRxMasters : out AxiStreamMasterArray(NUM_VC_G-1 downto 0);
      pgpRxCtrl    : in  AxiStreamCtrlArray(NUM_VC_G-1 downto 0);

      -- AXI-Lite Register Interface (axilClk domain)
      axilClk         : in  sl                     := '0';
      axilRst         : in  sl                     := '0';
      axilReadMaster  : in  AxiLiteReadMasterType  := AXI_LITE_READ_MASTER_INIT_C;
      axilReadSlave   : out AxiLiteReadSlaveType   := AXI_LITE_READ_SLAVE_EMPTY_DECERR_C;
      axilWriteMaster : in  AxiLiteWriteMasterType := AXI_LITE_WRITE_MASTER_INIT_C;
      axilWriteSlave  : out AxiLiteWriteSlaveType  := AXI_LITE_WRITE_SLAVE_EMPTY_DECERR_C);
end Pgp4GtyUs;

architecture rtl of Pgp4GtyUs is

   -- clocks
   signal pgpRxClkInt : sl;
   signal pgpRxRstInt : sl;
   signal pgpTxClkInt : sl;
   signal pgpTxRstInt : sl;

   -- PgpRx Signals
--   signal gtRxUserReset : sl;
   signal phyRxClk         : sl;
   signal phyRxRst         : sl;
   signal phyRxInit        : sl;
   signal phyRxActive      : sl;
   signal phyRxValid       : sl;
   signal phyRxHeader      : slv(1 downto 0);
   signal phyRxData        : slv(63 downto 0);
   signal phyRxStartSeq    : sl;
   signal phyRxSlip        : sl;
   signal phyRxFecByp      : sl;
   signal phyRxFecInjErr   : sl;
   signal phyRxFecLock     : sl;
   signal phyRxFecCorInc   : sl;
   signal phyRxFecUnCorInc : sl;

   -- PgpTx Signals
--   signal gtTxUserReset : sl;
   signal phyTxActive    : sl;
   signal phyTxStart     : sl;
   signal phyTxData      : slv(63 downto 0);
   signal phyTxHeader    : slv(1 downto 0);
   signal phyTxFecByp    : sl;

   constant NUM_AXIL_MASTERS_C : integer := 2;
   constant PGP_AXIL_INDEX_C   : integer := 0;
   constant DRP_AXIL_INDEX_C   : integer := 1;

   constant XBAR_CONFIG_C : AxiLiteCrossbarMasterConfigArray(NUM_AXIL_MASTERS_C-1 downto 0) := (
      PGP_AXIL_INDEX_C => (
         baseAddr      => AXIL_BASE_ADDR_G,
         addrBits      => 12,
         connectivity  => X"FFFF"),
      DRP_AXIL_INDEX_C => (
         baseAddr      => AXIL_BASE_ADDR_G + X"1000",
         addrBits      => 12,
         connectivity  => X"FFFF"));

   signal axilReadMasters  : AxiLiteReadMasterArray(NUM_AXIL_MASTERS_C-1 downto 0)  := (others => AXI_LITE_READ_MASTER_INIT_C);
   signal axilReadSlaves   : AxiLiteReadSlaveArray(NUM_AXIL_MASTERS_C-1 downto 0)   := (others => AXI_LITE_READ_SLAVE_EMPTY_DECERR_C);
   signal axilWriteMasters : AxiLiteWriteMasterArray(NUM_AXIL_MASTERS_C-1 downto 0) := (others => AXI_LITE_WRITE_MASTER_INIT_C);
   signal axilWriteSlaves  : AxiLiteWriteSlaveArray(NUM_AXIL_MASTERS_C-1 downto 0)  := (others => AXI_LITE_WRITE_SLAVE_EMPTY_DECERR_C);

   signal loopback     : slv(2 downto 0);
   signal txDiffCtrl   : slv(4 downto 0);
   signal txPreCursor  : slv(4 downto 0);
   signal txPostCursor : slv(4 downto 0);

   signal txPolarity : sl;
   signal rxPolarity : sl;

begin

   pgpClk    <= pgpTxClkInt;
   pgpClkRst <= pgpTxRstInt;

   --gtRxUserReset <= phyRxInit or pgpRxIn.resetRx;
   --gtTxUserReset <= pgpTxRst;

   GEN_XBAR : if (EN_DRP_G and EN_PGP_MON_G) generate
      U_XBAR : entity surf.AxiLiteCrossbar
         generic map (
            TPD_G              => TPD_G,
            NUM_SLAVE_SLOTS_G  => 1,
            NUM_MASTER_SLOTS_G => NUM_AXIL_MASTERS_C,
            MASTERS_CONFIG_G   => XBAR_CONFIG_C)
         port map (
            axiClk              => axilClk,
            axiClkRst           => axilRst,
            sAxiWriteMasters(0) => axilWriteMaster,
            sAxiWriteSlaves(0)  => axilWriteSlave,
            sAxiReadMasters(0)  => axilReadMaster,
            sAxiReadSlaves(0)   => axilReadSlave,
            mAxiWriteMasters    => axilWriteMasters,
            mAxiWriteSlaves     => axilWriteSlaves,
            mAxiReadMasters     => axilReadMasters,
            mAxiReadSlaves      => axilReadSlaves);
   end generate GEN_XBAR;

   -- If DRP or PGP_MON not enabled, no crossbar needed
   -- If neither enabled, default values will auto-terminate the bus
   GEN_DRP_ONLY : if (EN_DRP_G and not EN_PGP_MON_G) generate
      axilWriteSlave                     <= axilWriteSlaves(DRP_AXIL_INDEX_C);
      axilWriteMasters(DRP_AXIL_INDEX_C) <= axilWriteMaster;
      axilReadSlave                      <= axilReadSlaves(DRP_AXIL_INDEX_C);
      axilReadMasters(DRP_AXIL_INDEX_C)  <= axilReadMaster;
   end generate GEN_DRP_ONLY;

   GEN_PGP_MON_ONLY : if (EN_PGP_MON_G and not EN_DRP_G) generate
      axilWriteSlave                     <= axilWriteSlaves(PGP_AXIL_INDEX_C);
      axilWriteMasters(PGP_AXIL_INDEX_C) <= axilWriteMaster;
      axilReadSlave                      <= axilReadSlaves(PGP_AXIL_INDEX_C);
      axilReadMasters(PGP_AXIL_INDEX_C)  <= axilReadMaster;
   end generate GEN_PGP_MON_ONLY;

   U_Pgp4Core_1 : entity surf.Pgp4Core
      generic map (
         TPD_G                       => TPD_G,
         NUM_VC_G                    => NUM_VC_G,
         PGP_FEC_ENABLE_G            => PGP_FEC_ENABLE_G,
         PGP_RX_ENABLE_G             => PGP_RX_ENABLE_G,
         RX_ALIGN_SLIP_WAIT_G        => RX_ALIGN_SLIP_WAIT_G,
         PGP_TX_ENABLE_G             => PGP_TX_ENABLE_G,
         TX_CELL_WORDS_MAX_G         => TX_CELL_WORDS_MAX_G,
         TX_MUX_MODE_G               => TX_MUX_MODE_G,
         TX_MUX_TDEST_ROUTES_G       => TX_MUX_TDEST_ROUTES_G,
         TX_MUX_TDEST_LOW_G          => TX_MUX_TDEST_LOW_G,
         TX_MUX_ILEAVE_EN_G          => TX_MUX_ILEAVE_EN_G,
         TX_MUX_ILEAVE_ON_NOTVALID_G => TX_MUX_ILEAVE_ON_NOTVALID_G,
         EN_PGP_MON_G                => EN_PGP_MON_G,
         WRITE_EN_G                  => WRITE_EN_G,
         STATUS_CNT_WIDTH_G          => STATUS_CNT_WIDTH_G,
         ERROR_CNT_WIDTH_G           => ERROR_CNT_WIDTH_G,
         TX_POLARITY_G               => TX_POLARITY_G,
         RX_POLARITY_G               => RX_POLARITY_G,
         RX_CRC_PIPELINE_G           => ite((RATE_G = "17.1875Gbps") or (RATE_G = "18.75Gbps") or (RATE_G = "20.625Gbps") or (RATE_G = "25.625Gbps"), 1, 0),
         AXIL_CLK_FREQ_G             => AXIL_CLK_FREQ_G)
      port map (
         -- Tx User interface
         pgpTxClk         => pgpTxClkInt,                         -- [in]
         pgpTxRst         => pgpTxRstInt,                         -- [in]
         pgpTxIn          => pgpTxIn,                             -- [in]
         pgpTxOut         => pgpTxOut,                            -- [out]
         pgpTxMasters     => pgpTxMasters,                        -- [in]
         pgpTxSlaves      => pgpTxSlaves,                         -- [out]
         -- Tx PHY interface
         phyTxActive      => phyTxActive,                         -- [in]
         phyTxReady       => '1',                                 -- [in]
         phyTxStart       => phyTxStart,                          -- [out]
         phyTxData        => phyTxData,                           -- [out]
         phyTxHeader      => phyTxHeader,                         -- [out]
         phyTxFecByp      => phyTxFecByp,                         -- [out]
         -- Rx User interface
         pgpRxClk         => pgpTxClkInt,                         -- [in]
         pgpRxRst         => pgpTxRstInt,                         -- [in]
         pgpRxIn          => pgpRxIn,                             -- [in]
         pgpRxOut         => pgpRxOut,                            -- [out]
         pgpRxMasters     => pgpRxMasters,                        -- [out]
         pgpRxCtrl        => pgpRxCtrl,                           -- [in]
         -- Rx PHY interface
         phyRxClk         => phyRxClk,                            -- [in]
         phyRxRst         => phyRxRst,                            -- [in]
         phyRxInit        => phyRxInit,                           -- [out]
         phyRxActive      => phyRxActive,                         -- [in]
         phyRxValid       => phyRxValid,                          -- [in]
         phyRxHeader      => phyRxHeader,                         -- [in]
         phyRxData        => phyRxData,                           -- [in]
         phyRxStartSeq    => phyRxStartSeq,                       -- [in]
         phyRxSlip        => phyRxSlip,                           -- [out]
         phyRxFecByp      => phyRxFecByp,                         -- [out]
         phyRxFecInjErr   => phyRxFecInjErr,                      -- [out]
         phyRxFecLock     => phyRxFecLock,                        -- [in]
         phyRxFecCorInc   => phyRxFecCorInc,                      -- [in]
         phyRxFecUnCorInc => phyRxFecUnCorInc,                    -- [in]
         -- Debug Interface
         loopback         => loopback,                            -- [out]
         txDiffCtrl       => txDiffCtrl,                          -- [out]
         txPreCursor      => txPreCursor,                         -- [out]
         txPostCursor     => txPostCursor,                        -- [out]
         txPolarity       => txPolarity,                          -- [out]
         rxPolarity       => rxPolarity,                          -- [out]
         -- AXI-Lite Register Interface (axilClk domain)
         axilClk          => axilClk,                             -- [in]
         axilRst          => axilRst,                             -- [in]
         axilReadMaster   => axilReadMasters(PGP_AXIL_INDEX_C),   -- [in]
         axilReadSlave    => axilReadSlaves(PGP_AXIL_INDEX_C),    -- [out]
         axilWriteMaster  => axilWriteMasters(PGP_AXIL_INDEX_C),  -- [in]
         axilWriteSlave   => axilWriteSlaves(PGP_AXIL_INDEX_C));  -- [out]

   --------------------------
   -- Wrapper for GTH IP core
   --------------------------
   U_Pgp3GtyUsIpWrapper_1 : entity surf.Pgp3GtyUsIpWrapper  -- Same IP core for both PGPv3 and PGPv4
      generic map (
         TPD_G    => TPD_G,
         RATE_G   => RATE_G,
         EN_FEC_G => PGP_FEC_ENABLE_G,
         EN_DRP_G => EN_DRP_G)
      port map (
         stableClk       => stableClk,  -- [in]
         stableRst       => stableRst,  -- [in]
         qpllLock        => qpllLock,   -- [in]
         qpllclk         => qpllclk,    -- [in]
         qpllrefclk      => qpllrefclk,                     -- [in]
         qpllRst         => qpllRst,    -- [out]
         gtRxP           => pgpGtRxP,   -- [in]
         gtRxN           => pgpGtRxN,   -- [in]
         gtTxP           => pgpGtTxP,   -- [out]
         gtTxN           => pgpGtTxN,   -- [out]
         rxReset         => phyRxInit,  -- [in]
         rxUsrClkActive  => open,       -- [out]
         rxResetDone     => phyRxActive,                    -- [out]
         rxUsrClk        => open,       -- [out]
         rxUsrClk2       => phyRxClk,   -- [out]
         rxUsrClkRst     => phyRxRst,   -- [out]
         rxData          => phyRxData,  -- [out]
         rxDataValid     => phyRxValid,                     -- [out]
         rxHeader        => phyRxHeader,                    -- [out]
         rxHeaderValid   => open,       -- [out]
         rxStartOfSeq    => phyRxStartSeq,                  -- [out]
         rxGearboxSlip   => phyRxSlip,  -- [in]
         rxBypassFec     => phyRxFecByp,                    -- [in]
         rxFecInjErr     => phyRxFecInjErr,                 -- [in]
         rxFecLock       => phyRxFecLock,                   -- [out]
         rxFecCorInc     => phyRxFecCorInc,                 -- [out]
         rxFecUnCorInc   => phyRxFecUnCorInc,               -- [out]
         rxOutClk        => open,       -- [out]
         rxPolarity      => rxPolarity,                     -- [in]
         txReset         => '0',        -- [in]
         txUsrClkActive  => open,       -- [out]
         txResetDone     => phyTxActive,                    -- [out]
         txUsrClk        => open,       -- [out]
         txUsrClk2       => pgpTxClkInt,                    -- [out]
         txUsrClkRst     => pgpTxRstInt,                    -- [out]
         txData          => phyTxData,  -- [in]
         txHeader        => phyTxHeader,                    -- [in]
         txBypassFec     => phyTxFecByp,                    -- [in]
         txOutClk        => open,       -- [out]
         txPolarity      => txPolarity,                     -- [in]
         loopback        => loopback,   -- [in]
         txDiffCtrl      => txDiffCtrl,                     -- [in]
         txPreCursor     => txPreCursor,                    -- [in]
         txPostCursor    => txPostCursor,                   -- [in]
         axilClk         => axilClk,    -- [in]
         axilRst         => axilRst,    -- [in]
         axilReadMaster  => axilReadMasters(DRP_AXIL_INDEX_C),   -- [in]
         axilReadSlave   => axilReadSlaves(DRP_AXIL_INDEX_C),    -- [out]
         axilWriteMaster => axilWriteMasters(DRP_AXIL_INDEX_C),  -- [in]
         axilWriteSlave  => axilWriteSlaves(DRP_AXIL_INDEX_C));  -- [out]

end rtl;
