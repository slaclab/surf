`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NkVjC+gdv0NPzuql9i8aCe24LW6WOU45yteZa46ADxveOShOhPPTvVxaTiO3hiKizgXWco1/GhmV
AgW/B8D07Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SAuVh2vSQxNJDP9drsSSnGrzI4YKdIcU3EpW0BsXo4dpylBAl8hyD8CLNY8ncFAWHs8+B/RjSpq5
N+4TlV9xttnhn46cHiiRycmLrOfuIC0en8/W7lKKpw3kiJCVCFOc0pUkrxY08Ko0F7yIrA5WLQQH
Slx2IylFDjIutK5RLto=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Vjmt7AkPM77hECJv0z5E1VDl/CLchylFRiYYY83jAbZi5fWSvK+9ywWDUu/ml7pMKcZHuNJ3HHd2
MawxCfueQyIWVC68ujhxpsqf+WEuaPN6wnJMjJAYw773MPjNqDj/mRCil0ifZ/4/d8Xtm1FRgF9+
qKi1A5QqKdGH7kaSzXk1H6IjA+gvJzQqKXumTIYHUla+Hfg08HUJ7pOjLwhsrnHs1mBs9FisgPlT
Aoc4AiPSVZuRvHzAFQvREVujwCjChw4xj5jw5W/dwYMDm/YYG7XTdKdouAMa2bw417Ymt6WK502f
WcMNiGjFqgM+jS4WGyX+KyJCrhyY3+yJFFOElQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dXfEjm3iPxQ/3WBv7Azr6xDxyHgVn6ORnDFuQKvDOEiiZrUkmKT4He1Eo4w8+NLvjdr4QiQZTUnJ
nKhfE7Roi/NsCnn8a+7yeYis/Upp8MZIIiRn/TEeStzxTfaO9WA6169Lz8gb+JJCwzuV2Vfoz6q6
VhQhmkk7FLOGYCBgZRo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CMCvjza2maFliO1h0UdoKFj5u/h0nrkpvf06XFCMmELI9oFLFYPps4+/fQJvOc3nNwDLHmLlh9PE
bfzzguMxR8886WL+U4VOZyvRQ+fZCpdKTqZhbnd82/7O86r+e93/Ou10Ezge6Udhp3ItAh38cOqq
R4Fbr5YLPuB9GEIgpeH21attXEF1F2c9RO6ielvrFdelndkleZ5pgT7aAoV/Myj2nNR09dE2tJCR
JYHsXMBDldR5STjRAVs0GamnRMAIOD4xUSwgJnzHuEZOeoWHAzQ7oBufeIMxXd7hDFGLbWzR8qZT
jt3m/UJBYjxVUJJZQmeLGYw9bAF6+jwiWzQEuw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Vj37nw/1rJQKkjze5fa+SU33y85qg4LAMf3tMlcwNwj6r0cz6hELjaVy9v1102AbIPFCKjtfhD8y
afnroOOAjbbJbAFOlShHk7iZrxFoDFMPtusQTbawI55y7inw3RPJrusXuPdyFtx0kafA2sFQSogK
g4+XsdO4WVS9hSv+oz2wLoN+OF+HpqvikkEpHeopQf+o51WnsWd2J1lCN8AJeZlWqIYtwb66xost
ckWwCThltWhN30RfC9JC9wQtLISBQkrNOsthHDrgiOilWcv2EE1VLlRFRoqJfdWH0jgTg5yZWPJy
f04lvPGYtkTkngOkTLzPlOBUVxN1OvcFB3fYwg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 598944)
`protect data_block
fBG+3d+r+y6qTIgpZGJwGZBlF/CMbzgKx3rmHFgOz6YIxtRIpW6yD0s28XihJzw1ibgEsk5NDFXo
sORLqIEfvn9qs9G3PO3Igjx3GH5BeBh8O4B2Fyy47gSvRoRoyJPrskk+oJuPB9t4ELd7b+8n/2Su
wLeiggjqAGzY9PGj2VLF+5awrNm7zJIbxVH+hF7g031uLzynasK40WHA0mzAI2oJ7EaCKuBGhSZQ
SRacc8VsZ+kaQ9hdcftAolisDIg7KixqcVoEMWoyfzk20D64Krv6+xzKc1dk28OrLtAi32e6r7+F
xgOnvPHaIwe5JrInwKw1YRgwWgZsuAY3OtxFrN5O7Hua4DkaGsjTPhiJMfb01J4sPlHbM4A8FpVL
bvX6v1v/ERHF8hucYu6LZ7piQt2C2I038jl4nCGUx5E4JmBFAuTYrS8gA/C/qVgwRve2/+lse7Ek
1ONFmzDseI5zIQXF7KHIjSaLSbHvSd1cYriqJExM+nIH2zaH7bWw+oNK7zHhP/IQmWN47QF7JDiD
BN6f2kqNv1MpDEh2D5GH54HIPjETX5mbm9xID6JRrjEda3m6EcSev/F85caKUtucB21/P9hTm4Wo
fjiz4wUrfVd+dDDZi9nTVTVw3KeTUifh3YPOy38cN9UJorcEDLc2mCd3JHeYqxKIRU7ugfej5Mpq
Cv1UbCr9/t0+hJPYLBgLdfZBvFRpAhY3anW34NkfvDFBg0fPxQdQkHgttrR9bRLV6jHNJGn/FwsL
skt3UZckUnAlsJl+1P0XjbAfc3L2nLafmm+V5kp2PVNv2kodGHLCZXdZlPrPnhIjNkCn/YOgYzcj
O1jK8U/B1fLHHpSxDvCE80GDbErq8Z073rXfY0nwczx4zBezMdDQzGh8UBTgDA4DPAtliPptKtGg
VTEM9MnNyg8Wxr7T1vp+DQkYeih+95C90joY9Nbab9DgN6Y91Nyz3ogMAUDGgyyYXUER9yhrFz9Z
LCtmrWrng19kPrav+obCs5HyaOIrpdOs2bEHyksdTwu1l8iv3JeqLMkRvMasGIosSfiJe1X02uCw
mnULvTuFKLGUDiuF7Fbd8ZsArh99RKgnQNaQt1s2HtRvmQacZ4c1rcg4iZjzgoNTc4S/8mXY7aNz
3Wmnfeev+2dNcYQuNpGs3NK2Ssjfa53saJvAokdGP5OPho6PtsR2LLOXYdh656HvLZow17ODaxZw
5NKc4xX/xKYN3GzC+92Vyd4ToIjgK3qoM7jT76T0pS6orZCEDa3oZTseMrxuyrlfFzPThBJb+BjQ
yM+rg2mrYks9m8D4pbropmoLU1JX8e76C1z4Iu5pOZEw936IsAKY1giwkeTwnhPJFdBNQUreppKs
VYGydHfE+N552WkerAR31ZBVg+lzTdxcsI/OMQE+ePS275JNkzogjDHu9DNhDBMhoERBedWiPetn
4k73QbwvNC53gvWSRFcYyE8chY0KN2gEm5uXlh31nA9Cd2Ck6QKjBqCMSU//t2q7Z86fGQxfUprV
EJ1rZk2Qq44App2LGvNh4kNkMcPcqW9/BeNc+QnTHdYRwdJNd/WxbJn6qycnAxABY3dRtvqUKKqi
1fKuaTxRsp0oimApD0Cc+Ot3kjjYbGJITpP/ru29C1qqHX0Ip1njWUSXtnSde6rCd3LQj4EBdjzC
pJ0ibt623BVMCAn/OWD1B0C2yCJwrHy/7dnjw6A4ZDaf8zAnayDitHEjQlpDczGKxpHVE9s4zEer
MWC6C8YBJbsLLXPuSkfjk2eG/ZNhy5VhkkJJT4zSnpxpac7phUck/8z8Bxe8jKbAJdCelyK4CzRs
dGY0eWlBEw96l+yV9FtKmgFXi2/CQE3+kL41uQjH00PNf5SKC24F64+hzUZ2YKtjl8LbAcYBzWIR
uvdiLQL67WPwuxlX/GLpprMbBe4bV5MqW+bP/zI+cd0NYJVcb2Yo004FGIBL1IzEIY+63qfhQ413
gq11M6ll2IYSLqv/nZbQTIH8rdMDtEOR/WcIpin8BkbZwWV9Oo/9Ay61YwUERBjmKc5HWDhKS9F6
KWeBZiC8/oyUKvb9J/H3JY6Hwq+7XomcFMsjVInP/pORKRVV+nV0Sta3RE4p8oQmcYbIe9Wf2xCm
lokJtdxMNYFAwwhdvAIagagpN1a6rF8IEZ42JxC6/DMDTC6Kqlm6UaaI2wUGr3N/m43JA2RZ6Iol
JZLm6g3r8DtBRiRRJihPHZ0JVr93Ujh6GiYsRdfogNusWOHc9zh3eauNZhwdXh3JLPCojgJ/Ei1d
Qof7xBwCXhBjwyteK9jW8De86VGCGtf9yEuqdgkEg+VScmyC1NLzG3OKUWpPao2cjYiuTEqABudJ
kKnIBw5+01kd/O1dWcfkLJsHCzc4/JOUiHNzn3Tfe5czjhuNphsuZOaOKmK/n0LA9c2gROoHvka1
sOKHjVLAxdnMAVztcM715kyjII/4wKqSMB7YlGN5PfVMiFIkUQgufkKA/x8p+qS8op9dvwwU5WBT
8iFt0gv5e1VzEkju9JvSQ4PG7uQgMSNQF+oKOl1c6Rznyktc1j/N8BCdNDo6pT4BA9/UH/xcrIwc
h9n72K9jR2n27RzT8wmpGOhoTtAR9/iHL6G2wo4KG0oU27sty9ezcNT3idD5OjSUOmOdQHv7ZxUI
6ZdiDQGvg8NDJ+f9Zno4V7/+yjOPTpebWVMBTppJzQragbn+061iZs7IJ14SSJivTnYmSgGecriG
3OfgQhr/isFkts7kidCg/esReu7z1J9B9s9uW//l2ylMMTVBmDNsZ5CAQR9UsgOtwEBcmp/SQPpa
EvblDsHNe2eHDMEkt1cF+czbNzlLVF47h0fA9lnqfkCIfcMX8lYfX/BFrNtEN68Q9vRmmx0NRvCC
SzirKG1UgCxYPTFF3xI9W2PAR7RsGWIAJ1Lz2uPEHXzmv4cope6JqsijqWh+CovCdfY+hGLIuyQ4
niQaEDKn9CiQpWVTr50lFRjAHHRVLMfnvULZUQVvwEkeIHEJjvmdtiOAhMj7pryouelQeBEeYMAf
QDB9gC31960KDP40QmbvTNApEXljkiFNwaJz37o+ujZK63G1t5pbGdZUsj5s9iMCQe3m6NCS+nOb
lad1opZWHF00u5QXzAQCDa4oXnYegjTp4x1wU4XnEPY0ON+tTIqXiaz0YDtIdJobSG7czd3QZWdh
tpt7rwsDxBk4L72r6PXJCQZyFbTAsVtN58CD7OSfD9LM3kLSFZOA2Aednc1jhTvd0xDl0FJbhG5Z
hAVrPjmcMXPTuIr1WChbp+dCj11cXojQmtaICCTxA8jthpRXi6pf7SzUUu+Qybf35VBvXP8shkfk
xANFGvsQm5EhRrDyG4v5VZsOXB/10ZiBP52a/kWZLj3d3AGQ8S10OuL7zSNpQhkOcBqCDKGutT7y
K1ymmclsk9Pk8b+CiTWHtYouyYWW1kbXSlgSGtOD/2FQr06azC8VkrIuqUJqGlAhtPw1QkJRGDGU
zY+po5NgL83kZso0sDClROzIdY+0Y6B2pBJrFW/G4T67a918ZMJL5TYx74UU7xh6PZOjqHcOoyxQ
9jU/hvalLx+x7uZmCnOBqpKtmHJexRlCk0TFymZW91B0sAaHqrfMnBxoZ2B5BeBUBB5f+VpeQZrs
cUvOr5uE6K44wkrVovcFz72nweedDnhRjUc3yvPtJEeuB45pX2xf21GbMF3cVNzmiw0tETjPeFl5
JuFV/vt8cWkeV5UYjGmeaLbg+Nw0gSMzz5kzFUPc03TtuiRLpneVs/0toLWjsVV8YpM6GCyW4cyi
JnJUPE+NJLmmb4oByI2ukCFpP6YsPYJLovseCBMFjZ+RIs8WXgq9zR2qPy7jMKFzJiQNZUIa0zXt
4hdzTj8OVk0xkEJvmCpXP+ixwXhRnS72LaeYbZFbX9TqdXtdagvnyTH4CECtDJSkZnVHvPzmMl0i
lfu4mIvW08wMpsRyf9NbHoSTAbyIPW+K8syNvtGjMms9dlbtRL6EVXAuG8Lt6uSOzQfeN3+fsHa+
BRPOor5CHipobN3c1Tx+mo5/GZvNtKVvXU6oySQrftZ8Oj8KJV7eAz/6Fv67Ye/9iedIUEOfvDck
TxSgzCelkT+apgSbB26xTbFjaCQiw5VAs6yGos30LxdJrI6HO08DkCXPY7HkWXBiEhxiLXAHHXqx
r7tH9uFbCOPpVZZIiENue7cpJxZKiSJIxgkkpDA9byCKqp0d7YUs/FLrRsXlx1OgvzSiqBuSX+Jt
dl/FcIvooCK2/NfUXWzfbCze4EceB1CwRTLUl3Zahs2/uPxLcBaKDXWqd3urKYkqaGlrkrvRIgPG
r93PYr86SvWHIexUbK+hjCd3smBH/LDa3FhnN0M8J4RSs8utDI5UOm0Cafu2QVvRVGXZ65BhpjyW
QU79FvBqlPshuboInWbkmOWxxpHZm/Uw6Llr32+0QdK916xhp09XGrbdDTw375VlkAYEuyISnB4X
KMZq9Ke0Wlwo9zXHG+EMlJeuGb2Z7Ekl5g4eon5Lt+zYVGny3V9uQRz1baGWy3xpAkIOCdGZ2f94
SktCJ9cMaL6YF20Ct2cygylal3/Wf0fsYaOhxw4lgLWFUmV2kd8ZLqov5B4h2YUzsCeVBqvOcPVt
34HGaAWqgOJtgKheihu+/pcsM39fuHOPI+YIYlGkw0iaFW38A/1QWgJQiJbsHYMwFyTCIn7GEqVm
fcVfV6A+0vbOplyZFvPbadglJI31+HBMXTHuG8Uw1xViYNq6fT7b+jhPT8iOz/tKYVwMWXuuXfXl
ZWWkq2Ca+cFY5A0JncwV8LEssG4bbJKQ+TCy6RINt8bkuO1N5oeE3qK3O/IEANe/kIxer5h72H3q
fuo2mCCbM8KD3QaAn88rJcqrTqXrttRPExP3FHPU+MCcFk8QDGkFH6EGjW3RKgAl4W5kgu2ZCwYw
g5cQLkmXRxcALif6LLJ0A+gEVxxcAj4fCkhg3ZnLNPISKNG52MV/qgQHsfbQct2BCfYhgmeuAc5U
7CLQrHn5bPjTYl6ffJvC8XqSJyq7si99k8e4m/QQYUtqztqYrAksfHv/gJC53lefibNnb/hF8CiY
8+qq1sZ6n+X3ro/G04F/NtKTEXI5S0pEstcg+huxf4aTvYjzCfT4Zps73qnbpOe1J1Dxh/XniCgA
ekTbgENzEPdeFvnSlda7B6RndubK3MkqkmaUlZUpGNtxYgC3auvsJ8aa1ZmdygcBnHce/Rr3BFa+
Fapvhjh1JCzZQPA1kxsY/E9z0KI6GHFjcJWpdeNtOk31g3FNiUZ+M35JKh9vviH/UbNrATuAQ2B0
vKo0eKwnpRrD1xxhaRel9zXrzeEXDFi1FCZhrZDLCFg9w9MbrCLy8wu9oIjOvNnxXJUEKVwV8I8R
Bf/HrXOFNoYL8B9QwT8zfVal56umDn93E8XJNTYRhp69qgi0XAvarasEjEM2Ahvp7hqhL0oY83Ie
uxVrqA5kIrZgmNAC3+qePSZgo6B0kJzeYFWbl2T1a/fHBfaAiF36bq7g023pSExgdKh6suI48CSu
tSBpEUZyZyDNgqFWn+mzbm1GDkBk7XYVC0MszScHOVpGewBzlRJiwOmw/BesX4eRZHnHaDLGNMi9
CHRI1rHlHCR8YfVGJUl0PlNdr/RVGzT1lJsbVh1CphpX+FTWT2UxaT2wT/6iyjJ3IKNVhMlXcrSq
+0V9R6gKF6L3FPH04ubEKKmw2zD8uToAOJ3R3gj1fktbFN2MSq3ggfZBe2YIo5JF1fMoQAlxmhIX
Ptp3hfp7cONfucTh/5tdszHDqQ16wS67ev0xg2lgsUzznP4cpraq+15UlMd8h1OUmJi9KLRheWHu
a5vJHKBtYkfvs7izZ29aW7QSXveIvAdczYcQP9xxArC2WF7eRqwLbEtxtHS//mjWHuhFSv6IEyFq
Cl2D1UD6QitdZN8kWUTOOvDLIxjtonBEyioCR3e0YNk4rPsfTvku4o915RpEhhe1WfErB0uMKDD+
mp21EzBZ53MYTsZ8IeesbL9gEnOkfXNi50gHWi45rU12PVB8tfw6VJsH9CD5teWc+tGyzancs7xQ
AVtMoRr7cnKLxxqv8IDBmWteAuXvuQhYr/JcrCRDigeSAgZ9Y8R2Kto2j17iJbeZg1+tVe/1fhSV
pm3xq1ccsWgf4x0Ju+HxVmL34Sx1UXjJVdzEeJjWnGeyzD24Hx5Ct+Ty7Y8BjqCHIBodGoakchUD
/cB6pHHoM3It7g+8BUwPx7+sPT4NuzrROQP9/lkgbbC4maWvGzqcfISD8vi9NZDhZV47SUkJBZxl
MgING2JxxK3i+DbaZiTjouKgtEKIx/tjHvQkURuAstysRJGkZpvT0pGP/dG15qbJStsLhHKhKVQ8
gculD3NbUC33XagEx/8iHpIz+ogGJ0fpTcZYnyaBIM8VzyiugOSXr/+DrAUoBIL+VzlcKxH+CvXS
XBEv+lvhrc1sjfrBfweVYJQDaltgVGLGsYVt4VzrNyr2khxT1uWokAzRvE9/S0v+Bbr6pw9c7JHP
E8+72wiuwC6xNcKFd0/STzp4ZjHUkMxTf0iSfggEWGdKCYWiblWzCAnem/B4B9ZPNbCGF6Bs1EvX
+4qQIgnpe8dH0TmHsLKf9FDI26w7RO2liSML2WW5rSe/ctymNuWw2BHA0kZmQg9KvyCRTAAouNd4
n3k/SkT6QYsnxOPUzjCLH/Y1CvpnlPa7cQ7vStTctY4qw83so2JazE0ud4wePad7G++ljHZmqqKq
2DZWISJrHTv83RTYdgml8yNhB1D8v5Y7h7CYh7KjHRFcxATchj8jOdEtoCV5dtr4WqPy5bFppOvd
y1F60WglXFAfkqfQ7PiozUfbTlUtS2tJ9TtjMSymVB+y219XG2Z11y7cP00WZT0j+nBditLlfmGa
QKQiNRKDXAjmGPjoUSxSbAB4yIyEtQ4Bnq4v1YdprIjG66WXLe/WfTbrEMr9Spu/Et4lC1yLkv7a
rDq3asoZWJtw+V4GzalVoe9KY1KJHp+j8r5gdheE0dYati6J/iCvP4UZCdNnNKjpTajkM0Zj0PkN
OJYcpHdpVCCK//qEI8rEBotldytScsBf++wVIYVWUEuPSjge2GD646jwEYlN0ADhwAxnhTt/xqaj
pUo2RfLEpSe9OtN7SJGPWPBZHFqy6Ny7gB1S4cfpm3/sdSKk58XIBLETlcFf81kEER7oOC6Q8J+d
Bk2EToA87bfRtofpwuEHkpaCApFiQgfsILI3y7v4lKaUV+PTtYK+DDAcP5EVyiITTweRkIv7igH6
pDom3O3QmanwftcWAe2zGlJoPCkj2daH6YBw/wFS51lQKf8gjWPQfSi66jZX6tygN3pQ/tMsGJW2
LarGCkih36+ysG0D/WxU3TSZU6XLsoZo2TrthIwdVvUJqsNfYqdBOlHIhtMjPFkJ3LyuxdgEtSbC
R+p/y0xh+see4/9pJQqzM7fvIrKlaj/WoRD9BY1uEfI3hIg94k46F9R47EBfmzwe/VnBDnJDJQdf
7cxAidot5YvZs+SG7XkeFmBT+CcBviOUdHipcMW5dYt1Rneko8mJPV2SLxzHmQ3HwMRcAQHKSQEA
JmlwR4Qvo2w0gEGy2u8325VGkS0/vo4aboQ6TgIh/d1Oq/6JXbRkZrHiwS7Vqx7JUklB4J540LWk
bJ5e+P98kJsPD5i8g3v7DMI9F0B3dgKqDn216LWpN5RqdV8DS8cRGtK/8zNr7urNXJHdKN7eOR39
eO1TQ5tezNgGV0sIJt1S4auIdBnBSVmvuQJ87cnADlmc4xBE2fU+nPNWG/oxhJzfuSdmLYiHDKvF
D1lD3CbiUYniusDglhqCl05lrU4zTE9z5ejlDrdJmLkMxSft4r//6Q1xyV1gdDlp4LmRgumNrZqT
e0vpgR2jYMJsYrWs6G3E0sNRqORtsILe8GzpNcz1lua+I+fe1CFx79xzID+wKQRRp8GehgklxJ8p
QEv/5IeWHwNZH0HPkx+o+p7W7aMLP7cU4xSuOP2OtaxpgD+N0KC0vEXZpY1gzHm3pi6Jyq5JQm1V
Yt9CgTR8gbu/28czkmwZcUqqiwtXx5dK6qFiCISqP1OPSx303LRM2fgtmR35fB4RM7ceHboJZehP
DCK2AZk0frV0T4tubotzf42aNII1ozUPdn2gfh4wsyocJGQE/LVgYUzOKI1fW9QFIsM6n62gfxr4
pNQLi0HZ4tiVjGx6Xh3N57Wq8aiPzC6Kuy0ES8K+HAA74wMIUbtBsPauu4ncGomTbL2q2LMBBy4U
cKWU9HuurjsFRQZYD7AscoDR4Tq95kCY0S/FdubWPQ8iXu8C7fLcQuNuirQJCzwLfQjqpe3x/5fE
vB/mjU1eN+Oszhff9Bbg1mToQKIQox3HWb91TzA8QRYDP2JF8OPPmepAVTkw92LbH782/fVoVVgp
85BKoBEIdly4AXgQaFT8WWCmdeX7C9Cq0du3OJwgDWzj+W9Fu5orELWi3eOyyCfSvoK0BPBGI4mg
1TJyfxgBIQUq5OnOFo86qTQrRc1QVNy5uGscP/t8n63v3ZkIA5BU4wDjdBle+aCBGujRxPE7ClMm
gXODcEk4ibOstXTo7HatKQuptfofXzMxXjhDK/y3NrdodOcuR0Xb1ryZUwi6EuSwm6z1NtE1h2bv
G2kK0AlZAxKYUihD8x2zTSMKJnw9lEtq6L/xnEKl0jd3clqthRwTvxyEAys659pAS//ByZEBFBGf
DUjHkC1D+r/geDtt+CbXURWqcpC5cjuL/5MpMtRjFzZdYKCgyTwBqICutGoHnXg/MDgYOmce4B5Z
WyamkTok3/Fml7rdtcqUL/dZ0s0baMoVLEUTbZXZbrB/HNSjGftObErhTtLzC0a0O/KZRltVe4Rr
AxckGhxaIqSBbja4az4gHjDSHlE4+I1wlWSZh5o5P8yy5KUrn6x/pYtyTXhyyUimqlgaPx5ZEcyd
f+lajKtBT64qKDN0/TNwnApgay1WorUdP+x2psiDUQMkYYl51uvLXM583A9k1/VzuyouLU5pGbfJ
st0gMKfgXZ090zFHNr0Miy5nWBkGoIKKaW9co4du1pHm99mzib+4ryRFS24PT3gqA6hevNF5Z7pb
UbP9t6PxT9bGvrgUijz+8/etf0nwJp3ZvXKNRu75hikjcC1x172B+ES76VDnK2e7Nx0SlqU7fQst
LLqKa4UJgRNL/0Sb2h/eT+4uaNnEIFXF1VvEttOp9yaBipNWZlWh5m8i3kBILpey29x26XNqyu8X
RdKO55XCEDURumCf8Qw648JDAR6yuPVWmGqwT5gMcDW1dd7SktDjwkmlDnM9u+OdkaKW8Q8Zy++Q
k9w4BnREErda5iksCsCpWNT/z0pF73qgh77xBKfPF9IkehdVNl7EaKWKssQq0FEgP6IZcwn9hHtK
aDLAUfRdN/sF0BPcXfbO0o9dxahaw7uMnwuM8s7dtxRIjvuLnuNvt2kV1tW7Cx1hAmnZHlfuk/ge
x6S5scSHQKfzUFaXTbZSqT1HCVSDmos5/hWmtEyc+aUyOxXrbpfUc5CnmvljFambJzePS9iCVkul
oYIR42/FGKjn1+ZOFALCpL2S2NqRfy3AO4yFh/q75bkde142UzhVjS5AeVN0Nh+nx1GOOIsIWHvE
wY+YurBn9M5cfu6an+lSG56Mj8eHxNw8T+3KbnqjDs3mz+sml4+0veeZOYtdZa/d9qmOzOoEc5t7
AUcL6F5rwPsD7LnjSlXRLlId7o2/XtzwgWCGFXHqy2fuOuDTonQ/d+TIBGvvCxtR1R8pKd1o1bCU
LFefDT250dZYDMOkYBHrSYcTTcOn5qynkpfgqps05D4UuIBy2l+xHILH7XS+JVJjaHv8UmIPOQKp
ldAyskemYqZZw5dhaRb3k7M2VQh6KPc4mwffRJqTmNYAMZMfxvBnOevX34ZLeqXb2KY7SfDB+6ce
mH3ius9lnFnIJU4nI00Bn6d86ymVjXliyZho4SAf9pznZcy2uJBfPJEIbxSmgIocIwlFGW6pZmze
d9fmkz5QJdk5cUL9/KWXLrkVs8i3nqxqgZ5tPxMHO4nOsGWIs4G04rvATUAWaXS8+nxVcYdecG0I
iqS+wDtUtWTul4iy+kGR6JMraiwCXERIcZ4RrOB5BpCpIOJrh0cuOXZjYvEHB9n+5T/CKOuUR18M
jQI0LZu0C5nrntvYwapj9iVtnc9cIiZEsnw6w25oPa1zwlUmx2vBxVoFAgu4qLQ6TzZoeU6RLxwb
fz+jzRjJeN5CcldVLAD/sg7pTK3FxE5VwyUn5gIG3bB1qJHhD/imFJZMd+IO/491pgQ53YTjMAPl
97iHlzDFf2GMFDZEBH8MsIlFPz7K2AjNIY0nCLLYsnGiSUiZqUAufyXRlaPux0/DBVvNnSIApw/e
k7bTZvzXDl+6f20vT2YFlg6vgKpQXwE51VqjgtNOmZ7na6VUd/A/uoc1g1NjbSphMEnqqRIIubwZ
wgkyYCbrr/OWG0rhGn/RDkcXJZcLLI/lJ/eAY+GRKoSNBRipL3MeoBp5eyQw+vcuvcyZTYBF7Y3B
4QWats1wMB3NIXCCyUQwh2ilBA0tQaBjxIILIP5zw+u9YeJ3H22JFciBQX1V215eRvXnllJRuGYL
vhNQEdSzR3SZ3gGxqUQkusYnCHJDT1wf2NclQizU/ovCUxJAAY14LhLnRE1vqs6SRyCV56IEQuwn
mcAbip5Tl0wjuPxaosB5ASCfo102yelntn2/o4T/PweI3Vi7npsxkhW37XPw9v/88kw5lNAiYUF5
A7oeMPnGROn+6j+vGJXQWdlodLEXPuJsvs4U+U8+pfIPac7Jii7IW9sax1ycUASuV9UmioSa6T6q
Wj1R8fnR0KLOQ0n2aDJNT4xkeQPzJAUmujmR0MxNkIG/JoTy+RaGtzms25pWMimF8B7T0j3dxT0/
+Jypnr0RPiGUZFVPh01TZP28uCG7/cwJm+oc/8/eqlddjdaA7i+Jh7zIgwTZHRSgKcEFGuOyg9Dq
Yma5ykT/9yNzH9JnY/qpnO2OnYtx8znObt/eMvo3DbLCZFReEEwL9QZdKGjOWgZD0jAP7B6SvkkO
BJRddpzD7Q5oLzrqpg+p9KMMcJCuoPDmapkArW8/XDOHrVwqvo87MSUMsqNavjZt1LpacyHvI0ON
NXu6864kzeMQjC5hZXUnoRWcrhEBk7JkXbEPStkyDuaCZshrXnGoK9ngyOpaM7B68tCNQtDjskVT
W7RzmPzoeNgXbkw202KqHCNIN3QBSSJq5Scg+bGO4kgz0phBmio4Y38+MtGy7jvtUKdzkSTxPqof
hL3GJOvnL3pf5h6DX6mF0MP2X02Naziu4tR2byERDvBxmZkiTyFdu+xShoY5j/LDxPS8NXUkTddW
CWp0eB+0WThxqEzUsiasU8nGP3ng2o7Erf9OEDTLTAr6BgRrIdCMXa+HMRmSyWc5gdmj0jjP6sfH
3GZaw82Y4d0F5QbhSTMWrDejBq7AUfLLJC4qXXtTLNJIA35KpzTLlvg/q4Y8nGx69jWb9x/z4TY4
OPoYANaoq6SVOUjWDB0g7zSOOWTFeGwVU0hyWQnXl7aBEDIc2CDNorskpeSKuj72fCenJITG5oxN
6aVspTl3dcaDDLzoyA6yu7QbAjI8ovqojWHSSJQC2/1NaQDFo8mHiU/eqo+MvIDY+s+2GHfZBm44
TFvoBgvpS8YJL+r/LUPIt6v1QbeoD39R7TjraRwab3Uq/6HAIHL/HtpTY7a8kQ7hr+dwufeVw91a
p12PD7VXrpLbqJ6Wzibdojfx7F/+QkKETbgBwZkYBXywXC5/wu0V7ju5NNRsgYlEnvMtUF4NHKJ6
JJGRo6nu9jBLGeGpGqertI4HaZCMYm2IUGzg6uBx7Y/4HhpYteBwlyCMIUz/6gC/0rA8wBP4qANn
vEa5OhGnLOZ0fNvvajMb5GhLiQ5BYpxSHE8VZNIfFllOeuEK152LVB/BT+dhMFS40k2YbJDkqhS+
dpvelslCT5d+hW+7Nql5nCJrg/it3a7FCX5Z2X7QrN1PrZEmPZ5wP5gO0leDX7UGGQAgx8KxUKtE
RNekDLC6u3RKyOc6Mq2BV5lK3pnZp7iZF2g6svxt/cY6PeRmCNUq3euysbEMxqoyUZC7+0MAjGdU
9EDIipPZZd8uBPlpVw+CLaXX6XjoypGH0SdxjTmMPXkptcGHKe2YQkydBqUiJaQ7hCygk/y1Hgqp
7j2cAD/Rx4H78NRY9dyXfhNRvu3aIx+6fpj34+w3MppJ1Ip4IUZanUGXPfNKBWRpGSW5VmRA98AA
bfhqjFCsywbZi0o5NhLxdLxsiZx/8Ol47p9YlktZawKXGqNBBgjRxcVJb8kNWZmOZKKWbdysQTga
eMoezRGyvFAXUlX4oiZrVPZvBp0tMHwqGV0RVjSJbNvSxnGyC/0QzUM2g2X5yrkIQblLJAOPDCKp
UXiTLD9LTqf2OCJMLExVb6p3Y06R+xJjvm6O2SNJyB2THngXubdVDd3T0MrjZOwnWvIaeyFepdMH
BVPmkgqdjrXwcFaZhLF5q4ZDOsRVLUct35ax8hUwfKr+M4us41+V4nt59DI6PJjrgThwvtMhtIu2
JDEjCypyD4LV2ZmtsUjmwfkWlxH2rn3nGlqwSSEtc3DgvWHml7P5nLwVkOca0WUO5Lq4xgdbDvy8
g0uPS9w11MpOyTlsNOusDF2vBYNkJt+huFyJge0lifzY0t6zZflfJ1WVRVbRI7brnuKmRwZYB1x8
D3nnurfYN1gzW7Ec/wtjOk+yDTLYcxrIe2j5g9mDFEAxmm6qrfgaIYJBi3qiJEdzCZ1MReILKud0
Xm4wBf4dEI5MD+ikIiypJkhYgguhflHHQVfYj6kyM8DRL7L4h+pXTjho5m1EnuiLPSmnXqRBiO5l
48ghxYEnY10nI+fEc10xdK9tFLIRk2VyUEWVMBzTT8YlE5H/6WtEPzgXmGriv+W0OYWmvwvP2CwQ
nsBk6Zg+vnlvLnoGWtypbxXC/O0aJXBNHoaNnPyT+8hoHSQ2VDSdnMpiz+skjH7lisOsTSuaa7iF
GaqoNJNAhF22kLjdsf4C5ZAc2ZdY3ah2fGhhBCGEul2JNlBxj2rZjY7f1Zs9+ILZd5dwA8oxSKCq
6eVgM3NKjSfec6dl20cQq4XAu5RciROMskesJD/bjCwq9V6SIYqM8SDJk0bk9RifDxc+3MLVGDtv
YK8n4uGhB+59yuuTkouFrukn8noFHgWP/eZHvsT5vs9e8CVBnAw70g4v+LhYX3e1vKd4Vzl9kQAT
TDVkhokldn52OcNO3EU7tqDtwMsVKzlTDh+7ojsKm2WFhGopxEPTloI3k/oPKpCd6F2QZfR93aDm
g4DzdP6OWn08SQfBgZhOBu///cJc4mz1aKrL/ub9MMmGY6Q6IH5gc3jckTI07Km9ELEfrZ92s7g3
9u+crQ04cpSs4uL0cNAN7b/8pRSYT4LpyBplXMek0aovX5mVMNbRw5Lf+L2T5TUkJgFxf8Oz0we1
tGVaSREwI5o+myK8AkgyOBvle24BiX3I+zvf80LjEdfGjbu9a7nrOaZdlHbOwrNQ7EJpFwQGNd+T
4Vm+66pnWcZ/ZXVXjxnNPPUmaqGTVHEc0jSY2M+XfeEF3jjjttL18wx/D77Ci460c/qCvAVShl7c
jFYkggRUUo1/F9Ysovj8tBtyVw8AJ65zTWeWl3wdy3V0pjSMUN8D8+kdc6giQ7Ds1g3gYwPGAESu
q1T4c2tggEUvsBN0EGKHjHgcIRo0euaufFNxCn9BNtdKQ6zX0TNAbGHumovOECzgoJFdnBdOrvUA
75FB228/KLLGYLgPbUwsa1P4eofkyGsG/I7UF92OJRRmjnQ0aXHDe3MNZkJTQfpq5dkSd6M6ExcJ
4TbAEEvT4HtzSO8rkfThTv4bRo85QAJ8yajP+RUa91ahRWfZAevfGU95S3mUFsef1v6/uxU9KYTS
wcTCqiYRiRI32v4vdrcykpLNgvDnFs2oUc6i1rKGaJrele9D40eoUqBrrfaUGvjgLrKx/Y5IBs9N
k3jDcrEVw8EQiYDRhDBt+0TpMEvux8M2qDZiqCXaOxDYi0wN5rbDwRCCzsfKf7YahAyb7nCBXL5r
Xo1lgf6SCgX9taz+7BBZTx4mZ9txkPClaRvY9hUpqBdbxq3fAtEnF5mzyQSD21by8u9YeIILU8lL
9xxHavYmIb3e614n1m1dg7iZ6l4Cx8YfopRjAkuWOl8vp/ms2jILibP0rJXXukikzKSJEQudYDm2
WVLysGZFEfmjvFCQ0XbQ7bCQWk8dUEwUGU/NDR/TAcNzpayx8y8yalaS/76E9ws0wGrHwGKEqPXp
MfOTWvydjRm5uNzHptOePQRChRCejgXMB1ixVQ6C1Ky8lPZCJfQPibWVyMnxT6SaFgdxdT2y3TFU
9omQyh4yvcZVoEt4BMHb4PHpO3KbTFYnccaFenF2UCItJ5eH0g/qAa9lx+WHxzM6GuxDR39JQOzK
HPQF6yvW5ZEmyEEE55wOjdFUzJEMCUHhwpFAtgaV6q/RVNnaI6e26X5O6cSTUf8/PLomCIrDy8iv
Gbt3VmI4QDa/WF+GZm/Bb7GFnlXIBIUEgW40zvgQ5YyS+BC4ww1XwCLVtBHV93XPl3vLKDRnF/l2
CLcNM/Sx6uKL8Mif+aqB6uqi03xYugdLCs4643sUy3+dFqAcwOsWPGmfi4BlbrjpL/oeCEgT6eYF
YPsfNcnYo6lJXQCVgAN4NoP8EEvGaXf/Avp8rkR97Gki/ijoDHOaldhGC3F8+30rJIPdgFcNZzDs
Aup92bbCgxkqM33DDPSRxSx6cs3bpUukKF+zxG7f3kWQfSl0xTXU3lhSyikN4jGfBVglz8MCTVES
Mdg5mEKjw0GV2244ZruAgfjdlsIfvmH8jFdx1br+pxsKLXOr+xG2ak5OLXsjAKJ7w//Pgrv1Edsy
U6MTsfNnJuU19nodz3Z305orOpT4a2U0LRuIjLsjXv3RQp7/tHqdFv5JLtbHU2KjMWxSI6/NHO5z
QOwxakvARg6trl/NqCGM4AQpOXzI+b/ODTI7Rmf0zjkefTgn/Ua+r9Xf+gj9x+vLGLx33kh58+9f
RX90kJxP24qnD8uRmegawZ/1xD1GQ3QrnK3GfuHcdiWKkO+WH5wocaqiG5x7qLhgk83eU43qZEi0
Lg5VMXTRlU5hiD42TbiEOuwlg8S/UhbL8CaV8hfD6jyD6F25G9f5iYuJP7gQcJFnPfUg9YGLxDZI
aSeSPEI9Hx/OtQmaWVpawKCsQL6X/mtuQmJ+/T6SuK4do8Dxv8eE5tnXnhsSoZXj/Js+BLmL1eEo
i5HebENNcVLsjWdkgiqpA4d8DGesCcJM+A07EKgImDedJjP9OEk4nerfIE6/4v8srdziksYXwGax
cx6auPfL6fiAjTRTUjRjMfDevk5HeQMpkIMXwb/dM9edK0RoDCF3Vf1nAP1wv+oYNBcoyLHQypm8
xh1hP5hiKbZ7WlAvIgRQqcThQFCYjdffN+EI5d+mx1uriX3MBvVO9pQEHkrsXeY8dcvHag0ptA5M
A+k+ufzFt43VftI70Lrvkinxc1lUSvW0nxQY7Rz9+bBgAKNUKZlznv7Bc6Dv6dUIpcRhgh7oLFql
8JTiud3TmBdOX+YAxsCEABE6Px/jIieuRbE38+hVl6DZ/t6OzrH75PpFQokoctwGNH8HKpU7V64G
B6T6cFkSE9l15aBMz3HqA9GgtIaGVxLLkr5+M9gY7TBKm69ggMpxcn9gsF2NbP+41l3qnHF+QQU7
tGQi3U0m2OYQOjZaIW5hadRd5g+swiG9cJR/QFCTbGmdjamzI1ykPuTuDb390OCK+6WN8gJgeIp3
Ql7tXhby18iq9p+2hU1aBIe2iHIWvaELvFEQNTIzvR+I+Q2Z/+TCHpT9PaHMsCeKthYlhu28ECIn
b+LTVBcJqW3avYw8EtJqpZ8SNmR8TWQ+zGa9aBfWVc2blV4LcLvHXj5VBOE2Duj9yQf7n+rCTAH0
LFPcOU+BSoSELRSX6fcJjF6gXFXH14RG8SupCcPUPKVdsU7CpQa7rXBytHlBBA+LFn5RiJx3uxtu
3RCbfiHcOayhyIJpFPNQWhSAGgdpYVsU+9XfFbRStuHrHwNCGEK+Q6gqec6wokYC4r7ZZIpF6BhB
CF3EV8nHbfPotL0O8WPXJqXpHkdyR6x2/5h0cIBuhyuAZWZ2gchf0ADfMdPS5mTDbIkrisp3EpeR
zWMM2TXQusMYYllEcLbfJiZTV7IIq7Ym6le6VdTYK+7aIpoRO2hnXEcxR/A11DJOWC1luJhlfq00
YbYWPV54aJE5suIOrO/llSibVyhA/RJpRv8aNVxRwli7REyIqyovgeQCIUrO/mf8yqPjy2bTkhbk
g6SaGp87yYbr5L8HhGRISQSMWimtD20Pa2qOd/FLg57XlzmExby4iSrNJfgHAMAztmn2zb8BN2gP
w6Ws2X0GibotUI44Bn6A3fecrzXuYHRESay/xx/P4j5ynB8+7cOnTkHhBcU8kd6+7DEhQSnWbm4+
9mNSObnc+5V/8UJUmzEJKlvKzbs0vDFm+qy0WzR+ZkH4aAzMmwfam2updckwg39K7hGJPZqPUAKu
eED4XxwSjkTnTfB20I/pGPLXY8EKBYAAjDmjZKvgI5PMoGPXLCFL6NRa/nWAlx0qcgT9/o1rDNWK
7RCG3y+mFk2G3giygv0marI4pZCgWYDieDe0PuO1iRcKgvZdCTLjVaxBz+U+tOa5IRd4Y1PIJmzq
WGnAYdoL9NwfsbQ/1fJZJ/EKDsVC6O21hqyC6UTzMt9VoJskNuZB9FRV21ndLKYvBAifiuhgXSuH
WmVEicgpJ8YofatVCqnZuZ0qWupahLxsqCk1oe434mak/HwvAXmAU4YHFhTzLAeWbsquoeu6YdOA
6eLr321kuLREzl4rS7diW6LWOR4a7Av0bAn1iIUeb8NnPBeqWmj2BMuVXJDqAbbn5RsCmicbBk7p
6hqpYxtygOUo9jJheTi59+MIpLP31y/ttDC9Fkha94FkEO58t7EO0iq4f8Gu8l4YL4EHiR/6aamY
XYPiS6gDuli77hjI9V83JvmHXt3RLRD9FtflhLpxIu0ja2sbqQyjA7D3Z9aYwST3XbHxje74NJz8
bLNvBFPdLsnyOjLZD8pj62MI8eakctN75GwJuJoEbGTfv0RPgYAD8qkB5LUhGrXUb4Rl5tmXTrOO
1FFWbiIp5NZ6Hlu1I+Vbyh76QoQ29CsKcDxlFELSgJRY+BEA2n/Vzie3rOE9Rh/H6dPZECuoppFi
v1bLXrlzWWW+dCAgj5zKjxnC3lBlXqZCAWToo9qI+qHlLiuxc9e4tWl/3MjB7oOtK/0mpNaS9ujJ
+WkdAHr9ScufIcXIVGL3SAP5MucZ0U0YeH0lpYXCMNZRgNxvYSVU7DzLAjk9IepyY26IKeH0USdP
yj7eHBXwfncPCkVkSkmfbkkb2gqeE4qBn42iVIZN5Mgr7xu3GN3l3IhOm0GQR4PsJmktkNwjUCMu
EBWSYqqJFsvzcyvAs/Vq69ARbutfTfcIcQGG3YF2ZN5kvP2Q+xmHXW0DYO2KqfncwxpAXjyCXwAA
jUJVEBug4fC+r0LYKhZnXHr3zdfxkfKdFwmwkPEC99eBMLRI+KOVtOQ/049BcaL0wXn6lkvd6zB4
6nr7PUdMAABwT/stT4OWWfbF+ultHfCMdOGVzGUoAfV/DPL0aeoj2PjZxTTqQtHX3zjA+m27Go1f
PpEuAuy0uY4U1T5jb2XJvKXtPljHHxbxc/wKIU+uQ6/79SB8XU7yJeH8msns7uwxpTSN9TbdNOn2
SVmgwnsZfcJakDoQbx7EQ9QGuPUfHG1ya0sgtH+pS4VeunAg+MddkVDwjX4EHyo1m0wCO82Lji9f
+Zb5E+WmIzDBNJl2tBPfXp3PUs6927nzEcorzPUvQiIZmXBR4+YZPg83StJlR9F+mLT798ScPk1/
tPH9Djrl2GFufIJ3/ixmS5Qi7WKH9viJ4uErArZlZeVHqus07C3PH3QppDafX4p43xAMCJdSamLp
W2wbtJv5KJ8Wy3/kNEjUWwtbWkqSXjeVnq+ApmKFEBQOxIpof+6wbKnkIMNaZJvsp7Jndwf6uX0P
DXrG62HIVOJGTL0F3XAjnXBI5eO6OcR4RftEgXNXZJx+O6z786DACadXAK7pjaMoMRml/d/hb2gC
eRv00UYyabh4hYpSTjD8ufEzm6sLP31g7VMGftia3LsoCwx0vnrtJ0AhNRjC0QUBr6qtMYztmszx
fxGhLkRe2so6I4dlEX8a4fLHingHKrQUZ1B2m72HBp7fbiv0HrJWV+ewdf0NTgetejWwS0hTzhk9
6CYoGmAi91ncqnD8MXtJ0OQClddOiFw24sMMkiUuh/MYq7b4KHaImNvTKXYwn68LLhAmMmZsjZdG
KWqPT2IZaazwSAbSfIMuYdsc9rIzm25RmoNyRWletXCxeHuTjJoA83jNcjBp/WAdnVddKiYp8KUj
s/QZqjN0IpAFztIHXE/dL1JzRchzxrbS+p6W5mFUv5jeO7LHStoerLICmrXteUmv7HAbMSNL7/6K
s4djzAZvIYckEHN04gyf4RaShmisyytvG9ttlTYmuFsmydwMF46BJgMb91M3qXvLWoLz69BS98rm
GpHLe755FE+zlpHm8SEEz6RlwUb+vkBfxC+tL2LSt8mtsphoH8JE4Xs90BpySGS6vqJ5gq2PDNe5
bKCKHBYNrW78sVDVVpROa52cFsmX+WDOI4EYB7Z7fRIugN/azSvuO14kUcrbiWj4RZKtgYLnHUbb
TRK2va9cVO+pN4NZkG7TAZmM7lEzZVS/RWoWvc6FPdkhlqJqV8beZakOeq4Aw4U0d0liGiEp4YD0
6Yj5f3reEnJ5KE/s9JuJXsQLPxp3tk1zb3B8RkCQ3L03YVsEqG0WJjpWZ1SQ/IEBFEe9+MOCimRH
msijPFssdXGbXXbHPBMK381tM3RTAJC/tQ9GBzYSEFXmKl8436y5FtBbsoYjNA47SI03ulNYrRiu
47GcpHNACH/3bc7zZsk/wJr9yX1UbYY4TqfFEpPLaZP2XntU2NJShmS2vuj2rjo4GZDUEhmco6tC
NEmBm75UpB1UMpqN0X6Xu86lJUq7pEHC8MCmlkIKbGRr5PgqBd+HYZOxVMJAyMe9TV7yE2w5cZpL
NowiI5JZ+GDkx/fgJ4vmoNCbxmGaWh9mH0WEfy8gPaM6d0D45FxkI5HBD60C5cya76OB5cJ1xw/V
6BUGud2OtER0GIwZE+SFavuRUP3aJHfHzCIw6g9FFfzqHIJTuQJuPgpXezigk8Xa1clpPtPrDVpT
qlemVimCff0DxZTvF5Tdq2AEC+aAm8p9Mp785IGh7PnfzKY0aT2wJknAtoJ4mFskwCNqaDxIrh2r
eifpNrZ/nDuIDtP8eFoXxpzKUr0poEh4NhP/DKV7hgYNMpKMQfTmv2QglLZ9rBQJL95iW3wZVn9i
4G6FXI/Z65swvji1cOpEnb6PCB/NqTBoxZa5x+CXZpA+qJgxzjIUOQ5T+PxZoRsuzi3CQq4ROPdU
vVmKQKoU/A2XnfGcUYGb9r16/3udFzCr3Qeu3VTG0xkIN+DqY55oXW/fv5cHuhnAtXFm+wgT+kVZ
UNl+6szbkDMKGLmdPXOxQct7yQlmjvHZy4BHOUtTA/+tqOD1IW0uKvTEr6rI8212wNZDACnyLCvs
j1PZKCAWmFRyw5igD4+u1fNtSfmOG5uSDNfHexYivolz+wneErJAmZpRZrouBXh66TlJx3e3C0TT
X53dqbk8P3Crdw8E4VHXU4jR6bKXjL/VDe/V6jVEAQdJn5zUiT3hHVqEx8IiP3ThdGL3s3eD5/ll
MGnN+2oiMcCLud/kAV8oTHwmhfN9eWFXwetgZbMw5LghfzhzEvhi6O0Hn9xc+sDA2ziucMm5DLi/
m6U+2sXCb4b9O7L59Kf6prZ509L/JbaUz1hzHkKMjSKdq2UWQUgPoOpDnoPFDhg6zog9/sI8URu6
Pn+qJi9NomfweaqezWF+bG3VYj+ZBpHbr7ISvuhdM47S/9vvAsZYuDwSAKfxg+Y+tpyQ/+dW9421
63w3aN0HtjJMs/Kvd4bHYnkHxz7hbLudrPJ8COvgiT8Vb2fN50JhyoVZrUlnB+hG0OOixOeWh+oS
Ruf2gMQ2qD1MaJh0LZvOUdGlWr4jeG46lWmwMJI06fA0oK9y62x7ps8SmdKJfObRhf7n1QFiP3XN
QEkajul8dzwNTrnbx0+h+DanENqhrOnf8Rc7o98FnhVw/va0itJA92cW0gg8QlGFnyckEdsiDtoX
sr7Oq+SjuJoOYGNBjfMIzcFIm+pNa48hNY/XwyBkLE18lxUcA28UzB+TYgVp+fIvFg5MqrBz+dvL
GH5gBLHm3gLd5SSx3AihjbZM7KcwoqU1aaWxkko1dvVJCGDD28KGFbxWTjm5h+sjA2zs51XC6SPK
JNegc+5jOrMJsPNI3pycZVxn/3lCWwxrnaZp7sdOvslMm5FOt1nR8u4MTh751KZgtCFzGgx4rK8x
F3utn9r+zEtbjc6VGtKMmtUY1/lKuo4RErzWjy+Q7AMjtr9tN+KOObIidaaDPsDd0ktOydI0chcV
gUfSgEhf/JfVnvg/jVjwtoYMdlhJyIsNEkyYSmUvMXTacbfbT2PX01LigRiB6VuoxsccS7seKBvC
oJu2nqsy/mCB7OGGUZxCuw1L+7dqYfWV2SZCN5ZIFXASPHAfcagPQA5jELsIFcOQwzxwJGKZOfWR
39lhds6AqEIuZZ89JOQ0wumclP4yi2lf9sF2+HsK/i4xxy/LbFpWSIPlML8kMGzqw1ECbEvAWIt2
5T1cZRDkCNFVDpvkCMRVS0Zf2DW/LgUyUHIGYPnUuxojpB0vUGMWPeqHHhvH64seiUwDfdd4gcJt
AK5X7ll44oFcKuPyk1ZDnMF4j4UgNZjw0CglZhTBdaotGM59Q5YscuN+SHop9Ioo0Xy7nwZ1BWVD
NlP0CceUSUusC2s1JVsVsCmiC+E24pZUEhaHNRToGFiQtSYAqJSFQwhPPEfQzK0tnXCHpq29vSIJ
xuSDz8ubqTuqkhoszf80s3FUEX7DVVUP0/abh6tAxjZu+3Wcq0RTT63rHysA5ExxeYFydEYE2ry2
ivin+hr5aBJBM8idhBzxKK4oBWycnvVHSi4rvfx9vsgEYaC1Vfn8u7XSVsvFtk0JTg3Av8Shs6PC
hAI5hw5CBAz4DJIQobZRH++OZojUSFDgzU9T5sagbQl+feZEq9ZQMyRlhkrPC+ZGj7T7VKKsiiSc
w7/jzK0Jh65/6prvugngzWyYiu3SImwsGvqZ23ulZGkrVRkgw6TrTXIPTmUzaSK+WovMbtbD2GKF
8i4vSyBYgEnQ/qpwuvesWl/GCUTdc2Pv1SeF188IVqTTOUzK5Cqpbi7WgV+o+HDti/exnrFKeqkr
/5MS6Dq/nEiy2CR23wwcjMIkwsjzkll9DhJV+sFT7cfcSjcV0A+OXcfeYZ+dWFc/mtRv/OnkXz9A
ZrNo8Rm+MA7c17K2VAmb9w2QKzbPclVQ2cdPqiuxtnMHbK1q1TOzf6Uq0Xzgpv13hUlkONKKO3cd
yFqlek9bnsErEhSDR014/bradv4pP0qzDB29EnXiyqZhoFwCUtbTx/lCY752QsMCL0mYX9ijCYiV
r7sP+LKOqrAIpWKtXl9WVcTk2FhXsMlQW2Ypv9QZPXYZ1qMFuEmtdmDXoqoyptaaoXHQQgFqHopb
6psvL4tdLFZUkEleqX+KL3KBNk2EEEWGyC2qT8rOanb/5VeUBHj6CdhybsDDx9KGwyoDZFYP9E6k
V7y707lVc1N3exzTZ8cc6+0latHBHHi70fp3HjNRlCIsFmRzH1kLmd+VSmhn6fvTvxwdY37zUusw
//zU7hLCgErEXJ3EBHZpm5uzhzG/ZouTFBEBqA5qS4SHjn0MCPR2wYVgtNJPinsbdqfrEaBkZkC9
kULvMtNI4BiYk7ROk33+2nuTA/qhabBs4ftpgSKoWPHP4o8HdT2eVLKk5WWM4lwqwZh4VrnCkzHr
xGkc+6OfXo3eqkZWwJGE8UZ0QztqOo62NFdnYTc9ztNofnxZZeUaWxfe1Uz6UOFdoO7In/ECz8xI
OaN7X8i4sMQVwfpuLf70h6DZ9rS95ND/h9e7pdVq9ePPG9YpOBXCcIpjUmyOsMWfYn1IUyNF27uQ
DcV54kLFdTO7EZW3UnQ9N/RMQcJQbC0yiXp+iYAmZRH9KDISnk6USeOBGICKgD5zo8hfzbl5W9xo
CE1tBa5ll+C7PpX5Bgys/Oa7a/uWnKh3HQ4lyRjCU04jjUuX31WLT3Drg9Qo2Ot1RdzsW9Kx407b
lVloL3PdjOFyXUdyEnPpMI1KITPjRo8Sph1ijkf5v7eKS0gN2TuvB5c/a/CLgV8+N/1bo+ES0a5m
Skp15gj8f2u7DnNpRXKQWuA8bWu2Tm9+9vDP5MSbbB1MUrc2HhEEQDgiP/S8HclHFD+FpUlja91d
/TFYy4zklPxnViH0I3BG6Ea++bD9O47BmPiPggWtX9xA1KwyCAyrKsAZC4PFfRHXWcniLptepQAX
kiVx7CmsqzuiiN8lmzwbmrturZyxKE7cEiGJ8a+RAfDDnlXYoGGE4ill/PufZb74tKFBWMnOsWMT
tu1bsTZT3g5BccNIxz36YpjV3kHFTGOG+xXrrkNU+xhR56/z0/76i4db4581ph73hzfHSWDQdLrE
B+VKUN6pYknmF7lqHWMMKgL7dGE8oZR4eI1WfpWDKeU6Yk1gm+1gEda+67nSQdOwLsGorkoD02CR
lLzR6gMif5GuMex+sYV37wf4fBkD7R9GEReCOc3wJ2UE2y7wAFBo0a/80uVXqDy5hEKpCFMEiYPZ
c8k20jVeHHKcpYaO0qxIxIz/hBokysN1n1NywVPNfrdOOulYI0RlTD6HgVKxBjJXgjhJ37NOqe06
yNDYDxgELwIzntpLQhy73UwYNd84equ2639tWCZnAMJKlEh6zIqsohKeI94/ZGfcvJwLTzSaPmGq
koLwr6HoCM5IWWqYj5TZllBzgyDO1fUGT/FUiHLZIwMR5HJkKIWXFJ0syJFrXIb/oYhghNnah44P
vOW2e6wkOo6cn1NWb6fUQWFoKLzrr5AeujvzVo8knP8lDaTv+4zMEiat5QmJo/L6dEckQKlotiKC
n4B3pNK9b3/pvvPwhSCgHDIGKCHohw4RyPEEFybXa2DVm7G+cCtOnY4xKbqZj77baoHFjJX+jWpL
ddHtzlmZuvBo6TirSZtWwSUmfztcFnxQbxrnFUOhk6QVLBjU7uYSynx7E+PsRPmCvTIO60sN5Bi9
rZpr7UTDI62OncDEKMacX9wbF006rDPWHL3qXJhxVoGAHTkfJNtWZpQr5GBUyEUdAHrAxY/rgjb/
v51DyjEEc1I320PhjMLQ6oSPzHJCksyF/AcbaXfeHtyVDaRemlVr4gRrnAGfxx0lfRycqQeuuWGh
vEeDXdu8MmSoIkfRC1FxCm8xb5Dcf+FtuWGqobocndnqmj77zKSMe6qTSYxgnAh87hf+adDjJw7v
iacY34J6gVyLZpNXOhfZZFq7sFAi6EGQG56vWgr86XmSwosuOhWYXrDV2huUXju6/Rhi0wM60I/7
XfW9oZbR0She3IexwRURLof0patUsOXzev9O9Sb9pa1x83jL8ZmbKcoduG2n2wLCdr4SQNbn1xWD
9LrMgfw6BYZpRCL5GcLtYmLqnVl7VwAEKkaX8bmPBrNIQ2uDWTyApgMHVur15akjo/EYZEJlb1n4
+KoBtbVvQYYI6fIY+iGrHynX/8Q7e0kZsP+lEErhEssUJ5OBClMTb0g+kUiUnoXKTu0fCBMZAEwc
DdUf3bYvz63rf+7K/9KFxGsDWQe6IIb6KZodxB+VhC2ZtMJGlyXM4ZoiLm1u2+qLfCYu+Au4fG9A
j4OQcAwUE/2VDXTM1gRSG+PFrA+pvVzpWRPILEQFl5GeZ8PRq7OEJECZ41zFYKVBCE5O4MSlxqhN
vCpL8blSsnsJqHxSDL/SlGM7qdv1RG0VLjjP49x63+JzjLm8ae48oAK2+6KpqA9Mxg+x+J8uzZZM
rTPjTiO69f03iNVr7pmr5jrYrlJMOQRzaHK2IFww3P5+FSGNYLv+VExCa+WV8rrvr9Md+WSFvzK1
xIw8BLpHri/1POh1q0/J/Rhzsp2/Ye/TxxHSYdRq/5xX5TXRQJphfxCJfLb33MALKHWXYHvDyuHi
SfyU+iGESBfGHFz4y4QLjxrQtdI4myNLQzFgl5ylcf62mUEZ9YV6EBIV2WhbV70KPU0j3oCjqIMs
eGry8Ui1B0sdgKOsGZ+Z6qRc9wY/B6Xodt3UTaynKUOsKMDLdrOL0oE6IhexzJbE+6WTzhCZS4+F
4qrqHkP4tRFk0AWOOVx2OBIym1ZItQognSMJXAMJQWWiL6jBb3s7sW99SN0ayF1XkOEPRGcWeL1P
wNujXLx6gAKihRv173RpIRTwtMwlqw1fQRFZU8cp9XgWC5iW8bga3LgYr7gVyct6EEB7AZGVal7i
Xz8X7bP1Rt2Msn7u/PDo7jg0q8Xfd+DRS7X53rLhbdpqN11lFXXJRN9Ewcw+9zayhT0jpf9s6zPe
JgKJxuFDk254R7aWbmF1anZbfAC0ezJLi6s7WRIPf+bf+y6ZOoQlAQ8T3xOT5kka6clLRBSluQYB
j6tnh8dEC9FAY7H6NYv6/D0mmrhDzGj2P+o0gKiK5iI7PtSoADmvnc2gdFrEIu5za0vPjZ+Ze/wr
MZ8vxOTtMVgL09JQ62AGuQKVWJxYzaJpdrQ26VU0gdWF19brLBY80KsvQOHf+kWm93OUNFKQmCMU
Z5oZHPDN3XNSgNeuZOsa5LEFDfWKCfA18h/a4MKDm4vMsZvsYg2zyrerKd5gltPqkpMQxGwXE4cb
cfFDpo3Ogk/jmXgdalzq+zaggbula73+IYBtO+3B0NSu0ORJIgabliJjUAtmBczZ5nElOCW32IK2
//8WbQKJgSlI7+pWWUDvUMovCtcjXlHb7zBMQ1saglmfnbic2pNstGa9sBVAz7efhZG3LLWvj4/K
567ZLV2ZB+3O+L71SJVdeDZUnlY3/MUTFWWwKZfKOGSxD1bHIJSbiAggdcgGscxwBrM/0oxWoYZ5
9dmi8+iWRR+J+qRa1r6hwhCosEjJ9lT7rE719v9BTK/ESCpkaWg+TMFWTxm1WMzIEWIf0vzmBGS4
y/jmQQ0J2RCklAuUHJAcO3aKP288PGN/rpqRP3FniLMDSOOqTmbaHQr73tsVr/jQtxo2oY/b3SbK
wkE/5/JmIHl0QzkfZLYqCqw7BK1EHScMTajjyYpV+kXj+PlwDIs+rgQEIAxJsBzKJ7RBEOm6NNdo
agEYpPVVB6v//rD3t7QLbEeVNippUrZxrIoBto8HTZUHI2eN34uxYNLge9kbdfB+Xz2gDVKgCK6b
lwa1J7Rcez7AfJ6lxE3f0RpK8N5NaSEanznr+2aIDeOmlY4FQ6w9Y6bkiv6dA2ZGs6Ri6CPB+3eL
rr+t3NGT8pz1HhdmSuJnnCiJxvMaLIIjJ21/09F5OIysx22IgCHNsHJ81APgwwlHXK7aMFrA8SPM
ywXY6d14i+0BQ5Ij9fKMlfYfET2w1saak3Ljr+HDWoNhJgvBcqFv67pBbJoIxCnsddV+X2Ts7WPu
yk0JBWoiEEbwdKCcPlgy6uP6AGLzwYbLt20J4xj9/9OmErP06CVR2kODHDy63lQ9gedIK/YglvWx
wnY0am5skwLFVUw3I3R3HpldeUmji8rLTyMPuve471tqoOfRSRWikw9/x2ALTmi07W117H6nb2Wt
qyCzZhRxPyX6Hd81gzJY2dCfkXtKQH0+bpFhDOqkgYh8IxhNGKiUfqZqM15KUgcH/UVeDpmWjwwX
MaFvn4CLoWp9382G5kDidd4Vs/svBuDy5CrReMT8cMSf7mKPPSClH+KihrCGDr7MJS7mjbvI9UM8
VwSLN8vwQ4JIj03ySd9f/Td6n/orkr/guQZ/ZrbkNZUo0iNC637kBeEyAAGzJuj569b5veyf4/Xm
M224a29YO4UiTjJe8/nY3P8zAsYO35TgAdD9xXXwCr6HDdedCNvp0BGm0zQSOhiVumHtLXTgWWGX
DWERPSmezXqnlndVpESA7fodhgMNK4qhkff4kWq1LOFgth32HjJaHisemOO08v6/sfJ5pnUURhKq
OlTWPOAPVevEtp7PNlwbjFMD3pEdok/woe5+r/b45wYTw9RGzfrYlWqbUl7hSBcljCfNdKRaxypM
pn0nO0sDn1cVCe8WfSWfhq7CKUcg841Ya1BGeSr38nCnUWjIWsnb2kW7h1Zi7ZSsi7Qw/cI6miBr
LvunAn48sSIymoKOeIjMrtqL89LkBVHQbRRe5uft/g0Tf0ksYxEulIWOtwXwuardPMSdeWcu+YcZ
LsnRX8jFeVfN/HCm4nNI5rYujDSOIbRESUmpGdgS8Etwr7BQQWqu0aYfzm6cc3gOb9nWtSxsMXJ3
r1WG/fgznzHr7n1Ghjg4gZbrsDhtHpqqMDqDRlWmAXU84WkyNs2giWUKuTx/1K67hVF1LIyNXj5+
kuRna7t8T6Qr5h148XUsAPMUe/np9H8knrbhGo4fXXyRZCmymL02Pe9l/JUw3Nj1xTrHvzMyRDk7
plSYNT8m8TSNpSGdjFSpsS4zK3+WqnNY8DVRbRmoIBmvqDm4zeJSLYrQkI1zsBovgn809Fa+nuNH
7+ipgFhPJusnQJIocZrljU5y9dCFtK66qXEW3I5ZK6EaKah9LGLGx01OiT9x0eYkqz1wY7FNI/R5
xLcvwJr8vx7ncgiUGnGGRNQvZjdMXbaHnyZzFtyuaTjJAL+L4t6/U9u9LOgsMc2wKd93/h07+djg
SQhgvcpoEH8FawHiSkzYvDBZTCQ6lbpaWkA595BCBABNgK5eGbVubaODnZp/1a9if8AXufGXRHvY
xM7v/YKwNP1Oiwt14hW6cq/p9rR6f4RbK6CVJ+zxt/Xs6hqe5Ux4RMYGqLaYm/2OwvuC1Y9IXaSe
Nh4uitZEqlXQdRY+BN8uQ5hytGo5freO1B6mz4Rq1Vi+NtVdfscSjFW50JAGX+NxbPtiPhW12ICA
FhSbdex1fPDtUyc3lkXBl/Vdb8g86ZV6+GpId3ljjRToHKpKkl7rHvZEUALlZp/HJVcjuARBVPpi
sToBlOS60qBzJaCuyBc7H8DNxRgtd0ccP4jpwc0h7Wwb4nFKowKuecYaMrERn/sN5ujrQbAsrkhb
5vTCPw7a2CGFIgpetekWgJZkqubZSWsGf4yG3djePuQeN/1hfn30E3GuWrMZk7rc/NgMXLi6oK2S
6Zv4tArvQSAr2wrX++igRpZlZks78PkMSkUhtXw+z/bSo5npeJlom9jPFw8gz6mBg9Hs/4ALk716
EdRqpWXq+sTUUvnAxspYtF/S2gmJ5W1JkhaGl+4fpF+HypYCtdPQibB8KtEuc/yW9JQdEW9+phRV
uy2QlBixBm8KzdKKoY3EBbI7NsCy3iOFd4H3K0zcC91cLDw4VqIc4Ci2SudCVr1Kt8LZsoUXZVtk
4dFco3ECs0RpEzdpWC04tEC5QJiXl+Y3V6ng9ta0RFxnkRBjCp1FqzIkJYIektmqqZK3kT/8m5ID
cVgQTSRUzkX59HwbOAtYCG03pUmy+katMkkrSm96BViVZnW72nNfEN4RMvQBTSgIcBslPMeDFjK6
102D23zLRG7budVi4JoCGn1/CJUgmlM1eL9ZwRxmgUIQ6D31SsUQx5VIQW5tI2bSe3vY1FH2gukV
WbOkE+MxjLx5wH1VGfYqndwRmdElnOkRbrRFfoWSdr6SdrAlFWCopCrswuryHAC7ivdtufijrEE9
4l4+pGrrWmJV2ZI2Vhgl5PBokN+GaGfemWpUCYZUrETzxjKuXJYaC7LR9iSrRTRZW03Ho3ii7aq8
MJhFt1yvWdydLz06Jm+DV7mLdRWN+CtezFzcA71V2M1EWQyXLNZjT+nvbmZvNxBqxeE03eVN9K+k
y/XU7aT59m3RrcqpNI1FmSiARQH7SXq8MCi/U2LUvN04O9fMgonnI7H0StnbVQUmOYSReGfrM/tB
dI5r3b7YQbYC6VsWMTvLBiQ50i78mZVFlMypMXak4N6hjlIGCDRMF6cNXFursnwS/VhlgsFyLvdB
ZNp8ptgOO5fro8c2orsgXJKfq1+z3DsacD2J/yRSCn0SvhUx6870dg1GAWJHhHll7BKHSsSuylso
OP8eAPSNIrbF5JY/UImHJGziQplvBVmtl1AAiEIiPW8W574K1Hc4utmgbNdbTvRyf4OkOKXNhrX4
T0hq0rBn1Bbj08V745DUZmvclEvC5PMHDV9bFwcEZKDV8VyiDnuvLEukpxJBcUhLQfi61N9q0aZd
SUImaRloVvB+2vFaOC5X5/krI2MCv2rFYv/bhCWwFv3VzP8tM6mOmdlmsne36UevLdSyvg20xgT7
RUYDlpg3BXD8pUtkaCqoNHGWORGjqPxE4oeJHcBwvUPTy+m1WQBzU8D5qBnGMZYbpYya+EazI/qT
zi1EtHfQJQRbW91WLbFGrPIcIS2jmmdZa8TC8CngZGZMqz2xEdwpyamlg9rHU0pZnLd2GwTSMG2K
9o+WA5mHMzQuSB4K9pDpouI3dkh7+sTh82or9wCVdznF9XZ0uMGqwMRy0ps3BatE6+D7s4zX9G2w
caWmGeDxc+s6G+Boz4VkQx8R1ugJiYOHoqelhyArAHI522HIAY3/pDPJFFGfnDIaicbX7RUxwQS6
Rkv+fn4ZRuTVNkO/qfEJK+VP1E/XIHNAlMJRoqGdqH/rMA10zAbJ+WKWC1h7vZmqlpuqRieTr6ak
Fo6b6KMOFcgjx4oavkwSMahK6ZQLthkhyOrULg9743bRauzFSKpdSaBEDv8q+4A2VLnrypLK2szQ
zL062vac1MZ1nQkasqptY9ASoNy4SVinSxhdzwsoHCH2bADZRHCcMvS8jQe41vt2DDSh42iESFab
oj63BLVzlcmBu3HDqsvJofBhNpiazvnlBezO38ROsbMyiZhqFMsJA9esv67qf9XXxVdMO8m/4Jqv
TiGeHyOhSiUK3X8OpSjHa0uiLWnf+HK37+tSjdFDvxwCVlQgTok2FwTtcQBokhUNfF3T9zQjAXOy
gAPIbenKMgvMrLO3U9e/prVN6C6ai8/KS+EkEq+G+ipziCdLWsMWG9uTUSQUAOjNZbSOxExLT0/1
SuyTxHbpr/YsV5IKASvgwPIvkJULE6K1J2vV0zXrZpjqX2IYeNRqvyrJRF63H5a6U9da7OkjG35q
806I3dxx0x8B+zCTlkd3IdsOryUFihDSBpd0w0pRCDvLd2dVEfO3DRwTeco0P67RERFePFL7EYab
lWCOqPTBk/ijFR91kqAFoRpIGfMS19qarD0RHoru3pBTDYryOQDPKYqjBLLDSp6Zbp1A/Eha1Mn9
XakRX+8atHYa/oOaYs/PUB/7zY4ROLTRvA4bEX2vhwrGs6vY+EWTwHwgbfJVwZxeHFZO3c15i/uy
0Y+nkvkWKlxaDJPpPhBFkOwdxv5pqeTTE0zSlj1eUBwF5X46HGV5/P/55B/deJfsX+bXXIt5/It/
ea/EklXaT6KuuHl4I7ldaXoV+vz1Njz4BNo+/qbDeMxO8i4FI9FJQ4hdHBefa4UlNkWFqvvXaBwd
+PW8bKtwHCovpn0GHIQqd4pymKHKGRSFivDCc8JkcrZe5HFnw98CqWvT1pTiyQ68i1EWLTxOJVom
9/w7nbXVC4LBxPROErymjOYNTkBo7iz7rStktVXr5NTz318L76hc//RFyeIJOi+7t0cZtxLOlhgN
c4iR2CybZSZZkQR8qW5xBJ9lq6fmVHqXkma6fGYiExs5rGB5CJ+Falzlph5edj0H73vwhGvp1O9g
ILsqtrH32VONh+3QI/9MJ2THvw6Zw4fBlOW7+KIe1uVZy9izQ4qZCCAYL0OhI3h1sqwPQChQRIUR
4UKW0nl6kx02kGKE11cqtfEF/t6QQ3U0nTt33ua0yh6sgLR6jSIUDR1HTG4VFmj87p2/aI+m7ojs
fcMKeFFu9vGaAuJ20uig7bVYd09wYv9N1fJHN4af2UuhsbZYf/87a+7EGOrh+gkNOb7hAXXHTrzv
/ivbuLnog/mcChHI98uQ1vDIUZ6tUJiEP4dOsXZEzRbyrcqqYOlJU0YSrhvfj5hgpVuR2d9Pm7CS
cAer8RxHhZJdJoagwJK0C44xiw/P0FYyttszp4lRCKq4HAxYqJuU08npdrrCjLCnsdSJTbPEoaY0
b7+FjeTWV11e4H+f9P15CuPVfHJ9pRYbmc1Y2ONkcZ8PiSYlQSx6e+Fe08PXnGea/eNqaIzs8iYE
HnVNWgi8jK9hNEUflX3PAhUJ6agCzluYkUVDe+J/iCuZJtZchBzdgPN+kp4mQfyHosANivcI2HyC
SwLphCU9EkCtjAuGYHFK+NsCr9W5NjT9B/zgm7epkJ63TasJjUYdopC5EPq45cQfEC6HygmliGIV
l57CQpM/y3ckIdp3SuhNO8c50J36nxRujLlJWujFZosPyy9pUp+FvgehV3DoZqq605SaqUAELJ3O
G+FE2uJ11PUsic5dQIzkUP8rRHK+PCsuXZ+3Bbxlqtdle7fC+tn9BHyE0212lgvcL1tDdAONk65m
MBwFIZ4I2BUuk1iEgA5lBsfobEHuQI72wZzZst2Pa8hi+w3JF1SvdWYPxhtn0x6BZXOOx+ib3eMI
S/CATnFDultxqoknLjWahY8M0NfiTCMV6vF4YjOUQYo8Zqbd1nFYm/JDjWuOJ4KevpLjMinbfY90
G5/0N5LlkQ6TQk/EVGuYIyVFt29fIkr8uhGmgnLcwB7h/d4McYPkHy34LhvsDjMr5wlJI8TBicPe
5OlVFceZqmT8wZ+S+iHCn1vNc+PW6gsMdMba6lsChK24ED+2LYh3i0uRQTt0PmJDaA6W89bO59yA
BFQo4NYJufCUYeUEqqBATN5psc3RogoK1hDdzIaIx6eHfa/YGsGn/H6mrdDkrylcHUZkZ297FTrk
LlCccZDYmM7/JYaiabZpuYYanVWlPrZl0foOkvJCf/CnJai4xzh2suauLOSn18mDrTaJt21E8E/g
+GdpjO2tqPEhkb0rN00j1AHqw41DSgZpxVLXT7iseQ27bzIiG/ZOMq8aVgek4uSByp0/vlATvXWw
oQEcVooDjd+UcX44JUi9vjW9fY6wvFpdDz0hoNQIKXw45KATO98RKVEG2czg94nnUkp9ciGnOA5Y
dMhXXNSWLeA6WPLOV5wVxIZku7hnUVdvRc0Sv3O25d+ko63JAAolW7g9Myb7eKhgd85fV+chYfty
2RLNmfoAp55xC/w2GyseUGsbq2ztZsgfpq0z/OZgqR2gdozHR2A5MQiI8k3GksJcm1cHxSr98bzK
biyoolmxJiyIjBpjMYwaKp+z7sPM/n5E4JhwsxFfJa8bkSVh+zYX0j10XJJTMOzFMbic/xriSiYk
c/xS2TRWXWUW0akT98Ibv2qJ1MrcRuyxbHcDz1gaooAyfZPOLtVT/XqbA3PiN1ASilFSuEWnuQkW
edt5UefETzlpeEmjND2ySwJpFnaC8/UvlauLtgOBJQuoNNmnp9b5AOCjpOMGM1ms1ZDqk7vixn5M
2lpzT/4U4+WvGN3FnRpRiTY6a9KkFRH1tl3/okCLzzKDBhnqq+ZxB6yTb28LUEnmFfit7Iw6KPHw
Dz1Z0oyW+OaDRnmpos3jXAO+VG3X59K59hRnlgxAeVOE+pDtbfB25eBn/VJDorV3h57nsANCbuI0
01gIK9IxhE6FcG+1mDmO2JgFQOjU8EIb24TCPtnd0ExIfGABFuIZuUKSArOb4bXbVN76wTMiZmy8
BKunlU/6u3J2wI1Pk6pvwM/fQpYfpiMo/OTYNzRwhHhi/I7NrG+18t8XRrMHtTq8zJJIJHZhvzJj
HSYPACPJMvCD0hMJ+nryQe/LCuJ2xQyB90IJh7Qc1o/tfpo3OcwBy5UB5qKlN/91nXRSTdwQXKie
DsqcQnQjSX9Dw+x/lov7vk0rG6YjVpa6Qq9dYXBbUiu44N1JbaHoz9OOqG4p/8E6t1Tgp4RboAIi
8Djrp4c1sJMKo8nyMkK/Shmr8pstrEgwNQtL1/O9wxa+x9UQRwS7sHH/CuG/RMHDm/D31XFzrZwj
lz6MZ4q48wTsn+Nmop1x4Uw++WaPjuTMMqSmaJ1vLQhsSoTe8yilKY87R2lbYCVkeqc26eSxU4o/
WASyftB2J9Bk+3QTHc6NdCShN+f+9jOVqOJV5aeRJMlmYwD55bBM/v/maXp8mDXp2JDFjcLarkf7
GNtuvlgaZDKBi/YBU/Q6xuXkjIbMrwEwYRSTSuTakwOPgkGcCiqxgt8Lo/WL+lQ9u4L2uikvIUPS
YJ3iCFSceatcMB8m62WzuG1EZK+UaGW/agXY5i9orFgceex1nJiFq9AaKmivfpq+XwGYrDkikgFN
+rPXN8W9VLYCF1D+bvQy9vWOi7uAVmyOLFhgN5Xy2ostcx0e40Zg31vuOfTtycWkYHHrTxJ1qWCw
njgjSTMnD/ay3tJ+cKmuEhG6kYuJqm8qZdFMyLrUkDIEJqtQMiqzhuEo6iYSieSZCVtjPC2beADE
CXuCGFMd0zw8HYmi3reOcJHG2s8NUwkO+nTmN98c0vd1U+TngkD6r0ZzbX5I4thlbNoo0qtRLGIZ
TWdDnvVSf2ysIiSkGSPt/3VmWDgQcesue4tqtcrnEEzfM6qNxEuwkipBRsI7q7C6Y/afQP2spHMO
1qgrbaOHN4cMUbbE8ArInNRXAduAElB73JBKHhoNxwY3PwH5FfUwyVzJTKoGLTxWxW2/6fF/vit/
wsi8tigqK/QnBKZb1PlQySIrq7AOfJAeOrXsYJ2Uch6P6dJ/AHRGuOvmpsA2TEibCkV35VkaRBX1
jh+5i8wRST2nL+cK75Uijs3e3sSaB6uidI4zwDvH5xnVYWy0VEMt+IKa9IU3NqPYV8X52NnbUgJV
bZnmqBXhZekt07sPcpS+cD56mFQLvXypdiybrBJwGUJzEmtlG7gbegE/dw/fyXWt34Xq8bQTh8n3
oEQGa2XIr0DELZIECvbZ2znxJNELfmW+4VGOW555wOWG3JJs3sSt20ADZh98sPEyk8dARmEUKsmg
I8fJJnjFEm9x/hhUsmLCiNQ9de1CDRjIb8KdkKxYBOBFV77nq5dX1thX8/HL/HBbEqT5YYGx+e8h
I49lF543vGzaIhbFIgECXMkaMLV9QJX3gcti3GuXydmQ3clyG6OVhSp24DGEEeVNaxdqwPNC8QmH
k1+Gl10kP5bCvn61wzbEDnthtdiiQF/9NJmvj30zU1VURyaZHXkZL446O+CY5eCafr8BKWTk6bum
kRqx2WzQUBdRkh6zGTGsuhEJOfrRQGIrIS1yBh8R3IPBerwIC16A+C/KFK4c7qubN+Faq0eCpK2K
26mA6RP2zA5QNvs60snXkYkWxI+0j4Cdk+TADIynPApr8WQxOCJWdXgNk9ywm/BYaDU6hxlIHOWt
SV6rP/ixm5Ki9wPRwYQegds/M+RKbVGdSf279whYUw2/STGNi3YLIUhziQGoKeo8MkHIWgvwKoy4
HgMXcrpNZiY6I4kLMNZ6la/8SRNZcW4Goy2btShABjN0Xghiz7QkX/prcvEvsPvB1u3vhpCSEN7q
+MUV3STl9vE2TyJYz1iF9lCT6qcF3kx0fTLqcMZfebZeYSNdsUlEOShmv6gDRUxm0bRLG1iQslxq
FYWWN4BA0a9BizrHd5SILCksjq2WfMFOd09O8P5rCbZbS5/VcF2UU13/yK+A6wy2TBC+COa8FjjS
qVcSpeQo3PK1cQYyYTf+NYFDEVdMHDWz0Z4jmP0rzxq6w46ohr3dOTGdtafFTxqsSZzEmeb8qVWF
j/hDJULkGedGAC37VCtffjNmpw1NSuMrAU7jH9N/RAHbJRHgkooIMuWIx/hNhM9aQvSFk9AIn/jl
tXhj8GTDjf58t6Yt/OrJ9RXUD80Nyh/S9umpYaopAM6nJ6EG+HfiGYcJK5dfwXOm6ZdDksQ4KVBC
dzx5JjByY2aCUMZKSz5XQqxSi7jgOoh9D/0oUEvH6Z1poHv0OhwTlhOT26kOu/PR457igsfbODjk
el27qqKO9oNgXHq2jwEt3GV2gzxo61y24Z0jIQk4fr43UfSdBWUAInzqDkGNt24glsNzm6Cl1lVC
iHvZrh6HPrDJwCqZoZ2i0FSz1TkwazJr8KSOS7CLleA77I4dKX8V95bXDBLltEPUdhTuHKwDjzVt
+lGgd2+q18FxcuhtCfY2f8CMPyEfMMo1jIIS0yROlYeQ2lkntLJ9h/lESCPbqeYikSpqMRCMLvXh
XbJ7TVhBDxY7Kmu//kUCeQLW8vuPzMWHK9nYPnpioP4Z3icm6RWINHzhgCokIu3CwLkvZHTjWXbQ
0OytvfM+rzx7q39SWEKbklgZ2WJAWu7dPDSlcAcEral3GjBqmtTP8Nwk412WyuVlg/xY4GToUkku
czxpOJQ7BDi+IwoBQ+BgfGzjw1UvyAypOh6oMz9uIX/W75Q9lZ9MCwuElIK3LoP6CM8oGzBNhyw5
EQjfsClfVhb8EmZt8sQ5vJNktWkXKe5gK2rMR3r2zLenttnf9awJC9Jq6ztWpvlHt53SneiJ86+g
hYTbDDgb5jt4rsLrXyaqyusYjdsK3UeWAHm4sXqoGkoC0jInfbG+tRVaYyZnCzlmGid12M1VPU3y
dm9R2/sK+FEzFYSA0XmSTJvvIQOYXhK80LkU48V8TZBEtYdyq6zf48ChGQN1rRxZOYfuB62Bc5mE
/AbHtNOADC0YtgBeiD7HvxYS8K3UiL5+qy0I+qlwmb238Hmct7IiKOgl7N6Wt+UE2vZj3jAdsXQI
91hdF/sjQiRoNRcNCNbAdfnf01RXD9EatNbPkhqIbtuXuqx7/AWx0tepaukliC+L4NEEiRnGG15M
F7LiAhmHyjASGK+OpkR5RGVPmehEmY8R2ttrGbgslGDxD2dqnIrncXa610KzBjp0Pf3plN8gWXWk
hTqpcXIjhJdn1rvjiPHO+QqTl45ESg2AQFav+EsyEJIIS4++BY/zeWuwM69AgnJQ/DBLH49BCAq4
vuU6wfEVpuyT7mkaS+S8fqP9oWG7v0GRluX2ocS5eg7kwzTKFiaIPetrO7SD7HbVUMi1UHn/sPkZ
WM8MxnVn9c/ZStxn9l4at+x3VRiIEtn2r88xjvy9wlSY4eTRFmm4pq51vYIvqBpYbkXU2pNOpTOl
0h5o5FQWuDuTI3yHfJUK2JzfqvWxhL91tkM1cY8LqZZICHmZcPS/EKgPq9hEYbpxfPLDMM/VqiUv
d/vdaYpnLbaaY26q4g9m6knZSSz9UCdTzPFA5NzyTpCJ/EJ/tU5RmFOAa9pCiHpnS0/8nG+2rNK+
AK/fBihw0pZQshLd7Xp8PrTrQTsivC92omCcG/M6OV7WAbeirdVUCUGjLyUF3Qpu0upmOGmI+3Q5
K4abWmKbPcpa2mscsErtqJ94Eqk2+i4/RqjlzxbHIWP9kW69rT+J20kUS3wxX08cVln8wHjeANwP
68IWGN5JBCObTNwjzWD8ZJRxN01ojx8mCD/Mr4Qn6J91oRJOdrQtrY769o3B+y3Tcx46Xpvt2R0e
yXck/u+UggPtqXNq+RYzqjH6HyYDJ58eZwAn+/D72n4XxhXdzTm3JhBdQsW5v/dzP44aGS99151y
VKpX6Vy1FfPoD7mTQ0xcr89xS0nY0lqnESvpk64yJRCDRZexHPQ0Evcaqwhh3vvBnY0LagofXckl
iwlXgNJkdF3GCSjYIlJI5n1OVh75Egox54y/+QYmBb7icQ7fT6S/AmBeS9ft4VhJP6SkgRRNgULG
Kxjhh67hAk+KNaVtUOgC36LnP81qL7CHsCLM3RwsHi0OxEd5LaaEaLQHtQeK1UKsLBN9ri/ogd4E
KkPBDTgN1GFnBat/kFFNjql8RxhCaUmuHVVV2anRBQUGGMZf0gMpWJO5U1NcEZA0qankcdFqe39a
ZhoxVODBCU/kZ68fWu1HXfsiIWF97FT8q8eUQYP1TDZoP6FS7EzAc9iOZatXythv11vq6p0RzDHB
2TfqvXxe18Wj5gmNf75F54HCprVwKk90XxDlnopRyoRzaWdPOQax9iDYC0l4Ussw0hOtxEbXHtLF
T47+mABDs4lAbiKdNtoSQNiaV2Wax2qN4Ra+lV3qf/hLxAnewnTAl0Wwpc0xeZZ06SF8/ZpYCpRo
lbVMSaDiShA45cvpczPdTxOLAqDsCQiPcos06dh3fBoQQgaWhyBx8BcHHLF1xcU6DpTbvdqQsm2X
WasK799RNHrF2+qo/QbPasamtolF+LUZT2MneY8FlA6JhnuiCdafF5BM07yQJTkALWIi4zYG+zNU
Ys0873YNzH3OJDrm0cbxGhQybFV6S7/l2yVdkXVGtlKBviEn9rrrHXAjhxDenM7tufEfdAXzAecT
IjkTvG4SLZShb5Q0ijTK3zpq66bjH/5PY5x+SmmGj6Oqt7zr+wa3+EpLl7AP9iPUvAFmzZaI9EUI
6eescgncdylqSUWDWrPLHHB5xZGU5ui+6xt0Qj+2iOHoik5bL5bDn9ea/BnLgBNP8sXZYvyt+S4e
BeJijfy3TF6k3+h3+me5mGQdOwkUOAlAK8Rqf/4sIUdP3bsR1TwtWM5ostv2YkXb/3hQW2JXKpVn
liMf4ZKMMK35q0e8L2QydN3aVaGCFpyCe+dgsbHzcwKS/AXzrkifIRCkbtlkN8J1fyfaLUus3Pp/
sRnvelYyMFQXJgL/8yeRL8skZQZWBdsfFRx3UvbRvatU6Zh0NbgLM5UWyRwyYGJuO7b+P4X9pYeH
iO8UfS69HC2YsW1vF8QC77ghk8gl8zvLrLsLDFce5zs7g9fpNYVDRM5umbbVH9fpV91GMn0DaaCQ
XAZjYZuYQWFS+/IpHkpzxgmz6HVF+X9egSMqTeJa+ag0mpdeqjdVm5ZWPDlkUOFXXsD3eEIMauLs
xeZh5BYR60mdTzJq0DfPmlx6ko0b2HI4blRuhoFH4az0Pu78dsM3m5TbS28cjvazbxB8zwtU56ah
urWB+NLrMahf3MurjvBbj6LUHhIp9eRnxADf4BBsprxztOZpmrXVWIsDkvciZ04Gh8QgNqCVFJ+T
eRtemVv8OsaSKgZX6fU2tLDOc7k5E5R4lZEcFXRO5373kCWzHfE/Y3GhPGmeMrutEubZ9i0sTbBE
JgzedxaoTgr0PymWg17umNkquSM1Lym/sIS4pZcDrNTOt75LTh1o8axFq6wjz9nvCpD7SiKKPRFJ
VVl0uecfZJiJ2Ritvsb1oa9bHfGjvSMr+iinotAB1oAWyGsqdoOn7J9hNA8OMkrX6okclRdd9Udt
yyVCZhcrSCOQwJ70VC9F0MYczBoFbUYeOqZw5fJs58iEMXacPDXo91asG8GuW1qZce63amavNGV7
0D4TTDEGqCVJUSb5Zw2nj7QdO69mkhUUjHvoiviXVSj6/zUdA+0gkxw5wWWtpt8akgX+4PPWH/40
gLJzkzh1MrtDW6EGDV6dhmTY5tD+j2UvRce4IUcrVoYwrW4bpwGXtHnwejZPyOml/Hb7vvWNqbVV
qGvSAsCrtlPbPeThV/L8z+XX8VswbTvva/HS8aNmDqGCa/n3bduP9dLOmgmtYiy2bX2agru0nSvE
0HQFMb7YPyDWodCFLSn6irq9mSK2KV9ZbeM5QmDHeA8d0u+GFhvBdXLDgQMGy9OrTdYN99ygbMcA
s1neKH7CL+VzLkam71HUL22y2/gOcKiHHCNVaFdlqmVdq16GCqtQajGtuPrPMmWg4fbwKLwsm0gM
BfxS8T1ChDym72n7jJmGlJj1kv+R9dwnLW7OKvwYrnM47wKccE5W2Bz5QIK4Ywu8KDoSe+Zk1ema
3cCYTumFWfIeNjhQUFSpjHKjU4fDNOtbvK6UVLR6FUgPbWLEiVC2VoIuFk+6/MKyynWCbENknmEF
kqYEFxXk0clBELlSsfkvIbRxZmjKeqXmpXpHsCtgc1NIKrlqCds4EDCgmra+2ZHfJ95R2KdP/AFc
eUo3S017H7OF+Eb4Z6ipZuRfbvzJGWWAkbEV5ALBC5EYbVEe1tOpDbDabCQO5ooBc01pFMHDxJHZ
B6OIgCGpBG/YLBGmb83VaXgz+17UpaNRhXWPckywjOvmP1l4/8Z8AfBsHOAr/9gzk0TQxuZHqzZk
vWIK6Cngj4a0utMb/8x3rqt0AI5Nza3ClU9GoiwbiAVyJxssJ+L8GE25j45slbEmMKxBcrY2XVI9
MLoKtQYpbz6XnZVc+k5lq7cDEIYt82aCTJMYOhF11QIbgtfLGMYd3iCAlLqrUkZd+cMVcvX5eyLv
chWFIuISEwYbM0L6AVF6TY2hDblkU+J10z+LZWXRDVONnnwbAi7nR13max4M/doWGJkg7md9JoHz
pcxgqO0iYwUDRhFvK9nrQILH17My3kLplUuzJ5wMObHYLRK8ZO3xQ9ae1hbS9DSjms/JqWz6tNQ3
EoxC044LeaPn0szLUvxmshvmJAML8F5vK+ncby3Q2/Ogt5aotkIaeoRaxTdSVWedlHghGMbZS71A
bLaFYNTX21dA9xqhD9q2EgBjvn5slUvkYyZ9qI4+lWOXXjNOAYVb4iBpag0PcT/8bpJ0aHZano1V
zA/oFFlj8N2hkz/nnM2If/DOWdrxqWoboiakyx1Grm1FpNXBBzB+ZynzwlbOOBw9XDMbxfCRWf86
Pt4NQg3n6SLPx32katG2Q50aP/ZTOnw+OOyDUc9N5RUSZqNjSnK26bQUznz30vq1uwfytCCl1VaK
agwQWnKedloZam1u2mHkQVYgDPPFL7ygZDOygNA82T5/eLwzB53FrrUXVgZ5PT6tPJvdRSHRN9aA
Aiip3baOmzd5jHWxk2ucEJ4HGyjo08xFOwnDXRmFdUDqX3k6F67sCMRqFbFYRLW8vkbjX/evAuKr
Igj/yZDzQ6+IUd8fsheo9qExiM+uSDrNKWEnuzHycufASF/rw0s0n9ZXOhiwX8qrAvGNelsXJYPx
LUUxo86V1k3K7KDFMAmD8twyqveRbp2+0JVwyk0H5N9nDzgG4E54oPWLl+FBDHUwsxZuBZhCb9SR
tHHBl9gyHdZIqyHo//dlv+rXMG8+O/jeLZBJDsk5lg/AYgqfQVqd4lbl+9FJQUGpgCYYwnElStvx
SLLDISYZcnad1p2gX6yIR4vy5AjOuiZjAS3Y0PhCqpUucaqw9Ntg7PbrtxdjCFMx6eqpH5w+A9qA
3ctvUrIkrBPeXRdHlekrZGTTCi2PYpVlUXyx6zkDwr86+bYp5D+NoyGshQha3WTUwKWim6z3q1k2
y/iM4RlN1U/eCgsq97N08Dpd8YHbvfRsrkh9QyDOO9H3tmuOQzhXvlEjRPL/H68TIasDyHS2hOVk
vV9N8Sj08n3eVx1If9+Wi6ZCGAyLUW23Y+Hp7zwlIeVY9Edz9YbdaTUyrwMYT2h8TlGWM6MJWSxP
RVIW4H98zT08c6OMxkgamnG0qUr0WhjDSc9/7GLjRY+IA7TOKiDBGSJorifGqEYuR5YQPOdARTTM
o+ckNOXULmpuxfEuYHcf5xG+dnWYvF7H7tRFJs2F6u3UNk1mGt2yOzh37nSN6cq+2Qdm60rf9eor
qACDIqDnS3ZOnu+BiUXMRjsx2GNqLpe+EMpN/G8aZbzkQTDJEF8F5f7ZHu7WUYDsq4gqAG99GtJW
MfMqi6CcLdAjRLvpkoUcTJDFgOQUAhM2r9EDvqpG+zAKGcoaT4eHjtU9pGbifXpJgrm8HOtFlz6Y
eLaZX5MvF0QFj/MCBzHo892CYLoeQjkhsxKdgOyFIUHH2d977WS2bBmPyJx4HRnwlGcboNOPUsL+
pGxjoHQros2BA8n+h2BEESN/slP20JhYwbFdOJggikIeClwNK3z+Qo2BwTb81vF2znIUDEhMFI6c
6jsD+DEcA2ooX2ATtrTab4P7j+mXP3h5fMvfT3uRwDRhq2uAISB5Yhjn19PSssXJiDLdiQJ8Mc/2
tvyTJqkmkAPbPGxTJpmzaxDnERgs0xML8PgdsDJWS8Hoz59YjUnNTbf0NEMUzMzEcGQcHeYVFrSI
0YzBMmg0g519GL9blqGedZiZbFR1APb4a4kL4t4U8DUXEOXPYE/Lq+ruWfuB2QrqcxN85StppWjn
a8GwUhUzNRwLUEEchFGDLoqUKPq2BTvPxxLe1HgqnN1SV9BPqfrsHmHYx2GDKeTCjUozLggXsJLP
vpkbVv1iVPEGiWAMPmmsb2Hr+7pKiZzLYvNVbK+/DglRnzKZHwx3oalK5PyogN3NxCtsCmv0nGFN
TU0M3kOQ78/AqfqhHWaiWviMRgRN3GG1aF/glweycMgdz5VFSbizFC0ih3Ren3EiHbE48lZPh8Ak
XGsTGwxEIjaiTGwUk1rhhPYV2ZpAWxjLNQg0MEqdXYvzXGU7SisFV8VBsHFHWUurCaNtkuLm475P
PukSSQpgGYPbn0EL8Ln7YUPMv0vILmNkMf5mzZyzXVW6BbhNo32bYLvh9Q1sCDyoLfBxuhA8fKRF
ZFCfMONkI3F504inFHwBp7K5ycqqe02sp2dfyNRl48BYqJX5AzRYhkakoYwURNqqFnq/pLhpt4Yw
kCasip1LHgUKxy5ZgFVWftsbnmgqxm59SnmT98YchbRTb75nN3EssjtIz0g1+4C7pPsatLR0iQ0j
AAnrZOIAP4Yr4z7PEV9GpYicTeZK+KM+39/CgxEhhyfcurEFP+EMQ8cfAnBuEzNC5HODJlIfI7jn
eK/G5qVh+Ff5rRr/nBf3F8yJS7efM7Ip2gPuqRHxw7AsuUirQzUqUHZ/BeIwPMkZVOVhDwa+xDkf
EInt7naBL3zQA2pZ8ewSwSjjaE2FHNfJNDFhd0UuxBiUili9+NXTo3NIDzZtn9WfWi1U9IbAfmIa
u57zRZfSz1JuzlSpkLDK9QIrd6jIyiNfCK23hh5tZ5vpWLmEFCAIXGjsq920ltLE7NGbTJ1WMzGN
1XHxlE5wpKyExiYmBsgPDUfPd6WzcSMNBBbRQlL2iyVHEWWLSYApbssHUidxR5lob3t2+3Qmc92d
38bEbQVhjtFjkg7CHhei1drlc4j44swCG8nBtOsFCxRESuYyaHdsXfKyzQVMmVO9dna8K3MRf9o8
oI7lw/opTDsw945EdhTS8xJ6nxpgh8VYv4CAy0faIBHcedoVYBD5Bd8s+Lj0hM5FXCucsVE4gygg
G4yMAaOdJTxfGZ6I5HnAcbjuNfxEqdiBtppKFWMWZG+wLAjJc5DXMRYa8jSVDTg4/9ZXeZpk28U6
ptPWf1C9/MWB3TDlaskCCpntGGvf0NsfKeFWQREC2rzWx/kcoC4Pudu/OzQ28/ifd570OXDrpnjc
Uh50gfxY04tb52YaydibRvZY558p1sdCE7Psv0vjvjSpKwLLyG59tCvOeT2XPYgo3UASmcNtqllj
nQVr6VUocAiEpKAgvZsmsAncmmDoSBYY2eCy6nClH0woKLvQoeU4UsEcISH3vlPFe6FIRRC8YJ86
3syJ2WNxWHU2lj8SDJzAXgjFA2NAaMWiBtgqz7b05LHVYW5TDvUgz1gSqN3yv37OE2La5ZKhHLJL
JRjtR3FptqYcHLoRj73IKPDVLqrUYLDHyGWI5haLiwoRVSRoB74cm6b53xFz6661AYGU19JnqBVU
vaEPe472oy2tRKSYd3o4STEFhw3GM5z5l2HofmPn8Rwml3ZXFDdq4FBVvRu6uvSGVpa1yGvxhD+D
nwA/HCdHKa8Tt8mGRBfuicU6mkQFKnNXdf9Xd0hcZfFyfSj0Yzpk69PPdWU7ZmaX3KyRvgEGqjlZ
D8FJgH8L5UDiqJXVhuv32ZvlPrfIcGQHuH9g/YqrfATSLUZfiInEgN50wMEp1872HlK1Rl3QEYjg
eEXm2ponLIsQi1Nk/cHtLmtKPCLVHAEIygaNK9mXfNUWgauZEfQZ7nsmwgB/BVsrk6MixEUQzbur
GS8pp2sB2oE0383gNZmFQllg0bcB2clV2a1x/iHXzznNn6hQcZe3pxA7QBTn2fpgO/W9tJPNQCe/
YGRK/Dx1Xgqtpyw3NscL6nYZrpB/TGCi+kBccUA5GvoYHRfgciSlZ5bL8cvPLxzFmdWFr0ImkEo3
KbY9oOZwWtPgNOIfUPKLfC1SGlbCVem3uchX5ZGpyzbTqRjBuEZM50PHjrM81ZRvO3A0BQOEtA2c
QgSBWLZZ+PYFcPj+VyNWXhiUnUEbw0yGXA71Rpx0aNtWH7NlJhNJ/FpTHMaGbhQdxTVQbV7ug7lI
Ed5HpbssJqNPZi+azJ6TubVqunRwJMW6YPWQc2w/mbb21hlgajz7V1Q1/75ePuCz2On6mTH6IEJe
Wuafn8ugUcadbVGaty/XWY+/6M3U7utxb9UX6iQ4Z2jlHeTKzhf0AeH7nfjR9GXIWh/lIr2bkd6+
aP/ZHIdt/dXetJDn1vFN7o16IDyOKnQYn5jOTxABWbpNKflXN76lJWHuF10TyLZB+YLeBJob+Pq2
YVHSz+ie9bXpsdUMMfKGMXNCBAZkqJh1TsDqg64u/To0iG+1SRzXC5RwqyBG+AlIcKl95/2V843j
5OWZMQoF53hv1hxcSRWPEt0XBIX0h/lvX305D0hat1QducrB9Yr6P8PgJOiWexS1Kvl+nLpNa00G
/riNgOAevvtsn+XcWPnslCFi4mxDepq1f5aLPh9Xv8cLTMbxI7KCATHaEV9lK7Wa5kgGrnVyrln1
6l94dqOkb+A7ercznzHhh3AFg2/hdsNNwq9URYbWe9G/IfQcEyu0zvRhT5tCDZRtyUfOiMLQUpz5
oXmpetzU1GviZ3NhD+miFeKWNFGwjxyoaqaDg2AdQ+xuRzL2StdXZg4Xy9uR/3SdY0CjzMmaogft
VSQyMuPOLlH+evp7+9iGMO7DjKVUBa/4q1P8EA7XNxzl5Pqdb7do+AOgTA614VfTrDOIyVt/FNIw
cyxuUAODsjLV0ayiFkDPyg/Fo/YogTP1Y3pPj0H+Mj/ETx4eDX39llgLqPKsylmHPsq/eiCu67PD
Ntj7sVCc3i35xCYJuiTMP4MAicYcIK2vrIhFr0QUeVJlMmKrGOA4a8EsWlQ8OZ8C0XAHRkKAj5zZ
lwDrXK/guwfv2lNfuqOzm9SjDKxf8mSNLJ2I5ygYBV/y5HzzXqpy8ysi/7W8R7QZjCkdffcPLfZK
8/1VEewB0ALy37RrEmiFzJ20B0YV2SyuwB/ik6R4bMQaPjVvZdRFb4wHEm54uaRGldp1/Diu6fJ4
5aHMhp3yeBZSdOcVuWEAG1hzeVbycVLgxIWzZSB8nfHU4LxEPV6/I06p2JQOPhfSyYLxk+GKtmGJ
N/5nGENHF8maYlRFNrIXtJinpsz3mgVGu8RV8UTK3c4YfUIRwhSh73kSba5zxsho2WWfd39GlKtE
1E7rhbNhxIuUpb4XQbY8nqaRhTJVyiAy6OEjiKmXoS7DrTOpdaC6PU9STVE1cW9rCS/nZGUARtRc
8YXErIYuLO5AftZJVlb9JfYrUa9Q2FEwDGWgIPY4Dul7ByPl6pwTsd8+FkzDJAXriOnEBxYCgZ8n
XfvpULJAXGk1SkOmC26A9bhqHsgDGyjAIFnsZ6QqgLLmcQZlOjoG6sG6efssaJ3aiGGrNW7aC73p
yz5G9MEk2gsReflQ52MK2p8bdY37bumylAC5BmYsRFV04UCT8wUILz9Ap7I73Yo3nfbMMSvlS1RV
2RIXgJtNePoNx79UqKFWpwilZITtURVB4LA76VfUP0rzdBIlwEnJYQwBbPMFNnnrmuN+lzzwC37C
ENN7Euevd/H8NFwjjwv2tUHMZzYLYFK0qSpEFbOxutelbIb+i5MFgt2dPchGEZJGDh7WulXlz3bY
2u/OfDsVh5avcRcXapp96uJkxUuBaBj1ZM4WfoYAJ43b2zWrA1C916Vm+/HaKM6iyvXH/S/yiRz6
4ym89Rre1h8nLXV/IxUk+ysnNdeFoamZe2KvXVLIV7XzRLOiQ5jA8X8jSFZUFrLvGKhNaKu23ieA
ehp9kAh3XTPLWhZJuOwiC+pjUt1uQT9QMcEU6B/f6EsGm74oLyxL3CMEouGsCP2L5uHehsXEKwZt
UWnq3RrB4icFPURD1xlqYEwa1ElMHaeWdzhlTcxpFKQ3jMfnkO/9QuUfvOjveK1Qu7n3wlG+dN+t
66l0vdglBj1zm4YjV9SzwXUZScTTfwBoBx+IAM1rJ1KwWPWf5vixQaGwf2km5kG3+DeMuRMrmCc+
3FpWQ3dp60hNqoVRvUFeLh/4Z8a5zRAE+r+QnktH6JRVIAK5oTL8tqxVW8+vnzkRvALdK/eCg4mC
ITp1gaBrfcwXe9FTDoMBmSAYb00q3d4Wf3YJS5tbmBb8y+YLqzzPatxWFojDbPwh+XEiv39161fY
D20URB6z5xO5kM1o8TQI/jjX7cCWa8iJ78GmjV6awvqi1xlD3dBx74/RCunf0Yax1yj+spx+ylGR
W/QFr3kl7VGZ3IFYQKRJY6XiH8KGqbtd13mY0nSuagfsxpj5Fj8Pviqg9eu2pJCqsOeULIM5gbZP
PLQCHzTzHGDNrV6hGpZPnlmG/i8DL3IgzeVZ9+vLFIBGqSSxjqsvYOUKNykQ1GMVtPNdpzQPVGjk
sJox84ET3Bt4PDxEEg0GaKbGPHnYr1XjBWQ50f6FyoW81i2c8DA8FXwEPfJUTTzXE52a1CuGYrmo
LURtFHAjeifeBJgWvIJV5EmkGxa/+un61ag3nsxmSkPY9CeqsedgyzeCJa5H6SzXtEFX5Io9wJGa
IRMqL/ZoWD9a3pHJGsSXbmr305VH2dfYy7dYn6Wupes3eCg0JUFPpB+lR+re2e1LQbKR1Zr0FQlB
c/tRifq+EFPf61yWaFdTgneyABfhMUOofNU29n8cUv/NfdJMsN9jFJkysR7Nksbi2GCtcs4wppFH
PaoWwfgdWHHtjY49y282KKqZk6A5Yf0PSzUu2S6M38hbnON0dwql0IM7+OpMCC9h0oz5hxGeD9So
Wv0lYTrvbp+dpe1BT5XJfiZDOGFtRDtn8RB+ozF6ZNtrTxsb5jkFulP1xiCSP19urqeInk2Ib6pC
TQQmKwsKQAMF8gfEqb9xoLFeFuSmBVj3Na0E2JyBm++kquKYRWvbg6kOIzS8nuzDD95C1GL5zeBO
IbB8ccbKgA5yYGY9yV4m9NC5rzKw3I9ZC3krPdmzDGWODsZu6enHNRcYd/PlzFMsBzpOrrI/wPX1
aFlYbAQ6vuetor2zjhkQ1hM6xBVqEn+rDXn/Sk+QLl95xCSwb8KjmC1kZZedaNPzP96PwVCN4gw2
pLzar8CyHg9BCBHJf1z4TkmdgFGA3LxqqdLSsFuP8JVNmsQaj4knZFOF95I5Nq3qLE6954Xa2Agg
lch8HAcUsJAx87en7Q8/3I7cjJbF4KGot+GZU7DWSQ81bEiTb12nXfSLnMZcEA22SMirSr/nmGrr
XDTJ6vyZHhLiZ99aBvztsOGWdcHc0v7/wzWTVkaF3lt7HhlEuutO2ESLqRYK+S2OIjEOxx5CtpmX
fPQP7MQwwnOkMLybDlksNNG0oas17Gm520K4q14xmg+jrT7pAb/7BwG8mb10GJZB7807O/OmmgCq
o56+sKgX61SIJAZoKvYe20e/02ELo507J6ACgknaR3NioXAdohJ545e4jey4wFP/m+KANf1o0HvG
IZwO7AzpN1o3m0S2FhrvqN1kaz7XruKnB4zIJFL+IM3/cCVwZ1Ppm0V/g4abDlGy/WpVejjAyNwB
5ujqkS6teJhqvQUaF9LCnq3VkklgAB4lvM/Pv2h+2qMWsgnqnA1dkA51tuWaJ/U/ZLCYOYnPxjI6
b+H5pTZIGoOYYJ/wBE4zepRzyKClXVRy2WTU+s8AUqOy51QQSKATSn1rhYqXwVb1K1cIgL1Zr3C0
MDyZTN3LLFJdL61+8IqFJMNsyiLsoAg3cnNZg8uTNhCH8BpYp/iBcfYfXRfNkwBee8nn5yZ7JM65
T6HuwZDiTgdh21RO2tQHhWJy5mTXd3TyqPg6C3ZF7uJxLyp1YEHgwdNsCyLRLMaXQpayWfBrC+T+
fdY8WLt2/y3cpdm8Bb6AOOxPZgcBBJK4adw1l2/P4AjPQQncF6OK5EGSCBfTbWMqmjG4f+S10fHo
0EAzajyENlugrf7a8v3yoi/2C78YtdWPKCen5Taa+yEdYXh71Xf6D6GgeiOibiTkUrg7yFw06BOe
wFhtUypmomO2OaQwJ17kEf70sPRB1W+EURjegMzTHU77vxxJHCm9YO/AyGGUTHu78eFIhfe+N6tD
WjuhxknyAG4oE9SvjA/yYF+tSocHVgtt1NZ85lcePeYJzF4S0nHOkO5d6m/YMSCwEUbXmdtGh3Nl
7T6AWP0CBEbZ6Gc5kTRidEikkdbX3AG9/AhrYudzDIgbRXKGkh5E4EN+AB+6f6A4kFD8f0jA+nID
K0Iia0yYiTQQ+6uxzPNfYaXYRU8aVcis63t+pLSk4aV1+oEaqO04CjYbuxLk9C0Ggc+W9r8f2F6P
paMj+mHVSg2LjZ6vXnsGhRT6pQgo8w7Atd4mx04GzHsj1sQQOW7a3/oNQ28mjn4vANLcz0S82WSF
5gzojODUYy43gsIpKbU/qELoJWXC/TJ7tmReKAdQ6vXEWn7KWGb0CT/Grf541JZvPncMD6tEs7uQ
L1GUTl0yb4PFxIwdAbORNuosBoEikT4Iqa1JRr/BBVt+DeDr90EhnjKVPDoW0KEav0RjvpRyASZ5
Ldy/+mmMXakx19qyCnjOMwagYR6wjHOOEckacbqS4wncNIzrEAYjsKSBLyclddKECfDDJVEgdzfI
IzdQtWaoN6Ut0Qf5cs4XeapIvK/5ml+Efj79/Dz3FrnYdy558IAsTnLG6lOmXLrHr5S03btxXJXk
h1Q6ohUBtT22LPBTgXw+zSA+6f8ERt39yJGMIwzc0D0vK7Bz3oUeb9cVHliYPq2aVR7XIc1UOLJt
AupCQyNc+t2Mgpq4Q7AcwikRrJR0Mm0vCMbvU9HCsZXhvrR3yZ3qrcy/VyTrNQRsFp2fH1yZ05eU
KEeMBWsCjdrD5Mq9TrdUMVMB2ZKkEmd/kyAPWq88MhYIAy3IsX8UB+1KWsa8gYGPWeb9rGWUuiU4
gag2u5Dn39BCoYffaIgi3cCkwq14l8CBIthKWo2UX7qChXyUJqyodbnb1sqpSi+VazPQrzp6MT5b
DMUbMno9Ta8v8v8dW8+NWIBRUxPWUWk5j+nntiLSzdZtMxsP41EsELum8bvFvgc8ida4pZLeDv7v
CbS7EpbbFCxDsKvnS2mQ35nXYVFUvWMzOAK/DeYVuXbKT6hEx5YJpMtBheVXR9un+10fjZWwiGBo
KiMhDVGuvRwopkygRnLkGGdThJWiG+lpV2cXOeSqtIqvkI4GSihp9+IKn0KM2mxh/YX8DLJuzp/K
fe1TqLdSjBQU9l1Cfi+AfXGdWkyLKgY+dMS6GESbGOY0rR9pW/QUkVjooJybHq8BQsNgV1xaePcK
LH/K5cxQmp2A/q+YuVmGF9i8H64B6799JAD9j9r7abesgvPYcsOubBRnZbcAd2FEsZlicW1Xi2Rc
vmTHVov8e0s7VOEGmB98ZTsXNG1uimyUZikPLLJ2bxjB2DQwEhefrcJ6bqve2/C26kdaG3Hs6TbX
3HKtUBlefbUlcvHcV57ZtXZAS7EjTIYePsdXVb8ks/IkA5z58hpFV9VR3pwTKaGupqcRe4M8/YrW
kH8OrXTRaJ/2B5GXmFT9y7sqMbJiijv307hIWPbElyOYOkq1dM1ACvcIu4EjAYtNu7Nj/d8UsGKC
4NkjJ6ZO6G2e1BylGIAZzYu0ypvuAq/xpYYBxPMTdpRGkJ5fYO71+MPbcudAj4XUjkcrBGy4vEcL
+Y4I4FO01o8kAbSlhlIwjS2RS3UYt1jOUT+vChKqFJqdPfkNPwV4kCAQEGsk7g3Dnjc5AAK/JWHb
JVKYkP70qNMggOoh+5BHjX3uybHmIK7LdHmn/4X1cSB7jv1kwEH6/VaMqbVQF4FKHhnsLLPGKkCf
xthz0UNaLJr1Cjzc3RHcSBuDL07gIt7Vlrk6QoEfZyeFBCK6fRrY+ZCCjfJUNfkSoRSOOUiXYrt8
qUYAqDn4z4ms1z6gFjOfZLpshRWxN67G84TUGEA8fz/n+gS2wrI+mbytb/lK5bbPQ6A0eliDupry
1h/1L3QB0tZqyZijt9FGa9mMt4Ai9Ss0bosygF2PDzyTxa2EoX/8gztlGPTOaTfkaChphwxXdmNv
TQmZ5+QGwCzdDrWTL9OWqs7ZedTrOhdhS9IMU7V/6pm1DkYhvat3ySNpM1wezSkfunKMpY+uqMwl
3zI9KYUFes5KlfyhUeTk7ri7hF+q3uXISKRY98deH9FgdyBBvZ5X1dnGyJkHuEcPA+1QYqkyjJTN
yoECvtW3p9l5WmE3KZHfW9iU5dmy6Ma5aYFQIcE7xKIPlkT80rLqk161z7QljeQQQmjygK2Fa77a
C8FwOAGUzeNr9qj9Xiy8wn669OHJpCBFwVywLNHh1iqAkbtHYmFImVajygOIJYOf0apGT6OO3ttb
6fsDQ09XmqVp6HJUYHhpJVFAhJyyZjKqfTkEpa6hnoYgMQ35Z6Qppt0h3At+JY/7dXoCER7ggpHL
kw1NA2C0CWe1XTknAxfPqWIBLB6MYGinjcbwpQh3NRB/Nej00Fo+fAHS6MdPyyaRtED/ysRCUWrQ
RtSoNmK2FW3rArkhFvknw8L0j8JLvq8kvTKX9B4RVklQdN8tPRW3qiAICG3GJi5j1rpJpgmmkyl5
sb8y6cdP5pPMQZdHNNzZO0mrK7Wd3o09FWywdxg6/QisrnI7bFRo28kNFfiPlDlXKBajPJCccgLD
1vkYjdSPmlvihIYVxWByJE06/3aI4b6vI1DSg4PpRx3B+1BBJi4wON33FKT6ZYNdKps/8RDaMStk
lXDOGkh5ngWM+RYDO+AuV7KTOlVyfONYsb78ckMupei4TNHmD74IEmVebfOf5FzwNPl5UeW+OSO+
EFSk24CJvT6MYdFgzaD265l8j8UCBeKdg6QvwPxCQUZ6pcqP12i9Pgxl4FYOyV4+Tf6+nWiqTUiN
UC5h0smhUG/TkAJ+vF2YKtvrQoXdEDMxTp82mdDkamj6qiB9Zw6egaQ4ZYtJPxpLezxaEUfeeAlw
HnCM2tN1koDswb4+vQjH/L4C4UGWHMhy+jKCHqAZsKNj1Cy44xXC6qhQY9zakpU7MOX/2Tv/ZYge
hFv6eDzhXlvRjY/zxUdStlC9aYWnJt773zNu11i5hjNr2Gzth7L9ZIiqSuknyTLx+HDCnBQ7PfYD
5yGMLG6QAa5VvQTyrqCMJOpyGxhvOIIKNLAuOrvfKlAF9QSy9KJR36bjaNSn+1wscXGKCiGNY3Jw
ZwDzkF8wxWH/+ZznhMBs9x1fwH8SadRX1ijbbeDNabIPbc9fQIoh8y7o97EDhLnYM0JCC2GQyePQ
hl1EC36/OiwsR/H8rWWy0QrdOlaN/JyizTBMLDI5I6oyI+DutS5v9KfRvH0vFh56smej+vxwGRmG
XQdRxEmbUsIDb21GfR419MWHK1vXVLJ2QKeuy6zJw6B0YFkFZ07QnkiznBJCWlFXY/IlZWfN4dHY
OlK+B72K2ZO4jbPBMquAbtxOBslqAdyEl1D4gqVcOKc2immwZkVjz5kXt/n6Ws5aBtTYbCWomSx2
NYmSpFHUAziC+Mm5rbowSo8aSxNE5ecMG25BcA+OqdlArd3LuMKfrzQHFsxDrOuNzp13ehhqz0C7
6JqnZpYnGQvU1a+VhnyBpwbVpC+YdpMQZnzFm4ODH8WGWZOT1XFSEToTdkL86ON+xXWR/334tEHR
xbIUHe3MRA7HLyN6SWHyDjjXjIARMBTvwFN3/YFmYc1XnKdSimlYnj3utKZqKuLVSzzm/kmUKFUW
0Y/eBqkIYNMGtDXc5AWh84HSl7JDHEkQrh82T+t39GOPbfbEzYseo4KmLc0TBWGl3t0ZGR6vCw3d
MjEL3nn6TWa2YhO48oA2pchekstVqF6FIWhYxC4vZ5JGUAftbG8+pBY9iUl42f9+YPTW6E4U9j59
jrB99tErixTvGhdx5Bj+Kp+ZU26lNxvfg83+64Tjj7OFCLm8cMVa5LoSomG8GC8Fk8zwkDfIn4v/
LQ3+1MmV8ESSplCJY+Xz8Qke42V16aCh/mD+zEVojipL53u1ryTVONXd331NjuMEBJkzGTNpZ3yA
C3bSzlQvCwsZXPsfQg7dSpJ+uaDH7CF5Nm9J1QypKxxzKld/oXQInqpRFu9ELfBfDVPS6zf2dvOR
EqJXa/7hhOm+iTV6dvTMUqq2WETSmzJxMjOQp4dr63grEyq3/Uy4t2hObwCJ3eRtDrC/IhqGbqBb
UKzn7R2NHl6E3vUFGcHYLeSXyUl1j2Pmw8iQxZZseHJ96k2X1xmBQQ0uy08W+tTzC02MilpA4eUy
thUpD3MG1+jT7d2hstTvxua0clt+goA/PPyA4JXmBbO/di4+cALnwR8P7gJOW9iUNuCnweMYQ8Qj
fuZ0i7rVjk0aS1HPPFZ/CbIr5yDFY2kxuMovwNTDRTci9qRGYv5n8hvHtn8set7L80oD8RKedpnU
7YEusgKCvgZn3hEYw1hmH0VpBxWhSupcNPY+pAPB9YrVVtBsNZSRcXRBHWa4sbSKAZDBDvLQ1zMK
b08xYski3AjvFCGOc3nj5fsdcw6OkXpDsBVbTAIS3Tf67VBBBCIxj/Go5KdcDxFS58kZGpKJ5LWA
3IbDVvONO++zKm4sAhryioYZBMKxRmHZnOgKy7yCiOJRX9jT+d5Kyvk3DNm/q9Q/K/0QsFvowKQz
xG909WOlWwzxJjqIoL9Fl2BBkW3UpGpHgVO3ch0yKXOplAdmSJhSMJpXIfFbgv+6CEdN+izuIydw
dxnMNwHQhb29EkSNSJ27hAkQUBILMnT4jW76b9PFyWPM9g1z+rjbmhBnkLwijjMuycpzDaCkIZFr
5WPRvEKw+YE+N9ULR3DWHJGosmHWy7yTVS/Z9TUpYBJ4oKMWbZWXrwTB2uktgrixnfLIksMghsdX
fgTRflGbxN8Dwq+y8tEgulCfSKty4FA+N/U8tFPNVkzpmX+b45wRzM0mRpCxr0yxkELtcGNjQGoX
xHx+jwqikkxbuagCwiQDLVQypQL+uSL4SS5xTAz1SVI6UFzLEL0wa6bJG6qrvzKjiJ+LOc+n2TG5
+W3JQ009tHhL1NQdk5wptlY9jgbgtPAiUhmPUk1EDZ4DEfDE6698qahw8ix2N3dcbcNowUtIw1U+
E/JAaUZxP1LbBzm6riqV12dBBzSSKp6/8yoWUyFbKYlqm2Rl2c6p+Ges/slALX5quseRiDnFMobS
STcaiPl0Yh7BIPJp9BXFFSJUhW+n0WFiaFtyiAIm0Ccq88t/3Z9SJd1+FgwH2R/Qn8tz9idVANZp
Uz6uwi/eUZROG4WzrWbdSsrG2tlm6G1gn7g2N0D81TK5IGw5faKLfxjwFXFjJ+GMJ5UcQ9CNCX+O
wmXM2enGG+va0mw6cPxQAl3PxBQOTVsC12xz05/sDgxcX+RJEtXfyhDvvHN5Yw6j3lxbYaEsXSCR
RdyDrvb9QowaftYHTJZ4ZtKwBhHE+bV68KUR7J2CnmB31Rg0matFMOfZNmR7rhcSbKMAyNEE5jzN
cIsfXhH+nYzl9QwRwEgZaEBrrdhK+VIEyB5IDtAfoQAqgHBCbz5h9eq32IVQCBCwXq0euQXZl9B0
25ng8N71P8Tbgb9nlkh/uHjeJrNFus21SAMVLwEm1SGHvg22bv/q8gxvlrneaqX/3GoOMXfA75Fv
2+SlvDDNRWi+McZYfNLYLlWG0I+kNC+ZtZkkACYF5oiQPH8VQ+ZQyH3ShnZASDrwQ61w0yT4GEyf
bm/a4MZL1pXtNHSRQ6uI9KcXpDdDshdt9aGwRWOGicTM5Dq/t1KHAwj0qqMnppemgujhnUOvXW2F
kkjmnw1blgZQXZrbG8B5ibg3gs/sLW5XLX9mmB91cFBVuyKV/v+8yivM9h+PKsN1AgVxw9acv/zn
h/WA7uELcTwgHsOWl+FwEoVF3vpEOGxdprFfki5pcyuQ9HE7SJ8M+TOp8iEJz++0K9uWt13YdnuI
nRpcjB8bx0DFpE0HEEkrF9baB6pLUiJAqmUTJIfzPMhu6NLPKdHD2/Qr6SzUEiqmc+UaHdU2MZtW
qNjvLC4D2FTEk4j77AY+R7KSLTAceyAARok2JWMvLeqv8MTdwJs3ntj4/Xd35wP5MSVJeW9ZlnPF
5YQx0ipPvo5O17lehppAeGFQx2iviFOxnTCcWYfhMoFKPIeCeKgYg/2+RQz9qTraIZLSDAjAWv3M
q5hFovcC+8+EqZMM3dM8kq+ehKYujCX34b7Fnp7xyHV/ovSVFU1G0ZgBe0EBth5C0IwM6cyXgpaC
Odg15thxLvt/CmGfS4Or5WzIsx11m1sjbjzF+CezSF6yYLt20GpQwt0oiFHjsEVJ/EU8nz0XEgjf
pw+Y3R6nH+WYWAhjBedNFueS//hjnFtUDW+ElEBRT2F8/ACPrqTEIv+l+ASLX95lKl8ClZAQWUzS
KLx/MbZGW4og6M4Vpx4dDnKIs5+XJRGnSRcamOA2b6VwyBtxuE0Az9xPhRfBhC2PA30L0udt/p1m
yiqrT4LxZ4eHk3dafFgveaBn+C8flWI41NKqM/+mLLOL5dSnfEvuP8ZRZUrBHR/SQNMz0noQzt51
KeZnEgbRdshLLvkC/1RLV77BLoaEkqJGvUgpa6OKBVwKhie9eiUsVh5gTALzZU8fwnKTrSlsdvdP
zP95RthXCVsV66E48L0qgqep8ZEsGhTwjsoii8HcYt4XUzD+XjlnkRlQihaS9T0j8kjzVxl8405U
zwcFQ0xc7VVw+c7nNeyWmykXRHHsbW8L5n+uXr9qVMmu2MHYoTQfSawnbBdavWr4TtsdNgAjkHIq
bAKsj0Euxu3rSb525LvlOnnhUr+4bjNMloPj+fEvC/2mfecY9xaF/ntCGHkoIu2fHLPBTgR+OUP4
Vb6JpqApeokFo46+cxOOQMm32gZWJWFgBRB1QMwG8Ixr55nhQWQNPrRSsMGQDF6SA/iZaJRDb462
LSTJpQvuvVQfcljEiKjsefqdiPVvnfMTu+5ODWqYAIYPGiwbs1lRUeqIv93GM1D9p2LaLgZ+ryJm
m0yzSxqslF2DTvHut4/B6qJXzTRAJO5mAArvADjscdNa77xRtOBQ1G0xkESJ6zcjLCRLm1xWHVHU
ZyYoY4XKyg/jJSotx0OswOmU12dxN8fjDBT2ypUVGSU1u2AG3NGbRijxwW5gCVlIJYA5GwN5gcEH
Ics1DnRmVaRUKQprh6cfybX9CWDI9tlC66/fm8bOedkJpVE7SdrEJg6JeAGFfXUs7QckbyRW/+xw
J+PDrACUbdT/tATiK9X19ITmRoAZB/fxeIlNrv8xQAIUtX85TBqc/e7OuGwYbytmWos99GoBT4kp
i44PB8ZQw3xKP6D3Pidhevoa/mnNf9hwrhnacAf5yLWGfSsH/nBKJcCPhXXp5hZDoDmRY5SeJ1hK
cw0XRlj2F+8dBYo3Q0w1Ec9kO14rz3ehsNHGgRKKM3YV3Yng2w2erGBGAjIjlPIZLUjFok2S8jd+
xkgBMCQ0nYgiRKTCriklbSsXjEljVYdURE7je+R9gmd0QwRgKpTh5aNC1HM792kswBs7MfSbmhAo
/rMRZVZwd8ydwLuUQPeb4EFOHzdeIuTrGKWDq2w1kEB7mfT+GLDKieXo00Z3fAjyB31oEVHgxong
UzIuMP1IWFHAteMLHDiQR1MV+R4RO93MbmiQlxRRzQ/qGOhcauBpmUYV6IE9uEtxUOyWoFUiUSu5
xslzo3nCQ9x3ZbaUFQi0q02arK8pLOAvD4FRDhj+39jc0WD4Lxn+doVUr7Wg5+6Bbj78JMSwCsHY
6i/0FjKQ9zFnAMd2KMU8KmNueNpwjN6cCgDnb62PN+9utpd/S6jdJ69uGxVnK8eh/xvvGdjzWIwE
TAreF5lR2Hku4ATxvuiFjG0hA3eYMU9pxtru/+Tp204so2vWvhduj0cv0KaYohpMrGy9mmQwJPmc
JQfKHZIc3tpoJVcxhAIRIP07PqNhVKk6e2AmVNUuylTKax7ZZYreOxRHTTIhepZdAEQm/6Dg5cxX
TFdY+zlRJLl6Zzh3wo9cqJG1CejaLGeGgjIcXbIvo6Yaw0bR36wT8a6TPLoOHsry9H0Ge+ypBPQW
bLLXamPEEl5PUwNLE9XATZaa2jCUaxW7mX7P8H5zGIf6pq3hT/30T0ujXbNlbtxPhd6xm8RyPb6L
fFxSnGeWgNHVNSM7RG2l7VO9mKUnuH8Jka1kyIXlYdiPUEyT/UY5q12suA0nf5Rm2OBZFPzWPFu7
gM306Ijan0U1cbrL8dzcyuwAE77f1bZ9Wc75YscqR4kPOczuBvVi9nu78+AT8STZOmOULhSgb5S+
R2LEJ056Cb5EnMmIdpKjY3yfHDy2l3Dwo/waO77u7FEQMqrNk+Z4jv+cirkg9pMIVYS53077gpIY
/x+de0N/N1mpEAVnyaWMnOd2ujl0MK8mSl483mI4BjVZpl6VrNSWfhXU/HqmtNSZwjpqS8BbPitb
sUWJZKI3LYbfxTesDAV3SzGDivtvKkNAHfTtQbSZDMxLRRI59zabg4w55WOvw0vEGvvYsUlQ4EBy
VBQXEOXtgDGqnviEQFGxcm5pRoXM9cyaRGhCrtRguwHuaK+pK38HUM/Qsk2pEU40zoJeMDEVpE4I
Mad5Po72Hs+Rj+CMhpJsOyL6MjlzRWvd3T8ucneTUQc3YAmUrHsJt3XEZo9y8HtYYiAbAuKDiQTz
QFmrJwoQECCm/ZGE4jeSDJsrL7DgFmr69Zm5On2UnoFG+49w1+Loh8LPTFg5mBBYvO4BCEwFwVkK
5m0Wdu0XQriPnyxbD3P/AmNw8XWSsTRPNFqz93Ra/EYEraZcHS3wQtq0SIBKUBZozOHTeeK7bpQ+
KpTvMFNznbJq6dUi25JAgDQE1LLbzh7YaX/9X2fKPhn/CA03FNryrnOamXD4GxtzqgoIXegjlZaY
gfAUxI8hYV8boRD957FbP37jVZHuTmo2Pn0/dTb05Inixn5oyxyi86vL4OFSKc2bXBSUQMZEsEqC
118zW1IWDGtgNV3hN4RwZPlSve1zn4NZsiAWI8riqmHO69rW9zsXagREpIE8Jlz4NMHD7QSJxJNY
yRRhdmxqfPvGfBccFqr4084pSr9JB8h5pC1tJ1LgOje2ouWEjToJNKsnzoXHAcgkPOMNJfTeTNOf
sc69vhF0WJaf9HsVreZqSU+FowjwoVOaPQQcv2hlvkkt2zHSDWHeFAOmTVP36w9QyDxdOA1aTrfM
Libr7XoSRm7n8BiOena8YKnzhc+yWBql7IjEGby0Mfe20ytBiL4ox5X5RcoEGacMMSdh6T+11LcG
If/zMcILGxzA6vkVKRNBHfN06uLpOCtCvyI0xVTiDMFT8i+1rkh1AvFIBk+Zk67+gW7l6uEXYJMY
bs/ZJq9ZkBkFOwHQKPT4WEWqDil21/sNmhVydrNUSOiormmqudkEiYT6Nuiw+4tio80YkBbLdP9Z
3quCAzsF9B0qqZCP/xBWeIYS0ci3j1x9+T+j/0z4VDrdNf8Ji3fb5ESc7VvsmJlnEWD3RYWj4O5L
30fm6UmUwYDyv2fnlgF78L8lnyQZ9A6nSRX1Ss1wtmIU0VMJo2gkrm1K6vk0SBx6c0pcPk2a6pmr
c+Ca3rlm7tCK3C9czvCW1JVP+4dByWRIjDG1SpvpDh63TM/56xgY/eETDFFdMxj91DKkS3qH7+6m
W0g5RpDaXPlCZvAiM105Z2s2dCyshTo0TUNt99Hh3CRMuy1Uv2Z7dh37fYDgOZ0eKrwrA6o+l/Sp
at4DziO7EceyNABgRZQrSq3KHtFHihVre22KmkngCFWvWOuCVjATfEqYPuK0RlWfbe+sxdBMAi9v
BPTwPjEi08zXfOyfBkaQnObNbkTbAgrqeJs5VFc3seHZhl1e7s65BoOFySjYfFspwlvDdRqZ+a5o
+jDeSilkLWrk7Vn4DwR+LhLhzjbiiGbu0oGe9muyk/UQVuhTU/WaquudWIf/0oYD11cObrPDe3iv
7pAXZ5ke6Q7i0CsJoTOSCJWHjRHO153GPRzDN5DnYd4WC6WhKotelY30u7cr2ZtPmRlKNQLwQsLa
hgUBgMN81cQhzk/Q81ehEcB70qApzIVuSvf6i88dHd3VkL6u4MpHp/cDW9MT2N9BLjfNc5b1Zgix
fNwd3HvC3sDjYUZ6Fwpu8JZBv1ZqfB5xujJcLHAUGZZm+zWtv0tqOi3YSucuqXmbOuKZKWq59y/v
E0d3eYbzzluX3QqgtQBOkzOdu6SXUnL8R9ONLAzhbLatzNPWJIcTcp1yqxa7DKgDJYqsRiFd2wkZ
HzBndUVq5kjIlGRFn3+DRc5QJwR7spQLKloTYxtvbRx/ulE3mtWubTG9GVMX0xZN9fPcftZSd/WF
2HiQvEbcRsdTB6IYgpv1sOaO8um71zGY6DN9C9h1gmthA1FpOC6UlEg/tE8O37FSpOHJATE5nBgh
En5WHZzvXKjZzL5PPW+1Jt76NpKfGh5BRFlBbcXO9vzmuY3XRgJoDrHG9qNZtqHkESsZkOc/faSO
NxDuUD133Q/5Fwvn6UvNfGjVlqgmx1k0IBE8ytXJf2GzVJtMhEjQx0dxUUn+1om0gi9viNGJuEpR
bruBfgGEfwhq8ylzl+KrNUbFJzh4bD3nvRHI5uBM+dn55JGGb/Koy3NYrMvEotdj39FZV3RV60WR
0k5i8RnnbMPgnLb+kECGcPWlW3/1PdyusNVsV8UMJU+8NZQ7gIZDVrnabw52wO4KM144atmvAXjN
Cb6hsFi4PM9VtqTWnPp8YFkGaMZVNKqXhfnqWk1l9sd943bcxa6v3wK1loGVZkLn8QYeM14kaIdv
Ac/h5X69VBcZuUaZEOz8xHNAdP2tYTWbqv31hW4iVJWlHeOWBFJPNapp6p7unatKlqAv+AjyxhjA
DxR8gy6RCT2V5L5UilY5s4NQbUYtivTjAwg9/gq6KVJgh0+2nuBHIORO4b9Hqzjm/loPXTyhQ0rW
5onmjyjUbP1e6/uZtprHfyP281jVc9HNaWimnktdiE81r4uDSGbe1pj1+7jdXcN2PRiu8/yi1Kf+
fAV1sBirtpcc5/mQ7MaCBXejVojHy4RRwKPvd7jtJLXgfbXRZXsCNJLE8XExPacZhibVYd8cKBpH
eAeXeGDQ74oW16Z/2ydJ6I1QQig8av+UyC287e8Fi6Wz6iv7XMkv12DyUGo0Bpk9N7H/PlZeCjZM
9BHxLwNOtqeO02a0b/bVFNRW4JJXGuJZiNekOR29nIpibOLb0+f/YfiM8TAU0lnhBZBaw1ZBc/3T
jA2n4/B77vUEMfI/icGdPIjnnoPqmvLEuoodA4EbdhctO7p349vwNp58g2vWI/ZsF6KiM5JeJfwD
Xztf1szLUZIobIGM5ORjdJMoooSGkq+9FdA9APD+XJWu2y/6zmkMdXdzNI1zrJnfQrFShQMSR4NX
5Qq/EYlKgEpv66uzUvECbPaxjpogQFX0LEdAfmsenKMSJygGlMsODEk2d8WzA5O5e/ifGQLrC2d/
9BVrlCp/HyP0M0bINZRg+FlmHesaahxXtFSGGizhs9UXtSS37C10IV+moqT8NiIBqgltbxti9b4w
BIhVcdSTmUz/vqgu/+zNZI4dhtn59UI1qINWkywVjL+HZdW2ESNMGq6/7wHjUKGaCNb/C/P0o0+F
EorVE9D47BQmjcPA7YXbYne5rrAd07NwnWJ7UY0U9njYeUYeN2t9AX/KztZsNzX5KxmRg6vBkgzJ
SX/KYr6w3xTStg16KRV9EMCHFaLTq7yyEHGLCDWOfF8J7muzbkDKP6QQJC2grNkCDSKO6XLa5wee
TGCUdZ9IqF1OsdQyzePx0WqiwAsCqf6u34taPF517HRIucfHQre4doAYEZ3GZTLWPkGu9REQV8vn
30R1zDLS6URebyhGE5vnGclLNSUQT94AZDgTT7Va7YZCa4JkIpToAlZRBbCiUZmbZQ1t1wzhwm37
3Vm/kwWPbpPqRc3Fj0isk0Dk31thWLTpDIAn7Ye2WG3qtyWm9jfcjlL92zbpBroI2JPKEuuxlrha
BeLCeZUUq0HD9doZ8SaKTBAK6AmbpQAyNOpUoTX/XFHGAiLxs56gWVBK7TybxInNRcOR3CQCHo8o
zKZ18zi8Oq0OvdXlcPcKjLkr2EGgEIfXeRz0LIBOEpw4mjtvjGQv8LdP46TWk1XmGT/NeGPuhF5x
6KWzQwG6TcctqoZFJJ0w8h8i8FUhlyv6kqDNeItxjQ2EN3igafRqtNCEIWeJFqKkapKd+VL5tluj
qFLGVVUx/8ZIPKeNSShF0kv1OvSBULSPUcA5Xur3d3ft1pmBP2WxGnqm6jngyyDM9i4AfNxyHJtf
nmFLOuY+bH4gJQ2jEYSbKBq7pgmeEa6EFrYQDCouEKsTOyB8LWMgwDNFOKcb2ONo8BPgVTCNJ3/V
S8Jq62ExsBD3VxYT39PMUIu32DU0mEZJOp+aEvSqmyZbBhqwT9C8XfpB22e3+JmgfHI9HuwufPXf
j8BmX7bWCayQZ4tlUafhVcal4Iab54S1Jfln7OW57BMFVsfZ6VS9SfiDwimuCkdMk7nc+Sldeob5
xylE5M3co8jqbJ5BNKwFYffOwUy6pSvnb9trh3u1B0T1kfh4CLxxsUib8sWFlND00SDE/bDkHrgE
CroAN54rNzvnQGKjRFLBwoQV+JSgEE6LtJS1DWwe+6bbhDQrDRo7iqPX0bdEHKl5ZzBkRYQvdT4Y
ws/TtR9kX9u9Om+Bgj/6cTYuI8Jcq3Q1P8a8C8ejsA290AzSYRsjhgDj4Xy/HMXo3CtYHalnDOtr
7zSPS1/Tpg37xaju8OdyKxDO6X5tZFYDcSLOA9FOqEDFNiiZHpmbIaPmPAMLowx3vBTkxaa5GegB
NnkWRxbUZrz+IMTtXixUR4BfHz3HrV6VjHfQRIOqeFkBnU8QFsMJT8SjT+akengrGRg5NRk+k7L9
M+9+EW4TCqHT8RApcHEPlAe8SWbnI/ljR4RTUND0RHaJW7kpvf51qf6coK+Ktz/m7foOIgmONFkA
Oi0F0lJwjZqnhv2svH2yXwJFHhrH+z+wpui3Utm8NgmOjwXqAN8xBSbmI08Fog9rmfS5Uu081jXF
aJKbYxUSy9nMlYKvWg781rrLDP2EEbshHk5XBUhhqsnCOQaBPEMRicpJ+JdgP69UPFzrSFCKSVQj
7imIJ3btYk2sLJVvNH68LjhPYbMNSs1h8Am6dGk81ZYJxic4BDCT8V4fAcn8VOPPP3wu7n38aqmm
TgZ94yszY69S9Tb5+ZwOWPAjepYEGEENR9+FzCxguj3qmZ3SMIqcCT6VcbnTKcS2IW1cwEBGhjyO
TtmaBIivDfMnLDnQQOK6P3xgXD5LwkQu7iLyDw0MbeeJNl4rBVqwJ8aeWhNpaEu9oJcrDLgp0G42
gC6x98fgT16ELTj5Jj5jSzZjDDVZfbrUl/S3MtxR3zBYfJQD357GmsNs44nkf9Dy6bE5ak/ICXeU
T9OSbKdV69iQofR2crAwL6HiwYgwJTQ1ATflkTkgpRzL5NH5kvf/S/0IW0bpSxm7mZikKrOEp60e
7pqNqhrKFxASJtZnvwBln9uIG44SzKNk83ne6V+PiOREQLqhuQUN37uquoa8+gP7o/geKmjc/XoU
t4JjR85KccafxuFzfQ/K4RPE9hvCae6TjbDBYf3GWCZU0CXhlvRFnVtRhPcaBnq75bGRiZNdgMjt
SOyAZ/iJdccaRrqI9qHmR5WxBYkesrAlBE708RqLNftz4ejQE2hZNgjRibsInjJqGTYMhApCEFnF
Gs3Z9Cq0pNeBf1ZT5NB6TtjKanKa/MQud8gYZWjeKmotxavD1ER2Vgru4iEiTme6bsvdm8AALUzd
WJX3MlKDqVKtyHER+q/zyB53cakS9p5DrziUic2HuZlC8ghYHPJdNXnLRI5C3IKta1JSFAWD9D0a
apxdVv0ZfceLuXJso9Q5qQoTvrauVAooxhTbWrfZ+iXTuVAafeWosTVWRoA64tlFscw1PVlAw/QZ
0w/r5/Jx26RoUs69bcqaISLvJNgiHdtlirjNpZBOs2nJ4kbOUZnlTHEEWcmglXZE5W9ENtbcMLOk
Soohub/lz6pNaWlrXkbuWCXm4u1cinIz7OyLZSfDs6Rqqn6EnxeZJLTuFsfEiDdEd7QX9dTxANKf
k+6jtr23lMQ6EZNXCQHmVCO0+UONwJ4BYm5D8QgP6Y6Mdl4h443+q/ZmtfaXCHRcYobmh+PXpyP9
QO7wImBQS+9MWvQhdNmpRDfoyB7v0TU3a2SZ2K8zEUhxXFkEeo7lCPX6Hoh/m7zg/fx50SQIO5F+
UpZFTpv9SjJWMYkYsLhSBozPQLUIwzf4PNrmGlAmi7+3dcoY1qlIxWka5BWawBT9NLMYb2KBdrc/
RGRVMxXvTWZOHNMTybd/h+zYMU9KaX8YDfUliXFhldh3CMac1MeYQvwlf3ZXEfvzFBtvbXAwfiRB
t8e9tZkxrjRGKGDo84QHM9eKtRcaOXsJDhltLBpDGPmDuOp5vM/Ny42YnJyFPlx8/BSxrHWttTJx
d8OyEhjzZ0grFNveDDoJIbjolwD/s4nDSC4HKIhtXy+cV3km/IDUrGApvQh8DsKC73XAK7fvEaTh
5Q5983RpB95G2nLOv0+6zRkNnsAoejp+eJ7fPiogauLZtLSIvlb5QI9NLOQMMSXaQqYFMJFye7eK
nIKjHTmr2scViz5CfY2U4KLYToYh/3U5rvseYxjS1+UEwm7pMP04kKoigktWNi9srR0YMHY1oz7U
IXy0/a9xy1YG0PRsUPCyK62Dmuf4TV2EE2c+a1JgaKPMsT1d6Vk6F2evss7BZ4WgZTxZA1utrB4Q
V06zxUzew5f8PIcPtPoWoj4r+2H+vxpFK64xRM5Y+QysYo2SBzWXhHki74EcJQbh/bWGi6B0/Gsx
T1b92KJLmn8aGIHIbMzTkNIIX/zjMdl8ukoFgpOqysEGW4YrUbch7PZXt9rgQClROcdwoBqKgDZo
iPWWY6rkWk/QlsjXh6FkX64r9JMXQblszQrT8OeZZQngP9j8TPp01AxxjIgxBMRNMDmHpOYqEiIa
2O5nk7n7LoR5W9YMg4324rHkRzUZEXHV3j3il4I88c9Y6EilqnNmNg+VKXf1fuflGK2VAkN6qStp
QSLJPfoEvuZkWg4sA9NQMq0Fu9dmYRPyxxav++ZXUrXxiJ/ViQ0F0inlRcMPVsQfAM/iXZgjnQ19
BF+FMvDB/uxGpfS8XOhBdoxn9weWRcYJnkTjSuZTZ1NNZVtYkoBQvyNicKzyrVgL/b4xtQP6Q1C+
9cWo5A8qDMLYYwQK22jpZ7Jt2BFHjDiyk92FsXIhaEdkgOGLCxPt3Q39A1cP8I2kjxiZssTJIUVo
8NnjFg3rk9MTPzTGn87HvlY2A73UrtILnlvcBZbNrA6JPB7NPsfxvgrSnYX2Oap0XbFnAAJuVZg/
QcPHE2Pq8MuU3TJgsqQGiEN19q4KnmNJFLfUrN6Zu36mB4SqGpjOgnGTH9HIfD2xTD+sWVSqWTE7
Yuj7NtojIlNqAbCvBQUBnW5qT2KmS44D54kZSwyTQPbKHD2zdhRHSqHl98rVSFCulQhi7GIQjY9x
MODB612wQzJoAXJU1a+KHrmUEjfwj+0WVCQ0PSja7ebJlCSSCWlBBxPfQxoCaq5h7Xob2QmlUB0P
MGO8M0b0fyF18xeA+S21yok/OPZQOYBiWMWPCTRPPXV/gcFJq602Uk8ktX+q7SoDa5v8Dsgs02AF
shRCwt9QM7VhGTlF/uNklom/DFUdu1tVzjPl5cJquxIN3/DPR5O+HFeg8ee2wBgQSkD7ek6Llgwc
ctWDjqYOJN7tOh3D35+C+jZoWiwq7hK7WFZmRO9XeEw7mP6QHRxo595QE+AOK9Y6nedJmZ+wjkR5
fBnsW8rkGtUZUs3V0CoXAR4VYGBZukwFp9WG1kyj5YCUj7yrAUcphZiPyP5tOAvWcLYTm/BNid6/
t85cLib8uWDJJUAZ5KQIwgbKtOaIcjgOMrvR5n+q80D1TSDhf0K1Tpny0p13Q3WVPRvv+/FJANSe
pNki7nKb5+0S/hpJgnLGWqEkxkGOEue7QmqTYya8dl5NHjtDrbEUXK1e7uV296nH8tlw4fHJaCdc
H3qhb8EIPMGBRK/D14PfyU5kk7r/6RB+wraGBwj3VE7QMlT4iM8ylH+fiuopijtMZxJB9EXkmn9v
ZCE2nKj3R0hBFk+0H31Ur7O3AbJoKGEBU8kVdqg5R5IqHD2aP0Sybg5toxX6ALd+9Yq0qiofFQcM
86nvdda7oDeAABEoTp/MKAkMHHGxiS9YTDr8dRMUEqzNM/pm4HLarswCcxyGezaR3rdHCr72oNDi
GrFA5BwT+qs65Cx9jmei+X2VYT0Pwr4M07uoX8tUEB7uJXtqWGm6XBcyBU53L5UbrlLjzvMNv+9b
WhXfaXRf4GTw9GiKq8Kf8pgbnqfXxn66a0icsKniCCGKM04I6iICwILfOCAsgfZw/cZuTCzC/Gqr
33WM98Pc5KH+ralS6AP07nS+Of4Dh4jeNwBtxzHsskw0ugkqCfzZuAQPkKE3Yi5mjSdtf0QmsV0o
SzTjK47X7CAzgsH1OQIaIBTBMPza+7m3KSxTd2/MrIJ5xC7aLzmRu3pcl45hxvu1Bulre+SHQIqf
3v5v/J8fIt5gnKbxtOE4nOWoNIZUciaLMQS7u9lq+zU5q5K28TfnKJ9uylLMqgDFru5Ejn9onRZb
E/7qaI+KMpPp2FvtZ8XePLp7oQb13y9mlZimFjMh/DtLBfNG7Vxw4KZeAMTufK9JP7FZWxvca9xs
jD3BkgGsaJfqw6MND6OPLcqpNlr9fKtM2EdE9PsWn6ILzW0Dzr99A7vvSHqHOiRqQ+5wbofa33Ls
83t/Q5uXQG3z6Yn7Ae+csSXhkZm1mk0T21MBSxupnU9ospxlRgmRoOE0iHuDpaZ1jGv6eQDxkmrN
Bl1Td/aRaItbT3mn7ixfBeZjBt5q+rL+hd+lfXZgasltBqofeo1MBKm5XBd80vgha2b7IwxzDbmr
zcU0e3ns8b7oKFucVbqhWUAC2HE8MY0loByRRNXXFds0mG2FbExYcf6jJ7GvjBt1TvdJO28Nvp3D
penTxaAeD1KpsxRYDLyCb3FuDHsqRUY8zk6LrirRVVCjLM37r8a7nsrUfItHi1YaP4Hrl4wqpICQ
BTbroEQK5r+RGGUNTahel2JT0SN19XSHG1dtZyXOI9qu5s2Xrj23fY1G9VRGkVjRUl5+4fO/yJbF
FLZrXZ9DN/bh5yl8z505i18RgiscKmZVF3rQ3u/rdbrVrxY3XOF64PJF3eWukKpbOLxFQqt2TsFq
6iszmVBVavAzYRMvC/KafC1JtywJednhJ4cvTOq2VqTAHStPVzOJIPFaK0XcOOizarEfQpEz1wIO
ZdeLWxaWBwxOSbnltU13RVN5vSBeRd/5hW2H8u2yjXpG8Xsgfz9cNf2DOtCtItdOFd82WI6oEhf3
ZTWDqgD/Gug2wNK/BOq6quRp/S4vpMDgztXbWBaCyHpZDohzpB//evqyKq0ONG4LKCME2oISN7y2
SC6/O7W4t2NVMH5mkvKiYEVW5iHHUrpnS/bHcx4nNyWSx2vVYeDUz1q4WTb2nII5rY+gxPUqAhNE
TGiAEueJUTk4rhX+AfaO767VN9lm3jIty+whzBTktrBayhV3DkbduMHqx7Agzzd4bbVU//Sby+as
tp2Qdj4kfcEsYLzk3kB6b22Opr4e/fqWp5VIhFyeirXE+sNDfkTD1rI4BUI9eyAJErasEfDXSjSP
wi+kKwHwkrQOmyzF31rF+1raLI5ttrMvhWUDqWcSzN4BPWgtLCjAvUkvITAza1y0zhUkvp/Wsm0l
7jEv6FZGTOx4QzZbAzCou11VJI1FpK7vbiLRrMaXzUykXuN+DuNXymDTESSgl5dGGauW+tgUUyvO
WOIpd3u5VxCH1eBCBcF6S+3yszp6h3cWRnaD6fg07MdWmwDZCuy8FwHfXd/DtxfreSbJDOgrbeZw
eXvkTn+q99XS1Ai6SHjNkX1iSNtgprCla+w7Y3WbIQ2BYFKx2kK3pYmJ8C8R/i3s9TPJwL0BNr6i
lnQzdLj6qTzrADrS/q+dA3Jp/A5Y4AxCJ+4fyDJZSQY7n44XrsQ/21oBs4mQ0dYRFvyUHSCHI40n
2vVJVlqGJ4sZG4/vfLmHykFroMw4I2W2PZHWdNu1ttG6i93JPr972MLxnkzItZ8GmR4C116HWGdt
Jw/iOC40vVN/vkZ15Wz6UVd2U4D1lx272YvkRHxKkhPk/YqZ0pFXYz9CVQjPIFy+cNU1Vzcil5SW
ubc7VBY1CGm+NH0FhEOwJEmdWIE/zZeHn61uwGAzaf8Km12eSBEgrh/r2SrtCTDWAHiFkDmNHwN+
ZpbRJJSnXw0oqR3l9xvLPHddrmXKWPHahB/c6sTpHVFg1Udlit4r9IcEY8ZnnQsx5+a4OXdIaxRq
kFYH/wb6B3j8NmaX7yiNkF56HUK7/jQVqcV3cpcaDcTV+A0hCCQrZJPYr3+hBXk6ZyLhEUNYTtcL
DxLADKkfqVO0Dl489aq1kd25v8UR6mnbr7Vg9e+Drrhq8kqgm5IHLYzfTCLs3lisf6H82yczbmcv
rnV5zgj8Pf+kGrSKxKd2cWQhhTPEqXjsrUOm7USSaarHE0EO+994jZoM7xVf9UiMfjJ2ZSvSJY4/
7ZVtJf1nifyKD9PMXvfDE8xaUndLJE08GqYFmvCSuV5yBKPHOU45pBJhq1g9HXGxYZjXEMiQkOZW
UAe/s4VibsB5Wt8pI65XB5ONxX3D15bzoJ7dqHNoccwRHYXnnHb8J7WgDI8pI83G/kytKoTpn5SL
EeTl5WfpvFZGsTPoWKrBKNpe1VDh2BUln04gn2OVYCTsBSI/UVGf94WweC0XeYqTTjn5tllueGJX
LuknUJ2sBvo2DM/Nwp9E/YeTrc6N+cfHrhzijAJxRIWSXszL+eEY9hqowHyst0C5aBPtyCxjKzui
l+LOrdCb3M/ZHevgMV0rjcJYuqPnpOQXDV5zkW8ySBiF4fRiyMmhTqKAzbm602M5xxqB0JZ4OG/n
ph8RRLOZIh6HiTcfhXA3xeodqI9tOKeQFIIzg1U1eAwpua1+kqmSw52e8y4zXf44rlDEOCNvUxzP
J8dQDIoIIfAfUfoVS0iTAyM3UnkQM3wJ5G6GNicYNMQmJU5zGofBuE5G+O3s6cd7pJqGc9JieIZR
2ry/5+BdQ0OE+xDRhAA0oD50+Z5FQTh1UOv6L+JigqYCuwh46m/BSGM+/6vfbmKV1cqWDnoABCX8
yR2kq7DPHSU+p72PDl02iNlKhWkQvdDSZaETpUT7AqyHaBJX08/sPZtkvKYPhbOqsBibnigLwzPd
e5eX765kW+tWyhgeyohkWRPjnM03NFHmk4qVE9gNe4JVP+CvdAAFFS1Z6msomWWN72tBmv1Gpkkw
AC4e2nI3Yo5n31m/5giCHkYVAINitBDOwqte0hzW+VVuj33J5lqlB30vPC6HKpIEIJ1IvqDHZM11
pxc8tfCKBbRwsCHMEVLsqBAyHU6CD9aNZzHxcQCU13as6kfACA5KT6NPHdd+0lDDxEt84RBrKMJN
dK6090DPSw3tEJcPrj5ZjAelUH58ZEkMeB8mFXjkGBpzOsUes88MbZoVM4j+dW/Fn5WFDOev8OGX
rdGs4Bq7EgYhK1YpPWV/95Ag6zDxTuMHtTaXvyEWW+1CwNuhYDQv8r47ZOSsbpeedVWM5rAiWeB8
ZmZ18HDGDsC6Za8q2yVBIgx/OeWFajpECOs2jOyZF3xYEYH5huD6OyI5T0yQZ3DwVxtKM0oQBH/s
Fj776xkAZkAAji9iTIxJXF3kHREWCLNTNbvME1YPDNjFK8yzOAVvygu0DjRroAr3AQXnS4z1Qp+Z
vDwfxsvtVmxjOzqaEluwTYEunaaIB1tLxjpeTToSwUnvDpk3eH3cBFDla82dK+QmJ7jWEXpC4pJ3
t7qyfHFdvhCE3t07bNJOE/1/+ThfYbYJXelZ8T5G92IttO8XWDqO8aQKqagViDPii0NZXTQnPJ4n
csd6EKpVLWGvo/u846qCUJZyU+4zaX4yFS9dyzlNHDGOflPRkFQYOEhufMj7sL2kTk3OSFnmp2Kf
JeXS8nPAVjfwInbY64jmLENZOsnSd9U0oG4yH+tYHd11nDdFdl9hVhiPeaGydD61ElPbv+7rnUgM
IDtK3lNAoD9SkIoPE5F0GQHBbxD6npVW2cl7OpHPlorVBG75Z5b0SvVqkrLZpVCJaVyjk2PZr70z
Wi8IWQXyWZ08MZHpLa9PGd22q7LrGZ8xcVVRUc1n+G6QD82gDhjSuybaW7rHcrXsHHGMy8LHOhXj
SUw9O6inKWiZcOuPf0ymQnRoC8BZIIOgDDxTbPPAdZJQpduWdahhOwsxvv91onsjudz/0RUmu/6S
ttmHsKBNERATunlZnEIs2X0kBh+Ko9bqp3tZ8Eal/aNmmVIEWfoHy2aM140AldeCZbaU/mEdIo/0
GD1e3c8sYxhtoqR49sdF1/P8B9dZ7JP5dFhXAld9EbRL0hbKoUzuls4X3N7bq9yxbzY41HI1OXVk
cnc+prUVGTJX+CljImV3fFoDox44YWPlLBL+4dIsrKUIwzE8b0xI9Z2wplVPQaGtwk/RLg5Ia2Bk
YMJ0FqjNDD6LXrQ2bunAIfYdVO+UCvvrIohuJxyaJTTJhJWNAIjwcbrx5qw09Psea68zDx9WD8hH
n4KCZcKOV8AmMB5EFd1Fdu5Dzm6pV63VQr5+1nfy7bw2yPR5qJ2kcDAmdAow+4ulYanWNd1icmGx
fYipi9ejCPFqUsEByG1gzp1BsPc8qra5D0LT9hRjF+ylcEdydrYKtGv6P0K27giB4E5im7Ul3BzK
DaSbLeJPGIsJFhvYZbv0ACVpfyiOr8Y7TKx+SKyGRv+8F5l4zrTuYMT3J1UkGMvg4iM8k35GkkOg
crRF7GgnOs3/B22thHxwZgHtmi9w1Huhh37LIDMHHWgkKFXWQaExKbDZfkQSX3af6IAOfie6Qjpr
noU07VOs7BfwSkEgEkt8oEmlZl4COud+Rx3g+uDQMKax7cD/s6R+sBAv5gSTUzaHfyS7nFXumsRE
tvaADIvWAI3OM8eMcqKDzPHPNesQVJ1x61lyMY5qbyvi53nFbqTYttXsOhQ6Ds8fenH6SzoDc2ir
qnpuoiFa4H0wtNM5TIAKTKAlqVWSzde4Ai90XpA7YiqkosUDUN6bizxwLWGotJbmf7gHbI36rIx7
yzJ/dO1yRTDwKVhvTQV1L69CA9plKx5dFuM7Dir8CnuMco4QyPcOc4jeKImMMYTs75e42LkaXzJx
GZuz8IW2i6+hCow0Ag9AkNekD3PGvvEpBwtuE8YIDxsbNuGbV3frLrOC8mgf02OvPCSlZGjYyD5v
VjT4KbLsoxMy3nfpBkvqWi0y5iAQWQWCx8Y9OOgvBWPR0/VFCdkLUwXyDaq/mLzvoPMPgB4Gls35
SkATlA7WO6Wmucf2HxZISIU7uyJy7Qik6awOyqDKByLGMeIPOHBgvIlLUIXHVUZOVq9hFwIeTccZ
ah0zrHctOd7jcf/w9UvAN1m9l3+jm0VUC/0IkXEBfDjxTA/ACmYvm5FMuzUcODybFtZYZdtykP1R
vC7FvGXZWXQbFa/ED8ACmOTwqM5aSGpdW1RFQ420OycdDXp3PbPhP9v0I8lDYm5F4efVRe+mEn4B
uwVZFCshNShHto52tjKl7cwiuxZS0FFMZwbirE/2wdFYvjMnCOaqLzlXUlxfVCYHCiyR9vReDxeD
Adv/4s5F5JzZcLvqkfGjasZzkeLgJQOpr4S43fPI7LyDJDMbrHmM4dp4KAQKRJVrZlhZon95b63y
rDGgF2dZzfK+RqUytYKdw20bbY4vY7XYu2ZNmfmor+dvPjyUGL3JazoPCfqh4uq4qXEzakFXFkEX
ZPvIgSAqT/typorIA6fcy7rM1bAwzbyJmL1QqGEr8GL7fBToDoROVC1dp4jsHPCwxIT6HcVr5xkk
e7SFIQz98rQDtY0+Slvw3SmmFv+RGH/l9dJChkwHFTzjUhVWSqu/ofCEXBWyAVmiaBwY8T0xq6LH
9BxATkNzqahSpFwpOc6Z3lhyKpPmeD9W/rAVUUcCAaHDeX2/4RwrJ8Fwl8y8yPeKfCScFI1Llgo+
PQJDVDH+iZ0s+mCM4XPZnyIIQ8iOjJOplntgR+t25AqJl5gcoVLZe2IB3EjuYT4JgWBQ/x7EBK8y
ICuUM7iBfvn68SrxI48pdTtHB0Hipg+Gcg19VDW99SPcKbNGm2MwsRU7pQTaqewuseuEW57LcVzc
YLT6mYeaWBsRiQ+gLZNxaU0oqWrVnebRQqqhCag/fynqsHQb7oJHp4pFucL3V5KZXXOpXx0AF4jJ
OTKVJZGg15m9+673+GbawTvlDDWPOePYf+FBb6v5pir8kwYpvOou3E12i7x1uA2Esuy21qi6++pM
S+9hh/Zqczd3OwZmOyGf/W+jLQafl00s9q9yP/+UPAUDOd6eKjFCNJrqyvdpsYX0MoAIY8K/KfDP
SL+CVoj+hx5lIrqNu4VKg6PQv/HYRP8sLymVKIeYRGVBkTswPKusXPp4dmmXr7DIL2AMKVs0VSho
zLMxnTSIGF+8xv5WTGzXtBfSTGytZ59pR8RWb6lt6ORadantRzvxQShaq8WV3nJH+VfiEzkOH3CK
E1/GkAr1xjA7eFlFP9ZwUEsAPRUwpOLWC7xTRAq37P0+Y4Z9kAwIe+jER1MuvWCdVssMxNx2cUHo
sL/QucV6Y3qeh8PyyRGlV+UdpyyqMXFuB4yhJaaZDKU9SssZOhiUa5T4Z0RDNFrqigd4+Lz+2GjV
o5btpb/0yh2WBlvVzjLzexbTdjoTzJ63q3tBRoH6/04lNJLR/xkLpYdD9/IZe9+FPhggU9J1xC0M
h1fCE1MNePzc+mmACRzg5vSL+JTEhPzRPKoboKqR8tMBRW8NxXd3S2HtVmsXcnJDzrk1BqLyFqcs
FDkEGXJkzHekBFztL77uL1atMkkbMRaPk7XFmC9e1cBT8rNNsJSTHVdDQGOhMKdlGV5JvekrVGmQ
dfGBH4srt9RZe+tiqQyU03EwKSCDDR6VQ00Uv1qSyrWn7MpnsBqJorN0ca1b4Z1yw4LrxNrdI4NG
NQFJmNF5K9m211xhne3TuIPFczqrA9NQqszIRMDzFil9ri0uSGlkXyxAOKUjuM2hy+7paBNaFXkv
lADuUeIiK/0UlwRyMwJ51Ad8uaKMfxrgk2u2T7MQw/A+PIm8EZzLU0p5eNoqtDMpf1MaXW7Um3GP
Sr8Sam9lj7ygXTuUDBOEU0tNWfcafjWxvRajXFCQWQhjnQJVIE6RuWt14mD5CX4qZTV2La8+T3Iq
EXKJOMe4UCtLHX3gAtNWiKGQ/f+7xvVe8vFwOguYC+Cey7+Xe6iVfMq5nIrQ2RXciAdq/oMzcFAc
Mh7w2MppuVoJ5BMKPHlMV54jIzXsT02wnspHlH3JWUcKOdMFjEuA8EkGWIOrq48wMzZoqS5bQumQ
0AAG4eD93nVIPw6Dc/GQZd2C4U20xlkfCbzFH++FD+1md59zfyOMELV/A5HMpp6U/EWWagOsTWOv
pCpga+n7u73OLF3Ohc+xWUSf2J3LkuZWzgLRVZ3wM1sjqdNlJWHOq6JMl0JMe/OEssJxMJ8KCoPm
fOfhcbQte9mb+bmOSzGsWh3j0sayyGySbpo+mMZWfFVSaPq/LJ5zHx9Xb4Mwo8UkiYDAQx6XbRDV
GQHZujkYNQkn4803VLn+JxVl4hPmq6pT5pmIfRCKwtU6xA0HFJAGcKAnteCyagtX+teHj/Ni7u/2
2Q2LFOG/T9+Xj5APJDU1WSs5RRhZsWGOkq6bnj64ur6N7ig6erWW8BcjBejktFlGs463LnJawAjx
B2cXgyWMlYGlMb7/8H3aqQZfvADyS9SopO0KQ8U74PCCy1e7ic3R8PPzEbbd60oVgEb+snbirWZL
s1jwc0l4WiIwQb3DdqnY8p+8zzh8j1bOmAWP4Pg9sxD4cPtxF6iDOl9v3kkEhc2Wy5MQnpis7F3r
ZDq2472rM03seMHdRECRll4/aCtNJ2Cte92iLGjco0NakfjTxJEBp4WeXWQMcZLLrEfcFAHwoPsi
7iosq9a2vW4fce6+Npmt9PXcx6QYoyRj9ajpPRKsitW4tpan+KPuPJFsd0tTBSEmyeM1g5AzxEIe
5IyZghejsp7EP9A8VI0CRmxCZJNky94jheKpRXSZJZiKMSpm88gtWuylF9dT1PFDxiYPrQWrlBmD
buP47PF733O3jFINxoVbWNO1rQCLDGU95LiqoAWJh4xA++jTUOQF2eohcdZSVfbme90hnaDVM3Vj
KAA+eZ6kYuXYsbiE84k0fDolsWlaobLBBKk1GFP1rVVdumTSjbJ+8EuuCmPf9NVQQnapsntMoWvE
2SlNErnZk6rIJ7eQzI9uq/R1Uy4BUWj+aTiIurnSQNaiY64ToWv8JeZlpKAOUjik3vlAEHNsH0Kf
eZ9/u9NyaOZ1kdAVhsUBkG6fTuOJ3R0i4SHBS7YRcLLOud7l1RrjtugqdZbDUdPymFacKpjY+iBq
d6NZrsjVJ2W1MLwDU5+vCbStnx6FlGJvEN3xPyn6VCWr5az/Bcql6uR5o1hMynsju8qunSy6I1Yo
0MFgCuR8CYmBXIBrtE9gX1k6h5a22IbhWOLXS2omYdoHHRYcdO+3gBk/dOysjkI9fgde9TWwj45j
ORy+prFpdKHH26hlrYP/pExkAu0+ESwRN/XAEmkivpzM5Aa1gPOZnhFxRGnG6nbfyh8YMtqM0oTN
RnQRRrP6FsEY4y7YPVHSZaswpGijlTUBMczoP9gTZiXTdP6sI3OmF/q3FFTQ6U4wSfmlzHbjLqaW
qel0jXBluvn4VPcTk7jS4qBHo12LbdTI5bXVSSF41slyQ2QSoWQY6Hbg3K9DbOyOPkhPSfAgJygG
ABkOsgUPS8Cidf9qmRWUGH5E60vkNiT9lKAkscrPyXgPlWxduqRmbi8PiGoQIjMQFI9dl1gmmGTJ
0Neq7xCynDs6tTF9PiGhz07RKLuUni86lHWQYrh299cEhLOj/75g0Pciky6I3bIXQg0LRKaXBP23
Rm96SjLEix0uckbqdZ4jqEOkREW9Od+kBzJwvFs5Q6zIw4llIpTraHnEcneNgup0hzrnQdlyyMu3
mvea38WrC36dBMGzkA+fyqY1Dl5CrxEOAV2PJZ9m/y29XjvEGsr+rU69+wKpe187WO6zKJMRi3yr
vzZyI+o509HfvScSWABCYm8/EkPGEL6SoSLQfn7slap44hPU55S4NIiJ4zablyAQh3ZXzX0Smroj
UXBQy5YufXqX5tn8C3uYoPu3OixiciM6sr+ghIOUI4o27kvUvDaFQAMRu4sofEMg6WUvTZqMXXp5
3uaTlFEGeUQgZnRbKQm0oguxBq26Dq8oYD7uwtF3gZSh4h7HY6tgzCv3zcY8BqCW2lnrKTeXRBGd
iE7n4+NpFA0JCjL+jdvBlbV7ur1L28yrks2LlRHKiq2AVb5VTtadxBCNXBkgBvxhknJOKdcXP1a6
BfzG43KWp/TSpUZx35gb35Tw6NvGKiJZfZ0+Gyudea/vnNzzd5goRRnC7Zp6fNI03ce4pn1+oH27
lC+lncva3y0hbSLMzayVzYiOiJ7LTCsHM2nnewhU4fZPqubcytfNd0SDsaGzm3KzgqhvDDH3CZNl
aEZ9Xb6DYUjEEbr0QRP1/XUSPEeGylxDPCzBsG2ACLGgZNbTikMyetcRym97lvoTTNOxAzXT1gte
LooGSpshlzLjKYOPlRppFvxn/cH57gK7kjj+tHE4oeL/2VhVxXnTmkbP4OXBnkmuSt5SwKCmJgC6
wvvImLJlLGVLIIeHCRslRv61RPAO+3zcJ2ZFrz1Rs2rhh/CvxnAUf+6kS4u7kssTIvIBnDN+V4H5
gFKKcoXMb+ty1r63oD3TiP3zOOkYO5W0ZM30Ys/VKWooGWpV8Af6lO/FgG78Dm0YJ1u7AadEBMDb
v1gWPxHj1c8LJCFboGTT3Q3MyL71XVxOg7qL0sJZYVfuuOtTElplAJFZRtwv8NZpAh54Axlkhuky
4PtO0uJI4vJOuAvwb35AJd6s42FyZPRHf/bgc1ol5SbyNO/AKimN8TnFpMlePr0gxogt9Maz/VyT
TVI4zsZTBr54L0SQBolkjAzTbUlyfMvs8byVuStWsWeW442fX1lyYg/PLDHMFVWdiPHn49TPviO7
775+qkwkCZf7hX+cPHlj95seKVzMwzHyvFsSd9mKnzwo89INy3RCQZT4GqOnrM5aJxd0peTqp2TM
yCqWlC9P7/POlxbWoQ+hHJjqnV7wkL2Vs63lcqMHVoVx6fj4yo64dKGvKwqD1I2KHVTQvOetexTH
rZqvjreLoZ11SpwJctF+sJbfKC5MM2D1MWA4ajXeWSEqx+Sk9/bEAt1f6EKDhyewjbsmcu87L5/F
WrULr3e/INUeCnRvp86lxezrk0i5ufasuFyjEiZWoflGOy340VNW0TPDdYLYjIS0fczNG1n0S7cO
b0DIj+AvCd/f2VmJGsDbxdxV/DMJQzyZ68CpnQDWC/uFAysl2HGlexyKCPKN51Gd03LsmjfpmMeu
HnWfIr3GoiWZW0W5cNZNlsu/FyiTnpLP0f1Vv5n0GFTWmAMPKw9R8++YeoOsIe608DW7foo0joqB
5hJqrY3cJf0vSP8GnVEkyhH8wIKVsa2SR3NbWyWQpdQFhceSfCA7GG/LUfsN4Joz2PVidLSYzjVB
jMM56QYI1A8zxYiRmXuQNG21KNojRjVbw/KZsTFwA1vPooMQrQP73kZp1oSn5dlnDC2pBX7kE0Q1
KEoB2vRfmSB5dTdJNU2GN5U4VaLAxWHpqoxlXev8DJnyI81pU5jhSa/SR/kqFAe+oCf9MxxB4e0M
LbQOzJZnquz5rRzVcBYESK3o4rmvXAU9zOulnGFmnh4+Op7MP5VAEw+iUo/Q5HmozPusj0BE46DT
xTKG//9BYwim/9+I3sktP7x+pMAWC+khWXqwLTOBLg7RWaxLe5bIaKd3eHTfH+crAeKNYBns9uGb
x1mdsxaMwkSwpR0QZzDMCD4WkIlC3/M7/c6stlH2ravxyzz3LI52BfLJ/cwCuru+lLOckZnDrtvC
reO3A8ARGoXOSKOp2ouYhmc80OR/xrgmDGdju4eThkxQ70MOdBO6mp6hCq0lQuzo9PoX14fmFbWS
75mzBUwvSHpXccOe8K84aLO+O0oqvV9PjkDj3yKSwtMkKAcu8yBNw3xOz5WG2nF9dkmXzTWUVefY
ugh0LMv1snP8y67h5yAzhUpZJ2J5kiZ96VQrEaLyJ4c1KCy/5vVj1pz+kbwKDMU4mdc1HVVuKprM
om3+FrKPtAwO/7opCMvDsTVIM/zSNuCXq98B4shctyFEu623zIoGJT5L5AVi4LIGUFfn3mLBbT5x
WIjTM9BUEKdLY7BCui8THL5f0hJyQejqriYyjMl+qEiJ8k5e9fMX4vyJbVMRFTD5X5EIZihidLXO
21tfTKvYxy2AXFksqM47NFsC+v3nbRAwKhmYIGfuZfjokN3RaOzOgk9YGodPtAuolOVWEgkGTzq3
iVERPaeItiVWkzY53JUG2ihNXkTtxTbLqQRPMLOB925PQGx4xIabxSPjMkSgeudmWrrMI/ggoJj9
ygdXl0slppqKI61+Z4A+MEV0ogJe9Qa1z3dLmhljJoDJ6t5A2hjs/9DLCLCjbXpGVIp3XGjKGnr8
hw+ATESzv25QjMl1Ci5UQ6SgsR07BEptCRv3siOg/G8isYcyCr0++AdLBRumfx54pQVh/alsJtZJ
DW5y/p3P6cJGxI72pL5nvhtr6cqO6Xrb02Bs+ssO4jvKR92gzxxykwO9X9WPEAwrt2oY77idNJzS
31XQC0ogbwB2qJ5DHglkaykqKPgUHvGiw52Oh2kI8dil0Ia780aRC3kn08Bp1/XvX2IQcDabPMQ8
9Be79tb1PXuRtVbjwB6a2rWAXbE3k/ST8k7GvfYhhj9Fnw/t2Yl2QWeAB1wW5Vf9bZTMqc2VVoqW
Na4awc8gywnVzqkXDMm9rS3SeVqsbqGsA15jtff7RldXAEKalZNitlFbHh5mErph1ww/EefNHki9
erWOPY6zLl0m0g8CawkoJQqAKGDUla+neMukiEo9uDVVSEuKVOCBhrajeuWKAPRoVDosqtOyxi/U
N5sKKArQzX1f6vK25+Ka5WepafYLL0ED3bCFLFlLonHnPBAbOFaWSdfeRb2Zb9UBP2CBw3QwkgC2
b6posIFpVwY8GlSjn5yqt2k/3b4sLE9U5xeqzFb1OeAg2GiDZbmIVYXqO/Ki49e7NW22tbZiJIYe
+AnSVTzRvnnamOjhwYJ2buuhWOtEpCEXUgXUmCIPoX/B+6KdM33OGfCFsvpGOpw5fNmD8qkD7u7X
Zfb4BrkBQqQ1EnOd8syzQc6LNnGp8A9hweQDW9M+6CJ3G64FrUrO6FRac4nHtszO4yhEte6CHA7P
nn6VUxon2XT1VQyAWQLPB/0PnUoTPfajnQF0zDIiHkjH8V5mSF+gWEWcIdiKmhwDpwSXM+VMXXxP
svnMHSh6ChLjkie0Cn3I34diOZnBzfuQJrMdSUwjq1tmgPLdaLTN3zooFqukjQTmUg04yuTlPObJ
dTrp/PPGipW4voDYGBE1wX6bPuCG6NKjgqgcrzWMZcOIdkTnC4W/MAkYUGqpe48M9vymCXFpjzwG
xdMxZXFR4KpcBL+7NSqCo16P3VY7fjO5Jnyb/KTLUUcssT2YH88L0zobGoff4XaZnlybGxXfTjKZ
LWvOBh9ZgrE7YHs31Ofc5x+mQCIEA9smYjc1Phw+QFBWg/IJwGeokTA4Yv18AX6e8UWFsISOjeCi
A9yw3D7VXSndwBhhSC+njo6UbHSv3TWIJehHrgy6MdxRCd2HbWZ9FJ11PMiXonVTN4fnLAUUyC6C
HslBsMUYg0omp4PfigW+dXU7pRq8wqgZDk9Olpcl2NXPGo7nZDU4zxSuMD+MCWNVrkjmOmczq39S
PsdPjM3XA/0fjZoKxnBHjqeB+stbVLqyt64ELQH5gFvK8hDr+MPQgBPa8RMum6jxIaOYHyaVo/pR
WggNirGg8pzug+8o5W2ogSY4wymFQ01AEUtD0OnkPCKyrfdq5qtPcHJlF7J2s6J1j7XtErX90tsd
H2e4GMKj9wtfWIJOSHQmlMCpmN2J0wuqxn5ZwaiBdg+dMXnGOexwHTcXzzv1785jzH2z+Nor1VUe
F/CxxCNAcQ4kWGxomXqAa1R8ljdYVDAt/fVqnMHEG/B6BHBhG1XYnfNvaE1AH3VBaK5u7lRZbZzV
4BZea6znITm1HItK82tPbKr+v/U6VEMzlLp+ocsZ6Xu5pj+eAqAEm91aer4R3Hk2DeSFkPRFFLip
tZY/QaweebLeP9Wa63pK8y/pbtGye2bYtmcaCCHiJv8HKxVnrL/TOZlNxtvIPPfrEmXlufkDRzZg
v/JpIdM68bRBmOWplQQ4M7yw+4jcS+lkxGZdseCE5znOpZMHGFfaK8NBIiRy9u2G8bw3tm6LQg6N
TUWneqSXrM55VQNiO7C+CLt7lmZnx8Xg2zY39Zg6Oq3CzuHeRoVsnPIspUnHRTeqIB+ZKwwOv6zA
CjUfVb+6V2NDxHarSJsV5H4usrvUF83lpL94DH7JCl8ppibx3iLBIGPU7BPCDdfV5GlcS36X0Hfz
72jzdbcjg4vbuvvAPt7i3B4VdXMYU0o//UMSZJGjejMdCfGpcscVgWropyigpDVpNMQw8JNor10U
Oj0b6Oh/6KpjM3K3ZMQT9jG8u1NucbD8TbA8PN3hyBJtQEeTQ2a1diDt9DE0LkPBWXFNVtKgPVf3
OrJ0u2VPhUj/qgKUxcJo4FJsR0hSz2FvK/D2691o2obXcACQihKEtqmw6Ses10LYwxu/wAiSGb3X
QVJr09UdGa6DwW+KhBQzPlt6h+D8j1+h2fXLA3uw7UH9wnKCPUVof6ybxTaxFjcQAkmasAPivfHj
VMwdFTsHWxH0+Q9o7mOlzfe6EdQKfGf2W74lUvuMggsOGGvJRErI5wgHM/k0WXhBr/WPrcPTT17h
hDoHD26STt26Mz962qBwKVusUM7pmyk7cr6LIrBniD+EbUB56JOzUvmzTQaqqhG04pOeK04hc4TW
J78CdCKVhEqCGIbdYzSW6HJtrWaUwDtDYmRzNZ/I73eZBWXm7+riSYuhpVoR3ukCTa2EVuWVr8Bm
PMMGo2ClkWdXEWSgyiRYAx64a2p2q3euxV2+TManj3B9j+jY5FfFZ5LuGZPlL7dJpBzpvHUfk0fN
q86C+JZHuKvCzW9HOmdKmzovEjfsdXjIFqfndllj4Zb7h6IGFMLJ+pm74UYwWh5zibD49A3xOW5E
SXRzhd881Pu439BzKIXDeDSitn568MQWjkyoBiDj+PmdPcZzA20CSi0g3/FUY/wophH2GWJzTf2O
FeKd9ymYKkY4KFaRmMSOzLzXveBCHqAEXTq0FEOEp/nRmma6bZVsUJTRzf3dlrdxm8Cy3HRxhO1U
Df/LtAfEnDrsMcTNE9xfkoDWjj2Mya7A5mMz6922KO45r0wsuBg5dFmGiABxTubtmHXG22yO0mEX
tYYVVfkuaKWB1AdPSQpzt/sXefkuNu7pMnJYUCHlao/blsiY7+khMBDZr/Xck57ou/fQ0f7TbwJm
h351zb7UDE2eJUUlxoP9CT7simRLBCAk4EQjIKyBBJwT7OdhirLMqFEsR5RVBPWOHDPg8Gc7yLpt
ALEHf6JIOvKz3sT7qj2zLeAhqtTtbHwteUtMDJIpmu2cLRdzZmi+q1EnC0+wX/qWBNhk8gTEhQ0D
pAjSr7fmLyQT6QihjGrBwrgrFZJxoPK/lNv0z6JvhjdC8U+MCVwKkuNzWGb35tg69iZf1tHUsSSJ
PXEW2dZGOFYtyNt9A5najWopUcNfhSRyDXlNfrRkqEBlp9DDQaYyY/TCsASYlrsI9NNScxl15yzx
DUr2UMQUCwduc0sNhgVlwZTsDPUUEnClkUu0egIIYSmpxI9c3GN5DLKkxhldxhP1krHUzVLZM8Cg
a+2Q8zlKIkxojSMIz6r5i25Cw/ypQ9jVOGixFh0I2fLD3P48kDajvVFodPcSEcVBxk/68uw0efCx
t2YluYpbbmm+3KkuT53l3W1/Yb6gZ9vbCT6ZYkZ1jd89z12rMhItfW+0cob9NYRxUzbnmlsVH7ve
XPE0ORh3FHN9MSBVfhVV5Vj7m923TSvklmO05x/5+jlPh7XUPsulMGnECJegiDkIaxCDoYHotXq+
ayftfMhE2dMIT+/DaSoZIb2/BZD5z3UmFqF4PIRjRwSpCM2UulJaZBli2CLW/KbBF5bqJAwDCcSM
2TTanFokFsZwnSAP5iEvzXjSOBG81C7Cdg/arlRuILZtGvd+4xnxjBexq0m3XEi31mm69mJVkVqo
/SScx2L+IBO8r7TjFp+7aWkPuy32wTa0dP1UfnW0L5FzxvUIsrpz4WCE5lq85DSGgPpR/cpisbLY
1RG5WTd7BnRWUu7o70cITjwWoWYK270fTf7p8RWhoXqP777QKOu7eHpnQ4SWWIB7+OCaO8O1gvdA
NIjyc7SRn0YTGeOZ+ovcsN+IzOzK6vIOyLJ0L/cXZ7Ic3gO7ZPWWA416Fkx28/hm4Qtl6h/iR4AT
qhrIPGVKw4Y2DkyqrTAqy72BQqxRnnHMmMBuMSGGZ9frHsSUonrmQpaJBZNmCv4PxeGO3xQTo0tb
pnot8NHVNSFzl816TQTdmd7jxYqguKQdEpJWPB7UR+Du7Dv++sSixMkocCqh1sDnMACQTKUNdPnY
Qynp7XFqNhysKeqp9pQlRd/0t6MfxAwnEhVDQ/JBB4Us1sZce7LPwQCMCixGBzabdtQpTGUFdhBL
Wpk3lH5NP+1NKCSpPonYumW1l8L2fet0I8QebvsUAcKYbIJO0SP61VSU2xrllyn9y0vAFEFxOS37
3mu16mxH2GhFzRxrkAZaWM7OfKkW5BDy/YCHOOJQQ14eB9BYvo4dxrY2QW8yyUydZ1t0S6zsm26N
X36mphXqbkxmNRgJz7PT8GKXNgfg5D9PjpfcLxTE4aunhQc02e6cHTl3FXRBRT78hF0VBdnX/9OS
INZII6WfzwLjX82IiyGUOkUFJsd3ffLb0UtG+XadyQ3px5CQFGNPKz4Kz4mwProqogjoJ5f7FMfD
JFFkUIdozIKs1Vrv3Hs8b6P1LUPefG9vOd1S2To388DOay8qsluUxDpLsWJc7RrC9Zhha9l8QGf4
7UkzbUEMqStSyN31kjxMfl9Ito3pamGco68BOyoa/UiuSDThi8jDgJvP/NPMuxLdRtk1KwM3uuJh
xBmONSlQxQkUBFLW/k/mPk9a3xHU8BAi8RCNEr6cdIH/qa5zdW5k6BHiilVhgGIL5d3Hk+mXKpng
uru/ee9/3z9NGAzIE35k55sfy7LBA8f/o31wk1jgbJa6CCKSShQLDjB1FVNLROQQ7rChZwbuWWPh
OysRjU3bNSd7+TVFV4jN2Ye8e8Hm2iwEQkYcpArRftAcHVQM6dOzk1fgAgH3KMY+vOXCgk8u6/CD
K6NJqwPL+XA0Ec3Uu1q4y12QK1CijqttTDA9VDN5nGYBft1hpgIq+dRn+D1IaW11Sc5LuFECYayB
D8Hrc6x82RdxQ9EUygevOg9eoJieEX/vEKS5jZUuWHEUVz4J6KfuM4SZjthYmQ2GUgAzWJTmBGUf
hhUxwfWpiIu/tbW8dQJKGG6xiVu72WDbfI4D7LA3poSGqNzd1axrUlcVyRqhM2NL3uCOVXCnkTQw
jTHwWBH9QNwaTc8SQ572li94vJ9am5VgK2ZYtc2sNBYH3x98o9t9JhXykMxkllL2ck+d5+j9f/0J
lz0poHMUFUpQtMeeHoaYufiBT/xc7XDEsK0TbR+YgCDIKPX9qup0NGGb1SEi+97Oqy6CzC4wiVX/
TESrWzZ2rPwMLYHBBEBxfdhy5vjMt+SCrgIRi9aJa5A37K9zbNw/WqtNmsPBhCo9vDYnIRNIYTuH
MCmzX/aSoLD0IzAi1hwMSVC4Klh9ebOpQvGd813Zu9H7szHyhOWAwKaN9rZJxW5Ft3NEK4gEimQy
PbKDv7tRU3yeb0p6LXLWSmyg0aOfUIKW+XK/zROVTlvztoRLeA4x7p1XQ0A+OJTMIzdCbZxl8+0W
+LcvyCzqU85OcIv+/xiEq2FS/4LxEMiSxpkJUs+sz7b2Ktt9l5fAETSV/PZqX1ayhtmw/VQp2qdN
yNvyFBAmHCYj40M5mYn8HVpHBBdwylYeUTc00tgXgeSNfYcbK74Fw2Xqix3E/r3l2Qn1xlAk6OZB
OK1Ojo91KvPas2V24c7y+IKvtgdmx15UaF3lqmOab2zQFKEuX/fg+gDLySCmEHDVYz2agiiCgGvD
82rgiQbQSKw8g0OQH+cPJsigmwYhBkuSYy4UPEHG2mha8AUggvn+vN14NcFvfEdzN4EbNC2Hbz3E
EIRHv19ZKGaYBTEeTO2BR6NfTPRhPeuwpsWYHqCpa0w+KnTK8+IoO1HWiqhSXHJfr2dHM6P3I/XB
wD//7qxHfG/iHYw7Xjf6Oed06/ITsRu14tGqYRDO214fg2ToteYILrObMjVhvKqxNu0M00JxnF9m
bUJp58zhAH2FnvuG4Vu3KB3ANeeo+KZRYnjz3WXOU5/kOxCBzw7eCQ1DMJ9vyV/Cj7ZfLb3sYAj1
o3zOzqZTeB3BzvlG0bFJYwIBRpe47wVuqMaJncke5/Y8M+qANRkbKNj2iThfgPHTUQ6a9PYWW7M3
SbtzhSGUH7hq2fgO/NTXiuB9AjZCjVyXMwwPbhQR7glZ5lv/9TcMiq2g4eHP1G2eKyTtJLBogjM9
x7WYpYhWPqNtRKDXyGLgEUigkW7kLuDuu9sPHy/j8b2WHn5Hwbo0RI6wgJfZawtfBzLsAoOTgl1S
JqkFucDXikp7jwVHGSjK2tZ4zYHc130CJfDnc5V8cUnJwpI/gJqcANKvQhQW/5FtZI43btXN8EpW
WQ9mS9mmtMqIj3zWZ1vx8ECuoIu5Frw4XBJ3NHYW5zTlOIQz4QlUgB9XOfJxpvzenWQpmTuMyZwD
CaAhg7x/J1drO1Z63IYvl16SZI0nVm+f051ksvb8Iaou2KqsBbs96rtUFkYnxhqIUTuJsr/a0w8H
Z9DIgPbt5FVuua1Qizmht6KJ9IU1Ubb/7DydEm1X8d6pfxUkmNUAJETDbpYA7Djqk60ppOsFOTJo
Xd4P/A3tlancG8RTIPhfTy8HQGS5e86rXR/J3gbKpq3wdUepR5WQkwvDGCAuexjHfpQ5T+zizD1U
5/aVzIAndkuCD7UT5vJv40qMR119O9BF+4m5N5bjvtWiBoCBiAPDLtEE6TFLwHSiT2PWyu5VAzyb
ldKKjI9qVaeOXRthhOQ1vmc/eeJ4LxQqRt649Qht49LaKJ6glz7Adk45pR3Df+t/foeLFtbo29Gu
LVIL25vMxCWq/6GkHCPoxBQsNfIugcK61KfNheWQn8yQDooTIICmneLk2Qi4XYePvqaFBENf+cOn
nx2rYGd6EjX/Kb+1V7oD9jqVP6eItq+LZbMtXl+Ec9ouE2HDlXAJOB4fnoCRUaGNq8YeYMBP8w47
44nR+qpuJMzdL0iAX1w+sHhraQPWGOh3rJcrbeCjADwrxJ7NaapwfGn7VMwyhuLUpp0UcLpVSdqO
LlMjnxWYcDPJqxA17D6sT6Vry9Ys537Yhdyl5ypO9vbDpOYw6akMLXQ3wQtinC0ZnG8Gujk9w9Sy
dGutb4/4ew9Q2RCpfM4aAm8OkOJv8SAKk+MT4Hd1UxGnWHC+HPyYNdcoqSFbyXtk8Lt1BEj44tze
DBz+ALDqL4zX/e0xgH95USyw3Xj2cj1A8IJg8qIHxRSIH2O17WYhygCxG7fcL2n+KKQpgYZpSRV3
FO1gW597wBlQmwd1yYN51LX8wxBjXs2J2diDZDtO6iquTdi5yRejxNabpEvpzsuzDClf+wQY7xzq
cGTNHVMIWqsRRkpeop1CPsrYNiw3T+bI01x1WipcdMJVPiI7GnwC/c0029rYXtqoSrNETvamqDyJ
CPqw9VxHCzfiA/iE0UPvENlJhCArlzliXgZ90jS6Ei15xZDzHy1pKEpA6vP1E8rFsXO8wKSaVcQV
Y7cNJzzw0gXefnquC9kFmHwyB4RaixKsBqmgABNtanCbgPFckM+ZyNErD8uX/PajaG7BeGz9Z0R7
mjkRdVCQQcMzq1K1US+UVwBGG9vMcTZBHZ5fZ8Cl7UGzBsCo/FEc+FSkVHK+ILPKs5dSGuBrb+kG
wVTqP+Ea66tXRXaGKxc1bQ3cEpxWbNqNM381+I/IjRFJOeLYlB7s2lCJm2KV4E1G8A6j+qKOi0ZE
pjg/42nNsduCAL/z2CrTZIqC0e3l7skIhnMqyg8WdKtx6AcFGM+5ZOnu3ASY/TiBmW1jUUNHVuib
LeALI4EdjDY+QS8VEJdlHJU8aFi2x4uTSrs8AUHCzPZB+HTIkGVZbfBOW6l2j/cdcsZyklBcH+mc
pNQ8gyN0f97aDnstxcqQccxVd7o1HqlR2GeANOYVU8cnt8ohxhwUAvbOeKOj9FZFmLyfUObQz3Ln
zinpfAXK7SXS8DmyBrdBhASHy2UvlWxjS7rijYJ3t8N5MeqEawNPWqncIyEeuGcOOwi8aWctAb1Q
e7LlpO+dxqCpgVgMhYBuXMcSkSG9WiqaAnOP/z3LBInpXWUebBzbGYOH/PMmPj8FLVxOKhUEcops
RMLJmOWfKg750lkEXvFVYB1ITVFzeXskKY/On/A3mXLSmAh4BRMO7A5wZRnY8dhoqi3hw8AJaXj3
ahGA8cRGLAY0auMb3VAFOlI2pNDRgL50MqFYpmyIQUJeiSHhNLS/q8JwraqzybCUvDoDhZ58xuso
C1e9e8QvnFTt+nv+Nsvcbb8LZ8N1hr0Cyuow8QDBTHsoLqvr4ChpOBAZlN7fDxu37EDhuxWqWANU
941t0u0KwGV5ucCKUA/gf+VRbGw7u/Zmc9VzmU5anYx72YZwMg3181VPmFLVyqrSI+LdfxDS/hmX
kc0jTw6337SI6/roBk++TZzn7qYmVQ1jm8f7yIcfg0KG+orK+DskJ3OEsXjH+HlqUh07tWWf/UzN
KRTASBifh17k7ueMUm0TMkj1KDmfAp6qzSSMUEvKGighrjGGSC8LJNrB/ceCaS3nLCFsDTpezV40
Dwf0wULDxgxp3Q9JIjTOHfXToag6QjlDfDadZcNjsmxJcTtRP7qU4UBtwatxb4T2zXisRVa5DbGk
1wAoA//3iX8WkfS1kmicNmWeX4tQtvyXmrQsERUbWS8oI5q9UhDM4QEiimQtxWpCoU2rhisCQFFm
sfyorpCpzoMKjdQuXWkHuLLijT3d7/MbeFJdiDkeJ/7+y47b2JDSP9BcP8Csff4GEfDIKRzYEteJ
mRPcOhnEGDAH48e24HrYl1ozlP5+2wlowW6av/et6eJz7EyqZMn6maoMOleLo72AdvcN1pwTgMCu
9uuYri6r3kBMLWAzZ7kROrG0IxtqEBTFs6RDrbHeI0tnY2Chpx6WF+4crOw5H7f2NlITH4L26Ddo
GbwEa9+Hz+7ulZRwLJZQO2X135mZCx8IfI5f14RTplb0CV8f2ECeT/pb2w+xRnL0DwjG+ZxjHi1i
/rBCfR5ewiQLVHxQAwVnXGzX+pZV619BjU5NdvOsVyTk3wzFZX8VW87uakDHv/6DLHO4ywHG28QU
R9WV4CIOzL5lwSbAD9p3SQIAJU4nUAloJNp9+lOIJsS0jX5HrwtsOWhExrER7EJXC7R7PU7bFWXi
XnJ1WADmS+z4rqafHrAgUB8knB+PRzHrXPi5057CtV83NKw2pymOZMf798eMf6KsV/AdmPfNLuWn
fXJyH+y2y1GSp54CR9O+dAevGlST1BMRvA9nVNlZLjIMy+9XqrwNIfQYnG+TkCArDdj8lpDSb+TR
G4rFWe9GS4tVH8Dsq20Tl9f0yiu7uJRL0BuzX3KmPMhuwUtQaqCWWVez1RyL52whBBT0aDsF5YLd
MwqF25Wkb/1rTGfbYpgaEZVxZ6wAh/CzBZ48XV8fDZL50DRWwZcv5Soy25HOpM4nX5BE8DjQoO6s
jwgFDcHMddzHRVtK69jwDkvXzW1CvI/pUX+by+YrpvEWyRebNM1STc+2BK0D+pjNhOJ199ss/t/K
FNuUVWR66YEPFkqE0DndWnpNzDZofBDz5wbLVuBASXFdRApr68Gp5Dqr8T1qUO+n1DJIeCQ1YA71
avl9fAA3euQbAhwsS6kftsqW5p57VrqQ8kVpY/8KcEm37nFXytamp5GokqrNeUV2lU23sbAMKoDE
cX7oaC4lF2iVEiTqCs8m/2gQeujKxFN0Ux8Z2BLQTVmUIbiHhT1wrbHyAqS+F3CNHe+2Qfyb7sbc
7IwtZjBu/osgghdIV7YpLsCGNtZS+9CBTHAY+6AbCVqS5WviSEQ5uwTEo2mkbwpES+usYq3Gdxa3
/anXhSFwoxmSDg3JVeTjDB/eEKxVnqChq2Qg0ORu3D1vm4t8R3cXtFqB65Jf/ud90D15k3Opvevf
s5ra74sLNqvJoHyl/TVFYLUCPybhyMPO7V3mPiV2Wg8rcSAPVuvek7hVEMHblFJoDsV4ugdItREW
5YgvVItipBbixqe+xfl3P8cwJ3CEAxMfRdqoulAMM5Zh5kxVEJI2MxzDfKqVZHjVqIOCbm4b6QYY
aTakPRB+YwfoBnjzVWPqHtjTMJuMwJ5vk1zHffRBq5dGdetpPa6xpVEIaAdPR8seQ557SWxfg+x5
Sxt20Ritwa06ilwOoAk1fe6FY2Q8/mGpSkPs8wiBma0JUw/aZnA4+MFwmwzSYl1NBBbgl78Pf/58
QGJuQgGJZcV1ptrBogOkVM54OC+nhNj3byNaqQR6H9OHffFzbkp9L8klY1Z+NjkatUWfXusg3hI/
iOtfpSdA2AtQmnnGdJsSIwuOL4LGaOru+BHUqYcKzRsN3mCkA2MDIXBuYBUUmTEVhHs9VpphCf+1
JBJCVCzHzkb4wf0Tf+mmZuq+50DpbzAA9R+gagZJCqbDN9wPRSMKfA3WHRdxZkS30MOxwJCHg1rh
670hiWij7wlmYGJVAomXeYblvCL4hvRQyNDVrcdYnv7v7rHYG4s5+mtsTfwjOo31Sb7twBOKC4af
P63wOvljotGCyEdmjifFAJS2wjv/kDFmhWhPJ91E53CwjPTgFVAJeLYJbw+MxuYIwt2M9PphrxXD
ntdc4MllzldIz7ZX8x+w0LEGEyqJwBNJpKogn+VBB1oPjDzosDheIQYGNqN1qln611QPhrbqxWg3
47owDBorKh21+uiaU5t+fu2Ek3/qcCYB+xUHOMw8u/NFuZOc7L6Auj6ZhLO2QV9TFqziQic4WWB1
ZDGrhIDi1ZfBkD0cvnunFbA+lpazP7fhz1Wzf19OqSfT6emSl4TPGh8AH4Bjb6UmtLHgt6qFqUzI
qc4r2iKrL9LzMjNdUwUsm7gtXCDFtPkZ5TumNs0SXR5Qyyu2Q1rDVFJh/Bjve2VCop8US146y/jO
l0okPj6PKlTCrxmLxITSDO04Nsb4zoo3qWTc8vI8bJXh2vkccPdJQqXtkEta+370hJbjRGgtaNDP
c68PuF4TQFoLc0nxnP0iTokRi+96kAm3Yoowe3NgQEzur+95AzrYeEDBmDmeDDba4GXZphE8qOrW
GlO+wjbB0Idc5QK3yi5NkcZce7hB9ZdR0hMLxyGViUrXAdYNW8ZjtdQ6x3SHOdv2RduhoL4RGZMP
v9Ojm/IMCCbHllJ2RZuW5yTt9iLZ6Ja+A1MFjJgFkwTwlR+08VOPXj5Lgj5rPauOkpggITEUfkwZ
L5nE1Mz+DK/SuF55U5WHsikOUNWevj1R/NYTNkcR0FWAJZIFULAkgG7ocR1n1Lkwy8kRFOHSWmbq
jtQtDTW0TohVHo1wn6R3ciSZ9GbseIsQh/EFLfzyHRGr/LKuGlcaLnzDS0SdhVBLPi04ykQGgV9l
tYoluDhivRL1eCyAhjXh4fhrJk4VKtu17T8bYbl+cjtkj5szfBTe41e2bojDa4prv4SjMbMX/sZk
BbPj3JSFEwBo3y6pZGZSDkk1AJEyLFL7GRZ3b9cRUwniP870Y/3wL+QNf38QVUlQiZGMH/g6mgpv
np/k0d8I1nxVCzs8AP7VIyo8wAfFFogMpiJG5CV8AG+aAKemnnWgMua3/Dw7agfK4OjJiqrWiW4M
tuQVYGGftD5fuftFkO4M067+wTfp2zcZq60AJJ2aZfBsYpz8G6cvv0F6zi+ej0/gbS/8kOYNhnZk
1mKVV5cQm+hFSi17NVswW9YY7cI7UxjuASb2y6cpIGj0clizn0GXyTC37tbDFt9ajRSljqAXpECL
RWGqGyUEF42AmYNunpKalWqaE4VOq+m/8h3HpqEuOkepPet1aEJJk1nHsSCsj1JLi8cpQi/EeKEg
voeq3VXklpyJorFwOI53zHpR7MZmPsfUVso+xMqWCYrmToGm9etxjJAYYfzpChpZGLQu5omuP/Fs
2DeRfWTfiUjSBvXaiBGwx9X8a7yH7ENJDjd2OttdA6sOKXSl+oMRI6KhTJASfkj74UHNFQGSgiaV
KfwGK2cv6ZmRk45GD8HwdxqVLAh1RWlyMCIvyjTXUYLZFiFKra4jdxW3zcmDHh+q6DEEkkZxkI0x
I4HnGdLVlyN12FPdOPAsFU6paqDL5QzarnEG58B4F7XcOP4o1T+WsmB/rFr82YtNWIQDAmw52oC3
Lh1vBw9fVD3ds3MQc5tzrtQsklX3eN7LINgana6weFtSgqgjwIE21EleXRGv4aGghqlxKGUGL4ML
3fzqWJCfqGa551g6M4BT+BcAucjAigFt5VeNRBigVNlePueNphBcgl6dNXvuDWyD11ZWuvn+YC0i
b+j9QYQQUGBVuFIO6/VQ/3LOwuwQ4KSyqTnLISc5IM9Ck3+juvHyg1Cabe1WFSswNqRJcxQ723mE
OzaNmmDTLP1/BCdHHIv/WuiKSMCJXp3dEpsintlAEzh1BYdU9C+7m16n+X3crjv5mf3459wuHGQx
r2rWoCAzqSV/gAuKia7trZkjjytjvDjyGTefEU3+f5SzH64F28QD9gwxmz0Y9jkESdPTnDzocAKQ
o7KS0Y6h1tjS7UjVxJKaHUUsjJzNOTxyEHGoclWqiXobl3BvU4SzSOcKQJo5VdmzTlxbCfPNk6ve
cnh6LFCSWeE5oTx/NRca65RXQo4gSbpqv6c1CqGluPdgQC2+ETXihX4niernjqjPuCpC6XQO+qSZ
l6H2ayEc0lcf6umrBKrHs4jvjmytbLveYm7+H/KX6giz2h8pLGhZpQee7CX+ba5TKvQkTxz4+P+3
qnuPuu2velUygmXNlFQM6zx4gUkOCKsYWzEw1ZFra84aNAA/2wod8Hhs85Mfzvv1rf3qN4zFeLJ4
gc/bfocGi91c7Q9+CGjGG+ZeHJUxDs7DHL8jPPMoVC3TuVXVWMVzHaQNX+NMkz/hUrP+dEe4VzSV
dJvqMMiFARKN5twDZz0aSHVrYzerqbCNaB0LTpxrYOxJ06CphevCv99GVrtwOh114IK3RrIfeoMz
cHF65wgl1ixaUm5MJGH/5VmnuCfYOOfetwXZRoYqFDd09PXY92aT/1CbSN02AcExADrlrF717Qqj
xLkrAQHuAe47TNJTCeSOVzRjk5Vh5gPo3f32OKZV29peJMAuAhaho/I4NgPf3wloDTFVG1d8M0+a
JiVqD+vEagp3BAhSthk1HBEW38gh5WO7n/vNTTzTG1TkAu4Sp0CphZAPpp3Z+Sek6DcvHNOhnvB2
w8W+3TEfjkV8w1HrKTcdLMz9+1B+FW2BkAkGEYT4s2v4Qr6EOpn8wdzr545WRhlWldz/jz8T5m0r
pZB3r4mrDsaM/g2PzSwv3jocJSc0zX9DzF85uTGSTkxFaIAo1o0EOoVtvpfdsu83mTkKQKnsDzic
S600lfJ5gOALUunIoCxui39yNBQOSmOrQ0rhYKAoBe5DG4JLkk2oCDB+KMJBkIhzwj0LXPdUj2qh
v9EYfkN5KVy2DF2FU+dFTGn7hkAtUAKaimEIMTEEGgY1yNjF6gzN7ZFNmHltWM9Ajtvh8yImOg7R
7h32EJ+Ei9aAFZaorZPdEac91Dtz7qClVLLsB1hnr9Undc9ABpKACrTaVmRuncX6VBMTUczrTe/X
KDQ72bFfzJjGqLl+hB1by5tEWAcdbpXq77RDD3vGnSZD4plPsOnPAaOObg7zQxITXiDNi8fjU2Ie
ieWIbYpFkye/BOr2e/wwa9dhoxVpKaVOAPmP4t6zAR2wKas7EnkMcqclpNLBnIQVo/pMKTO+Fhm8
eC7xEWQV1CytdDOOjXaUt89mh2AIS1T7BUAd9K4o1gfus7RNIjAdGt6gUDaO3CZ/e28NZihpQ0YH
MbamOJZLa6TN+Rn7s486R1AEEIIWIzArCE4w1tudPtBfNoCaFslS6R2uE7F3mrmtwBX+51dkXaGR
3L7Z6J6o7Vej4ukgwR/8zyhIIemJieegNtuxzsCCrMKdokAhH+g8BjeSeZoHUEMAIK6ZwMbOK+uF
ESJV3jDhnZ/uzo28e8ydZVcDl6NIOpJ0o4wfvdIO8JleFuUHfxu03bbCo/41sPyAwQEs+/U/SdcK
YHBYRkUVrlxEaUB7IJ3Ghvc7iMZ9qX6YnU2JMtKPC7we/7mpkCKc1WigsBU1K0KRnJWx/0f3Ts1i
xGMddCLwv3JpEmP3B4oElfNNfFWXJjTwoKd2VpX6JSshQ3H+lhyUmhr9FdqV/+tBhGJOm5ZBktL/
wkDO5xUJa3eyJeB1AmoLf/I6RhHg8IDaNGdwPHe1qo7xrkwxohZgexmcAP7XDHXhj64KrIUZQSQP
KqnTPggUKfrHHy0QLbL9u97xr5zo3ySOglBRdNdAjasR/d0GOeZJQlA1pXYPFQVFrCJgNKGIWFUC
aVYGZGW5SUT/WVOAtcFfFFNgOBiTuBKQY0nwvPrVJsvMzZFINfHoCHTGPcgYyyp0LLK8fXZYbDkh
Sl0EOVw9eYtDG9uGUalI4GbJ20feT3uphYuI7L61lYyAfeK3lbD9VbtLonJdAMv0oAS9G9hC1hPw
t6QiO4XMgvzRH7ltudwVXFpNUPSe8Xd0NtjA7eiLILQ8esMkzfesUmuITbUE+21rp9sxZGDwv0vh
41N+d7xsIUzsDeCqQy+dxSd+T/JnK02a0JTQs6MdrdLF7vn0bAHWDW1wyTSDwWE9wUzd6ehpEkEY
RFKIWc4yaC0Q/lbJlSbHLTdITIP8xg4MTgxxP/gNx49kPcoPh8dxnYg/rczbhiTQQ0vm6eYHlcBR
qZaLCzF07vQHFT6FWkw/cbf75pXBxjoe6SXkTOwGYEPifT8Bk2McBqKFpOgX8bQw/cXpCbIyaYEp
A51IeHYus47N8GXeDSMeOAvZEyfqVntnMpWQSmPeDIJ+EkNECYTZcEWIZDlDytyo1z9MEnFnE6co
y/sDhJsjoqV6Ys0fRFgxLWPP2CWMMaXL/m1tw9BB4q8U4TKiFKNxGT5hN9lEbmrcWHRjEw7xaETX
0ZcGpgsYoSTrej2X/8KomwZpJ0Hmw5RcovGvGXt3e62WIs5ZM+8tDa9Hpku7ziSTezNgqYEcLdGr
UOaZg6PAjJz21QLCfaWtxB6ByYU/oMzM5iQprDlsPfQCgOwXETSLot5BhbLFkfURErAzhQRW1qqp
waW55tZvewY2xWVGj7Q63UllGDYnU4X1k6YWBSgGZgDNKAnTqqQXrAOWHestUYFLtAPUK0fV0TWr
THQpmYxvQztmsaDtfF0j+wfb+0B1Vk6CSYoVa285wRhKwWQZ2pLFny3WcXIoR24Dvg0VEsuns4ZX
rwQNdK1s4g6ycOYa1Zsn6cR+Lo4EkSDq5/Wkv613VAoh9b7fxQJTLi90nRPiFcXdqaYmRRIqt5as
3sisk7RzckrV6uk0fZfZYpjbFJ66tZ2CirhVpa81xNDgc8SYctGabjMd4a6Iv9PxfAFtrnbjATwx
wKMSxUbQrhXMZPbGlSc6DrfdUxaOw2J3INnUB8WoOK/qd2EOnSFV+HR5XtDKj/+gA5Y/glDpdYUK
MsdlLtwq0aCvNy7ts3V22HkrTorJK95yH5ryB9cHRxj4nyBu9skBj/yNGKDuPA4Mcp+8m1AYUe+L
Odb8m3Sfgs6eL39Mz+EhOhr00J1p6WnzMhMyM5plfhRGeR0M4Ygh7/6GK2jCistRfLKiCEPqc/JH
b7t1xYq8dferAh39jWvKzBjJlSZ4IlJwwNaBXFbL99U3XmC7mxN/9L+iMDczU0OpXKYB7/Ro+hfE
IufeOldAtIRkUNAnt9A4qYrZzY4ePMq6/Ckb+vsI3kPZyZJ7LYN1SgMB/xV4AFjrPTBv4ernsjoQ
9M648LI8i/dBEu39YbkQBu6O42qsddv+vt8pyntXCEySvbcdxFQGzfzTva3CvoeFhz4bZULUYr2m
s7Q5qSSuM+Tymc79BwZdhF4Br7LqwSfi2zqcTGS2PtnSGDM3CIhk6FVdIKHxBmGI43XKu9ZBfyDM
oe96gvH4wHQvAapamu//a3uERXZiVRuwObxaZWzwF80RGvnhpSsMgXS2BWWmZAMlJIgGW8MD12WA
EXsGUV9uCLbSpaqn0Jl9O44z6oAbbfZDBLpH3CP0eJyKYiMEMEAJXfGyqKeQUzFSs0MHXv3VcIhI
7z6pXuC7ut/8nKLphYuRvN91gJaeUjpyaMEe/Dzrvm0HPSUh8zEWP9WzYluXn4CooYLdtZe4QmM0
ALy3ifQa6/dQJleyp9nhLD/PuRkvsROeI0A6GkMk9RckX5zp3NP7B4jDypYrpXn+AbgFSziaSBT9
xpVaubF4eKkfrAAORUgzyQobRw1lCD8SW8VpEd2hD9GQKMr0HfHQgv39XyjZGOB+sNlIPS5VtPQD
3a64zdFPhLtKJO10YDgdYUq9ZxTgrrJ9gkV3J+dBePzN2deo9L++mzVnUflrv5wmgruubeEwm7R9
23e/8vYcuCmy0KLd76Kd61eT/krYFfXNg53xJotAvsaSRApkLNcjPhmyjLEMhrk0Ja8v5dUFfD8Z
GFV7cMHjeEI483D85nuhWOizTVPHnJZGYLnOJrpBzwu+FGh5Nbzlw+vlzQ81ilSSfa4sbdI8hNVk
z9ZVzIsU8T31tkOFmDaSxpjWSo+g7OnM/52cEfM+ygBhBXBGNILv3IPrP4yqi0Tv03iymwMhZCSF
EMtBi4OkZP/py2bRroCWwnzzsWawcH387qBw/HS8vvzL1WYHPj8evyJAsgNnJfCB0xOgwucMoPG9
QsGsGXo6n2vOejjm9j7/Ksd108kXDbuhkcc74HVbnv9cKDb9LcJGILMU6NRwAalCM1GzsHE6ut/I
C+v8gH41scsEhirduahSe6I56pFk9oOz6H60VejhmTd/1TU5XHbHVzDArL/xmPIX2X1J76jNj4Y/
9m4WBPxO9AjDQvxavm7UjxHvy+eEnJzQHSzQ6niB+LifPkcD1lol52nWL+M+t354vg+YUrwwf44/
VWwLXNR6kyEMhVWuNaBBuHSa6zS5k8OBcjx8+B5o6JwYotEQX3UBEW+ahlnudhdJJL4tvSHmmQ+2
ufSvsywkgnlkiQQY0WJyTj9/nlQbuo1kFNCFjEBzteC1It4UPjoaWsXczFR4qwsPgP+hpYdFGpL5
JWBr4FS0EMBB614yZ9AJI7V/CM2Y1c/hZaGE1FB54OwnUqZCVNqST0vjVc3H7kb8q2R36q7P6Csx
jTVseJdhJHE1bPEEh+EMDRVbUqrDZxiGAiae910ZPzmM3TXWfchM/mKM2Xy4hTJP4QR09W9S3YyK
D+8gVwXW/bCNVq8YT9gurQYqNV2cGRYb29YdsFSwYyqnf54lXaEgeCbjqreATdyc4NXWScblPOL3
kmkHXSuYYCeSdgmnLSuS/K2NGnOANFCmJd6iCEWyQqEa7UhoSedyNE7DchNQIPbYub9mduTJslkv
WmKMLup6AKIz+5Bi/L/fMRIjC54W2Ps3c8LgzfymH5MeF5w657HBkLct5BbuCSxM8oYM0djMB0NW
v2i5ee13Yvg2Y7BBkDa6z/QkW1hWQFPwDnS3EakK5dc4vXUCcTNp3z6nBB1ILvwWz34HPtIcJ8Yo
PtoR86nsskd8z+KsyXho8ysceOXdSwcUavvSUqj87Fi1UDpPwbIapSZxicUOc+VXu0pP/FbNuFfd
24H3BMdrjUPQq5qyjA9ui7dGy+PL90up0V9tZNuCHxM9F0qIbdhEimuEKJVaDSel0QyGMbt4STzW
vLb+pWnNt7khE8HlzzUrq/70qHUfZ2BKpLVurI//8Mu+8wzOHRHAFKtGjVpsxstUZqMXMuQF8L0f
bFAUX9qGTOAN//69ORf2JFUO4u/R87o9aCCflFOrjjJFSyzTBIlG4OwrmJUaFpA7yjYtEBTndcRN
Aq2uyAsGLqhrtvO+3hkApqFMO0G89gleU2q3DysrYb1SnIEUKQWAP637vxDkBJoHHO9NBlDr09nm
s44DCDYYRNJZPgHoOyi/EUkOcE/F4fIUJbH7vmgufTLAkfOZKWAXAnPlrU2sqCEYDRixx9KAuyGL
mm59J3awwJX/Cn5gWnlNQuAkzjoHhxt2KTpdpEXkN3p9OUKbYNfJbAsJeVPYo51hiqKcnaOtVWpG
Jjv70kisiipFn2RHiXLBOIizjH59mcnVbJrzK/Q36/8ZxEZMtyhJK3zmqeESHYDhwGt+ySBvmfK6
pBZUr8u4dfaOMYRLENx8fbSw66PtXI0lDG1aeoDx60w4d+PAn4tChFliLZzyLAV2kSGyhZcmE4JE
MKXta7t2HGFaRmRHU38QR8wulBJfrIhNQpL72rEUHfzHLX3CX7BNTXvXkj4HkERgVeGIG5YZFcIZ
i8bAWl2+WmAuWCDhMhVBe8RiE9MhZy6oEk8SCv2F1cG8CKsBpwmknRG9vKUj32AuOnnifYQpGxIS
KH/hCXUUlA8twZPCN6sgFU6OTVXFc4w8j0Tz5HDhuunBdJlCCHsbhtYXdXtMJJYcon14YzI3Sufk
yBEphb51f/ojPkb0zIM4vTJ5QrQucj3pGVm04QXZtcc650aNdGXcI1Z8hna8pQoOBekTDOjQ6ur+
3YGixxXcLPiW9z31e2D7/q+/rxPguCPJZhxK/zGxQ9QAMC69I08SgLIX2hMZrdkUWqc3IQnj4w4V
JKpHB46qpO62XDwiJ0yPQwcFxgU3qrTBUSBVDdq6Jfdk6w8vLdlvcQDatwT8dc1rxK5K9L/fkq4H
d3KvCp7iUMlrkGII6CVuPHzgA0TYoLFdJYUR8dYhXQN+XPS2Zl+XkFKRO/z4UNeF6uyQ8cLtpX5x
8XmgPThdRBsw2slipjrKC40EmJuFVgb8o/3obAF/lzQ9cAcwK1fVNc1sj4wLiG9vB7xv0h15Fcpi
sGqe/AovhOWWbNccikWPIlwkEsJwVaJ32HdLVnr6aMj/hWgJkJbniO9+0TpXsMt/WrpEgJSVYrYz
mJa7flcDBi3lbvckoZJkz2crGhYQSBdbuobGQGSubV8kvADzP41bNfcqSXcfnyBfSdEn1sp2eJz9
6Y65F05wxUZ0VgtNTsJpYSU0kIKKx6UJFY2JnaSSZ+RUa3UOsb/SwX/3uromWSkOEQH9kIciIfFo
/p33LFoooH//ag46QuFiVCweWDzYgetfhuOYKTQ5A0SLCUrPa015KD91Za9h5rMCJB6JsxL5q+bJ
hRTf6roIbCzl4my+JjfWyrfTh1hpf959Mbn7fJjKOPsvQdMyX3dslE/vnHI9s8bWJQ4p7dimx3gL
JIpAILhP/jc/7dXMV2IykZBwwB6mYbIpJE1hpLY0pJaN8TAVyqFpsvK73qCq1kCpt754u3YSXZMe
wuxU5psbsafLPn3re78BX8cSc1tQhT9HUl9jcfiYcLfAFyHFdj1b97sf4g+6OifhcrfqEdliC4wG
P646LJm3qJOmOwehEaA1tJ7cJZFZ8HvQpyvlq/AsefiURrKWx4uk89bi4dysGKi6Zv+V0irEQ5wP
Q+BJeia0j4gD8Yj/HwNaHLiRUBDz2ueGvy49uxKvTZ30qxopNXlHOb1DdEpuqOOMKe7y2JHEtamQ
hZwy4Cm0adNCYhWPjklvU1R0nPMwAskOjzokJq9n5lIripKnO+3tyA5fqxvJYAYVYso+2OMIDyEY
IkIOlEaylGOolFmHVVvotccjzL7s7mruUzh2csU/1LOIcmbrMwPzRJuyl+hbKOsmxtdIKp7HSFwC
wlXT2mgty6jHmuUpiqYnCYLyEuK3+iENE6CUg/4SYoO0IbJqlmJOTRu6XS25UgmzZT0Jwu6HcqXi
c9EeIb8zUKhoWu1kyEQdlay5K+cxu0aChuUBvfxlMNIJL3jTIP79cIK/4CMFRtD5nWMqYTd2XymI
Wdm1pX7FMjTJ9Km2qCCrrqOfmhnqeXaU93YfxTindrKEaIRB1JzFmtmrM0utmmCNlPdIWI93IxXQ
CGX68N84wldnxx57gdfD+LaN4Yes7GjU78MEl82JJsQ1kOUhVa/AiRDQX373Qbig7h0p0TWqTNjU
J/cj1Da6iCC0R8YqiojYTF7+aNUDCC3h/TajC611WjJFf1+Kkp54JZm94ioPBogfwGek901MQp+c
Mw2YMSTMoe1Q3gAw8ztSqtRy1ictxSXBXDVjYAjv7IlaTLsMs7VffQ2beRA1RVwnrr6tiwUhidES
oLqf18FSAI6cwL9M8jZW7TMFUFW1MpjC5F14CChw0MYpJ28SBTHfefmGJGUNSKIibjtWqmSV02EQ
P6meka64WUxuaoSi+sALhA64xjhTvs4HQq4Cb6MNc5GcB0mNsIiCU0sUDOfPV6UEKf7gvqqwzMok
YivhQlpkdaFevbHh6h8Div3Ug6p6Gd2YncTODXfteBwiIBudV1xkeNmFNfrrk5yxOGxlZFDWHcNt
bBmENwqdjZ1WpWP1F0nrxHlbpUERYRmKjE6W2gFjfpcoqBJlcKcVaiHLZTSyE9DUVIA/XzR9ESK+
TP+U74XIbc+/bmxDF8VeEM8+3GnRwYe+NzNREYoH0yc3SGZhQlzXcnAKl/SaZ4+6OnhtITeZ41Ld
5mstJS+KDxNDXPSh76h0+So9Y/NwkcT/gSSD/WmKg/8ie5cLH6rhOuqsOq5Af7StnC5u/wZmlg8e
NHQ4hd5FMf8JvysW38iwh09VCvAtJ5EendOmU0uBlmmdWWojAOOoZpoJjxt1P5Ax6xl0cMBHpEUj
73IQCd5I7EM9WT1fx+sycUrBk42mc7rLS7sOfKaRSzJ3fq3exVaZFHWySmZNUP8QTHa+nRKWy+hT
q4WliX85UDtJeCQmfyp9fWpN3ncn5sGnxyQ/bL17JtyHRLHHYkh5ry7epTGxSZDZBAxjQsr6XPld
oG2Zjpv4/uM8Xn+LqptjGDz/MQijlFISkt6UZwqMWvuzfgtHsMGzkFpOygUp5iVNRDVj8cTXBj8Z
MwGPHu0TAh9g1RCoLlTlPsgEU+xwP99FljIkDt823/J/yU1Lc4CVhMjqwOc2nZgwdN7ljzuc9NUV
zEe3+nzy2pwstsQomciNo5PJIbC5YN/+gQjLXWNp0et9XspsqoCImD+irzFiPW33XZX7E97bvzla
2cXYJj3Yj7izqL5Q0vCPeFI+TzUl1L28a8GdSAW0RYd80Yr5Q6daQkBUpkn9QveUgFPczCX84hUD
QlN/xeuuE8DEdbVq15DFoeeGpTdEv/DNR1PfY4MWNcmCdOC9wL0dwsvIdNl3XpNeSHEjaU625Wnm
Pt2ztzOsfW4MLeo1CCB8XvlqgAcqezYE8eYxRO6klP39u+/U44VEyVQHrYbFJ2rNK9XLCw/ZG9oB
I5nUz4kemwTYuhZjUPY9P1Hh99nB4zJkzkOnGwAlLBcDSJN6b9b3O9KwtqQ52hGUmekdFwQkoWc5
K4kQZA2AwUISFbVilVElR7g6bbN9HMAipQTW+NI7ZJSBmsPqj51LF2x/JFppLDoKrMR4AQSvuOA5
c/Q/HrORJYuey9IROJYzuMfxj6rqGBxPKYmUiXykX6h8ucJtsfSNNS5G1f5YxdcLsvtqSOIjzTDV
lU8YCohk5GULEMO8orLNmJwGFjdOJE4IE1w9aEA419bdHsraI8mf12jZRmE+hUu/Y8q6lkmb5gjc
hYmU50J9FEEVFj2gchNegZNPk3q7DaNTCJwyhdx/CwMZWyUEsQ9e3jHDC4wmmOnWoBjUaNvAndni
CVoe6v+e/fQFUhK/pSA+5p6RMg/eo9S/2iwfq/wgnjPda5N/PzLT0RF5oQ8LifOG6n01dG53yOQG
pI21dc4rFO0+4W+FW1JKUJeAzX50mciNfreaLtujgdPKFiMS88eOcz5PW8yarCkbNZAeYlr7WFNh
+6Ax0tHNNiwV9eYL/ftM6YG8x85GLik5DBxzRbJz6/Ssg+B93JPCuBue5oQqDGHoOQdxBH4uu93D
rLh19izQQoC7tL4BWBK3gLLTGyaRE4U44vAe1pX5Y/uBsvf5ahx2aov42jpX6lD7so5oPT96E9Ok
z6StG7WoVyn5VNz40cYa4gNldSqy1v4cE4A999Os7i201NqfXl8xrDvVgQ6v7Hs+7KqFBb+oICXE
nOTDwLI5bnwlQVQx0e8NzA2B8PHwe6qkcPjQX6J3p8+LbTUfkH+j0f0fuk5lfs/iWmQMHAt4eZsd
6AOtSUx6h52+q8fNWFcVGIiY55dYMAiKwYGW7uIfVEINoS7SIJb0yrL7IjIxEJsORAAKbmu0CYzp
IESfE3faOjGWjVOqb064cU8D/v8//GL/49N5T/Enn10mDJqoltoUU74J+bcyUpsCKDUA5fKHMYY3
aOM36uCrTaDyn8RvHxXD5Vf6koX/Qsp0ObVTdBdjav4raCne1iQFuXWlEnuZelsFKvNo9DwrI/sc
I+Rkj4/Nx3MxbbKluxEmaSMq80rjCQVhZbwtPrtbNj5Rj/wIcvUDk603twjjz6abRDUmQLeNxo7L
p8WqY4k1evNg81M2L/QQrDETktoG3/k2SPrLEOfHZiRCqhBNYNxWuzZjGs4Q1qLXfcbdTEPmUp6o
ox0UBF05ORqwpAORwDtSh/pj6WQ/JKgrWv4xowt5f4D5HiLBLKmtPd3wYQ2HMeVF7KNKcCci/5Go
LmZhRpZ+EuT9EGG5D6PxWe9RSvGFKHmpwVAgEmeh2IXtU8dhw08wLT8RqQ7fban1eAwf20NMm1Tx
U4Jv4iqb9LEigipdc1nyv3no1wpBfj4tq792j1kd9ugtfY9gzYeV0O+RQqeuoErI3jDbF0SyhJwN
YDroucTcyU7NzjRquhU3SeFhm2P8YBn5gH3yoCieRbPXwVbSkvzelru1FKY9A+dCxRV3uXTvvO9X
2irSUnFlwmMsXE9obUUhAJFWU+JNKGntnIH9a1Fu2WMuOL1MJRTd1F6EGWG1bwWTo+xzBHkaFR/w
4pzfPqU+zKucOclxJdi0bBobWues6v0sZoF0y/ExDsxl7ZKEAz2Ysb2xXTFAA/pViBql42kTazSU
QfG8wrATN3YhyKHWJsmCLaFPEo5WKUiyeKFPdr1nWJdpwoaVAdT4k8s/UmCqQfYSYYfT14atpysV
81cIKLSwCzz/PdvatH6trFh6XqOt6b6FcncHbnQKhmXNoz5chGhzYKahedF1Xw4EA00gw1VSOJDo
t094sK/aKJij+hWS5pZqez8zTX4f6ghDg1xZmyBmI/DAI7wSIjBV5kgeoYPvuoSdw+BRAPPPzvgq
cgutwrIBNXoxGcgJ6yRipCXEMKN3yjB0rMtyTVCoeDf4EHvR0+YV5RUd2V7tJixtrdwFQA5kd4Gx
pyb/p07VzHlBJJEYVrNQntsbxEhNzSEA4C/qXmkbmlZrlflKt+vI9E+AXzxIOVZucSJzVojqblzN
Ij5srwZvdxLO5MSVkJEDoCtEnA66M5orMXPTlyGzGsRDbSD4FgD3pok0G2zkhz5qMNaeuBmix5Gu
RZtwXn6xesGazdV2sPn/BpsQ7DzipY4SIeLrs76AZPUXD4vxBD/pt/mHIk2l3ApHELmsoKWpO99p
+mV+3HsRPu9OFcZ+MUXlMQXm35ouum2goQ5Oe2SG4PC59aYZqFn666YGiQ6w3zZ1xIi6rXQHRfIo
CagnFltFH0yDYlCz5gCGcY92vFqaZncdOVDXhyeJFBGzw4v4t5sKjyzUw4Z47rCueOGi96zbMRv0
n5yuJpgOCyi8YJDBJjnDaMCVggZzY1j672Yqa7I4unJnv1xOzdlmSv4ctLP63OMZVkTVWehxTtBf
v0DEkFY21NtPR2zHIwTpIET8C2jz2nnUgop/fpPpKB1sA2iVjWmygSrMmXrtf459m8OUevaOh2D5
aIJw8Chz6VpJiunjshzCUcqRWVHdaBNYF7h8vVEgH1zpQPPI3xlm1vP07WpN5WgXGR0D+eRq3ZzD
eBUC3jPv/cv9g+5QTyDN6W+wldwkvTre6XXXrtsdmge0WiT5I9wI0todD/n2/UUJnoMDPFjJeOFN
6+A3b80TPzOW5M+d3YPOawkU9tBnrUdagdd7XjwDGeth9v8fI8mh/SxWG9dt/+3qA1cb45fHqd74
ZLnwzXve/KpLWF5M2F5IUL2mncQ5aZT9IMR+Fl7LBbZloVieDe5FYv1WfOsavJKSIpiQMxyUI3ez
IrkDPxPfcAaj76Ccj3OzxWGnHZy2efQ3sHWcTGMy6rR5WLCAXDAdF0UMSjzpIfzD7cO9SNDZjz9/
TNpGK9FbBL+bh0Mcxqp7OcPTTrInbQQydaAuKBQEErX4XHg0/WVcUit/3usMhcIIVLJHe+szp4Id
goOrwwT3oQu4FClgmwwlwLSquk+NNLQJ30HqdSQByQ21X7jahYvGQN/ywBC6kp2YXDFV665sGiXB
8p6ON0lgwbgO0hHBgVP3/MvfOwxTIAqmV60T0e4l4QUKAtAyTluBAJb68Ke3mjzna9WvdI0Z+v5I
/STGlJdyudNUxnyBMKU2Pfb1B7WLkyil+y+r56DrGPGjudROyKkqQLAQ1ghTUedkP0eoi7yPBBHr
TRAKvMWXkamT8JuJ7cZUEubCA37s5q9h4v2xgjxHFx676I5mVlxi64ihcDT0p2xA7uTyBbZn877L
qVnpEj4ez/VCR1IGO/zhWQfF30WHftsyJlH7fQwtRjIPYhAYVZECDS3pExA76cCz8tAaiY3I7ko0
BTgzmOsgFf7eQTQfnu52vfDml7xlB0qe9/yQT+sqLd92IR8NPB6JlbjHxR6MOhUtaxLW4zkL1AF7
gW7md3sr1ZdNIGJ708cIDG5rXZDN+qCtt58Gw0kYN2nToia6gmgWTSj9utQyDvVwSXhcGQTKBYxb
i0ZwL6El654dOciwSDELOJxyeU5phrtoEYFozp7JuZJ/EXeOuldYrYH26Yw/XQlOtNj55bIdO7u/
G4KPYWKTJ44iq5lzvrfYbZVBI2OInM5V7bcZ6GaOnckcyi2EflzHp/JFCfK71L9B7pOqGco7tWkd
puL91JqDGsDVECkqbeKenr3AScOpPVPtbfPuiWhMUumpCrFxBzg1BrtmgzF8Fe1Z6y55zTjPoWoW
Zj0GqaHuuS9Jehpt1uJdShPmuK3zAh0T9ZIMazaD6b8AZh7UqYlK1wAqYfb2FGyekZ/4jaZ9Rcpj
QnX1M9zYqPPKgUaCssBp+DztlB5QWycyEzceOPF6W5mwp2W5GZej7nsvWcL3G+bvNelbY4oCODxx
ZqPvzOSbsn2AXdHjQ95Sb5S8uQmDfNLXHRTI1Pi5MCphYfc5iUCR+zoUkJlGn8L81hoNyUHCmmtf
w1gHlqwEghhGYRjfRXhAd34JMQKBdzF5AaRWg/Tb/6TcRwbILP0T2gF7UNfaFPAI+cvb/VuSDP7a
TBsTMnFR64OrJa9FilNSNvT+8eXSRh6XmLtSJe4qcWg1k09yC5J9K0pPFSknZwFieXo7gHTDPeOx
UZ1Wg9uWDt4ckMzS2B8GqDUI3nlgmakuv3Nt0GRAOFYT7TAeVmb68jMfXLSQ2LSh2SMhaRtg2cu+
aGKucFTa2fxiTBDsbXOtYxVed4rm/lbTNjW1ftNc+0kq8HccjfkyC9z8Yo7wo7a8yPhlmNT34NUQ
f+R4znJi3Kce4Vc8tNbikOewcFXhiyrMrOkn04Je9//cfawhE36D+11ApidBGyfn+P3CSSCJ29yA
Ft3ohf/uLVuLut65pohvM6lCbZq1GJR6qOvh8U/NxnHsv5fmh7ykK7Mj/K9ru9nU3FhCRBK6KU6p
W6a+Ad2U2eZp9ZAMc4hCDLNfv5oacwh6ucZbfOn8H03mo3z0iBRbS1ofniQP6l3A5wWnA3nzTdqn
iv/z3ETvfwAo1LbDBuMWuFSM2dEYPMlaOGMABMsIpbdxMyyJ3S08QWfx1ncTU+YrmNNzEX8+OqSZ
4qFOYIGy1ujxR4Z1VY8CSkBTB/JloAptKAmEiQzG+5FtFqZB670yQtXm0PVd53ity9G5T3jjkkRV
ArbnOH9x4VcfjkKFnWlhO3ozylQIayUxPbqXg9Y3PdZCq2npkh3vnMNaKDnfNHIkKM6ViiN6wLt4
6g71S3i6qs2VUl53CgiP7Ly1xi4VT82DIytmYVRCQIBkM6Hilcv2AA4Whx9WJWFFsC/Y0tmL0Q0B
hRIjVN9/cQ0//Hlwf0I+AMOqM/hb0wivCyY5nPS7eNgMkchtvVUhLb1yoMgDZyKDryBdV+TKIB20
B6DsU/c3nBOieTQcmjEP4AkLDo1MwyeCPrV7cRXix5LIXuu6opoYTH37XH1J13FJuw7qpSfv3Fau
SJJrz/KblGpp6LG4IOAgS2RM4YXShngQrCoTriKgsgHKERtM45fgUWP6fjFR8fQrHckYAOph7Dw4
o3vUHOJx+6/FdH/AN1EEG09HOXlrLlVRNViRE3hDJA6KDg4LavppbaoL++n+ua1+MqLnDYCBr6OV
0MYbPly8WHD7AkEjxRpCe/ADcgkxAFm/BLGhNZi80Lxqt7bLfca+uuBmFwcE6lwOurdzxFeN0lxZ
FFJX8eYXTlW/83aWRbRiwXjqcE4Q/OZhY0+DXBL4irGzby7BX31N58VeVE+s//4yvNB+pPfsLGsl
WcfJSpQwsznAN4JCEMmbVGBLBxFV4HUfyIPe5DZQTUFYG/YK0eoQcPviY2mK/x/I1vGJFdwSMnid
kEtz9E/3BYN/VyfrfIWpVRvsbLBC7rO233SkDHvItGgLhkVfevL+mtuomwt/6dFBsok4xrm3bvVS
MsombMFUoN/oowfBQZEbmPbqtG4PT1AJKhziRxsS9nUobVk5YIoyedEA0DQv636OtvSvNk8sZtSV
nm0aEqxtnzvcDFAFWJKiJOG/+cEzQS1QZzzFH+cXCxLt0JCOPiZx7nfZLZor7MlEh8y/eYbdgWuR
0u0kADz3eDDidoiSyf2K34Oie4U/iImxRv+GILNmEm/ElD3SxsUGlAsadC9wzlptdMnp8lB8bNRa
eJDeMb4UNKiwzFMHo5/9HDP8TvkTYvP9446HFOQ3CZRdoHBvsQfQVuZFPdIUsn2RsDwjPPSPYmbN
334canPF0g01NDLxuz3RPEVhXQj84sAPxYwkvMBWol3AlMbhrNbWk5zLtLseXt8V0yp7hTh8yI8n
oMVBWl18xncoh9ehNnOeS+B1C4UCjNL30vJCNmBv4ZPknBWKlgCMkT3xLLbN4J6QLvRMD7OW4oYC
WCWtaQcnU5lqlkwvggA1MbCtFwCwUMqOEFvjOIZ+FXgbIHtV/XW9ruad0O+2EXWySwLKIxjQB5vZ
LiaBdiySSE6+S/AKsU3wZ2xCThsH/2li52Y6NbnBJPlDZqLxxF08Jj3wN8/SLhxMOQi8LxFcxc3B
u7kypqV2pky56SOyX5AqqnT36rfrKeP1Mu3sS1Facrks6ayJKOJy0ATKlbFH6npujXwWDt8okAw3
RDdBcr4BWJ6fMS6JV+lGTOZ/cxM5qSv7E4MOHkOsWAO2pD+I2lMEXgiiMD5fOnxore01RR536FHT
rRgqQWbIkkvjwu4um3hNPct9YWN0a4pwSsrrcnzyhAi1gLBLMsPJXG4ey7Vhdxi638/LGXV7q6EZ
NmaPVvi89rrRMWZAfFkagfy0U/v16JMIUPiiwiYp/MuLnydHt3djnkriK/qRTAhVkSnFHxe/XEf1
OJkfM3pyV7/oRabU9HqOCTUi0UoPoJq/+xGQY9+0NwNnV60tVxrGJwhwAb4zBXpM/L5WL2LHxzr7
iQIo4EuhMhnj9lZGBf5hDG7EVRy7lNBmgcYKOSnKRGRUBUZaLSxWgESOAMuRKNzvdlbB7htkxLHv
BMa6SAE8gPG69d0S13li2dn0Cl8th4jn/933fHkD8+g7pczp5Hkb0AaWr4WlQ/f20OzfzXarQ2ga
9rXkmRPOPpBAVEUaTsp91mnjVaahMyf+SfIdPaOAJxA8P61GoXa4ly2yLLvMwh4xKFX3wWK2al0E
NaI10aQI8W8Dsz7tCVCR3l/wW05pZq4LX2DBs2OPSUru+dXrTE/ZqPeZ/wNSBabuw9gijvhwcyiM
ghEIyvfoPuiDmDSzVknSTd4q2aKreA3VgAMOQu30sM4jsbn6Xtm9bJraRNFKWl5Mu5XIh0KNok7H
PW72qsdrx8Y1MEnjs+59GEluDEu6aU3JRcNGYxVCtY0PNnp69QXzYL2V8qbDZnfLVKXLYM3hlFo1
P8fzhMQVtpH+ef2IIT/ATshX/V28L+tLs9tWIIGK74csy0EJ7FgHbla/d4xroEP33A44pNV9t+n/
DpD7LuadnVqOjhEb07DdnIDiY/4U/REwqPAGOs61CWvMMuv2YN4MP0nmN0vSZIfpXh+UWOzkCo3x
20wgwj1dRHZRgy6wlEKoi6hefb2JZdWkhYqJ7flTKMfOc2ho4XB2Ibqk8HuPpf8D+yB8YH/2sD6y
nXhCOuExlZDkJxXuTDNMFQ3rK6EiIqKeAFal1wAlNa5sqQM8m1a07mUKDNhkiCvJKlQimreMZin8
MpazasLEGABbaAiFZ+Fsy2S7hsWr2YMaymYFFkyxakeVC0wbIUkhao5xFgLxAO9vs+uii4DSb9UO
mIn+GSx7l8EIflL16CNW+mH96g5H6AULmOCT+a0EgyWjYtzo0eJiAwUMDvlOXuuPNx7WmedoJgkF
ab0ScT8jQ5IOsW+IBGqGi4qLk0LOzdg/Wv6Dnh7FrWggmz6Vz0G3Et7CGaYbVMLSykiY3MYnOYVH
t258eZ6kEDR7/qO8g8W/NjxtKoX1kaVs6I5VhDgPTzWJ+aejSgU8FcLHbCR88qO1UbEPA8EgbKCK
f33Ep75ZkLITQzzkxXl37F9gB1z5pbn5ueEsYryUPHspeslzdewVznfAC1ArRIv15GnaxBurKOOV
1il+8jVl9duTyEuIwDdrPUzZ7PRXwoavoF8ioGAFjlpA54j26RlH818EdLJBXsRG4id3DL5BXeLR
1MFvKFCYZHUk7uAgTwhNXqImOMqEDQbs9lW0Bdrz0ICRSz5rlugdOkX/YF3qZIiiEUJL+16GJSKn
1Nkz0slibaMf3ryUWUS952FtosxOdc1Plg/+KgV2nOrB8cdOd3U7Qf3pLnhPx8OoTmvrhi1PcP7v
9ZNbXFBs9VQis+QN7TbviVzyJHr5M728QUUFtrIRkpCwT4eTzQaSOJlsK9ea9/cKdDpBIDs1IwzX
3xEwZa30V7UOZqTMFld/JPTLtbewVTBCVd1DtfuUhE3h7Q33ubNdj71Wv2g8YQ/O3zaYXk21mhYt
MzNraYeu/MBpeiXL1PRr8O+VHZpCE/ixAP7OiGVEO7x8QJpv8RuAmpBwFAczhSnYKsIWdOL537YR
ORSQx8p6y36CZZePb78FkwFwNYUtnKzn3nbgHSyIvRhSwN/AwAn1MeMmiY6RJySin8r9cTE0cp4P
kLpABu6OXH7/Yhw9bEO00YkG9uaOvwwdL1V54cNF/XuXCZQxvTzt4qvZZUfHWWGmc7Vr6RtbmlGZ
gMgz+U1Y56fwBmU9JyW0muzfwzUYvHRfesJUITBKR/0Itjb6c8ib65wELS1Ps6adHukdgawvy3nn
HHJEyGKs0avNLVCUaqesKvtZJmlzwCxYUczu8XLVbjQc+8virEKYr9ZpsbGPKpjHy4wUbwbPmcMs
TWcDLhw5fFMEqphN/6NXaaFRd/8b+wDgtn2mVhN24ewQL6PiT0aJw3gxihQEG3Rz9OYC8/mEAChh
ZFnpubAowPV0Fyi3Tq6IZiNvci9DOPy5pz+tRu2FakB52TLsxGLJfvFsobJMlSYBDLDQKlO0yrfz
Rv1qxzxoc33eTbzzlAZ/p5O514XiiR35qHJLxQcxoKxbDnfSEOgasyIFL9RD9rC58xAnNKNOB57z
9JtmTIQ3kVgnGuzUVuOe6D+gOsVKrPTiSvKM/9S+anhwzuiiGLCK20rltLHT5TnjmACV6OHzj18i
nX/CnSixvpmkuRLk50GDmXY4bXnGnLAB0e8j1tUUlI4rxZAlBsRCy8FNpIckAAcjD8F+haBdnNsZ
dRP5SB9pxy5HJwaw3oI1z6vX4J87/bRpO+F/eTOriMb9a2p+5NjQhFVhNF2Wu7H0+7dg+tRHl3rb
cxRpvev7lsGA32tR7iZ2iZQ/8ibgxr0sKEQ4ku+CFZlKbHH2U3/1peEULCOA3a61PaX/lh+rFrBj
omvPNAdAJVFY/uTavZQpY5bx+2fzXHZFABxnlawMWi1VeGNHc82bXbXGV2R/qxEF8RNGha2kMyyh
PTR2mTf5yT1kSSPqupjUOw9WRXrN6/7e06eR61grh6udic1p7ubyCB7k+ZGEnNaRukkRe0TZmCy+
8Vxfa7uj35oUKLpTGhonsDuXbQi7xUF4miMW3kjYU4c56r4dHH8F+9SLnzxLaA60633UBj/+HnQQ
SiSTITTQoPA9vuO2cfUHfE7n9WAFzdw+LuvaxPPIadIo0Vk82zi8L4X9Al6bRzg37PflFgskqQXB
hVJO31EDrsOWoRc33NfMfIuD8Ah8tk+CS0JnOAa63qGVnmEvYHJ+AizoSEF90nsnOdY2Eoa/djAf
+6cLNl6UsIk+VgM3xtOqRe7QKRzmY4GBRgBJp6Vt/DN0jRxIxOeqE93tmA70SqI5wKk06IXI6+CR
gEQgxpa0DQK9YfIPQO78zDJL0gHEuxiezW8/aiUAALRbuqVtoDmBuUVt1cza3l/APdBD8Jdpam9r
YlAbQZU+h9AeRqiAqSpjEw7uIYIlZ2YWMbxQB/wNcnDYCxBc3DuiOn/Zo7YdbNigSIvdW5lw/5Rc
3/ybvXzvUnlTsSZyEKFWg5LOWSKrApLNs7wAZxlqGzrAxmjqMqZUB0D3DZM+PBHAefgvGQ8YUtCM
omGmIyjzAUldlDUC81iAAuEYi3Afjb/K9d3Z6Mg0Zopc/t8F1EKSxx7HOryhkoWnrZX2DMRgFByA
GU4aecLgWYoxIW3puTxlw2quX3Gx5+zlxKfD3rFub5yzItOVuBAMZzbNKWK8v3G6mItoEsPJYjnJ
Nbkhx7vq5vAGrmlrh2kk2rDTlLvPB916ULA2JJfuxaazFEqjrnhtl8tL2sI0tR5mKsf+/DDMIgbt
dVqK7715WsIQdqKBKpI8HwOIzHgOUc4mvvJkmWjvGoiQ7Auj6KjHC2X+dCKLxAbuvZUx9YoXEWRo
7zEK98OzaXSes3PU/tjMz4gNj6+OwIWZEIX2q0sGAQhoM/nntmiNRFdcY2h63aPts/LD4zJNVTKK
++upKM22cGMaYPAZ2lQUEvfFqQO5jKeILQD1gYCVOMgvv9ii20HF1yUHGUOw2FWymZehVZUEnFbm
zhArm2M28prDmRxEfESQ2TO9g+hJE6oWHa+UB0f0iJIsl65+7F79aUl00Z3O8AEmf/bCNTDbA+Od
H1ltrS+EICMLthwooCrDU0P9iPerEiCIH5qRBIXT2OtL5xxq1ETftAl0hPH3BL9/wdstHpsaF8gg
033ui9cDSRA4r2mn2SWzvAbuxbtzVLhTn/u1MJLnCxMlqsQhfM2KZ5l5e7w90tsdb438wc/F+Ij0
sZEwj3kIfYvq8hHBwbZYh0nOaQjZM9yFWnip8SCOLrRW28I2yBZX53wavpyvDOkyjYX+/Svhe79Z
wnvsRYrO2dwSTgHvFHuIwJCl2Ab5sYl4+6j3/gTOTM4jPCwYw3HVBsqJxJ7KYg9NVN5+pDkiA+MT
AusDkMLBRGTwUVz5LD3dNN3yE/RMiE/04A0Upja1iuK4Bnocs+zLDIv/q0L9cs3ozd8XO5LiKTtG
Du0AbM3lCFV0Rm5QZ4sIslqc2rHup/ywP0afmj1Et181TPsQGMw3BvP4KZXtqv2N5/2SJok/NN/S
71x5f8pSl6BSdzwD2WbdfFQonqte6OGpclRdfQGubrdMlLhFqork4vPXUPiK3tiqfyCJNs61B8IJ
ZtbMMUTUbl9crItp/2GpT4aaZXBGMeHNPHnEmzvG/rIViDy8embVX/FqQ+g6DOefQU86h+zWdTK/
zu1kTrF9KHNAcPX9l6dIq0wmGuXzsOxqPtd1gKhGrl1x6Q8M/a9Rb/f9JLlSmolTdEW/CD6TGh/d
BOwqzbNyvS6DH6APt8pHjB+O2Pdx1G2AxtvL2p3BNu0ssJaUiQEofs8Qw2ZxLTl7BzlT8HxVx4A2
xqaMoLw1hL6HUDxPh38TtzhPll4XQjq62zsJH/F4OYaBriIKzAT2S2QBAWVEh9wz6FWVVe1B9AsI
HcrO5hxkPuxU/ZuWGppN9YbND+OQ7n1irdycvjhCLD+c6BQ+V4C9r2XrJ414TZJICWSL7R1koMnT
gsbji0SgTB/He0LMgOvy/Zz+ZyWtd3Xqmt0saw9j52PG8l/2Eyqa1ZAInQEONmolmphzBPFivGnG
nBR8tDP9Ryk6+UxmNC/4qMEyD1/J8Ma80Ic7M711ye7otSMZioa+/oNtowbvJr1FG7wtILRN8hoc
M74/5JgtrV2+j8F/SKXHaXpTJKMiQxph7q+cY6d5xwWyn0HMeu5JfZkyBHjZZP+H6sZ/nt3w3K9U
qYSAVIcpxtYobzr+/EbqVC83IrbPRFYNKheV4NOtDLIdaLkgoJddza/TpKv7kfHDVrMPH94BiHhh
dz4pLNZuoHPyk/WW8OzWYiANzQbNjANhDofKkzemwUf7zw25spsqGkBJv7QlxarCf+NdJM/vpMXj
QTt58PJuH+yPvLpTzD/NJBjeKqIExc1NluvQKGdWAf/IV+JKj2h7Q6oXv0c5XCZvm165iafxuavi
MsqwJyt0ujhrnwZEv7mo5lnbE9rlMPBMpO5es3M/VphfS4x+dzx44WTikmCuhwRq90NhKqXdVDqC
7Yflm4z6ZSi64SiqwjLd0KTrswciCaO+DYBrOhBFdBnAZAOjk7j5132XrKmYVQ8zOUAw8A/GBXfw
S2E8hQsPcxlAkyalny5Y0TR4RbWLV422JRLGO5l3Uve11OdB2BOKz2ZpZ80umXVpCGup79oSFLi2
ICUSkN50qr9Zsn1zsKYBUM9r7BZ/QG78dTBO5nQEVVqNSpHJP6qyOB3XSSUmjtx9E844Cgg2ujTB
jB5UUkKSWM1bovkKGaGzYIbx/fX7YZ4HlbbYNz+6sUfUC1Uq1HQyuZQUZ5JwwBzVgZaUFUNykHG9
Tu8YBQSMfYbGaWGrtSVm+UMhzbuiZHLUgfeRjWeHLJgGZyHxlCEqd5Sp77moAK7Bqhp2umvUAZL3
o6LRnvxAvqAkSRgQbrrfxBzpKtkncn8MUmK5/CN3S1XLza7a5z9Cl5Zl8AsKn2Ptu8RytVHEXyyd
AtQU2PWg8eLo+lJyeBQ6gwPouV/LpD+tkutNe9lm7kI7Dp8V7s2+ExaDwtlChs1pXlNTTV97Otzu
v3yVIwmLWLixKBD59myBfHrNE2KRuXqADw/CIaYXfOPlnU25H5PAOIyiTdDjtxWiGf+8PfzbzNvb
GLXWepn1jWvtPdZBcyZLo9vTIu64knKKT9+kaYvnkAb6q+2JJPeVRWshZvgLgeox79jIBEFxbZB/
kQLv7xHp2ReHl87HfohS4hEcrmOLwzltPWkriVoUkbM4GxXtwVtRg7ZLYGlcemeV6n9lZosn/9F+
2JmjaEPgFMZTSkEAc/8oCpcaxAvpqHKTpsiJcYH/ruzXQ6tWoQ5FokK142OM66TrC4mm7hX/iWM3
EnU6rXJUVtPkvSAEn5WBpDTTmOH83BmvT5mg/5676xU196MQJgZazVus+Rh4E7tMz6fMxHLqu96X
oPWE9JeJ9WUCVOvxw0YNsnWFrDkBvLeumYyM8dddS/+S5ucMxKL1RNReeVNQjweB4KcVHjvqq5B5
WTsdsh8i7lx48gTBKTfB60wtISDyS4KuL5ZwXQOo5yzp336LfWmmcUs1UuGq1jLnj8BmDv/+H36v
5Io5UQzTjXmV5aKwpIsTWvVmfXCuOnHW0iPyYCN3BDmuGIG9EBXb+MZcUXqrRCDzdV//f0LJmbcp
OEEqySB8yjk5IF4PxJGevmfh8+wio7pXXgi8tYb1eg7rSPklw8NkmbgP7YZIknUQwm89VceCzRzG
w9RxrhzBY/VT7DldHtI6GS8qT4OmKKvFgxeujE4+zjOp55fmEps1EcgVMmWNoVipptUzgoNPpp8w
ANPEH42P90V1HJ1iEq3r8aDm1+gBylzy9astukzA2v30xm3p7UQaQm8m0Z/PjlZ1zAz0ZIqmRn2W
KBhgg9DsGhYdYPsr+7DxOCoCjH9APVSkpBbqme0I44vHYnk8/qvhcKRFkPggrmS9Ib7EnR6z7L9b
reodTgczkm4qqXT/rUSusJk63XrNj64SRwpROH93B/p04nSlHNIUAfP9PfDHJPpCpDCFTFAVW2Jl
wN/OIeCwRYjw0L0hIqZ0eu4Ch3dhFm044SeKZjOd1xC/lStbP2EwnxNxUOLSUhxJ5OWnRvkN3vYJ
TUeSGadzupCozzYXMvwjRK26SicJLMiFGQtRW8MC4McULX10UJy6CeBo28vJVH7ZaHJtIgs1odpS
lA418uvcxbsJhdny3eCrkFhac/wXxLVXirwwBrVTJGcmsIpSVxQrkc+AtEgG39cH/48Qy4SN+jnz
WQbT8AkLq/Axx1M+wlnO6mn+sp+9n+c56bNyS/+RWa/n4Z7Vl6EmCTmSwmUAV2IQkbONJZfMOuO5
3nRlPckqyo7RNZXZNJ14biOii5E/PvIMrtsqKC0mjvOCKKOquFhUZSKGkyKpXqvaiLX3ckzeg5er
RTaVTU4MEdfk28Bl5ksZQtxDHI8B3F4rVaRLS2EFtHBsGV0x9YRTn0a5lq1rydLENNqddaHMquw/
AI4Ua3wemLg/TK/9DAUEzMBu+5djgMCGcj1eRzMh1/qw6Ztrn9F32F2yBA65LbWWiZAU1P72XwiJ
hm3SwCIcsuqJzb1eC5VXz4oLLsvVtW8TyitlY82JSlHVNd5GEtDw1Ad7IQ1KdvyqQpieR/hQo3LJ
DaxiUysXWeVvFoYpeas1Ms+oVVpPyo20pCRfLZhBgMnpL+C8bXGFYyCcbN5U3sjGxMWTn4AjKuit
P6/t93CB8UhArjUJvuB7cDNXEaXigxdt5mC53qAEukooid8BPsD6gRbhBOjAbzwQWXrKJjDoiyPn
E+PguTzCyvsFp15uKJFkOIR8ne+XAANQXlruEdpiGcIc+Rq4XY39qG7csHUSUU2yDaaXYXItnT+O
Me747pmxnuEQMj0gSiAbZBM8xYySRZEGATm9E/HX3X2V06SPbPdJP/ysul7Wx6PINTXJAuozWzaH
2HfbgDwqT10KrND1ZB7DqMTzW9hwxBQYFc9qUrk/rj3J5X37zfrYmVhGMBbeVuShVzSLGN4C8u81
PNgcQ3kXY1LzkUQhfgkJMwzayxuQm5vIGc+cUvpnQs12l8BmMccMaieoPzZJDRtwJ5Y8ixyYmt5t
ZXBk5wwgzfZLsRx0xSUJmUUDjp6Fc6pmsmPgYOSim2xM1mXLG3prf7MEMggITr5Kh6n45fMEcYIN
InURS6plG3YkReiokUi0ioyLQ5oj/VBiUYCjBQG3XhlXgNkFHt4prCyXRNK/ul7Ly0nhO+xH+gBK
wwxfoYgjEVHWZfzvG98Ze/lR2MID77FqjR8DkN+6PyZe38sGp/NbQi5tAcLbXCWQ5DiwgcVgD9W8
EmNPt0Cq7qn9pJLh+8Dv1WZkPOM3APX1Xt3nmwcxgcpxSltttzuxxDBEGbnHuRgTCynIlweTUk8q
kphM0dV9rXkIiEPA3e0wQnEesDeIZo/2VC/cT91IEYfXZPvUw+EF9cbsZFh6xzuSEG55RzgY0kiC
IcHSMoevFjH2Isi/9jAFqKynSfs6zCjjf46YZSO4D6LxgVRAWn3WwoiHDK/GyCy3H+nLw47ctVHc
9BqqYI14iH6kL7bjsnTBSNFeEpP4xA5TlxiFc9P6aHHonnM2EdRyDcXs1Gbt9PHy5LvlZ7lKu376
0WZgU6xqAPEjPyR/suCpR3mRUi6vAnwc5dJoSrk1BJoCDv3C4Vx8mSPn8/PkM9l1MQ9apIZCh1s2
UIqQIq8f47rpX7jmuto4UpOYoK269fb6kZvkrJ4FfUPHBnQFPBojYHsRzs0s1868t4iuwoGW0KkO
fZb9xrMjrLHzFz6MZYYVS7LGE7aVPGsJeM1hLl18Eg/BczxVfFuNNwaqXTWH91rrIPmmreFWHSry
3hFfKNKyT+laqkZCF4lWCIRI5b47uPXTiT+4tXCvYuM0MybdiyI6A6oBsljX7NPLxB2GIg+qWInN
nZ83rvJZT0sStimn/hmxbGK9IASKn+QH8wmJkoVwLcKEzwQ4R7QL1LjX+mJrTcRKnWXuJsWKFEum
lRI5URbt8rb2b6q2rdOZ/G20KeL8Xz0ohNO2eCBF0MuXXb7idZTJ6PXsF90HeNA9C8zqbckLu1wq
14TInwXzkDFG8CaRVVDPcYrh4EZqfLx9NTOZfMUoHN8PaOfx9Puyztn8/pD4cPO4RZP0FKCeMF57
osQBcQ+23iO5fgwOETxOaXJhm5PGfV+qC1ge8JKB0C9y97Kvr7BHAgarEfC5uP/S4Evcn5TRmA4x
Tz7X7WsAhgi8AyinAOONXkVrVvY7BqJSzfJ/5PZNnafGo85c5LQsfYPcA9heika88owR85jjFwzn
drqkl1+G4eiTNZ+5yvawc0c8/hW1yJEpAvbcQniaKfRO5tLXA+w2+NqI3fi+8gSRB6wO49ze9JlN
R9Mn0HPHBAwSZoCFXRmM2gCz5Wu1KBvaY2odokNqxJpGNyefonLintxUiCQV2FjEqbM0AAcZvMj4
H0Gh+dIAk+bqGqCxN0wSKvB+SeeJsCA+o0pg5BmoEEaahobVUAp6y1L/kc/l/PZqIHkYDAPOIwpS
I65Y+yC9QEVGqWvy4rRKdUp3jQyaJWDTF0nSxGNFs8GFCBJT7rrN6WKBa/zAsUHEBnNRRdsIBOld
BwJBkGFhA6JQrFkNN5YowzLsknzkuiZ3j6pw1R1DZW9l4vwqT70CL4ZjsrQBugYYacnd57DiIx7q
hNhUJfNhM5M0wyFgjarkkRl+J9YSCAH+IPN3hGorprA6u15h5P8FClnPC0PdztArJ6dJ8vTRSDu6
DJUxLhWwjiBec3PC/WrosTt2FOqaXpIvpmb3b72JFdj8v0t9jrId4EjnXgKAeAuBvP35zLrh26jR
xqPcw3fTKFhIZO41+xDYoMAm4dJuZYVzrzET9omnELzzBU2LnK3YUqJFb/EoHU7ihn5+T9cS5/sX
V8B8rSncpt+MIaUaUZ86sdIJOhjzCwaBLy9gjSJYso9fbYvts25d3SGJZASLL4I2LBJddDu7RTYe
mcETtKd5wJZaXtJYwBIZCCfN5tzdjF0JRLUaweJhUUSKfRFkA4Wd88THSXUOqwfhZwLEixg3uyTP
K9KsSI7Sj+c8Qxx3OhFQm/xAZbXXSzwMAUBfYMVine8iKIO/0k3D8GVGeeSd6jDK5ft963o2Wwl8
BEEXb8fqe1dMeSGtbwdP4MYMXHDP0evenv+VKVHCuajzHuVOqQpZATZ3onMwMqVzVGhC6g9J/zXz
lQfJykxaI5IxqNW/vyY/vAi7z+J4uNpcc0AS/vX4Y0a3CqwOh4Xqg1FaD1xCd5GBaIIbOl4CLh9k
MyplhVt8CsmimQ2cGs6CdALzr6MKwLqFcMZh179u1W7R6QSMvBRCgOID/y1XGX3izLZAJmYQW0Vx
UyMTl0Zyrp1E62aUQ1gmZQfDAJUE9UlwcB5HiKXayr6aOEP6bU+l7z3GcxdiUhgN6Dscpk+Ea6bL
k+bzAdgSlb+vcWdN489J/NPhYISTTfM+46SGAGs0TgMNu9qdZB0BiZ7+pEDs1ZZf+4XBMefEmYoL
iYZG3oMyZgI41NqDxrLrO9bCSQZAgOjct7LYgGVRHZ01WJxpuTIF287USblgS9VG+2lQvbmcEH2t
jSCX0NNS5juRzitjPo52A8/EErzTrRsCxr+cVA2lEeFfcgUPtdCEIHUEQarvJQf3UQ46o5FYkEAM
eRvq970VwSiuzKI4wNaw5lapX7ofhbcISFTQw6+BHJTKz4+/F9utrqboot0wrjwCng9j3bab4yrx
F5KfP38wF7EpEsE0tgWINSaTu9gwNlQBxthbPA8G9KFN8FrvfSk9XIC+L+essGJ6NPZyvYWbxRUH
FdEm9cjF+zoSkqK5wXzUg8bPycLwKUhvv9JKrWLdgsEdWQlN23AhLA6Tac1gEXGeLwuYqYDhkP36
FYUEVoF3iyXB9SFQbyL6Ys/570or7tCpO1arjKvvNKwQpK5cavftPwCFbvm2f2bnWMtvg2NqqljX
oAKHyENr7xXZ82r34p2Ne5mH5551q1UqDppcDTaKQO6CkzeVgCaL57tR8tShlzHTWD1mdvd2g7JJ
pni79PB2059aBPG3prtYzfDFitbBN3Efg/3DgPtiBR9zPOkYOvMT6d+zTFtJBOiohBKPvF8UteFW
U7K2Sqk6WKfi5ai8APrsSXFZ/CwKaYCAXGoUyqn1h7qFnGEZ2aA7v6oJ/+k4koPGFDc87vhZ0w4+
tt+1l9R1tuAVKbt69IvfvL6ribzZObBV/RKnnWfCeU6rmISf2/gicqfZxGdLa2c5f59C5zptM2Ln
Bic/yvPfwrdfa3iiP3uRWcVEoMic2pVJpUlld0FPXyZhjimIKMOjBn/QKkZymnrrMJq/u4UmabSV
qxrUlgYjORAyPMLd9G16QQipliQ5kV172O4unR2O7nFnSb8AHGO+bzWeT3x4pqaR2sA3mxZS/96k
Fzez74K+4yMGczb23SUU53gtN/2/mrbnXLpcrK1o7E1cUvfL8RsjUojL75ageDP6MNseVHPqWtaT
KquUULmnrcJigI7An2BZ31ClPsvT8lpwy/t4Lbd3wTxrtT2oXzrHsVVVKNlydwrHqdKgvsFGWPnu
brLay9hjSHbKpjdASdZsaO9dFtSCADukeVyhDM4hSEw3MAN1j2HIoSQ2MIIucw+nOCqr0/uuUTv2
c2eBEraWi/Y++K11bsOOOLtv2h32pWU4gwfk6scCwlspwJORiS9n59sJNd0SJlU5vAof+/UoUmTa
FLMEqnIeM8gpnTKCg7pRwMWnxNuPipbuZQyslDZc0Y38e73RexWsf+eTnOqtBppFIT7mu4azg3fm
W6W0wNEPRd8JgiR/0AbswHbv57mq29oXSVo6FKOyzIYGhrl5D/rr8kGlUcV5Z6MKyWdPWSp2VfT7
0+66FO0PnZ5RDPgTtWgerZJELVOXvgLqxhYGiKGvc3JPQWPwnQtmHmkyQJLqCKEP1fc3ecnaiNKL
pua8FLkGkqyp/EZFp+DrtWtY4+4qrCyp4iUBzWeutzPCRUbiEqp28/4RUf6pRakj+jE/KKOcL8hS
PaZk0XJ5+UGnwvQFWhXsUoAQvS5jtBX74x1abw3eVKZYOHaoifJOX3IdTf6wD/GrUuUQcsQ2guJi
8UgBAjzxyUVTdVfylF619RlJ8N0cp+0X+HT8c9tjuyRfih7vzgc79AesbXefa7As0sIEYJfCFyX4
LR7DgU3dKYp23ZqJ1Z+yxtfTlYVCYHpNe7an+BcStkUddmbOy9+mkuKTssW+A0WAcpUIAcgIOrXZ
6FBPw5WgxD4cpuFXWeqNpFk2bembBiMZUoj65H0zLGOBj/ik2pUl6iVXUHldRREsJ7pKI8DF92pn
GBcC4TayF4xh2LANRQHLd+Gx+X3NbPICZfZ5HD0hOfSrGtmp3Xl+By19lPrisDRI8MBt0/A0WuzW
WrsRjmggSbzj6my7Q8uJ2WHzDsP9mAnzHQANV7DkzwVIL1p6UjD/kACb8Rb5y+zSxLvBdEK4JAHM
qwQzWrmM4oRguDnNhnDRyu38hD8pjDQVJJ4jalJAG9YP9vL59mNT9F2MjqAG5gMFON6TtiEuv4uy
E2vgh1jGXQF4G78hS91cyj1wadNPdXu8wtVnaoRxdJRYFgVi0o3zQuZYzGgsVEKEH7+onATdyIVe
bettDkKf9+oaJi9z3BwiccCoOBnKFBeQxGwskmGcRz1FWLtnCnx0uLIlzRIdw4mU28UCnmDSG/6X
noNpCAU0VqbUJMnNfibJU8jFCDzHDa91XWNWaudIgvpKAX6PNQhQ//1Kx+zhN16YrzjX5dXlgIT9
CojGZ07UOTXcBkiXo3uaSLCEHjkW7bdxPcCeH8gCwn3o4m6LZB1GIDqRpmzqUKjle4KcUJLPSmPi
F+QM40d0GlJvB5w8TXNip4RaJ3wZePou02i8AQQV8oBMGf3ECFYfWBgnQHpJ4ujhZKYXMH99jGu7
cOxfoy8E0sG+dxfc8E6S9+WkyCWI5+paea8Fs35DVW1CUiFj+c4OTzzpyhXmmwUN2X/h8qfZ4koK
Pc+Hx6T/HD1aEjmCT/04Cjos1Nn7bQm/JD46Lbf4EFpFYe986QYbLyMrFn1q3ixm11c28fXzupMD
54xh6AidiK24vZ+ew9IssVgIZLXfoJEFs/Bu2yOx78S/OSXLjER05FNSMoO6rvJd5zWQp5vg1J9A
NVQFWvJY0bGCA/HtcMk293daX7x9sTp4qGjPtxLllkXK0NKedb1YDB3zQv6+gautAyEsUUeIog1M
p1bPm5Tz1o5boJoZs+xF43E0LNGPyVhmT7JKfOCylYBcUOgAPn/cd2CXXB5l4cdV7CoF9ZzEGl1T
aVKhNCElv7vnQ2jejIOmhIyocGGq9SusUuniD4YHSRvtxgztJkuMyRVUT8WadQpjmUdJMTS3/lR6
xm/KWv5Ojv8Tg8N3BjcxsFfJuxSMCJas0/DenI6Z7fe3WJp3mB5ePhpI48KNxMCl/SvI6bHi4uA9
U4DCfeuNo4mT/haNd6rEYLkB3eGAp2w7n5bogyRG+CxNGh1o8EhfqnSQBgdZMZXuiCKILRT3Sh47
PhjHjH92YIJmF7eNwpO6OLN2e5L/Oref23qN6nogNZaPFAcIHevEcFJ+6BDlF82u3c4B+/IwAP+F
Z++7ptroOaByO0xhyzGmAPcRDsq/fCVthfB9gQpCExm1qUfsMTchrZz9wn5XwpS19zIP0/DubPbF
DplAqG2DETipggdWnlGhmE5WpyiuFpNhDo26Q6YnsDEaFPU7Rqzr72whFBmmrKx+zHBJICAnZN07
iLiCVYZrDCan/2v6RqKiyw56I4Z7vx+BSx1cdwl79IU31HpEDe5gs9TH13ZKFACbxeI4p/p1cSI4
39xU9iVDvGgQRI0iu7XwZ5buiaLc3pTc1Oqwcf0E5rJ9SDM1VapQDLlwIW4ebA9X2wIfB1Riz9bO
yWCzPfzeuQycJnHdlcC5xR9qBwiecAPhk5sbx2NksFjDyYbWLjsfX79jci5jdTk4+BZxpACK6Kjs
+blZ7QIrckq+kDJTQhOnLL/rMIXNb25ovQMiE/oa/x7R4dp2wXr3R2fxDOrbnb9UHafE4JKL6c2o
8/BDuG7aYXqlbhsAMtGzyshfni4VX+VdvVwlW79OoxJX8rakkOtfdCQ4IDn9Z8jipiQ2vU0mn0D1
eOyyPomC+VubhLzz6yR3mAd2ypdd14DeJDGiQe7XDyY3e8CWvjHN6t5z/4RWafP1TVvY8CzN6zRQ
jPwkEKOp/Kw4vTxQy7bGUG/nYATyg+j5hBpV7bsv2zJS4RXUnd0WaGZVB+Orpj19hHUgLv7VP6Fe
9m3jrFASxZFzV65MQowQbA9a8OYTlOBX4MK4Cr1qKPdu86LwXwnPAgY1mTrap7FEvDbcZ+PgwhN+
cXR4E5MSgGPn781k/tvbRfgaOo8PaKFHlIBe6gtx0varkLN438RspXIovqNIoM9KV2n3HCUKk1CD
zO3ke1w+SDmwff5mCshehaAUrPOxebC/yk5kiQ9Ey1K7EYY7YzplrMrOJobuoVnWbLRzFooSHfnr
aepoast5FlOBc9KJo4BnJiv/BiWgAs9nCboc+XBkA7Az+mCHuMRaSXkF12Wht/NAUhCer29m0wD0
nh/vtnngG3bcOdUqDEVHhPKJV24WJCQ/KzvGXiRggA7U7uWXdyprlJnG4HIrJInia9UiyHXzRJd0
Tywi3fn/UQny2DJeuG/liYOipq3hS0J/zFFLYK/prDQAr/3ic+WWgdE+7+V/HwtH6xmJZ2fGL+qh
qVBWKHcixQBweogxgsfxvuddyGr9jd5KQ0o+zp0sEIzkSJx6HPeqNRRKyWGCQriJEN8k01xaNU6M
DXHFrRQ73cXdwNJDM2y2CUN6cEYZRynJHmi20iQzHmC46y5R/5zyJbwxR5T9Caew2L2vqeP6pwjj
JceI+ssMGr2ykZpdOxOH5r08V/xfw7Lfp41Wh7AQT4I1QFqciSIx2x2YDvb/BtOTbvukxUVw/4tU
nspcAgRXypKfBB52XqjJAotby1PWRpZ/zoidO611hZfvGAeINLaRaiqBZAGXFDev7ZvtShzA66sZ
SGdZof3lkUXGcnJscT4qPOKLsD5hmt28dX2IknXpxY0UvvPdUXd4nM3Gvb3dSGVfwWH4BSb8Ah+b
RZ9wx7UQWm3g88l8g6866XiGrLfeX2itLZsOHLiqgaOODZLWaLdhRccWZr0L7X0gzmjREjl2rsft
SWsT3h6cICdYUJ9TJbhNJLdFhGnFHpBzwk5ewSg+8QfCIEHbXm1QnuCfYJyuyxnfK+Gl1OPmrObQ
6B3N3j/eUJrDeF8Tm2FizXAj72uHseMaDK+W2rCRD+mxxXBiyuEY4zBpgnD0lJRIwpXnQzpkw5KV
JIG7feXnSVRNFUmuw1M3blB4CL2ZdGVeDOTFKwTLf+5W9oDnOP8Vx/t0fO9OsiJgSfUyZAWWD2Ar
icGRwJ/p4xJlZaJge/UEp8JTHKsGROIzGMSg9lRt4eGv2IjFm7uQSkruuP6qS/khcWPs+ZBpvR5K
rp/CW6QVJNoMTSp1WMgRVHiwhKP1AeS4d/4+XYSw5YlyWYhM4W/tTZ31Bd6qH929zBIG7DY5xdLX
zwwW0bAZqVKJj9nAwAohlEpFepzGxCeW35niNmKjfuGE3xnW3iLnpzyiAiVG9XTUBgW4H0A7n9ST
KRscgumQUu3Jd0hIEoecvxOmi8LrDk1CqyctzZjDU4vihWUD2X0ZFvfk35Py1B35mY8veCPG+ReO
BIPsiqAzliGONaA4l6FN57W+65mwBmNs5sml/6tVbC1EUIyRP8Crx+srBVc6/aLNF0ayxhMSn31d
n2g/gGY/hABJ22czDoh8N1xusNviHVWDCGb9molHientI+ufYPVFzD1bm1T0TbBfG5ly+b2U5LRr
sg8VTevMIIMHMLm+tssMZlTgOxfLPYUZGAkE07jxy8m9SgE05OG/RHvrWZP3HQhqQ61SnQ4sR9D5
X4LrkYVCmaYIRhvuRvYV6O87LSXz3plKSY+CRfPcD7ouF0QjWuVT655ElNiazSdbdgxN8ZI7r5oe
3aKLYHkD8FL6EjBRVqoFWca12LJZiLCMILgju85YKDZ4Qci4pTJeAYfNiCRggEqdNuZdshQ0uT5p
RwPUueIKN6GFpOqsqJt8CNTuz8JdTtsCuVZAXjajKtWwLHDOEa4r+GYs89DR4cWpink5xZ7EQ/9m
qsEqG7HApDZ/ulhk2dwt9w4gyKu5dKo1qfo9n+L10fkuE8p4nYfI9mjI5uv8NGR1jsTzdvtb0J/K
mrxBfl/dv2RtxdXJVn8pDS++WsdQcVdQhIwU+Bwn7fkGmQ7hFRmfwWK+dRkmnCJBxFyxfCunh8e2
cknZbxps/5zxrz/F8bcIbPlqmYlJYxx+rSgoTDGVCWtd4Np54ZVPTR2S9n2T1HE8x3jqXDx25h7I
174ZEACsC6TIPb9NH+djpoFPqxf/YV0dQl5VedWWl4H6qhNXHI61nYpD5GToz3oLvuG9EtPttHRq
v1LHrl7KiW6bx17y6+ztyfX12UMKxNnQG2VGy2IB0Uvd6A3S5vyopMDiwtcYdF2aSET+NGXljPqp
0r6mR82mdb0jfLdcYAuuTOp7NAye/ryTpXwVokC8P7lB+99h7Taj6GZWzf1eQSHE7knDSYQYuRSd
5iwwdNw5QM/g2VLMEi43GhzlA2Fe2j/9/dmQN+p7yUa4rWn7aXzyriBhOCd9+/u7K2o3ajhsFC0p
vPX8tmUQwF98nS/LbdBQFS+k3rhBU7+0hmuybLg39d/E53dYIoJ9hzCKnUCeRmA2TLSlTFntQWkB
Lfteq5X6acO2NUsNQzQ0nFeGBuas4/rjby6uPPiZdqQelipKZhN1E6QTzhnqizP36Zb/ogSXwpvz
bsQ3tyM7xEQpUAEIv4K8Xhtq43J0VR3SdOU8/yb3DDkZJQDU/M+QXnL0xSo7VAccQKL3yF198H55
H4F7ph0K78DtYjFzH1J4HL+a6y9Q+tL17i1ODKi9K4Q+kig6zC4W6sr0ry7CeccxbhHdx16x4buv
DEfKMRfEjqu0W73UFTxJGcqdkuYPbBzveicHWLo5dg4Ik8r4007/sUPpZitkfWRUf6C9NmVIGQp4
ELOYpycb5uXcSP8UWwv/BydXtl99zfDgL8NFchs47iiIhSezp/G2zHCQFhzhgmw1naE03OFNtTEb
VpHUpYByuKZ29mm/70ZdDzXazCV7Q4i+8j8mxIzcd7gSRl+pdxlraqwjxOF5q9fnJlxAopmZyM2g
GXfdCqQVzBxEBeN7WIE9/0Ul5hBFzxYNVgNd+D5ahfotCf43IzWB17FH7qVY5CaI/DsZi2jjvrNm
qwe5qI9/kP2zct0+q4R6qflEQ1boXrEUI5w4/2ZoSyPjeogiwuCWxsMSkE7iQbhJ7x5X0otZ2hnb
cmkZKaQ/2ss9oRSS3Z53ZjGGi6l6LNzXYGBrFT2rVEZmf/07yAbRMhkuR59R2UkVX+S1F0vnafK2
EY2cBoX8OVwiBab/fuqPWRAzOd6sxbMbZOoaUFDmH/oNxCVJD7ZrkP8xmAqCWTeruiX72gFInUqC
heVXqTab9/LxkOhO+9BcD3gl88uTtNBenWgAcZFytFEzdtdR8J2EG+pfrfEIcA+pz269EKgDYyfQ
z8ZHQCRyJ+Fitlcxhwz3tbYX9G8iokrU1aJxipQyWy1h3c48rK+HGXY89FQPZXS1fqQLwKAe0PF0
wOfpG6muEk/gvDG2DXzdGBNRo2F4KHPE9hcp2TFxRXLAHkdEkH35+xsDs06M8+5yA5j5WCCQ6NZw
aQMFwUt0mV+92GGex9WzyPyQtUS/rjZUVK3SfL/c1Fu9GzgNjb5Utg+I/7O3gQzqvEe78vVsWtoL
2V7OhdmkDZxSFKv4BtylBlAwRjlUfkPeJXXhL9UtK0o0hmFTiJI2KZ7KMM/SJj8UYrkiDGdM1p8f
0OuveKK2pmeDmF5OL3kd03MfCGQfhL+NOkFNlQ8OoOK8pmITR8hjqSoZLKgL7NfpQ1ukVbvjjBth
ExcSZ2XWI4wcX1aeG+Sg/Y93IgM1RP+2VQU2FafxU/S2rIXCvtT12hwObAJNywLs3cJqdXfffQ7B
My4N2Z2YLabC8+rnlLRgAMua5Xnr+fwtT53ZtDnBiHtXnLLaY/ul4Junk1+gtkC89w0c4aGQuoBd
Giz9eFSJHrLg5AxOwHtwEZljHt0+PQ57wF0DReqgcoRxWLzUVRgSzMWK4ZKliEUVHOqv/KlpDeHP
GXo/VN+h0M0bapjmo/k2RzqE5Z1zVG8PMPxjKmZe/IwgNVkLIyHOnZDKmK1qvarEVf14GcfeKDCB
SgLhOqTXL5fqD9siU9UbYym7mhmfnvQoYexJ9lEs2ZFiCcbjTlugsFKjmGdFyd5vw1nBL6C8DWNw
l+BcUp7xF3JjUtSQYH/FV79m8BiD1yowkhtSfaK8J+ANI2/Sz38dfE/9dF+jVBXaWtDo8xmWHpOT
u8ICHVUiSXY8ib+CUWxub0VPKuPdy5EIrAs2VrWXiSyhNoJt33qiptiKQFkTby5JhltzZ2JrVk4o
a8iUKi693UAAhxs4qafD/mUA8Kf1pZc+LcV7nqaMNn0Psd1kDn7q2OpN0iFiMYSLfyNwOE+4iNjB
hq7RX7X28izmK3VCdxH4S7FE2m4ymK8BLLM0oa1EFUAbUb2D+6Gdi6Vmd85KSDwHeuSygxEYSqyI
D7DhiCLbucmLr21mzHkwMR5WfZkv29NalQEDl7bmfHxOg8PaNAhCE4rD/YPFk5/Ufa6HbST785z+
fJSVnjs73dnkCeOvDi8nEeX/20sgXL9w0EBbsxjItyC3DUkWfnjXbsooxic/LC8si+g7/4UUl2fe
+QZ7VWLb2P8LawqhB2wx0RPGooKeeDBs+PAACetxlZ1B3s2/7puNyBHqM+afFW6Tvfi45ck0BUgX
iDZ9wOYXiQ9D3v1YssVfz6EqGB6JJ2Qqzp4hsuAg83AGAIdFiu/gficKyl2hks5xBDPM51cCay5H
Nmj8I8ZSq1tmpE6OLKnQwB8Z1LWFeEwJoJmSqZvAm5phKFrbe3RND1e5BZ2uDKhwQlSiXtVCpZU3
Zn+cvwh2kC9Urz+aoMBcf31NkwLlw5LXptCBSZkVjnSAFTV7H2x5tKSPEkSpQPMXlS2pjAVcY0a8
rpb0UU/B8omxg8TC2xL1Dw5sSG4BCEuCoppB+PCvjAk2eVCoN5NJ19y97dDhFqKXGb5kIfTGOOz+
PgD27P/K4KDWxgCYqADqOtNSvkda5CTzUkiLGOqs4ZQXZECSvUkUgi05HBvU8O404vkg0xOp0f+z
C9oMyTU55uLYTcWu0KP9jTUv/mg0JQIRAyPbQeqgjP34ucTk3hpW+8Evrz2vay4cHpU5V9zZ/sl1
h4NCyBIr9Js42jrc5OPBrgkjRAB1Qr6Rli1KcqqhHX9iGYAM+Mrwa/q7gEA6+0wChxydFXO+AcNq
zY1MNL6sGBPPKfR3vElpDdVOmoWRq1nRuN8bNnZmU5jhe4k34f/THNfogkdaPwDYSfniO2XHR7yn
QyXDVTAfd123OETN6utm80ALFCAR3ou0rgxKLTu2npH0oxd3AaHwDSwOEmcnaZlr135wRLd8UR7x
cFg+Nk95Tc68AgWxjWVQwM/HLthXhIIlW9XIlGtmJSQ4XOPOBeZIcW/ieOxAycX27/OPzA3yNytV
fOFdW7VBqAFboJj1M/JfzhsJClQ+VsL5wgznqHg1jge34hsZNT9jhOT1Axbq+RDodfM65uno0ZiE
wkSNGiavkJbdm3Xrg3QctcoEAl5WMfIrsgufTTS14kLrJIQ5NyRRAemHrRq/93Ee8w2bCHE7IxbY
LA1gjAbZnf9xFT8c+//DebKhXjqPlyiLWhbygbhnO6+AdF4/x2agR9BOt3FEBPezXaRcHKlCnlry
k1BSboceGWtS5W9S5rfmsW51mcxGfkU1bzUGdSd5eVDgpifqq1FK43VKMG8tWKjlO7UMkS8VCe9P
sbD1JsIu5ffINqY1qlJoZ96ihVwnYcQ4QxOXjSfMXIbD2BgKVzCRawDjhJhRo0UgmooFyMigqOh/
Vi67Z5U0Qly0/bua+59FWIm5AQo2NiXWIIz4rEcvuRsxg2hiL6pKK/oVnROHjwY4WB9/mU2ozv6/
ZnjgI5dcIfE8SgIOdq4wag7RjAMKYLjE4M/bUSJJ7JK8lpfG95V1zsJ+0FbNjLN9KqRGxefsrORY
wO6urFsdDBjz7/phzefZjr/qm6Yt+mx8ppBiyYJ2WI+OHw/3nc47T7wqRAC/sshuPRE0C/0nHWKd
wN2QnTf2X8Uwi/66wx8EVP7EY7vyTupSX4+tlyf39B5QK3kk1Hmcz+4zV+hXfcp28Jq0BUatkF7S
e8BKDJNRMFLUxKRX6nanV8oz5Paj86N+HRbjtMEHmLcQJzxZctkDpurPW6HfX2R09ocKEaWawDzE
Q+aeuSwdfddLsyI6UPRaQVgyAKDXfnZKrzGSZMOdj6IW91kyEoeb/eXEqjEP/cvv4fLj+ZE17DHm
hnH8ScAp2ZLCy+5BHBuxEPShHeWASHbqXiikP6VH8cnJxcK5Zn9hIgc+7KNxDEPd3B/DJXPmCGdq
/D9z3anqx4om49sBZjRQr8ZtUe2ZmnG1D5ggqOoZ2opH+w9cT5Sm0LoZ/vxK+ofKMY2rZES2eoi9
wwZ6sFqxdi+BFlA1WEbKFRAZAFGAu2lROT3MVzXOx1cnk/wW2tiikexYwrg21lBWTU61iABG0GtD
7ZOuUpQszF/U2Q9yf9Sn3r/nZoTuBALUk3i1HTgKLc6RFFAFKmAvRHdUw36lys1I4uCFTjK53SyX
ift5qDirhQtBNvyX8+Ir2j4VLRndJov3vcdlk67zmeVvgTVCq1OMgZ4D9nr1CbyqdvWnuU+vJR0S
NC9JZrJ7gDyUVQX7zH4HY3v088M+XqL3XwhQ/UTATP07iaw5TiKx6SYVo6A6RhaFO4wVX03wTd77
eUPwCEi64lOEhRX1LWeYlElJKmFG0dqAs1vnn7xwGvlsFhycwcPHoBvHTTcUZv9L0hwXUIXmOnoS
h5QDlKQpcSO13t68z1kOPfbVtDX3bKe+1Bzhf8HN9WN1VTmUY7ihYrpjlt/zGlau8T7lpHc+74Hp
ZBKu6CVpoBdcnEx+tTq0dRLb82dmJvlsPQcqUClTKnrDi+lDi4meBfyyL5OyFM5sUz76+fVUtAZn
2X0dhw28ZWFyQ/a1NAEkg1rCh64ss4AA6N8rf1RLFJ2zy60jBgyC3pN0CtwjFMc0aMv8bbfTGY0k
ZAsegjOGVAxWl9f/V2M4c1GBoIjW78ffi1tQ/c1RNB603gAn+iLokqEYi2U7cYOHsmGMfPtyV5+u
zb18F5sTCcfzMLS5oVkC/Ne3WNnPXY7U9eC9bq7FN+HW4kmdjw2lD0eLBmJfixA5jrciNMj6SXbG
XW3I8ZokMRzZfNRFVMT9i4He/Blz+7y4No8Egimp0kN9EMId17qAGwphJYokWrt5Jj8aktfY75UF
RPgnjfR8+yac+pXO9Qq+usoGxAAKKld2F4i46O7tDiPuhrLFoLXAzbfbUdGsTSc5YmWkLiREvhhB
W011OX4FJBEJuQ80mz94otwEVoYJ2OWUaX1z9UYJwU/w8w2dYUxG6vVQ88IVd7OfG652K8TJQAQW
sv2qYxGzdYhhHGLF/XaUaj36625SQzyWRZQRjgD3peakNQhO8uA/r9SphWRFclvSscEwHB5xQ95L
Xh620GmB13Z5Puz2NuxbCMw45liV9jyFo8bjeuhPuZECgE6WpvizzlN5RNmGMr7Xizkk2hcv4KPo
h5IZauEuENmKVvUs6EUTwm28dhDWuUpupB6XkXYz3bSzZQIaKcXmilFvxYbtEM5XFIxApU0V/62O
78Cfw/i2LfWTQ3VAIeL0jrz+jgq8DPpI1qoYk16/SCAK1gFNEYp1GAkLLX+Soi55GdRgqUuJ5UUL
9NvXLI5Pdc+AvCVSZEG98UW+kT79CL2rH+LeLVPZly+SEZnoyYhjBlywbnEjv1p0CyREoTM2VBxD
/Wl8cCMp+sH8PNYmXSSZG1rS2UkYBLmHBiKCNHaZIpFsRaQPUvR1//kvOLJcaM8kcRQq/tuGXc0O
Vp+qITujzJ//62kprbHyDiB//y/ke33pGAcrNC1aoWwpMqaF2E2eSksLsmRpBOh2OyeaBIIXASUp
pOyoRbtL2suFMAW3tvuN/iBhqmRuupdGJ2UZECssFh4NnsCtz4YbwWsRK7vxCyUseypPZ5SA3gt1
lcJ4NiehS7Ix2bdONQqY8QHFJWT3oIYExxalAnovgvUodrG09DLbXuVoPJupGR1BdA1U+je3vc7s
91iYL3m18Ybb8eiAsnBim+fBMbk/47nK+DU8q1iPlJ0MowHpQD42XB0dBMnpa2EzfzGuNu+NcZC5
QdKwn4hs+F6DhlyvhEZhaS4IQCUSajGTBuEedepeswiNZPYAIpAyr+oYfkFJ2JtWf5HXqQ57Gyub
th+9SiGvONmEpY0rAHdHraM8r1xBnrWqLp+zxFfQNrQDzbMAzi2m3fvhNJND1UyG4WfWxpq+uC7q
keERLuf93URxs0+TpRXwgzJQHoFt5N2Be2mhiw3Pc/ciQGtyOaOVvRcUcgSsXqkv/HKhWcfQ7wA2
2Rxz1a7Cmmlpojgei/KsDdU2MB5m9U/oSaOHQtSQZ/hRiIn/xkj4S/gE3QtktOUSJYQ85IQwVVnt
SUyDIT4uw9bMqMwo7jyLVc0uTgpqJDu4aYSXy5uAXBVO/5PsyRockpGM4v3PumhMYgLsLA3QnmbO
1+7SyKNhhkDIMqHjhccbQNvJcs9fYCkxLC4r/sv9i7wMZLVrFBv7BcBVcfHIRUdn3sYVDhW8UZef
K0sOB4uPS644rr1Jxbwa5by7AWOP80wzPO5xIBXoODHqZawnt3CabPKjFbmpeiKGZM7fmqvsYGOO
dcoQkiIkUH18aFF3RFH4ok+qYnauA9PLf62ekzf6oaZ952heBu2oED+wszWvq6u//QVKJsz2Si0p
4L/siTahKRhg/bY6AOUJ6F08LD/qdIph2Ak9Afd59+tTV1NYkG5MwuhLDrbxGai6RVmmuv2Bk08n
jwQdWa1TXctfJ0azMajP8QCY3QI10dIs/4PVlch4r3AOmwnrOx9hOnveHdtNcXKk9J3B51BoqMlN
tEkR10AYhE/fUn+Fq3Guqn6W4lNJoojKlNOv5gUrMveyhQKFH19rUDPU8UnwHZ4blHIoJ2qxvfty
UslSOwSshcQ5y2p9yVBTzUzuKZ+8NVlESl4zm9GtwMXHpo+9r1PFyMyoQXHQAWTbY277H1q9G1oV
27825I49gsY91F0uzDbSLMvCgzdUsLCqSx2ZtCloQhirzB51t59Z9c6zAcbq+tQKfWjVMzJT7VOm
9QA22knk0VIcn2X6FsNbeLpz4bgI48u9lzyFlDbhngEx3YDcLxj08OG12S/vLfYViv7LblRS/v+e
SDxlnDILd6qmHq+S8lT0KwzYAniRmcbWPh+aYbkaGHpWvRXebo8+PdG+q/eN1Tyae+WfGRRaHwpA
/8nu8JVc7Bsy0qVn68qC1TjT/aA/NM4FpzFloLd7FxXLQrsBLmRSR7+gP6fgZxysCcnD6BvClGlX
o2j/vV7tLXXL7K9xacd+0dKRon140xNRMXlQqbdxyxKs+ej5hDlXuF1yOlpRimdM0WHvsXy29e5Q
Gf20we147upBQ4VlazeQUsc2rx1J6WWayJWVGzI5LgKScRQ56S/5Eb91MWJfszK85pi3AJ/H37Z4
GaCPvPdVUXhXK8sCJiz+1rnk4vW4fE8sQb1G/2i9So58A4niWGOf8rP4XnH2PehViRABTCfTh1iO
oCmab1hY3xFbDmwMqNE9PWr3JH4qYvJj52oj69tfewA0Az7IfZgxToe7QgCv20DhcU3N8dCjNrZq
xsc5fPiEM8xsb8EmpaDi7B/dHJwJ7rjyeIK9UOitYnzt0PTQrchQcpORSK/vom9LR5TGpONuYC99
5rXp25RLH7UCjTcdN5xGpO/bgAG0lI9tpmfLwiHiEPzP/jHc3CCBT0XIO+xlO1yWa46Afia5ded8
E8pyj8O+AyvrjdMzQrA0rM1uofDzwJVoJD2z5ivONYpvT4mO5KoJWjLmFKEQqvaOAS2N8Uqpc93V
EDLanIMKiyh0leSa07B7IuMaAihtIH69TycvXuMZx4tVHu2++sYGQ+l5HujWP65s+y0gqFE2uzjf
ORJFwLK19HFlQ4vOCcwGfUeqQkjR+ZEQI4gOUHCpnjy2eUVDRsVectWxxMYvumankEgEJME5smex
C1nWJLzMYrDABDUA1qa4mNPaXZB6YbXNdUGQZ2kZNUzTxWj3ZGni6tmLjiLxWXpwHc0f2r5hYZj9
Sgq0dOzul5any4u1Jd6xJwhyXq5LBjAepsJNYQ4Gkc/3yt6W0mZEo1NA29ldyU1IH5I2F4F4dGrd
WuszAP6OMM1zi/VBMNER7icbZolux2G85Hdyog/I/9P6tzrJhPk9S58L0PIEDEmKfO0jy9OT8bn/
sjZpzTaFuuUmR80hcAm4rGm344ya4ci77KDSO2solnHQ9TiUFBZqHYav16VG8NZ3kR83oLzqqLcm
qzqElKlUEpKdLgt9QT5GAlPAr/mWK/t+R6KocjhvOeMMp6ZJry2qjNdSIKisYghO9LM7HlxlJYrA
sIneSEQQ+mlktRoorcED8yaBxSJYdw4STTEfxcNhUpm6SomTbD0GI6cWLx32W9gSWF3VdQOM9o0K
sqeYEp9aliRFRKjUT/6t25qbA3nC29gDnELMlH/K6dGqZ1hrsZyW476vMo8VtbE4a9W/DR2lxub/
3DH3T7aoIzRaroRZtCBz+X6ai/8HMS1EQlL+sTEb67kBTcg6wMJk5ae36swECES+KGbl4uOjQNqQ
gzKPiHRzr6ZMyHEfp/2uCwVH7cPx2a4UBKmoBqEabtEcbHDxCIzgU4joFmgGVpCAEtBtuHtS2IwG
hBVfY2EEA9rS2tH7g7AZ6Heu5JlyN1dpJSzrLbPa40j52P5RWj66waZhsRIdDZIk5cL7yABNB1Xb
SQAf8PxNoAJs6gbHtHN7Qhd5IhWE7v3LUwzuJobHktK1ii7z2MiEjWFImR/h52Sz38urEIffWxxd
x4P2Xw54+IYYksMjAna0wguqy2HFu1P2bz/Ys5tD/TuKsHjsYN9JSvdpwzWhZ4JooKLqKDHSeCHv
oFFuMQYO0mrkXSZR55p3CoTQlslMKI6MmScnwnglGbXjSNQkgULb1YQQ9ofiQjJpGy62c5MmDDJD
BNpUGdUkO1lvtoVaDShJoXBOu5gQezYTWtUF73cmVO4zgex7RzOO51Nl8MSEz+bqF87+S3e9iVkd
9MOGk97mFI5K9UveKBbBHZQj9a3WRLsZiOgm78di4Bz/yPB0qH2xrL5lJm7lNw2xNn+kpLdUWgxi
QSaS6LTQRAtn97kciyYTbBY4cxZqYwc6zCYaCFMVJkatGAa7b4s2ulBIra9QroU3CU9smcjRBpgn
j2G897jKT4gvc8xy/dN4/YuMC02fsPuFAzPjfxXIqpuRFvVfwf91YbmjffNAZb1gCS11jomFTLuZ
/mvILY1mt+SW5yPebM/+oQduwUyf2tpG/jYmg0hK2i9M4o1vEdkQFwue12aGR77fkEeUTRsd5IEp
XStBNP61CUA+/fmuyOWUrrbCrEo6w0qfsSlnqKEnL8O/S/inD8KI42LWhCLLD6TCSQV5rSr/keT2
PPWS+YRmvlZE6pwPN8u33ExW9/6dqRGntiiraMkpLEXDoOuhpurq7A4N5f5y/KucrpLkp62wCSNJ
ZUWbRiXeRjRZph+WLcpEL2qPLXAulU73GF5tFKEHg6N3UHO0j8VBx3VuEAJ0bpfYZ3TGmyqLXZv5
Eer+19mjRwBYfIeyICWCdp14tHoUjDLQ1O351UTHDFvbtofBR7yIbrPcyOwkGE6uIeM+yx63UUxV
7/F0I5kvWe9jTEIZR84t3fA08RtwKgxRzOTqVSy/cWsjtzs5Ld/0923z6sdGUpIkMtyETNKtnV52
hP21OmWF09DKNx/v4S22EUjnZbYbzSEcqINivdUqm9ezerWV5TfdVP/BoxpQ5wZtSo9dRwJreZmU
C1rJfDxRCJEBTsw+Yl4xLdORcakQamfUf8PIKhzQLNdHcTMQKN7tYZf5BJVfGn4YsAGfylFkkgCD
EFljlgFYNbxQRnW7Y55NSXIo+JKjnTc2pkFo9HXmo6wMjv3+QPfj4gwqNDXkbVLXASbjEWmmIcQh
94LIVIlk3fGOpqjePOoY9IHAyNcTXk41H/9vlKl5g47C6kvdj6IK0fGEp7H0iPyV+QvJ+ZsEFTtU
0uxGvwJCXOwILdvLe12i2v91qDFHYoOE2xW081HakYqvxsLbbZpOYB15bLZqgCX386Lxdwh7d+vW
IWdp26MU2/oNNgp4QT2tyDNC0XgKs7VK34HF5PnWrDBer1nOW97nXG6A9vBk1Kchx89Z72iOl+xU
hYLSYR4bVJuIdewGiANO9UYNU3eRqd4oj3nd9KlUUaG9Jt4+2OKYmowo8QnqTK+c5AwmN92iKS4q
zV+1jBvl85AhI3IReCAFsc599gUUCpj/BZsxgLISxiqAjPicwU2gDPb6GSBmMjVbKnI53mwZy/Yt
3bb6rBTVduO7tPkP9a6vW3o+q57g+0Qgc4hJ293f4VFF+Jo5F0I5638oEIzq8pDko6uu5jhy6EXt
arz2w9XCh9CD6n8GmtbIX4wV2e/1te27auXFF4ath73ylWmVQXRYvjnmOuPga/JlERk4NdGix0x9
hlADAQOGliHz6GR9Gst4GcEuFdcCJAeCQGQNYqDh323FRuVL1vVZWpmSOGa1mUR2FCr5GjB/ZiQO
xI4xviQ+svTGAxEEmZ/1QCz5Q4Nz8FilMgWUUzhfhI9K9h33yKeRi8ndEv8wGM1jSX8hZABCvR2x
Pr2w+zKWalftNPUXv7PoBYaBLCSfJmDIn3UG73j0wzDgxmLMsrT7PB4RKpPUl6iRHtTK+imeXcaE
0EUyis5JDDA64dx1ijBwZ/Sbd19TQeYv/MlcRP8fQiEJh/l8SninIKM8fR1XMJGd697WmbBX2quZ
mhuos4NSEaA4L1dKUthTFJpo1263OQd6kpy8MvIjEQLsp1Ywa0BEvawKbBiXZl+bmrcHJCi0QI0y
mctgQZ/BXKbR5PxP1+Tp+GNuIyPMHNTz3drLacyAMAkrSQ0bxDIpsa/8AT9sjWVhUUqCkxkF+Mza
mFhz5kTxkVgsovoqAcb0mlBx/yIff2Bq6FYMatyKs+Ye/P4C/4jXvA9HqsIkk65C97esaxoXJD8P
2tNUuiF3s2k/z7erzvYXtikXnOCqZM/UKQ8rW+q6LCq49O/zF0qhsIfgAvTeTYhBRwvouV4R8GK7
/UBjVrS6qDT61iMEHMB+yQYZ4Qp+SwmfeDOthVtbrchkpfDVfPldrhOEgly78rzzHi700h6hhLs/
ofrc+9mDnSTZV5hxGK3dDmzuYKDxWSs4yMLlsq5+k6mwFzzC3shMKoH5OX6yefxHqVj7N6cRtCGP
yksiOkwlZ6C40wgyVG77TZa+Mqwn5RMjFDLTilRJqJb57V37zp6/NAi6TcDzaIpNPdaC5wrpfJHQ
hoYHVQ9qWvD2hr4eLGUbq20BsgS9n4K8MKA3wY7ILxYgK+fPq07Ok+qRjh3SijlUA4Wjaowos58/
ViU4vkbRl2uNvNi2vkf2A9os/N2vgWeOCpxUqhKqGbwUiGRoRJzymZaA24ZGKsg8NreEotrd07MX
WCiiN3ZFkggFhxtrhDCMozU38ntNMGlwlUZyHW7n4tCfq2MlxAxH+slU44UGYYZnukCXTF75L+Ha
8DjgK8cTk8J7X5w7Aaval4X8NuAcOdMTKF5qPKYUVr5NOSCvuTgI8CtGYtIopKwEt6Ssc7zb15SA
JdcCya2jr7TInSVyluzgJPePCasVUIDwp43ZAp6P6Zgq0mW6xMEY7U5eiL16/8KdI32J/ViOlqcI
KH7Q8sFD/bS1jdLEYCSMQs8HoAm6TuVWUUILrbzPti/5a0h+0RCfOpYAVtvQQLPzjoz4T1Rqy30S
lodpUvEk2Bj7aDdiEVTHKVWZGJXHCGOkyraB163zEan3RmTyzMs6BCvZ8NeV9t60DwnVY8KGENWT
xEZPj+lfCqbLtCV6wsqNg6oD3xNcJczE0mZRXybAbKC8Wr/1aXJx5evp5CtDhtxeNBT24R4xGrxQ
IgdyX6yVp4ZJLAbERz1L+hHUIIcPmxE0uJIXZxBLTiv8tC1QXNawvwdQiaJ5ZLa9Lt2SbBUkF1K2
zJxa+EDnG0CTImrN/oiEVRVvrrrq8Lf0X09Gen0ul9Pr+gBwjDr6qGvR9EL0JwXIxlTDVWrvymL0
90+ep+clBgLclLiqOVflHgDm6eaM5VuYAJus8x99OGu2GuBlh/JNxoEAhscZDL8pqygVzPDT/+v7
sWyjPGVW0jl/MbQRVb7WhF48zM0954IbhCuTkhpvhhcnbC+qOgDkYF0t+amfgYtgh3sEzUIw4gUf
4iE9wyI6ESXwBShLurEJcQ4Y/lKPcVYwwpd0LtMNhq/BjXO2RNy+J6tYV6IQlwnlEoy45YcrJSpQ
eITtEsp58Mrp3muZumMLDvPOMuaJJpN8vDTJSo9gauki2DMhedonjS9gnJbbGSmEGNKuDU00kiML
UWdyGQP97H1b7/5OWRqIIzaRrSVIVUZi+0a+8YzfcTKDPrdLtdr0PbPoa9HIBTe236gq85hnIpSb
ob26iTL+5oZjDM6Ffbna0ADof/tOtYsQcb0FgQZO1d13yHZJ5AD0hzBk9s2hFMa51H4SwoM7x2S+
sIYkhVhqh+awM/+tuh7FSx/2q1sYbxGIDxpZwBhbt1PUEJwVKP/LPjn88fPKWiKKJA1cDzX41Guw
cxwf4SgQRUFluER5muytD3jVNlWscPdh2986kw6FCo6fbM1yEZ5Kl7Hf2ezk4jCcXRS7e0C1j0l3
kquuu673IJgH+QVlrP2RuS2sYK/OTtXfvqezKI8Ve9GoZtS5vFj99u3HNoizWso+90TnS4AZylra
GaFI+s1bEILuohNPE5+D3pY1snZyITiywKmlOunC3m1f6HHgy6Yt65hcHFfbIEk6RnnZnQcaHz7C
aHU4eDzGh27cqGMXTtY1BE9lBbDjSC2t0Vc1oaYbp6SRe81O+/tLNCEeltQB/R7G8ixbNtljChAL
JglNXT7q8t4+3uWJjp47s75sXUy2Hu1o7b849AGGabGc8bzAvlJ+4VsD0ORJyxct+1p8odyXFu2g
DU9Cz5SEKScdhPJ1hlsdcYeGjdFao56RYCT7TdWREP9hs9PF/nc9ZHwNraOQUZfyNoiZEJsuEAk/
fsY6nx7oK6QbmdEjX20OaoRTlyUkebOVtfnPWfXtvEUrNWPeVZkvYkjVmgWuWOwjnWht+BUYiCE5
6DaIlCMSqkbDM7i1xd+RJ8T1Df25RLL6FPuXGVD/+LpCZ8NgGjZx5o0z+jkV5VkXwvdbM0OmnYmf
QyKg9TLhEbk8N7rm0PS1afq7Ay3JuSn406hAZfS8lRQnp6KXB8Qpq3oO3u2g8rMF3Q0yB+p0TMpT
ZifW4gucUnG2oU8YqfR8f5dXNDR1JQw1xnvYv19jWVEW6UrmzktUWiEy/AWRbKep16DVb8gB3jKN
9Z0ob7kRgoPF8DTAzS1tSqwuSxow5IO4tw6msB2ZSIwsEtJRhQ89+C3lcKIrY4DAi/u5aglNoVKl
FLeMFtzD9ZemzQB6QpPhmR727E6vFfeMduY/EeVFFmB6+usNf9wNCfgCVmAu9RG5ZTNyIi1W7Rew
+mCxIvhQVk4cUers5uVQ3sp5ehX6EJzmi5vf7g8cKhnhFsDd6le+0P0T1RKUWrzEwBWlulrnCUbJ
wk3S/udHQsxNdbhmZ7UAoq7GkwAgXoPnXrUk+C5Xy4a0YU89cHIdXpwl8ZSAzMs0aST3uOH0JAfg
9kt1Rxa8rvl9NodLKk7+aCukTmQ54YuWVWK7LiYHH96CL6VRiOo6EUfGIN8++WhB7VIqJ1ehULst
OhQn6xek4Shx+Uz75GGP6RTGjhQHCHxe9c2egsmBGphlR90W2v7lFjG8KgVoccEUqFTkbkT6Jls1
BE/3LoRFuJMFlf5sGROrdIDiE9btyMiKQzoRFrLUIsqkYU46RDOQtWcaIV+Ws4GSdWRe9qI0V3wu
QAG60F+mxW6mFIQD7dgRjUfqt7hZhCSPUCLR/hZvvHg9cp4GCzfDDR+tyPFXRszyswMYhaWrOKqh
oDD9tVvU10tksuqb4GIMlLggItG/exp6xpZo4OUjTwnw7qHyWxecNgX8EkMXI05xLKPnQNkoQ+M1
aPLb7j+X8KTbAOzZoYmSLdNpRqbzeQnd8ZtzlObfyM78pL7a/8UzEYLnuSfVhZD1TeNs+xy49qsa
cZ0AJ401lPpzZY8R8jHgzV9TJRkjBBNzlswdfct0j7HzDp6mTAioyu07dmafaDLNktYIREfhZ3su
AQSefKjFpZ42fnJV46+UFf4CtxfOvQ/BF2Mw9MzoQOHjzq5HyrQ8CArhIAultzKvkbXQl7d1skMd
adde3b8iPV2uM8hPva13jHioLuHA9merY5NYUE4Fzb+oLrrjORubI3dioyRXfDPT7Zt4eytTTw+H
yfTof/obLcq4+h+2MXCLrZhQ90nHIOFVresBGv3ET3NYjbOJ/xw3BVY3yPPNliQJxjY2ginDDEFn
ntTnTfj6E69+FKMKn76DJtbW9W7odsSSJV/U+F+8T2Y5Eju/uOh8OGWZweBRdd2vPJDxoT9385pp
07XyMUgVgEGAsDH6r1IZhtgWPC4Be283J5+sOSwWQZForkqJ046kjCFEJihA16Yn0OUDRPPy1l0U
t/P3xJTjRmBGDYDiipFtphNe+hatsAY6V6kzogFcxSLN1MxX/YCTSZ5Rp05j5Mfx7hWXxFfj+imL
tSBwxpHutKMbwiajKmGrRlqmip/WzZlGyGgLwDtHONXExgSg2ngPwkMRKaYXZFkVzIkIaEOlYdiP
D2OBKr1nw9qyEDlLuAn7CAdJ1Kezx8w97O8uEuQs04a1jlF+NEbut8l5tT7toj9w1TulaDq4Hk8N
OE7oVyhq+UNLsss9lU25v+ryQ0KkHhqjASMerX2mHTIXIrOxwgdWwk9j8rngnxh5rQddHl4MxHfO
lZ11xozQHpX7L1nD89umETy3o7+gTixYA8Sp/P5nKeZHBY4Gyg7sW0X4ajWW/FuP3erhPCQoZUzR
sw+y9vv0GcrMTlhu7pw7dR+oCogaiLxZhz+NcTNoh6JlwgakuSr4NoCta/9754hAKn/c6YYZ6T90
0QLGL8DOKZDrfURJgb4u0HPv8/drkbrdBIVDlIQL4pYazbEFpeabmIglRWK8kjU3nvdCA1nAuSwT
m1kyzIEQVFppRgrJVd1VH3S34DuKN1UVE+pGwn+CAxoKemA2cxSY/DQOSRr7j3gc2XxkSR53NfjX
NpO/J5yG0sC8CmgP81K9UtRgKSmYTWibAjLaj42sxjvSYXq0zs44X2DpwS5j7bFTTA3ShKklxPX9
ivenMmm6eZ5SfiAZ9BYMl1Gp6LTxxvumG5f8B+TnoEr6BZ5BcK/fTHhwe+MqaIXtN/5C49ai7YWT
IxxVcwtCewbzDWIKfHMRdMKL7iGe3dCmgP/n3Rb3dI75qJJkpeF7EAPlbGqM75JLRT8TeJiAY6Fp
ovcIVaVvvrNhYbAV+vdlS5y1eOOQ5G8ksgcz4llPDRWWc3v5bsndcv0ZNoD9xe5uYhA/+ZIYg+Jr
mqxzDkPeotkOjJwWyGZfoYdqbGu/d8dShab8Y5Ov8apc5n8hSLkXvPl88NKTrTv01k2qJnpTuy66
55p1cW40VwzBz3pK8QsXStdiDlne32w1wVXNKUi0fke9Z/KcClS8UGWOEa4ZRPk9pig1Vi4R+GOx
y2Kpe6UAAYshnsg9BJJ04Y7XM+oOlqUyoX3YzOUrd51MN5s+a9+69kq2NAn5J2Knb00lVjXW/3C1
7hVlQWE9i4/4nf40VjxOrfSZgaPAgBwAXEAdhlZUcHESQ5UdR9yxPq1RzQpx83pox23G1fx1Pcaz
Moaw/fi5MwuhXMuV5x+t8duWyK6yo0mAg+MSxVcvPXOwE+SjqFpJr2L55H8iRrJoMbGJih3tZkif
1TZeperR11GTLQz+nkFkwIelL2Agd263gh55xXI97A1ixYMroTrWC4mRXS9v+vigrCb5dPt2i/+f
jCBYHjXQNw9aD4OUldwFtJteMNUA/bVBV7jVrjD5ijBXCYjs3WV4oIgspmT/IEZyVPp/tF0Q8JXg
FlEHptOz6rNzpLcB5hPY59u2M/KHooNs+vDrloejObOpUo3RWuZ4Cz+RlzwP6xtwVUQNxjPUsmqT
AmkWQ5lZXEni4bPW1kN2SYg2DFBNbfS3RGDwCBsbpLUiezAf5kN16pS0RD+2MNptV4azBd3BsLTO
/YaPQ3ExOKH6EoLY1Vngx9JoO2XHPZFvzYGFeMnhcb/+ThABwyk+P7ru0ozUqPSK9fYhWv6myZiZ
l+JRibNvudmBSEKUbFr07LLP6E274Vv47f+1Px/E1X9nzL5MFIInsWVkCyOFL7ERd+/iSMazcwNy
NJeHq88dIVCre9wEMcetjnwABXGE34xL3qTg7YBF6O73485PNf9QYLxkjOiS1IEEv0v++cZ9Pq2n
WWueIBAVX/KrNH8mk3SxFbJrSyHU5tNaX3TenRvNnExm6ovcTrOw9ULucSsWqGofSjaDvblYmxVP
uVdu63Zql58U8MuGdvYkVnP+3Rqevm3cbpPETdkTaGJPLlREKYeZvFPYysF5+RZUOaBiGOnA06sT
zXT97ZRR4CxJuOJbRn2ymMi4nc377MajcZ0bx0QpVOwlu9EzkzOGDby9LytcDKvclMT1y874XPd5
haJ4e2q51NLnS/VkJtkAi1W0a4km53j42Ed/yjZKUXTYenil1FPnfF9JjrGTsHPofL21WpG68bNs
PXBtYGhnh+cmAE524CRIf+Poet4gvrgj7m5Nx5pEeeVoJkhbGnIRs6TzOGBgbTsJG1u2lYNEQ4pC
RgcYc+RhGc50xWdZXW/mzw6Oz1Wm+ZLl6QPMWIuemh2+wwDSImo9fD5qpqWIs+iy2/mVyIUKp0Mp
TxFD9aItO4RNaQ4SeGIaqyuae+Y0kj8a5/TeAiiBYOwh85vXhqzsb+GlysKK7heQzFqnndewOJYj
vQo0J7fZLQcjEcuqqD7ZMIBu+78PPVgPIt6yOPd0DT5VlyRdGu0ofIh/cAR3za3m2RXhWJiY7Bzg
cogIDl0P7j0wyvIZB5SOyJI9hCcQsqMWvWJjSN+RW7HP7wo37OpTvPIxmjNvQhbq/8zCnvqir+99
D1D64RZtzV1MgTbsyA80wYbm43LlNlLdaJG/wqog2DdvZoflzYk/wUrzVAQE7A6dAOdZkoCqUK7t
BPml9+SDGCCZiF9z/MKJZ3VW+SpxtSkdPE4EPhIoyTRj7OXUKYYXBKix5GsHBoSHsCWMuDNukrSK
AORJGZEs6mq7uvk6nyu8JGbwPqY6c2smLCN8gKXCCjqCQTM5nnpIQTFr7C5MSXpQ+39L2VcbmHfo
D17wRVmJCqhFO+6J0h0l5oC5DmPJby4gFz98g87RJa+pskQ8A/MOLlVh9QBauEwbCeMvr0wcTR5K
Mpr//v+59OWai2u75ktOZeUr/S+qmDEGvWk/F9sXex7fEIjZFJiJ5XHxhDHlcjZCjktxt6+gji1B
bePLnI722WV3Ec6ucZd32JX3x8iFDL9ALFL+GLVv/cN8v1ueyAq1Z7urw7OzfT3il4QHDE1jJ9rM
qXzS8qe8uz+AqKQcKBaUqnSfj15v/JIbHfbXD/FH2i/8fgnc2URch/cijKFOqGvE/ROU+pSmENKs
DTbUOk/pzSjXoTwcDJNjPlT6blaV/QMNH1FkpSViefaF4DwA41+CUWGodBrVgOq7znZjyYcWJZDD
PdlEdoH1ZNNhtog6QzyfZ1DmqUe2DE2o06zzPjakZtspQABipXzTDoy49h28aS6HXOHb1Q62Ootg
PlzAF2cc7LwfASOo7B8vzynyQDqu8fCyYLLsehCjdfVzbUMXtCH3rawHh8D+b6fmg690g6izQ6Hq
KmBT5KfTqtjvnqNZKsMrd2DhSboaT2pHjVw4UUtUNsqGExCjk6KwL1lYZC+DaWuMSjOUcU1NPtCO
dZDd5Qc0Iv3bghSWqJhgNTETDT07YKzJRGga5Bvun48GGtUa1sD6nqxa4P6qrLSoDgA08obZT+fv
QGy8DKLTdUcsjenpnATeZfffIwLi7BAjnGs7IFFixlbg+juiI7XIqgQhZyeuPVb4RA7aZtM0rWjx
1x5GsyQ0VNZ+KQNQEI9El8dxnPdyoR6cFxirMeL+jc8qyA+Ij9StEin7rdR9jQmJffPP6QlPr0Qi
NHBp0dX0/4y9cMXJs31EvQZPHxTbSMY/Yo533dBnb3nglxAF1poX0zh/VohPGtmBfTOptkbWVrB+
PF38iDiUOwpzgwz4LGNv6i/zvwwljyKB15ZrbKfx+zY/dAeCRSMfPGj+ORWKpkZP6+DOQo2IHVbz
5BzxMr+F8sqJrORtlzsfLVKPJkicKPF/E9wuZT5z/P+EfREsx5qSDcDYKgTE0I4O4hGjAntD13CL
wEZ0zhePeSl4vN0GKxPJrwoAROzZshoWNK7g3I28io1sK53/QSzfTmrDn4l808mTYMHDknoHWxwl
RmnWUbipi3Dwo0K4wL/8gj7q+mU6kNg2xz2l8ljFYDe5yOIiht4823y7Tf/hOaZqLZQpxdinL194
V8WeZ0UwS4PSTx+h30R6EOXOts4ogdWTq1GSCLXf1fSlInN2bzmHc2JIu9ZV/8Bbk7XyXajT+LZN
ci1Kn5mCXi642BOKsNH9DDy1Lbet+sdNdaOAHPCjvrwIho8plTvgxCALtS8qqKyOetEH5uAYjyhn
QQhEqNcRnZ2lyF0+wlzQnn4MSfTSThF30loYNQgDnbtgm2iD3NkgTsjook5FRi1+912vX5lxWcUt
vtY0CUxejyencij+XOGsdX/c7PoKW+13IsphPf9ugoa26MN0x+fA4Kp0yfcamOvSM3BIo2vSE9yB
uuNwhbhxHr4cSYEpE4kWoJLuEIZGp5FFmhOc+Sj+L2PjcibSn0kIvCMCIEZvjmgJMs3AwkKO3DwR
SNpnjJEAmXkeXAAAN2JqWsdY30JxuneZ5MwrWYpjx+bumTEXFeBWoeInP4RQOWn6ltRxQb7UycU+
yjCs4oGm3nY8WWxbs+UU3CKE3OniIzAZQHc2RGFy6exuyKmqY0tAYN9hxrSp+Qi2klVPEXSJlEfe
aTugsUnLMMHadD8ukg6Hts1tsKaNsm9AmLfU/eNtMaocS0+TebUlz4JGBmIqIEapll0Vb/yzj6CK
lLHFXyZo7FbcpQNghRLyruo3p7BAeaMBg6dY/5OMWSCbNv/RnjCJbzjVqJhdyF2j4BGV0xkBZNSx
h6kz7qOKM/4/Ld7k5xTXT9YMO8RbqpVE3ZbnAyMTB4boSJuQSkU3taLgI05kSx7pQyYWXl8D8QxU
aiqHSS36ayEYD0uBP57PLHc+pDDV1NTnNyUGoMatG5YUf1pliPAipj4mzAiPt9VmbFPQrOo4pjzW
9AFZlt0drC4/eyT4YeFt0Ix/IKXeT5LWuE9a2tSBErttsW2FZ2aqEbk1rlNS9GuBSEX74FbDCrJe
IviCrb8T2BpHV7J44kVF/809GjK8iXMiIr5z5L4ZdXeW6acjSH/qeIoJVcGr1ucud6g9nNqaeYPc
+Az1piqHxJDo4Irbuu7EJowevq4Re4CC1tc1jj2P0QfD+Qr3VeyfY3h3d5TVIArlW5sorh1ce2wO
Di1YxdEbO/h88gzUxOsflwqU4GVEiPumThLFc7pMPzqh4AuwEqsIUl/wgBPNg+85KurdC0RUD5Xb
orqqW2Gk8GMxtQqpG8ZeAcRE/F1xnxkcHE/SgZYEG/UsxILET2sBtNbWsIagIoECaRbUoyYIr0MI
e8qnerOzt5yhV/4hwft1bfY3haw5DFdgNKiTfEUIEWAaBbruPmoDEtiIWHVVktkjaTNjieorShnq
QQ4b4Rk+lXcLU7wuzjVxj4hFJFww1mS1YaNUeSbSVF0diLyFfFJn6MhDZXx6L7FwUcFjSHYzbdpe
TrfbCpUiWEL2fTvlklYm8klg8rPNfy+KmjM7tB0wK/gb35Qw+oHmq5Bcn3kCxNj5OXlXuxgns85P
djms95KQecv5bgZVPD0OVpIzpNPZFlEv25K/IPAp4+gsfNgyNCRGiq7PtMVrysoeqViksim2eEev
LbqGKBemw1QaV1Tye0cmYo8M9/SupAfK4qY1V0PMuMoZOkXgUpGqUeof85P/bv2tEATiKnciqH4Z
WBFPZ0dJ5z5msIQbg8VGgf20cVDVHMYUuJYQozK3Smstt7+HQPHThPZyiywyFUzFCEDB27XLJpsp
aebsrtiWfhNzu1UwssNs1MLJvo6DrB50g/RdscAPloLPVL31S2TVsXDUHDhX/K3e6VSzlfPl6gK7
TFKERDPgRFQ9tUF895LywJmoY6rZt+YzBg5r6CHP6aJfR08O5JKsjAOdsSjBQwpPCyQpPo9UlCtk
dDXYAPHvp6aks2nK2UwVAhTOmEZ8pN+b3U/jCldEepQ3kR/ZQ9EC5VyTlSTjIDHlaE1+KQ9HhoDn
qWlnUpx+R7FNRPVHaziqbZCNK/RhnzUEx1iFEKZnLpDP8Tu9UtnaTDcNbnFZHIpOeupMamWn5B68
yxei81AyLx+rPvA1PKU7v6+6UcT3Xby50mrqd/TC9YRn9IPUO2MBW8IHlQibC71bUaAaVmhZyheE
cjDNNIYTMa99UiwN+2Gu7xbG3Q17CKGEoyjQrfbq/ti1vHsFg70DR/ySf5Lwg8royVOMBq+GfTVm
7oUwGo57d6bVsiFz1ywIs7qZywI6Kg8p9bY+zvMO9id7yaTCsv0iAY1XZ0v8LNOrtl2YwctUsdt+
QvZkdFTDNQn4OCjJ7qHECjnfZm6c2pQAxgiw5xgH4b7kkqd24NsH/6K+GPzcwitfTgL/8IgQqxpr
cIxDmtzqYedAQZTJkmV/tlqEWchaXPuRrNowgclzPhGDKDe476yioo7hldaV9ABxVWutfIzeRINh
XHoEUNhcas6saI/ahEZvj9aou6hBd4jZfYwyzAzaKGVtcbb6/YDiOTNfcLAxhTYoZPGl70FFyAtU
3F30wPYWOinLs8Gam5TuhNZErg7rwjyNcCNdmjwQrBvkX9TxzGlmEn71zk5XrXcsSSPPP9Ruj1aT
SzxEMlO0T8AKnDr3YW+QO1ieisoEpg9P4WPQDzYsKCdDiKXsKLFFgBMoo/dbA9QSealgxcnKgv2x
8BMtohdel7qT/lHT2m6ZuD4YdYm0yjpW8uAL3DCIYTBN4Du0EG3aW1L1w4JUexsqWpq/Ipl2RYUM
1V+/So0ZjV2Pi/mE19gaFrFBt+KY6smRsVgmJFW3meHXrWya3WGRiVkW41c7Ur6/JbIdIOKUrNK4
FHWpJdnUPfXv2WOIi8bVlonbSj3oBYW2ho15cT8lm4bJFpT6JYWxwIhqARZBxCP4F24x+fYc93Ns
/6keqNvNFF6/stDO18+ldUealHa8SgNejlO3WcRyBCDnXT9yo0OPikV3Khw8GbuHpgPIq8cEhHor
0sg+FTmCz4AmTrVzMae6OTJWe2ScfNWSGouE1VVwSiTl1NioCvz4DxSql0N/FnrHZvm8RubaSgLP
EHh35Ns/N5/dh9//RFsXMfmwZDtP3jV3+0JjbUIs5heW7uaSZp5etOAFfYX1EDFC5A5/h3Fpj5SR
EBN4ucEIlSBWZVb+IyEGRhKpqqPfGLbq8+29OEiTWflOM2qhBu0hU8GrGpg1nC5dS7QgKiopJBKE
Ir4bvCn9MMfA8Qv+2mbNoXUZtpo4kKHpN2WAL04jOdWDzyTp3qkp3hKp3m5FJlsCXIYkCbvXl0NI
hhHBn3GJJ/Rx1gnTu78bvW9kkshms+lvwu+ByLAnzEZdTzEbkQpDVgk8ZYUwxisF+qARom5GqQpT
Cbxh3piCBVKwLul+qgXwcQ4XYDTYdGFh+dkBRPFKhB8fEZFRVglLSb5IswndbwXGRE+h7FGmDC+I
dX6ytRiPRxCWxM85IL6I94z2i2Ij96x7tGRz17hjGoe+d2pO4/Nx+3df99ap939xYMEuiq6rf/m1
kv9Tz8pTuiTDVZfuMslbQP5mjjAV85mQ55B3AlA+rd1VxYCYou7okjzW8tAuETp3cOJWjXbXRd9Z
PznN/IihJKPmtRqu4+uFmtqBpYtlbpGaUY7zt8PXbRqsPwSsEB+L4iEMMIEh0T3nxWqvmoUeLk/X
ohNTeicOq2JiFmMVxbBSbNOLGkAJEkStNPK7NL/fsxbQMng4ABwMROT9QMXq55S+cwh19fpZr0tY
2wSHvNJm5rt31pOspLUE5MIQZHi/ZgW2ZxfJRGnCFHt+ZHEBx2pIVH0Rk5FDsW747oz2zRFzdV64
Wp7kVPVO52z8Nbi1HeMRvXTWPX+M4EUlTy3kCzHSSkSYdFoVE/HO7brbKQsF6qj/M3tyub6b03d6
z1KP5QYLlNShGYdCjD0gOzts7Si9blG6Ziq7XyQLKn7mrK9UxzKo5DOROnteLyp2TBN1xnT+FF70
UqJCP0+qJrQzFZpZU70GgzaRRJna3jX62E6T7Er17oTiz55aNEk1wJ6BMz8PT0oayM8OM1HLeukl
WIUCV+5PbWwo3W9XXbIU8IF3jv63B3idIJ9dRD+BaRqOvp6AyY+ob6gYg7/YnF1C/jM3Q9u3X5mE
WCe04MTYoobpVBfFOjCBTi3EVHQk9s+QT+gVnWjo1S6JRm9pxxDK7zC1215vVjt/Pa5T/7iQ+zkO
epzUoOGGbj7lQ2aleA7ncr7KoQj8XpHldAeOBOkRsG6t3ZqmhkJ/8GByWDeFXkO1glBWRAxn1u3j
ziL8Hz50U27++YmVUyjiiBs+fuHkdzt145Sr3NQZKZdi5eGP0Kcdc+s8oORtfaLLj9DTiFAhs46x
BV+iuA+UDOa64Qd8ml/+eitXlkMDWb2snviipFw+kcB5bMRXMOHH9wpL19mrVVla9wjm0HL0NId8
Q96OKu3qXHAL1aZhdw170JWhBb2gew5dlcGHVmX7jvcyXYfEokS80lQ9B4uG2pXq8m2JQMkJuwzo
CzDdOh6UJFH0KrrpISNbOxG8X78hpn2x6C38CBmFjs34L2kIo3eNRYIAQponlzpSpbR9LFgul3R+
PVs/pL2ttemV/VnH1ELWTDVD/AoF66vsyrnsRh42+VMLKjKSOn7zPNHevb+cd3s/hx3fTe0M5s0D
/KgFrta+UTnUogp/BwgcenLBVQicoANUVE1T0GFkGSUQBOOMUwxw4XWmFxOXzhw0W4VejTq1wXqX
5VFDt45lFv2joWHRvubB4CN8/DuKiz8HzytRbOfvl2m4TH7+RbWJthlLYazIT85+JMz/y21WmWjg
apIiTC1V8YFLxKnZ7ulqNhInmH75KcRzBlM81BApTvn8D5R2Hd9olXYEDDVrwXF6OuR6HC9xbaNw
zwWtQoe542jVDwXjKhZ7ihjwfeOK61FNGCKrg30B+1jiPEnPCIKFnMjQ29MZ5+Qiq17l5j9yrSRG
I1E9AasnQg8+dQ/f3BAdeDuLoUTCalFrBITQ75jyG110BhCMdazfBNV8b5gylaHYFIaBYgdFcCB2
Q5vpZUyXoRQZsj+yE4GDk8VScmhdyoi5LP6Tx/dRH80uQHgRaJfoKHnQqwpv1m//DAdbhIM9oplM
vHJKPoFFxzzc2mxm/0J6N1MjhVmQp9HJnV50ieRssRza7Whfj4zc0x9ZM07K9AB76oG2Rp/j9i8f
kQpIg1O9EiEZHPxmKlGcC5bHKsOGsT6bLWar5aoSXaLNqGCaODUAYkW2WmNthpux9XRZ39YGgzao
LW06hDrn2zKT6Xcw0gRc4iNKPPo8xNg7Z/2XNc6hQtJcUhI30h2xvKmo8RLDMjxwfoQhXQfYAwfQ
DbgQ6rd3UBObNhh/f58UUBbp8++SmJ6C99jnvZtJdKgF4Ro7WIm7OQb3NE6cva8j8CA38wNu7uvj
r+Bd8XP0UQpz+xRiKhxvYvbSpUv0sL5fNyH12O7WL7QwTob3yOhVYxQ1QozgpE98CxpDO2gdZpg+
TqfF6Dthxv91hugctqUZRqSiBjm3WqZ7976RsF5W+u8I7EY+Bq6+VE/jRU9Ery7WCAANiC4NOqMS
qw6YnlvLI7bCHbudIR52GQl5/DgatksImZ8g/F7/86Dy8sPZq9Vcjv0gwIFYLToQO0w9I3BnMoyZ
8fBm8qUcyA07mtaO8H2M6kXDtjbzZyV9s+5oe1aeCu4K6FK1DbEfEIgcxIdvgqVVtyvM2rEzVKjd
Rh0M/uKezZAeXkj1KQP5mV5YdzxW5kFgSMYlOuXbvyfONSzD76UDL/ze8DDDNhEfPzkDBcsEN8BE
ruu/gL7Y3T7dNtCd8qRA30wmjVNizOgAHM6xG+JrcuLB/jAX9Yzc5z90ydMr4Cj0NzxaZCIHUQlu
Dp51NEihV+ZkRLldAPMybY1feHeZhPcA1LMKElx19MQF8qhVdoJ5I3WC1k/bXuPUU9dz84OuyLmP
jf59ZuA/z1fffwGv2R6j/Cq4z/ORSMnoC3wUxA38tLQUD7ut7dq6ch90uXKgJabJm9QouYYJK7mq
JkTAyZEcl66rukkIIPuXUvV6xTmQqzeItev2XFnvP15RP38OvcUniGhwKgBxS+7zVvfIR9b/Pcae
qVAScOyCXu9OaZD4mUNGv3Fe8PWSctQTevBuVEQDj26+Ol+rchZISty1/rkxbU2xkEYSwaiXyxS6
6LuGhrx3JLTTrksqCDPDhX3LAaOTKGoI4wFRk7rgr+pb8LbleG/ue0EjCTf4wLZn40eCNp2hJWWy
cETaRC0htUxUTnUHx8xg5I60yepqGQguOmFgXGbtrJAiPXgnlrGclVny/aa4YxAynEMTG81NhYuK
v/+1ZYovKd2O4dM9ljQYkOqU2bJwN+IgAtUc57UcUrCsPc8S5ZRfpMiuRE0sHrt3O2QtTJBzQTPB
PoVMT7IoWnCTeOdDQSiP8UdO6HNoC4QBWZTNq+XLC9Qf9pIQAFIah9wWpqIDwz68gsJoWsTIl8Iw
34+XebceSbcKS2Exn4k+WEMMvMt48lJzJbu0/kribj3JLAnWgAfXPFotsm0BHWMvW9aeLVT3rCTu
eO6ChW8aCPIT6p88VOEvLDreYwlUVHmvT97bZD1OJiXIfUokKs9lIzdo4wbiSnRwIux4nBMBnCtM
4jVYbN6t0vnZIhswnDfnKmb4+HxPtN+NXbd+4ncN0iopDa6gv5lapmf/WhQZ8dWCY6dmVo8paSoj
pihKroGPq2uN8Nw3dIsZUGuTXLMqEoaXA8mHwi2BOoFy2fepoCcfd2WCZ/5/hKWDjggvgs7JBQ8h
Bo1QvLKpD6xvAEF/ySYF1ETwaYnwZXZLR00rT8PFkh0YykP7FHbJKDB0X3VezNZvIpEBjPdDFO5W
8zh0ukQzd8omjCMJqnP55jxlUzCfeRhYMJLtUwzty3m6Tk3Jx/yZyBoRa4bmyCQSLVA1bXCnWO0H
F+PyKfFl9wmaCp77UaJ+c2sLGrOUI/IqhauCCGcpItuq+tEoEBOPOPwAc3Kw71SOJOHvklI9T219
IhAaw1iYc+X5ISK3lokplVLEv/MkvqDauJk3t7TPojHRQiqI0BkQQ4CLzPhUIxplT6ruGMBtrWq7
qGKO+1MXZmzWkfefXC3d0NPBLlCihe+aREoR2g1yvCUws35xYlZ+pJvPMnShqZuUDc2K0gnAuUaH
rXChtchoMSQIBSYeQosc3b0bdWe+jL8QZMFq6AmrQLXn/D8q4hth48wxJ/Z7fyqFbYg8mlIb/A2B
2K5FZZh1UgLrJaRBiIrpZorP43y2PVMKzqDFceu1T+HbEnIlVq96trFIadFwK4tb5314jH5H0glG
5MFeB7RheYTqYdpZZcA8eFYYZdcJlMKIwMZeCQm41pAynJ+uFmRcPS+RoUhBZfQgDF9rj+p2/OQG
u1LUcRMZ4Tlqe20FKhFGp5UHi+i1AjnqcGdlGQc2vynz/79Q/LloAcXDqwP1TUnmV3eQGR98j1Zi
/vq5KZhCt2CGpJNSzVma6EKMCJte5zqihakpHJe4pntYqI3oy2cLs9l7+QwM3RaPNPpAaWWhMPOw
8uR8U68lQ3vBAn2SC9Q1fRfsxOtAYQCEJFlqp2Bq7Ka/uHOcHXfydutqaPdVFRVH1zs2HDi3qxMm
1j5FxDPVs8UnOTuWwliP3SJOv/ob2FPYkgry6AU7cQV4EybaM5DvbicbfYaj2TfrDV9aAKDS5L6q
MtqYgOD2j4NzHJ1wyEcRGjY7znFrcFFSF/q4NeOb1XxfPnDY/35cdU38OrNvdG88biVqbPBCujWV
lqM9u4eltZ57BvxZblo3MqAkqniwvmNZ0gix5g0w/MLeF0O/+yXtsTYIRdmKh2uXd+Dy0sW6+LW7
IVPLM6PyJuG6jl+0CTAbMFaM+v2qUQMcpVN2XNimn84huQK2pJ0APKVWkxQvNk91rNnqv0CF+utG
gO9wK3+ITOjaJn6GfuXATHxCC1hVPNQO5fSPXoR0vcB3HGhODqn+NOS7kMyodY4BCF9mTwK6gYjz
Oq3WjlIavTOr/5IGuXulkR9Mt4a5AhOCw/UTBokO1YXsGH9nG4p2ACjIkkvCyo74IxAUYKrWQU+w
OHPbFv7JhlsAcxge2aRKo4igObf8uxHUbHsgFoQ2u3C7JcAt2wojAW1JxhGKzFXqDmHXSJbs/Wvi
E+vgtTeJNfcWnupANlwrLMkwEJGnLUWrr+SW4pbTHBN2HWWYw3nX8stb2emWHbQTvOPId/yjHZDI
sWW/oVA3iGigZugz/J5FDBkz+Kth2KRUojBtWxxw48mEhlesjCBuv9MJ2MDfLHffENXuZ8cdphoV
mB7MBmwf1u8VQ6A6Za5NB5ib7mvdWyH+SgR1rnXsMSPguol+WZvVtVGxrUOq3P3BCNy0k/9GCC5G
SBkLrHPBmytHmBErAqxgL58BhBTwzIo/tk42KflKieCZ+eLsiPg7hIlNUrNHrOneNnJEsSvxRdnP
5yzIC6Q/OD/l1A5in3EZCOoVl8e2q3cNrOGd+/sfiivmewpgAbL9vkqpB5vO3TXMqcKd7rsUqqSg
ryi0ClGqKxzawJDRobHjZZzFGZ+riPpk0g7/Djh1/3wB581Es5z9WTre87dQcjQj2G7Ud/ZuWwSi
fFHTa/v9DrpfrF+U8sWZmp3Octv+VCojVZMkbaKeiKHg0mw9TXMY88UhFCt7UHrsZS3Uu+HBUb3j
JMoz8puvldg1T0t7kNoGi5Q16dEoyEoLhNEwcq+7VM3oZWdsUekTwBmNza4TZ3Ujat41Ck4vkZgD
ZSgPJ1sB+gxZzaVzA5NyN9nxBU1OgFBdr2rdS0XgMP7uYX8xiUzZ2pIbBTeeE4mF9D0e+cue0VS6
zDz0pH5KW7R1m+P8GX9LGFUMZLGHxfuiQGU81fI17kdYcy2S8eqC05bOKTuw7WcG1X0StoqCrXML
oCr5Wxdvh5NhHj/8yihGwbjdHyXk7Tl0r+yG3Xy4ohsjkoeZ0PdtTngx9bwSj+D4mJblh9lFvbtG
vnvMnM2pudSA3zDDGRBR5CZDbQ/oAzcq7gYDhqF8+HJu1kKDS/6i6yslY1iyXzQNLubNR5pgAG2X
IRvKi4IuY4TQSQ4fsuuOYAPGQ8Tw8OF5c4glU6SE4J6fEFQTGySeqDhXqpVaBE4X3pfm/P10F3v5
ad7RNQxvr6x632vIy9YETpN1qc7mFqPinn1NgVEXpdpC+B1qqP/+8Dzy4ll7IfnNAKOncmkLopM0
41h3tiII6EcXvkTDq8xjW+ZzdH8EstO7phLOxmIAYOcZtMDu4Zh6XTIGDcaq4d2VHLJaow0nqxlh
vtlhtfy9pi0Sjvwl01Wyyaa5UGJh4H47GuYdr9csYU5Sigx7wKNdJxxvCwEG1FImhYUPeX4Y1YWf
nvHLIt8fJiimYnD0JrqMzDRSH+hyka9St0TZbeHjB+HCUal+BGs15M5E/RX2kPNZFARf7sX0Jt83
8P9Z129S+D+4yTPaTWC/XDfwERhbluewKqXNBlt1SlslYuYRfGISo03BXaKFBzAK69Lr8Q9M5vmI
vHp87ZzVuu5BSjeDQq7RSuLm4j80zfY/e1s56iV2Oga+RaNTN1hIGVYKEKSX9KQ0y1oQzL62utNU
UQkgxUXeToKsSCFcsKQM098jZYIPjS1A/JRMi2+C2EH0ZZUTvJeTRJwBnz+REN5mq4zKgoGJikfU
Yry6xVuVabylZxlRVrLGTEuuVuEhrxyPzaP2R0lkSp4JtFLWrUF/EGm9IaWkQGXSJdmt62U5FBqy
FPKNhoNMMObrtvWa4QQ5ERc8O2HRWce8ShBKTj2rCXOY5w8Q2rhku5NMCHRLWwqzXzPRokR8YMqq
l2qvjh+xuUssQtFYtXWJgI6FqTnBtw1pIfSvlohwPeKJqDIKZekH06qcd7ME2Ufda8XsVQscS3HD
UpH2JYFVzoDgluAf0axb3QrdX5omIDgyUa/gsx3t3efACen7KKIX3ypIEyDs144dkXhJfb5CAN62
E0Vr40tB/RhL3wXv1RoGACZtJ22z0rjUf5GxJ0s09cf4IPDfixhAkwb56gSTM9NC02DWNIuTebb2
DLhX/zGbm1pL2abrXbmS1PJoWuPsqM8CZy7U0isUAgEFGDP5J1lO+UBl3yOJgKeapIyDfQc1SMso
RXlOWojZV9+mnmry90NLAOC9SYC2V6L/blvLPwm2hnWtRV+dqyhfDw33dLbCZA9SkiFD1MILsA50
GbAl1mIkv7Px2fW7CgumSxoYk5T1cIpvyFVHDluU83z5U7zuIHGp7cQLscm/JNgWkJkz7WF3jJZy
IavUMhzTGoy45gRAdaKPzhLXyd5fFBW3kB8yQB4NWSRjvxRwGxcFqs0hTu9DalErUgHYauH+T1iO
P9gAT1xT1hQd3PcrJ1R0N/2nZfDK+NZzcl9WpqVmWrKQr/uUGnDk6g81VjyQKcV4GeiV7fKoQBcG
rRJIc+R2K3K+KBYG/Fuf06XKurHZGkHW7zlGxOqPm3lDU4TJd/AzYDmuJK7XS0PIpcXhgAwxZm/w
yK5J9obNpmHk0WePVoz5xWKLuaQg614AL8fbaeNr/xSRH86D8+9ikJu6WnNae6m+hcloQ6CLZyJQ
OwHXeW1YPea4CT9P7nW7f+C1TP/7qWrCwzjJDHaPV9Wfqb6fk0f94YIJMsHIOZbt16Obk3FMaYKt
kQuTtHnJ5IOJlcIcTe/tUaulBgPq2yK1yMgavY0T+GryVR4o/nDCWxvvB5P+U3t0TzLaqApVlfl6
Sfa/Z+KPkmErSqQvvTLv0TK5rHlyIWqPS8V8G24Z7JxM9G+bsOcqS1vEeqYVGcLnLDg9RM/+peOE
V0PqKawe6VtiB5SYeAEhMjJ/pgGuCycv5Tlwr1aEK2/zmE7oRsGP9f+epiXQMWkDfIhDLYEMwbwU
DRCLbLJz1mma4hv63YE0fcEsVhPtWVHU2J/G2V/J18FaMxJbDeXHjecuJxk9lMHxa4x18QhqFJU9
C8NUSFD9+PQC4jd90oQTAjQdPWhj3AKi1kb2l1yHjWhTpAk4WMv5+wlGr218laCNRd4XgAH0UC7W
w3/cNhYLG9S2gYRYrnWy9Iv+5+24miLd+2PdCIcrSQrsjwh6WWVMmAsO1Mp4BcGrCIUyF3/MJiZi
65StRSWdoE00dYL/Cam5gYUY8eHrW24TQekNfbeGbyxLOPHvNayfrPATn/rwA8F3z4QdfUUZyT9c
BNdt3sHBKQ+mJJ4Uh4AL+/GclYxysyV06hxtBEAH0ujN8+dBK6dbKnrMwAZxYQzSFFNo/BOIr3+e
ouk5cCKlB2FwVZV6pRDQPRsLOXSw0ycE4JxF+ZL7IlRzcvrSdS1WUjeKz8TrkajfE8JPNB4b/Zyf
Zvfko2Up2cFarSfV7JRJphCOf/DBgCqHRj2lEdAkYtk3J7TI/I3RCGIcdAg43GK7LLgfGGDy/5O4
IKoxo3h6w8raUPYdS2OSC8sFbVWU+xn8NVnXbdgOPWWb0+3SjNJw6GFC2m+khOLTb5xcYV7kYPlK
T/bXlIXkJums+h9K6gvnYwi4oHGAb1yj95JGl1IS9WVajGylV+/ptd4RzmlrABw8cYCjcbfgDdv2
DBZhhtkfIx8Hl8jsEpItPYIhTqDc3F5NkFFqNtHbqRAy1PMnmA1OAiZ2I2tzgBa313qFjf/G1YgO
qscRT5h+AVFs6Z+HRb7QYdjjcGXwGpX4JCaFdwy2pubFtq9vV9Xgw/tzBz/CAYWcITvZOZx7TU07
Aj8uLK9HfYOnAhbNyWmGx9SZDyE4G3eB1wl1Bu07sOVkmCunfkhXoWYjvKoiq8GLIqQw70tgdZKO
dKa0dERsB8LiIv7u7wGaaosq2mr3TdmBC6e710Mqh8M3MtmkhI81gBLtk5ZEQGxUpUsKQiW++MWj
30dIRKy5Z65WTbxv5O4urNCYx0pg4b4PiAIkfVVSwhmwHkI8IKxKGNr4IgDHpDzMfdB8X9z6LG96
49p4eX4pVXnINeSs3Ug9KqoZPFC3uNQiHsa4qx57kh4DZ1JKHovJKKskArFLRN0w7GYmUM0T6idt
Kv0PI0wY6eTioB3TD0frNh24ZXyIk3fwVogqLRCMam1cXywHbrksYjYY7/HUACs+zfIcy+CAKZte
buAuRy7s7UWSvUZJJWD/eKC9FebmSphIUrOwAXU+PQhYhA1opRwrJEQEbvR/NKiviHt828QPOApN
f3Vm1FnBOmGk78ITVVmH0uS7rBcxBE/XjN0S0vLnyVQGVnAzOREd8Fpd+TV83j3ZzFXuvaubHXfs
vjpaw3ZulBjk9TNPkzoJqxGbs53XPJrC7wrNyNS34RgSvilDbdUUFyr9bhAgK2JRC4tJTmTOKBjb
Kc3BL9X8BGFe7wJPimkpND5XOG8ppGhyDgNaOdAvAZPqkAINEEtrGmhkRBFFwyff0ydJnaK0G4oI
L3fCM+Lso27gyGmUdmtsEAqi7S68TF9FWT1zyK8cyglBjIw8tqiKweqOh0Ta44gNVFCQIEEXr0fj
zZxHkqc17ZLJd0+2t0dkj9Eyned6SYBEeyKUFUJvhybWHfbA4w7Z4OfvE6qXtnhlaRguZ0c4XLJ/
nyYStT78ZyLele8BeP3nzVUcDkdLX6WQLPEUpuJnzy9GwBfnIMiAHJuxbGBn64VMQRSQpcT27jYw
i1DSuisD3D/09HtDUO8IFwlQD0dQa/Pg4Xw3+gmJgRpBm6Q7cpI6d+8gJwle6F6tZIKlRF2WYq/S
Uj9Vl+1Dw/31RsBMynZSBCDrcH1XzdEiA3O3EmvGTjaX1FdjFx6+/FMmDdNER0nYtutJlJb7Awmn
Gwoolj9ivQb1jKDpwnLT+Rj/r/i2EoVY6fV8OJLuDdQJoiBJfcaYYPV/eA/FPPJiSeomOMwA+BcH
udWc9aW9B4oPjxCHL6EopKt6k3BncyIGcfzlhiEP/E4/TtNJ8AgCaHj8ZtiKlOsRtdlGOSUOkkZT
zyPuMoIjZdo20GBm1MCgQ1JixQksMgy5B7oMxbe4UEl4R4mr3d6jnwk1qSZl2IBSXBCXr1WalCwE
kI3HpdAAUQ/ET7urPQsN5ztVU7K3DjNyKkITDiSzectQn7fBqLmf7FmsEh020ado/W883s0WQ0EA
v1K8Qs81SBf4tR2CRTykqcFVbO5Q/Iein7Hx75yA1NE7z04a/QZwbAX+q9f0JQffcDVuXjJXGqAc
IMfEpeJ/5SBVcSz8t1S94DrVWDOq/+HjSVZadEi1SuQ4j2GyYrF0bfpyhPDEgh/HI+5ezA/CZKQ1
tCTWSJPtYv+Glq5GNreSdu/kDPoL6Hs8qMEK/540Aut8UgJn7/6e7rJrHI2IbcWwshnfmMZt15f2
4CCzig7SqQw9lqA0wFzWz6qSizSgK8mtZZzW4y/zEKaGhUh58hgwraQ5rbi90pJo/+1DULeMT0Tb
ToM49IxrRV/lCl8jYyiPe6ITqQeR9FPJ0pJTn8tZ4jfQBj1f9iJDRGJIvrDNHL9MddCS1i7nFquG
uqgI3wKJdM457VDJ6sjiZgCMYvbLkvxu29R4a8PxIAFJaI+d6A+IjDV29lj+L6A/l3M9+zT2eDaL
FP6lL814xoavs22xDIEYxbueYGr+VaKrKE4jcKxuOMGZkvsUt1CWEtQykPLF+zMwk6K+exTEmvDv
SB6/wgPZ14BcJGwHrSilMHWiVbXocKAn8teVDdKiEp+1QYaNGt1MY5HYRIS95hNaTfNHaZ9AtgsI
GAexHPGPNrsPydAPyJDy6RBwpTNlsMWVfSAILq7Z4M1yYinivTE0NRop5w/FTCSQVpYuqJWwHp+H
3H/2c94uN/NeSPDMDMxbBgOSiPGEI72xAsuoIKNpJusVKBcJ+2DOkl80Y3e6w93AmuM1SyvmGOiR
NWjMsNMuF2omKJwf7GjEY4QbIu5j+UqzCYinZfMETrzfujcBJmFB9K6JA4AUj3B2I0VKSZj4dVZD
3woTxj0XeJCvwA8Fn8NSTVOuKvxwIBiaIXVD7cZjIswDzlDlJnh5qAuMP5EhOw51wEm/2Rhm7ctp
KCyh132s8Rdz7t/onRNzdMsL+Vq/Cg1BJWdhDT9O4zabhEAGEXyqiyKXnznwTmMctJlV/Fw3Dgkx
El749Zk4q6udr6zMLHep/pFLignGyWNBLkf6Ufsp8LAE8qY81E8v/WEx20sAulgppcfvmj3gXMDo
kCdki5DXtg72UCEu9+DV7+1VhBhwjPsj98rejaDDLrouFtJGK2zCjKyzyAeKCQRs+rO780Xt1OcP
+JDPb7tK/v6e7a/nagIDiDVBszbqAjORBllVQsQ+SyWUOV6do+QoOO22attdEmF/z5MjhmBNX0Q7
88aaqwphh35QtL2kAxuxQvYdvN6NCuT7hPwTvWKlL/KWuAF9xooThgFjP2Ej8IG5dawo9hQY0fqr
LL5x9CCHFmqoWQ6808eRHlJzyDQTfj0c/A2VePCtBnegRRnHo3aEp9XCB047fq5YDoY+FZZCBv9s
ulrpdsHWw5zAf8lPGCnFdbqMpWAgsmjXTnyxuAeDud5KwkGVBzlrpPTMTOQAF1CJE5sEPVZ0jhAi
I/iwIEZDEKZg86Ocovq1hCZxrHvXRRJv6XedKPTSv4B93n0hLr0pVhI3dWlfqsracOHKwuMx+y/E
hLWzpOReLFucU9sIS69/DF6FvjdErHp+t2vvD9VFGJuT7gDE3zj5f86Xb8I1Egvg958Mup7lfdIZ
+lsKiiE9765oqEdtDY0qFJ/uV43s57gh6IwsirdqRtRJcbYeUAVzZ+e/YzcVBudOCa/V438PnGr3
Y/QEYd3oSQmBJH9ZhWTADUZqyAMPuvlwQGbuqcmu44UlkIml8MA72UoFG1VL20w2gnp7QaHgC4b5
YRwnzRLmMjoEAy9IxBhhdhjqHoQ/wathbfuO7zMKNe6yTdFyWzJpSpfyz+q1PD7d0wXEcFRDag5h
GTJcL3in6m097zqZ3AaIwp9Js5foEkQV2e1RnLPl0++x7Pqhdby3n0m8H4Egljd9yYCMLamwQwPO
FgHk19Pc7t17qzx0Krng7jYZA5k06gWxQBVLvOrqXFHtMOle2Cb4Lz10vNz9O/NUOMVun0mc1mCh
xji8mwA9UCf+k+vMijznxmCBr84B4TTwIte/SeXhxl1iMho674kf+L9aL/MOVfdrLW4QHwb3qGLf
NHUzPLTJMQFUXAQ1RMUQgVkTBg6Rwuy9AN9u1uFKfYokOONIw63mhIEb2mXy0yIDQ12asRIzjrcx
L3TiUyYtIUDs/4w3U+gz1lduliT2cmQBAffttdVVJ1nRBXkPdlQstuNyFjsa7Bzsxl33ZtdRHR79
jzamOkveKAxTjM/epJyBUM7mjTEQm7QZ6xFCMAFn1dJWVDB84nV1+TS6yjXKmXpVTGo1sd/Wiwly
7kZ50wL5zGxz6M118J291vG7rB/ZqXAUi5eW2n4CHIQnaar02UPq2D+RB2TejmD+92y5AiC4O9Yt
HTL+VXqNOMyW+QVsnWZUHGq6k+uE7uePXYXlswORog48pt1NoXAXExGl86frr/NwTnUML8fyIcr9
Piqj/AhChVtcNCxaM8D/IR5spR3uaI6OpNMfeOCCIWHjJlJr5rMznO3FMRYEScUz6qsQYSLSTpBP
n+KrQcjLyV/RtZuU7VzQG2ykswQcn/CmK2nnumDP1x8ormIWhfH/oydjClmeiR+MIY94abfQRsJr
n8mwvjWZzrXIqTugntkaVzCLoZxYoJa5+ciFix9CNTwK3ozy9FBe/Bqc63yXSgTqa3MjlEV5ArzI
A2u/sOnXWO8JqHHBT+lWZTCqTbrd3he8Ih0jGwlcA6rxsJUScNBYHTHP34D3s9q/9yCSoQeoI59h
QHJ4YT0w+T3bhUanoEWGXKizaERnufAJFxwoY4MS8dSciRCwTvniqy2LVEhmlVYo//EzK7tbE7Yx
nZXdYudmPmx/wY8AcA/hl/7A3GBKCvRa5fwXwzwzkrxqyINnSpAsj+hjgd0ePFUcB4udVIOQZd8/
qUxDG01gTwC2yLzdEnZhAT/uLgi5INbvyZTsYU8tlKd8napjrAPlVI4rI2Bw0BvbOpB36/Qtdt0k
JLGafjRsaWrHrICuC55hPZt3klOuBrmhoMY6PbDU7BBT7Qu68JKWy7+uy1rq7EYXglA5UZjxCrB1
9FyEkSjJFmrrVTyRxoLpyVzN7Aufyy/5u5r3gOrqHHF0BCnIpxUHXcERTQmP79e1fLbJTg3ryIJV
/vnwQPLxVieM4/IkfdQE4sH9b5IisHTWwS5CHendaeaa40f2ZQZt+pOUlI5FhKJarL+r120W+mqL
6LfJ/9FJTvBn/cVbmO12LwMlPE3TpYxFCyOSGnK3QdCpLJZLBbzliqvF4dxKxSBVgDHyC2CFzofg
AwrQpqhGeuyP+h3U21dgZ8raPnAzOzgpBxCOUtSF6dCxBZnmncy7G0mX0c5vXa9S/mHCeY+PdILx
n0e6LuRi5/vWgmTYSaMwthQbsdVoDH1nW6pxavZlQNWdLWuWm0/BZMQQjab54TLmRU9s2qaqZo7q
qcKl82W74qF4pJnnPl/FgfGls6fWf67AeJCA+0jt9r55ppsoobObLNb92+YdEz/AZ47pjo/MjvNS
mxb5VBHAHFaMQht/NI8/y3adQp0ci8/GS4KWY3UiKuFGIEzeHBwYaulS3CuIzfCATJZakbIhgz+U
u1yXu/TbDhi57mEq6MoHL/vhfHK67pM9E57PR5YEeVrOGS8h3ODBZ6/uhL02KjrcqKMDy6wV4zXe
EXarNmNuXMYHl5TacfNOhyEjSxkPaWEM2iXuqr6HaxKwIIc5asCGI+RjjzgfMmgZZAK8ZmSVUmd4
KbIfz3IBLhNo1uHQu5WXfY1wfqS6aoUdkbdaDE+oexvaYIGVuB8aBAzFycWZsq2+a499SbnUF2MD
oV8Pg6sVOXHHPtSHxbdsoc6kOZi+fGsEZE6hPqXc+/OGqXCcXRS4m0EtcFCXPgAMquLBTnewreHf
v8ApA0WODLPlLA5nSvJPh91YvQLZc74eDBofoL4N2ElXC9h9bhsoiAD/uBZI/2K/d2dLrWTG72ZA
2/otCg3vwDm+kOtNIMg8pEBPBeGxSxMz3cY12VHgL/oeS84LHKPEUqhFqZFzLFH7h5bxusylj9Fc
7qDRYeb9g1ofI/O+/+CHoNPqxX7P745ypPlvc+PE9J1Ijkamm5ScD+b0RE+sFdf+7hvbTPSnus5n
6uF+tHCCoJRbXnz3ZxYGxuDwTyJvju1qxL5fPl28p3qZErXNuobXqSn0cSPOYjXjNbMaJiDV8KLs
6pU+F/RBD/SPLUrmjBv13C3Ay6I1w/1uv4A//LPJqTA9ga4Xf7OAk76UeMrq39weHs+am9Z2JlO9
gQQ8mgNaOSIcRrfX3migWRUR4xzpa5W432Pdio8NSRqmbQpLoWEmQffa5CJaI2ZGQA8lp6e2Vyf7
wIRKYn3VMYJLhJcbp+iRn6VasoxSm3JFdnSrvH2MSb6yduwKDZEuiV/ecRnAzj8hQFEWQ6z3h5VZ
T0xWkZ4G5jfRmUUC0XpiWpqqQiaS9pNXpPTTUTU8QzFjYP9O7OdGw9oW6iAtv5qh575n1RSFoT+Q
ZLMjMd99cPy/qtfZS20JfOaih+yVz9M5EYWwrHej6sFhHVxrr+RCkM14p2hFs23P0qzylj27QWNq
QnEx0TYQByXBNe+AO5X3vtCNVvWSuF4W8na3oiunR+2V882/1n/GhJGY5hCWmvF6hUmnE820nKgD
Mizmoz6B6m3LljOVj9TgI1RVcrtGHpcal/Li0VwlX3JE2hg5mham7n9r4kv8k/9uYMs0KQVj93af
L9bMAHA2aMYZplKOf1MGWq15hCcoiSXmYV+RugUymeLntwEmtGq1eyesq5/ScKI4OxlB0XkMOJej
VsNRKOlEfWretyo6hkaOHhEvlj7tISc1q/Wm+Kb+ovKUT1PiQ9njUKf1TIZFXxMqMWVzHjKSsSDW
XvzFp1jRGoOmheoSJESLJzGHPqgUv3NWng3IZQrOcz71665tF5qXJK4JXNAXjEg/DdEgYnaIp238
kKdnLZFDWjPFAmh9xiHzHNSEia+oLiax+kUO6wu158gD0O1lDsHSailNNDLVVMXiZ1ccj36bUGfZ
/zFc+jCzPWdp1b79rpXysDCGPrKnoTM4OM2zGudCyDloQkt8GNGJYVpMZg2kPhOsJT3Sq3C24JC9
KROPUJWzsJoxTFV0KTo5jbbHKzndwYmjtkPik4rG5VXYPPuymMtiWxl3oT4WM1rmkZ6G/BA7SiBV
81sBRp+bAqYYKL7WTYDF234ZFU/fWpUE92Wg5C3onz3wJK5hOs3n2kH9hm0/Ocl2vsGLbnYT7xTL
EMTpNlPHXQjzGGTcpq7wZepfO2DBdnaJO8GxclN66RU3shu4T5neb9FtoOrIKODFzskwI5vKpVQB
c/Ih9h73aNO3fXp2hIclM22ffE/ySk86PIZufd3JOWsGUR8bMYc1KrHvdGkd8lHg3vlr5Pfjv3mB
dVUPUWnWzCueCHCjrGCgTFA+yRsaGeGvLeqUJMHGUCuk6mHKgDpjqFWDkvflkqvPtds/F4ULPUAi
e9a+eqMMFt4c/inkpUBx4zBhWm6RX/wBjFuMF4W5F2sARvIYTCOTYQm7cmauBN0GqqDTW1XK9GfB
B4NwUL5UzbWOK8k4cuQgMMtfvYXBrY8WtXhj4Fs2TnD0iqepDIkRvNEz+uvO2jKihutp+2aNv4rt
aS8EzbQ1Eq7yH4e3ExFxAIvsw67Vsw6JyUIXpb3Sn/R9xlzQu+BNcFzn7y/MLYwSfL1Y/M8y06IC
/8DlU3guDlHtANjTUigXNMA3rjduCoAG2LleSV357HK6yDtzuuYL+3bcUJN2LbZGI4TorlfQM3hL
jfJzxKSMNNcyzq8rl8tp7IEQXjklGx5bYs1Kbx6E6kpbAWu03WF0whCaI0+2KlUOOsIEnWKYMn59
+Sf8qwDpfdqG06PKMTArWIu2xt2+CxtMzM4SAnq+GFadYuNYx5/RKEZlP9lp33e1Y6y+p7lbIdgZ
TA9Qfa2L/TCAQUKAdZ2xcWQkiPQzVvNQFja+MB41VDYqriXCEweZMRY+xab6DMPZqFDX8V6YIa1S
C5IBtEjLYxMahJPv/xhzSetl19G/31TnRO9XlQ8FxXc2d470xFK7Y17OwoirTMgl0fA6+jzHDXEA
TI0344z4emxNOe9AKzElWDRTByVS8iXEjGVIotfEx7bI54bU/PSvlJknQTwn1hkFM28yiPOPIeuF
VOvp34LOEw9uG1qhUzf13fuZX5eYSMSnC5YrtrkkJbgWIBITe3Gc7OHFsT5QE4hGAieDzBRFeGGo
9Y51Lya0RT0j1p4BmbUdvIWIzpgtqPp4J9AfzuohLI/rh1FSgdwUwtop5dnzKXVGXHwM80WWjSue
Euxr/RYwdCoObWqWTrTzazz6VPGU+X1zIjyTHbAWwT6YDozt1B0vVEMxlC5OIq9E1BqAPcnpT3ua
3Ltjj7oE45mRntDBMw0Mum1uJRbNF3xUajv3+OOb4g0zJksk+qU4m0Y3rT5ILyEpJ2Zc0HrD54VW
y2bokeAM9gvutDCxxOUkkBsLDGPttwTw8Rj2D3vrZObNegpNmFlepqXDL1j/k8tz/CD12M9/Do3y
wtQs382hyre46pTYP6xo0TFVQxI/YJyXQFIacbhSIFCjgpUo9iPdar36fMO+8h6dhLGIUaz/Y0PB
4iLNAOG1D4/LLNV6wGssvrjVOmNdjGLRvCTZ+Z4nMUmYcn3awWkQ0G97nc/2ly5+av+1UKAwAiIm
XSn0ybDeBA1EMaNj3JUvW92hb/oVziK+XdbgBL9XqGesWgYocAVg/GZAvqeqPpID2fG8p5t8vNrA
cEm4w0p0l2gZcyMnRTSiDx8A2dqcrO29c/QjZkB2SL6nXr72m8M5Ds9Ou4X3gwLQ8abmq/D7bW7H
ytGaEkGU+onxww81k8Mpxa+WDm79nT3xwPeerkediFUc2kRqvmGW017uTKOxKeYWEo4s2G+kcqXV
zJ+TOs/Ng1wUPWYiD9AlpwZhT6nalGkxTr8O864nQyuOMIQyGLJP8146t+XuLyHcm2XgvWvIi7Pi
/Ibann1DQktcVeUH69O2Es+HT28GbcvBorJbB/RxkWWXNnlySEG8MwcFhVfEIgzRfIUpQ1XcQVmP
QFMuaM9opGhjKyOjBNp37mefxOUH8zwso/wPcqcv6ll5lHOUTm75tfYQQlJ3lPg+1iKFknvC7ZvQ
YV01z/At0E1ktBQSMT8sZPLFGYHE7IBYTsu8DOVMaZMQttx07Eyc2G1weBCQDBoH358oJ5bCp/Vw
sA6aqjLZmjA8u92+q+2arpKAFuezMdq+2C12PE2b6kewq7svZEUQckCMkWbaqtrGwgZOc1JJKfSy
Ot6MIuHOELAClWJ53dHJHDD1kJTCtCehrbQ0S008YK/FAexRPT3exPhg29tOKjIZXfZ2Su+/xzNv
Drtsf0YQeSGpUQuuiFYJ7d7y1Z5bHaflELqC6NZehVm7N5TYm96syH/6s94HrEbMLhFquK1/bvs8
vIrg5tyXzqiUONE0QYa5d8ZBO3a96WfOJF72KIrzPquBVd2RYxa5p9Fx1x+RoFkjDqpORj9DJ1ct
ufpWt4oq8kuiA5qna/oD402UUMOnwwYAqgei8GLaJzObF/nUcdePENt4IBFTTgnuk7blq83i2pU7
3S/328ASBU/PkYVhY9Lj/9/tH1q6qm7VtRr/t/VcuPeWxM7mnM1a4RApv8/+v0UPNUWC+GX2UGYb
WFihmPsb7K4vO7YPXS4rxGk/84Y43bbaWpD2GTNNC47ZZSrZ50Ty7nWXZFguAAjRYOr+66QPk4SL
YRU457HtQ+Axq2BhjPFwIl27BCu9TkXfbWJzfAKC+gyvGNRGB+BiN39ZY84cvlj4h9pOnqESKmTx
AlikTqL0W7uxohglz3zOf1LVPCuxGp5xv0YfD9BzICYf7Tn4lZWmfSuNdSb4R45bbNp/GdPegPaD
DMjBi3VwXNJJc/rcUvCvkIVeAKhIqz7OOlz3SsL77PoWKdj16RIyCoJvdJgYUb7bY2tmaKuOha1C
DHFFEkfwPo0Xg58XSHVpGKYiyMalgM1X2QWszWxepi0d0q27Bf6DmXwyPV9pZe9XbuiCbJnafJXU
beseBDx/nqiiXs8lAdCLLEUMgZTNC5nphUK2ehdB+mG0bKf1KCc5Fl0ylxvKXkLjY/yE9NFKZ144
3vw/nsCmK7g4rxiYQmG33bVldCFiaQ9MYA2zMjBAFxWUnecKZRwH85D4G1yHFjQJIeHMo8K+HWZ4
HL2zNxN9HtYwD7YAjnxRksysUMotPb+BYXcIew1Vovog/Dt5+xSKofMZHbaxOh4b3/xyAnGlTQb8
MEriOm70A12ac95bo6yMqBSrrzUm74DP/x0GWuUdjXdgXvjE2WqxoxqLrxP0KPKS0S7/kn+w8LVO
BgEj5rGFH8UfP2+PY4ZA0aUsebZBKgcneyd+U/J76u63Zv1kQYa8h3uC5j/fOy9ijuWVbIo+d7Op
EKEz19iW4ZcM8MrblRLISimoenSlgdo3W3tMcYCFmraj2XosBcmb2s1Fs7FJSeLBc9uWid1v6tHs
8Wolahh6seyFnjW+In+WeiRCmW1LGhxfOZINvQTFmVHngj4RqG8xYzVLRKTN78NHQbRcmxZ5Bttn
GS7OsKfuz+uIvbjdtbeq2XEZrrM65lW+pYKA5LQKZa8QgZ8Uz5vmclipKs7gy2s9sPq3GyxgTziq
Wmyd3GI2X6pDg4upjmyVxRlE2D94/fP0v/5USJkNvDZOkgouf0012ihYoC0xgQzvfgpsmRNjpPv+
5uKYL87lEmDipbRy63+m19/5lms4RUAPDZazrJCZlXRGxM557T8RSYq+h7H/eDyCFaZHfo9VM03E
70w7ZQ1WrwqyR8jMxf72XwxdZzpoeAO0NH11+kS8NyAWFqwlIFLbfeM2P8wjXgO6NtZ/yCzuDtM0
5AZA1rurSZwd5tGQbr5+dwVyTD/OfFaQCEsWZ9OhU5jyUTb09Vymp0DoUNEg5Rzqi+BPk/5/1UKa
T3dpFj5yHZvC5pJQDauclJ08p6ZL4aWDC9Rn4dH9ARj1jE22+uLSr7j38qWA/5FT3tCagepdH8Ea
2uTHZHPSFXfE/1o5IOn/50c3rXWIzVCNvn/cSB51KuuRQy7+CmsikNl1bAp7QfeNVz4iJNt5armQ
owvN0nMoAwjoGZpo0TX04WOVEc66V5dwW8fIF6JsCLKnVyDD+/5DxA7T71sR5Dl7bBv03QZONAki
6TYekZN5v63WLx99x3HDHISj725FD1amDOhUnuF0vSsO+Y7qf39F23JjvOfeEVGazaMo6ofvMf47
xf1HKaQQg07SMNi89nh7B7Udwo8dAI3L6p/67JuVH1WkmxkT9F0Q9oaJWQHFFygaBc9SZyR2hdwn
e98lqthRwOYuy+4ED1T7uXVVbHFUI6zAormEAKe82Bwnbd7V1qbE5ffdXapPH+3xXQK+jf78RQRW
QNxBl1qhf/4lEwUghl8x4rFqESi7TV8Bfp/uPezL5RwQp3npoLzCfXdyyunFEw93SKVneFSBbWJ2
nlEh2XYt9CM2uSDO23Z6DMrLL1kpzJbUoMhPcV1aeHa7U/IJKPrtXljsjuRzX/jZMzXhoEIj49a2
i/Zpe9dzbbuH92lI7rMKXoVX3GAZS1k/T8Dni/Lr36LV/Ltx9WFkShZHGfOdhIIppkxTWfHaxEQS
0sl+RBLC6nxWcU/Thzs99ibhjiv/y2GseogrxvVHtgo2mwN8elUDLK6fVgSohV3aMIDB86liBvVQ
LuicIKOCaEJ7o+6JEv3L3/jik2Z7d3pTBXOwn/g5Apw21x+rVWC5AJs2pmgTX48V2V75OmmHIJ4X
+A2rZl2sNL3ua7YMM9/kX+0AoQP+N6wNZ5cPH2pLM+jozWgpk7a7//BWu6feDXHvNBaS0mvt1Tj7
ORxuQenQwgvm24PVM5o8cFBYAFsIK3Ym7iMMmm/8+fF64I6uvY0wdvaUQLkoPw3+2BJqjn+O8KZj
WHscS0jvZ+zJrO+dco7g2+ZUKrLRmCBvUqgiJKIC2OVeaYHTaUPS6o3oYG/tqSppSDhE2YV6GJ0L
rTdB0GptnR7e2DFUT45cT0KBLoCtOHMiG+CoHHWJebC+oa6ViwgfS2xKUpCOWH+kaRy3V7fEePdE
X9C0My24JV+FxL6YK+rPmXUH33fqKgqinrztbx4OlDCE3byoy0Dw7I6buGaTk3ng0kCQwk4yqsKt
OpLFygZ1Pb2dYM1/ZTaSaperlnM99lP1yJbc1C1SKGzItVPCOKKBuVl3uZV9XLBKeorVgSfjZ9Mo
W6lLxlALE+VnpB2QdUBGgY8QZgxgCwdWAkN+yeB22KXvCOeqto0Fj0bVH6EMby+nrmewqAn+DNIo
6BH+03uLDSYC0vV7I0bkdGcbaYAeNNx0CwALDz2PS/yv6/huP2a/RlcLlQOHx6VLKbFpy4fl2YZ7
BUU69zt/waklikz/FqrdLKMpi5wxnJT7ZOVp8UgybLRi5HLLC9rYUdUT29J3E6sb9+4L/BO0C9gQ
WdBegozzdxs82eAtZZnegMWN7idcFAW6WuPIpsjWplLrMcwsEd4xFlV5z9uNymD+UbnqRJ3PdDbM
nrRQxx3r9nuJddEYJf5668fsuvrZxPkgyqEjSzFpi2tJ1JhXeOlWp0xPY7/WJSTfZXiJzDeFRu1k
B+E4N4yyOHHunT1/OZwC1ogW9v0hl16jdfic/Z5Pi/cdzbjrD3xsKE4ks+9kI6XRI+m0Y5QlFtVA
P2M4Eq8UOjBvOeebDV0w1gotlAUZKpCSKv0rs9D+JlDyez1C+fvl4EHT/huIDmAjFT3XMcg6SLf1
ZPyUd38XcBiRW7NqsuOt1QnmIOgt3b/66qZ9XnBS+SsNZD004ae7Wxa/MBBcMfFaIexM+ldBmGet
KhHelPs5Xwu85zARV++evXqj0EkAqBogMUB/mMCyzWHKzOQGEF6MTLDtNqXIb4BBsnIt9c4VfObQ
pSi+r3tPXsPo4w2JphVvnVgdNKsdqxAbz+MGygHqoMn/j6isKGFHV/rowwrlAOw3GpW0ncsP9oDF
cdWgdhQPw0hGOfTOX2Bzbdb/vr1IlpkN7d0ZnNIua0GwMDU5NXOlKqwNI4jJfzeR2quxBsqXX2XG
LMgwCBe+hhfodyfXgUiHHM5Bqo69TyRUoOXVviOtQyvSe0t/bLXMkTuV+DXlPwd5pZmatLZD0XI0
l6hLpMINyYk0TtFxhsYG3BRBxLF+G8phWJ/gnNRwKAe+4RRlYQ3hXTNwUwDDanh2ap0DomSLFVlL
+DV9CjLEFRXVfU+iWXu5WSepl2adtH2LrbNw48MEXkDbBC/uCW9dn5xLX+9SEr6anMJF6ROoCzmL
gbERc4PMVCoflxhxZNtWxY3IVbvIeQB5Z/Upn+DB6OQCJSsAoLba6b5+AnrKZQjxZHPjplrJ36Sw
nuf7hgql/SBhIHy7tpd8OY5sucasngl3hNEibsrUrBYWjWnnEeyJKoBW1PwcHE4R6V5pqlDxCt2i
ewNHPogABiiBA7r9xKUmbMpRgOEUdHJG+FEs9O5+brN6ENmYdKHcvbYj2wEpnsSSNURHsMJsvlvs
kM+3UZKC/eKhGdvAMiA2aEuOfXlSoSXmAF+oSorAKDmVdLrEC8NfTr1BuFxuFNkB/0toQuDLlOGi
80LH0ITHPzyEJRYKfOvFHf0UGyl51b7iQDrA1e3Kag89RFA5+lURD7plzYp1gINJRSUghyBEC7im
aR0AMmjhqbsIAhsGTFNjJ+I0y9grgftQd9KqSrmODaWaUakG6ZjRHt3TuopyPZaOH4wyfU1/Qafd
htQtUQBRZD2+hjNloosHKNUGNK2br/GaYPC5jVgeXQLRUg5M/VKPPsK0M9/aruIEXYXQ0i/ujyfb
kyrLF712IQtMjpD3MnkxqW0lgi/cWeUthiXivjvcv/MlutdCVmuXHNN3uvBKvPKzXmsYJuRZUGZG
8gnys3DSlT7mA3EiX92kbORWGPAgqkgrm1BsM+7Wnm2FvOSUQvfsHpD2P4wjPGEM6s7b+2KThNoS
ai0OaMYVBwncrAGDzMMUA+ud3tmRY58YVxuLeBgutUb5F/1sLKZrax32GztursBc7RrpqleSgo7K
dPeMRmmTRxIAg/Qg1umull6rBWIRtkhi6b0kPTJAauCiucljR+HcCV7P6QWyvDAaa2Y8ZaaW7t+8
qdMNvsIWFmcRYugpSnhbiupECx61BV9GSVV7dFUjgkUgSllz7pR2GPSLy8SGebUk3gWWJaFoGI4o
KNuEnlSsBTLPlKzYYv07n7jk73/vJoAw+7NWrshAY1NkrIA4jJax1ZVcl0bPnzr0nA1tuAxktVtv
kiJCVHsNbCkUnF1Ut0L9uFB1NBSDSxG9m/AkAMi1fwd/bT3YLqK3xqwfIexO0UhdbM4zPvQKcldx
0/P0FK3q9D3azcQm96Nmo8Ty/mSZDRfF1iCaEWTvrLQLV5dngU2ed9AebLrGecekH2tKBiSlm7CV
1e8DBrwUXNyWNp6H7AFsSCr/7873BckgtQaLxCt1r7rQgNDle6wAZaLEQUQtcudI7ei5xwc8zODI
VRE8eX6/QMmxPsw51IIKFy8du2Z6TTgSQ7DQSTWqOMVelGA8EIzEkcmOuDNKCYYoZBNOBMptkM2r
TJSsFKDKlPluSusoMy2LcN9ZPGIWEKAK043BrqPsUfQYy6HND2PiM+V3H3HZimMevyhhfsC2sOKV
98LqaDyxSUFGjEzxzqfwSafmyQG5xticQPd0WFOT4uZstqveXtAotXkBFBQ2m3IFVt10swDT3Tbc
wdSqohlRwX5ZCYnaiZwkg0+2xodnJyZnLzAYHBnYXC7AbwsyxEIhwjNQdycsAVloRaAtipscMHow
3TqOa010zXowwox6bLV++Xtdq/HnU+MKbHdbho+uVwJnYHQ0jXqb03O/9KE5QBVEg/cuTk2Y0D6+
ofMb7G0p/NYNr02XU6pqXLf7WPYYs0VbmexJYbBpmYeCRNc1jWYkZkhT0WRE8HCEe9/s9UWq+7Ca
ldgeYDgdY3e2TwTGNi5f+1+Te88XXZ5ME4unE0yHhaOpaJTP6TKOwaJAI745wIR0kMr3Y7HMLD9L
lAJeHko/TrtyfyhxoFwWZ6vDlYcP9m6lpVUyO2+wB+eucHEibfhdQlLaBOidH5MmQPAA1YQkFIzR
38992mmvo88ZBAofMYCLpLIXl3tbDs2Zs7moAl83iDaoeZTKLwyPal38HzdcOyePLtZwhthPkRGJ
BN8pyxVT0vYZ7aKxG1GOXuycui5nDkH2glKk8PzdUCWufT3u1n9isHhZrBEP5pDydsSBXfVLDA6n
U280PUoQdKwI++N0s8tvSx9/Bij3T20XwonI59veDvUJvxU4/SXiNc+t0MZ6eHTtoT3Eg4fVqrUt
q70Eq3P588Fh3Udl2qCP2+3I5X7+1mesb5qjdSaVSwNca+kSoERtfXr3nCZ+y8/V2VTFBfL2MCsB
Y8XbACsgT7hcaLGiuZcgrnOSUvWMNjFOZuh+fvW5rMYD+hDi08eFwV1DVov0xT+dfE4aplcbdQIB
yYeHBburp6NGa6R6mqhyPIMqhFmKGi88EVjhttwQefEvDjQI5F2970disGLImI6N6sKLGc6tmaFn
n5lx2CdNuMAd+Mv9SUkfqDkRAdNygTVCFqvK24/3pRbc896/8tg/DfPgE3GAykp4Lr1pxV4wrpEM
9wRtZFsznalCX2xr4b6sXk1YoR32gz5D4xOOymdiLRmJphoCF+LpJ7Gr8FRAvCc7uqCbZCEHiwG2
pWfXn3ElaUPZbhth3QJxWaEn+lYOdiDYwx7zIpD5XmG5ITMXQZm/qO6GHzP6hBct+KAGaZxZHooo
CUP13wvKQ7Z954AIlxAl5NCybGnfyJFZOb9Rtr4QrlZ6ZkcZ10v7DEOjQoX17vfLyK85kvrdvbbA
4l0uRTut6PMSUfCsTXvBMXlO+K8SelKDdSrpkExgY7qInrILDWokqRgrEqC4k2Fj9h5o9QeMFj2E
lCj7hvnSSiHvIaqo5F5a30BKS/k2ivrC7C1mlgVIBQm/ePobhMeMH/q9O3t9M0tOdf8AG6FFVOQp
Aolo8lPbqcqEXKGb4VQHTpMHAc6BQophjzfs1b9cotjoqrQukWTizdzTc95qY7lyuxjIcvustQ9D
TPgxn4pVjw/Hh2W2gFcFG7uf5hLuneea6ICzB+vLbfVRtrePm8TFiVVp2XvXmPFVXVw7ZJiYTj1g
eQJTaPd3t/dnnxN384uTolYCm9mozWKPkggOdhyoRWhqG0E8t3VURMtcL25MIiZt5ldrzklLjKKX
28xfKSz5IVJ4YHAdKJrI1ORbu5KQTwhcbbykhTjjmvILPfsW/JVLcL52ktKJTlvXG3a09QAPlw/F
AEmeMzorVo3qFhZ4XUUQ+lTruRjCsRz7/ztgdJF/YggzwaHAM3sO+Uxgn63/t/0xRECekn51akTK
yJ88Bnxtj8PbEI9xJxvj3obxGMxcw6E7aOVszqzaP+XDbKXwwmpMX7hf6hb1wsKNd4+Rtfx9keG5
8+A+i9sepyzX+7mtjn7CLcOs01jORfnojG7F/rqv49DzSmCiCcyklsSVCDZekNKGYRBsWjXYTqa6
/PYYviL8tTLVXjOBAjizX5JrfaOUlkhK8RNKnS8rzUO2DOyMgbEY0ZaMuMsKbOMb/OEAHe4ZRMfY
0ATzR/ZUdqj6fIB4EuvDdFgm5TdrNjZwx9yxzbTSNoRToWUuFJ8TkZ0d9FUX4OlLYW/NpETyl7Tr
4/2miYzh4j84lefAHAmzjJAlpvwQqwxHMWzzyWRgN3UCYmtzMOTbrsLlm+6uzJg2iP7bpcJ+S6+p
jk2IQKK3pvZMlpScEMjthJsMl+4SGiv1iMNu6UDmvq5FnT/VPahNY9dXhre1LpG0Ga9X8V5O3lnO
vMIF5Bf8gb+4ar4wi6CfTD0WBF3zp31DrmxUexXDcuOQ5TDMXsuGbGUHJYihgAdBSkD1ha2BldEc
5Ep781Lvaw8xPeeu/LwXNZM6dQLKGG3bdn46XbFshBZMXWGeTEvqiVpBHx2/GapNOCeNI5LZ3ols
rUVes/fbQ1fzyHZ4aeMTeTGhRBhUyTArnoDVlM7PZR2cmGMtejq27ZoqGG37wTOfCPGyFb0Xvjj6
s/0Mw/mEN8ReByS4D45XJ5lB1OQNiwLg08mI/QCFWfdUicUrYJZOZ4vja1sapMSzYZVQ/Y07AHBX
F28KhTZ2e3udPJ4pEY7DMjHleRGH4rd1IPT/6hZ07LoF4ckiktNzoUAAfF+cWJRKYd89Ui9U4Au1
OPw906j49+0iefcHR2t7EY2oF3ECHwgHGDia3mvFsE6Jinda5OlrM87eXGQw4TNK4vtVm9461fJu
uVlKpNSULZd6J8JwIWHpiEwcDoJLQRQMuk2y1shceu5UzUM7NpVpoZm29CHMpe7AE5CwN1oEsI1Y
1JZ99oi+W/fCjChBy3G6y5XDdQl0QPmQAbsc+IpjiOtfFaieyM9w/znotklWFNmJtQL2TJS5ISqa
EogN0YAfUBkUEIJqD7kcIVuaLBwN0u1f97KA+z55WImiUeqvsnD3u+Ceq7cC5CnsLTChBzFT4qm+
Ha/mCn2RTWYqGIj6YLJJNSxcqe6+OrJPyHWo3EniQi6A/ad6mj9Clb/HCdkKOx8YVhrnp5WNudje
MLxTWI3SMWifSj2xwu3/rbv+NDRXjLAjfJ+EZeaXFtN8X57I6xO9q8ZEoo2Oe5A5lr0V9pkDacSg
2c75K6clfxIW75TpreAF4ax5c00ZQN7Fc6Up9B/SqY8nLeV70jziEFECRh67YHrluaqAlXKdisBd
ThCewdF2Ns74r976156unX5x5k8gLKC6WzP5Rfwcwq0+Dbm5VC/v6/JT3zgEb6szl43qCwFIgLoE
aQp4Ar2vyZM3XUF76V20t+4LkAH5w0BNYNISQF2WTHi75TSaiz/PRIckD2M8fjiVm9AKdNFVP9AY
aqDOWYJIkqU4mO8ss7OemwgVAwgXzgYYBy/zpbGaksaaTteVs/KPVvkCKJdnhgT5/flpPcme8dsv
eQYwZgjjP6vWow7mNNqrBsE2L/WfUnbD9r0xnFmLi1ej7V/1Yd4IXtI/kBdCmwKWkC7WZn5YSj8A
C1c0M7oE1apKNufVVLUyg7tBw2Abtz02wL2CmxKE8XB0H7ugWMVXdQJ7a2hHfiChSpReGb1idSjM
o8HmQpXOdIbhGGZIfcoOvziYBU505ZkKWR3c3/PvHQhE8O3Z+jwDTQUenv5UVM0WkcVUGfnhsYub
EwjaDtnXQGe/+wXQJJR1B2EfTwX4UdTrLCfKTe+6lHLI5dfee4IjETaCIoV9oxaX0gQWIPi/L0pJ
fjrFp0+YU+8bh4UWi16Ly+gfvI+Mm8SmyppzJPjQynyFQdWguHcwoBLc5Hkfvyz4Gs0nsKtgNAHS
jbuOI8yzOyXeYrdDNJgOE6NxEo+SG8aJqC8/uzZyfT3pNWwxbni5zz327v5j+Py9xdqp8Rfafyfw
Q/KHCyvXy/rwZyqepnL+T8EseJ6TQFJkQn0j7E7/fybUHI6YCawjIsgsKwbyk7pY3qE8ZcnysTqi
Oig1fZnFefn4b5nVr+UgPyt9xJ8mJssIfrRkCxK52rL+P1cG2nJ2qHWGpq5yRYXT0qwNEcVL6arP
TQujdlzphEloYhpLy8zYkdJt0f9x9xrkTvy97bVnlLVP0ROUcwmmukExYnrCuju0Ar7UdmzLjwG9
I061fAbg5oJXWZQBzzsSRwUg9Wv1JkFUeO8XXAAISkRWu9QndmiQUstofNXOdWAzTT220+7JKJs+
0m9vowgwJKS5VcwduInu8GjfJrw621LlrbuVnwiwuf0Tm4Dgsqg8XhljzPPv1IUcugc3gREFvEg6
gEXZXuwQ3yOuz4Kk7KHbxQVC+fsXy9tslSBhZsHLNWTKwGPG+nuBsXHlOrE9XoO6K0hTnHSWeYT7
1SfVz73/DrLHY9UYWVj1NHdw862p2F6Ehc7hSKUQkzVJJfeGUbj41Vojd8E9UTzw8ElOUo4gFuG4
/KiixVGST+E3a8kgR3kOkVeW/kPxMbzhZIXHAZw9993KUYfbmZmWAAFljXuHyXUEvS/DAS3ekXWQ
YZxrcm+ETRFNkbL/E8Hxv3N/7a7whSj6JO7VUR8l6Ku7x6awM5/A39yDmHrJ9gcTsY3D7tX5OXV6
JUSesrGXe9M2CxgCEcCCqcDnp9pHLVoU4BEptd5ENE3Bf0q9S8tS4TZpiLJSge9h4yffnPbiCa0u
/t0RP5K09gwaQlEFaL/mlmftrLElgqDZEzFPXN6stPeIdQL6+siyVxV7Qa8S3l1ad5yrBlKqlPmw
PBNrY2k8lm1IiebfSOZdTMnNvnIPl1dn6ec7CC3r/rGV54ploDX8dYhFi/mIKbiv5Weo5z49TsHQ
qEKCAfaVChBoiVlQrWmVk7vi9r1HpjCjZbehrIzsBQ1FZPEsHMXd5I2W4Pq4tqyXskDiIOGz5G0L
6Q9Fxv2kPadqVfFO6a3cvLWik8eLxRWFPEGD9Qc8zZakW2MWtr9SajAXC/V8ZDIMaBHj6F1Do7nd
wByJU0twGQPx9W3gKsCAtPrAxddqEM8ZQZ3ggZqjT062I4ilt8K+MuSEZT+f1I5YQBwt4k2jQQpx
mgxEoN4dfRii3ptPge7BNfgzWqgc8VHgPXOMt/YY6gpkBrDxcdJaGIuXwh7krKbCUlsBwaNqSIj1
o0dEeaZm3EAd8n0UaCHmk1KQ8+M91NS812jiCQDVq21E9JW1V3AJjiiZVoXZS4X0VLN7jXyuCNVQ
EkWBE5PJjQT1TTflJovJAH2Db0SN/d/9A7tAJpmjZ12mMTJzBmd+68nw9KXoGc85jYg1PdXidpcm
AmxPpnBeHzfe9fjcc0eyUTUbnfiOH3tSRrTUPJjopXS9HnP7AiFYFSae+NjFVl1kaJQUFZOkOKVj
Hn1UJlg9WGFC7sYH4cjIV8Ofnu1DOUxagFoU9hc+7MMaCdOFkn6EVRIjj2LepjtESPlEprijTyWg
z2Mp3brSSeNJWQjzd3nlCV0xzrfNFM6MVDXRQEkaW46W+jqNSud9Tg6KuZxlP2SKJzc61zSMCUvp
0/yMTjtlQrXZ0QOhyxNBbkfmVmdJ77jbj/KG6l8FrSecAagHLKqoEzCs9jYDCNgdAcpCA6E6qo0A
hvzMe5ahiqxhW4j1ChsJyL1eNNYuZW4Q6Udijoaj02F6RnDzlBEwdgc8vfYGAcZL0yYB4d566kME
Nv5ASzMecvIOky79suYTnyrgKnuDBaHuRVzY9TpFfZ3PsXhFm6qmaJth/fsagjfvlumBrHVdqM/g
14uUqUCGxUeAw3kL36zXmRCSfB/AMLjz2tn7Ye4LXAdzrA3ndO2mN+XLZ7auRQ//P5dAY3Ca1vso
t5eaPrw9Gs5tBWE6nHYBj3ux4TJQPeY5sL7vLbmCpirgbJofFPR16Iawi6rIeKsaEUtoDTll3yeG
ItrIBc0HTWA437VLI8+4VeT1bfur+QH2/D1awkvgosPs8OBO3kf3HzmATNB35OMBC3FRPajDS5zo
slNALb4AWXTv+XdHCGLVQaVeP75ndLIZc16rDPYAXpWNJe+8AWWIU/Mt/74YsSiT/DEpjjsTLk1S
PWSKQrq08I4V/QRHNu+5GbsZrOVxno4DAoik2iVirx2zicPjb2Gt1+G8VwgKN27HZrYIC7TtYTj0
Qv9M1CP3p0yIfsbMMmt7PbOA87IIGb1t3hgVbYLLd4uIfPPI1MX5o/FAzV3eitBbcpq+25fZuGq9
IYFA+zT8P4k0r2BFlwdLDB40Qm2Huczkxoe2wX6Hlj6LB/Afso/j3MBp4yzNpkBSXGQSK32ZJsYS
68Eou6EhN7FcQXCqS70wXnHWKOWMJTfGdXFM3c/D4Kv0T8q7PImxcyB8oOAMifZZe3C7oNwjeLdf
ddRutS9QCn6ARmW+IJfA0M8xjB83gbX/yHqDrruvXI34Pnrj+P+JZhG0nzrREqPCGcuZKJIViqzu
kqu+XhMW64LmeVfQJ0oBNbVXjaLka6vPXEnPIbVn0ynzm5F+ruFUq6PQYpkwGIK8yztN71pr56Ed
aXQ5TIseLqaPbWO1MECGd1Tyc11CcK5QP9+foXtdh2i52+nTNObZ58C7ub0k/mXd2mJ1OVKVm6Gq
ubyKcpalFk9N7nMQ/Boym9ax5TOV6tIfs+VyrD2euVuQ499i/pccZTI+BpvXsRJxgneRTvzfreu1
bBCWToIl5prehu1XDvQmPlzv5mF7r8rTF0LxgFQnJYyy/BTPdA+90EQrY+6A87qZMAYc0hDw6w+1
JkEN6M6tmJ8roFnOvpqgIv8RdGbvWlRyDqnh3iM/gFeUg4OSyh7HkdA0vcDqLQwcWCHElBw4kB9v
HpnidnY05MjfmSePi7UPffAHEkG487HxauwzuOQIC1nytXFZG+N0DaoNsgqpSpzW9EtVm/tiuJQT
l5L9ky2SDkZHQ5xPgdrsk2li2vooAL+mg7lUtQZjOltAZWJdV0oX4PLo+LokqCTdNcwILs1QF9Q+
vYP3S4UlB8pRDY6LtVrjIP0ZZjyUhk9L6VeTPSFHlYEKePLMTz+MNIoqoaPaLIcMJi6l9UOpRoRM
HDBJS1geuOFff+P/TVEWNZLWKOXqfcmaH5Y7afwVRN5c1hNos3p2YEVoYzdsONqT3sFnzEc88Hyo
0/YuCpn4YXjlcqI8qf+bNLwCMeZDtrLvj5cXRdCyxzzBomgTG61EsmXggF5h6g5vt7gUag3T32iV
xp3pLANNM4s+Qa4SqjZUPe1JbhUaQK9tr7+6If8Ns+FrC2HpG1eUAXydlj47xDW7ceojgEtWV26J
cQlXrEpR70tleYfPEiBei1S2R5a0u1x68bCtCgP0vVtBN3AgpvWnixdmJhU4S+rqHouGSd3UzVtC
Bn6yaGUCI7PWQdLYs1EPux8lwG1JBKqv1w9h+T/ykeRyYTMKeFi7G3wxantEzSQGYxNNtaQ13xr3
uNjKLv8KUDtS776VZrNPYGtlVrA9gzgJ3b5dsNw8s8cma1fwW4bRfmV3cASHUVCIbvEcMgPbtnfv
OEflNQI4zPNyxxGHki8ZxocYkeE20zzVZusSjxaRcA/5yIFxm9ipJhHv+FFVNgFJ1g2Cl7p3j63k
n5U2alr2oFKP3Np9QEbQgeYXnH5Xbk53tSX21qkupJySn+iQGSNR7bw8D2iV5FrjEVJ/u84sv1eS
VznZPdGMporBDPoJDMkFh67v0nM+UpgKbOP1j2LDMhlEETcoBJxA5Ep27KauFTfYD0Tg6jHbV8fi
ysSGTGxolNMcGmWhyvmAkssaYMkOzYuF2uHa6k35Lih5vBkxUiyfknNSaHXFYKplkYRJLSyVaPhq
UMyaMZq7QLkIQOnHFCp0VWyuGS4BzFKpcicOFrkI6YmwfFfIgemvJMJUl6T0LlW6hEzJkaQKk3Sx
fLq4T8ym68MpA/TRdVubKRdst1i9BicXzZg0H6lY27QQ/QCOeL34du/pJsn/9I03HzkIEyqxpdvf
yCnHkczTmrA2BSZRuE85fiSYWYKxUg2NkrYqgAU8TQwRDY++BoPONn7WtDsoQhfeFUfKtrQ7cGqk
LbkINsZZ7MQx55U8nxA2xHwpqSY/bcyd9JtJV5x4ak25cf+YJ4G7bg0wm+mPsF/ANDjYkZ2YT7id
f7y+WbrA7FWgUcKfBnjbPB/WsGi96GoNmsCwtuFbgJwgb8USRpYOUUQp6ZfQ5Sq/pvNqaxWtBA3R
b8rxPEtYmkKaG0lWCyN4AzuuOAHvBkzFAIpfpIUgZrQQcs80iQKAkNMgOXVpoxKoB67eC76MJIB5
80VKJ5M9Kr94BqMNxu2Fer5kiPLb006J5JKxU7m3rzGWNCfeLBPF1h1DbWqYJQiCXlFbU4VO6IVD
2DjXANYqMTHZtUBBRoWI4cwMNxSvBmIuERui946Gf3NG+cfeLd53kn+jKMhoLgSMe6bmmdp7Id8Z
IXqchUr62XKIWyM8PJq2RkanXntiX6WKobFCp/2vDsutLgs/QD1Ckc3zTp2s+M+sViC6A32dkmhh
sUr9zpHgvtBFll0b3xeHscx8bL4vglRXm3GOZ34TAswEb8hhHlPxUuh2jDQpN+VFViyAa992v9S0
njKyvQsNy0Lf3ksyPIx9hZirfx2ffvPtL3BQg+kHqcyNXeFsVq2oAwXBymX4crmAog+PWrDLtU1V
GzPKplxMck7jeoOVkFckbocFYVUKi8GWpi//Fh/XSxJZcqO1yCg+/tIxNaIHJitu0xMj/Sf60Pl+
sT6rQuYcKAqXhx4PrnZzUChFA/lmkxL9UtZSn+2iL00WGLoScc4jkOdnwfecurpVfeHWJZn5tTKe
WmGIODbEDtjd76qc4Qje6fh4C8bGBmEz4Evkrq/votYUDt/I+Ga8AztG5nO0QBqn9Q1V7QPoh71E
VwJuna4PxYHY0Awpcu7WyszX83TQxauG6my1aWO3vtK4CLnx5xthRxm+5bZV/Fpn3DitQkWDFRTE
Mx4S5MCIy1Cpu3X7Td2VvpIM5tglMw4i2V44bcCN+2GsYrRHtS7eGz8ULjBxNW6LTxw+ubpImXWQ
9shyreteDNFEvgU+XIBs8sfKvh61conAiajHwzgaYOVnV7/xZYzwLzvQwZUAU/uogSX+FdA6SPMg
rnr60tEdAo/tHpCqPkC3woMjjSdTrcDRI6HBFw0Z0Y0SZOY6SYuVkhh7wdpNlb5cyFYsfcSyHsvp
q+9+ls4WVTa3LEOpCmX1DPWmC5WFHCtEYn+qPTo26AzCtOIpAE8w0jwTjXFC/Q++kj16GcIvW4TL
qtwC+H1ufw3+qrhaxFFOXamwZ3YKu3fp/glOTghe3Nt94g5Lt35oR/pyhZb5//aR9eyWXfQwTx7N
5slo3THSex4EhL+vTsExa8h2DlTBdhrQQ2/aJNsG1FbIRN64SdQQ5suUDBRBSbQ8Kpa7c0/BzxPj
rbqManllRODSMody3bbN1D+KY6ypF3+G6GLk81+Qbg/CjOltkekFbMHxPRBtTHD8L5zI0OF7W4BT
SX47SIMZlMD/0EQG637P9GnjfnTp5myGrIzRVK7ALb1NB2jQVOIMbHCQc8R1by1Uo6ZdfAuCkrmt
Jr+UEvEPYWisclPjzVKegtsSavfj+Y38OrxJIF8pyTKHnYyH/9YrnJYHfUZqCgPvIGqLy9he7mHz
Co52M+T82rX/slK7TTH/J3YVYvd13GRri2Y0rw2hDSGNBTO7iA+mKOR2Im+9LV0qm2v76RTGXVhI
l6l9OfXC5vR8A9bkVREzkDJFHFkLPAsqglKyvObyZ5x87bvIA8B0YzqL+ZkwOx3RnNZRgOamhsEk
EuX3Ywp1pAeB15PL1zxLL+cybiQAHloSPTUYO2bJDSxdlfDIIWzi0N4ce9K0Z+x4DhhuIc5ZRY0H
wXfKBiIqcecXHj2wMcyikABOL+ostRWaxxX9494ZcdD2anKPx2BdQl7TtYlQE059nP9f3aRkS+KY
8O1O2lCrcFdpy0OVwivOGMz/I3mhwpSzgoSM0skkk27MPJlZfCy1Psb50LvM5zU3Ozde93k1Gz7H
irGlc56MCVMN1Ul0JkZ4F3X5DLxoibpUENXupGQeclc3D8tG2dqhLvaqLXeNzGSYaUt8dsH3Fqx4
VgwD4BZ1pAP1fXknfjwb+wOzzT/ijCw+5yc+Za1S3sgOHrZmTqrVC7S09HB1I78jBYK+8nO4g6I0
lf2aVjXMQuuj0+r+6LUauJNiabsuaPkXt8Ann8cs6FL+1IEM/5LMWGPSbKI5Zm09SQ9QkG3lZcYg
iKikheA9Dwj6XzNT/OLNJNfSINVLt7DZjsz8WblsEHt4iiSyBvKsffFbtLjnrha+3e4x8I4N8Y1D
bI0geQF8SgY2HIuP3a5PcBhCtxylkl0/8yEtyBCoehIQR/kXuZVzTtjrs/8XnjO8nsQNnscz66bz
jpjs1l3TF6L/hjkx7dNKG5KwFUIeCbbIz6IoAee/fQDn+yOuhtTWSapU9TEltLUfBMU7DOd7t0EG
eFM1brSuRax0LocKhJ1JNi1BSb9p/kGFp/owHdHJHw4LMrWmcZ2tWucmGyBo+UmSuqRX7o/dToml
MguBLc2WfGLVHT7ZqCJJQwUoi3U9/rJIJFK+c/hQh8J70mLgWdagmrwyMBTio7zHZkco5oXliZ8j
lHzrpOQ4UDD7tJUPs+KuhpWS8YD7uLiADTJmOCmWzjUuLmft/bI7slhJQKY3nroQ453FmqpiV4XV
UqwYed/1A57pf8LpeipqK+L9jHV9HEzSl3tutYMSU+sZFRfSEegMVuYpNYREpzRVCfXyR5Dlo3sH
/fXQsqfEiq3zBj03NHWC3ZpWnB9SZYoH4Z2mA1uNHzHEQXpCkg9McFW0Uw5SD8x3r9xCmy/oCbpr
vMUy9kiDv/rn/9XlMDCU4MftH5vWqYSOuotGO5f5k50oNm9YHhQBIXTb/oJ4gTUKx1kZQvIoM1kG
0WDvir8q4fnSAhHWLXL3+zqCzk7dcfJay0f6wYcLqvjFUd0Dzr3bU4hqMLfXO9hdPUxfHF4nzwBj
cJApRiZakwnLXlm1q/qdKeGTdApBV48c7Bwoa8nP/3mKVGLs9OHnvOJ4M1klzVP5S6WDFdcsBzqB
fThO9jgvGqHr5uFdOiF8hP6gLLA9SQ1ErtlMC9H3wv8PaTfaRB3WA86U+eGlVD1piT2xsLozpNoN
Chc+n79hyomqxpc/JUdxERxh7Ru6imjiqBFakAW3wDjchkFH0DKytXeSY/miaHxhtSXPN2zWLXJb
lqsiICyKgZ7qefgHIinvnPGzWYpFroqZQvzcWF3Db8lh6evnr3k4QtjhZU6Zfng2nV4DEvbGrrJw
YX0JdW0JAlezTV4EZS7z/nlsuZ9xyECZVrEXVR081FNQyx2FhZ80sD9Orsfvf7kYGVgOBAA1ARRy
U579WixOvQflHOuj5svtKLqXKGmG4z82UjMdehZmJobIv9dSv6MPfi9LHCLM7GOXFRXDQhuVIpEc
FLUAH5QHek4DJnr3n0j0RJ7i830LyAT0RayTjz3EF4z0fxe9cMu4lf5Zs9ZNFu6jaHk8Exc/yiAY
Myrwpu3IeClSkXZwxykhOWms6UnecyCYdoNbBFTttPe9TXHPK1GIlH8+vB3sKTP0eVO7ixqOtKyr
ZNhvZXXZSuM0BScggo89jmMqgE7FQCkYhWPB21TzhuEmx62/ydz4QjeZ4f1L0UYlW6GLrvenJc6C
rwLlxZ4yUf2VhwbIwZ8Fa28gxV7j+ioTuex3UjzYhEdI2zs658153CuX/kKRBEoCvYxYQv4F4KXn
RbZhvA9jDVXkXRacmRCJFumm8V6y2bRIDUFrAkMHBoW2Gm5fRAGMpn1NY7i4EY4cXN8aJTGcpufi
NIGDYEQBxzxrUFIu2SPUQDrQ7z0vIHBnhbMNeEI9CVYpKnB0079sPgLgKBBeI7aCHNKgmKgZvcWj
PH1rMU475oackpLHAU0fppy7FYx6fXQA3wsKgbDS/Nx8mc92fArPAsBX3Br7xMKME4YbuzshD5xy
d570nN+ZbqSZNIYWKCFruV+R/Unof0uX1ONqfaeyIrtA7MO+m75NXmlGJG3nYWlOrnq0QqwfFe9t
r5XWJLU+BLMA5SkbSNAHqGHcOMrrCPzwMHhoAzB33zMJW/LT6cQv23hIHYgdppgndBuHDnn+1OE4
d9HTJNpwyiZ3IRqYx196R+u7TTR6MO8EUfBAPP6DpnSyY8LM9lX+pmqDcRAf0UuXwPSZmfkLA6Ld
u7UaHoexXEKPgGXj2sGRGyodRpWfBOBlRnDMDLeRJ8cVtaE9h7PMlLoTFjAU6HVouwTfIyvS4KlK
UUN0MmH1zwvjodPPhg+3TtXs/qYVnXJYoMevXjIjoLZatecAx4jvqMR82pXPnPvro4tWCLj7ahCu
TGscXZYHbqGhpq3V4F9PbF3ID07kTqcUAB3KTMI7waY8t/Z2G8xVuYtbSB1j7JlXXoeEn2rbZHBM
JCIA+3z52ZEYdhnN8VzFce1Q0sYtKgFjd3fQLN66ASuZFJJysJNOYfiMIzjBKpxol0yjC2agxMFF
NxylZFJ2b+p55S5FvKT2DcD1s8hhLspxIZjIpxRxGbsS9qRq1bx6vZD/js68WJm2r4XbcchWqr0w
JmRaSzyIIZBmlsdCU/RZRdDd91BMkxAmrb0Od6c1C9C0npQmXCZfaFChTLptzospn2CFj4jPwQJ4
X49ZHwEtlD+UCyj73Rc19+dWQAZvl19iuwtZI33LQU7WP8Lny+4IAnXMS7uI2ueQKAOKTcOWOF/X
X5BAO05Eu1sBViHUrJ9G1hbQ5yPKEE+j+VSkc5PotbIPMblSXkUuLWONNrshlv/lsUSEYeQMUwHG
oyq9+XjQG4tnu08Gx9EpgN9oNDvwPS2ZpFV1uP78PMSFz3W2Pgh+Dhf2mDvNvZn96IbD7wXe0G29
L4XIOkG32Iav/w+U31viL1P1p0myjhwdplTky4/JXY9F7od7aV/PgCnQfoyqotdIc06khfmAm7/4
q7eeRqV50QF/k5VhfaoT1u/I1VB+tzO/Oq6WrCLDk2wwgxq63yVMPDZfTdhITzGgl4Xg1TbSls11
ebOahJcYeocH4oDapqyLfgk+h2bRHGcBlVMx0emank6s2n+ifmuEShVN69L6WnG3SyZTGsZkXInP
sfK72D3mjamGHLdiobJRbtkcDFgk/IUiGgZEnN1tLVcTNkWY1DEZ9UGjBNNvmkZDn8I8WiLYMiKD
9sxLZWGP4ug35GDDQ4xZo/CtLFutw5TjRg81fD/r5vaP1yX149srslPjrIbF5D9jAivGPhUhL/9e
ldeyXtYGYxgSf6ghM7Z//7PpYKWen+S4PlDgeZP+/EAbLiQWo2CfIHYG+72sQOasc4Q46Y9QJNyt
He3uEyX9/T5S26cXkyhQtTznjuLq4/bqKpyrkRO3aJ4erNwTDq8PU5EYBytaSNtZic3/3LcGaZqA
onzSijz7pqc+cgEQ8DKqKKVNDMO5fnLwGBbdatlpwREWjm4fjfZ16fLNwJ9G/ebASsfebPX3Kl9c
7C4rd6B2np5unCL7rBQD50ggKC2W4TZjnboQcgLnx8ZEsefTj3jLd7ffG+g8cYbRlQIaGIvJ2Gdp
vSR2SikrFfaRtzjzxcrs+WcNjDrSg+p0Z02ESyNXGeB2OffTtxi5UJiqstXdtSTHqTxjRZfe5ZZr
6wnJgg5pknmstNNgGPbNDOWDMeZ2dRwnAjHHXzyZ6r8pGdjUajihSFsLSuvmpLBI1mZzPKcpNnES
th7R9bCMyYlD4dlS9/1C3W2a4NAu+mWM6F3lFzF60XFAx6eoE2yFw17Xn1tLSuBZCL5ZWuUkxvlV
X7IXSqKaJNS8QTI9riPnSpLCq9Oa/oaTQdIBJm+FaAPRwYFh9zRW6S8YKmjfe3VWRzkdzaUMooiB
zIQslMZqNZeyYHLmGUzadetQWioD/gVkMU932hYEHhGhH3yqu41RWfcDeHkpXMspbrkI/Rf/EJH7
xBEO6YQnm41U/vlVk+KQcOyPlUVKaG0tVaGJUJccQko8m1s6j0ARAM0dJAgqChR21uldfn3uuHFT
AdLvPZsOoV6zct8/BvYzvwCTmLPdyJOM0GQ/4hJ4erKu35j7ZWV6VAUEDoTceKIX65/3c4qAyRjN
QFUXAXBEoj563t6S5AYDRughX/il4SZJjywzuH+4+P9/xQjzErnAgxGhOzFeXLZmN/H5VYbuswYF
awOFeTUNAj4pOY5XfDERTJSgp0ksTSl3rEii2xlUyKnyVCPKby6STkkJbRi8OUJ3gXEUNZo/r4HT
yDVvT5n/F8cmVBemracRrIW8iEJ4bTXxTMcqpem77UBNShk3zzYQWYBXdq+97DbMaq3GrvbRLJHG
r5SQXO1AXoYM58IO7yUrZeY4jOioZuGPPSTxtkE6O5z6tviAiVE8+l+TU4TqgTjPxhOKMwacB107
JPZaRnH5i7AuAw1RdtBgk+Z/kdwzbFj9fE/mBIsz1Qh+qiMOPryQZLunFEYBjne/tpfgXIWi2IUG
RFsZB5gDx5z0Kqaw0ZCV8li6w7HzKlusc0/4WfK4GTKjy8oFncsxCJG2nNyQZNlL1/xiHW5QUF1E
zxQFImj9qwPPOZBV1CPSzZMvgu+Jd9gAu6VE3/ky0GkP/DaehqHrFN+RJksY8YqJ+nEY/5EzdvPU
QAOzYendc+wpMFwiu0n1etQ5GhkQnW1F4ksc0oDi2f56d9pGGbkn6XBadZ0mk4+9ME2Xw/B43EGM
eFPCnzON5eXRjL+rNcVaLt1vDzdVPpdes9yFEUOWe12J9BK5TNPGB4xAudLDAnoOPbBCZ2j43mlQ
KVoe4YMV0pFQgvG6veJ6gWq/3mNgb5k3rVu3LmDw/C+EXndNgpalY0WgfaghUDYsjepQVCzCwBUG
d+3loXZvGYU30PqX/IlqrSE8jCY6xH1ewX4VLqDyCK9KN29oyqfJe/okJQ8nW3opaFOnAZtjkAIQ
ajvWGoJaz6buEOVMogTm1+xElVXzFHAuWaASch9oy7rnBlqiM3Md3/vD+yd1RAwj8yZdVTaTpski
YjjNLxzc5Tt7aEqlsp8+t6QUHKTquXy1Q+xpBiN5HWeVx9lAW7M/1cWuMtLRl4ipqYpUrN39VQYF
t5dseGoqV5EjrvibqFQchhmCWh7MdxnVErWQYk3sfwHtQqmOR1FkogV3qqms85SMCEx5huJHZH3g
jrvU57Td8BY8BqRqtrlJSO62NzKqeqNBGtaXU5Z1YWm1YYEXIsCk5OZRb5fdL2ZUQLtVCtSlTM3D
R+EqEq66cD9dwk/rwqqWsD0GhD0gadBelzaJVT8lPVTCUE6guzfcj3/q0yu8d09syW7MotA6fgK2
ra3gJ2VbjCNAO3EVP4Khtc5ydVD1DpNQcd5sxWxSoXC0+KSR7M2oS+Z94xOC8lP0/MaHrBg/Ljd8
lGZLTMSNZgEYHho/2sbhjcZa582z95QnE5JRkc0+F+gkSS2p0T34VVLQmRauSKa2CCx7WR9Kuxk9
ltQjoFJh0/3/gVwWUNb3VbLXxnPvX587UuttFcj9ZAycVzcoF3XOPGz7FQ9/w4Z+kSnilZqO8KKW
JgNjABUIMBYcWxETGhLtJo+2pYFftmfzwklltEOwddZLlpyukANg9yhg19eKvWV8J/iaO3Mt1ywl
AVtJU8sxlFyEB6kMrMQSCV0rz1tS6/mVzyRMS5jPXADGXlvlykKqV3kLYWRqUcG4JkOJo97KsgSG
ukHYRS+58U43wdUtoofaWdOFisVtFvn9JcO8I/kjzvKm4aJ4lystcVm6KN6yrsbkTtCAaOsKnz9u
EtEeaafRTuAkcnmVa9eg6Fjgb+OhfmsGz8G/SnXrsq25M7UPSIWdiXqzCtG1MwzU5xcV3pn+oewd
ytfP56hgXrXFs+mu6yb+FwggbaY72ZkJMCOswqkVqF6ce9znIq/NkPGPwmI9dFZpLQb7ZDOrXLm3
Jt4AqFFRAWr/vNO8KyDBsoFhZeYob8LOnF0HYkmLIBH3E6SjYb8qKWcKNBDPlQu9IN2KuE6EV0tz
pIzBV0aryE3T/1Mh6LPblW7b+B9M45nhw+0irW1WLPdbrcfM/Og8vM/XZImxc3RhH1r9S2m7wHHz
kHL23DCY5Ra/7bRLwa/TI2mtMIdzeOdQoYHyPQ2X2BHp+HGDmJKm0uGfiBB8QXUMvJO/RlvNCLOz
S5Cu5M1mcz/3wlZlnhpZ9BiIHyGSMFLBxtdDKI+EOrSLJBmHF2OKBmH/H5op22VVuzF+tjqoYWux
7lmOZ2dtGNh0Enm+FPRcErCNUCkk54e3iR0FtApq6u1+t4yXhQ5O4bJuD/FaDqWWlG0u1SkAJ5Zb
tzMPYN10q8aj871pFKod5nmMX9RvZxAgnJ3ov+XNw3hTah1LdfxcxxO6I1dZnqhofnMeLN46XJNB
UOvgaaywNhCZ8CnmY3t8JmAZCMIr2mOJV6oXYtxb5GwL9noM8TKtUaUjlg4pCs8s4Z1cvQgUKAMW
9eXl3aO1peu18jqz8DHPQuCcvS6xeMjUVKIofxETDIB6w7jgWHicYikVgWGk4JOWH64EDj47vvkj
r7b04xkwWItNKv7nxMLTZaVNvLGhCEmG1Gc/KXDJaUODlExz0V9ox436sSSofNQzK5g1S86Jnqa9
gFgFjRjlodVvl9wRUg4PHsN/Ak58bh01eyV4wBMDDN2xfx/AdUUSjuTPdqP40CdZo89p6xdVD5rp
yBu8CqatymT/6FwHm9kZGaGyJ324hKuq21A4cYOQwl075VKKl6+zAWv1AYmzOgfvbRTLGO/RdnNF
UJjKUkbc3rTjd3Qcq84huBEcHWSkUSsueTZLw2dmovxaGd3VhqwD6Z3VqWEChI7nCeIEKcyUe3LJ
SqbxLge1mANGI1YOD9K86+TtWS33XwXJTdZ6gFSsTzfafzm4taPlxOpO9R9kh/3DtkJLEMRK3/mR
pduLHM/cNo2M9LQSU3WsHJq3o/aI3Pa6/aihgktAf3aXEasqzMBl9E2TvjgVgfZs2CZAHX55Rwfd
RoOoe0RbYb+4m3dvFE718Q/NTDghAM0o/su0t3zjLDXodlT/twIZn5CXVfOHrDEWizdvATIxxbuE
y80CbF2tBfIv/so/TLJus+r5EYjgjxnc6KBPOhME0h7ud0iTdNLOD9piboJ0p5XKSG5hok63VExP
qbsrcuCRH3vSCweCteFY4d1R/IIv58txiyO3eemwrX/fDuPIylKX48PjX0rVgLcnytgbCj0QiNqt
zTMPM9hY8/rSuKb5BEDu/i6CemsFAn7gSsXZ2MjRWGc+0CiwIMV3LjOpoeizEU+UJUTRdUnvnhWf
XCkundcgHjTkcepZr8p6Hfux35Z40JABArrzM0JLuTLtuHb1amN2tv1KbsaaMK/J7V26Cp8IfSZI
OGrCj2mMwCwNC444ptGRcT8CbDZmpqCJz85COmFNn7QD0A59pwdZ0j2l6WniMljlqWaOyKdA6skj
X75IAxK1GPX6y/OJq1Ch/WXEWIgb5tc+Dap7DPlNDMG2VT5ywDGAy4M84pGvjRBqKYs1a+PY8rrZ
8QFR8ynDXkh6ijBeBfBQJRdYgyjTBujaR4N23AewZEqtY6s9uQZtP50uj41qoFwrMZNrMTP4Qnax
JcjzIQiXDGqXvHvwmnSnpStpPK7P10ypxLnq1fEaixangq31MFCJ8DsP2hNqbP77CWuilFTJGAJR
/EYT0OrV/iNRkbNmMUa7MqyX4EjqUCiXb1arOScwud+lce1bNeyldlOUX9Gf/lExE+9qfFqVZYhl
sTuQXx4WnVz6KP487sS0gEsY9eqzNNfaevCgg9G06Uq+SWtoCRvXp3nswvX0fm1Rzfg4oL+TdLlk
SJTDffF2GVgZKOQT4H04xpbcFEgxniTV0VJHkE2NuiZ+eKMt/EXgoiNyrtDcoULjpXXPHBWoP+TX
A7Eubn+M96E+tgqJoGdswH+5edgMx4/sgnZnetiov31vuufRn1T9RuNW8X41gH5ikNy3Q9/lkayW
BXBaqORJFi+IPvbLdgiepYAk5HpYpMRip14H1E1HY5KkbM+8X5BekGC1CQT6vJ5Ah0Cknedg90kX
Cnv7KgCfSU7ErN9MxYSRlCjVo16WKrs9KAQah8hdj3rOiDmjK1VfkxgZ5g4ebtfKGsztp9JtdITM
dCvSDpAvdov0dF0p4dwmgeAeukOovi7on+f3s81YZ9IhWPEAVleGLF46YjWPRXD28UeMaoTATYw9
K1n274e2xeeN/2Y595SNRK+yZ4GKHgZAwPweLtgAanJTMigkqVlt1rRtp5EYMPwVTD+bSDQCRLFu
jrjV4z/AZj9axBknoYDwO4Max/ZMYY6lF6mhj+GRfja4e5LP+xZ0Go0y5Weu5eZxptV4qHKa9e9F
7Lh870hfSUnhgiKW5cuCEvxCC2nLXDsllL/Fyuri1wdktwOBHYujwCZdpu/aHlXGjoRaEFkOUoDJ
i83cgdm+pPd+2UAhgYBAh6699FVCzr5GcJWhq0V837fCb3EEKo90Frs0SUhjsRkyQWyTo9SfEqAn
IkmIbQAIn5Y6zg6cZCo4L2UQlgiQbxCQIsjI/POFzsWF+kCloNADUeJk8PjtJxz+FQ8fHG4ZKvBM
hXa4jlBkJJ5gIWjWeq0bIUtCG/8IrbH+R6blkd5i8B04yn85efQ+Ks8iGglpWocW9wAwuLLi3FoC
P8BmhoCzwb9KhkkKr8q5F4m6LksbK85KZ7wRX70bN32ByVs2XWTFME1+rfR6MBmXOESG2rar1erQ
rIwn6EFuedelnUXCuaxP6pWflYFAduSXrHmkE7qqX+MTD91Z+ie9k+qGlhFvVwVWRh60EWR3tMvT
n5pEnwj8qLXdIRCtDG2K7pOOed8+CvS+eR62OulFPrUzbtvG1nhFf9OxFUlD6qqDbVl5tne3dC+f
VGpAho3jVlFtgS4Io8Hp/w5tlXaGcuNTSX54vDGwIDSj//UKpLuwpzrtaeZOWl9D0n59pDWhGjKp
Ac+uMu5MrAaBgikbz1s2VS2VlOzCaLJz/dgQlzdhqv0GSZ5aKiXyYso9/NcNvzN2mz+HMPu3AEO4
E+Y35v1FDfOwF9sL50S19TdPnrDcOFNiffe2BswXXhnXNS0+uhV64Dj1+dQ7wwiZm0E+3/vsZb37
I948e/VtVvRqvbqzw6dM/L22MiREhyABngikgeWJKhZZQquVfubIxQhOK+A9Ytn2EVsDfEmkf+AJ
QEJRVuKC8JMBBQYHMkFkJt8Okh/LsESNN6M3V5AHLfkFgtdmVLx0QEJGdPfS8KzLhFfumZRTqEU6
vTqAR421tHIozZwoFXILhritst0XkpMvfsni+5l9kRQjLOXWK2xQTSAN/uyNAlpHeL64qgyqhVD2
Ajj/tAAXpzghyM+DMOXyZ8KqAMKALEhXqe8/V1DTXsq4XrjSFsuFbLO7XLCwRMG4jioHmxqT7wv2
tratZHlvGWM0H4Ql4sXdWVHwtLPqII9pn/E7anr+I0RATAMfdGaoOkJGy01ty54xBUKSZnlvjRg9
yAIEr6BCnMsYdF4rjQ71xBQ73b8D+n5/dfHGgKn9nBHUGcgOKN+406CzXO+NoZKHf+KIEeGrw9nC
vAzf7adB008wd9rK8y/i0qSQ67P2M+y9kcFjgUe0Us+E0SZ618A/eq6yJkhne/vu96LTsPpyi3g5
0XJZ3yyialDu09zvX1HGCcW5UEXNsfI/9wOjIDyMWdZ1D84YKnkR/aPr6E0iSncs4+8nZYGeiV7G
VjAZXIJOeMu/StMY/TR+Gqe+LPNNCev22n3JD0w+P9Wa3Oa+VetFIb9AvyKR5lenkRs9+BWAmg33
19R9UsaaoN/5Bzl/Z0VdbAd2PM2uN3Lxxw9YUMETw20ND2yH5tsd492ZtsPF5pnDRQwHtLxd7af5
TyC8RoqqH+Evgm4W43zP1ekdr4MBPLo/AyFPgihjgTARDEsj7atIkQYAkb7J3Iock9xpnva4+S5r
dUjvgLqnbncY8ePmTVihoFbkVYt6jtcwNKeZqERdoqmnDwZobUYcgTN9eOHVMP4xm3YOhuFpUvE9
C1Tc+5vzwtxh1WXkfjZyDStdngfS1OUmtZeImL8z0eAMw565++O3KolPUn77cNhloLQCzDc9cM9e
oK/CRzNJLQY/SNZnfFrIQ1wkxJ1nkuzrbh3Y4kYEfPAtzNxNlyXjfFUXgg4LbEZdUtEeYthX42iY
iTsspya6Q/gMtwAc0J2T9vqB/VV8tDGzGAX/NXJOnJkMkKHXVceyLlhlaSWskYs19Ce1zsemLPq/
bqXK02kgMgX0MGoiTTPVGr3t13q1Bq26bBtJQaRqEdIJB4DgWe3lqYMzhq/J726s4gYG2yANm5XZ
TpzZysfUe947HUJxRao0WroHejgMaY3bEhHMVXr48rk7gv8kDhiqx/0lLZk7+i/hK88eIeEb3t/0
4zYFQRJ5Qzo4FQR6AdCNgC5cwQYHBGRWECWYhOMYJ2y11pyMLgKofd7eJ22Q67HBa3pDPJRgVDoT
TUWIcZIvPELtxELN2Ma9xMV4dFL24238Q99hib0pKwU0gJoJ8wU9TWhUrLod4HL1bW/It7Tw1PIg
VrKr7UY3QR8ZmDGCxsmAjR/RawRvo9QAc6mdAA/BDnOqzI+phC2PeAPgMzVx+TD9A7k1hGx5r06N
vqXCc0cpitXPBlvMPRE6DJdO7j6JsoKFiIWoJHnspBAPSOF3/VRYI6vlHDeIhvDIaJY1Xa8pe5CB
0x1HcEioDQASzuKscRHJT6YiYsT0XbAz7Clb/qYn92a9TJxrAVCthZrjKnxiCy2JfZAyamkZTMmA
ircZUYx6H/UnCHD1WL0K4YlHftIfIyGtqznEcCdb90kmtSbIyEraCBKrIi9Cp3fU1pfUzrzPfgaw
4s6yVnxubBx4NgZ5WW68EwM7GGwUprDdAjMCxeq4+PMu797dTnrQypBsxkaT1Qi7orXysYF9uW05
yvEkLaCa8+HRwaBaTF2DwLUewGVhSL6rV0/PXmsu4Hgy+H7wd7NK5TLaAswPQ+gHuvYaxBizL3/T
LOTu6nEJnULIxSUWlzHLUo32kOFjy7tpONSc0kGgEDdCB0HJ0HGapCOS2xzVttYBXeQCkUREXbz5
8P7Og9CqIQwqe/5eGS+5hMivvl+gPdaDEstx7SE65J08lSlWikSsqW7i6q1xszVfuscjV19A92vx
SqFD3hJBvn3UfOjaxJDN29yG6dffKTUVcB+lFz3A2sSsWXK+rHgTxXEZ2kYkfWOr0OPKYuNTUEA6
iDi+oIVku9IHxmU0sVbaDcWMUI4a0iIxINdbhrU9ytDG+59hum+D3whbssCxkWJLNjwszLTt32c1
kUb1Bx/S3zTZ6D62G+NjYSjsse93dkg3K/KsGlpaAGEg5nwPwuhizbA4S1ywpJIQaO494RmZCkdF
0UmDtvFqJZ22oMIXXQ5/hl57mF/0iBgU2dpoAMpb6Nvchn4327xUFl0fob3IeNamD6y7Fa3xG7Q6
dFZX0eIISkI04pl2nQqOyRB2+XjZ4pD4s+/pp1kzZ1QFZdmAQFznDbrEO1fejskIuJH7QdXt/lyE
rncfsDEcetcWL9kh0nMxf0WYL+IQ4t1mSBtREfmjejASdK62KS7LVEuFhrIFq3ibFBKa5zm6jpkp
/WtdLg3rbTd3lZkYEOYhQULDzcuyQ46nNvlvfWFnuI/qjvYrkbmjCwJ3BDuk/W1hYc1vJLrCidmK
nW3J8fEsnQ8Cj1YGI5rQe65G8YrjagjI1z/3VTMkv5ucKU7TKNPm4rJUZkgjHilzlm1M3/j9HZ9p
8X2pUsohsakkvmrRfq9S0ZBnzx+kQFuNjD2Zm6590kGnGizNR2ospaS9GdsvE6g2jjZtYgNwHmZW
TXL4NWHAZnGo+y+BJCz/QnsnZhe+AuOC4dp6LC/FIDrnMt7Ddqo2YKgXdJg3H4OWQFpCBiLoPtPp
VwUxXuVnvYytNdr31MPLhDN3yssbKgeq5ezidewQXrMRJmg2/qPn64ppUwLUti6UibfutAYKnKoj
ieJexB22h0B2aEHwRSKPRbV8aFC+3SKYhw2j7XGuzXwlibziyiifJccAnqjBBUj4mj4HMlURQW2d
bONF/E5pVfODJwDRufySiZEOayDJXyl6cYPVwaVuswLQcWdDBsxRzSGxaDOypCU1qYhtNHPplU2i
nqPY7dxI7rK/1BgWhXWPFT4Oyv3hZqhR09dL7SP/stKWFqIFZ+HPDKkGY0AEsKOnHn06kvqa97fr
9uLQ1NDJN6dDMAuCMSwFIZoErdfNrkW+MRxeMJUTpV8n6hFvjbfhiZpHk4mkMWEUB+kJ0WJ47CVQ
Pz+OFcUlJPcB7ifuko7DJcxxfKZ0RD1rT9Hn/ZXbiYB6Lz8YWD50RAw9JrvLdwV2Gn2EUtHJNuMx
gKuPBwSFbUqB8FVchQejOSgJzbhwbSX+QF49ljO9zhDMWjaWwaLBS07qtohxVZoO5KfpXLnQhhiv
WdzSheBLEQHW7XMZZ/nBgf7aIvmyE6ODWsUma6kIf1mlSDpzm4UBkGoFK1OGvN47MXMb9zZAi2Op
ItijTkH17R1IOcwTyPtcSUoZJC3BwIfqr2b7wpXsb33QxmincjO0xYwcThPHD2orQi0yVH+ei8xD
Bpp2cZPTuut54ueWNKoQ00RBXI9oX+si2SZO4sYonfTzqSk0cKAbvsnBapcrxkqGekl/WwZAbFqD
zEzkWArj4Em304ei3lFE+hhXmsvxvp6pFjEV5b89TqgeyjDfz6wWFdnwfjJIi1dmd33B4X06rZJR
8wnNkx818qWxtxqo5S4HBUnFE1LjOe3snPIvOuga2cs1Bnl2Tv+3V3yvmwyKGIG/3tytNPg3axz4
rUFvAsKBV6TNBnvHC3qc19reb+h31W98CF5dvqjYzcfBEkMdf7idx46kNA44uT8TFxItRKALJQY6
Hzi1mhqDAxaqqW+TNEKoLZXHxl+VOaehuQYWhGjy96+yTIKNQjZQ/muaeXPUSRkBQMABZoWX+ImS
s3foU70j9HDDlPBjZYHywSsNYyo4FT3G77HYB6swism8uXD6AturxjzXNA/dIhdrugrYCIr/QmHu
oMZh2aH0f1NBioGsQIbbiUrSAwK20/6MS8JyCtH3Yw8AVv9OAjhwcDW0wBJ3zEn+hcBvbfMnghpG
TClBffsm5q3LW+5clMdS613yz+beDHaLSRWzoC+2MjNT3iB9p4vvsUtiu8Nw5LPdeafSJPAIl+nN
FJhH7UbnkZd8cFky1xRQtbU/M3IiL5NEwv1u/w+Uv55/bRKKoC+vbt5etbRWZUfzsBYg18dovBDG
8AIDsczpMQk6aDVmgsOFtfDMi3t4b7D+FzipB8OlyXr8v4lctard3G6+ToY8lgxetFI6yY/V5MC0
yB0gnimAYyGBaTphfa8t6D6er/NKtCLRurNBun+UvfXFQgiybn8AzU3slMDba6kRcHyAsQ4YwXHV
pRwzDC1CEYrt5bpwClJkXdfgLPyVxf09Ua3MTEy+1pjZwtgq+IbYF9K4epiSyvTU7y81rrJSjraH
Ej0pwtCPLriBKCwrlvl9qKBaNdhnDhjtPhWkkKvJnQ1q+/83IDhaJ9clJtSe4PPKH6VIHRyhJTCE
gxS4hHeIMJkX8hPxgVLDFPwRCcl5znn0vUZvpiZ1zryZGfu82D7jDQoFcR8fGiO8Mz0Vu9nc8UjG
/401UDl2P4PAOmBKVxoG0cP39qHKs1hWKzxw+VV/wG0akm0c2Y05ZPMT+LJT1Ej/uvvX5oHGJprm
Lmf4FZaRzCk73kIYSfi5nU4Y4MhO7WGPRT9Ty5TySQq3/qNylrNKsGHzdKWLHYyAJ318kSvSQJ2D
GkpqNGtIhsxr52bUREeOA0bje9rp8TVqFvM7yZChYlIzM3W75PdUY30Q0zm8MO100l8/q1BYLOBs
H1CdQRMd0qCSBeX10QqxB0HPLvsnc2ctFkxcok3gLGTCam64G9OPA+bjix9IghUojEiG899WK5+1
fi0XLeDQ4Oi3BLKJlt7+cP2aXdhX9D5exEu7MNYMw054ik7f8Nyn/xQeknOxAzL95mYDVO4r9hTZ
w5q0/1Rr+W6xSt6ANubX5B6ofXxpgerKNzrslXK7PIvCueW8FLLG0dcRImdjHwo3y5utMn0JgYqE
g1t7K4KvKq0vyCqsTDzRrsJCY4I/5UDnxj9oK4DkAIWo8KEbDUWyVnywV8sP4UvuMqEJ4Or1w4Bz
Lg30vBzfJQh4Y7uSjx2z35IJjMHFBKAmsh7lDNgPc1o7LgudRfyeb2SX5TVXufQf9htkW90AlNMg
zUXIGGQ+hnb8aVWp7ejiBl8nFbEA54o9P36rgGwMtsowFT8+quhRAYb8N7oBzwHUW6XFbXT9CQra
prg/TctHhkN5YvjzV5IepsK9Q2qCFJcPhFKTofz8NuIAClHy+BZYTq16bSKhPLnwa2WQXPpVy17C
/dmPKwy4y+ojVTLN4BLoP3yVztWI6LuDoJ5J7OIrQQ/6/dWzFCUQEfC0H58DwaRuTa9SslZ3k1w6
VS1BA+YgL4BB+Fnvhn9B7pqdN11glOSd6AJRiUbc1xHJZk1NfQj3PNfOVguSIDmnhOAqe0ei4zQR
gXFi37ktgmf+hG2WjR0en1bGuUm8M2JdE5xa2Zw5ZDfFbEFMB2X5DGOSSkWCXaS6jAvb0gKYfmnn
1paS5kW7ZCznwbfUXpAKw1B+BYnqkz/fXpX3xF4r+cTjVJMEW09OHWL2LoharBgHtGJlFOE4YCZi
oZiPPtDWlQLJgXOukag1VDrIPXIQ6KBYAwK4nCTAuFaGLYmxfim7pzmKIu/B8aOdC8C80mcVcZ67
w0Tudn8l6QTFQnwBuBerNK0pYvuwuy5IUuEQLZWEyJ7Pk5fnzW7Rm4Rum/PmqY7p6iVLup9G0AEA
m6tTN+EjI0+Bec6qmPI9s0BHgA0wTa1gLRlu2TAC09kqW8cqePhXxqyLEALxI/NX94N8c4k/aSIA
v4b+5+dOp6pzjkCu8ex7qu2DtAwh6fW73kyg4cdwvFyGWg7wn91dwSQLNYazvxKQELsN2CmB1kqS
xosTkJB3UmKgeJDOQcZLzV0nrq8Eb3h1scoAOq9vi9YdlUnycP3QPmIkqjlYxCchUpPUeCnwczeG
h9pm9ld5fXBe9wmbtf0TvrOwixqGVRSclCn4ruMV08bGrkpM38VTd4t4Xw82Jj7apJMgUM8Ism0J
24aLRGYgYNDX5Fi8lU820zbWMcT7Rz86+kobm5xg7W+LQnWRycyI/qBG0lB367gUQCkvwsSKdCBm
aZtrF5O1hjtorNkvmzEkvBZjEozDFytSY76IgSGXGc/JJl8ur1Fq2rsRkvzP22m3NicvS3UT7uWe
ktsknylU97+r9iFBq5CA0WHfGtDHkDZ7dVyCuFSFNOT0+ssvMH+w6myEfNcv3dfsR9tBQ+oBZKCk
hYTgZQVgd7SYPpBOC1ds2GxAMRn4rfiS6H29YoKPU0lA9a7yOkXeaYC3GUOtVVPevVDGvBRAoamr
iy1PGjWTlTnl44fHIjyhF0Q53J71dzmkV/FAhQXAgFfmJxmCEACrEpAl9jg2NflLz6eMFnsND6vs
rC2O4aG5w89GccgiAQ2bclnJ8bfy3eBz038eoVzF+DD76y+tbaqpnP9sFV0Gqp3674tvogJUcEvv
RTTh+mJhjWYUAqOKFDk6LioWywP4wobDClo3JzQK1LXZWdc7KyKPEne5TQiW9ljOHbetpSZ9xzz+
lBP6ecHfgJNgLbG1dcpOtDIr/NIdDWQqiLk63Yrwp8koYMypLgY2als7kNYqf0Grwu7F2EfScHd6
e7AZ/VZwxqUG8Uu8juJT0nfG9ZMlyZJP09tdAzmoZsmZnCTtmHbmDiZWcjiCpD1vAoZJy85ogROr
+srngEWJ8hzQ5cb/qnvMQgv6iih+13FSA3dvyfVQ6icTXnx2iq5+K8ukY7RN/8CkDkDmu0qmELjD
xBpKblcp8tnzfV9BMWEB9S7g197yAuzDI9Ws7gSeB92+PYLiMWR0dy1QjD445xwAmXH/EgZUjU3v
/TnoXRnagKmJPyxjsStcwGua+jnn49RnhLVpJgbsjunhu7Pb7ih2grpYaQTxmAfgaDuyn8qd5+wj
xJnVz2oy5k8xZpx6+pG1cDTzoJaOT/EHkkRAMzSHbGurV+N9Mp8lUcz30RsSKuIbiTE4vB91nXLl
XxA8Vu4bCO0Jh25kRBUywvKcWH39x18S28NFvyNlsXLQVTRId+NGwsdC53z+3AsbY4j1SPQfP6iL
xGSn4LjYCUqLpayOMCcGQjIddEmfGrIUvesL4vAvqNRpeKq7XLiPsBUhEmsr8wFvRh5Nxx9FYwIF
QhZbw/YzW1Hy2UY/U8D5sOG1yiN4MgHdJUAt3o497UD77jdbyM0mjQzqbxCMius2qq5LGPwdDUeG
pF3CG/QSIeWuPP9jg3/AM5JEAmsal6PfSs82CPviyMJCfpOmgKC4FlDXa7UMdXXp0qLgdj1hG8l2
rQX4+Z8GNxIbWe+LnpW3N6EoxoGL2vDb8ID3nzDX+K1GDCBJdZlWq6xRo8Kb5mOdho5hjnizOeD+
PywJ1A6/Iyg/d7YNSAi/XY/e0EGwZnm02J++AnmVSZdFBBYpThXw+ksoTLF9ifceSvlSYVWMNL+N
LrdO+IYnUwbhTHRnU+7YDm+fu8sX3n7YSIXZaLfpOZSrc42Y/1z2bUFqOF1ewhp6c7Bci/L578ah
rP43ybbmxXz8wglyHfJSgibDQpG0XjqR6+NsFjJxwt02/22nHYvKJ8By0ItJCOoaxD2aQi9UZRWH
qQ1C0053H52sKR6w4Q5LbBQRT6VpmbuGBTmbZBP17MAasENyw0m38+0HWHJaomQQF8SVrA5tWSsZ
RRk5I7QvgJskKOA+usck5Vr9AANvdjtKfgPmMMBUzAvuw2N0waGMkUD5wOTqzWR00g1464OX9B6C
mnB56nudpE4B+78iqINr1f7+4EPD1Ip7vEZtzyfUX2Z1WKdSw9mN/CYvqxEWaCbhtz+yrn9ezrIo
iHaTIidz+rOtmfSF4oQ+pqLMbkEfwE3owG1jXuTx3yF1/0UWzIUdKQil34KclVQ0x8eFqlCkAaGd
fwl1mxVhwDdDGSoY+tZoUEiZNATizpDUfhzPADrWPieBydkHj6whW3pHOhb9GayMts3CPHCJH79/
yftI2REAfp0lQ2Xmh6hkcmLRpxNm5tUh/9/oicXrPWhba+9el2xZj/UB9Lmvjk4MEEMLDbqees4+
LpxN6dl2l3L3m1lSvgSl0J4ZBAnAsag/NiefLG40yETMCPg3JBdIPnkxvOD3t1sAnKEaxaoT6RUt
95d4/YDtsWpgXX5o8qpAXuXEJoNSjHlPvZRQNklKGDIfs8rfzF5j57THiKGeD+1hbPMm3AkBTfDA
DhF7e6Opka/A+SLi9BpIreLE0C2vWIIwq2dqFKAoxxo3yP0Vyfy7REjMWQl00XS2eMCMHCmt1s2V
EvAtPwQRZMiANPDLmhwS+IpNe+NdHBmnkR879MH3Pk2mI4D9xbt9JxcIxk0wCjtAFlOyIqWJpVBn
toVRZg9f0FUHFsqMcwbrOYbaDI59ZLqVm2widX77zAbfK7Plf/dCCmdwUE0DrH9PjElkN2gECZ6t
ln2T69tIarEx6zjAaDqeVtMuzv91LoGlxwFXrdnSWlXB5Gg9RgLNg5TmWLzI/Vlr9c7gpJY1gmpr
1KxZq56rGD24T7OlyNvlKK+MIrDHBmFH3f7RtID0KNtgHfX+23Jz/Lps4lU42x27NHcCo6wr3PQ7
YUwgKMrwPz6FhIshJlq31mBxBdWm2yGgczq7ZyPVTFdZnVI5+424LY0Pde+dlxkHpKr84G0do+8Q
/NInFDKZkoxB6fRaJjyiaOxTlXTKOkubcJkd9TRlBaPTdVv0vBI2TuJlW0B6rcb73wjDCUClrXjK
DLbkoGIs0HHzjwGoX2CNm/K2k0EpDLv5BoEFkNnxsO7C45QAIBwMV+TvyAxjano12LXJZeeDUNdj
pluvNd8J1QCkXCPyyeikGB8TNSKS6rucP8fBUYxIuUlNtVvQhUF6SetETAKoPqexQ6jLuYnbNbJl
0KthpYcMvekNiBcQBryM1TVvVqQ5gPB6u2IljBJF4u428etZM2o19pAMUAy/ktpyM7uWP2ra/fF1
E04AIr1aS4GCpioZbFruJQukCwyziBMaV4/ViL7rnyNaLqSWMfBZp5Ze+ENCRRRKSsa609R/tOv0
Dka4lWbIwi2dVnfQ+eNJ7wP0j6I0qfEB4hbepq3GdiBL+eMGn3lzcb80bARnonJXpH8XDj7RCXa/
yA2/iDo+/PfKAQF3CKD9nr5Mi5al9Jg9vjnJjdkeMxSBuzXeKEG6nNMXIrf2FiEtBeDHUExz2j0v
1ohf8mnPXxlGOATvQL7LnrPj5LBb2Kf0xbCkvyd7+58/SPtUcJw+5kOlxpf5GhBYgHQZBG5Wb3WH
G0bRLCriQN4DU+S7w+2uniB6pUFXOOrytFfjz1vHAwsjAI0m/4FbZkqdswHsgbj0Jrpc52tcFWfP
scIFIRJNEEOPtIHjfIswrZgzH5ESGL0sK9BKc5LWw4ekCFIxzRFzM/z3v+9xxntAuLgdPpySXLkK
MHKPAGbn+NCOPLr0k+x7zg+cXMoHZNhqKqC2U8Bqnw06EpzATJeDbXx5lSq7rzhj99OvZLUmXhk6
RLKhj0wx3SiMJzepaR/tVPh8ld7vlsBcAwxWrKVpl+SD6VWUgX06/rneiZvtPPYZB2ShN+4R+S6v
wPjiF9NyYoinOQNIpD1lLjgTtil+2U7bqtgJESoRFE8fKlKt93lwJC7c821hTgjSYI4GNZO2qCUr
WS6ezBxmNoyBIXOZ1ndTlWpr1ULb7d6TR+j2Z8GvJDiRaAHfZyQGNxgaFy31PlpkKwq3u+jnw+lk
WXJMCRHQriySca4qt1UTtbjxVD5SrawYhf8ZK/HLEjofx1C+gqAfMaPPTDX/94FoksiEaEXMYnCQ
wvOjcqLZCMZg0nkZaRmSp0M1qSN88xp73N5ct0bNsRFAHoytInUuv22HJaK6Kx8BnGw+ov2G0WDn
xnXepd0ndaZHYJQWKwiIkY+1Oz4Z2W/iIay0MR2SNQQ7WwS7q/jNA4QyC4V0nhOCrjwYpJLFg4za
J0CtdC9losQfLpfrtkx3Qhbqqjsbwn7dWKU5WZkRIEh9or+pcVPMmxi1gRdgPGb0AByXrcTwZrBX
UlfHQCINq4zLuwotI0QKuD+k63v3ovb0KVPui4sd/maMsOJWqFWGw2uKJ5hH3DIfOZn45wCPyJwy
MDObu78juJ8LzbpAoTdEnf8OoAtGWc0spitcO1Q4/Oj5Od9WSzg5TI0Gf63/dVOkljfqdNx7URvb
HxnCIm+LOUONPW5X9g72pA9YO3DZTIuakoH561ZdlDUfMnyeU1BlWG61sAvbw1W0khjvEenW4aON
Vi4CWpCZjJBTTVmpKKnX7nN+R3CfkdgtflfDVsO/mnjWDes6xXdLbihSiJXA2NDpktq28UW8UfP/
dERKMocxX3icZV72lZP/DtT8Bz0b8zUb83vIU1ayxu5Tqkh41CbIEAn5lj2Nb8Xa7IIfrLrXXPJ2
rwE2gAr8vP1Pz3E6wjJs2j8nCkSbdsW4T80/kVMq2kEGKB4b3XbBrAPOFluaTzvKDWInxK96qVCv
YnrVA9nr9ushsgAFaADHN2QIEXDaf/q2LEUMx5mXLe5Ft622k/zlfF3ErLQOu+3Yb/Tgp3tF1am7
/bCJ2Y30CNd4er1z06c9c1UbdWvstcZ5Rv4pQDTRq6CA3B24xX2mmRKo4SdOxpnI3j4Utm/n+aIl
HynE9QCIOM3mON0px2eyHHuZQ7PpXlYNajlMqQAkpGWRcXl/zkloDC+03mT4H4CXH35vv38+fB11
zMP6PMV8SJbdlYj8+PipScXWsxm1ljadY7KMNCOhu1Y+O0BP4YDrkq2O10dJs78tez1JAfhuZ0JG
TQWTZMcgUc1NiLPiicySXDS28muDkT/A8X+wj7Tkt/QI/orP4zhk+++SrGEqQJdmK2L08+MneBYC
VkmAS/Y5gHLlsNEnyMgLOUuM0q5rOyOAyk+5t3ZiM8I+yY+B3u7UEpd1jzrPLR6hcBpOHS4grhG3
FyouT4NDUX+GuSN2oYAHkNaW4igwNhMxeg5BQO+l9y2Db283F2WbeXsb9Ik538u67KkixgqFYgJo
Rk8q2AmNJRpCQdrz1YJHBsuTrOBi+wf/HHGYVIv4Euz8F7bYhIa6RkI1+29E25HgAtqGO+3mue09
+vV8c+2vxg9PdnBzxfNfMroNy7nN0yxdeJs9a0Y6CP/smwtHTwmhB/XO3yS/aZ3yDCIt0Hev5y6S
1odYH8GkT0m1bb33QRy9M+Z2td6dk9x9cieVx/DFdN2QNuPySDgDfBC3lchPiMh+MrtKBoUYFLjH
D7tvpPbz1rvzmzvmIlVaQg2mDn9wwncG7Tx7eemnwcCYY7PDb4PEYvZhOWvIgITXXCLZ31/x/32R
QpFYYCPHX+Vgb9kuVKHRo8XzfG1gO4SoCjV6J05YJl53XnUs9FKlDhZfqatKilngra2I6unqwLF3
Rqaz3Gk27BoWXJ8xjot4pfVapBqIJs0o5FHTwTPUuY9FHZmogvddkkuCpTNQGOE3njrGhdMpJwLY
xWGtMjsxXZlxmi4TiYnlMlnEA1momrhz2aVca/W+sQFSvIBPWC076mYAeivYAeyZPdslfSfEY9VG
EV9A0muUkqVFYCfKMQf6Qx6ZXvyII5slKPslSE9UPyPJJsvPUZKDoTtEzJuyx3I1jXB7B5Xxpmhd
r6sDmm54PVRGMQ6q/VTe6zoGzfArrD5mzy5cLBP26zTZi+GKMv2Wt1CRXTPeaOB+YIMNY4WL/49O
PzW1CP3BkZCBYnukU3PU9ymsIbc1Po9qs1ymqQrTux62yK/A2V8YdVPvBoOvFfQ5uUlP/Yp/FpSy
FhEWb4PXd+lWWu+ZJKiIKS83cgMqTWnUG+TQjb8P44RjvhHPNc3soNH52evfiD+XAYOxXX+R7C6D
ti+4cS7YebTbB5U/LGroxAqSu7O8w/ANy+OJeurk3P+sltdHfPhTAV3gY9Tj4rRDKVQgfCMzDyDd
fmX6++YICYVRxHGRbHfKMpfBVOJ3PUXaNkUIrAWud7Tqvfcdv5kehWBNXOyPN6A8QIG19ImFsSrp
u4S5cGzMUwZbA7vswilJWCoyQECCEBSVXcA5y6MCtMNjk9rWxP472mT/AqNiooJsRtc9EuUlelaA
KD60btE+teM707dm2aaiVttZLlq79KmOmRcM9rFE6JHvAYG19P8ZwRID7b3xKhyhBrLGN1GnMBLc
F8I41JMX3WXwzp+po1u/bSjSPb3UYStA3uFLfS/aKOb67hCODMeXr7mC8GhY2YAGRqYhZarzndUx
NexURVxoggNNB2/DrBUWKgvfrTB2vQKyPAxLV+2jcF7sFmmtZYOohdUZKNuSeRDvOgH8wvpJEtPI
bk9r56gwykitSGzqqk+npmws6FJFtnUsnzjHIVSTnGj67I5C50w9teY8nvMV52fkoFBtTJnDxmBC
h4zUcSsGz/dnP6xJx/DZSC+gttp1HSjAHSUyHZfp2385PzOWzlbKd6kduVD+5j8Z0HMtPNGkdYYM
IxHitHID60+FALpLJg2RkYwyv7AxQOkw2FzQkiNh/0WecneK6ll9crN7WlTmgnfTzCvcyHugft/P
RL31RbbQfZjzicvkWpXOyt4wkCGZdqnYl0rfVYEP9ViItqmESD7q17z2gZeEF5PB6g15FFx3dzSG
zK72O2dsH48h1Wk3NOHQDPLoxJipQIcMOjtbsU+IG0dWQ3MBi127mQKyAmAGxR6F8Knm//cnK5Bn
a21Wv6YPO9vC6wcJWwbP6ZiGIYp9mdbkL9wUljPo2AVDeBvQkki+MT6xphFThj2cb2wCSs+nfCYm
1yabNMGZtpb2RGkAcJp8SUroWhjRysxzipW2uDRWdeDc6Rmk7sMDGu0MXPjEgigI+6HZOMvPv2Cs
V6FS2SlX+Jv+/IShZWqo29zo8duLjIZC2ExRcEiFVw8p/0kIALt1+eLBPQS23BwOSIfBaHCJLDPG
1GvZCEIElkAUigx1egoK6OvfY2TblD8qDOvxPFwsGFO3vENb3xAzv6zs8/YQcOHe46lYk2LuZm7V
erJZVLiq9Q9UqnBuF8aTWqwWWBSG0ecnlimSyKh6CAWZB1fLMxMwLYav66zRz+oZc6job121/JDM
6aXZP8SDi/GDsg0EaS9Oa6MuihFcAPMOVsTi0eMFqasaK48+sVOJoTHaSQ/XY4CbWOdAlf+gZBR4
bmeoCC1CZGOJLle4mUymom35tdRocdvoOaZjrCKtumNqq12kmaIWcmQ7vXYAL2InxxLq9e9WFn/e
Bn6EFrGHDD0mFayFXJyJ2Emoq2PpheHP34dqIrCaTcZKIADyQnRn72QYCcagvEbZ5zYRN5ai0iJF
hAc4+wPrUHfvTb3AuD3csyMk/Hze9rVkS8hIKKaF7mfOsARNWchyb1tFa0E6FrGTGLaqezXdDpWH
im8fTGa1kNJEsHn9XmX2d7kXJ4eZnSXpPBflwnwJQMYZ9/epJ1mcEMV1Y3guKSqKpOyntAPP2umg
FMqPMdKFD8y+S1VBPPNFj3szwJrKPMt8VQ11wGwSwQ7yKnE38qgRn061VwI6wewARYAbs3v5gtcR
bn8V7eisiWBxHrNXQNRtZE9SGi/dsfaHNJSULwkNM894/Sxr7o64ph+wzLQwiD6PC82djdXRugu6
umD2RslcEEqJP4jr5Sf/+JtsyBsaNQkP/T8AtEspQw8WEd6uaKDmG15ZKZj8AMIYxAAN8wn/lkpk
79P2YirVP+GMRfEuymVSpUGIaIVIn/k0e3hPmZIPLQlp5uYJDkzCQ4E3DPNZQKvharH8AEnP9UfF
IQ8CT1vBPeN3aA9TozoelP2A+VIncPmR9nEv5kli+MU74Fr/iluYdixWH2DjmC/iEWumRZ7FBLGu
d8Yro3OzkbImz3R+0jwGmykJee9rI2SC19hf+yCmHqd1cjyI/4SVDNgdf08rR8Mi5CBLU40+FpN4
9cZBAXRpM9lIi1ZFZ3IMiNlaRkf44BNrviecDienXBPfSgQG6Etl6XdwuU1e9S4vlOy1E5LQNAIE
oo/pZD4NQja1KS4P6ULqYO8lu7DcHK9eFxOh4LssqHFQe38fxvpxvh2lScTvxOHYRk6eru3WatUu
b7T72KxfdU5IsAfJUg+82Xk9Q0fzHNxiGUcR/xw+tyU7UpkeVYUsgnYNBMustUnRSrVC6kZmJeVH
5qJpxfb3G5vZvh4bI8bSzXKGEl/95d2zOI1KzaWwyp69bKuUXNfolm1/7k4vMmHA4NS1USyzouy7
g2KDe964gYUXQO4K3OHA15vDEmJtopCKcFsD+/hdbW1uDo2jxAgmj+UNkJEj4LwE4q2Uk7UZtDhx
eC2fUjM6nCh/XzRu6hVV4GhdOK+HwoUD0FMwMi+NY1mbTJy5A7PoGnJxH4KmkJKKaRPt5gtLrelh
ShOT5gDI6M99Ia+teQ4tfoZ2kd01evllQsyBe0IxRLaDiRuSl6OeqOYQjuUd23VrGqiwIMi6ZDxR
rrnQg5051HC+BHCil7mfWSfT1kdCfEc70XQDpjQWrEHa2R/s0kb9XBf8qQ+id2O6Ir10CSAPAzqW
QMVtMVO0C2f6qe4XJmM+cjKxFj1pfMzmOICng4ULE4SkKJ47rws6u2sgRQk/NXu53uqJTjJBVXd7
17+LiGmrdtqIfSOaag5ST2nX9KOTVtVpJxTAnvQW8iNWdV2S3lodE7rXWNTU/lZKUyRk28ttpIRk
mgxajzCZZy7Q5LUBOaAb1rYTXWfOZk45Y7ddYr35Ing3dTQJd5ewG5QugfDP1gkN6i5IdK/QIc/M
MmTNJLFpHCnnP6yckFY35YyeZ/77Y8u8GPcqtAQBRzSNkwD9CRnN348VPFoAvb0litKsOKC6BGJZ
M5PffKPsho/ntRcj60TyJxEqFueovepOIg5d1zwVe4wjbgZoft1x0rH3MpV2I9JwStf+uFjKRbFK
j1TMY1ciqqMO3yDsPgdKtXFb49MG875p54gUAqZj6foP3DsBBMCdF3vhu1KllceipPJ4y8FDPauJ
SlKjWVAjSA2eTo1eBK8NKtj/kxZa6arPX6YSgMsN8DkHgX2onjwz0+2OVQBV37RVe0wiMJHV6UIv
vs/D/Zti6YIo7lfK11WeAq9+dr9/teozP2Lp1QlsjZlHO+FO8bHnt6t1O5o45Ka04i9i0IqF/PMI
1cX08b3dG2JzHornr4sdDOLEkcoR/iR9ZPaww1ztVsBNENY0vPx/iSg6u6Uz4nmGYqivJxR4wlG7
eFV7U7xb9x2h7GBY2/rW3ey5npK25aL5yqOS+CrlGJRlN9tj/8PkJz5teAaVjKHeAJPyzETw2iGN
tiSYcINckQB3FnxsfJAsTw/dNyDFEiTd+Wc0LXKQQaElnp89aTm+A/8eTD9aUtaB275T9blQV4FT
XuDIuvLCWFf2biV/XnFGZPLzO6k+T/uJtkE9aoQqX3jp2pPyvzCgfgeJ4LKvEac1u2AY8PrGG16J
u1mbgaakpfrTAMJrdkIWKCxSyCs2VXYBiqzUZ8EY4cDWGsx8fTx8WlVxIST0xjK/S8yB+sISMGIj
lMuEIfSY0u5WeYrlrwIhrEp9rdiSbu33D/dnZEet3kWyhpcrKaS0P1TgNQlA8OdoCJcX47SGcVNx
oOaVDlIXIW/bGuBLYVlEKnblZoZBxkL9KQD+/xSGsLlsH4KQ3FDU3nIr2m8+Cr9E1uEX2gAbyJHw
SFzmwF8rLWT5XQ7X0dj9b1y+n9sn4CZ4ufab2PxgUkwd96DIeiOlQNOdacBRTNLTOR5DTqoFjXrO
1jbFdLAOamc30eYoOLYptDiVL8ssjTiSpawEgtQZAZefU/y085/iEBzsPi1ar3TFOlBXypS1yUvP
SBaGZRnSZUZZ9F01vtiUqr0kSscs+PGLaEgfjo0d+xL213hWdl42NovPxb6u9whsJibC0HgiKqTu
KRUbV0D40wwEXhuR1g06slbpHTWnXmwjpwrUg+VJqutFLF5hgxJkhkSS86ATZq4nCsc2VHnQJYpa
F3QRrLKUhg04kGBfQuXoqFP+eqtS0vwb4owLoIE5EBNbnkCLvwJigjG9Lq+RtQMLJ952blUTg7ny
TKxpZAhI7FdAPHYJGwscR5XL/zS3IAM+A/PvRdkURzDCfn10dm5j1jrJAYgCy5e9MWcQJ/cPNKQp
2fg6a6eHBZlGg9mplwT75NdcskmSfmFsS6yttfi3zWqUNVSv5jjUIqX+Y0jn45UN5Gmp+78e2jQF
X20sR5F3sM9+PAGt0HVJfyC+l5uxualBs+kyzgvIG2ZPX7vTl2FMe538K3DJS2KtP919UQKW7gd0
mz2pPnN0jSUZyt/zhDnFIQDer16xI0Wj3pnEHPwS9A08Rkv4YSYW6mbGRBwB1Mt0cGiJUGm+LX/O
GpMblw4hSSNGINq8GbvDUDGNUnRH76PB37esKJfc2ZD8O1zinPEHbHycro1qgIAvjO+iOXW+2Gtu
rvtLX2e/swrLOEPBUTHTHf3XqQYHKcRR96a3FIvRpVrTvNPPSezzt2p2AQFpTwr5AaCaZTkGk8qs
IFwlU/S554AQjLoMGpdf3lfrZUutdp1oNQnkrvWjpvqvOf8RrA8XqPj8sGpwu/US822seigefQUT
mpV2VmrC/SL4Nku9o/CNCGX66RfEKk2jK0ssp1LEAPlzCprhBh0lmjHzyCGgFrU9M0Ml9rv7V5lf
YDqyIZnOe3V85jwRfL9BsJByNzzNUtwUbLxKrtZuxhvRgAKPRGQi7fVYv5kijvnsDLsJHccJ0poM
vGEk7eLfHdLNspkcGMwVRfky/EbvQMzSGT8wLWK8m2N7O3ur5BlVODhcKNkdrcd0tL/r6odFJWga
i9opFeMeKa0crQnEKUWHka8N0gkdWjQbU+I8z/b+XuzExdtlv8HuDAX/TrZZfAc5biEeHLbp2PYd
APhQkso9UKs8i4Fl2iArrfdod1MU9Y/Wh8GeTlJFvgb+PXaRvDW7d7yX9Q4FFLNNVK0k3Qmrg0kV
1tTEijS2LnuSZXeImY4OSwdScW5kGCsVygr5Q6JxoCh1Gk/C4AP8SZTI4Wq4gKDK3a+g4MjEIfO0
SL/7fYKgRPY8tpgxCPI8S/bMTGe3vyHaOEXU0wgAlFbo/5PcosiBhtleBaTfddIPAORM9RIEFEyF
HEMNahoNejxMYvurATuQ3J6IaBvJBZGkhOqPmzj8FzHJW3cMEKnS/c1MmgfhmfdeQmmlUkfi8a5O
PYrFOeDlffK3arb+fuY6Cb0h4qV8vm9iO23wKrHzeV5FgdZWcycOZbgC6uRs7tQD/lxLMcgfDLmF
V2WK/rDjGEGutuSiGH7ZzfEZjduakq3j5Ha7W9OcC9rVca9wEqahuVY5HEw2ACIZfptGstdj2R5L
Rf0V1kDgjUeQTtwYVyC76qmurqjpPHRM2MJkX2GL7aLXoDoH9Cg7wdKdsMDaJRcAenJqo+J5iGPh
lrPhdm8pEAyfF4ZwBdS4duVHoqKekWBcIefucNWWSpjrrDwwBtVFuqQ5wVTgfp+3tyFq+feFHagf
WaYg1wyGapz8utYEMgHR6MrLM5nV6XbfOvQ5rnfQ63vjhjyWfpMMtt/w80d0kql5rZjNbKiMq8yH
ZAE3jhu6QAgOfzOjTLzFhRuALCTS+mY7+NvMMXTQoTSSU10JNPlb11/r1HYQcCbkPpN91cXoIERY
UuHMPoAn1ieGfOULpuujrHyAuOksjC8MhRn5gr+9Ft0fpyvH0ILgGBLVtaTv5rfrujUMDCQzDFXC
xBfTAI+xKcbvPyYFRIJGXuwttPWaVfG2Pc0sS4yHXOvtsSnhZqKlrAWc9Una4WxNahr4fd9bJUzF
oSJDiTBHUJ5Sw/rtl0HbdalteGE7lr6vIGhbaNPfEDr9WriBKJdw73cgesqKufM4k/+N/UQ9Li5f
Y+RI64RGTzSq4PHkLXrjHJHU9aD7y0VsOY3v+JSNYaPEIGgCADXX+tdEItDc+/WgyAvV7qEOy4sY
990L4rqLGaaWUYlVZ5Ac02uxxrpX1QrI/MdwvdQ/ssUFkEo2kDGctLFtV0jZSi7uiwxD9jLcZAAO
+dU2oqN0Np96fhYObJBYeRPXpVZEP8wzflteVuXCXfYPy/Am+KchjK9LrjdqX6z1m8v1wFU+fImd
pkxn4XQdK2HYmP6a8dWLKZfOnjb1WzcFqqmr3eAV1DpLUgwc1MknEAebflMuCRkYhX9g/+CyJxuQ
L3WgO2AizXR2r3gl/hhtJYfZutz1V8QXTvJVYbOBnUGsLMbQbZmWyi2tgyzwwTgP0loZGbbLaYSU
7QqwT1JtIhNs88A4KgVsKPR1fJgnM9oDcwAk6jLw5MKDN7IGHKmKt8WkysRVh+mWhfYdNK7+YvFz
wojruw/hNf74i48T8WXNw+AzagICFF386oZ2QR/14S26VzsBImN4zOlNT2Ii2/Nevek3idVWRR9x
A01jO6FHEUSdn5VBL/5zdkEoIDsZaO1jv941OP6p3vBEeFiKcHSBhJVY0A1k89BuKis/0WokWdFM
ZcOMaADg8u+upAfRGml+Im42FvZIjDJu6/Nv/fxa5GlKgYEBw8iHDiXDJKEQO1EEHeE+HufLB2jo
w0slZ+2QfYs59rIv4eGDXqvyd2PPdwbSeALdqd9NFOIQ8UxOzADTQ7aEcKqSYSEGHhLgPjkYuC7A
vU4m6Frb+iwkK4qEvcHjbtIf4r14yTbBYlAvjewwvri+crOrQFHyKFK7tvsglhct/FEMF0WygZie
fqYMpxXYCm1moNrZzLOmBdnlbr3gXs8+ROgJF9FHZhQ/z59yUwMP8G8z2GSW/ENO/r1/9QMB8LfR
h4lrfN9DTpH7vtdkH6ZMz8iWPgKTnx8FNBgIPBLLh/Pg6bPlETxg8klvtRw5CzyQIz5UMwSGpW2m
TpASz08uj/Fipuh3y/wPrCrv+aiSqnvUu5yMtjrUV7Kr9fVpVK1ohGMjvkih5oUrMsZINDPhcOXI
Z0k1BIJJw46xisz6xUpSBcbF5RZGKmHEdXL2hz37CQ76zlSUIeNmYellMZn1navtbF/iPfQBUG2C
9jMGuH5iC1a/qL/YBHVdALoPt+09Kwktvw3MvCBal7guurpXuDDYJCwjPea8Fn2nBUfC737s9fUR
NklxcHKfgfuLmBibZvqlVTWpTju8KqMxWQvTEh1mn+mJLCCtU139Ds3GYTcUbOm/FfabXtNVMo10
HYqJd+Dpagm99OrKBI9k7A0qUX7Ui9iuCN5aU7COxTiVJ1FImm00Ytu8SoOxomfW5GfBHL4IMqJz
9PeXP8peoC4o/ufhq6ZVJU1m0pyNNCIvYPT16ZG8FVpZqimcE3d1v7mGUw90fVX28Dr3rh1jml18
We1wp6ffnhxUGh4pPZGxDTvAgHyRZKopPH+1+1FNbIupYKXFmFkwRhKmS3FhcHEy5gPPKkuwzlh+
WIR/Db+aTnLpB9gO0Mon+r/WgBANGlc6YrhrVZIue/PuKMLhglfF1c05zfI/QaoF8YNu5VGo3X7P
r/a06jLFc0Q3ZG8CK2YtT6fewcc016N5sfuSaI5GtXPXHnP/Gs72M3NTsuTAIIhKvXrmjdtgHy8b
gTRZ2lOR9gS2ItVQGaI3G0wbL9tjQkbJJnK5hqnA17lP8SkG4YTaLBPQGoyQMCXPqDXRQugt/im+
lxWBz/yER9gxyZ/mZFfdvyq09LvWPPBfVv7/zRScAYKdRS8FPSoOZqecI19OeDsx578d0bgbDCZH
j2Q1OKbR73B9LaHITU3ISZK30VHZhbm76RdH6Ha6noy9cYYL5XqkhDniD8xylXiYsS9FvJZfJDFK
SwNyNeeOlzyKZloCBwnVoQWNX0+56zHWuzwg2qcJgECpl1MIeBP0Ucmj0ZgXSTUOkCabH39EFHHi
QY0gGQbMp5uRixX33twBI/veCIubbOCpCQPWZsgXeGOkpFevzWLzmOmMmm8lZuAIOsagKI+x3drB
v0qlfl2vAXCAJTFXYPox29FY8q87aGEXUWA3012sye6Ke+XKJgiXpgArT1rcjD8tWEwRH0C/XFLd
GDNrFJKENVTv00oJ+SCzrewxrQy6nLyYz3vLsDy/l3Joj/D6KUwgQQqaL1TLayt/AvdrGRCcPF5X
/uf6p0ne1hkIsJe4ExbtYGlJ2ZwAOOE2UTKdPFNubPZ8utJdbwDG3AM+5anfi+/7zWktC2/xB3kz
CHLCy3bWW6GNO8d0HdZK3ceN7ft+X9nyuZOpyZplJ5W8nXj4tHnDzvsQ8Aepw12EqMd27i23yqRV
m7OPuSXxRAhQ7V+McdffXbdv+yQqUZLFAECNgsjKqu71G+VbF62AbE3hskvWKYDL9R6G1wBO4j9F
GR+wi5IOkRaT1klzQDYQGHS7iy9+jkrLwsPOirgeyc/glAFem1x201n+O7x593CnUhRDqpeq9DiQ
CWMDSKsvEJuYhFB7M5t46QYdF7KQ8wxAybK3frl2oUhcVBkHjJCf/C5dlagG1wtSCh1IrDpShTvm
HWs6esH9B+DMCu10fkrI7P72PWItlK3Y5JK7nOFW28HaUbBQawJ+ToiB4nPdZfqo01QuLr0q+bYq
z5HVMvHlCAWaSGC4tFyq9NeTb4HsCvsVrIX3BBAzlm2lWdpIbSBpjUolyxXcxH/G1YOup4ohyE+y
gtCM+gfZstZahFoaCg4h/J3B16e7awopnacV3/VHqwAuYQtDPQ3+Pbftn88UxzFUbG7dV2f+OiAC
HrB4Weoqr2AGeHyGFs0gpPr17kMDaMGciacP4VkT7+90ZoV0jkfgHtk2Iq2pyRRnLQByO3q73qvm
xSsaPIlA5UQ+PQVP2rjU6iaeMWvXk3NT86Rhd51vQDnoYxWgV5Bqvi4zcIRpg1I0P4ffJgZO73dg
eelkT13148FX9MU/Qx6OQAXHZuUK5PDhNH55udV2MHK3iKIoghf31xPp+dL/nXk4a3+6PZjiFdPu
ZB9WRltN4J/J2vHDn4TMSQR7ADYAFLm0oaAiVyLkGyQi1+6AF0mPe23M/D6QJXltHM3En4De3pYI
Ik0LNedc2vEvp0KuF+9RvVdlc0Soo8NA/oWv/F2Y0oNQkTVlrzJKzguy5eo/G1X9Hw9cnBWuE+5t
leuU/N9C33aN+JcuvmZ5Qx9Rm3HbjiWbUgrAOHB1ChtdXN/PnmjzBykXSooaP4S1K0D8ZuxUknir
DkYhuZaC5Zn5/olmOG8SOFzpTpHhG8Ygf+ndSwnfsWrLnLNExRBNh82EgziSQqxsrSAMmqFbGGDj
Uvftd2mTuYouOatwQOgoL946o07HDNEA0PO5E/PH3+MoAhWsj2O3O42suhT5pyaqaFmRy3kPO6/a
531slKlWyuVGjwLLCs0d/LW+IwFCiyq/wh7JF1WUuwmua7yol1fPWGXda4VGlBJWMy7VNTXfPUiT
b5FNx3/Bcp+OtvsPPfqWAGUQ7YK/d+WFzDn0tcMyhiwacxlYinJceIu5OMp0HB5HKrkAT2r63fRp
wgzQwpFc1X6lm+3P5zUBa6E1ZEv5HS2iWK58Tl4HQGDJ2eMyZdr79xH3DauyxhhlMieiB55A2FVi
apZhums+X91ng2r3WJHkyyM81p2qMa9gltFAIoof2lYa1+wyQqTxGPP11bu0UUncAMxJglqmfYkG
O9ao3K0Rh3f5cX14VCIeEIHSTVYT5f6P8DBnrflolaVI/cQ1KQEZqs90GYNEEPm//WBS3vK8Cqh6
bIJzUGMPuLcztUY/N4g1PY6FGSJKZh0mFzrzrDCbL995pqAa8VlAIYK5wrs3ipSLL+wji3eQ4Aua
OPr/2zHOGIyUKa3X39vbdc+RWV3QB9DNKSMMTLt7A/pGm3kB9KtEImDqwhmJewSjRtZPQOYVmZDR
LR9rOHppT8WBA/lmveEfBYh/XslVwntlSLEaSzJ3eG9ysrRodqqotIThuZdahTDuAT1mu5P9qzyz
SlS4QedawQfxwbrcLoI64Ti8N+A5B2fIixNHQmu/Ej996SlQX7sn7RhdTHWl/mKxmJTTwB0J0QJ6
am0ky3537ZM5YXp0B+ySYurbyMDoQvCGISAH9UzkOPHkSPYyKTaEIHGpIy4J+IU8h0rL9H4kR+ej
0ezTpMm6bkuNBokive7bDbmnhA/3vy9nw0VfxYqluKCKZPXdVGAOs5yYtUZCDd05NzMNwN6ET1o/
qgHah1ozsWZQfqdkMRC9pwXab6sh7KVJIPVcy1YXWrk5WjE9svucZouU/i98GKbz6RhInrHdrb+9
dhXnbktDPXBnt1iYqlj5zqUKWWW9I3qZPPRrjEqcT6vgF5zjISeEsjfSREpbm0OHU0df7wG1ww2j
exJ62yX8VF9WsyCmyZ0TSjEMHeGNmwcQ3FsXFM1ENU6oqhd39fd+znmA9fGopABj0q97jR7x9F59
wT0vlvtHu+k1k4VNqcPnxfc8qurhbYKDRyNb+4RC65MS8qRwwoACMo/Cw686Muv/XwdrCW8UqTUu
9VjjZbSjEt4MSFVz5qBh1NRRpxz9/8T1oPp7Qe0HWmJ81EY1UqIszSoXT/tKlAvwrGj5xdx1hz+1
fuLiPqxshLEyAUdBmOhTs6aM2D3vhIlEu+7ehabFuh3qIqaphvVETtR22ECB1hTM5cvXfa/Ol341
lLI8sJzQSoSCRyUDrshdkKIlHy4XN8uuoUDanjS+mQtLmdQKGMREXPCHGG/nr/SDb1dzAdpN9DT1
KyVvz8NqsVhWIZ32wdmBshjJl09z+Jc/5cLmVh4NbRbVThbaLBBJBijj7w40mHg+xIhc2uFP1JPu
lzcoLHQUKxN84fYSxPcd+8mmJ85Ji871w54+50XQ+gSRFqFqZZJ5gioYzkZDlEYUuPpIqlk/YHiQ
oEHbsmaOdNT96J5j5FPttqZY2GACZHdMnnPT+rwR0IIyZXoVaM0hFIM2Uc5QaXru3LUVKRTN8uyY
K8js0oNa2B3q81yeJYSb1K21+1i6U5WZzvq5NfVXOcfF3lJFdqi4CFiKVBVqKZXevXa51pHSDKpx
t3fufBEp4z+AAdhY9z7D6og9OJ1hxu7uCr80kUxyqpGG3gKYASp7AkKPeqTho6KfddMKllX7DcH6
xdzexX1q3Ihcz4Zet0BTzcAZzeSj/cIBS8xD/kC3OZpLDrmHTlbH4ycCZSHvpuuAIt2hi57MEhMU
JdT4UYFpcyuKeHZ0i9fxGdbJJGSdEFcHCadSGKuIZ6lX5rqF6oiFBDPL0nyjz3+droetJWsSsEZe
QYrBVPJXlLcQN+F37ZbAThxjzvRFCvFqGRtOClavarGDPmMNVSswkJxkCTxWud5BenAyAvBVpQaJ
byR761is8eGy5nEEPWbWwkPZbGpvGMiynkkXY9tIwuP9XTYYwdZxCn+Yq3EVJDMSO4AHGLUXsbU8
tGxDClmQ3fT4kMAi8mt4bhDOtVTfy0g4D4uMSNZplrW2znNMyitnOJBE0QuvQ/dO0csz9b9OvdOR
3lIINOOphzstc4Jg9S8lZU1clxff8jocjNroPId0f6jS5rgxV4Bw/RtFIfDNvv5Npgww2glO6ajL
cw8RapbV1nLw+tG6U1cqAEvGl2QCtXgj2ciU3FKGDl+20cULEvlyWc3WexS60W/+9M3nyvPJTwEF
YCqdFAdvpOUkyeQtp9IPzTRxLNwVa0Sf5UwsiuPRgOQDa0DfH8kpHJqhwbtjMhTDfab3liAIafo7
I2q9uKMUofzRCh7WNWJrXgBZwV2f53vBydNXMOyHxcqzKqen3psEdStfFYigD2AoEPGxVaoHt89M
6ArQuGGpqxlO1NHnjCDhZ74iZGndceeikUFu36uVWVDQ5u6jcZFzbtp0OsSBIiZ2jWx21PMAXTXo
WpJt2FVGJtCbGoVTQEmy1x7ufsMlSKBsFNN4/gY0w4J6ItjIKiaRkJwhY7FboaD2RnoPh252bsQM
shxz3NE9VXlZN+zAjGSQMUXGqaRbvfXzUekpxsPKDFBoLBd1IiGQgFIbJEcQls0AllMCJN0xaBpv
Kb7cDViEL7d5ba9WL5nVZL22KB3EQP0r2AnIeXTyFGl+207NEh2cnXSamSlygTyJb4i78tkNxbya
u9CHNryzeUHMFwd86636wvo5eFWFPBJL9P9VWdd8e1MirqQ0bieeKBoBSWr6bMyB3Kmp5eoqjeWV
1KD/D5yrQzTDkqqINk6qftTPTQg2DgwL9a3sCj27vdQcQeneCVZA77n+1B1ahFpXn/We2jwPbezN
WNRfjoRTVjaBpHiCFtcyQcVosGjVURkKY0P+cBHh4HAa3E1nfQsGPQD0/DiI2lbVpIMkF+cxYaKR
4YBR8Po9xG0Qg272dG//XmSleLfYpIv1wvSFsrDz66JFUwClz2GTpZz8GhJVx96VlHU4ZblAUsPY
V/m3jN52nahY9bs+LDjhD+zCshaTAswnAYNhgF+4tD+R6Tci9MmkKOiQRZWLi7mS2CMfslH75L8+
iHuH49qU0EQJE2usndtRuSvEE6vw/giaJ7sSHicJT0xMsP7ymI7Antr2mkjpj+KeElrNmLUXmGGd
FC+NSueEx+cVPb4eZmIp17YG22dUf86U9Ll6Mw2A80TjC/Of47lRBAlhoNb5cmLjYeUYyDM/9JQN
rBXbFva0ebxMEi+oRC53p8LemKOETLi3t4sLuD2k92h3BlU9kateQLmen8LLVL14GCLS4qchWF3B
fZfXOsdBcnOz33XZlKa7+IW/nQXULr3K/SdICFS8Ym71qkiV2KWkFydI8B8drMiKz3VBQCs/QdJt
bIAtACANE/Y5CbpjJsj4/ZsjF+OYA0gZgmYeHvZLcVAOe2eNEhui0rx6IC35uRx6lDn1YybnBxFQ
ZxA+tRzYPz1xDQPGv3RAbOJMYLeRU0L/S3bSzhV1UGA+wW94BcVtPQP+j9iEjr0A4lE4K/2ZQ+EH
RNQxRvMcsvBk0OyG8S2wyEg7fJFBlxYf2T0ebl+TK+4QaLOwmFxQteqJy/JUHIgbBXyqGP9HG4hb
B4fNy8vljtGrcLMZl3ohIRUCSfnHSp5fHYRlATAVgpVN2VybVN8zLk8Sva8N2TKpyVdsp+ZpM2nY
HxdjK63I7OSs/hZuoblOsUsmlnDBwzA+GbNYQoDSH/fWP5GLXyQRPUdKAMlsx/Y5RxWGkS/9SNr6
sOyat/iFuwrAwlj+1gkSMgmpnA8CzfAcUZMPTEac+I0RiF/TUKFQGTRyjJzGXqSMjLGQzgdK+E9u
CbN/FDDCHJeGoEg+3++zZennHII4g7YSH5piYgj1hopxLcUuRizSLfxLmvBGEGxLJNGsP8t818QV
6Ghs6pjoulGJx9Hx/cOguxJdbuoEP9yLvJngC7aPtu0TfiCro1qgwu1GVpYwe66o5kDZVqN4wtma
2LM9Tnc0Eby2W2M9C8mCnqT4d4WYLP12Z8e9rYgAIly+FNx2PS05/DLRo+ahW+ZxqS2471qLRcan
1hE45l0G5acetZKADVHLHpbJAHUOG59fTk+WiiKQ0Svf/O/CQ9loJjp0cz479LzveBQEBwP6laue
dOi7nIttQrEYM7CWyeyTNGV01IFSmuDR3QNI8GrDmDggyxBR1zlNxFiBvYMh5xnafBF6ilLkkL1V
D0vSrkrkWYTOOuMn7MY5ASxCKya+/Y3+0/ifII18C8uKYPG5Z6Wl1AqRsty0798uaDSrMZmKN9QX
2Ia5pvmLbrGIHgEtwWkl3HBlQUThf6jUaL5nUsUoeff629fcPtMI13RmpW4CScZkQ32AYMnqFH0p
mOdp8aMjzXefMHRrwoUeQVcJLcBvId2XboaCfrjmQiROSjTeaHhyaOYwbZI9dHtqtrRfo2tx2IxC
2ts9TCsP0PEMCtuMqvv8VpC6ZJa3Zkn3pjOG09HVyBHaAjsHR0PlORGBXb52ilOgmoc718EDXlYZ
FE05dVstxUKl/Y+EZRU3U9unl2BJSPYqhs4cQpSvnqsSfMB1U26yfRZDlEHuohgAo7i/yngQ8aoI
FKPU1esWg0d6gBYx71ZCnKVI9Kr1GfWliuHgjbY7WU9ho9BBNEgwvunzehTgQwnKya3xfeOdE+/a
mTL70+E2aSWZuOdHiyMrsT6zjlJtvMReRfOH63Hy6ezqDdt7I2A2asIgVnVmOfPo5Z0vNE0njacg
aDLbs5rLjC+Ex4jsMBGABo/6bD7m7b4NIZDQEMLM4liUWHc2FzjATgAlRJ9c8KtbOjxLTr8sMOzH
R3wjEjNugdutx1qAt56LtZhNNTYyQq2ioHaQ29pBLzfLHCNpDMEgvQ8nvUsFJxnNPVOCg6pzlHj+
J0N6ZpH1vAXaGmS6hcgNe4MZRBLOKWZQp7KK2wodE63kYkSAyTBiX2a7LUoTN/rUYwplFcivxftK
mcLx/Oku86k+EmU8tMsMSizIbxSk8XEvsBZ4OaRblPcvBhexrkV8l9fRKDAcotY5Fd/79Su7XNCX
a4RUXzCiCibCbshBSlCJiFiN/wjQxflH913zqWqBXHxQ2qZGe334UkeZ6Pp6kRX8hdhGjrds3edV
Zz3GZ+zfQpbxXefH9GAhsDCK9KBc/9RqhPPF641Bu+uhMOqkLmlsf2wLxxpjTMJXHAfOnjCDqhXL
bzgOYXjI842yQ2Plf/lT8Fi3N/+AGC2rBcxv+bQcfU/jYswotnXlgFXRkpsfnFdX0IhNdoFVfZTa
i5x1aQrZkEwJaoVyMSU61RKPyq6PwM08n4C4IGVIoutwHRSUkZNNpgR5Fby/HCpsNAM8VL+uCe8o
Lbw2YYFbn+FJ7IJvRXbkJVWtzOv98e30kSnGV1v2Grate2RfX67xHokCSqGFG43uWYQrugQNhfLD
RoRhxhfwFKTsX3IdEy3a0jhCvMI5nEqIrwpn/bfgPiNH22wn1CczHXYhvkj7bWNIO75p/esCF6Ko
LlQAmFou5WsLi4UC+EeGnrrwEqNo8EeJpF4g7BUdr5zwORuwSGMrC+5PQB2aSamNikoR6E6X1X7d
Ct80d4xPlWY206iBCbXsk2tPlF0k4Og9mQ1bl4ob9WUoUNhORUu8HBCRq/slhdObQTnFDAH9rt2v
trhGxUAdnFB8kSl16McAscjoTZ0tpV8UZYxKsfLGVPbpIVXrkzHfVXBTNjwJw9ZVKFfk3q/p6W/t
0hZX4GDYLAgZ4Aftvh8BfIRc+VanEh1wMp3XfOp2vMpSoSUzK1+qrcOctYRhvg1/fBKGjU45LCkw
88Zge40Q0f7DCWb/j7Z3xm++BmN2vSbIN39bLXA3x+v1IIzVb5U42me5IWHYzQrg1bIfwl0Q8TLV
z0DgX/Ob11GQkZ2I02fTuDg8xt6iG3Q/jzJX+LMtngRjQBvV4KT7J4yAmSgLZ0/qnjvg0rr6UbRf
/oSpIuec5pjLklR5h4a+eQa3hvLYN8pbMuEPlhKX4FV6HwcXs0TXLNXAFCfCWkbt+kIeQdVbF8Sl
kWc0IggJE12hy2sQMEMSkcwqpuMjE2cqU9DCxqso5DpUQBJV7PBsvWOYApzw3Zp/9Z7WQEXJvl+m
5J/nrXxQ3xcVyoaHHBHAAcgTtBOCH9FNXT3xqRchz7YbWKAJdwAKqmRbP5mPtIpaCqY5aDwojBEu
yIpgA7GrfjRhsFYLv96yO4XWz31SlUudWWBz0jKZ/ejIdZo1FJrfLAlPnQkqeG8qcwY+Ldn7FLvm
dlsb6XZcO5PHLr25vt3mvjRw0jAiEjg46KWW/U94K/CZFk1QoHR9fJe/TyBAXPsh6iAnEl6XJySX
edpq3hsQj/XQwXM9rAMQbMLG24CpbQ6586LASoPnrKULWGNiloaFit/qcwEB/lk7bCfmnKMCz6ax
Gsm1WvC6OhZ6AlAUeAnpkThFkLe5p6fozQsw5pZpmtl9IWK4ADRHp2SCt9/DjGvvatDozsCOghln
gR9CUulMZVFqHJtSqeGGdqxUUoUwPeZs7Y61FfhGLw2sxZ0NL8IwTE5jxVHfqlKCfz1eK1SKO6cz
9cdFlFd6ZpOVI/ghRjcPT/Xof8x63WJchNShjHFARwZsdssYmS/m8xdFhHjaGs9aSorlu6F0VS2B
9Kh75MXfM75CBi3YAbVRUNb/ps14K4d1opNiK2zZqe2xTYkHc4mhDim9gB0TwXCsi9r+zqgkW5Gg
MD8Xui/CXa9ki+olsXHboeX9CVXMSBaUt4yG86iAOaUmf0RhsgXcQymrAEzBCJWBmtSll4UbcYAg
CUSSH5qm49maqOSA28f9SHvXE+YJHmv3PUhW7MUUD+sOuS9dk7/CNDyLJ9n4Oeoa7zKooPSRqWNB
p8RnndFLAiQ/PqHW0bh7Vn62t3GraO3EDQje3xeMr3KCMjlQTFaxDzFuq49M5xwE0YFuU5das8VB
FHIrI7n9OZbipChodTx50nmY2LZZznalB5gF+Le94+MYdT9/XFGpPo7KaAUDdq0Ly+Eu9DgximyQ
LGtDtcuoBRlEZ4XkMcloDL447TnwnQonzZ4nlKOvqx7FgIT8TYLolDCI1D9Apv1/j5dekGEs1a/w
QEpsul3I0vG/bWCQDq2+JHvnO7ICHHBRHAHF+LDIEozAItQiLedIm49omlmpII+mO6zeeC+YJpDv
LbJuPkVyuLAXHeBx/5dsJjJdxosDozGxl07+w7XOU23YP/T1W052Og0Hbyf2LS52oywd/BrMNVwa
rP1EHpuRvdlA9SidF1iSIUQfU8J+8sd5YK5WnkMCyXKi5ZSb2Y6eM4INg553sXNiFsuAg2ta5nub
TD95S+xt71/pVgq8/C+bScPdVNqgsoaE0azoVXdLLp60sN+29BOdc/Exw56G7+91DMeJnn+fy58G
5KqBHvRMpnV50HVR4Fcy92217NtW8HsfDOZxBoFOIahvd1vI3/rRlc9bJY/N0Vq+vRG9F+e6COS9
J2ixoPY1IJZvCZ4TDchr70GuJMvIl7gqOK4aIrGNQLXFTGGCyeUN6X/vti4CN/7awHZ36GlZbwMf
sYmQ/GK1S/SIro9QJSZXr8GedAi0CKBYKRvMiNVpcwx0xOGkQW6+nYU3Rg9ZaazuU0VShrruT7fw
Q4Caj6EvulWXjPrIwbz33p3EVNHbkB4YhkqbZBGLvqhA+iBYudcA+BaouToj31/FTtb73mmZsith
GckEtLrOlAKO6eSmfpDsbgn1O98ZHDdoeApHja6s7CCdw2L/sRkSaTev5pBKJI+/M/FoGZrAGmTe
yMTFxj5gKMf7l81qvF7pfdl9RzLm1/3zLAJ0kZ1rT2+r9+bRW2UtJP/4leifsLIPy3LaEWtlqmvr
/9377HFQcSnek3JeIXdnz5k6D4W6BzFsT9CFbfBHw6mrjis0MaF/mPV2rQXQGyD1g5l2KayTgiqF
TY8G69In7cuPWreiN54u7VhR35TLg4ZBdBBd/fuc4hstYBPWFJ71dXJMI51t1V3QXRDMHaVBVxV3
O4rZd0EqVyAiORYHFhbmwSIBL7fZfrBAiKjSQU/8kLdkQE3voMbjN66yizYwuwEhW8MDj4hZuLf5
FC4fIzYw7aYI7dG5piW8ILXN+ZQYmYF3ZmAa2T6eTzGFvG9ipTORJkJ6cjAl0VS0eAORKSnCAc9U
uyqVze+HZggorlVoPNO1mdzoRfp1bNBUatNlewKqM+C+3rGQQWlui41ytlvJFGweMnkkH9oLhbCq
nhVPta3JdBe3aakZVlrOFNoCV/4ml/MQSN32egCkh2F1IflZ9iNKvuEVeprnR+9tOK5M5zBD1O9Y
HNh8t9rmyS9uBM+nLUz9EzHRsFmEchu+Mcrjm/1wfqmmmc60v7b50zASV8HHJXbchgCHehhmt4it
a/yYB4NF4Qpj1ZIf4nT87zAYrkwRAEZdp/EBoxDfqFffcbHPUUKWFILekKr8KhSLLinoVtnq1x3z
87cD/U9D2nUC9J4VQOB5Da4ALfMok8laz5MENXkcTwILbozA4GfCuNQkf1UN5HpOUTJabBA4ytWr
RoSNQb94a6t1UqaKNH04sqA41eebpQM2ifwKqD8Gs7o0qiFdDL/I6IuhiBhrQefi+lc5jexPexCi
nxTRSfTezoz2/u9qfSW3J8y6Fya4BPWBQ5fQp+vMpZrJP6QJPa6pZ3Ld9LfkgZZULHjA9OxsEKwe
TdISE+LJm3ti7qQVNfCGX4K45PnsywB/Lp8g4Sc/HbzYHwuGCmwXww7N7xoSIbvuvtuq+9d1Z9ZS
nF1/Qs1+qjdwEFNppRXFb2u/Naj/kXEUh0NgoDP09hLsf+xRFZLIWlN1+9fv5azHMwYAIpOPRhL9
INbP9lgOKjtj2H6DT9uxjPfJSrRLWoZgxYQ0gY6h94NEjtzNENo4/H2UKF5kTOZREJFhFV1YGgqr
lb2iqyyOMv5XqERsoSJr0kzKvNgTIZ5N+93ujgRLqJ3WYC+9KKtPucXrYBSCz6VhrNoG6PQW0aWp
t9FFBRTlgOwiErehJwxTPKNXDW7aVfopQohDJWNszSFmfLQ1ihcB+DtW1APiUdC/bp7IAT8eBDZJ
krFYwMo6x7r8zQhDrHRYu5pl9SUD86x3lPfu0C4idbjUuQ1tVh7d5qTRTVuCJp+Vpb+g/PWFTs/Y
FgmclDZfDdIsG0MIWFoBZ5lLeMqRZATZFuu2BcWgl8rEgVL3kzkipv+QevN8EbK8fyOLpJfoCA9w
/L2od6wfViUdbxcSJhQc6yqrh3F8lWNakMaXILTD9/aCQrg8pA6e2Pd+CC2nNqTGipHl6Re/d++h
lhd3UA+70Jr7o3NRNj6ra/5x3ROdvpyoh7RE6b3/VXazi+w6aMdGxJ1we73RaEyk9PXK8SusEFwk
YuXSU//65RetIbIYreL0KcnHZGnYcw+qpwe9pOXIRyMK07/l9LhkXHR0iJ6JYVwtiOIYW7m8ldFo
ACqRhsj8bbc8r2vVZbQnc/I6QUvlQCuve5c9xWkM5F9WKMKhf2TiqvjF8Gs6q3qmKacpmNkF7Smc
vX4RixK8U+LaEmtxhzl1/b4Nhu/f552s4Doe74NQsZkzqkmuCkT5tMnOISoKV/9gmN2oJeLYozYs
KNup/qnhVoXhp68X+kECAaSFXILXJP8/sh3dFq8BvYKFbaEO8In3Cz4x0ylvBPagzlt8Ayed4w+a
bsr1tx01tIhjEmwnqLp3zFkH9DQU6XRomJdMRCTvWX35k+8I9GuwxqBRcENWkdauWGVbDvLBLmeZ
lQ6uk+7l20ojfe+q+MgJOunSI8Y3uUtsHB4tmAOpWcQv79X8+mtlcXzzGBUPyNVtTzC582vJ0tvC
ntAQBIMxugiDxFYXrVoeCWQiDjaGdDHzTq9FG8Jc2D29iOvJNmNQjrB6C7kJexM+Vv66LhH/6LwY
i13PiG7a3+0BpSRNhWYAXpG7mUqm8i6sXsbglu1fYMrybNekppEr7BA8F0yGGPk3PAdyiQZ1SOBV
bJsCPwCf8HWKsLnLQiONgb4XBpHeNOx3gQ4P55Img7vt0LC/CscmJxvd80XCff/wjnhIIo0YrLcR
efvFxfkuVwSsJk7zs9I+TjkmGnkA3D8pAmMK93sOp5pAgN4dP0gKdGuCkbWlBp/amsqV+T++W1Hl
f3Om1VYuVg6LRJhGQx1wK95XnjNhBYDr1759GFOopYeWp/4NzKS9JBy5C29kGuVOsz/hsEb7BypC
zYOGEok7QoEWNxaY6/Lpu+FDGKiBj9ttcZa7CZ0TiH9242OVggYbFme8Adg5pGN1xymLyPI3j2+7
0BrdnBQOh8j5VrE1DNV+JErNqqU9CvBxpbCzl5j4ssMxNJZVD8Y7zrAoo1gPl1Kqds8vQVfJwOUz
dfuyaQI505qul21oagnZnXEiRLudqOqBjwcivozm40GJFtXQ7+XuHx+Q4Djk9gC5LgsIS24xFBAZ
Ca6L37+WO3G7fYrxe4lJJF6DBjsLvwsCSObgVZw5LvsjJyuIWClampMUaRwv2cKlUc1NINInbDuc
jIkNVCMFLxydA+RM6KEgS3+OLr52GNw2DUaBek/C3gVBQT3JLC008oHCO9H1BcKrHP1ykZEePehy
cZPIpQEAb69IxuMAfpo+I2Vf90ZVUVnipa1+8aj36SzpoFTK4dUpn5DRsTgzpImOq9V301gaO761
EoBiGz/RRiRrtYZxl5ieNCAD4WfAD0p2QV0o5HT4oF5uJFXlZf8JYyBNoS0ekWoAMUyboY2YNOnX
NJAmyqAjQ6YtN6qv3c+Gbur+FiE21+xUWTLI7WY1TRM6RGXBCAGRjINkw61nG0t7+f9kJkPudjfp
Wvxbh7P1FEMQl6wKo1HEChHhZRMd76E5EDD82ltxWQyQIYz+oN6whhGbPsAXshy0Qk1v+hgQPdtQ
Vc+VkkB9waHaMEK5CEpXLX1XWtzDTHnZKfIuIUrnUkYL/0kt58Ntuw4X7hggxccMuUFaD5NyA4Wk
6fVH2tu3s5Uv3nLc2K8DmPDuL9tEBlKOVy+5yFhx+hXs8r/DJP4vKg0PhIuS9itZUSHYfuBfTLBY
xb/sj24LVvoLu3YIsbURl4jD8NNZ5Ws/c/4HKCzzRFkgFfebiT3T9L7RjPkX4C/CfDESiP6vfjjk
qdHCe9ujilYh0FOSl6KPT/FUP9GWxcaMBvX6xwV7rlt+7xVAqkLZRPkwk5U+jAunJLJiSdA22ddy
2wb/muG0S5Py0BVi2b7C+XeVgNZtig32rj9mzeiQbtGG1SRPnXm/ad9k3VWzsbWVIH2LzE8SR9Fu
sk2BCakH2jpqG2kcd9FOddl7I6Qx7vk/xSzh69mk6UDpa+MAddhytnNLUpI9JGeE5rzX0uFsJsdL
vGfpKmPiCI5iY5gmqCxJskSlpFSyiNgrT8gee1xTphzwQUvgrHiATWGHhgwLzz/roDoEc/0H7P+o
CbZQx5nBZd418i4BHO8vxSCT4/O7QODFRhOlhRFayldrLPDpa68pmbFvZy7AR2xY47W68ndpadjb
PbMSyjT7Vr7pNzgESLmeORcSOiljE3niDGRC6UzACO1nbjlMA3BDTBaXOzPtXKPiZoxekpDF0A4X
/yDA4Ph4tnYdIV64S8Nqy3Q04FN3iMFcsmTnBsyb1V1seiUy2zxsmxu/isyIsBFuPCt4xRjoKCWR
fw/z0cW5kS1h5R3d2ZAULB8zf8ldiGKPMuegnXZFrpwWU4o5GTBnQwh//Ic9QYWjJAB6/LV1nJ3h
rF0MxkBNpFXyc5wvWAZMLn5T/eistxWiGT04StAOeKnZqVtOcyVlV/R+oc/EucoHPF7KgEfElhUs
2t2ht88pUl2m4M5Jfil5QOTLh4ry2KeWcoUA89eUZY7RKrHVeZJQDmVTEDwWh3Dufk6KZldl0L7h
0GakVQGX4VSyFGhqsaYYbofTBwhidHAL26H5luFKdPdT4OXd0pBAnc1YY8ViySXdTA8rv8CtFzRF
bEW41bza1MMEP2LvOWX73QJdsxdcWGqvjXKVAIoadrp7Vxp3eVNX7W8PFWLTi5c1lr2Vos3bNAtt
3ya9ZL4UOqXhQZkzM227bim6MiKW0dA9OcDdXhZQGfP+zQHhsI2E8AE/4irFaTH1/zOeHspLEiyY
SpRfZqQWu2MXsRjFP72zmmWtuIDHmqcE80mDBwEMkWrnUrZFLwttDL3BS1J1FfFX3ALoTSGcL+cW
E4Ygyt1+8cShcWcud85rEhWXuWH7R+Bflcyk1Bx0jxqT3lMcFQ2VxqhRVcjCnlzry8KL4YxU6y5N
qtBSQ5qKwUqzfpZctsaK8BvURLn6z0neo2O+P2RB7IxjBaix3yGtT8C4Jhi/LL8aS10kxvD/WDRt
dGezeTbQbSFFeEqCPHwb0kZYiP48pXO/Q6HbT6TPynTw9vsvOclzUsgv0Os4xYkVHdq9Fp4zS3tz
OryyySs0wDELyQHZWlHyxnm6PHTdpkfjABHRKxAJSWKnQhDFzOeWH1UUot4f6qR2am4OHRzeekVE
isGiI+PENhuFi6k+3sGBd194471Zn8mVPUSi+wLT2f8OKn57TY/5O5sbO5Ufq0wO00JsFTy5Af9b
9yRvZkr2CH1e7LQTmZuY14fEPv6LWuNcu/iqPZOoDTeW71diMJfVb88Jz5FbPD+AxZL04nl9Vl2Q
ReQl44OzsTcJ4G8SR+GVLLR8mCC2Z2M1odMcJg+ugY1brp3CBP06aRoENbyi2YmrIEOpRYI2ys2V
YxM410NwXE6BGCI6BzzWlZngbU+AxOWfh9HpqT7N1bgyksRC28VlmSpWhV+rihjXfyQPnUPUMnfk
OB3cqjIz/S+xN/e87ADzLQ2KMtp6OXDPSjwmt3HT/LkJOBhi0H6wu2SJ3lJ34m4qMZSSHZuF6dMA
6BFfZO1KCMQlj2CWdg0cRzWh1AFbdXJN5cwtIC67TZ4zvmNG2t6Rh8gdrqaNMuV+FCpOTAuIrw5U
0kRH9lcbQPRCedZMmrZ9R5iTzWpu31RP8kAa9FopxwiuWIvADfitDunmcQvAwda5O4yUnUSqU5M+
ZB1OJ+hwYTF4PM1rMTWi3Xl3kN6FZitHN8SkD9b1gtUAaJLEOrzlwa0/cRiGysjOuBr2pPzLSvVL
Nq7B7tjA6aVk5sBfI/J2XB1VhRqD0P4ef5RkKGBTNS4Z4IbVkrmbAN5RkRVAjbR1jH1uzMvif1Ns
77bpa2Tm0a1YkcL3sxPXfsdU8hCQXVtz+yp11RH4eqzYIjf4ea4WZT+AX8gMDemfcSrhmP3ZvuDl
plg0Ivr4nmOjqAc/XMRJIBPwlr8UjtlrM3m+srLZHWUO/wFKeLsXKBX8mHOGrbKlo/pmUa0q2HBW
Yakp46gKmXASW8fZC/Mj/7nWQAIMpS1qUwPA+yJKUfgbKu7LpW8x2hCLLRh9Rhdith3xdReAZb7R
m0qABRwwKVkZwfa0gW3lBWU9FZ0GliVBNsmCjSvTr/aR4FVD8+sZQdZHM+LCsP8txhetR860NNHr
TInfSkzyfBMENf4eErVLxRvmABCPyWVDbHQaLh7R3mNHVUS6id2UTnFvfJpt5Gy1YIztBMSxnYsf
WN2A2fTPAqe9O8RF8VDJdLmH7Zc3uG5SR+f8Cd5h1Q1yGHF24MC4aEk6Eo1CeeU69gZcbkXFaMUg
mSPGpvZxDLd25ePyERxgW2EU+wjuD3m4hfCgoI8Lt3tLeGc95Z+RKqU8MvgG2zKBHxLdBM8flOYy
q38OAr9MXwGVXvnlJLVlHgTBXkt2+44h1p4mjtrvUV1utUfBLXynKM+DMW+9NNzg63pVNeeatvQy
rVIiwqKUY6fnfgYb9B4JvZ77116boBiOVP+XUZjSoGNKMFfntUD6e+oUxt5Rwwn6gLA5jp23dZ6Y
St/LnyFkYM06vVEiEnsIrww/AtpXjpEsxvv2Xjk34J5NA8s7ZmoLP0qn+w6kmmG3+zgFFuKtmxAK
dfIDMQdWGnY7ryH61nCBAks56IYiguYVpXH1DA1aRijubKH8aXg7OMm6GZ3udn7Vh6fliVH3FMqd
923W9MO7Zu3O0Olw89S6Qht7y6ObL16gGoh+6U91drZp3bZFmLuNxBEJr6uQelcuYpcr04csCxHi
VQARuXGRMXMsbL1+6HW/uBnAhWdOC9Cji0PreN2vgTSoDFg56JVTkyY4zI0zhe+mLZjz1laH7oJP
lgmE9IGPHHOz44H9IPg2PqGD8eCdb7/VWXiIYN6TRWlnpbNCMn+CofgraYtORKPNezmz2yuOdpCO
S+Kfm3llspCBy530Yxhg2/fyzgvPSDheOKWDRpIbeGr8oU/I9/Pnag4V1gXoZcj52KfEaG8lL5MM
BMFNBjBXYhOdruFQkyodK3KFmeVdYKUmJUH+iHWGhdP3Kyeu0ikLljajG5UXAOgru8x7UyGjYB3B
/sPC1JwkHqHP8dSkLEfo06ozKK2t/Ixqz5FntM7WPaiMAYPvYcg6wh7dNsdab1Zvh862TzJMqBgp
yQB3AwmE+LCpPi/7X/RAFy/hKhjeFthAhy2FeiI1hpSCvs3uaKHJ8kqP0MOiXDIRrCKowEBYkXjg
43HPRMx7rjD78R2MakZus4NNTbR5Q6MSVCT4eauUKjPFlt/DMLSTgUfo9z3ouyvx5GMkVqPFt8AM
7BcJRUDp0kBXR9Xfdgg+L0lDJhy0v28ejhQckA97f88AKcKnZnR6dsws8XprEpCkmX1qPY+/tXQZ
HSlH7dg72zQVQKFcOGlqcxhfJLNHtyak0TWGn6bl15o/wfx3rrvQFC8Wkk8NS51AI3kS6wMzHiPh
/uU+3BP3r8Mjxt3TJmBOrXcDh1WxjV0WPoKxcQFUYTk/QF7R0Sy+Cq8LED9AHcAseAlmj6kSITkB
cNhAzOBA0+AL9g/DfN9LJMqtTw1C7sbT5+i1YaXj01zrav1h72UPV0/cHdFoS+M3c6z2P4k/Vfpj
KT8vnRKt3FCMu9CpqBvdwtredTiV20rOnSEnlQ+TC4qcFsQlAcWTf7oFDhq/ylK5ELxNsfTiTI1e
ErG96lH7IBMcYMsybv0LIHEUbioDCr4tZMBcekuNJLornAdrHMltCV7qzf+ehmJ/zOVaP1hU/DER
VSxbC4lxxU76AIguuxV8Iyst6HlQavA4y+EmBKchFvna/aJFfuKbkMX7TPbLpaKOjVqknFSKUKK2
TkWNlpMvnlB1uW633ZcvfcQ/DKYZ4/BW9YDNTAF3y/21srrbB2vkN1k0mUSpp+/Kdq8B16v3+0+7
2IFRZSMD+aY/DLHdgOupQ1iy+CrJKmuvFDD/DZONvNVAzIVdjm/i+oemGjFHvnEhV1QjZBSuMp90
vtchNxN1Tnwf4Chd9WZvQNv8+71rQXXFGooS9BKl4wVs7L8V2ofw3GSplW++wTxrWgFdSopGrWf1
M2AchVwAmKrZTY/yjs09IZ1nFl4AggKb79CtbF79gnLqnuOywH6/reNNhGb6LZ1EE3jMyjGFn6tO
sbnu7tE3H2eN+AXuDiWNSzhBSl6YEoR4KrUd1rhUJbtiq658CCPAGbbxhjGqQE6ElbQg2JGgRcX3
W0I8OxGUXmSUoqq+c8KDHBpodApdiWs7bpWQCCWa80TOuoBI7ZZM1FzOV3M91CtwcZtR75ghcbXM
F10GoNK9Lw0K9QRApDinJ9i8m/ufBPhQdiJRiptevzHg56ZpGB0KfK6hOsnz0DgfquqtLgBP9V1K
99Tu23XGo9WEwpKJgiK9qqdZ3rMq8sFK2uDd+daayD6mSiD5riCDwAMvxOPFneHOHB8myjkEL37N
EUIxrJlFR+FRv2yChNdEkyAL2PjoMZ1t7n2Gdy8jIRCvt/fVsYQMhVRkQMvRyAAaD61BKuOAFaOP
FnWM+xCi6JmFnGdU8++tSVFkrl9ubLJqEi9eVvuq/QzaSbUPb9462yOo5uSgAzkgIHRNW85pGNB9
o9B7ZAFH7SNvo9YNFRFUiCr0DhJsrq9fn26TYgQ6bCZ1Cf9n6iKQ3z0X4uStuHhJGDAa+EOA4zry
tA/HS5GhUoKfR/NJAPn6QCkO+dzopzGxvqAY9yFMuDU4PPExdKT7Ou2oa+blpDpIoXUiEb23HivY
tNyeObWtbOJosTNblcuRSVBfVhCJCvtBFJjY7s6+IIB7sE1qJPoa1Bfd3Y6ywF1rn7VypM5Vc4zg
k0UWvJz1kWlc+WpcaDzpyABG1rmP1TypU++cpaY9fFmIYBYReeuFiPXHW3knB8JB24k3h0EGq6KY
sQgGFaSaIUAz7EbUhuEHJNnkt8ZNtb3mA0l9RSA3CqNN8Cfhd6COmh1Xs/190bTt+P21du4iQSop
jPvB5RGsy+R2PgYhWhnJtWbt4oMAsg6DkDmM7Ob8HVjnWFc142Ucvx2GHpLDW3ekSkg8kJJzj+M2
k7Spb2r/qdQPMmn/+sH2SB5HUJAzgmhehb/bfXmciYZZal20TEIsZjo4PMdsB/IHCLINUziEReZO
qjIe5VRheSsYGsvBsYsNFp9T4K1DiNSIpz6qnw/Nqlq3lzbRp6DswmbJzb2MoFoRaXBrEHkKQp8r
LM2D0QgOuL+o+EdF71XsXqwC8+pG0+F1Kf+JP2cidQDA6XhV6N1XMHJ2y9Bv22oEtJxIHL+lr5Hf
u02W6xu2wfVmwc7ObJeByDdQhd1V2WWprYAQOCgYj9t6h7GrYzoGMEI9LXniY56krBIGm/5ialBp
zP2ZKWk+HQDX46er7sz+D2CpM3xcL2w41YB8/HtujIWO+2vuKTYxgjDkrV0KxlUV/KF6AJf+Xiax
2QEyrwU1req3ZZgj5NlT89utFNSPy1X0LM26fH823XFIZeI27ez9nU5vt0l/0FmDUI7spwt2kuJ+
A9x8/c8TFuZhATXrPKnAdgoh5w3hc1FS6KXvRrAxfA2nZ9z/WCPLGdUnJqh/tt70ghGfKIc5MdYm
SLN73xUnHjBsDuj6M0zWONzPDq/HtBh9fCs5cfSJyHDaVYQ7xD8Lv8UPLVkdFWZbqIRmNjRwsfSX
RHzPrP7tINq//H4SJ85aP2QZ8ixFvXoVSZxiCGmm7KEbXdMueXWsPHUv0tMRhimeYgkD0KaiALWp
jkYYQhWtQJ9+RA/0UzmTVAou9FC6WUDiDC8UlbUkfcQ5+0CB/Ta4Q6h0NoIDkL7f8yNgQoG5zOku
sPAgvmi0DdlLWwwmg0A61dKgdPIKQfJPMaR6ZhQ6Q6W/5OUlH3A66WWJ1j7AfQgpbOiE9m7Pkqer
VYkMeOfyKzbVmoK+GXiACTKpd0xfxhN6F78fxM7evGA5RfON5KWpnf34iVy823OdtsghkICLma+R
eY0sB+efIDxZ5NWPg7WYVq+jVxZQWJx4g3KjqZt95AW9IHcbdtoEb88Qu6whXHlgWfuORcAAbRnP
OJMeQNQuKHgk+jm5Hj6JeBzi4V9DzEPsNjviW6XNExDyqSY22m6lB/ny0qJhj8iZRbt/ensurskL
4sNzmmWOC9/KaHIyhLCmuTVzM/X280wN/sFsUNKXboe4lQWqilwZZeTOj6x2QxYURbED0FZgAXeZ
Y92pUDHAZX8bf9FrSKGEcJxKuEkTIq2SNTLARRJ+/9i5xeXLlQQbzJpbCsGv2OthWNeWZa+fjA+P
URoaCPh50slktpk2HPgl/vNgMUQgKpfHgTJ9PWArA7WFFhMNn5szb38rq83rGSOqgLNOAUY0gwp/
3M+B+lxHZNhYFlQ72TsSm+DER57NKDPywmLUWUg8mem1lO+y73k3SlbuUcoxMWRXcnou4q+zhsfI
1qmUXSiNungKDZD0hOlE9Ekk5vcOBAcW+ogu6DpcCiAtUXg5RLUgQgy8CCuYvWEpzwyoR7Acc8i/
CNJ8c8XBYvLXaKXFe9h2RG6HvLlnq3b8E6yMaHZ/HKXle4K87VRwR0L89DLt4sByIqTAqw17U+T1
tYBovT2A7lyNUED6hT3vjl3TRhgumfzZjsIQEXyVzcZ/wRV911ueCwnXnH5wigN+ZyPKO/mr+i1P
t2Izkh3w0hWeIYAzVeU3yEA7yXwEz2BcZrnRWBF7K2ZjCkf7CfOhjW2odpQ9LD9EUomfFlnkNl7o
ILsiCqti5dWneNsrTs1GmsIvF3qkkMJRERCGKIz3u7uNwNfBe8NKUBcpXbnjXd6I7mEgXvgfoU1q
X0fRkyCBVmdJhzT/0eVYjNob5szWdEynjwHtREh0iBCMd0opms89mAvWvj4k4+WDpgm05nPLVSRr
5MFso26OcYXggmA3pq9CRwjEOCS/abf4l1RxRRnrevlkjE4pZXwLGBbHR5qtr6MR6Bdk3fRRjC9u
0lHiMdPeC56BdIWt10l/fsnfmteQAuSIQ24XhogylZ9hz3ffw3p0nqO2Kd6nz6vgdE/aZmQLrWQe
O2rVXHflokWsFa3uqhh5BEE2MrGIpAvUkWQozqDUVBvSatlQGZDa2xp9+tlS5JGCmXw8zR9A2xHQ
K1ZcTzN2NdLewUSnk9EFnmrduPCi5CsU12zn1i15HK32n+JEJ4OUMMjDmraL9ZIUiuX5DU86MrU4
JoBYI1KmpT0dR26iWYTvmwYp7jnlWD7+UBVkWLd1/vAa6TDDxL+9j+Cg2oRucjNkQMimaz35/zH8
dbE6MybTZ/YHM6uju+M2O1q1NtChT/173JPwTrbmuMboHX6CDXYA6Gtp5RI7lydOVERlttHpM8V3
UF34RXKsFM0SZMa2JKTuiggHSTFknYXEbyMrlAMLrMycWIzoBH9h0ysh0vwnTbAsgRNyXiZE7K/v
67JSpJshO9+ybnbkoI6Ir9ogGPR5opeK0cj5U0FM01E6px9GzqIGznx8MVlU4mIFgzXpoGI2T1Wj
CCBLf9bfgMVfur2MlCGt5xZyPuaslGV0Zj68HUY5b9F60C0ZXDR52fu+4aAms64Wz2u74iL/KUvR
LNFkqI7AfwonxZPRru8AW73JeOHHc0rdnoKlJqzpKS5brogwTUz+ercML+NWYPzWt01T3S6pe+LS
h7LM0nJ9CyIz3OULCDY/U4K+86Jw9ySXrePUqxW1CP4EiDosv4ey8w3Hw69EcS4WUlAHP6RBj1H1
hxvjxq7aOptSjTo1lxmS2tcsYL3VO7JNT6leBPKW3GepATZGu7V2GQoGJwgcXsWR9JtJJ3aAapY9
bee73RCFY4vKnU9QD2mOVOOybnqTDTuJAb40EQxiqr5VfMcnbTujdpung3OBKkw7h654Nqs9ygOk
lxRv8JSt+JagAw7np908x14yzujLaGYSfTQ42Mf0FPCMiWz6/wdKOgnvcoABdWN5Q28/ahd6qzfk
FUoSNXA+fqEhEkG0WHXqRE+7XXylQx6Y1jA+M5k3hzS2u+WpU4pviaaBbQ+EfodeyQnoQbT9fwfd
BPtkX6VnRAALOb+HNh9SldCE7mlEmYw1Sm3ZQYJ4+h2QivO941d5Q5J684KHgU6Z0KweU6b5v/g0
E/9JIP7Ztu6ZK/ezJ0ZxcUWa1nK6SIBRUYSC3ivf49A1RHjYLQaASYnxm4TmwsIvCCDjl7hnF29H
nO6ugzcb/z/zWmrvLGpJn/IkrJx7W06LB8N9f/0L+MDtM4NZbgNR6Gw9vowt0AUHNoGg6eW9OQ7e
YPSGmOhRHRjkt/rjSX3GFYY0Eev9NeDLvf+N3MNLHnhT0B/X2cYOqnReBlKfS5j2U6g9ULeWpzF2
i/gJ40K/dLfPr/8o70Vi+PibeEDsRcFUl9lOK+yqYsRHTgXGu4WU9tDR7FAncC6mI4fbaPItJkA2
XI0FkO3aQc7Lbglo0qsRDww8yWHgrQ7vIvrnNtEWozx8FTy160KqiD7GoBAJnLh0cjT6cam0W1OF
BOfLT9evubiheoHgU9zOLacNeQ09oqR3ZOWqvEYDrgPdUoLYfuiA1spXMALSypmPX5e6sjRs42nz
J1Ln/DKo856F5prP4Hzqk/yjjZzZkCOxXcpYuN7Rlik9UjtXvt23jA4m4uoqeeTJXcZyS8p1jiTb
kfE2H2MmIEdYeF0V2YnVPjQRvees4Laxw/ynIwAruS1Qu6IppCofS3696kCZpkNugMHAbEqpADtm
FSYyNvN4PixE1HgmTrdBSbs1AOjhpobkEkdn6TfauGS/f1A/dDrR6AJ5eM8Kypg4TjtisvNdtvTh
rb49L71+e3v1gaCxHl+rgj6IDbSwRxS3ZlaVdZj7w5OcZbofa3yNm45ibujhJyV3fIsASRTFDMlz
EyZlTdfeZtR3ddinWRi2Vm2K2P9HOgaWnYoKGTK7ixEm+GKu+AO9WGydONdHy+oVU8KmDrq+nBSt
eSWycFlVxKitmSZwY0jvx4c/Z5q024Pt9DtNTEyIfc/BAO9zf10SLt2iFR09ZodvqOchMMbWJZub
pw2HCtmGLM08LZl+EDFO659pJMQbx/y93WKi+dWJVMlpqXtYuto6hQYVI+P1GMNB2d9FXR3DFSyi
PR0ohXHHGmdJKBBvN5gdCxf+PPIwExaoQUjj9KWRgjnb95HCiErWO0dQWKuD4kgiAGRYzQxkTCSV
YE6xRWcaWElKFaYfbTm5p3IYbDN8vBnY4yUwYazjePXSP5XGPKOjITswPk++srFqQlx3HsCx7Rm4
EzagIoI6CiCnhLCZJNdmxkHr50TVskV6Xqy2qL3h8TF+vX6CwZTBnVj/DDt6clNJuyrHbx5kMank
+OltjT0YIf170DnYMMBZiG7Zm4/vbKPebNoSPkaDBbEVTnE26vitQv3GAfcTBjPGgR2m7qGgxpwS
lBd8I2cRLnvSkcsIFN4DTHS5EYpjSIFGoSScY2TtmTLc/nNVm4ynvCgsas6PpOmSF4rhVb6ArP4h
pAJMqmwyjiDl2NSi8VXKSQgn/7KstKBqfu6covBp7p6dXURdZ1sLML6pxUyS/s8c8/FC8zToliyH
TuC3Sy3T5SMFZwq8VQJpv5T+F+aTnMufBTvCn+kKw9qqxq/US1XLxHIqQEtHhLmIzf2qrwORR2gs
QYiq8IqrhjvYiWZIcrocj+zUkNb51WKJqkxUmCaGFLslxiJO2KAJt8FsuzXKwC82dGpDdWBB7cBy
NL1Wurp7yXAl0UCd6S8VnjGlwVGHcWaiQe4ANjjR9Lua/kZs9vqvpzHROd6y+CIPrkJVXJPw3odW
18dXTjMTh8Fb46w4rVgoQOu14Huo6758DAgZBX+L9Rex5NoyY2atuD9UxtNunmCmU1BGqhIBsdlq
oaVOCO3yk7SkG27m4Pqv08wlGI6YgUHZchHcRUoleQVmUAf7QliAtkIen4d7vt1N0Wryhq267X9B
YLiiHYtjKnXStn4Kw1YTCqQUyzcPYqIZnA2ppQSO6CIwtlPvhIXGFGiPvt0rZSWejoTuVtGicG4c
d+zJSLsW++lmhVE1vem/Eib7IymrRWreqNB17TI7JyBQUSRbVgUZlCfDmK+rglcEyz+rD7+08qxM
nCL7nxySV9TXs90O9XBudGSMSSgJ0CNnRtRCshMqJvkCjgs9fgH8n4MHDWB2MgMoqOKuLDRIBf2K
XGPnSAmnGgctKpy0QOSXUxH+fs3NNQUFdBpBH150vrMWjZU9DEpIPABsxInA7ji61Y79j/1yY3FK
eql4UCoazOu3rsZx+vRWeJ6RxywCEajFgCr7mGYvt0GEWvSHQLc+Z+m1GhMTM041ARss4R4oVfiV
A1ndOGVmWRAbQBzatCPbYG7C9StMtYnV8kE/l1FObz1hytCowqTtLkdvN/1a++RYizGdxl8tAS9E
KnATxc3xpkSp0qrkuKCk/4DwLJiNjqvSztncgTfMjLRdzqviXHzxtKGoQq9+Ed0g1ihCkVwfEYhR
1jAm5Z/P1g5kXiCv5VolQmLO0yD42qrbUy5XPz6dBxwEJGF1L2M4jyZlgBUzXun1+qIKb43LXqZi
tHQfVZGSHjwPh3dn5jybE24kai4YZ5Mk+HTfl92r+MCRF6f2M/kxKH8luPfTUoLudUEpxupU0roG
hqNZHebGk5NVpfyQQOHRaOf+Yffmo9VEy2fXh7qnt5MyGdjvs8iU8qYrA2hr+67Gom4IarqTrAYG
YiDBPCLYHEuaZQlGvMzSFrZ6BGsffGLfeyB9e0Tls4plPDg3/AU5KJ4Ix1QwLPoxrLMHI1WGiWL6
U3nJKwHIuci+kOLrcjH9Jz15JzsiIT5IMif8ClxEFe0nCsAPYSIknxjLv2Ia5r/V05DfcGUgh0ko
/WQG0ChjCwxP320DQRWHaSbDZGdlu9ruRtTMAUxItJrTrFZ0e2+HCGQhZOfB31/412lgfeSIB9Xb
z5oeczVdPxTO7HZ8BzMCT29L51iaJV6x8/8IXalK2gE8QZAZfwercNKoASxWhnhFBJBe3MPVNgoN
2XMGcU79Vom+p0o1WbvtYlX/SdMhHHzWQ8CHnJ5bji/W6tbeCT+wqX6e5ZIoE1khK0psg9FCZM1u
LPZwwDundCBM3oRLYrDLnOdq2WLBDSriT6a6Uf470arFpFO0kZ0UpdxahUaYnfIXqFPK8xS60foK
q2eBTbSe6g8BIjuuYy/HjCqdJd82qTrxL0073LezKXCzM/CqVpEpFEVj9r6DT/P/R7WHfOgcyvkS
FAXhqf+IsMwrY1xqLD0CkdZ+BCu4SfFFPTtV43kayr39QrrwA3SIPlhHgXmS7KzgTQWwyiGhRheZ
dBe5HsM9krl3vt1zYNFpP/Fv3R61WGTuHe/I1D5Z7GzutQ6yfp6baFzOFCKDKWbZXCCj2zSdDMBK
sn4C9yjkjY4waDfXVf8uNj+/esSJ65B9lD5fdmYnFKS7a3Gs9/snmHA5+HLJ2GZD9EsDZ2Vv/2B6
IlE5jMNv3Jh3ALyDBKmVhq1VALJOPYsPkZ4eJ9AiMaqTg+yKhdKsT+3HasDhfDpjk58zLGTJNCa2
1IWIzU/gRuuDZYpmezmumAv6zAW7OBWoYWGe7ytL6mNzCXdZr3qQsygVpodgoaFLbQq267QycEqm
0eF+nay+QQ7s7r4fuh/3NeTS+w+Z/M8IN957B7P8fOVgT9pw7eHeQFmCWagixYJWcH3UMYHc6/Jn
FLSCTrtYwi9SXAvzl72OYOM+2+hw1XYda/qHlXW6UNeXY6dNFZhn/Ez4b7PqlzZRjMdeKuwPPSbg
0uP1rUFwLGqRcpslcMIw7sdEu+6xVi5n74oBGEb5Mtkc99Is4w8gnZ7b6pMDUgzwo1+7vpzleXk+
vylgDgjkSqWe+/oAirnV37ZLPPCDZW6Cts6Ll7TpdwOckV1b/fsnpI6XVroQtnffHdbLDNvxiiMX
4ktKlHPo0Yxej0hOZreUnCsLV0jB5LqaESwVuCPtbE0DHLszQrrZyBYtUffIkKe90BljoFh+b41o
KyeYu8FaL3v4l9hYEFF6sKpMMlmjI9ZmCb6rxEL1oe/+jjM2GhxjOrX4PfzBkuBPnoNNkC7xwIVQ
khzY3XC+1Otb9B+FKTMqMp6djlGYAPGzFaIQWHAO0UHfHMCIFZjmz57JJOggVe4+qEHO3ZTyVPgR
oRy7jKnpjImGCIuYlQXdT7jmYwR6/NLvaGI+z1TS9tJR3+1z1SjYxz2ImEQmLBVVIbcP0cIdSCL7
ElZZuSwRZmXacRmQGkS/e4xwGuh0LW6Q8CDwtSpqYJ47L7at34qEYRi9gXX3+pCBRSZQAWdML0fc
RDnuqMl45QkCS6jXgTQxt9Vtl7t7IKMnYmeyPd4DwREeUovoYugJD9owUAkuZ3GHjJCbPcedyvVM
mo4vaDKCA6FumXppMT4tMe4G+8xiaxlwpoDwNtaYBPXYdONJsxQgKb6j0Mf+Vnv6IA1klsbJD+hp
hKbd30HXPK5/ap6VdoDAaZeHbMfaRaYPmqM+h4fIDvqBHB2NhVkHlorY7CaYSyl1IzoVAopoerUo
KSAr+XUEK+Weqshy9gSRQqltyXrqQjA9LywrC7tKop4Ptx1eUd2CXA3Xq1ML5/l5wQAHROFxOuAH
MCMYQTmO2E2l+dBMS13DiqdGT2RVE+n2bcgYyD8HJRcbzXxdt5S/tsMHXO3FzdmfeILpcCsLNRvj
jmrf15IdCJBIuYdjSlYQUZK0Ro45vmp++yQYNwkBdOAvoZi437ghu6mObnksgT9ZlLL6gsUpo4mO
p+dOo4zWvoxH98t+64FFzArTlHiZ9KlkEuAfXfdWuOW0wZ9ssGpWjh5K+WyzYS+Ds4RHvM4yrcs9
Dax9LIX+7cPzCMZLWOHq60c0oa3xiVD1fszA8CI0+5ZK0FaeQ119JzuuLs6nthOtuLii9VTKTr9b
pKktNqeinnUdVU3G1DWOY3hCv98zmcc6M/JE0HPRB3Lk8mEw12vdTL3I9hb22IiFJkx/Pmo6KE1R
N98Fu8curMyP+qh/wi6AFoTNJ7j/civNrpyLBNzrvuii2iZqvyNLXyG4Y+JH4DgYNNklTRxh0clw
fVjLsMFQUUCWYZg5LUOg9gsSxNk1KGrUurq/P0QpEY6IQxHqgA2QoukRqeOPjZbEyXLis+/y0lK9
7AmlvDQfiY824kzdaHFWRfTl+cnKNIM1xjPUl1RhvdhZSyWme5mAX1aC6IJCTmpo4fb59YkaRNk4
RYCOmrPO9K1zy8T+KIPQ8d6OAn+/W2SlS7wW9G5S9HknSrAyaUlhicSmXInFemcvI4WHwb6WvqP6
xyLYEJvZNtEeXtwqfOPdR6HmBapVNpKvQrZ8tY3zILIMmAlx4KiB8DF78K6PFKj2E34TYn4wSSym
wXypdLE/RiYxSRqpnKXQ0NcWKTGS8V8lPUVJSZ2kyDjhegNHkfIlxsU6hJ7tx3dHA2Tuyp8p4zxf
0y7j9ENrtpw0r9DIYIj9C8DECzdu+7PZ6U4lL981+8Maz+4GkQnThmSsKh9KaXODz1QovYuKoZnl
RyibE18Ln+eLjIGW/MV02PlBRVw9s0Q9hW7FuGTl9/4dIyKJ4z7cgSB+LH0C+rk+dKdvZNtsHukL
D+kZsJhKyBuT37nNQFcdVF9f0A/gPlLLbgD7nHN4lOZAutJyy53d7ihcLyxteCPJ33Iv1fNQyTsw
rlkvalRtDABmN9c3SVUg+3JzBU4oi2I7kmODMVqfRXpZ31smHXYaKlM53sciczPCiQtVhJXZV6uo
MjMNy12GOWDYz63bX1i6PAt8IL0G+1KR0D68FtHjWHRxforfKzdPz3EuCgrBfRcZMWTSyMt7fFZH
BuUVEK7VzA0fMs0PcpRq3LNR2fysfKmR5I4mDh74aatjaBOxB/wKy/R+e9vXf+labzhbVG13u/Sm
zJMdwuhncoyKgPbUyZ/Bx9MGqBFoQ6QoML+vmeW0aq59laH0iYdrFuyKhhiX3uf/V33pJZWvSnk1
uj+ji2SAt5BaHf1uE+TPQCnfA2hvorCq2WYZiHGnTqthKyhSyWkRxzKzjIWJJIP6lrjf3qZs419i
N1whfPuLkhbZOEqloRcmxxy+InRm+YSysRUJ//wbeF1H4KdU+UUd+uqmmDUMaDdxmO2akqqb5PyV
vOdCWRR74mxm0NvG1GA2S1QLnuEu02ZLePiql5YL7i4tkpI8ELGLtu5WuadM3eAx+f6FwadcMy9o
IIIayfLvR3wxTp7hBOWqN5kx/ejAuKu3kQRYlCJLqcn6US1EU1D2WwsALF0kXS7hlbNDvIeNaP8x
exVQ4AI6ZOQC5T8Ypufcm/9Mz3xF+KVkabLyPmmYSdqnTeY/eOWAdrCmjrGPNd2gCyClvRKL1Jl7
mgpxytmzqoCUEsm0rNK6vH1fs7jlNevONR9bueV5ran7HMBGUWmtm0BTpWtpV4DGJTRd5nq0XPg6
eFPAyOYJn2kw2+gsvQxcqmnnFF5vy7nX8g1I7f86SAfeUCeK0uaUfVLEj50vUKCD7r7+HBbzQDr4
mewlFdkK9PdciuXk/PpjZTRBhVrgMfWn3jnNOxcyeFUqtNK6J2RUBhPmBWhQ7yDJnhWTj0tVUKwd
/3SxnKN9+UGdOvX1sNSZMIghu38e8eYwhTn7NaPkz2JLxjDDmT+Z0aPrgG0Uu8Qtu9RpFSB200oX
7hG5PBvs0lf/9taTaX67SLgOLxSNLocJJqh5/3KDkS/OS0e3UPSlZkHVpJE6RG/qRgS3JtcZ022Y
EqR08PYEjEeZAi8ud2k/I7nrv99ryd53ktFHVkxJ83WwOZ2n0N13XPuH54oez7EF2iP2Vln7pQia
W+dwz5V0B0WCJbyih+dr9lXTv0I7ErcP6VzScafk8o9kQzCPoMLxf3xs7Mx88qxiNkoBdIta1tWX
S3RAr35hRcI8HtRiCdCDEcHzBZXkNawn9LCAi1/N7WZWrdfVq/6tfIFFpAHLcT7FJZKTu61CjS5p
3Q265blGJGGmL66/6RIayIynCF1KD+S/yz7I0TCT3phlJTC1O1C/Z+g8/16X20LiC+3whWdu48TB
sVDYZVLuKa7nAN+oAF/fhCBF/6KEdpyfnngWlP66D7x+9wR51VQoLLpIBbflTto80NgJSfy/C3hp
+45dZTHiuuyTDByYgcT042f5EGrljQUxiPyEvhO2sCj9aWxiXTAz6UKuffpCTfNXZMYIgPTON52E
Bvenbq3RIE5PQaad7w0S+zW+KHUxbhKXHv4eyEAbN1faqNmIEnps7mlNitrb2d6XobinYk6LLIra
YYzkXXLoitqiCcrLt0v/tBtkanrs3O1NoOGcRDZ5E/94mHOY7v1jQDC99pYnyS/idb4cvqM4E5e4
JcDF0VelrcyR57f4yaWdjpTt+GXykR1jPq6+UmeXDU15xYKf6gZvp+0GsRh2PIvLCFmkt45eeCeT
0WkA6OzuZuTxT3Q6fBNsUQhU3+4ebvw6C/Y2XUE5khNXUJSX1suZo3HEUr17ttTXw0Q1jYXtz9lh
nvYsEFgoATFjk4aLDXbCRMPHA+8OqbjL+i8TqiOV9f0bDUCUEs2HY/Vzgfrx3WUnYaLSaWGeckjb
JKwXNds7v6CHx1hiK6LeVlnIkuUhPUOpXBF3oDkl56H2B0mL5tzDCpR64s4KvnDDglNX3qDlhOIP
E3sWXkozQbV48hlbO3nHvQNsG2Raz6ytDYep6pP/21XVDwN+9I9Ltbxi88e2ezPn14Wcn67U3aEZ
uYgcC08iN8dKQ4gzBPosFfIaKilEYcC5Q/HlWUBoe0XWHzeNbh+vs1hKnPpDXlWLUV52/pAD9MS4
9lY+Qv4Etl/fSfvqLjNGcww8tcrrDk/pX2VbfOUgtDJTW4/ORY5jrYbImnOY1P/CzL7/WEHn95Y+
mFuBfLONok/3fh5n1DNCi+VGlrJeExO68SbynOv6tjXB9q4rBAnI1H4XY8n1II/OyAkr3/zBQxCJ
WxjNTWY/bgcxauO0uajrYbYMNT3UZzeG6fvjI7GIixnF4UvirxNpEVRO/f68/M5haXst+kwvTCsa
Vsb7FMBspO9Lfnglrb3kE+HQXuzprYuSA0D5XdoyzT0HgB2JB3yge98Di5S5tOdPZ9SLFZJiDUpA
O4CwnFciYLsW4xWjaPz0ZiszzUYzWhAKtTWKdsY091M6qFRO3kBOxMIIP5iECy7HkDcVcFaRiaNv
IRMOtjVlmLSYYR4dSgYl94qj+yNvNCh4cfNdsb2K5axxaBdQIrzd7Yj1zfx3Siy/Rd3zEFGXM56z
BfCabI5+32LK201HHUGXKfgQxiLjLjPASIgF+sESmstE3Mlhh5p0EOvFgIcnLQ60/uGjtjbB0KXJ
cTtJhOc/drIGtvGKq1KLbFBgauIxczuRnChPECL+GT6/tEMvY31kWwdgtQKpZ0phxKxzu4nHBrjZ
Hu2hpVV6ZjnCFq7MnfQjw8i3WggBatd3kp8NnhRfHiBEJXV/88u/Q+BA7LtyKuKQd1b0MW64hEa+
61GJKbzvBMdEXMy4RThIpXfPscBAbtByemaS5QNHFw7Baog+nh3OGPZKIk0IkuIZCrWt5hZF1pGu
OQ/Fa03xsw/jKJdJ0qzeBcZocKE6eof9iAuoVYnoAIiAnHbJx0VLCXoB9MpiBAAxE1gOewoIGV8C
5Jv4davcsEYD3huYePHE3w6egTdP3Ihe0kcEqWFjWGt9qpT5Fdoaw2pimGvbjSQLVTkpGl0Kk3xQ
ftI0lLm08wHyDfWINOREIKUsOsUmtr4z5u4NmacWWrpPsYhyHYWltO+BBq5XeHbItZUlmDfwmpif
1zJSkOdw3+RWEYz4vnt4oIgRm8yd61vvS+j45KPDT0NT8QXwB1zhyqw4h8e4cB56SZqkDwV6J6Zd
fbZtUuYb0EPYvbq9v1+AYg9CI7F8l4VuIeVshoyh3CZ6HyoXHbEl84FEdLb/yY7q/PbZh97lc7Hg
CVeQhgP9v6JB7bIazRnKKskeOsXs5Pe7iCub+JPq9c2CPcXIvm5D1r+hKT8UXYBjrCL+RxyJsWLM
6Xx97ouQMWawwhtY4HqWy5xAL7YOKasmJy2SaQ7n6ZUKfqT/kAkKMgx99W8AfT+KreD91BZqFoqa
VhTJj3NGF+Ttdcyb/TNh/sd7oIX0Jl/SZGVVx2K1MsQBOpDBeGbIiL2QfgZxemBPOL/jT4qu13DG
/B2d5PLsJ4jz0ZEVvnwwk3r+E+RtStkhV3EVeA+C8zjospMxOkxOu7idY1fkERqc9YhPTamCuleS
SzEaTRUY0qD6vv2IjxielIBJ11FbkQBwZvSEJlM9U9/MVA8jq9l7OtZUEIH23E6jDneaAIGNk8pS
wtB1Caj1YJkeGkFQa9JNk7spySBZAxml5XAGY2ysWbLCweR56+a4Jy4Aj85u2G+8rnBGKOtzJcSA
WImaoHgy6ndBCR/2eaW7b0bCYnPMJGWgJ46J/9nDiwIBgcDBBY11CowEpoafCT4R7FKKlN4G2vTD
8b23xt5cbIM8TVcrcDB031MP0cHi9NEi7VK6SxYUZLlTr8pA9JyilkSvIl+z0MGQHuPMXdx2zir+
UYMCSBmZ7tw87FhI19sFXPeZWUz5N/OKLLvhMlCciX1r4TM9+kxI8yE7cK528NU+ejF+YE3jJ0xM
h3W3xS97T459qSAX5Z/yi32tGqtC0nwEBvUHHR9IR92JI/f0qL7xYAm7JoZ5MGuvsf15gstGrgHm
rKHIsMe4aP/IDtvJe4U5Czj1bxcJO2cftJihaQb7yOCTgNZcUeoM6Togg9cOAufK03lTWHbK1vcS
ZNikyzmz+rVRubY6rBPtFUdJD1P0vF+CFZgoFzZQzocfmiRLb7UFmQEF/Wf6Q+XgOMCHs3FLJVsk
W0i2y0GhvlJnvj9VCdUmFaeMAvL48IzMPh6Ln2hDmipz8bKheG4gnAf5y9rxafgzP24j5khq/SJT
2+9JxyAAZ64hoTZhSIRhKeGIndKZ4/g3CbSqlE8rfTYf6Jf1DxHn2mZbchNe8bhVNKT3k685bu7s
w4pnCXWe5GiBpWrYbCwdsqBsNLBpWgRsyg7ncq6X3qB14k06e16fRErDfVJKrHTO5mQMxi3c6Pqd
IdfhQCrCK6mwtMDXbfh1UoMMFo7V5Va9OJb5YA2jgEWC3ZGJOOdLpxs10DywLKlGDbLRlaRg/MNc
O7TySFzwqGPXmwvQlOF1a1jqgxpbtKdaj+lg11OzQ0tpC5I7ZlssTetwKXhUP/ixLgEkJy3fkfE0
x3NHXJm4Yu9FVaHIARIxy85zlXXXaasKo4BBp+Qw1ZUEbDBeRZLVUsXdnM4WZpXcaVpINUNQwISE
ULg8MB1qyWF8+oeifSrblT6gkVWtS/ZMKCBaYKt3E5QeIU7Y25lLZ7OrtQYbOe3Ia0IQ+sBX/g6v
LLHsbDVv4SS99CYFTr6PYB6vl0nnClhIcZfNKUNS3bUIc1RMfkzh5z+iZX+W7TGUTQRWyJWjHH8q
W/BZeUxNEztSGxpJiKxbHR5BcgCGlaSjc+LPQOvE2eZqz6nATEYm0JW7ssqLsG5ohMj7k6oXPk+7
bmQewsnEB9LrtroEteZUXtycBIqUU0k2WTF+lXXDkx1fUK5Z6Gsi3+3fcrfv+nm1mdGTtQN2maWO
f7CuXPLeDZ4y8jZUrOUsBmy2JYtcBxrLIg4BoStUQH7TTgQoekzZQd3naUP0BTvW5rHq1daXmnoT
2dKEUUlpSc2xDdIjDb0keFHQJ2Y8chgckG0zawOLuRBfemaY24/9VVPCJve2YeiMjO+b+iP3wAKq
A9350KeopxV+urmh20c0dnQcFbR0qii+7Ur5rnw/Fe/2sQIX+LjYwTgpZSiwOsc5K1gCKT24tggt
8TO/PsWmvYK6hZXvutfVtcgsWLdpKTHf7gj/Vh75la11m49mwEg1+d0UWeRWbIe5nKfl21WA3GLL
n1j0j7YexzAEuG81C8xNGGsjSu8vJbBxQbVXZ8IQWapmabiVdQawTUTcZt4yDajcv9uSj+ibThTm
i51N2EzFE++oWDGlYFIzniCshWuDRHNj6ATqGj4ME/8TO0w1wzsXIyDfCDaI2Gjca9u0Su8w2UnB
kYvcW7ieJi8d+ELOHc6AHz3dZ+pts9scUTx5bKEgHC9NBysgXEtft1gmdjF8JjlSvBM3bN8y3Pia
okS0rBKwv40EE6j1enfrtb22TU3vXSD/SZuwvdUk2ICSR06QAYOD0FHlSwObHHDI5oppIkEvzBQS
vi19hr4Pm0xpBazn3iPeFBXGH7C62TEM0pPQxQUh1FBhrfJbksCI+HkxtKV32s+P53sTHA/5FSzn
iy8S1Ls07NdE8mREOXzE1iybNG8AvY7erq4Kj0CrAm/5pXJz3gzHNey/VsuaLDH+CkwJGNcF2HaD
48E61KeU/ITTVOEqzdeHXEMaojgSsWBZdSdraBL/jGdsmOb530yuoAqZ2iN3xMR59lhiHXNHRd+Z
wU59opVQTx5xlz8pQDi8XK5znX0p0m+Z9ck1p4bFV20I6gbcPQtU1uqxaQE+Zyd+jDEBd31p+pZL
zOPlBZPMHGYd2VC70m0iijlPGXs/tt4wT1b2J1lwKKJyOLGfNkS+5HLXf3qfveQ8FUPK+ezYiyPI
20xQqou+nh7KGArGvu3KFa6DcdcIoWap+2uTQpbVZzzHC4G7X1gUef67pjZB4fx/10vfqCEgH1Mw
V+7yG59RkXChDgc1HobrtMVwUqQ8OEGgt8rxwsbxhPeerbBLfkQQeNtZtwZubTTH6xGhl08TkzOS
0a3qpHDU34FU3/0H6DK9xifwEA4F0L4UkoqjaCmlN5QzDeLjLt4U4i/B/1xWtCoy7IzrkotzZ7xr
4FPYP75rsIsVDnP1G876WtsYOjSI3bWPueNIT3CLiPAqFXo0/99HXJrisFwDXbj8GUltU/U+YDv3
IdrFfPrFCtpiI4q+0e/fsq2ZwfmBSJB961ZemotbhErWg97Hn1zCUEoMQPeub5GE84Zq+F3ABX3q
+nCVWcp2i0RC1cepIbbsvi3ObrmGzKqWXdRMyh3Gb58V93kIJ57KJhfRlRfNV0Z8h5BUdwsTbXzj
+B2jx//G2S1BYZxLmjw9xF0NiPHoX3PW7Otby3yyipGHgOerlD4n+rQ0Ixx1EEVJ77w3lAErkKrS
z+iuNz1Ladf9DsoSSV+6SmcUU7q382wtJh01ILUr25um4Vl9HCozUEi9nblCuEat7LTeNVIvfSWV
zE/PbM4FWB8zkq1HrtZcP6VRtpDvP/wggfJwSFN08mC6FizRzG3CcVHMxLoJ7IX5HK06fqA48EMl
y7y0H3R+xnecCdWICPpzzr9CFY+KArdrN5lYklBhCyECOc54Cx/5VVIZT9PWVGoI9tO4jA5YT9gG
w89+h/Ju1ZxJ5iFBwbPfdd9KhcD5EjWVxPXhtlIImZCv3K3UyRdl8j9jcsXUvDXsWUdfnsyrgZq7
gqAwm/zagBtJ5OPE5FrgYljl1cmEc1lx6xHn70jQp8C1Z2cVjw1zBq0gWF0x41TXN5OM/pKKMiGL
Lii48VFkMAddIh8EvqUCehlQ39GuncKfl/nvgdcmIJhxsU2o1FtL3CteWEXcKzJM3yneg37+8gZn
hQBuR4T5tbq4niPMR7mJZzJo0K186+vGMOSJT/e1T9MHwPZP8kXvaV9afk4N3oYSVmGmVxHzXUz6
rYaadAsjqta+HKENjNV1T1XonW0v6BoAIwqD6TIyzBjiaS4XZ3tsTXV7SqkheYlxJO5LrGGSXnck
7l6F4ts+AkRh52jJi09xyZ1/V2pjvPUm64ZPmqtI8t8Gzvh6Qxd5JNg64PmzxOs8h+/rcdyqYz+C
R5d4CdwgXwdCrgqJpSiDQD9ybOuqaiICIFQkEUd28HuCVqI4+c/0xXATa6+oWr78UL19515dCn4O
fGsifGnysOYTxlFbirjf43enJrRFblWsk4iWzhz3mHmhEmhbTY+KROzyRuerMRYVC2pO02cmF2Cs
JyX1gDghyvwlVilN3mIgDR/b9QPysKLrBhIlTzIHg8lVb1oQi5nekudmJCVhOCBt4Bm7tOcNkmN+
NZ/vQ1I4KY5VUCNVCH/FnOmYWfvEUt2CrETvWlqDzHgoC4Lj0yx8w1p6Uz9IzI/k/2v7+V36TMGM
HpA3Azno82g75IZ9gTO7/qlT6w+GVz5QTFR5DokkGX9sKdk9WO4hvP8mEt3cGz2Pca7AXLPdN4Mq
My4Kk4OnEhwsdVh5OKv60ByNeEigTqCNaCdtgpbpZU1FtJxsLe6jCSdm/qXGxtb6pNzk1yL7kbyr
RywjmuaXHy1Iecwksy3h+AlibhjlIPZd3KpJP7pFxj6UHPNOXNDUjF6scF/J1UNRWPAwXcMKXSKv
kxQjXDbJgKs69G2KdkL+q0e2VMfVDEXi3s5mVD3K6EcT/Q21HjXmsuJTdi1AhQA6BvccwuhLsF3u
qGvNQ30ERDmFXUBxvMC8EerQ/hqWMHP71sjLbYqfyO12d/DEdlgYL04VWuKG8nKCwPl43ZQhwG1y
+Fh7yE4CZx+kFltMGLYLjt/HASEOHFbCRCopKg6gdlwDlBGflXkiw0rWRXkELCNZRxM/xByWdx8U
9R1A2QLbqVJGyTyw9L8GlMlcWGGWIYoMzMK6m36Eby3cRGbeDHwIvu3n1+q1q/4kty/7k6JSdlgm
B2VCYe+qR7d15ZP2hrNdyPcL6ds4dYVBBqCvPUe0NRG4xMwJXPS+s8mtZFkQycPo3fXqxdQyLUfO
7r64w06iny9i+dZsjkk8LFls/muN1PLTQBaDrREKdFrjMF1vaTFdiyUBUJ4yNEzd94Yg4iSMU1E3
WQqW6bEKMzNE0vaYa0NTqnDoxvutLrgcPxLkl6gfrNsHcc0IJ4S3Bli0f0i7PJUMUcxtUKzwsLGe
nAdueEfQ+KdW1PYmXYI7t/uWdnmEmHOBZDln8xiFdfAHep6Ny3OPlLdVSM7KixlyVQROFrAZMdWv
+1BWhwi6xD2Z6bK03gVGIM3ZE7BzRvFH4GibpHJOqGS1XxNdvum0Mi3KLUCPFgwgMwh4dDSNH1qE
zJt+0fosSXB/ks1s+pzFSaoUOsq5rT7XsTb7Be6aYB5M1vUUcypmc3Hhtqo8Q/y8fvP34TgQmlnC
ntmbzY7VDwkhwUUxEF/9QCCH2YqBcpKsFa4rjAqk889GXBZwmhuPqgdMCi78pwTkvYX1Y0GPmX64
1IBtYRffuRTHOmOwTx0mpmLDuXJO9HYtavJ5+jJ5GBf4b3O0M6ydz/bu8+YqP5gilJ79z+JnJPXH
ueDplbixWZ9wArPAs8O4JrgDb2SgSBXnbwiSW5w07QIb7nrscVUjSX5Ph2TGBHRjpphMZleY+fvI
ZXLB6LdotUmYlh8OCGch3X+vdpme9pttYE0oBsa7jKFFSHIVZeHnT/Lw5HT10rQ53CwUkce83LqZ
ikyQddEX2tAX6ORGnLzpWyLsTlVGKOsoOC690QUn0SFw+sMUjFFF+hFHaVpDuyK03/WqYllxMTsV
qE0Ex2gER9o1ZpFrv5pyP02z2FSmMseS99aWO6ji5+a19CHmX5S/i38k4fqUIpq+psHkQIMdKkYX
tiY23GYHxFgaTLvEmMxX+BqmuLo/0Rp2TttsGTvFjac4yTCloqM7YQXR8Ahj2qxH3vUFIy7XWE/t
K4g9SOlHNhsVjPq89wrQI22JAA8hcHMHbR56sCWgC16dxB0olxvOdtyBtY3sMdPXhuoKgS5MkPUt
19U1uTNj+wVBz5BcLAw62WyW1eOjJr7Vsb7zMhkcsLfu1CGZbgyv2Ybvk9KN1jmEm+ZqGkxD8Ilt
5Zk4D7cjHZhQEwVpYnCGHZsalRjjKWSL20YFEyWE8wDNW2tNjcfibrOivULN1ug8eJ9YJSRePm9Q
HoUPyqXHgEC/F+2HsXUwtMKFb9H6l7eUrr1hJYtpLiNex04D1BzPb1zQpR13g9DWkOAhMTb+8fn9
RiNWxZZU4btVq8IWT1Vq3AOxhV7eWfZsmmy7Zp1KOaWop31dROAaNrfv3gpXlCQ4Hkqvpx0vtY3S
jNqJ+cgM0pDZ2ACo7jadz9RCziEiWYVwgJImu9I+VIzvPX9BtD7I/BimYgAUbDscZdDrQGWkDPrF
i1JHmvDy4AID//ZWoBBKMgf3ArtvyD+i2cQOynWckkzWsJToXYrhb2WUAtseJS8IPyijSBgWCEJW
bKB4AnUJlQZKbW6CAVYrWnfEavpTna0Ik4pkfieJMMPgvMJmxj8i7VcctP76x9A0/UFEQ4pMzh+4
3c0I5m8HHiNIZoMMaw+mwDsireNl8mCaztBqO0p+bcuK8YNp2OHC9JHJKn4w/jfS5zzUBCNuR9od
ujHPCnrEnQSEwn44Vj26o1t9dlL1Az4UnVrHCQNHEXvvDDG6i0mxMU1fuUOVUTAKqpDvO7e1BycU
4ohre6m0FmkjTfXniUrmKPpUQfhro+uMWCvv5w20c3SbdOpn7JhjnKh+6z4W+YOc+rp7jAzZV9Ux
1vwvYwCjWRex2MH42siWfnoOmir4XPusTDKO6wJJphVyuoBmJlUB3BNKNr9vKq7fkKpQ0hE9qnpc
+9TMPInCBvH/ebDA8SFVsyxTiWAkP+IhDlwykDbNtmsyRnX1QRHbIi0dunWKEN1FTIYJdfEPEMUd
LRS4gaLRo0ss0FFuXr+zaXa7fl+aXgKEDwbFvtA0POaamV+V3qnf+mmHBoVSnpmgUEoRGCK4o0kE
+qhKVBgSesOSYB2dRtgAvU1yQ7P6xWcbi2NdxZnt0VVUcIHvDsQyUG19CRJb5CMr6hBd6Qwzax5g
dVsaa6CG+//yPi3ce4WG7qXACyKC8uiHfppzqEY06SKgTRt03v6FmyhbifgbXqBSvLTYtfdrwS+D
wwpViXwqZKAMKeyeXYve+PlEmtAjyh/qKY9JFEa9fifqOuZfq9uAuugPnfGWv7HSWZWxYFobs3vj
DiTyPBSrXMYipQjQMxfAapkFl7dX0xInap7AF5SD/Hcm3RU7vNf1GmoWfDA4YSowiv4FCwGRqah9
GiJ72edVCSTjVw+WfcZK3iJS+aVfWBlIqm/1IQXSQN8CMT/ezrPxuqR+41vyTV9gdnIqyZS4K13z
zq3uq8JNBKHqdWg8VdcngXPhyQxftEma8Zy2Km0qXmbWTNLwekXjDgchz8jvbyxI51BS5lDpDdPl
fSZO8OkTi/To1OriGa5v/4Utb4vOGBV19tyVcg1CnzyUhAz4dszaQFd/L++ziM7YxuExnqPjR5mj
S748c9JtzvbmNLgffzQ/Qp4yZxvxoDOa58DV1Nsc+g3fMc7vrgTKWeA+WzZGiDUnAbFbwO4rxVvc
1HE7fd/0xrARxR4lGQZscikUNZpqLc+/2kJ+6keG21gJ5bY5d3WuJoNdsejSC4itZqu5teWmiOWx
6ZfIVl214uhMe7sHTOpFnFrcWZOFy3J4GxcySoMGiq5XVZSZVyFa/svhur71kBPc36kUNcUAdifP
6aqid8sVhXQa+xWuyUs9RbxOviYktTnXeI6jWWKW6ABhmnN3dU66kIBCMfTKlymmDbMtCXOwqg/K
Tb+kcrMTjM4GswxDUfx/23MVYThsADn44QMLGSJPLxXQWYcfOv+EoFnz1+S58wqQRCin9zBTSLCY
3/H2O4bKRN15O9pdCYmLjpCdijBp8T08VkfCImgqT/izUtMM3eLStjtCIdvaDJtH8m9NBuJTKrLu
/sG/765DlI4onD3s+5jlBUDXX8a9XXUylBt1JRwNtMX1LGIN3AVrTKQ7dx90yd+GGbw5VFvLCzdc
XPO+V8ehKrTq0eO52QAh/Wz6esyFFJJZtjvT1Izh+8QHIdsgyr3Aar0ralObokilZfFH5KwoWEBK
0K9ZClE3isHb1YamcC77ZJuKSfJk0aK4Tj7p6p1hDXcZ6HBRZ7OZGYoqk9jgyePfq6XltN2A4isJ
lFnObYdNcP4SOmJIZsV3IOgPAerLIoSofKg9M0Wv7g3kvUCTdIhX+8v9RK8YMtr5AJSOMiwmlIuA
8h4hF4iZh802qLcHvOvH/clIr+BZ6Wgq+aocUWrQjNeG9d32Ewt86Fs5ffA/GOrMMEFPdybIcsIX
O6izZXnMyMTUhcc/nebkvHbpmXMOwM4Qe/xjU0Yr+AFq+ukznFQjP7RkhuEklLVhFU/KVrY0bJK7
ij2XTvMCaY88J5ESvW+Fjm3dDCcDqQ/z0qGrIkPBXFDecsqJKAU8gg3IbuY6btkblZEByqQoylPH
F61A5+4lEO+5S6pc07TnlP9Y4zXPHuIOxSEwjEsYbUsXgIC3P4jHtqNz8keoKSAD0fYJ4CGDoHb3
156keaVSv6StrS6HtwlQo6UXVdDQ73J/7JFVTOgqsz7BCmIIJdXVC8IjPxEhxvUjIZeiCIJTRgY1
ZCkDMjoEQy8ZPLKyFg5nWbVyx2f8As+21MxsSewCW4TWlsqWERBEWee1Ha5dq+ICPfrILo8wJgpe
P3FT9PDr864JCQBFktGk3PRu/PI+Ok2wRhYWYHt9M0J8TZF1ZaaqkcFhzwylPU17auNR8uMbqtoJ
SeG29z3Ejy8eZlyu5RjqEeuxQhG5G9b5TPCxVtyvkPL+/wagdWkZxRunAZgsRIzda1fhhhSlZZey
VrvXVHv7AopiamuzDapDsEwwwULSnBlkrKNKDsozyItOy315elvRGyZy/wKkTm0Q1EHj4goj5VUu
vss+aA6YN9u9xNJ0Qu9QRTWcyZbWyh9+gHpumGsLA3iN5ZonOTBHInudrF1XY/0p+vfSnekSTyTX
TElIAuQzZLBhJLJvE91ycog5zxnDyjcqKz8i80B6PTDiuQTjWV/ieo77WOA/s8HHM7YjwU8GB1n4
C/dqDURtXN13O//iYVgAFLYuNplIYbnPxvT9t6VffAT2NRP+95DyoI0AWVoJqJK0yCalLtBt7ksN
Udv8g87Gf05njcl6/hsCkX+sX1DDAz295zuLB9uqpStdbcLwQQy2I0XfUMFHSrBf4NTmVMrgofAn
wU1n4udB2GvV4ga+tHOZcT37sfd+Xd/rXlQuc/JZvk4KPPBDjaI2kouRYB0nxl5zWQay3GYLkPNQ
W0fjBr+vOKkNXY3NVTFqEP4MJqfozVnmxeIUyXStP0d0fhSiDiToU+AmWyKcFJFOssyWsNJdDBkk
99SzFYZk8forsiqv6EsCqATgBLp/x05V4vVUytgBQ9KwpArIfVQ2k57so+Ljrp/0ASCN04eu4aYe
v/L4Py+vZk+K0O50PXai+bP7hNpK4cM+bDU3cHGDJvRQDkcLyJEWbYoxuFr6vWn8Rln2EX01hBuC
hKzercGVdnC3omHt2kFrIrCnBALa+Gj45ffr2h5X0dgFhvNoxdgjn5zCHBxMdLQ9QZBybI8psX33
3APkejS+3VLp2CUqmeB4zazKMg/cOnJPL418FN7y3El5MITkcY55KtAyhYgrcnSi7VainhX7nnX6
+T5MBBeH7Wx5GtMNo4c2HeOMfBA7Ck+t+VKEmIBr0H5tzdWnox7DaWPfY42HtVESevSEag+ct7sW
+Lb+kcMxupoSBII3igA26R80p6K4en4Jj56FHj8ltQjnDKIHtlgoV1dL7zxmIorjx8ZKUCtDdToB
wXCGk3L1dsG8XcmKWS5S92TqVI4XfYbmd5l8KVrQTNPbbERXbEcNC7VtSAQFH4I+I3t7mKAEKknd
IvpTAjLabNuf+MKK/IXvIQV+jE+FNGvOeooxzYuVP+IZIvZeYml2lgZqahquQLE/8A52nLlRu43n
iRLryrZqhLVhXEeFM46D6ONMnBw0porZb7hoR7vmNNkf98J+8sp3NuBMRUreclwmL+TxjkNa29KO
9mVyd4HYpD0qJ7aW8J7x7JXSoUDv+h5boG6grPObyym+MpJ35AK7IpS0D2XomF0m6+86rMk7m89T
1C2OYB2OHCP05j7PCV+sP/hOwF0c5Iukt2y2pta1FFDwrF0EXHqj/fz9Q87RgSVIzrZSGRrAesF2
BhKey7zSJ2frigVgPHEFXn38uVJPweEEUDsgu3iLEPhVkASIY1UJkTWo14zV1ue9FPex3t7mSgTV
pGKuVa7bE2I7zFwMAlhE4+GTFjD7IxsDLgSubVfWhMIE7BZi7anv7rAa6YOrelsFDWUTqIPPefLz
VVPTv8HZcqVk32pstq/pCEftoPhX8zdEnlQNi2nXlxKSAi58G7rHZwHtq2SQVKCkIKsOT7HaTIVX
Y2nD2HWjMcSawboqMMzkm8sJz8y2EsA1+OFulFh2kCN2GXDcY2JcevYIhdZV2tdn4+fhAgeVz+Ko
L9s7Lk8wI+HDzTpYUWZulhgcYziN9bUQyZ/8pxGfASU25Y2zuO6d0X+6Fi2WnRU7DM7T7mexsyMI
5OHXPZkCzQvK9YEOLv/coJ26mKO0N/Iqhw2kgujERekAvHrAoxzMa1lB6sUVMYtJiNUT3Z9zxeM8
nezrBPH3nJWMUKcIdUZfz2FRW1sEPCAm9fX7WD/JvFeUOU9fIl5ZmDM7cWCQ1jXJ32ikSlkWHGWz
NTZSVjmnDFcjpW1WBBaqy+L17vmA8xnAk1oGAMQ2a4Maf/UmgA1NGsPlQCRNcs2k/kqWyMqH9Od1
4lKQpc7fUNx54AtCnWiPQx3WUpDJY5gagwQ9OHA+pRRhQtfJrE7kTFe4pX5uWgvA8gwxEnbXiMof
LDRX+hR/kkOitMOrQh4Ws61U2TU7ECOOrz/+xT7tqIpl6rY51YDsFRH1FrX1RUmjvXnMPeqODUmA
tBNSXS+PrsZFjmpRKy87QWBxsfRVM89YmQYjoV4/62Y2IEJlp8lTZrHSpUSfE3oWqCSFGDgcF97R
4YhgloVxU2FB3bwqRlIIbLHSR3yuX7zXZuq68Ouk19qt3KpfmKwsSfky4hfiu2MhNiq0owkn8mXU
R+6n0Uu2wXEf1VJM9G/Dt7XM/6EkDNaUttA4d/gfC0X/Zv8USGbWFPORpwAE26M4v91+X+ILK656
Wzoq7QzqurSf4gwpw6DxU0I2WZWgf0CESM40B8BHhz3EyIiaDUvY3RE0MaYTrTvKpOflenNvYjUb
5H4z8AWhTgbWRAx9ldlXnOgsy7oF0vU3o5LP8Kaza/z93BSiyfJWeQIqRQE9WFhV+Mm4tg6ALZXV
IJIYhsKVdDXN0QuFg0091IYzQd6qDfzW9tB8vpaCGuG4gd6sNLUXThGLlxuBJ2jNBTp8mZGYCw0Q
nBH4LuC3pfY7X0hDzbjZSvYS5AQdeUpkw8UnH/2pdOD73AVdEs+NsfH097i6EK+S7cU0B5ZN66xQ
MbdNhmc8lsgOneilNXiyJgfjVSpXhxN8WB2N9cqPaCNK+FmdDPdCntAkg+MpaS5M/O7fg6/xBMeO
IaOMpAVttzL88U0qaZ6jbanOluZ3V36xe8NF3yVN0FVw//zHJPNPQ2G/40BGjvIGItKEy1hbNCvC
FwwgsYmzcexRvcBh2k4YUJYaLo7gdEOyUacG/GFRuceAOQNtoCtPecf4Of66hHznPlBvpSKtI9Ma
8cEhmMIq5FR/AeRtF0GV4rzTqhEY/dxn5q9rCBMYGWgvm6HXp8PW31eYKTfDWW8y2ncRQhXkWs33
hawLyYfkNW2cH0r/7gevfEPJ3ZLomNgiC/pd+8KqUkgKrbZcvFP1c58xcpcYgD6/hGpXP+dcGeyg
XU90NHWzJ1ImK9degxtSvkOfqyvztkRHm5cEgxxbZOC3KaXnjnLGErLkyU7GcG7oKBa7UOk2j4B+
3pyHo+RlLQpRazxi7OwEtvSqbaIPVcDYNewLpFQAIDAZRAB4MFTLhdsE0CQ+1CIGrUjyU33EwvPw
oaQ1XQf1Vs0icLXnW/m5EA0IBIzqwJIB0lOVCJflGtMkdADlvRuuyL0s3JEs6pB80oDmCBPPXaPP
y6bIIj2eWW8zSQQ2jISi5f36HRC6Emf1TMlSRq6EbOFOfjdHTktlsnzjVnzsY7Tqw0UMI/1sugGa
2KjVTJuAihfQDFR/JHY9oJ2cB7zfYlRLc4OEHLKNrpS7s6AFy/r4pwUL1FUx+DLcw6p0tGOos1Dt
Yvs5IFwC9O6gNsYvR+hAa/AE2WnmN1r90B5FYXGe1FvG7i3k2SKNipFJsQG0prExLSb33L59tTNi
xcRe0Kc0wblfSdGrwJC72bvdssi/g7paij9p5dCRR5X1ZcejiQmj02ed4M0jZMjVhH+tVtjoMZvf
gl+6EvUH2FFpIItl69rMSlnNh7/iQDU8260TJdaJ3FXb4mSZt1M+CoVPBofA1EQKxfKazo0lhycb
MvzIOYvdTAaCsjoMfemmkKjXfOCvvLzTeVzW5G8IBzb5CeGsNW3RslLUo1NR49mw8xBKjXitMVSW
YmGq5JmXiQ9DOBrW+BDz/9jysm4vgAq40BNnQi2bAoZveUe14dE7vYnv2d/MLDmETXNO0xMC/c2g
V8TVxehM6Zi4OBGdrTXXT9wXbpgdjJQF6umXMgZrefryBS+F1gS8DJUpHYvxERAcoX2N80VfDY5V
O+506uCLhRKYZomEmm3Wno/244RpxnPkssQ0KGnWkyapisLDdD5CWj3T9ne1J0Q9xNcgFbazdRzV
npYEwd79BzglPMDJAyvasGCR/nFR/M6BWLTRvZTPh1ZyjO+o2FnYfWt4BNq3JSgnWsSL23e4WgXJ
U/O0ZDkjrUOmLIdlMlcQFLu8Vb3Aqxdk0wYBjktZXIH2xlqwX4WWNbf5BBGDhw1eD9K+I6gNLevn
7eGeaNsD7F9oPaZS1oJtE2DGkvfk9g9PWrN6ZLGcyzrBSZuemihZ0/e5AvBuSnGtEUWHeNvjLYAe
6y6NxiGfyAgZ8PC/K13lHNxpSQFWMz0MfrlFBSnPONejtt+5qu9T1kgbFNi7+p24zjTmT6sP16QX
3mq+WIYCV4TD4Y215/WxInEEQKdDghvYWCZwF966JZlBqH6YgivL9y2NseHW8eTS+tzcO1N11iNl
EgQql7g19zEqOa4HRScrkIgy2GICDkLaZgztFpdyR1gosI8m7LlMuQIKYb++2/ap0RjTr/Dh6huP
C6lCg8bXCszLrVNGR2uXM6bD6HsvVSQ2WAZKLcqcjA8BhxNaSVucIDwLwEcF+hs6/L9Hn5FHq5rQ
Qr2iDJU/VywVQz2o2icjbcSmr+gofMpAejZu/ljweiMRFme4yOdz1zKfhOWkNlAHYu9xQXp5Dlcb
OsaOOsDmFx+UV0nzeRVuNng2092DIwzddvL7gTH1jb2fkL0FkdFCOzLrvgYNx6QHRZQlL65LO2mX
scdnwHou/meMxlBnm0uwggr4SXBeVRLClgL7HYYEH7b4dDRD6siraMWx7ikcEPidq48QRTwmPh2G
A5EqHmYVITXFVDrrVjfbMglIwPJag6YYjRp4xoL9l2f0SCG8wu66IyrQN8CPrljL01OrMQZOpzqs
zxNTXzNIYaioAX7Up6q+dws7F5CqNFPwrGm0WWyS/BTq9fT/8U6ET/YD3q7YxBO9/sBzoGZrVnsi
hIvUeQGqdUVA3aoKu+TyG1gAj3c8iNClOEh1pSuZ4XtCUXMO1nWo5i4SwwvXYS8ah8RYKlKWeVfk
S0Fq6aENvHxIpryaNiGfoYnTOfIlFxaSM7wXVZC/3JgoQaUmNPp1PipvvCYxtQkDNjKHb2F7dMju
P4d9ak3iYA9ic9guu1Rt229zUXB5wgKRgJtAZYtXFvgtcs9DGg6W5b5/XTBAHK0eOdjIIz19dKjc
y4aM7zur8wz5v+EDN1RlBdox2G5bILiagTE7XyD0nNgpWFHTCYkdbVLjZPEoYkSpraWGRUT9iv0J
7cMrA9yRwLR/ueL8vODV8+KbXnCvonzKGotSrZLDeGCs6GTmcH38pUjOxWKIa6D1O7C2/YzA+ztR
2HQsdjo5YwuowSehzF9sdFuQ7QLdpPYsUypxLDtHRuvDbtIvGK2qXH6GF6Wh4dm0gB9lJC3BCrK/
AncZ1n94LlVKv/t9Noz0ahC1db2eRrBPPoV6j8xGvovYIQJR3rJQH6NcumcUx/I624cyRsFZ78iv
wNlEF2Said3R+NcGhy6vYtrnek0CCBdtZU4/6wEGFfTmqf/lFa5QSjfPEiDrvUby0PDetn3MzmbT
cRxutdpm5HuCsXZ+pVBsf/gHos9sNnVFjUM85erE1nA3qnUuEi9/WgkyPY/g+SXXB60VUeq0cxvH
MJOR3mnnPQTSO19Dn+u7/ZjdXna67CmQ1Sv6z7XQdwOyRES+x8fGaXCKEuI56X8jug8LqCRkhfcM
t9lrdCaiN7viECyon6hJhIgfy3s+gPqm9CR6+0sRe25Xqi/mJkNzNAuCEoRYtQNDgUWnoZ28f8VY
pLb2ci21JO3WyZikHXUeiaLnMGKnJwUlpKCscpX2Vu3v+DluaAl6q7AjkYtwFxW1lyhDZZHi8+5l
9mo7BS12F1T14uFOMjJ6O19blfoVaLVvTrP4BLQcWmxt7+HIZGc3NF0L9QJ7JcEMS+Fjw+5mXLsa
rWc6X/2wAlWA3Jej0mj2jZkMzD1WnR3fjtYMG0dbnLFOanzl/WM6sYUUNTDFFcU1XoNr0YSGfAkV
L8BVcMCRRPp5Vt8ZfWCdqn6VFrjQO9nw4r+H90BNsUlFyOyggQpxTKxhHE91cv16rAFHsMbaE6bI
hhOvVqWaUF1vcstLKDIUBl2ZTliaz0Au/wao9S9NZWEm+HNZcoNKKDN6Zhvch6sMdLaL0Hl09TSz
9ahqX3UxtMuAYYAoz+ltECQEyAc174IN80dcg3gfeYSNxd4gdGRbIdQ8TVcbAFAsBH+8bNXl14Gw
W8VyJZR21Sp9wBgeL1uR3zZW3oLx6KJze/xeJIWl3epDmjGwryMOBRb3ZEXnNFa0rsZujSPoS2B9
dqmEi75cTwgf75HVcfcOSKWAbQCGOVUVr/WjGyurIeUV5eUmLlOJKYb4GCrrXLhrdWqfDwP1lBsu
uEbZquZ0NXyEa1g6RzgqQ7QhBMPNDQuKXb7eN08Yq7zdZ1f0UIevXZ7RnfC2hfcfi05RtPSAZVFN
Lp9+yn2ePb2Ug51Rh1a/C1yGeeb603JTSX3t1sUQeSUds5RF5dDIqDAMjadLIkj2YBxvMRuJl6Qq
rSRX6vRKmOaf0zqKI5HWUyxxY5fs2W2OHZuJzidQDjHkmhCZiZ+q4/vloGBQzknF/uwwM7bQfDEH
FIDO7Q/XjnVtquM2AvAwytVuxMdg1c9KFh+NzUvYhhCp/92adyHmm9s4z2d5zYNd2Mie1KiS7gXr
Lm0BdH6yTN01daCKAQLPhFrWr9A/Kb4eUQ3YjsBgExXvh9Ik/V6gu0GTSQAyxqy5a849A07gWdgJ
goeJOmxnfzX/AaKD4L6E2U3JRin/Wwm299q7PwWJ8u15wYoumQGUW/qmOOgdq8GgurLnGWDdRyIG
4dL+MSg+VN8Zv1Ry1rV+j9ICjCe+l07nR7D2slNgC2TImx3YWCedT1s9XmUDplKRiIbI+efqVUIg
BIwKNmLdahg7x3XD7KMWmg//OmGRNtzG4jGQYG3duJJkijVR9K4/vTl8mxZ3MICYckonzh31VrGH
Sn7DWmVqgdScFARpcjJmFkWxcAts1m9NtQe2G1HBV3BjGOfhHzBz7/PBZApIpyFbD70uLkVUBvNI
DSxO9skaC+EiphkhoCDykVWyGT1297RULP+RsqtfmcXwHkib/AeWKqHiYfBQfsUy0FzORAsyeydX
cIBLsYfAT+Z/eDBsepz+Tmgk5XwotpuEEzC9T6EHXT5lw+dl8EWjdVeJJjhK5/pSQfHoIxlhGkCK
fWymDTu06A0wxhOlEAYlz5ZdblX5Cem5PWPstSruWWthKpDldTdvRHY7Wtuqjr8nv8DZoj7VrUrJ
NzepBZ4hMV+N4NY/w3QYmz9p/fGKUZxpUuQGgUzDboaXA0uSVI1cTzr6djoG6Vb4pYKxcEXPF8dW
wAxd0nsXlVUkHxPwLw9Qt6YIpl7d2MeEefqZ064xIFbhiggm2DDp5UrsKRH170IuorAGJUmESbhM
RoxsRdK+FhldrM3XOfLDFnl/uffsiK6/oDTQIrdqBq1u78qsOlBNZ5xXqiqCoFCQiYyZXAk16GnJ
GTxTIOynuxrH4kX7iz1LDITBCC9M+9Kp0u0xDahgRHEi+JJMCHwZggGFLV9PmX4BEmDvlwgcRrXZ
8/ZSqnwuyPUx1va9DCEavCJ6nXJknXO3am4FkbmNJaHULXsAxse2Su+1fvznl56g6WnOjCMj0QLB
IrHDXQRZgEffYh+w+GYuM8UE5Z/wgZFbf9rgxXQN3dU+TVUYK7vok9I/AObV9s9wuc5+l5mWUbf5
fSxMKz0Uo5rsDPTpa9oL2Wx0BYNTRvT99bSBLSndLL+W1y5wYUZYex5NOXDUMSnQGbgTdQERE9P3
nfjX//4NmQCDg7Lg2//3Zk6RxePJXDAa0anBd+x0P2a2xymYofpl+L8ydVkWcmqt7AovOGl5u1JZ
bXJfB25xBHg5JXWO1XlYEpnLAvjAg/ZuVjzCpR5y54vK2TfgqC/fOw2Y9uqnTA1K8+qXIONY+N1X
t3xahNVcZdBIoOa4Oomopja0Q+Eq2enFNRnijOz+SvuH3rkIkTLZjUCqDjhV10dogCmWCswThzv0
hyE2ZS4Mj0MdPe7PzvpJn00zgCs072dW5ksnzTPxcoAuvzE03g5bPjh54VrnrbdjijzYBmXr0S54
kupMg/eSnJRL6sVbQ90UxrHMZa8glYUAseMtGbqahRrhL13NO15Ip+BuIdckGYccnxsQpXEoiaOF
pXyTrL4i/oK8fe18cY+4gUtvzYlpSYb3l2F/ppktNkKTfmacft6hv55aDFPJjSFOnzwQ5kTcG8EM
gb4TpXEG41AsM9HLdUwpFj0/MnDBBlFVuCxSdClvMNqpJjkBME/zpo7TaxMP+9mzQgjGjz5j1JUI
+Dp4PFsIMk5TJOCXw9xZtynvV76pQD2eCckka4RdmXNbW32ffi4NnNRakkrue2TSud6tweoLGmyc
vW/x5sHO1stOTdPvOPvKh4KhGolf1iRyUmKeoZZM+65w2t6mayUoqaq08xrSBSm0CvFC8x3uURC4
ftmk17mY1LOxWnUi9lfRGNmFFOcdnY9sR6Zdg65JOKXfIVhiQ18gU6Yodn36NeJPm2cX6bzHAu62
SlTUtyQLN/KsF/T0cAWcSvqXyrLBdQtWUMwfdfDZOhhqGQo0ZBwsJyPoyr9oxRbFcxmzYANYHeS/
+P8sFsK8+Vaab/iBmo7Qar750GfFYQj5qvlUOdg2IyeZ4RpsWnoB7m5Q2SAvrTeNw24DpAHrXauk
7Vb1af3NPXXIXI0Wq5tpxDv2VvZ9hZewty4WGWlZnGj53robGH5Aug4BQ935uBvtuPNsRaevJqzI
p3SjIE5EvEnE/nEb/4gdFiiC1baOeSiS6c8EIEdbr0XqkjbuLvvf4DXS8Iob6XsW8sh0M5eSOWSC
sM0aVGHgVdBN/k9p1ZfEl7tTcnwC5/UrS+GUarbFhtwVIHjyQliZwCJMTd35BbPFTrpotDycvHeH
5u2iQacB+iB/MlytQmZFUdmLFK3vgNWS9zNjPxQkEpCPWhDdUkQg3JViUOg2vv4HTBnb3LxRixjW
RTU5LQ0xtRpjEuJ/6eMVFoITaatTtcEubTZ3deuLAv5Q9ipnL0FBWXthufbB1WdN+K0OvOSXAcaK
wCb6z8YixSZR0qqySq1bK+hQzqca3wtLNgoXj1pzoNWMFkDW6OA76sWPE4ZfHjstdFmJ5EYLF94b
+BhxynQ/f5B4VNSv7vR3rXf7DIzeqGi+6vKdUyjtiNPSc7bID99Vjvy3vDkyjScRRtNn9r6fXzT4
SJAZV1IcFndxdYygHonx9ILtwteAtmFXtr9lFN0a7OB9PUjWKdoy2NH5YQ1WC3dW5OSyQ6HGabPV
pMysZEoOg17fOc0UPlbm8Za8hOh4QSnJUhrNhc/529ujJ9nG5NuqInRU+dZhg+LCAg42WrYWVUnc
CnmZf1VKfUtN3mDz4ljHlttrzPDF6ttKcYM+/SVe2rpk3AfjF8e5cFPpRzrsGEyOeJAMkCwHFh7t
nWYX4avvfAp4LSMdO3uWitIQOa5DHaxsEKQx3PDimqksv8UP13d0J/2vAswy0/JVvPMgBQaqF0QI
KpSFvPne2jc2bHn7ahY6NOHtkOFuYrTerUsn0oNj4LIoRKPXjVdEFsfEJ/Nt18wCYLRBROVzZtv/
1/B7MYsN4XGPx0W/vtLndvXmjsnuriT8rLqSakXxmyohWQVuwifBxLEXqhu1zFjTIS6A39oULZg9
M9Fa6iy6DWZXoYt3CtljiYDWm3Ud44JzG6dwnNEi/mpn05mGAaBWrxOrQzGjafPmE8sjvYo1p6YD
Idi5a/CDz0m/Wh2SZryOcf/1bmiEs0zxYWw+3BOzk7++9pkcwGCbIRFNwlFemZ+86H9iwQd5//a+
BZ8qgJYmSsdoHEGAXKYviLDEyG9GVVqz8MTpwSWD5nhzUX2sWs6HmqXQPC1K7UwRkg2npUiasckt
8XmnLDqtRJyfbzXJJfkUZsju3dtGE9ISgrgoL0gwotW8ahwQXDnC+vuHeBOmmm360kU8QbBNUA64
4FAvyeN71J0QKa59c1A3QINhZrrWtnGP1YPsJM/XW+oLgv5NMVYoco4ou7oZkUtXQnPh1JAMRNta
7GY7TYsgKTlNZSktTREhgii7Rsl9bywrrUlZM0hUYjc1s9DA2HiFGoPDogO0sJV4lMk1kpTU4+/s
lnL5jA6ntVSiQJ2NuhqAbjLyFkXoiEukhqfZbhT+54e3UFNUhMdA1GlaMRzXvNhoV1bT9Zh+2Q9m
ltyAdsXfGVGooElHP4gJ+Stmn+dN3Bx5rsGk9DbIzIx0Ft84AjexmnuolBctMRtANAF+8+t2brtt
AYuPtRehfQ52Y1dky6sHOt2yR8eEQM2XwITKfT+tYKPV/7A0YwbzcFO6ayNxrXqTIqWrfMYl0knz
RnfOpjKUEY0is9w0qFab/Coq5R6oRLLmNrxIYGrxfKWlJx9cFJIliLzZ03cwXovdvOvuW7ZIMIz8
EKC1J0SJajNxN7S+UE/uJuNhscKbRcZ4jr5DcbYTlQXqT1cgm9n0KzgaqiWP07HmlpHAbMjl/OEn
hTHpSjyR/qR8VdVCGzoPLLkLmHzn2Klm/ZcLrByfMbbpzvF77XvWf972jEiz/CeYQQwfmUEkaBuL
NbJC3285iyEzkVCcf4SO7aC6V8lWw3yy6bm3x94lQCLxFBJfQC395RDeYXnmd2uZVY1o/+T/4zJj
uR3LJMEH7D28yS9B5gx6CSP6qiRBhY34eCaD/FVNeGexzj5mkLUw4PuWpLHLQh0toNsps9fHVGNM
MM7YYbl1DbOvrO7neZ8ZNHLcxnVrJUO7oLkT4HN7xtLtUHnv2+4Yl66Is4wrtQP30VToMC3YBoFo
o4HeVP7H4Xw0pmOOsBLz4E1LsI19zogmKjnKs3BiFxXmAP7rrUZEpaJTcZtieIGr9+ypNqr6fkb5
7VR1Qi8VHXJmopX1sUFS4aK17VryJi2LfXa37w8xjvw4J3mQJ271UeWCgJYDTrsYEqyQEpKyzqzA
WWPuiuSa6MnqcLF3aEU+36Rdjvyie4fRTlhsXNq2qreP1fUsB8AdG+9uC4W9ooSoxlSMlarC08OV
ENhHV/qXAUWFapZ7EyjRVzLJj8abNW2K+cToXU7bFXhULcsVoUJRJC6AKAskhEROpWH7XWzEf6/0
mfxBBdPRlJq68f1FAu9kUN8B32sMblavTfanFpeWT8N+a8BRf1CuQMWLXHFxlVkc8EYvyihRAoxi
fc0mBbGPnXW1+b+jqtSoYILkysDa1GkhI3RTVBIGy8rZ/6ji8cHKl04OtsLhsUOhLK5SJvdHkg+F
A3CMJprHdnPM7hl0WK97VMElwDJVJLdgz3kt+OFzGqJQRyKfDTxvaXDwYhwj7gNzNdxK3hkaxsu4
3CHUDEhe6JsNlBPl1xWiMrxwk84LTPbXDSckYaOVi+W5RiCtTFOdk/FWGsoKGuIsK3ZEXwBtVvUT
JpyIM7PUvaxBupKkueF0gRqm6ff5WoGGAkbTXqvSkJ43ExgLGDt0M/iICSb36l/Nic5b8sMHAknp
D1gfON21yNF8+2kFWBdzpb/1WaYcWViaTW4r12Sag7ql8UL7XDhgXZgdgB4dEHel6WV4WSNsitEs
1QkeIF52lnK3pTmBIzZYpXDLebqQVdHyYleqijuhUcpp7hn7Q54kdGVLi9CGj3rQ6I31aqzKJYp3
OfOPILsv+l207h030ybFSX3u8g70tYmbChDqa+6VrsrtBwctJHZYWTSnRdykaqE/qY/2sOaZYoom
Tmau5FJGKDHASm9CPhDSkQ0khEnG0SAIkBLnA5WEdVTUWgT04pDRr8hEdabcNtGcZmppl1mBpZyN
qKrTqtgWEAZQGY3UktHsqzRk+2fa43u5zR/YbZ6UwJUpndU0EG/53X0cpqwAhN6qujfg1ar95zKV
AIrCoBtMetexilYNe0isBDodiRITq/sHrr8aHl8glGVlIs439f9MMKgp/+d1Nz+y8WE/OXC4yHt4
3UD0fAjpvrCws7qBKFMK+kJpyLS2eFYx9lIsh8gSwqU/RVALwahV91b7ZbdI7xWmsb5KNkLQF0zH
GNI0RcMNoVCB9CT1KsvY1aImHUrv5cSd+RgX2A+QQh/NJDVoir1oEAnthWMTiaJLEpI4LF2f/X00
+vsQtYimGrPUOqgGkmPUGSUDlEuoJ6RVLPNWtY+W24eWqJbndZF8DlpcmqvYD2hzCzSb7RocZc/v
kZ6yy77jp2dMuKZkwIhkXS1tbRsGgMVxm1ao4XxAtswrfPrMybW9Wyjnto0cnl5s8PMEeb0mTriI
yaIO7fOEEI6HIUNIDVVG+pMOWNDBHLsWDEJu2ARkshbojCCJVhuek77MIG++OKF8bV6MW1+hdE+9
2rS0eWLGBI56Fihk58n7OiPi3Z4NJjEivVuiwV0vCUEK+rGVmjvEr9th8kvjw9FpJcSnvgPBr7S/
e06UiZI5QnxdPd9WDnfjkoUNQVITJFvat2Vr18VbOH1Duf4ZVQtHWUvaCTRG5P180UJwJumiaW5w
fEQUruzWFt81j2KK4gErikujQ1TiV4siR+dEq6BY2EuAe2kKvDYumR4YxO0/PBuVL9J/cCFOuPsq
KGtPyob+V0X4aLbZyPGeJF/Z6SRxufrPpx9A0oP12qsMreLYocDAKZdlsEVZTUueAUKaiDC7ey+y
1Il4G4SKv23CH2QBSX9AwDmE7PQacBf1DSvKwfY4Tvh+euV7YGjq0EHsHef9uMe3ba6CE2tqtitB
ptqwlSoKV60W9/9jCN3vAlbfk4FsYxvl/6u9D1B0r9R3B2rsemy1E/iHEIoGwY4PeFW8Z48frJFq
fCWQxeDQzJ1Zl4wluXAgb3+6GudYeOm8W+xZNZYaJhhDILHuxR9xrr9iv9dKaJr3Upgo56td8r+I
OhAkAdDr8SRtRCtM3pPw4SpEup2BGPvF4+rO188rL1aZZFHwjY6TZIk3Y3Nx8dJcbHrKymKbo0FY
s83B8dxbTYYgkRskVb0bILpVWkfeZFmzDrSzcPY93eMGpoe3UqEPnyOla1tM/QJdaRlKYEn6LAwh
56JKTF9oVibTkDe2WYl48FuK17VMVmZGq0Qz5UgEUhi49vTDe0tE947zDnAxweTIt69TSbajftin
/F2uHBO4+thJBryRpbg6lirghJR/c1cJW9qGTTG7phVxTi5QtiLidX9jxRI8WRROWERnYr3DM/6G
oGHq+/PjbSLm4T2/ioMvuorucnEFzMiQELp3Jwdo/KOi2MGy12snELWUVOc9yXcPbGi1PJ8Hvyvd
zilP4WtO1MPF3+ztzx6YbeqAO9sqXOOX7h5yuksPxyxjWuAWa7MdGD9e7nOfxdTCPc5NShaFzr02
crE4MBPl4eDhOSke7A6scosKS7xN+iNV1F8AN7GB2Vz1AzTng0xgqEUFl5fxnUcQmJR0y888LN/K
AAx+cLSwgOPPhTscEUVV0YnVPICWr6cSkxjHlauUzXXFC/Nhw+eVKlJZuOFwUNCCUdaqjPU8joN8
k1mvKCAddxs+Y+XWBGJX9ZKBYjh4T32ZSZHX46mgz0+v0loxNqalc+mFVxcG4RkdLQMQbMV0SGRs
7ViJr/vq77vG0g8InnBVf4AmWYEbtNQdvqMDrtpuGXFVG/qgRhSvSHIHdgzqfqD3lOktcHK/E5av
cSXvCwXUkzACrMdUu3DEiN/WIvX1Uk8hGy8/4kB71SdolmGmx4oEYFh8PNn7YfeTCLI67iUcLzoA
ibJbZNXJ4Ijso8GnLuNyktDsccPcdRfRtMTLlDEscoQMJYp7D+7fkeGCIc7zF3WNxiLwBFfm4dBR
nAJIrx8bU/jDxBgL3Oy6b3GcUYYexvW5wYZvu4YlnM8Eo6QAnhZq4XL/WGPcKfl8lQiQJRBKILfA
LMbFP44j0dX+SKLlfD5sUGnMM07QNmI/p5OFMx41HYdsPBL2/YIpMYY7I+Esw71zzZ/h6kbmyVBv
JBJkAOQ1AxF1ibKggPxbM7BJziQF8b8ZEBSxhOw6yPc1hN8mJY3GMTXcmlUTxmhK453oosrjzd2I
WZM6DD5joI2A4dXg+E6aSvafMltefHEI9hXWfVzb6n+khiJSYWRC3296cnlVZCXhVHvIOGJTU7bI
DsW65vz4ejCVyFeNBlaUak413UPBesbw1w7GTD83J5hfE7B5d9Awv3waCNs2BJtQqUKZJ5667WtP
fOSSwAuvSVVrcTNVoEiXethMGvdHI8dd3DtZ0Ave7U18tmSKR0rENWwhJgAb9YuzFWRpGpk5oRp0
ZHTRqocajImn8dz8+RWaYlGN61pLl3LudYyK4e8DMUTL+yBgSe8C/XBZ8YUStJ2nFnVoQECsaQCO
0JgtP0MZfvgUSDsPf6Fyd5Tn3V+85KXPHYWSSPzAMSggC1ZSgi0O7GF3PXa1nBgWHH9mwy8mYeJG
dqeOI3UFYgW3gaVQ1N7Df6lWl3/qbONlFPIemekMWUCuRUBGTyUN5vWCAxD5qnWsUT+9CBmLR6CI
vafS2Bw9dve3YYF59rEi6qA8bah1z0waJcH+ChFHAJHYWNSlDsHo5drCPG9/xMco6jG6agpf+7e2
IZrAafjkC6WX8wnCQmHI434euXhsGZmteLucpza9chbR75uPW1UBXDnrG3HT3lZK33ukF/zhSkIU
JA6qbZmhk114qx7mEzT6mOhrqCyMMqxh4w+MRRukJfaymOpNm12myDIvClQAFUfkjJay4JbVyOz8
3GzzmVRT1mOYsfk168fuS8thvHEMe6s0UsS+4rQoNUr3SU+oNn4uxmidOgGt0xohwSBsYCj3INPz
g+fTPRy03mw+RkL4GpVQTS7bP4Y/2mGCpOdGLTXM+U+XeFXjTQB0zySukY1DZkbz/5OF8X+/Os2a
RzvI/TxnPAjO9mrAJvRsMrP5QA8bS9tnLMG9InWCDm+aBxM9msAFOtcOa69tGRU7WqsBBMDzZlLM
DwCxIophkf2WHHTyWE3rQcKHfRE00BTkNTeqDvkgZ8LHmXe0yl9wtHEviPdUiPSEBKAFkrleGJHs
HUHDsix0gKy4GFmWqAcNbt+rcy9YR73htffCmsbN6deYFfsYxzw3h2XVPt69XUzVc2ynr3zowl9a
X6Y7J93Zh8pblnhikXuhZev82wG7aAX/qqtchnS2z2zSJAPWa7Iif3mmhD4SfDsN7WvAMdErfqeT
YY90KbPGB/cjclOD3obNMTmZXOt4ie6Aa1RffwkWsNr6Q69RlaeW6v+J+Geo1/tYVgmS5cY6reOT
K5Wy0AT4gNyNTSalIE0O3Rbmwaxwne/bHwWIh4vNxKIr94fRe55qoK9V/ScWX2V2ti6HMhi32iCL
bT9aDhQ/q0WbZmaHBH1qM92oDkfgoJ/a4/Gyq+VhLnqXdq4nZorjyCW0z9dvDiRUSNPdGJgjEW5X
KVklGEgY9PnIX9X9lRim7wfdrP4gry1kzLUKqsU2hSEnvbgDoIYtDg0NdLU5VO3RIa5I4UMUhIpw
20SBP8eAFeVsA05to8/DcdGzaw/83OJ8R+Y7hI2bwZUZnLnBgYkbjJlbuwhT0HG3w18j/wVsGF0s
vkerajFmMNW0lW1pTgCur2zaQQ6iQQy1cyakvVsAY4/JeZ1z/+4u4f9wZ3hxeIOq0CtudZ18C4pD
fvVEgErduemgXdNjNbpTEnfzkMFreut2CARp6N9uE+W1b/7+l9KDPRmtGm/HB3fmmi/SZBgRYvGR
70HQyjZaRLnb0Fni5TmG3FpVdhICrZ+wDvZLS+D2Roo1ZUZbbXB1d2No1rv/ovyeS75GDGK+7fD3
GjrdX5arAzQZ8G/sy6BgCDdbsMBSOfmsavGHOOtQolKlgGxhCxtUfmvNRV8RS6f/i1qRVwv011VU
aMfNL1Nw/QqipoFLkXpM+sN7Jo0nr4PIwoD4DFSyQPEBL9nohtDAfwA5QLfoZCdJItSI8J5Tk7ff
99A8nop+Sf06DrP2Voh4tMTFp7CuILr0xeUViuPALhJRDSJHq6gXt2ja/fBFELHpHSThVcLNU0Py
XB7Z8ksJ/h6Z3rVZPAylJAb1E4TObbNLt1BZ8bn5Invh3i/jCwqU1aUjcfj1RRWVIOA0y8qYZFXB
4rQRNU9ball+JS1rHS/tqAcU8x10g7iIRvVVlNZQdoezQV4ZSuAZB/dl9QaYzqHhU5tChFWnYeZw
zM1mYhQdqKl+sETnlgVEPqtaLDOmoxVHilR9OPPgVSBj/h9oxOvjiHmOL0en1H95pGx3A1EAOX+S
t9gqip0U0QnNQDoh8RT6W5eay9HdaiXOmWYNTQHb88febHxeRXZ+NsU4D4FJz38VnUAbVTkDOUyQ
TzqcalIR2Ok6NcDCKW+6cRo6bzSZFZlf5VBYct98rBrYlJ5JMJonBX2ZgmUH7O6ttNGJBZ2AmfKf
No5Jiy+j78ky51zdcoUq7NuXfGfIu/GUmxU7XS4zIcDISbPoC+kaj8NKTuWpKH9pa/ZSJq9/Q56v
/8GbAvepb99qv96TdAw/YbTSK22UzlyNcZZlRPW1JTJsLXgMYLWKOi9rZWxLv9zRivtOwMAuTTu4
T+ZTfF42kEk7Cu1yoj7BcVBUaCBnQ5ZZ0BdpiuxTDDRbD1a222pK+UI4t/vKFz8tql5qfJbSHatq
qfG6glqHCJo10t2TYqLIwsy3vr3SIT5cZHFN9bF4OEgbNwWLo2gvFff1hoB/VOBZ09OymNbhPU5D
aBDjIINXctOxSPdpXqWde25TChfXKCnYZyYsYlg1aJnK5W/LWYTuu2SBuNBeM4kyZU2mJoEZMsCx
3S71i0ocbhxIvFQX5inDsA0FromSxaZ9/rqsuhddvZr/agM4EWCcJq5NtGIi5mhyhcOA4iVpxfC7
xuMKUQehBT/tF/5NxnCkeOETRE6w5he16u02cMTN83SUEeHQX+4xobp6IGYZ3pTyDVIRXMXKYtLb
mvJr/Q6/lVr04iAFFn9PKKMjzSERY+QXCsDznD1q9wF1WTiWuFy1wRKPkeWFpQSUo2gAZJDIEbOG
pQoDYNXWKIRCVhc6AwDXBszA/nPJ5KvzyH2gapm0Tzd7VIHnPJKHmN96fXhaMNAVdE8H3fGEC28x
6R1R6BMZdpoENZJMorrFfO6t4TKPRFTnKmI9ljyYOFyEkIrtOUVGuPqbR39Zi8/M6RXhIHdPplgl
QoCBY0LEpKNXujvHbMOEHqJK89BIkElr5jBRpR3vBzYUsYX7Rd33GimkgNBK2C6/un145pFAUEcX
BNtcuOiAK42DmUnVRpg2arcBge6LiP/EENSfbATYm8xDplk9o++8LrpgqwDalX9Bcp2dhFRQ1U6l
XlC+XjXSfE+20x1zs5ItWoJASapHpJA4c4VdF5itGAxvIJne24EJPH47bkK2k8699UyT1G5JEsVd
5HWZlzmpyiMEqBKKVbv7n7bYJS8CzkJX4B/4RpqwgHQ3tvjVTvgAgRYfqJr+P8nd3hBygg7aqFGH
E7yUt3FLq7r8AkymyZjYdMuPi3yKPzgJ38gN2lP0D9hzvuHOWK3SEiPiL1a7Eu5dWOpFmHVsb1Sf
PcbX+WN93WQIMuJvvmhZC6yr7sXBsSK018TyDwqzvmiHY2qgbd7IX424twoR31IuJmDyFyuANymj
jLHXwQ3peY90yT35TSagiZcjvgr2LynDQmmpL+OB5U/OftNcu1UHUUykzU82ad8jDuVyiYSLx1im
kVEmmn8mOyJFuxrf4lgWtb4pc/slTxi9juu61+VGMkw25RS+0JsJJPtLZWnIRV6YFtRGvJiEaiIx
bGv2Qyok2Xk1YgiVb7ceWTSDGdvZJHxKmSkcWIsk1fbGz+K8zgfeMk+160et/XY29k0lj1AvaRXn
iOGcjTfctWz0wk+KllwtC8+b5TKP0fgmIBKh2fAXM175sZTut9LzZZa0c84BRGWTZAQn14vm81Et
fXwOVMHOH1dkrWypV4FPZ5D0xAmDHmgGDAtpUfO84PGi7D8N1tcmr7WNRbjTmhDQzzVZvssP8wv5
aJPoivM9fzlt0SYXsdSOai3yPpazwZF4F8HBD24eUH80Xhe4rPGK7lw5t1fX0e5O8QIf9NnZyjWA
5zMV/3cunojfcBUol61AwpZpYgUz2ZsGcLTpQrZeXhM0rDwtz/3v8hyoMIPBxuM+s9DrrDh5ikAM
pjlCLPxJA4oRQN+IoWl+IxKTQi7BPIKXUbWuHWJVP2Hts7o5LlrHKqWwVbvfb19rlWhDMuDDDonv
EruXSK2nDiYgktJswnST8lZLhQbULWpX/zozTYu7u2IR+RUjXtvuCF56lFWWewKSjVd3Sh7ou8qg
UjeLWt4/Ah2wJSa10NlFe1Y1md5XpX+Wd7XLVhSEFyH1Tnyk0UQVQjjfDRmX0H0bvIHaZsYcIIfH
vEkmP7cvwh0YEwODJi9ZDVZ/zkuo/FBacCEJrcrPRjlbKIiilogch1c8U1fBmU4P3UUczFw/6Rlo
juANcqmXs6AXUOzEJaK3UqrhTxWiduNI6g78Qp6ico9XIN9sg5Ugjxn2IEeMpDBUuAyagMoVVDg/
xIj8Q3BZXBlxpUzrbFjnWTZEK0doBS/ZDEifhk4eGLL39zurnwVBFSI3idqLNB6rl614C3wY0iCT
5vS9to1TngtXNOdBNS/MawivBweS/km7SAQck3TQ+WZMtLka6LEjH24b9r83uOXNVSx8EEqV7C+y
HUeaNFDju+I6QDoCOugcdy/EHWa+QXcvzvkjr2+Pdhahnhmk0cWv8lkT2GAphvReOfyL4Fx5rOaX
AunixBbP4PEwCeLCzWT6v7szEmLbbaAkRoFIySSvmGCTEqsFkzGt5Eh5s1lQ36masULgxnJBPEsj
x/5OobpAVfrwIT3YmpbzzD1Q05MvA6dnxMQyt6HF1oOgU6Q1rOX6y/j034mqPboEYmVLEy8CBjFc
qAnjxB7ZHtC1FAu5DS4iXyMsxO7zt8M6nc3IlS6lgXjDRcFMze57hkTz/WDCLGAEbjoIhyyybBRq
oK+QGu8Sjy7OIEdSxcd+bcdtjLpumQln6Ta4mLf9FKVG8Y80CKSoXcg0R6plG0gwmt0S6v8gJjLD
pj2eYh1/2oEw8E2IowsGa5apSGDnFiepXhNtu6AfaD/U35AI6MK6TbP9sIQiqYAZGWUrfx6qe2LU
h9BHRcp9K6xmCo60BKB33h+2uWkHTrRND0rqkH7WZHPh42LHncqPXTKFpCFFKamElqMeyKwA57J+
kXMW7fNBNWQFkmMOua1yy/deAyXAOoRUddPW74Me3PWcnIxxxk/QSVVr+zAa1+u+Eb9TzBckR0jk
j8zaRQrodhejIgvALbMPRFC0HfYn6TNaBF4Sfuy+RnsEU9dsr3SBlkrdwRbz3Fj19PCfZr8rEe3C
s70gIOrFBva/+7YyO+UDRjzJRbJVDB+/petPVN8bSgEY/Q0An5rXgpXhc2MPh5HUNgJ7EqxT8Hrn
hD3GDVjODR0Jl28B/erx00Op958Z4a7r+echhp6jKmt4m8v8Ni7rqjgpAcId38os+krfpBCpJ/xA
VeTWbG9y1diRNziH/ow3xMqxKrs+DZyIVlkwAoX8Pjai8DzblAgXxiotkz5igw0Sj2ZRZofDh5+v
drgSL+gQNkylhXOq9Y0dHukJu3RUINXkT93cMUfpG7Qwzxrm1YYxka0GezVSEEn7nX2MEIaW27iJ
V3rb7myqpfeVWC2FI2XPsXI+NIzJKMwt/3PoJ4yQ8UOLh2rts18LxGXmKW+aHzZO4p196i/BkHh5
Xruvc8mHTyp8Fr0bmdMaKxEiOcx91pN0yUNzKH/O/kyKVshRIGTyM261EETHCHV+htpnPdPgnU8C
5YmNZTj6SuxOC4KVC4/Zyao1cfEESIAuiRzdlfvQXG2xdTD6mCuIHZO1t7hWlR2K/EZx8/gCyGED
I4FviYecTmPjDcSSTir0QG66fX/fFeLU7S0eOB4FIIWpFBqT8Nx49hg6mvVRwMJrvltAzd5CbUy3
5OBkgbeuUcazYFn4JpFXmG5xur3Rz2I7kyadFRUlDdPliHdqE6O7kCNHDz/fGQHYjJN0JrNZzNbM
H15CNsyPU4H5vo22sRzPNBjWZMt7eSjutHERmxr7NMPJwF79PdfB04BO/31JIjT0LdU4OE0zAzs6
kbhYZZA+o4z8DQOtVYzzd6W7DSWnH6ZLuFnCQY1LHNtY04trF2DyVf/Fs3f3NF6w+rLDOMnXegxu
H37a51m3vr1o0aPEpKBbsQPRCFV0kFBK7g3OVFLOdY2HTaQ6AFoU9pypAP7DmZ+i7zYFnkf6MV/d
pjmP4OVCjIDDFcChrZN5+NaCUq0sVYNCVwBKMu+5FUwb7Ff+1Q6FXDcDoisTaSkX74jopk0woMSF
FcW/o/q1cgIwb+aWTpX3jFoe3h35JPO0LcnxaEyVyz2XDtzZL4ciiMcsuCQZaYr0wPXv3my+iSVn
LjTnDLfHtnIkoA3dibDoOUumsbtWSMcsQl9o7ER25RBIYNeRphpoUs1qxGJeFJOMh4iMuffFNZhp
543Tlq9du+RkL1j6I/sB5XwWignY8xozLbUDiiXIqZGpER6GRvUISrV7CYv09bEduK2nYjur1EcU
9rU75xehWRHanrmqMrbaOMkvrhY0kP7mvFYcyZsZEDlypiCnuyFSKfuyBQ6ccFXxe7o6h3T7uLnZ
1A6kktPnnS8kEHerH21GhRfdZIg7BWXbFAVj0n3Cf1fJEJZVCg+eqpeHvt+hDTSTXlg9ZzoiTKfE
W4bBND3LkaGFLROMk0p+ZaFR4bRp5r0pMUc8MyIQH8TXsK9d5Okm5+IML5JtVQFDSAohZID75tPb
FEp/9lbMFe39S5yuDvCeXX/cJbseCDfgAcS3RyTYDNqKnTh2j8/ARuOEfgwyssItvnj80Dw16hjJ
bi8Y+/2CZBnNwgiJ9MuifV7bNI3f8jn4nIg3plrAXgabwp5Pqhe1UG1yIPWGMTktk71WbpykDfUW
HUsNC18DMo1iJFKncjxtRKn+4IjMmOJ04su8ugPuIUJVg7nP0DQOtt69alSA0aQqrObx4omvkYok
sCzsX/dIrzl6RJyYMSUV0oG8UuV4yZw09ehGDUIKULQc5j06BYnCgV5Jm1uYRB8zmNYrCtEx/dg/
myD7AjeEhchh4aeer7GPfLL0vXyH2HkInZ24c5mJe0cGaIardV6Siek2L/g15OsHIZpIFwPwH+oN
xwKx+9o0Kd2K9u3Ca99eyXp5ec+3dnwX3lzKS1sRfXhO2migcucQRN9vzg8W29dfa5JNUc+G5d9/
wZEKnMhSNP5fYvhT0U/x11wZ/kJ9AdRblyTT9mVKrTgFRwh3QiKFQBnzX9ZdzThyLvVHhYspMMmi
Ogtv+Pqy34Vv7Bexk0HcgdPCjJfBjTUgo8sIQqz0JfbmNrTROltXtkXeadbwTTjzp1/gNuaUEICh
iaqJXR16rJedQfqRSSYRM6vOlIFpqm7DeazwJw2kJiuoVYQCiArqc7ojULSQ9pWd/LxG4hmQv8ZR
OfF0zCR1EO1qiE71EXsChK67lbCzfF6ntWry6/LRbKiOQs4A5mMF8yeItmM58wzvTTTg4JZ6r7fp
vKOe0mg734ImMXWGs7Yn4VNSsxHjArOwDBkg/MKzCcnIXV7h4gzVWml2at+r+fNVipyDrhdnFOBk
K5Tb733b3gHvMHBIYYzTRTymfuHdC6GvFPyxj90mODuElBJf5tZFdv9mhTfQ+dQfQ3xXiM4KBqo8
eE6RrxCGU2Ngts0QQK2GvDvTJcz4GvFA0dJ4RZHeJ3WhEzY7pcNXY/kQvQRheM0MMK0sfq74KxUU
flGIVqtW2hqlDhhp3EVydld0EEBQrZgRKhhr1GdPn1kstIXEf7GXIfK9G310Ku0sCdI5gXkjr5Bj
iGi+/a8H301cF7wfsjL5oGQmu2VUyTL+LNiounYQQT3KWmEh9XYBFVksAdnD45Y8U641NV/s8vDF
lkgYjmCUJsKUf572kUChRDLj/iDAFoRBNpflG+AR2Ewh/GYh58WwAFY/Eje/0oYNgxd2HJeHzTHk
bXaZ0ONeowOkgrwV7u+SVTqWM4t3rSqXGbdP7vIOTJopqTPPNodrraoJUNtNaO3E52LZxp3nSBR5
vukuWf2VWEI2P2ABURdnzYVvgugvtLgrgCCGNVu6NyBSabkMiFaIvGWJhWZSZRmR+Um9yyo1YX8n
xn2b7qbnqRFEtuNkopxJ0i7DS4S7OyZQhy4PoOnL/c2E3ud82y98kLPNfv0D+d7OGkzcCwAtZjCC
cHMOGH/Q2xz/Xbu/g8H0lYVHihfvaRb4yABG257eZlCs7WLApkWMv+iEthUMZ+QcU8LwYTwmM53a
3duoh4vTMeBb336t1E/ex6o3Sy89ikICHYq0Kt9aKBM6jygMrnRCT4RGsyfd8ptrsjTiSkuJL6Bg
dbXTh/U5m0w3cLTqz6hFpYUVKwluhhJ1sREDBZYWrnhkzdxu0hp2iKh6A9z8TrIa1Frdzn5vTMpX
Tf8Vhm8xRfzhKYGS1uyFDYPmXcRTSLJae/OUjO4/YuSQMJyb+G2Oo/0n4E1TBUIz6/f7vGbkK2kh
HGfQ4csBej9qFKsXfCLMe3rIOs+vLzbu5e+a4gLyu5749I5k+xen9qKcOci09TeRpy+1XfGIFLX4
tMFnLcd2uYqSj4uWBhgFNwYAa43DyFHNuvwuU8dEg/oj44++KAyDVAoMYZJ/Ce3dpYYxotpm+gSK
JZZfRHTXez6mCRAnDBWKdAlbCPQf5YS0S6bHGdxpddD0NsZ78KNEtKSz22by2PrS+p6ykEFcIZSK
Sv9ZAzfI0NutMwBzvKdW2pVvI99gSYd2yIcu4/S8oewXmJSYWxChqHZ7x1n+6ZJqt6biqKEYrssi
3bZKuJEWy88+Fq7nA+TKr8sGLW7OaNzuh0BARt20Od+2JO6/39Xzo/LyzqlWMxqAlwK/M1rOJkTe
8u9Zya5sT3HQZE7XLlNY/NgwLMfsOiNFAjb8bjDzLFbbTswVDs4fAGPZqcQwxp6ev6iHBaQ5FxGU
qcnNFqSQloCttM38mtyfcjWXH3I0HilYesojmaBD2CyeP9nEn1BhvKayI9f89MutkvYJX4N15D7u
QnEO9eS0duhSkFE200r1gckb9I2x1GEWyyT+A3hGdNfLme+haEVKJv9ZO0grvGg0osdg+HZBsbJY
JW1R1IOEFIVYkVJjQrkgNZHkfpkiIB7qcwLw4VzDqj/JPQP0F6AAz6K3HC9zLuR/Bpb4PnydULmP
Zo3z2BtHWdmumA79Y65F8wx0s7+wJKwBhzZBZCyU4ElP9zarfh5hdfRZx9Ov0ZPO2s+lkhqScf/b
iznuXq5v++tf+goyDRRL+FRioNbhbIgX3IqzwrgXzoAHlWURFsO4msIjQ7PqYFMG2CyqWpzXHKv4
Mi6bYwBKxvUKAga5G6TUpUL52OPdiHZnGWdk4PqUJZIsvuuRZ+OHF4ERlbta2l1C3/Vu8i2YrFzr
3XcVhrqvT13eMThJoeomYhmGKc2kH1EjZccD9rKTAZ9nyGpDkK1zG2RzMamfbGek/TP9io822ncU
4j8gfZX1uVeXbdV1/88hWFnrrE2Y3BTPZawQIuL87jw4mbdHzXDM9IzhrSigBMurA8d0OjqHcGtp
UeKIkLwrh41W8rlJ2CXwrM2B3Vg490fabj8uQ+70CHzMWDVQWXppypFtUEwEFMboaa8TDmr9pH9H
FB7RHFO8xxdn6SxBsyK3j6CdAzWhtL/cO5Mt5usxqGAs9Zyh3Rdsm1lqn6uoOJWLcuA1RFbnAwIV
JSM58JzBzRXbtXEoJsDW3NwPeFdHZpHvv7w5+NfE4B6OJfSCzZTz9vwDEzMhggm3PzfZcHyxRvYg
H9IzIWWxw6cIgbw/UxLjx52ds0LuKwxJMYDO2EB7c4xIxAzqXWKPUTGB2lAsWpKM6AcLFqNzQaiL
w36xsxhFotLEY1FZtNiKPXccsB5mp+xlR863XYi8aHVFBHFJurwdWalr16RVrZpS42EXz26JxPm0
IcEXonH9xGookNc0Byz/1hCEB+W+RGK4W9bhwLYHEbuaZgMo87JWNT1y2QBSOETVw9a3vBuH2NMf
+pkCCM3zxiNIMQ0qGj1ccqZvwmmmQ1EJTw7doNEB1/djqK0L+MnV4tjgMhmiFq2yupOdnbfAmwI3
vvzjUC2fTbje1zjYyInpcoq0U5HPP8OgCb4W2E3tsJCF/RqwQo1aQ7/CWhah+KPklFmXSw3/Hgcy
cz7Y0UNb8MsUwGy8L0vo7rJCYVFvLjR+GEP3aBjDIiaGifBIA7zRPwODpc9hC58HZYTYQpqIpCmx
giDnoeGd4kTK+7VQ2ykCHoRKxGh6Evyufu9I16m+9ebVunx4nByIBFVhTECnJ3Ldz8Gt5msB1oWR
2aX150u31C/tVPKkMbNs22DXrEc4BPzZncnTLV25Iq4Vw0dTPXA5KWEsKBqGNCk7K6dw03aSMFv0
inRDCEXySK6PbkCNyB21ov44X8TKq8ebjY8xc8rAyVNd6K6JIfobgkizQNAc44Cvgtp67XVYkIM8
OlvKSxR1WzxW+EdzAFHFSnAIUIY7Q3+JxSGu6rIYAHulJQ6f3MB/8XCOo1BW+9l3D2wbQmxbt/G6
T9On2ajUyEdxANKxuVn2TniLYA8ukR2YbpIIHQUba0wk6FUw+0i+E+l/YYjWcS49gQnd4Xq9lzwl
tvy1t3Xv/uUE1O3IE2uUMrJQtmPqnXIYwDbUVz2IiOCOtjcyzxY6vfvUckMgId3QQ03tetxi97rU
qWjIbQa3AFvoYl4gZ6OEEqzYAEFzl8vzbCoQDwsra9MHtIhksPOGIwhjkV08hLlK2e3JrlvHuA5x
hwIca15OgL3Ql0V5HphrJRhmUH2y9vas60KvqlGUGBQoMFL1u/5DHfkCVyCJMQagKy4lFFxI+83a
DPMSNEsHPlBX308Bvfqht/mrQ7i0XjP4WJf/DjjbD+h7b+r+ITNITzOV3fLEQCIwZnDvu8kKsgzA
+nS0Joskvh7dM4gvslsmB+7b8el7loGueJ03QNriPdEeSGymJ/zaU/GM6mKAkMl1pl+LoATW6kRP
GQjYVl1G3QB1aqvc1vqAKB/+pRgF0A1xUvI0oqh85b+3cT4pT9+6qG/mpDpgMTgFOAR3Le0m+Do3
nnuhslZLT1vzGTCAVp7/qYMYz73KnaiLXdXZ45DwxbeZ9fTvGBSSPErAU0JLRq69vSC78zNvThlA
GvTX/tRgeS6OxKtTFkHIG0H0kZpPCMgdeWCtreoUTIdxiRHIih5+mvNUDfSWFUBVjVTZ0qSu8fH2
yqV6jHJSEZpuuzT3aoT2TjIlJkEEE0EGJbCD4xqFoz9ckXnPo3DqOjhmNBnTd9vbH09/AQgS9TgJ
ZHG8zcWZx9oZmWAxyCbBueziyGZ31QNCWzMc+C21ycTu3R4KoNr87gqggSTU2IA1U3cVwHTT5bfL
z1N/sneGs+kKrTbwy89E3gEdWCXZuD5pyo3azbS319bjQN+1gJxbzd3SCIJF3soGIx2VGBffV9fl
JX430+usQqTE8xKn/EyiMw66pa2GvILI1S42WpnOsOTacsiwIYWblsv+4btAL6kgYJdkw5oLJgSW
HC5ck/MV8JaCAeVVvhudTVhlySPz0ei1odyuR1Rv5B7XqbMk8UXz/uLCmlYVe6zhECuIZSRyhCJb
jW+xz9Jckh1JDNv77U6ChCC9GATlGSk9i9Vg+/u9/5E/b13ZdfmPiqfdMctAZALYZ/H6kdFwOFHv
AIrd6jUCubIemicuj775ZFh++a77Wi6uFr8O/lStlofTZBbneEj/EfJTBLNB65ILkw8+zMBaWC5l
SkHADuMayBFhs5m0jfn9YknBxprY4Yx0CnCB5x0dIpHQCYa2x0yONfoMVPSY1v3RjkwnZMTvWHZJ
OEsdsIQH1rqpvmwr3lHUderkDZYPKIImrm74BHcVodEL5o6ip7czsLPzJUM+qNkw9pEOQtiP10u+
/w/liBT5BHkL3dDXAOEliGCDVHacOiXRWO4/8dchGjTxifpsiVRhRdba4YOTH8DydnGgQi5cKAiI
KLQYDBSrLPA1mPpcq/6CZWEHx4VhMoA2ETjYmvmTVUSn0rmeYnKflrjlVzh8ho/acSir5IwVnTZt
tdAN0x+AJMplPkcgEqWbDAehfNPdoh/HbJOldE5OzhUhMohlmy9g33XPHa3tFW6+WQnaMiPLSr9q
RhjQAady+b+MROg+PJmBuNZvu6mj2V6rCkKpwp8Rtfur33KaKEeHrlI4k9N5QLk34Q0YD9Zt3cJv
b1oUjV4su5uu+ZA7+ZB9lNE7KzyK67gl0oxuT43tHHHGF/pK9mu5X/BrImojxttxcfWF47lgaWVO
PVt2lBOQ8Zo76RR2LQAkzD2CckCRbfdZ9Lg5dtcfIy7KJGtf5IWWiprzg08M5sRM71wgobMiXwdM
OGmABO1fFiqy6u4Um1O0f8VVziBB3Fdg/AKL5AC4umtD5ff/RHgt3uBCHMaeutR+zsBXksZeLR/H
oYYeuIVIFZ5FJXXDrJnOLJuXm46gQ5b9TrxwoXvlq6rWJjfmsLV6C1tLvBwun2+UGHCny8HSYRZv
8zg9xRMBXdPKszy7gjpH4ww8RxpA15qudxqi7oop2KOow/Cy6BwXgKDJGSdiInwtVNe9uToRPrIN
SiWNAZRnVTWPOoU9rC24h7yDRyuqJlZ11wfHQ6KYcINfYcYXkb0HlcdbuExScpnDuSfKdCCoq0Ge
Hv1nSa4rD+KekfX2LyTfp3vtopyEW/MTtDGY4Zwxnq5kfHCHjhQNyrfmScXL8rZ1x61P2eZxciJP
K7fVFoszNaPOHZx+sF1tjLsJCEvkF01lqrIMR4dEnIucp3Ko9IRrG4Vn6FUqI57z+Xza7+LehIKw
7ebCoh6HuhkfuZoSiKPKHMt6cpICuVUpAI5SGPQXnnMZpkH2wFY8IWTLVjHF3DuCwaCHWt9w+rWH
+NsNqwVMALPDoEo9p7jpzEbslnCJAYkSGmoc3qWj4VBeS0CvVZuRl6eKyB+7KVUxA2w0bxHJPUaj
lhtDR2LUZyMsRdekhX+BST5IGp2Npcotx5/2LCStgXoPlkps2t2NXIABBOjyDbeN4ZIohhQiAEqU
YqCf+gIJNu7/c6oxHnbg+vW3LfAKIMAWIZKBfzq9Qpz4P+4xhwfOgZT1jxwmF13HRU597xcpCqqV
dlRRST7DyMddkznvgPv467aRMsxwM9Yam+MldpokKQZFLuw4lzCQxjvWz/RC9aKedNXf/jdbgpxc
Izja9cHbmvXsT8TkwhcRXViZnFeApUDS/qHJhjPM9FvMymI/F6iQ+rhU9dz2VNeDh8yFywmawjwV
8FzrtO7zBQdB5mFjwoYhi8Nc6cwYCaVZC1+b1kpmiPKfXAyWJUkPfJ4U4N/qYv/e+EO7DSRFUXtf
EgZF5k/UbBv14TkOnclyvypqwDP14QgOgW4sVreiGeerp7vnuFmjm/Xgb0Q8drnqkSaYVy96IiC3
AQUCza7SahCH56pk0KLVAiSf5VcDi2c7woc1aPddGccGzZzpZaZNU/B7Rk1eWRbMyZqCBJwf4X8Y
kfxV8v+VH/IvEEdeFo6OFa4LMMe4O3uy3VHgPb/bZCcO5eM0gTM8EQSmZ4xJwNxP7+i5GS05PWJd
wmPGblvxnXus46+2zx+bEHrGx9RTPprsBRYCydgC4RxYtmPoK3KHa4fyb80p3WBffHH3DTpAAW6q
2RsTXx9slXsIBexkYtjAY/XqRVUeZNLhaaUZzmn4/6QJ4tDlnCdfyONAgI/9KvSvp5pqEVZNe+Wd
vlJ/fz4yN4e2RikGkFaNQe1ZtgY2CpbJdsA9lvdzEGpjwHBdrG27Srmuo2NT2o667tZJNvrutKOC
hfekrRRVIPkwanvfaP2jmjzUAVC4028NFqi+WUU4XZGE0KJIBmuq0e+BM7eN3yakpjNcpuKRIR25
0LRhfX5H+xLgPH47C7y/h8K+j5vdCQqtRRxx7kZIzsq7xR239ibqnXUIuKlMOkm1TnmiLJ314G6T
6XF8mXtM5URsuTV7SwRiTXP8J18c1sEJ74P5ZqLASgGJu/P2g2quAwz2DgD6V7NlI5WtAFuwYlAx
o4uc3N353aRQkD08p7C7w+F4NHmAGLo40ESA0CYedA5CBTW15KWVJ5hJ4YCx1HD5CTWoGXKvM+0G
KG21teNM+EFhfAeJmgXfusHv6N10OpmNpKoXmTZBuqHYOZboXzR9czPJkisZLnDgCkyROyWnvM/u
gUfKqTURMbmngj/+0WlSIv5pPIoxgw8i9yTk/Zf/nXoZftsblXTlQScEDFVf/hbMLVob71/T8wNG
U+98dnSxe/FGITWJSrU6t9ms4elndsFmDt9h24QyBticuGDCDh0l9+tZJboNUsZZ4981Qtj+qrz0
Rc5jj4FbvflNjVWqAMdtklzi3yKAI+y6KgRj5FAmHaopF/Kra3i3YN10FPhBN+oWH9WuLcdoglsB
RX23h4YGvaoOPdY00HceuHb8u0TdbhM8iqTgJpODOpumYyNKFE7jq2NyOJi7z5LtYYvE7yBKx3tL
xLr4cs6LrHkJkG1ryRYOLDOw8yBZ7jJAd40SKHj8dKrhhD8aGGdE/vUD4QSA6m2PP+9F/EimKvHi
sW+DNxwtLlEZ1ecrPR8nXpZgSyv3KeJnaxWfAxdQtzFLtZo8tRksGs+1wuspsttliAu8Lay1mgK0
4LO73GdrV4k+Z8j1XLz9/65NbkjPSDLTI0cNZ1z6xvXe8VrXJgj32cIsAjeupiHEv7GQTfVbqwLD
5L3t2qsgKcrj0nBCz5UTLbgnZJ50wCvh2c85jWKZ0kjQHLshwoY7Wjkv1bxJQpdgvSN4z78oOauX
s1VxKkEnq/CEBK+8pZoyzHZKXECP+qGxYv0Y7HnTuy6VHoTlHyENBeI0sFql4Fj0MsAsx7zvUFh1
VcrTXR6Gg8pR8zTWKcSctoTgWsZeAZtknF19W4Gtnz7udAiw3q6rWnCHSTKYWHnXyWi5c7+toRrF
QmC3w4uMydkdOve7DzTg/1d+oyKtl5ubAwGtCiemeMlA+cWP1RYhIw8iIemULeTCu+BjIaQC+AQ9
9FUkfofB7xxJ/RVX+0NoQ45AgaVHM2zxGsE4OdMOdZXkg7nGjyB9J7eHfNYggc0SIvn3rEbQP2uu
Zs96rSO4yTCKEHbhvj+/HmAez/3VvvwrPF5P3r/DHhdq1Cd0vyawRBnak1GgoSJA3fosR0Uw2FsI
XmUqLohwaVu2uwU3i7nhta5A+K4TY8GEZOjt9vPyPoCZlDG+fVENIAYC1ozIBTX9xxpJWwgLbdEu
oBhTyNsHXq4k4rm5IC6anZeTLnhZhA8oKaxI1pdwNzbHlaCEr0jdokYLzb/d99mAaQYGqpXMCmy1
oOX+8/kRDXEOJw2xjz6xR7gXAyjUJbQNHjtSj9WLU/BJvau+nKJGrGSykdrXTy2McGnT7G9VcdY3
bDaQlESrcXxGKWQyFdxmacaxso8VorWZnE72w/o4KD8iPnNbGhrhv5EsBvsCRQEeUNyubB9j3q1Y
8EV0UK+/enX7MX5YlxkxLa4C4+3+MFW9wHNzwkHSpETUbyjEj+4GcmGibyAMGM6QJazOazZ2yI9M
W4yxThozpKBoT+8EAty2knndkb2ymHH9/QmjG3eDt7esqDJ3Usojmo5e6F6c21IfrZUeJX+0bNIy
H5NZVfVtPe/L8zPxwQI3VgEuZT8zpS2gUBUtP7urBUqgJYRJL5Mkkbibx6lmiwLz3v0GFczJHS/C
2C9fPyINe0t+A30MTTG8sfQsE4tmhtK93UHIB6JldYEaNIraWrUD8tpYCA5vAs/X7/ckwWnVvCed
Rz1SdrbqDcgcU88A+pJAuIvrEWiexBhCzbzad9kmUNSOGhaApcOcGGTPl1pYTmbgdOZSVGZYPOJV
knPKwWZWzupVbXk5I1zHhrJVDGRMM2QgozSdN8RXOm4zarPUWbq59VPPiY5dk6IgbVFTWPEQM8yZ
QnRi/DGTWl7WzpjeJKmZu+pdJ/tC2NKFd1ZpvQyYWPFlY07xLxQWs2GO5f8YuId593xJVKxq7Sa6
3VJPbwFZq8P/HHmR/YD7Vgu3D28ucxlCSy4pBUzQoovqUIX1Ikr7ka7vPJkgIavfyJdZUKyf4FG4
zgchHCeei1cF1XrbG9gSyRFmIffMBOA0+xxn+EcFnOB1/0XkFJRkyPrhUQHtaJDWJn3z2aRZw32y
v0qQ2AlFy+s7KcidZELYT/0OMBe0nEwQ1ovZo7kUNDTrA4BegRa3cp1N3UgQXtU6nwUuDJBQnPo2
7Mapw7jEp64FN39luC83S09JcRgxX0XpkbKUS/xDMlwofC/KRBlpPY+Hplp2zcntbkuET0giuHtv
dHRduqJzV+kHHnckzVrzz4U2sDCjAXB1HHTAGulrutvJjWvEk+rMxHhVAxtmlyGP9jkcmoOsKGwF
2FhJN8chRTE9K+MWniNSRwt+clnZAqBPn3QDXFy8mE5XWTpSCsqUf8NHYwYiNs0goXn2UOHOdcvK
QnP4VtKdBBopVefr7uk8CSZ88+67Tslo1xYT4O58I80A5FPO33HGvLDla2f79fXj5hjGgaakUMv0
KO0I2EboHwpR86HPBbAjYrpUGWvv7SQ//RppZcANMUMBDv+noMKtDO5dI7s8nYR4UkL/jkI3IGWt
ih/Wj35Asye8RAnfyo4MT+vagsqq2i9qo6Ud5FhcRNtoIWNJGkXH2TSbt/5LAIMJhM/pUI5I4dzo
FhNqIIXhI7aDzlAXG0VdnKNo7Is7j/eIYFFTyD558df5BpUTmJy0cP+ylcZX47dzAYRCdkHupUQ+
u3NlZMAokHQLfLe2yZ/FBdgHUMSCQf0v5PVjB42mxzHu3E3dZhbq3OUWXssX1EaFRUMyjMO5nZhI
GJ8h8mvmUZ4PJ86qSF7iHggxOAezWGbJ4JZw4I1TauvvC4feSIQdQMaE6lN3KnjefR9nrxjTbEc+
kTJOVENeyuEDEcNuQVqjrJnHy1mEDK2VTsxWBtQSRyNxIvDOEEGZ48nFVNSmV1QPlBgeMUMCZJPt
WoUn1gYGWFwtPrgrNhViUDLXdgJ8JFhoW6Wy8CgshPVUoMis2ldw3xoxU1g6IWCIhl1crze+UK9A
ykaBhqBjT1n5pZgPzL00SN27rQWTFlxBqOz+D763ahJ7hG0V3ofVY73Bw08C+kPAngikLijbuiD5
ze7D1AtNKYui0tU9kTd76ID7x0jljB0RFg7psLDbpovLUaWYQXYMG1gjBRAdf8EL14VphCMsdGPT
gt/SC7J0nXL6lYWRUrj0u0cyHUbb1Vz9rt5ruEcKd94ldql2+jZ81Ta+fiB9Ypk3ljwFOSzA6Z/B
xdTvLsNSi627vUorRb2YaehM6kUPJW3r3n6lJwpvo6oQXJZbuLLj/bixTygR89aig7tYyS9UXmDZ
SkjlcaIwGFKXC6EF+gTdqM9IvSZUcCLpY1qfse0d1S5k024YLG4FAGx+FNI0bpG5qGboF17bAVxL
mXF7ir/jEgXRp1Z2/hS80TVKHCn0bf+VG6s63v0YzIMwXSrB/RTOECy/XVRpOHz1k+hddVpW1R8c
e93sHgffEp9kb64iSLcnFT/+33TtWP/FJZJHUhlFAEbbaA4OUfyFPs5y/zKvYVaLOxL0L5IFI8Ed
rfFK30c9jYrCFjU/T6vaD/uuDghoZ4l8BTwCLXn7RZ5gqXQu7iX6ellci224idVpMBFi6+ZpEVqT
p0ZWLjDeunL/iyPMk/kDzelf404YZJS6r6kEX47pWxxcbyyAokMsSo3eVTwExQ7+Y5j8Qs7lGPAV
ELtD5N6GxVALubWg43w8dgUzG7Pel2BK5KaDqfrt7BoLnBgNmo0i/iAadJg4ooUDuHoXgwGzzJG6
8wXerNZpJA95nKcWLKVmReBGxpA4/0xo/lk+hHVY6vgqUoeQ46TLYizJrmwYdC9HF2NOWBTxF7Eu
xx/CKHoZbVB9B3D4/nSbXWi+p9rUIviEhc+D0LSmbKLKqW2aSkhhiZycyf5o/mWDi0Yovl9hOEQg
BPAAylM2C7lVVm+4tQl8fiYLHFC8PWSOzz0ERpV/tn3JLkahlXljw5TXVe3G5fr9yHJC53ojQH16
LG43f1EZCqF2FX/4B6Pamm0uW3ZSZSqOXAS5NGxSRRCWKwy/FlShxv35YWh9y0ORW+OECWrCUvNG
bySlqqdRn58jAn/J5AYucrNc4BOqShgoiVpWFpBkmUrzMGfv7Oe7Y5DIdvGvAzAP7/SFPituhEE3
n7nBs2vqXI7pNp3sQfENOr1fNgBTHjN+kL426g4r52Ou+LKcb2UUNHflqKvbiXQUtPbw/we/0ulD
o62bAWymudnvfvA6EX0edfk58PBU+Ng+k4MVbiLEENElMEjB6qkz2zos/Di2Gj3P+pD9nuySPt8l
gD2AhKxRJ+Rvqxk83XgeKJcwCayV+2W8zWdD8pp/AQcOkhpIQ01ZdhjHy2Y38T1TGPwQ9qaILA9C
MiQzUlIRTT8hS/A0yJ/R23R3dZtfVueQ5W4+rV+izT0Z2cf7eSAl3nBvlhXTqJa/vqxVQ4913jim
kVyNmlsrFfO/XCcKn0IMwDfo8cneo8CF/Ud/SkeHQKHlEIp8cGotftUS8yEw66darIWHG9Nqe0zq
5ebcGVbGNGgCpzZTMvHYLG2y+64nvG3wbID14WTZEUklME/kbd4gaY5V5jcZ+Tebt++p2a3VUxG4
egxDbhaQ5c9GjeIha57H2P653iHVowPMx9w9h3w1DC4XjRsBUFxonx/02wNkqnmpsuGbcJshlftd
YLDpFs5xXiv0NHAlId54reTjeAysNX9z5st8zbs2KHIF4NyGlsPbqAlK3HD2nKbSlrtqZpR00gq6
7U5lbG+0vCGOV7j/3G52BuLtZhbOH4d3rUYssRwoYAeQsCUH7lMkqxEVrnEgqXKtHGO/zH76mBZ3
xc41fj9iV4zaXWVZ4TviU7nYStGlERlWebAkPxam6RFzz/VVRkmX90Q0/921AH5ylvA8ggcWQFm7
jYqPr2nTH2sz6PKhzUzVtbmAhTJsB7aRO2QcQYgrFERTDsHrakW3GbaRgwU4IvJBt/LoiCrKxUvY
nZuuuht9QKn/tN5oV9H/Ea/NYLJkDkq25XEormcZG7rBDEwOow/Oy2RiW2wL4yxEcUh6/s7/RJP+
/Z5qN4ptWUjjOOILtXqScN/j+V9DL2VxNCcQR+rpP8AHJJp+P5Up2OvuqaEwGg2AJ8J524up9Soq
7ecORNCiseS5W0EVvtVJJxl2yyqiEsPdJdcOx41qHJ8kKg0nla30Ke18EXw79cOzQfRTsiJAspMk
3hVIjFEnE9mRiwPns2goNgpS/lYnzu5S7dfb7KPwQJG74W2NQOv1Yb1vOydSOAD+2bFPheWz5Wdf
0FfvaWnlnYr9zsygiZNeCTWP5JBjq6MBS4A9abnPADgpfMdBhQLI+NCsHvISildyQ2aNgabISUjP
k8GpD6gHG0iwEmCB7GgxCwQDB5JCBkLNIF5Zj5ZRRSFaNvbNfRmYaH3gXk4olW5zB86Q9p4CfIA4
xyeTyCNpfXOu33bi7uCwomTcH1YqnbwPw+kP1MQdzMX4npt+6vuY206KXcaytL5BGaBKIwApq4RB
9s2ysC7aj/55ZHn2rr2vBw8qYszaQUYtQEAPxNhw8lUZJwtTlwS9jFcUsoHp+VNODPbZ1cNHtPtV
Vequbxh59zijxF0EM2Bnld50/a3j9mvL876Fh/fSCiZOKKZZHsxfa7bd/JD4kORMaMOEr5G/Ptuq
43iYaWTmhDpbqOgzmaLZrwWEOzUm+rtFJFugRy4VZoVAdBgG7LhHBAocrkKgOtoIMZolW4dibu8X
J2Hr9wzRpHCh0q40sTciJ4b/Rx1N6dKSXkZaXHezYyr5lO5n6u4Xbya5FYR/wmEPpQSdpz/6G7H6
+8WdwrvwtRjvGvUOtUhHULWidxbroRfmkuna4xr7rAAYn2E2BFS3EvagLbpdDyZWkvZvPKAYtxa9
4w795JAPhaaJ29ZsTSWGMZDw80Qvgw6AEjRUciK1KEEDr9Vt/HIlICjr6+sqRR7stFn7cbKWc+8O
knXCS9HDdnwKDaJQENdhYognIH7Eu0YwifTdHFYLoxj8RR8U2Ni0FRUejgrZE2SxId665TIHTj6O
GuGtk0YhC0KI4WTnxAMMzEN1mFIheXMYNMDPU4jqI8UxrdPYe+15IZ4NjOk6hiVmxesx9I5IJzLb
9kpab8pYv0OKBSU7Ld/f1VkeTN7M+GUGygIL+s04w/iU3/C9784RrouHWzmJJceMq0jK23ZcBvPf
0b40nsIf+WLWrGOc6Cgk5P3XjtF2Eit6RVH7cZCaqO/hOK5I9deiOTUf8XesX52Eh+qFWZh2nmO4
sXCn8W+mJt63+yqoQHeRaG1rOy0uyxdnaLVSUl5oVl+mqQTtzMGVZTyD2iur1+/8Z2KMk0I4w2he
+rEEVYcCt2r+j1wwpZVawaBTXtlKZhy891Al52NjM7caRXtDbCNLD5VplTm1f1Hz7ZOrn5bomL3i
Gb6SxTo7V6fCZlEkEjgW+Qj0MMxgc8MfbZbgKIni7VmViUYdRjWBehKZrSL7BaINDagwA7A+mrUx
vD0lV5P3AOUw/y43ItrQQGR30JjeAttRa8d9WslEflYjpCwwlM5bNsLo8R0d495uiaUQYYJxXCBz
2+Hehno5H0zm94k0k6/QYj/H8jthknLp1L+px9v1VhIXJtwhBIMb0nW9Px4chPp3YiC6LBPbVy6d
fhZpZHXzaT2TZ0dnEt1+A1Xckq+LaSF3sy2+B8OfpzkaCTh10HYFlokMKkMhpoP/NJ7mT70Pf5fo
HO0ISgiE8LKV84p7baDtweRi1fsjq9AnjTyRpUkdKUpbdvP+OAe6/5WSWTPY8ksbyJsskUUT4+JH
U6N9FUWvqxSTu+Vo/xdVqD7pSeOIWlBoynqBaOYjc1fE4tTEqh75UPJ3LUWjN811xC5lQaKzB53N
xH7uiXNQ/yex3LBOmdDCDyj/baq1zTm4CoH3JpFqukLPFsqDGt9vUUZpduCONGlveIAk+XWK7f8u
K0qktYYhvbnxUxORcJ4lTBh7NuSliI2Qu2ClqZxalF3Vm96Kp9eClZFq6SLv661N5d8JG4fBDbND
CHpk4HyZUyTDQkFoZ3ARJFrwchjbDDgiAYWzNTVtaCS2He8au7uP3+h6o9JYjmAw8wbiIB/RX3kP
H4gJQQk5xa03PfSI4jKiU5E/OzEuG8XfYSXnZt+O6zhf7wYBHrbI+yl0vsWNFnm3u8YMQtHd6biy
GwgkBbBN4YibJtoQoPmmOrBNJ0X2xsOlW4t+ZQB519BMs3qCXAyFeQprbjumnh15h5nH+bH0wXwA
OJV5HnB1ve1r35qKIA1JifrqBLvZ3nbVujnD0lf4ZdsZHRCzVqoPTrQkFjE1bO0Tpp/glQaveHGt
C3szK8KmAFXCcRwYfgM4eAfZtyyF9Vje2Exs3eDK838dGORYQEQAWWH1RhCbdSSOYMlCo9C/Zvv+
QVHBf1pGKr/b2jTqly1ujiUzJTTK4QvJTEsa5boGIAIq11uscNrfc+G+Pb4DIsvCpK8RdCH8n7ho
c4viZ1j3zN6FR/50KKiZTUA6SM/nsM0VZTVZNOvMIcW+bUSEYDWOnu8NuBFNg19+zovKJ6UHFtmR
NJCwioX4aWdJMkIXRSbv7qg/oA8H1K6DwBoj5nci808/nFgLmVX2MsRfd0FjO+gF71RPODiNZwVa
Zd/E04GFV8bNo6/RpDYAiSeyR+UdppEYG/DFZ/2iBh34JDuTTDXCKTKLlFn8rpXXMuyEV1rb6quA
gMNuSWLJBddTfOvBWEpT5UvGOtprHb3wuECwmKhDfhx2Y5RpHiLU6+s/JwgKOg6eRXwuLp54N464
t6Z7Fag1Wg9hegybDqbJ4UvowXZ2BKF9GfvLkvH++ivKfF9m3/WDE3bOiSaBs82c0A0abLohKSo0
dxflz1oDMtR4aNoCPAJQkjYqUrv/3tNz31c92ULr0pgWYSJz1XUOPkrwQG1cOkrLHl4phfWMBT5k
JcMK+LyTN9pQnlLbRNwaLdFrZxx35rMrMW4oZZ+SXOmKv9tiXoi4cjJy8aHTBxviT7S2SUElVNac
BOMlT359LaXTdruPQcQD6Vnm4LYLm4KEZEkOL/lOs3/g6pHoX0KgZAkfI4dpuo120JTR5TPBfA+P
K3/1jspl4x+ypfbXAhCM7V+jOnWGOThIXJE370h33jV+qm7UeM7plDzu8nqEHsD8LJaYldOK5lrs
UsCaunglogc+VrsW84nAn54TREUpZLk2sVDiawLPu5JCKWpexPnCFI2NaY9G6bY3WFe4/qKfa0A8
++7BoVwVxvz/HmXqxi8yGihouPyIqMPHRmDYiJ/zdaUhVTb60kFeXzenWjx+MExohyfyjk20U8/m
QkRorUf/XMJiZSLAqnvzH7dwDIkPMap/e7pfzqZWq7si6jeRz+HPnT1Gkw+ODXw0ChE/EGEpjXYI
PCBTBS6O/afyPxAbp0miWsa5Us8FwUM7FK78/hIrHTaIDlxKglcanmfc5VRirKQBxENkxCHdok7y
b5G6XNtNgrO9U8EcBOEZD99dGyBVpHBCnhTvSXBGwXsrbXmfACeADKwdFX/L3+dConPELLPlGkaN
AZNrZVSVzOQzopQFsHalJGgxDrvUp04rwprVfEaJMZBDDK1lfmafa97D1GAgBkLZj3mPWWQ5M1JZ
bcNLImWbZfFaZLttB0HwFHsWk4Brbps4paHeRmQOLLmRvO887WGw6gaZn4GTwszctD2446lqYNlz
At8XLuxmTMf6XAgtvEgpWPPHeX7hSQeC3Ec0J1ARZXlTiCbk/x1D4KmCJARLKfEktIAweAju+JpL
kaSUep8BZd1YQRqOmzC1ilUROHoV9Hjymu5Oru4Qqwz5xIJSHEsuR3S8hDi3a0z4xjuXuhylil5+
E9c+BwUoeMGcm77WBi/WRVb6L+cHmvMpUh5082MpK4eRrnD70QPU7goFVoq/6hwWKO6noiZL/SNJ
axoqvXPGpVE/W6RTXmcSspaEN1OmCN5ubV2ZJXyp4h0FdjKCYZYzkFX4OqiFK8iNwSh/t82uyML7
gT9+QhWq5joh4YeuAr7I3rJVlz3qzgC2FInzUtgeAbiqPO6nlY2zQkAhA3FXGzvElhsPFmZP6ek+
tixFelUWW3htr9s5FDvT+9veKqiuYf6DnLyBrdqFFxrt9Jk1sgYjfj6lXTnuEsPy01zQAri9nFnL
/haszrQB4oxIyT1WDJfoUopk9v6bL8cj0aQpMM9fEiop4FDC2hVHC87k4AIx/wk6pGtdhXSEcXU0
18KOgmUon9P/VI0iuxPIYY4s+DlogeCnmoKc1GzdjneQPhvwc8DZ62n3W5lS+t6iCGgVu0anXkLh
Iw7LxMfsdNybpF9ow6tUPYqt6yQMaJ4XB9HaquLQJDQlRFJkD54IoPTuWbFQ40YBKxGKhWOXAwcG
fEaenIGhDFNdALnEmZsoniL5mNfqUsYrmQMrAE3EQXUeOgbpGOgqvaT3n/bVNO4/RevLV6zUX+eF
4fYuel+t5HTK8LrE/nGmUsBrimnS5W1+7HNWk9PMFDSAvkYv94xK3L/LCSzzXVumVHVqCtX+ZUra
rVQjJcpx2SIOEKHVivRV77ClKMcphxIWcoUZgZpC9xi60SXPbmAvXKlGou9MckFE/ANZEq5KfJBn
tZ8LoHHvJ1xF6cwc1i/TWa+GeCEStLX4tOia6oBhZpXcITs83W0CzIxemVzcFd4tydRscNLJJE0f
cKebxIjc7XSpLuXgbhdt+ikV4V4fwuY54ZT2dmq1uYMw2Q1BvAgCIF9GFNi9+HXYn9ztdtxtHJ1o
DrV/7Hf7hDPCunT1PMEDITXZ+Fm45YvXr86ZOdtk7zZwCG+j7DeVAHXXOB7JAu8r39FglO6W7cpV
1wf7+KcPv2ln/uLqnlpvFShiXnnI8EkAZ/dvtM1UfVVNZIRPWudC/rLcf9E37OpQ51o+vZ8Lr10D
sgGOwyz/3n2yR0BhI3cfJKo3Plta6d0rVWB+NAGjBPhC8m84zB49nFerbelv4AZcJOn6qesgMYYO
W61XbfWZZkmMOTQZnZiCQnqFb/oEQYvlGTd2Q3RZRxzMZyGxvCoLPrp586Va0Y6R/txSVn7wkxhm
BJjpXeHchiC4It/febPSr/Lh0vS7XxyFhkJAgknp1ehSmkwfcScXAq2Zp6Smy8cyeJnyi9k02LJE
3DUlYtSeLYuPkXI7cSDmc7UIVNk3TRD8dOOqDwoiOGcUsVvmP2YArJx9J9bPYtxEFFF7HkXYS+J6
o47LAM6TW+46LtRtY+9c1+19aN806bRx5VRMc0jCYYM07y7TNnuHhUubA0v/2IqhKz5m4hnDZs+S
gzIGco6/OEFGaNOmF1mW8o5+ppbEcnQChmm3R6O7eKvtnN8mWbtDJhdWZtJPnwQkbMcvS5mXVuZz
czgdrYIss0teXSEO6TJ7b3CFkEVDpAxG/+1AJ78faADsxou2pn2cZZ0EMjuMBLQIdlqqFjcKRLIM
xrStr9VDFUajXfrWRnNF0SFf6cWrSfNR/nPVJhALdoFJp+eTifC75y/KuwDqhjaxlgl2buhGa7yM
i8I40e4ZY0P28pzZs9TbrL0smNvRnasBkfSIrIdKnecJ7D8h9p7e9ZjQ9owVfgA9mHXjnZRL+CVy
U7EU/JUM33tPQvVtNH99RpZggDdBZSVbQad2HCDtxXjdDmNj4ZP5dHYu51BXslo21xlbvaVb6uBa
8vOIRS9tSrTe4iiWRksnTsNDBSrpb+vM9Rhw4169hq+hUKHB01BidikMdYY0A7aCU1c085+p5ViD
6/r3PoGhD0DiHe8IWIB7KDMbXaNRpo0axEt02IMsM8OoiKp/MxlwEMV5EAUlOKqtcVm5XOW1Mz7O
n+lYN6/9hZzf7h3ssdyvUTOS463BHJ1UnauSLqIQc/joiAZU38PfvFDbRiFPMWwTS/jwK7mkwLzd
ZAw13u7hNAJnz14NG++hGnWxdvXH0OgC+Vl+dnycz1vfUopur+ArhaHPRd60I0rkEnkBqQBbm9v1
5SCBfo7UG66QJB0yzTkIPF+u6no4t2pyxDVRSWci6TyXEnKrPqLMIBnHFYPB7uZJCPDPfqUdIArB
Qf/Vkn4PP/eCyDm3UoxRFvDwvOim+hCfLda88It3/YdcrkEgnaC7pvjTMMa1njA6QGP3YmS7X2JV
qhpEqxqNAB0TUHkvwtGCEtHwxqGeRk7HyZkIVK479Ie+wKEm6oak3Zs9v1/3CywE/gV2P5XNZoa6
/hIcZ4Kl0R3sADiRV91VJgJgPMKgCSnuu4/qeq6RbTWhYbHSFBKNULZBufgkIca2J2bOq9AV/79s
BmK+n8YwSzooQFZCRCMMjBohGGU/4Gg6qvrxPEyLXmMLvZBdKF7sc8szfIeEHt4Um8ShOx/7ZZ87
8ZEga3eN61Shwk2W87NkBSMuXeDICkifAXtnLLjm0hn1dpXqFAF8XLM66/1FMlKD5me3hPWXkRy3
WfYkPnuJ4BJlaXnk0v7Y2oRObuUwt01RgCrG6JeGetug+mMuQnib9I6u5bk/vOstFIrjVbmmYb8O
Suj0Im6jW17zmIkjr8pdJqDtR7MiXFlZv9nW3IUTZP0kijw+95bZ+FOAs152EpzLJ8RXtoGEEYT8
fCmYhaQQJBjyoasYQDvCimMDVOoFjJr6kGtcTdbzIbJQntCkou+2QJ4jACqYxfe9Q/WLj976MTc0
eZ3K1r9Pm2e44xy3GuZZISQNhZHa90z5U0Wts1Ns66PS0v6WzjYcttUCs4EqcW4FvOrx3BczMDAX
kpehdRGnEwr38J6r0k2OEEsf6RUdbPWdYLVlMsa+hEuZOF0VOvoL4WaOaIylPjDmr8L8oEh0RFNe
qHqvZ3t+HNxbWfv9EIX15bB8zpCEHL1llQpJNKq5WFFW3NibNZtfrJ9o0b555SFID0NoSIpnU5Do
nuRotFZclhYRGoy/wABVGogNwzX99xwEgjASxUr79GG2WuVB50Ne5xunhpCm72+5CvBUe0l5WQIh
24Ud3Yhli6WVBcQbe5ZXjTWYL41axe+zKI5xaKDI0V6142aG1T/Y9zZVgGHZD5N1eQo6hmj5XS6y
Ik1AOSmY8BQcS5+kT1ZRmcxqOEeNG7Hr6w5QbkQZFKoSr8VCHgFS40hJ1bqcGQqbJDt5NsiXFLSs
8PBHGD1CYUy1fsM4Bdywq8asqkU9HbH+6y+bbqcZsJMD7URb7aNtk++c0FJJfj6L2znwHv/FXZKJ
kzLQNJwPrnu6g0RvpCYBll+ipu3Roy2NMHevc1ajk9UizM1YXrjk0sRAexiYnBTvwlpAkZ6FCVII
SgRaVroy4zcL4donsNSSdf6yJUplImm5vawIwXu0lGPscwDyUsK+exVj9YcWowyMB6zWiulG1Yrq
XsN0oJFqPIKrRQz6V2Dg6eksjM9mNZR4/JQ+6pAe8xjrVRQEW1YNFOIif0F5jQoLx/6eMqG4lzOn
KfyB6bgmoNcOmboaGZkaaujk7XpD/kJz92pg6n320PJ/VNezD3SIhYL6Ym0awmWaJqxrBPJLAovD
Q1gXshrRhSR9zNFtgfjmRXcbBacuMx8kGqgG2v9b0hhzKLjocFL2NNulH5N8n+UxVAzRbdB3ASoc
In+m9StAO6pNy6i3DhEd2LvRWG2ESEGQGJLAJCAnscSFdByV/JYIrntnImmeNCPM/uijFtRIPInR
CK+ZceIxCy7pvPayTPIMer6MmgcVrs8vypOpR2ncZWm++X0Dv2Iddhll2KE1HX6ECFMDuMdpsOD0
l+JLBbRKjpL7r4MKTkN8kp598bZ9SAPVlMjx44lkKaYaCJfoGAeoinWDaEE+TPSh9v5m2XFyXSXi
ySfO4mhlydz3CLknxbncNC868LY43z1KkuEZ8rYsBS90YKgE+E/Ymtm67Bjo085WSCWQVjLl/db2
NYcI7jtXXuxiH1SGDXx0gkKoGEkS4K4JPJJsTZFnsis1nOWmUrDJg6GmBnnNEom/0miW/12Jp5hO
dCMwp3MyoiR7XpOneh9Ro8LmcYlWNTlfKSFJXJg5u2sHKbxO+oD6qgUCJUAz5AXtv6lzMNGK66tr
sALEry0bSQq49cpuUcsTxp9wYzo41HmRbPJhGALYbPYWSJRKxjrXekCdcBc/w39KS1gI/P58/VAh
zCNue4v+0YK4k052psIHWVkDmfM7az+6BG3x8gXfQNP5taQ2f7iojgssOv8z4ZlmJDU3XFaVSAlu
XVkileO+L7SpcgpFPBhPEwWohDcYAr+crG1ITGH7Mxu5vKdqhGoi+PIS8kyicRJxl/Nde8byqfU5
cHDe0Rkf0lpFVdQfOzWCMrUETfS/uKGTOEh4Ja16UCLzm1GOiXD2ggKwDZEdffSm7mvhIlVahJbu
BAmzshO2qVNO5/nBqOf/Oz9tXzDkSdST5ODtHqTfarvT9ji0DzZ4YrZEE/5Uet5H+J/C4rP+jHYb
+PhAjKbWHGJQ88YmKoP4rfg3aWZhq7mZCWq0wMOxxH+XW0el+jwtomK/QMSneo9VSTYTI98J7zjK
ijtDJfaCct0YyWqqOB1A240q5pLXO0/ZkqD1I0gfZ909PorPOorBT3r61eNzLAlz2ozyYxXptRoO
ZKcEOWKuVSItWtULua65TIGBNwPaSLE+ScYTQDxFwg7sSdhXFh0DLBqxD9nrpnoZyZ9zYKnGlf+6
+w3VDoS89EJi2MVgWB0e4FzDXmDtRshlxOfaUmM8jB/ecjRF5ONjlgDbVO7CtzwrAtfB2GrQiY3F
2zKySCbMVR5WkKpMwzxD59MRUfjQmTde3tN6xGU+dHHMOXtV3lRFypGEuc1IR05mkjORXb6SH4b7
/RDzDh3JWvGM1nDMO5HcpcQ7A9bqvjt4GO+YNOkj6hwyTCqFPlWO6mdlgmPTXTvrDHARZBUlDWk8
tb6Wof/JF4i9rLD7ybJqdX/ISL7+gE01lqub+6etNKxT+/turW3kJfeteymU0u/16iKenZDEVsXw
S6PZgF8w4SrJiL4f+n+BXSNWru3AxxGmfrjUORYygTjtSQkDhx6ivA1ENsWEcFHCYgZsYAGkf0fw
i4B8qfqkyEjEr8XfCxka9ZDBb31K8/+kRomZHfxWpzg9tmb+ponOioIBaZ5alb4B1UACTIhtsPl3
iHdBuopGqp8CM+V9NYdteJPmQ6zGJ2qhcvXG5DAs9GBzd+e3uR9BjEVHz3Lww+W4fDT4soqSx2ec
GT7WB9YsNumZ8TRvkkAtPUneOwNIfwHcJdMHXS8S4bdQ1/CGUhmW6BUNteQopZfnzBUbLOJICawJ
tcnGibcwfnCSpk3tS9c4UxPbWB7jnOaPU6VOOOELW8AlgagKSPYGxWzsCx2ND62Uqgja+Qsa1fMx
gROxwpACLNZ5BDxO4Efpdd0L/SpXbUpsx2XCt+qMzdipR9qMRa2MO+w5mf4DAe8vo3Vbs89xPFfy
8PeJQYV9++kpkh4mYWQOuXH8OBLYiqiaUgidfLnAyDlvGKCPk0Y7722g0XgckBkrEUcb+IIpHw9a
8ap51/fjBHDGszyg+5RXwZg/y2cee0evTQTJuPQxBLJ4EiGtppTSC0ph16oBEuQhFb6jyVIKJGym
6J9pB43fls3OSzqhbsYW7/fL7ywCOyfKe5EbdQqtvUNiFy/AyUEy3cldO7IM5RjE7Jgi8N2sIpIP
BZymYHx8WGLprPgJizhog231WpoqnAFyFyKfby9SuF8Tf2et9hP1HX2gk9UmGCVtwsJDnwNdYn4C
z09FBXXE2GMAwI6rGAvMqikh5C0UPp1utSCKBDCbVyvmCvQlILkSTdK5LSjzIIBkzQldDrvKxvuw
KXTtpbYEQfkVNOSQD9M99zZWuR1nNMnvS/z2H4TfD8Rmc6kIxOG1AeBBzSApjnncg9pkr14GFCJf
sOkDwJLzRafO8ymAN2zHSdLaMV3Hd8bXG75tyyfieIk7VLriLMt6ovKBO1hQeApDP0U5KT/uiRvT
9VWgm7I3KRLGGuSMXHpwAcq2TDjHoPUbMdGk9uV5mki902VeWXLNEQ93Azey2AnTArj+iD3h0DlE
WBiYZrJC+YB3izzd+YbglDyCRzuTkn1JfmrxnnTuqpDa1a2/nMJCd7QpLZa4/DZt/QsrFdhDrNi0
Yus2xwNjpHYgYq9qVb4snJT3slrGfrPOKuNEPt7co6Ndcu4fmU2cjRaSFCmpy+4/7EkWquSV/tn8
cPah/CY0QvqyxFxrPAoAw+K1yL489AjrYy6Z2Fn7W5sPpR4oFTlH8Ct9JexItohSXGO0VteTInfa
atQdjntQ28lu8LYnTnt8heA1T/HaQuNPS0Aoutzez4TXeypNdgU4fZ5MNCQWP/C/jaQBN7QnFCUv
cKaVmUxxCzRRJS42HcEl+TOQpulEEUAYkACtN1TnVt3tS654l4FO2FLZAmfyAXILxWZMEQJ0gFIm
ZSnfyrAnxxcncbNN+UL6Qw/kCOhCo3YsjNeXZ2Xa7qfQFLvAXuI1veYT2MdZkkvnvjFKYgCjHf8g
zNrPTRDHDdm7JFjlqu9aBF3VVeA14h4zMU6yKKEgmYpR9h+vfNJ8qlI4UtgiJOmXXFVaSwoXGevU
MqSa2LlZO4np8sx2QNy3F7YD1M+oRycVZTpD4Olkvez895p2YHF7yAv08SS9dN06u+IVgG4YNBfg
Znz3BWLavnphNkwnVolmY0qKtu5d+0xYquZ216nn5hfj13R6oYy6uan4QK4FRjviHT/D0jdemPQ/
gQA/LiJnEQR5CCvSB3EbPYBEJPJogSE/zK+qTbJRuDS7vx87heufR4RAgNPPFeyoIKeFbEqgq+j/
Eyup8bMeXXICdlevmTeGx2jppxCcb0YDeWQZg8+MbJTsSu/QpiYdBTOkn0sBEh0RooSf6sfcncIW
VqZywP60o+ETHK0h6xJ86TDnNscLqkFnZF0N6K1Fb+b83icFjSCOpYa3E1BZvWCQpVkblfzgoddW
/LuhouOMbRI8V8YXqrJGnwJ9Y7AJeOc7/+N3I4ehE4BOA/U6p6RUA6yldXhhY4zpNO8tNnsYMK2c
Qk/2tGOV2x1eZg3KcnVJwLILVguRquh2mxijj3Gf5cDmEcEPCwjAGYzAbGQ27ishMJzsV6Y9B9Tf
ffdFPaxBRSz7lJcioKoMCi9hlLFzoJJUzzWetEUTPtXQJBJjtqAXTjMHESQy+fdJi5sbcwNgQQY0
V+KwbWeRf2ex7ICHUtcvpF59dORurEqh8wSKa/67B+T6n6aOuIEn15TaiKzBk0HAXc83OlotIJLl
cKASOv7RkJJ37YL9FDKUusG3cJee0fenXQfDHRwjd9KwU6+d5O95zfZRmCf22UEHjZ0iJr7Ce4sv
v4XxAlcOmbetLkyopvxgkR6VOY/6YgBHCcjFNB9E4KuB2ue67nOyyRR6X3e/0Xcw2YJ8LkSrekmK
qGhcjszyOrm0W8m9zboXAAlwGeycshdbrCWku54Q/6I3TlP03MGUdL2e7svsvvlsIkB7xb6wXrek
wGjlmzKl+DbTy4BNse3sWPWqlsIvANfC8nlbTsRL2z9mxDml+FhClRXA8y++XJw2CjIyYRoJ5Iuy
kRI8oek+xR4llwhwYCBNmK7kSeTR0Wy016pvl6b19V8BYB8rGitHvQfT9BEUrL5sZZcIJzs6wJVr
WtQqLv+IFBmmBU9SxJTAfhOGs3r9FLBSKVNNQf+zV8CiLoFDJD4UneOYt2AynD1iX7Jg6hxpU4W1
HvAS2n1avtW08tWkTnngMJFDRIyNFGE2qz1Kv3mo98SzY91OTvcEZbdBcz3+JReRMiE+t8bfuN1O
k6BDLshoDV/IEdv89MfCQaF3dPKxpMTphOawsBGouTKuDqzdIeBVfPtuklraN1r9zYO54/aG7N+F
jEKqZkiU9FcW/FCilgGFLvmG0xTbuZn8vn8E7SWvDAFr1rIeFlGMfSS4oigR4tCX5Dm+RpnUJeUL
fmyP+Qe/wnSpBah6iGta41S3TqbN7fnAZzpMrgN/tcaEU/RagfJNyIxgG5XPiqkilD3reE8f8l/Q
hCP5cDl10coaIxEEnEcBkR4Rwgqm7pwAudz+Mj+dK94CIvVnzLJnCr83VhcHiL+skvYV+WZ1bTDf
k0KOdunCYzNW2ouwq4oDorPW1RtgeiQXiV8wGF8nWsokcBeDmAJLfml4Z/Q2YjmP2na4B2MeuDbI
upkJg+yPVrY6S9Qhna50ZoDsF0+Uj3WuUCmgNuduN5DNXfuLQOsLxlOdBS6/ZEZINosmWChsFHeL
Tyw3xUY2R8q29Z7wfJkkeeKNKCSVIo9XIIQufaP08DWrFbcc5ouela3smTLTWiFAwuQQKFDCVQAe
2bLPgb6f5uewRrr8A1zXLOMNg8UxzNtChlCsleTwWs7a57MggJNIa/S7dWgR41CmRMRw6sW62srn
DXJdsTarmXu7JuMFjHDDKVAnnxSiCz/wKX1ZwnMvht5dGM2Kcu3UQ8p6oeWCoxTv4FDVe98qUnVn
asomYqPjLmErScDx5xT7FzLRYi6RdDjLV0pd7uWVmVDwh/6WKa/EsMJn+D/Nhd3P0FIVvzWM08TY
rGGpVZtqtm5yWbYIAgzqaWziVjY+wIli/55ZHuFJcztuowCmBd3DR+664JPUbK7jU5dP/vObVQwD
b+dPdsE1gn/XEV5zWoHf149/6l9t2/UMf45OevDzllR6HvaEIMoZr7Lm9hVFEH9tAppmjl61u4+R
E0NPZelgo0qQK4H4fQZ75ucBx1DFZNmd6C3kht12GIg4MGin+4JdbHx2YUX3oeFLQe1vfOtPVvXr
7DrD3JUfHjzGbx49kt3SFgzBWbFamTUozLtSLhmqh2U0haQSMpkm//BrZKvbjKToUr2ZpNuZ3Hvw
/VHON5pwUc3j36FW4Cpuk+mT91j6U2FCzBLTbkhWJXkZcVzYOdXC4rXekAq4ly+BX9o0Nmqd9hQi
V//3Mjmk+NgbQOWu1IIM5c5gnAcD669mQL38DKETrdUj/F6cghGat2gv7GwC7MoU5EUn/H0fhFNZ
EDak9K15yvI4594IKB9Z619C6GKFgSoT1lPimvjkg9oYZsm+XqA9CaVOj8pHHX5H5osr0t1tAUoG
gK29GvzComyc6Ka6oTml95QFu8rig5YU2S8BmoWmdHLq42H29gjTGY4F1wSZrRQ61X2+LJLRBUHq
Ct3IRbyzabI250/8PJBrppIOm4ohUTIJupSQatONboClAua2x4bkumrZ8OrCyctujEPC246hR6pL
Zl2KTn6yCTSxnCytIF+XWLlZwwyHojLxo2VnJyUlc9kodq9AmtnZxqgQIX3jptotUCNJfrwXZzDE
XGj+54qpdsksIygcfeocH2LTWS9qVQYEalA4bGecsxkyDEhQxQAAFB70oETeedCK1f0OOWIAkrw/
p1walB4sSbydwUODcu0IgenCjwPO8JILoxzOnHsnEkqk5Nd2/YO3apZl1ywHL1jUqmUDlgm0YGuw
9cWxePylsFbxcpwER84Yvqw7YhuXmIuWKDD/fcTuk3c3pdLCa3v/9MwZ5wef30zYx/Xs07yxhlVU
jOOWITygw5UsnRS2XzFWOJs5ysIKlRlik/9JqY9MpNIprG/Bfj4zTlvwLc9/A7mdCG5z173siSYu
GxWcrXYAXV+pWKGuxOTcy5BhnaNrEOKoC3o+Zzn+Z9DVqMj/mZf58UMPuhO3qdSIVFTvecyA7wpx
Kw7K3TuMyDeXgXLFoVALo9Q2exLa5A0cVBhxe6e2Lw8HwGAYUZ/uBqCWB884o23Dtf7ZIohPWLCf
IBxAESHhDLJw0x40EvxFO8in+zOKsdOP92Sqf8LlXz8Kao7UxoNRh+HSSTkoKeVj4SuSbP1GG5mm
DTN8T8CvAYEnx7jPe3SUsLNMdNljsktFJAGbAqNxTxY7s/ZGAD1A/KLlR9pA/eUCvQYWPURHNJ40
cjvLWGjG43nB6TW+FLeR6QJ1fB9JpUJQ+RyjbTsPPVEAPt93u7Wa+Ky+IJxVS7bbULK/JHzsT+7m
HN/fzlVGpvNFfViDwzg407iiQCiwbvXL48Sir0DFThpCQwDT1pZjiPnunr5x0RWs+x443jVQrZ8Z
Cvk+LLzpgQz2u47OoHcX9dhqTXzbecHhNocoaV6Cl24hpgRqkpBmMCEjDlBQzranDHzeYLwllRKJ
xA9UHjs20ESyyosvVp6ZedW0+n731q/4b659kuVrneVNQmd/rYE7AD8OvHCkj9Up6o8pWJ1hXxUC
qVkFhY4Al5+wXvTWCqrDuQnb/XFXNl7QoVPAQjGW3fAxoJcy3FhDGiqIJeOksYDw/mVF6SqYto1o
Y+NsT6JbjqrIXY+dX/UunJYvrV+MB9nEORUzN6qSwLiqQMX2WCFLpxZn+odI4xquZkLqV4bsVqgY
bqJSP4/XIEDmMrnELeED9+VmvbwzHaWAVL8WuoH5wOj9QFEW2pBuJgA+lBGBsceI3s4DmpHh40jq
mcPrnWZb81atoo7OKedJ0ZdD6L51AVelkqFd8C6OqZpovcJ1i4fhn4RDh1rpEgzxhEJFFRCj61Ug
zYUsctjcnFVk4Tq4D6cCbRJiU1GaukXTmk9Mn7V9zhsAc+6ZIA6KwV802CKMR+Ei+SqOPzp/4DV7
P0TmYSpo5Lw9E9bmwC/m5TVH+ndcJ6xTR1FIlh8OF8P1gLeTtqNlB0I951uHMXb1qWcUgcFWawXG
3VLOl9WPd2i08UV+66gJUb1Rz6Es20A8EWalMkOF+oP+k8xFVSZLdFuUnkHcAeJ7K7E4qG3dBF3l
pSRQ6KpH7l5ELKogY1uG6iJicd6VexPYBBDLj+k+xOsBcuLCkU5uBrnCcLKouMASy9kp4jtAtVeY
dZbbBizWN3MrgGYoua+OXt/vJAXkz/OIR/+yq7wJWW7ttOOe/vBCiot5tWU3p6BND2QbXZ+NNid9
OtUw95YZiTi3bmBIyfi/Qzu+ZemJej5WxgT5LbE4DFDqm8wPH1Wth//km+D73qHBqF6zZFG1JGut
tnzwBtcNdyJXs5EU+qadQLNSpUmuKrwHvy5WyBz5OUSKBNOseNG9QnDpX+fBBuyRqhttarFwFdVT
s6Q8/VFtHG94Z4iKrRPZuBj2yrYb0uoaH1RIKUw/sBP1Vxar4Lf9Ca/luOlEwrV3qIrxo19D8xI0
rz64cCXjb9pk3rtDXr52Fq+buLkPX8M+68mta3Lg/Cc9CyNQiKO9VZ0HYbifgxJnStmSczW8UOyt
xAsrynujr7nHhMKiDs74NNSmmz4zKiHiwkQh/V3n2sYSt+FYvAL/jN+rqcm2YtPbuii/sPe6zJPB
kjgrwRBG7Lftscr/5hLhXIAMM9Hv03oXp1b2ync++k6x1KdKHtE5ReAjNAbyjWOA41PvENQmh6Dx
8yavGIii0GRK4HpRSe/EOuS8OcZQEiordaryjfP5aVoBiV6rpy+VSbf8IgMDkqwW1saWXtWGYkRf
SqCNjMdtZ01L1mDSGQkJwQAEvZ/8JjzYiD3/czrcpB56+uA0PjpRoj474v/CK1LKrlt+gH1bPA6B
V/7TW4lrIsX8kAevrTKzTL5tiuU6uwTZ5WDSTSa7TLzOHOcVyLQWWp3+lHV6Ya4CsETRUPXP1iTW
t+q5WTXwQi1Dkmj4k9WM5+TgLcqFGqSRFyeT3jpveexR3gSREAri+OagNdLWf4JFOmqi6U/GfJyr
l/SavnLVzPVmPWPUY7oFJPHmhprXY49I699z3Sj8pRPEiNuAZvDxHmWKzdSaeSax6RzKq7/lCykl
QJuWOitIXhzbsoK8tLcPLSRWpxHQfizsmi64WEuwFqSRnqoC0VDnBfhE2O9inZkcjbJDSCYl7Z/b
ju3IBr12A7SlNZ47+/pmCnkidB5ufYT9+IOJ0AI43VUVUA5IwQX5bi5vDlKOiHEP74MyAKyzSXXm
HVtVh+30cyB3+Piy94MDe6k6UcZ3/XzgWrd9phNDu3aQ7ilAyOMd+LOBTJKFoe/N4QdX+aRz3ssV
dxxnottdEn7tFjudcKuBikUSqy5pRFUUsUKRsnJYrEXnQZks3l6itrK6NyMOoAUwic/0tT+VuU6s
n64bWlW6D078J1isPHmzbZMD6azyhS5KZWnXUsOBQf2gFM6Ew1a2DJvx/Td8FAy3ZYtZHnjtR4PU
EUbchrR1CC7w3KkeCjKextimJgCbYF9jxwA1yD0vUKFzsWk1PcsQdy7aELHCFoYmetUlXmY7Ae1g
fVKBYGbydXCjBJKspDb5l5WY07inN9g+uNMsGovmLuAArT5KyYReDDaII8ENUUZF3xZIBWylxJIG
Z/4pnpC+Co4kOnpzHBvK+TN+iX8kBwC8Wy2bCXYYvx8JGYBYVYRbQSQMoTe1XmdoHUpWZUcKkpWP
2DkSNbIZwmcF+nM3MW9pvXix0dAYWEA9j0da/ZxfsgiY5tSFu02qUCEyC9xuT28Pr5Nk7tTWw0uS
4twD1quyV6A+e8lwzG3yex3voukQp784Cbo89Y9JGwzOaZ6LeZdPcmLmkwPQvq72RnkJMi6g8naF
KP0XzsWE3RQf1koXAuyBvfDOeU2R5qzb36t7mrq8C55mFbLvu7/z5M1ysPS5Js48HXltzmhKwqqy
yi8F74WN1wfpr7/re+ll/Fp7W09oVaUfxo0VXkySWuO6cXjw9UuRfHZ/dzIhuch/ha7jVZ3so1ST
6Syd6x3QhLjw05QpQch/WPV0VHI7LoXHS76g3NLXwqjd2CiLcGm0TCyqf6qxds4yjb3wkBCRmpH1
4llLldGvRox+0gYbG7Z+1qe25fmrBVkxMQGtPj0TmDyOjGXp2o3lIYvOw3QVJ6nB2voMMCfC0FwE
xTdYWgsjf6feg8y6Z9lighJf3NWZcVWL4n82h8SgPmu4T3E4S5VkFMsDpZpbgo01UlTKr/2LUql3
eJohctptF27e0GKkFO7FI3aR51lRydzs5fdzFbDsCtW+rcTThjidJyigi9HOS7zgS39TqK0X7t8f
hgiQfAAW+cqr4StaJ4zK0Ec5Z7LVG3yxvSem5vTOwrSGROtSaIoZKfST6T9PRmvv1jJIoVa/0WcX
JmkWoDOwS7s0ru4/W+vKtvf6pXHjlQ8XXBdlrC8xvGGczqJCAUvxTybWKHQld8/dYterS0oHNyWW
gll/HCbiVdKQ1ysAtcYfbCydU3JxgISgVvrhliik2Ym1cs07bTQ2UkX/7J8iC2BmmfmJWrleDRcN
sQZkgKl7TTqjckgxctgVNc+o2oSpLtF1dFFPzv4OWiYkEhxD5zBbGedMsoj2/p16vcs1Bu3OJNl+
obN0afpW0v1v4hTbwJDpgTraNhMFE1U6uMtRzWt3MvnYC5aT8d4GpvcbHnfwQLJy5snM2sarMlmj
+fckbJ1flLbitCnu2sIEjdlWmhR4BGLdZRUOmVnM+7zPJlrj4AOM8YFzJ+OARbBjlJU6+YexR5dY
SUrD70ubqu0haKFWq7cUOqrBcMOC7YVmVg2RSqWT83m2aYfE7lr5WRm2EBBVtLNdRxftSLQmloUv
p8k7tqQ+Ve7cmT6r12AgXO4GM0su/rlteT6zuDCiFmM1RzoIDFgG2niPV+GDqG0NogSlrLfqRyXF
MJmMQrvyuCPbQO9n9CT3Ji9Tr1OuOrojTsrx25z+IsNFyZJfe74e2KrXDme8UMjGuK/H35YHpxIk
1QT3eRsTcPXBiBmZwlFSwEdOmEeZZxI08kRiPDO4RLpi8oT1pCMUjjCGjsBFT04eUjWL+QFA+Sro
+p8qFLZNxk6hlyOFu5yHfo6u/UIQHl6Cr4bGp3ybHeGRmeGA3wJt7zv7UgOo+yV+cp3jceoF8A50
zNmyLYVgP3MIa9c/1xD5aTzj0pYPj4FFzbovgJ5dro8HoB/CG1rTiw85fMs1orci44f1xcu9kpeI
8tTYokjwtLb9aNFw3gERYNXxLpRDwAR4BP4D/TLsxGFvr2yo6Yt39chNBm7PkH87vrSrTWCRNPrt
S0x93hvj1GrNyEG2w53UlFR6p1Xob0GYkVjuWA0AUbQIfcKU4ITnhjyQPLkc0Rqlnx6R9br6zW1y
4AF+6Z4RmInaZhCuIoLdDTkgtmBBQ5gLWJaNqUXPfvYsjIUxvfAHTHtoxpBepi57Oiadc85czmLl
s4eQ90Ft4CYZkob/cYc3X7/Dwj/qHJC8LpZwQGOBN5UvUgQfejRLyRA7O9ItUsaIaRMRJwbbB9CE
1+kq+1AOnR1kh/poXujQHt997UjnMzFNMbIYNZ8ziFlBe83QIr3OZWH7KrDSL/IlW5et28bZth8h
N01cOLn69zYttfVswJHbVkYmhPU6yYhExEd2eoEflDo0yMwtrqI48fg+pBgvknfAn5UQecdKOhjV
gL5UVJnC0gww5ZgS9pF5wYF4sUflZOykSKzT4lNnCs9eZyNlgEgaNVeYyVHjXmKwMMHsWVFpTRDW
p7frgYlfK7kCyWRsN7yOmEYTVxPFq7eYrezVS5dMaErSSunOhMcac2iug5Nq+rrJRgrBJ0I8lcGh
PYNArYNe5GF71EEgRoC2ZFrogch6hGhiErFALnwHuOQYSPCqmM7UUwlCgcjOKTM8U/DG+xSAXOyg
AfWkhvDyEZxb/pyGKCRFBp3cNqXmQLA00dT4nq5RSf4V5+qPT5JLmyZJYdur2dfoE0Lbqi3hQR2s
Zpd2EVDQHDXJ9Zwzl0SEjKT77tgm/A2SvKqdxad8c0NavgqBpzHtLX60EpDV11Odozj2yDDrP2SZ
GVrACU7iiXkkzylETvQOhH52x1MMvS016fE+if3eMVDSoXzUdo7y8jQt68xM/4phVrquTN2xx8px
wrzXRs8ruqOhanAGmSviFqaCbA3wHt3Td6skAScYSEnFOGwr+1nPZNt0w4RhgNkgSve8cNu6jH5H
xaXLX+jiPUNpIfoDxn65SywsFpM92+iMD/t6yRZ57umbtSQ8CakR15XRgw8NWVUvWIzZZJ9nWTEH
g94uJPOcaiQqcLG3gZXfbcbz99sVTkhvqNHkPjHed0kxe+XjjYgYKp+/QtrNU707m1IEnI7cVCSv
UyZtpf9xLZbalOsvNTG7cm7RelZJKIdM7llZNL9hxNXHIpReOmeZZx31Bb72cvY13/XVr38JepWG
4Zp/NpnkWb+3WILS1SVLkLHZd7b+ayMAKrqNFvJ6LGfiLGAyu0mCMRx2GQKtf+Yz9fd2Q+MJQ6aW
X1EpmoyFDTVyyIftCSDTBkKImIupDYeNaXV+ed0Ex/lyLiIwhmX9HkJR0udjmc2y9p/A78f1Gk2L
fAkCln0x+96qIIPkhlIOrwiTZoFLRb4MS/g6nMg8mLblCMK54QvqLFtNLXnG1mfvBHMPMdLwrpG3
d1p3LkXji/TGnT2n+Tct8+H26rvttnYf24iwQ+MnvYg1RN6uX5Gfr7k4GvOCDw0ABDXXDr/QCAqv
xwiPKvsMLZUqE2ry2kLdrFKt3vtsBNFPbKDLDeSf8wZurGEQKyE38nzsvksobCIjA1RhFJPuY7vc
Py4F1MunWDoQ0n0mCZ3faH9RevsL34/iRhzwyuNIwRyRuEo9ujQTOHo2/sNq83Vc/kcJesuc3w1V
XB5Zu39Ryqre2K+ScpuEfaHpFYTJmr8Nf5zEvfV4fUgvfTHMsaRvQUHoK98EuBKU8rkI2J/9C48u
LgJ41/XvL9JTUYI4WaJifhJTt2vQTHxe1IYI1Bp/8DJOVxdP5iGQG/RvPbQNNZmCu556c7KcY7GT
UATXOQE977yMMWaO1gxGcVu4FkGsMQVWEk9rWYM5WGPxvkdFDLV+NFp4VJHGSk2ygm4Ib724qpZP
LHfCfwYzCISdYXSE7AciHq6Jb2iQAWBcC40yuuezFiA6pU4BTrNTrH33iBto+DFoI/W+JLjzJe+o
r6RKb6modwVcxsk7KI7TtMPnoFhPchEke5CLoVa5KVVXYQyhUPGzp5Ilb20P/CM82In5N78vJQdN
JP7Qs1Ro1izlHxDVJ8jTaaoqOEybc/f1ttF3ak6axAgkD+uhMkQIVmb190J8YZJ8C2UTNtt0OEWZ
VTyHTt2YhZjfzdMBCCo/SJOVZqTfF/9PBH3dISd3+R2etd6cpXZajqzwBwzJ53aCybEcGDoKqAKh
magCc4K/WyovdeBxVb90MPRl9Xe4aIHTfBb4D7PA3pzySBJs4wFDqPEMYgQ4FqZ3miwgBlsNvu75
CX87OsDdYTXAZOAlQwP1WqvGGZlWTZZiBS6c1/YQT33H/H1eef0vVmt7xf48vpo7uZUcJ2NQFraU
wYKEKsMwkyFSVoaCzfGZxviL8m3RiUZ8F4PvFdJSM6jv29BV+ODIfnIo+fEZ+WSxPAKpF2Yzvfu3
ajxbP6jq+7YWTBjhw2/bJSlOY++OgX2K1G2O4GL/Q2dvTC4aQUmU7EQ8IHU2igih5FbD9VS1ObxI
PSRlStGp+RZhfzjBXpEns2/Bcjvt1sqNvNtAmU+joyx6clsAYOxqBhQaAagehJRYCfakSnDXNEmP
kyTiiG4EiTbo+ftvfYmQX3ALFymZZYvRm05wa1zqhgumFFjltwaZWAHLXtKnxGbBYFtNg34GvGQ4
Il2zK1aKkUs6chTz8DYF69nb0wvSX508wMCiy1cEK+STOjJNgkKynxceptrQ5f6yX4AosRLJMPcV
C7NA99OW3Dt/v4s31syE/PeZySWa01ReHyKjHo5lKT9FOo3YuedpZfqWYs9GE6nh7wevw8KxKt8Z
BzzNw91AGwK8sqbtEu+liQELMAIln7JvnLs+bsXXEPywTYg1i2BuXaZrmgAgLPpw/jAjR+solELb
i0a8FJ462ZPNES/YxiK4payiQngeiMZYhwDyU9u7JyuxkdtTn8x4AIXF/iQz/GufDp4pQ5V8l3p9
83PGglNfK/QxU9Lw1+FNYlNJY3Cjc6jNE0LrFMPEBzKXIdQaO0Qe3CZypcCvTd6655g+romXWzdu
KFXU1lCFegUG+H9kk4IT37imsClMUsnO709xGWkogPqAGuwRlS0I2VYfVQiwMjwtzNRt+Y8Equ/T
tBtWxI5hsziQNzKJxSpN1gapdED/J1rKX9S+VYuCrCve69xlJ3b7aXQwdb/4iC1HSJtbo3lPqs9A
yV75QVKYouG+Ka0LTJey5TpZRSF984Dd94nBlic7ul7gwI669aO7TPhgTAujRHQve10ys+tcO8zF
cYaGp8XT05tGHSBFtnQpMmEmr62MUqwr/ei26Qlg7LDJLffZDMfWVeSAssJfPyeOguLJxy0R17IN
fq9lIzReX3+hS6lf6qCZqgnzgNiUdOWaJg5+MMdRkzccjz7b/PCL0iRqfvWxR9s/zPxIQsASz0lW
M6Jl/V6nTACXc6FcF4oL0MvbT0AvgZSCSaJ5MDJe2oA6MHvXoMrsSqGufwH/20SLvPCC1tE2m9nR
LVnlRpiRNrptSqNshcVd8oaQRYi5i0bFAiUipxmQr3kUr86s3ewfjcJZUIGk6p+a7hssemTi0DLZ
6M2OpgeX+FjFSACteR06snb25dEh6k/vyDNFM9lO+DjP1Nn5QlXFbI1rtYRl/ljTqc3++9bHXyIS
3zNzqmVDR9AeyC2KwKolnA8OlUQLkg4zCsSOITRNRAKCIEGnxXAmTgTUav2uMG3hI8ZEarjmat52
DvJjSJgpamV4ZKoVci3lzKfUTAMZ+XaoMqczY/9IXcVtqbqaHvMIOS/atM+Js/hhvfB7wpyEcOTS
Zc0a+C/ni+oSFzX0T2tnv5UFdJeunzIK1SS0mChbPHIl67UJ4NCWV1pbFu5FdlgU95Y3pxr65Yya
8Ib2swzHVUCT389I1rDiOgreT682QiFrGebUk4ASERp4Db1PSfXzNULkE61kVTw5p5qyNT0T4gAE
Upchs5d8JAncr5NftyfCJy+eVzhYI1Jpud/vT61a0h40LIxIo06BhyJU95ElRShpfRhuBsRUT1t4
+hfJSZggg0TTqQRcw0Fm5YIuP6udIV/yivsNOkgAZ30Lyq9hlMh2PHADW0/afbypSo0edaoMwClu
RMGMgAFsBbdtG/i8llV8SJ8K6RQBCOSS+OK+/rNMU7kjdPG+OT+sItpoMoBDKmx9BuckYIszGibT
YPmDoJzNqG3XQGzp514JO3dYt0r5LFLWwMTY8bYkGuA5lcvQfkKGkF4TQ4nY7MHJhc8ze0kB3mSj
JF2qvGZUCmAzC/ohX4GL9wVYAjA8sG58lR0ox+pGZqgt4IwGqe6/6JIQl6NTl+NEW72jEAWpZD/R
ysm64zG/87b63O6eceyRlmqwbq+P7uY3sL6TPBI9j6q4SKAGC7PJRQ2dbn400/TfNtn2TigX/mwt
FxyuhJfI7t6UPstgEvs4TPMbFWLbhWasG7EYqFRiKTJjTdsWV7utVCHr8KJ7R026f92IV9gIY5jO
elbDnJvJIiYI2NM6VD7tv8HMBErsNUcpLPZl/6Wtt7tGRuur3s4ExmKQpeZWCGJBvM3n1DGkJlXS
ZSqTn76lFchiJ+MtUp7BpNiSxeeCPYQtYxPD5uIKP1UlrE7PsEOl5miDmI7R4/YntN25I2LHgv1T
e+172CCfsFNtyxrpbwp8RvRYc6fP8G9QFsXE8H3t3zLvScKgLIkfrmaiiETXMFVITmiN39GxyYIr
AXUoeBgg5Su9Ii/ty6c35JjzBgfyXbSHb5fTJfCnMgjFVosvs20WVxmRC4G6LHkYEzN8Yk91INQz
ZLaa37r45vlU7P9Ib1FKDWnj7Np1z/DdI8Jhzg4ZQG3xlE9Zahbtzqgk/74TPuCaAO3FvpzaekpM
F0zc5AUg6nfGAIKoEHeqRvnvwBCVcELXuM4HKrzn5WwB2YVzzpQ7cbmQDFYS6dHMUe1NUbNAad0T
Xq8t/tkkDCceFv5cnQAKSCeLX97/9imRTMll//enxMUhDCLtJCnTICiA+3J5nUdztujfChVCud5E
Tij+sYpelcD+AvHr4JmOPq1MftcgNBl1w32kxcgwLENrU77uWZiASQQ4MU/15h95BRFhwte+2jR/
cC6GDmEVDRvAyuEIVWqcFpT+2zxdoGgAuHphhsUr4E5jf7IEJNAq+vk3vCpIIEy5IWVxyoPh5ZlK
Q0QW+HoAJ6VOL5kNtQbQGvo3P4zfVMYgvCIKP41pPFpEhp3NA5VFcuCq54WQ0DIpF5gnFHC5MBfE
Wzae2ZlL4rdYZZGRB3pMZ23aXGi3AbNZxsD3WtmA2ObLtZ59QQKPCzpXwftEg0IRDEb8CCNnO2dQ
T7gIg+VZ2maSKsowhq1GwOa5bttHaBxjluCBxMhQ111BzxRz4668Wl5E3t6U6NTwGYhZ0SnOmWg7
uvmm4OG5BMShcHuC7cxW1adnmmhdAcbtX197rZyx6m54zVmC+O43ugC6fiEp93n0EyJw1PJsgcxt
DBhdESypoSJEeFjnU5mxBi7uJAsPPrMwup2KseXo3FQI8bQUhfYXAMBhRT2e3DvAbbdEmLwXqm/2
CAbFkwfA2eq42pEeL9rkPxJ8tuHJa2sQUYjpfb0Bvq+AL5J1L75YrwqewYhHPJpgCp7Pr6nd86aQ
y3ptusNMFO2gxE6dndwvnO+fYMHmUUvAOv0m/SEDg3S2bOWFVLYVzXR6FxaVdlPU/hwPpc7hG1lJ
1fQEj+gdXNBTQuS7Fk6x8luOpejElxYSbLgFnzVmv88tSgdd7dN6I8dW2j+znQA279nbBgAlTEHp
tqLk9KMOmv2mDpWRRYfqptEAXP7U3aKTZNw3mDeDDCCW2Sc2lbU18VDuHGlYmz+ky1gO+VN2HVGP
INJoSD0e9ndhTiYDB9b00wWINTLtGO5BgCwK8sfOSNwYScwVEXwp4FRCtR0r72gHliavIIteuxfo
RGJYwH8AgMTIbncOZO/Amb2gq3JLUiByOiF2VE0eLJapsuv+TMqRFhx0nPdryoyOz/aLCvxIlIMo
YAPxuSfkv0uOsniQBsBJPhQodnpmxvIX+kOSezG7zVkrEN9E3keRq2VtsTz5GC8HjvCaqcX3gsJD
Rqbn1BxQRWeGy1UOBCkIjCskcHoWbuK1nXkmVdg44OT+jy45kUR7XeSWdBGtGrSqqBh22mxe+6xy
eWyfu59XSpKl6WqQPE6Xd09omJ7f5RRmqtwEiMGXO1TN9/vZIVw1eODpHJqdR/JPmP7/trFJmKGE
Gqgte0dSlpedsX944rCpX2oNAZhpFRF/EqYsbBrImXx1uoEP0GGnRy2n+pMGIisy3yGmpN18NAnB
GG5fAiK+hE5EdCkkc34D2xi2ALi9qY1LOW6WKcKFpLidQfP34Jd4TiEVzaMXx02ByKf3DyscaI6A
lTTSp1FO/93JB6OArChPnbVYtJlCYAj5xTM1pI4kKmeOgSjFtaHkBpGuIDJ+s8vONfrVuPdNhQKw
cgVKvt7w+o8OrA22SWZWb2U0+MlPm6SkBuFdvf4xgsDUELoGOP7v3k8Kq7PlofXQqMsvqDgHKNPL
As4A2/iSH9twft6aM0FuTuCTYzIc1sWGUZKgl+HdBrl4KkLYpFvAUGjIx/jYkahKKQmLToNohw7I
Nz0gjPs9AjHbgTMdAwK7EZl5L4LuxamAz/jaC/XszHYfBpl1fIJ8WerBP/WdmsRV2RBhXleramY4
FCXXcu51c4RpxZI9dDsfC5Y/QUs5VEwPVh0IQWNIt4O2ChhfdWXACzrvtZgbSl4X5ERM5hpAe3f2
5NE00WlNMgEYd/09hlu3xuLmc85CljmqKwsNvbDemS2GS7Tv0Nw2/rkFNGMVWAuFqvlAHEnrxDHz
GOIwomqQUQkLgBMvQKonXH80E2beY4+Y66H6MdkuPY/tujBtQB/qRW8yPpKml9pa8Q9gwLt78rmy
Xy8aqU7IgSZPKNcfbePDjXMktHbYl2SMKGc+MQ9m3Keea8ySEGSOG1LGxRtPsb/IZrE3SuAxusGi
Tl6j7RHaindmOw+Bn1qd3wSBSEvPfEapPKMjb8/FUeURzEnmRa2UoYavrKbQMcYuIUkRrw8uqbNt
0HncKHYvtvh8QvbQdqqrY6IvzsiaQAwjlNVuwYdht8McA3sxp4Tw/34FUL0gV7aknHJE9xywCmJf
S5MiCXNy6Z996dSEdUcfP6ZvjroKl8hgBw8TQH+EiTqfp4147bmIqe/z6v3R1PLL7b+JIpCfx3/O
fYtx1TFYfXZll0pTNn8Bn+fGUxF+9zAbzDQZyRndcLu6K8lmg//hXpsZFNxXBhixSn1C4InNmv8I
NUl4DGLMfvR6h9SkVP0G6GuYtFfPI7VWFpuwuze/Q7zM/5PDeUrFQcKY1aKbSzAoZH1BIP68psun
n3O09hCbBghHZJPO66nKN/jAPR/Y1UPqryVrjOel/cEVrUCBYSfmEi5H4LsA2D3H0HawlvdhXgM7
RhEYzeuh0Cvi1PLWOs4ElfOywtvT9tAAfXiuVe+lbh/YYiaJ8e+k1UtR/iJFAZsiPCFCs2Jzh34y
NSJeU1F6CjioC2JRzgKMmSTiV+UjhblY7uJGBWf/wOsf6gtofgO3L/1A1V5K/WH2eOR5lHfXEQxM
wKvfb0AyZn/WW4vftg4C63GizG8hleHR1RYunKc6QVCIkk0UPkYATe8Z9/6DzNeIosQGtsYpVAuP
SgqiRzvu3m4D0cK4hQlYPvovHyxbna/vsaY7gWW7cc3sKauz4b5eLS0CFaWxifwQz4somSWzTAju
P6xcsGJlb/VoSdQ6X45OzDvwJZLX+7vBJyTjDiah61P9vsbRh48ApZcQiQtKQNYrCx1YRMFr+bvr
YlEaSdQlhbE39J9RdtXyV1Su0DiTwH3xLLVUnrMROmNqnSVIel4KQ1936hbB/19+cWYfcrn2UPdy
1aSRq1iuOIqczN0Ykt5uOFUpY5ue15X9IWdsW+ARmT8JHSsEtvOFPPwWpN6vDNEcpNcg3kozw16y
4e/93Giz0M4S9VQWu/AUIXnCJY1wojKJU0YmUIXoueY9uPTcJQESEVkIh33AzoIobA7lPXvwhLUq
NitXUowplvHjLhmBP6O5W1p5fl4D4BgMF4lvpsSREx6BPUwBEdUps44IY9jxE6FaLV3kPwhHUk2/
qn3BMwir68Ush6ltY6egjo5exeG3rcoWnbIOYZkU3R4ybQjZBQZaX9ynVTbc2m3P9odwISlGDcnm
f37lcOp8X2mEwfPR9ytncbCx9CJvNLeqihjbvw5+wamdjcS4nCPwNsWa84KlCa76maGVotikk8/s
4kqY7pl4n2GN7hn2+TWMBKd8+U5VMWUZC3mmcTQeQm/QB7kZ898oCzDLDgg235NpBF4iIUShiKep
xI9lysS5dWiIngUfa3ev81pDXx+wW8yvx//TD1fdXXgqVlQQxBsV7M/Cv6tuM/doQoRi4+GMx8XY
J/KQ6zw00RL8EtcWJA648UHbhA7/I8taY58EpgYUc/Z1yj9tsZ0nKA4apFWcAfV/l2Wif5Z4fP40
Wcc09Fd/wtfApX23qVG2ZkA3pNdz5df5/v9339KUXodWwQXHgYndaDQVq64MQeQeqoCnmXVHmiZR
fW3w3MXARxZt2iHWnTJQjnkPYrkQ+vCAFoxmROr/dTDtIndvI9H2KZf2ceFXxHw2ShL2sC85IX7Y
N2U4Uwl0avQE4goR/eiG7/udk3v4qC4veNNHuNwiL4+mDaJJYnENl4HpNrsfij8WXkhu3jizyCh0
G6T3v5DPP1xzFoPsUdYvw2jSRQ7G2XrFwuYNFbf2R+OXMTqqMvM840GcAyhwUAJeUMd4lpE7PG6O
5C/wU4xLEkg5tHHv4GE+OaUpP1XI7L8VphojCoVgVua7M+CJy5qdZVjE/hzMZk1LTxwBhrNh3CeH
GKQkg2pBFK/UQAGCkkkxoowFD4hAbRc5wi7Q4ZQ0VgV7mQYR2vTJHr1mk0OLVxgIppiXx1xEpd4W
a31vJ78Gl+3pJkj9HHLNTuSOGRY81wICMUeHO86pB13/c/UblgDitNr/EKQM8b/QkN5tyylkbAEX
LSSkx745K3OJvdaXpC70DByiuxHNGD9zhi2w+sZWXifkYU2OL8J9WI4TcShTl+2EuLUtjhRGjcMF
xZ58Xy5xqEIh4wRlOJ3+YXypmmp6UJBgoe2YveSolRU047Mgbom8zLjK6hVOIVl5OkMEnaE57Alr
Bly+UYRxzXE57NSG8IxNUr8kWh4Xe+U1OiiGatVcPYg4iOZMRIZMsL26d3HT0qRrtKRDmPQkC45P
dGLTeL25GRV5xh6Y9ZNYaZCT36HSSbYEV+mQnGNyUU2uRsDuOeqiO8TWlb9n7O31KuQ1Ks3XhBvy
6zLKm5+94LDPyH8429Ahpbg2nqXsyaNpF/M+9JVazBgpaCZqChFv6ykfEWt2Z9ZchrjA9mDqS4b4
C8g4ft42NohzwZUVXrHzcdbNUaRkp6T90+sKHas7yVBWUSR9w6pqwfR3Ar3PaWjSI4ZLxtYRhZJi
Q3osW9857orQNrtmSFjjsqh55pVkMrKXKvypRUS//vPodit00fMX1YwF9Vzop4COAYrLNqxY1Cwo
O9INrU7BiG+gdLLbLbhvOnd6sQ2Eszku6zZ8Du15fOK3aR44toF5itRaZyy2qg798TXlQ+TaIWpc
5LX/c86IbAmcncG0n+EE2K94XP246qfUZ/AhJyYv/U5rQYgd26mwJljpJJKHZchCjxtSscnCCZxx
r4WpKsvzq2SpqtN1UsITcZDE9dzqLuMwHoD/j518wt5w8Sapp/pD1tubUsmVUy3VoJPvsOZiO/kK
tWE9Y2HNucQIII37k30s2d3AQpQWeDfD5dPqkkjEPlEVhV5PCFxX3SeJ/+4kcu9+be5Tj4fHs4iG
NyBhdi7gtqkDNmSv40I59r6v2hayS/ROqVFJSo+VklTQ8AtpwFgB50gVvubtWs2yaa9ddMLxRy90
P3hCpXup2z7kWSUeEyx+1aphqPV9O8QKawYGlTAwFaMVZFm86NYtQoEG/F9Q8TcX+Q3bPA26RtIN
T8wrNBT25Ab+HS/WVyS34dCp++YIKwxUxWywUj/qt+sy35SNTOzDJmLxPc4fz21c+0WvUm0G9vjH
bWapuZX/IRKgtipJnTerYCby53tOuzUCxWH9i7BNdnqOkUo5ChEzHXVcI81dCI9zP/c2+2AXo0is
WSGEFX77XuUpJi2yKonrAui6Q0OArvT09/BB8Rb8AJyk0YyDQtJaMuuq8GCcltRkoxm/ZAJGKonD
qwjLwtS5nAJC4d2SqWbzsnmYyxUUSTz1pUaHSOmmgSGYxD3S9us9HO+Lpk8UKjwzsZcj16vnixAA
rl7NZX6+v7dxL/pFfX8W3G1LSxJM6jQcxNC7E12lmxwy0LmItL3Pe+kzB3fLSDuS4fbj6msY54j+
DiwrhfV8hdrDyVYf8T1Hy94u90ZIEeePK9pznV3jh7B9o5mujRyiTzL4ScxsPJbRufbIT99eSaIU
loPnYNDowZzUEAGZmUHdXNyx6Yl/zYf5bQ4k57QAXmaPeNOJ/wJpukAnkwH+DRLjn4d79w+nqeNo
bQZUaN2Zvo5ySMuoX6RKi0tLAk1p1+Ppzq3FnGdUyDygqZ0byTx0Cp6VYp70rzEX5DJCubv9woKn
1o/lqy+LL51Ub0vyBaCJbsYj0Q5UF6W6V1afRTSnAHRfMJSAAKzX3/N47aQnoRTZvRLuuj1hu9jm
zLavC+8FSZDTgV0yA/xVQT8uWeI3qGO6apwPJwKdNqFdvYM23OjGW4y3mm40WBM38Og7bHTMWVfc
TrH1aAzo8dMFC61yIXSCzUDyz1JrPgvbhEHx1PvIFH65x3cTYzbbUn5owJ6NRXJHAxzsmKynEZlL
DmCR06qZTbqFomJs7apfYgzW3ocY96YBPJOw2fnSHMOeyBzpDF77bMZxm8ypT4PXxGEUiI37wMQv
1qfrgbwN5r1Hyoh28ji3LbeWgag7y/eAIlf1N9FcgCVcteUSDxgbeGC4q+478e37O071bxzIdqJK
VqXptGIDmJ4f+LcyzAa6T0dA1WeNCe/m4zdMrtSKlgXuQFLgu0DW/l/lyckF+loQt0G/nrR9Ficm
yDJklk1VGlQ7dkBERXkZ15MHUQPDXM1kB7rOP8NSpexcQahq2546RPyow7xLCnxBDee/qEQVAk9g
swMr5x/tn2DZWmDXwWDju08i/K2pzLitRSdgCWy06l+RgCjlVA27fa4OarDNEXcanUlzC+M2ell+
aoo31Enfj5Qrgsv4mrFzu+8AZXKz5kOm/E27BiQfxIQLj7zV1dHi4fz7qdntt9dq8Dt7svdIYw8I
mi0+A5/p43P2gA5Cag19IHDFMIW5Bs8nnL/iRSx0N2eBnjfoRsFhrRxFB0lphduOBn+DYHoG0LLp
1WAaQoC0vx6F9RW0fPiexh+FH9KJsY8v1UAfmN3WBDTNHUH7Agur+OzykGVM0RvAFvPkGkn0IhDZ
/XOJkY2E7z2BdbcQkI/e+N3yizMeAIkFtfgvjmXdXzcr1NJNNIolEhPYbP4zj4PE25lIFbvmWDOi
6v31DTEr+YBV063l+vwUV/mqzqgM5+YoQmewCsgbKgikMx5L1f+Au+JTOOzm9XfRg7S3w1OjM42a
/EW+gWHBg/y5sRSiHAKBBc2qBQk11ZsHm9/bOSVmXNHczZ0r7jOxiVfoxhlRfk1uytwanYjPK3I8
rF4qnKxwkH9qyENHSTIWo/YLAWlQsonbwdWrM24jsKEK5zdL6FPFzp8Xw+m0LHAA6Bc51pZPh8i6
gHKa4Ox0uAq2D4H15GJ/YZFqEoAi2RaAvHy8CSBjGJOOAuVUy5d9vv/H12pu1NSGM5/MZbCoFcOi
KD74rqDMgBQQzfzYOIlDd0VxNCcWfV16rfTjnoJtqV5ZkEs7IJXVsFoCw4ntGpTwK3/etHeeftSt
ep5M8ikVYFKpQhbJ2x8g7x7Y24v3RzFjnKt2dKXuz+MlsWFoZ/4uQP4qHQCTognrJbWp7YpDnVcv
wT9YMu5vlC75Geb1MjtEEst1dsxjtbh9Qu49wSExoc/YQcHCOkwSDleZ+OtQWB1LaPhnAhAhf62+
ymGC6NA0SXsY0s6ApKpaIYkU0UhOvxQ7eP1lmht/iPLqlXYb0dXz54TxdkkXJn4vJ86Df04FZc4x
4JUpvhIRUDBwS1vEV9nDBSZwPmn6raPmk9YEb0WeqkETiWIdIemPKyjDlF1QuOMLbLz+D3wldEJe
oHa14adDiVOZC5XWUZs9IIvMPR/5O6JBD3e/vQBfwJMSCBpVlTLPsjgRc0LUKyDmxDPVUl3HjSlw
YolPdSTWR4fkQxFAmyWcHnJwsP5lSLhVwwMI6c8GQtMbFrcX8ACRrPkufvgqb27+muMe7dcIBIa8
SheDFwq86yCbeDV3NlzYifwBoMo6jtFzATnYqw9UDWp+iIyu3H0nCgCxfNdCbKfzyUzC57I1UJDn
JU6TkV7kGMtxVruo+LtC0Wt4yobKZ6oxW5hY0atMAt7DkcfJ37Ccwide78natXH2EiYvvLKxnwua
f+riDksq83mXjOT3l8M8TP1F8VVYCK31mp5bNl/ocaMMM1CWtPSp3JVuTTE6ELLNzDGBMz9J54mJ
ohNQftS8bpGL1WTjA5QC7N5weYjcIg3CbjWzwSC/nWi7zFv0un/njkKaxEUj1nGT93+1wHBop26S
L79a6pb9nDiVgPslzjOJQdg8pNrfXrx0S4KgTXPZKr1KS1EJ84oVhEyVQtadCUuCS/f4YZMJRlAv
y+7vU6X+N+3eFvTRQi/Ijcea3WaA19bsqUxNTVoaJgK9fVEBB9oFOhP2RGxsAYvJGFDC6YyyBXq5
Od6dBlvuC/RTvn58IWvUPhW4wRFfn08YreN83fAlYpz5/GusO53Ptl+Fp/RGqoLPzEh1yWRYC5+H
JNbA2mpZeNVxkyEZjllHkomo3Bmmnwm7/CFvvYtvfA1C0V1PokJokU4nAg+GUxY4a2GwxVxHMDoi
w9T0H8bfRNBDmwUvtovsR6wB6SiJOgzFKHNyAyyEol2mo3oUtUmbOwlPLeisenzayZDAL+jBzmyL
Yw0j90NTv5lzvbhrFuowmwx0E+FDfi3BWIhxtdtJtXP0Io3aakwPUaP7OkZTjjtEnG4WUW4A6vgv
V8rlg6I+26U6V+M4NBWd5J5yGa7Gu9mt8elCfAjAx+7O3QM7OzTXEEYzk/9qydu+kMSTRYps02bY
GGDDg08eeO9jxsxOuuPl3FHY+6Op6selpHPbMd22vtLAFUZJvWYHJHfY4tTttnpMBS24Fd1xOJTW
F5xTSjarKD286s0QI8CPqcWvBbKsUmGi4BBamxChpe/OOrBj/LzxLTVhUckfdC7+rHvS051IW7/o
gs9oCOcva3nVu0a7vM+fB6MTkWOTcXUKom+R2mQtVSiB7/8+E+QpG7r6Zb18FOfkTS/iu004sWZD
5iNUxG96FZQ3Ro68yDBgXegLT42ueNUBp44+k4VMrtc20snPEW1U4+R/Qask+OibrVn3Tc4MmiMo
VUalzJ6DsxbGDX9czfIRm2nexFyC6hQK5wGgoSANCav83s8d2YWn1CDawe/JzuQNToesTkDWH4ZD
OVyERlxYaT/O+7eSQSzFiTNOrg9aDTWD+RVqyqfwcgy5H5K/dPD5evuYsgJwg3QgGZIfu6nhgyEl
ZaerJ6om/yWTfq5HaR0x80XfXpB5ZvNqElDUYE97dkWDvB2YdnbxYDt35VThBp1yfyK08tZ9NVDj
+qxpiUsnUP0QvOOBzSUs7/PE4llRlWUL8UBxHaD4NLzLwfMcIXrhHl67lVZerQLhPsXEJgSiluwx
N6tN4+QwL2exqZUlJUcjrRGoxQvvQ8MJNsRaS7hL87pNuESDHnGXWzzHikDLkLiEozx468Nzj7oj
oD+aqjqm6TSVwcLFXjganTOKl5GKu9yeIsBvX8cgrwzDTc40V90dMZEgyPU9s87m5ILso9adiNid
Md18LocU0liyVgllRQYBbXcZ/Gnyd4tfIA29ydWpZdGFEWT4uQJrVOBF2dMu+EEWltyRsJF8kiGa
bSGPgkzB8cAqw5pI39YTI1qgKpk57eLlAt/XxrAg6CFPEmodlVg+c5olQ6kuUwS5+hw+KPbcGn4J
SieBcRXtgj3bGpxg4/lRQuqIr/qEkPNMlbZvzqHk25enZM7QjG6mtmhiDIYKVDcwIfq8/ia9z9Wb
RwCPD8Z4OtJOkherCMyrySOqMrFZxbVAyfGH6vunFcgA8Yk5KAbuzuAMfvpk7T84hLqTxAZsez28
OHZfortqibj+AxdxCqFPce1QO6HfO1WG/Lj/FNTYwu3rzvEogbfRSl+XpEgaGb8LvIU0J+/OL+XT
XfBBvxyQOooyOPdPPNmKvNodJMMik7AmB3tIVaUBiUxpiG+Z5ftXYMuExtbrqCgzD6YI7XgWRjNd
a4jz0b5m990WsriFy0FyuGfh0ZBcxp4iEi4VHAlpVasGlxAUPS+kx4JTBJMcIWc0cDohyKb1Olop
sjNv7p+iLTKgXeoVVp2d2EPKndxjZ+/p088p+1k02xyQg3XEU7tCR33eG7rZs4YrRmCMk8YkAI+3
bfgxfDU2QF0HzJzAY+aojp8BChc1reCq9xQFZN90KFJDS9pwL6/2n7H/JwI7k8/u4tW+6ziRh1C1
2N+i2CPvViUTZm8l8rEJLB8E7XYQqrbSrLRavZFKjkuOqtD6VwL5TCbUuqCHjZq5MjWLIiemDTWH
2eQzDVJi8uftLcFy2PDURc7PuKmSY8hn8YNP4Q1AHlksic/CgZQhSmC1RQAmY9ra8PFbwNMhFlAJ
CUOUqaHQhQOvprTGRCiD1Tzvy/oYtaINA5khIFdg/RCtUZCSYHi2U+u9Msxvv/mLOaQp+xA5w8U5
yFVq2YVSDd6oDr02E+dI2Vsho/UvGTAnMmRTeTB3TFAV2mmwA0nLl1+2LvZQFxTNlP3QWGt2KoJS
TSvd6pxGyzJh/Bg2aFAJfoUqRwuWoMUM2x0LkQ2wsKAsqbJnBMAw7BH/mLCYGDnSKmpBfIuL9iPT
F7KJR1Bz7IkMMCdIR0p/w8h3ThSeuRWz4viHEZz4cVV2W7VeNkF5A7hHaXTetxKdA0d4NIXLQJlO
YhiSiEHVUuMppv/unIn7Skcyj8ptKyMvAj8tRVDtS6jD+MxfxRrgW64DNFGdHdjpciKNw8cNF3t/
KEeV/QZn0MRBar9/bnLTUVWGeadvoYOs+prc2zm/u4ThFE7a1BdNJrRvod3CB6Ql/jRk7Tn2Iy+w
klB7rXnhmfC1rduuOwQ+Cmqu9oXrutRL789efxHn0M7v4owRkVifk4XIcwZaJMBHeLw6cdZ9310S
51ICG53StxrDhXf4lO8pblPRLsuFlnQTN4rd27Ap5cMP4a5iweNuyb23bxMWF7LmWpUurswTFE7W
9ilAWgQnaCi6CNWzGSYx3m7IgKZPRnznUJo58Yigx1/Ntykb+MQJswmWnUhwuljvgRRQ61phXPHL
Qk0xpCLxrgRC53okOskg3TaneDJf8RkWNc5fJ+5MtlhcBPW6IRq4YySExCBFVWsA7DW+mXff8EJJ
Kwhmgv28EOWemlHmcdVHfd520lRdlMjlo/o4SYUFbBokiub1MCdSXRNf+hB7vAoLPR3nS5tVN0iQ
QNJIUKqZlSVGjOS5GEmdLUurJfIqr6GDyU70cZNtGZcK3pSgFCwVR6QTfB5sMmL6z3ecIU0LXak2
QnGwvAPesDCGIGIIhDtU6x+j2wyfl9o5qLblRvKiEW9KDPQkuKRk4WKtHuIADJHtBA3AAgDdWk0E
+BhLe1ckFSJ7DXQPpetndM6DwHEKKnPfF+xtZOmaYdqWPheNbz6VdCMhR5gkYDq+Ve+UutEdxu+N
tZ4zyqIO4mNlnhlnHt+e+n36PfBJGTFYXCINjpiXWqHdzNkeJn1B+D2PG9DmryKscuZNjJUcXw9v
myeDe6mf00kJqzURkXySBLK90mfUsn6MOpDDU/vNYohT/tyLx3HK6MO9oU2skvVxoDXuwkHEstQ5
D9kNLXT0X1IMMMDoFLTOqLoruJSO67DVt7rvHglzzUlFhUpdyYXknbcVNL/hYPJvPs7tHArn4nNp
GCVEGH545UwkNBrvCCzoDUVUJcEVuNyc+fmQEBmPtdUpc+R7FzdiXijcpH5o+NP3+trHSset/XfV
W8TVLbKaxGakLp2iuz59E4pbwE4cMlTGo3/Lxk0HbNV1GD/ajoo3AlAVtzGVdms5PjaqP48ii+IS
CRXad2mGXrVT34quP+V7pMbI7QJ9VJys7lFHPldT6nUnM+y3F8j8I8XtYKmXNI2akjY1abCCcI5d
1eXbhTTk0nroH8igaIQng60PwtU97OnqYbXRtQNbEzYDckgG0BFNhtAJ7M3hRF3gZ1hqjSVVEY6l
TZmGlfkG12YeNbFVuUpBFSXLlQxUYPbdnAN47tnz3n+Rj8HmNyPl5Chn93despMqPA9OjFk1ANoM
B1uaaX5JwM5cO2mprO3au4/umRc9Wl3x/xjhiRJs0CF6Xc91I9uATafRzXhTpiflbFHtuDcbCxfJ
Gz4/VbWdFbhGwzuLeq+uMgKH0fUJn8witYKwZS0e+AsbO3esKjC05jrE1mbnsQKCVk6++NtTIm4o
32NuNiIZCaYtVQzPjMeWVklWo0gsQ1WoQdIeyWsBEkDULbjSi5w+cY+iOYDL6Ei/jQF5uurFaYkQ
/67qBF61v5+HZkDaECjxoGnMKDtDhXhP3JL6JthdM4GYIohS/sYZet8slDyVS8kyD8ST/AWrVOj2
xDXzo4Jn1tTvMtYbHTOHoekulZ63Ued3HfMiAOejPXOW8jDpL8a9KV6n5xiDU/6T/mpZqJWoS9ks
OUnOBTKLK4uUCRDaMcZYJLjNEUrA1IAYVatJAQRz7pHMnIdtz01rvvCHM+nYnMZPCAfmQbJ5ZtgC
4nrxzQPcyshh/ZgHrcWtGmI5GMhTFG+fl6Snc/VLT7FnqFnig2kEEyi1cnfc9CnM3HWZVDxYnxz4
iRJWFqrt1okxQ92PceEfW5cXn6K38jqYWuePsdhfbCQm3UFCi8vBDoMLOoNaXKE+mVpdpJHLO/ND
aawOkn93suqaOEYz4+iZEpeSuvBjgZTFl30WUZKkklIvnHNxibNMFELSyWC2qSF9N7hED5S3BmKh
NCytJuMjb26jeGY5GNtQ0xlE1B11/4rY2zOnXkPWbX+9s/NXJGReMNw8V9esWBcTh8luhQFtB+9h
R1osJRHH5XBrJIQVpWPvQhbtdRvZoIXhqrSnbdoOG0mFFM1J/edhhgJQIQTAhgQPRpteS/nCJcCT
UAwZVFb/KMjrI2Sb77UKHxOqn4LK/ZTN//csuipkKuRiwUdexqewLSfe9QEyGvnWIa0G2ZTSvvCO
qtB7007VFZJSOCqCqn7diUFHIDED4Vmmk0X3w5n3qqt0BCCIm/SO2wz9+jmbxBHfi6UkkexBnQmQ
p6tr8vjbR8J3jFf1nPAYvsrqDBCaO3PcBRiYTPyS8pLr2mpFC+FEN+tPjpdHVpYeRIoEIndDc3kx
7hFyykwSHMgT1ftysNfyBDTvRbL5rLgk4sqry622DGDG+HlOOhMbW8AheC9pMaLYuelh7PFEdYBT
8NxuT6QficuqvpyQf2w7oI4sm5u7dL13r/5sMJvf3QyIg42h71q1cNAipmlZnCPWHDy9EP4YpEOi
2HF+MnYeroVs4bQpsFgtjlUPKCagu9wOpxs62L0GPXM4iXWQfZSCIaP70SvaSVIaJo9rwZhpAHv9
KAsw0XtMiulGIFpTE3+8KbEAoFqyeok52jVVdZt3P3MByuT8CNvABTQXaVuFZAlmFWRu4q57VhbE
zslZlMLqnglx2KA9fo4uyLPrH2ot+hFSsUye5P8Shw+UVJo+quPteaiMxklRBI4XTapIgUavDWJJ
3iGYTNdNLhV5Sfn8EQZ58ZpvGlvyEBmz4srxZkYfPDgvHAcZPAHc4a+CLQuRZjMNxKcbE2L0CLV4
jSe7+6+BGEbE2J3ugJK0KbvGQH2WnMO/xFQ3ZZDkuClb5ePy+z8W9v04neE3R4rO4YK7zpjloPMy
+NsRAuDNwLMslTiUfMSswWobvgTFxv4UE82NLMUN/Im/aL70gbRBPzrVi/XiCPQFLHqXsYHNCEhi
u41Jw1Pl4kK4rIIsBiVrDH0fAek+6ndLSzbmDQ/1k59oa7Sr/prKxZSQOayPn3BFX5Hg8rubFynA
fkdzB4Jj/ndcquAfzeje1nK8BZnq5I2faVnyEI51FFX1VVFptG6uaez28yl7mWJ3V7MDD45ZYdkq
/wm3NtPw68sQvWU3J/aOAICJH1ZH2GjThn1U6GY1w9JQECMQtfN/TYL8HZij0SGWEnZQkhxQ75jh
ml6ErKxUARYANFIAZGTxX4HdxXayBXt3UzB6/TlvrIikMSYqhv5juzkNIbsMVWxmYTmV/UMc7CRa
s11Wunf9gAC9SQ8zLjYmvk3B2ABwSNeUsN6wR5KNJNsu5tY5ht8Tyfr9VLXibvNZwvLVW95H/vVN
Zngc+FR04g7snG9rDx6sWiYhMG6jIhU9K/nSimls2QU0z2b2yz+Kn5pHTQcHC7XhgQz4VlKRQQkM
jWowirCzNxFSuno48FLHf2M8PVvQhz9rkYM+TBPNwAUhxKfJI0oP4MzmKBccKOobKCLU/wwPZ9MN
QET1SblaPHTgzdw302kd/4QTiPQp1HGaOxDE0vR4jIDiGw0/YLH5oJSbbkUxNMzLGTQRxlypO3no
DVvFd+fwnTK60UAlrrWznfhrdOA8eadFPFqvzzU0zZ0/okjqJDkmpLi9e0Vmg8iBL5HFc4GjX4Yx
Mz9jnO8yO/JafJ5GYvtJqnYvvbE//zZEOGv0NDAhUZd2UjGQwsMHyMZIxdJrf0MVKOlbg4NCyxwf
8PGYYwSnM+9kERhMiCXYC0zUgDcmOz3pzaKcTGGmy2Tf9Y7EROVBdtipHuQxMwo35EfkUpLvjQI4
FkXjfszXlMTw/117FZAs1Ftu8aHX1e/7GNYUH6G4PI82TbodvDnO+rpKpFNtJDJMmomJDOlFz9ov
LyMiz+NX7lMy38RubXWgZEeXyp0g7J90nHP8M2cV4ZsYrMJieQKFgSQmqVT+eGxXxn5g2WRQNI6+
oeLo7rRBWAPW1o9PdnBGW3J1KwLG43Jr25lboeVZuaptrMX/Er4Cq3TSFXTGhcuiyyaSjaey+pFf
8NSCWONm04WR8gqCBCgCQfBS2X1nHcrn/IUcyKl6u8mBjduI1y5FeZAR+HUjuK1Ww1PNdj/o/eLG
Jyxo2xKjvR4pBuCGj064X114nwRAoMCuTbi/ZL2MRC4npN7L9cRpjuuReXVBEciYCqA2JRZnc94G
wR7lbT/GKwqdOwr+zZwIFBmjPAFVZpmdWcmFfAkIaAKNo7ChbbjGx8lfTPyiEYy+QL4inZnPjNTd
FlNVW4/vP3WGbQJxmQuN+5EKfZFgfYmhHjJhxVeSSZwlWBwWMb36TgeZ4qBL/CW+nmjB2el+vS6D
91UaKVuzkEp81KNAZCoNDx9bsU8uQGE5LTVdviaaYImAfE53dFwSW4KG0uPlFbCmoceZapvLBxtV
cr8MBMarDqb5KE2XVAg45IZApYQrIKltU6f1TNZlXIAkRYbJfcAW6CTgjzlfmo9OTcBGfsV8Gnm2
s3GSwXwI3VHjdbHUIYvUnBoqbaaMPNuijdfmBQ8J1xqCV0gVAimmbYKWD4xgYxxttD70ICbqIs54
Du1AReCCTKbgecm3261V5xajZGx6SuOOXTeuBlRLwpFPR7D0L0NIgrpJ066GCEZHKyYJg3dl86b0
u/kDLNvSAXj51ZzZs2iRUN3/XAIs0Dn9D30qoRMpMoj3Dei64WPizQ5EHCkzkefcNMDKkWNAiQu6
aWgYF8oFAIXXS56qyq//CDsm74/dP8LARh+IEAJn+XaT0Z6No6B5YSssmowz3RNfR7Uq8SDaGijD
jYEsAu3YaIdVROpc74EB58R8XKjvfgu9ZZFEHYJIveTNLlqaSxgHyanzNBjamO6oNfqz40o336nC
vlM2iVQzvOleNfZzvNQ600us9TsLM7iIGLZ1ILZ3kCx0SxBSV7M+0rqU6F0Wz4wzHZFuyisovdY+
VwJ0VTR6aD5DYpyPPA2urp1vwQaqo0VYubsFUMhNOB//CP2n2uQRS4Au3fk14tv59SSoMNiGIC1u
alP60uo4pEKalBtdHdZ8X2cN08xE8jvhtMglMEpcv+NKNA1ubcln1OQzp3IgzFS+KVziD6JA2NGi
qlEY9ZMMB7p63PX3lFjPygIuhvDT0YAF1VmL4FBUNV0uX8FnMxZDwejFmD/sw//qjWKNvstMohse
fCzYCTnZycA93EYcyqrxLYuIiicYMYABZXZCZxbq+jAiDrg8jjXUXMAQ9W+BgecULszcnyC9DrkS
9Zj3U2i0NnYqgHs9W0MM7yJ2vCXX7HdfjacHrE2bQ/7yuWpl+qqmtHhRZJzzomer4NMrhxKo2F+4
U3FAKwJh7CXKTdWLBdY5A1nIJ6wvfXu6piccQLDoSm4mZyn1BrH1wAGaNlXyVM9umcImmufZjUW/
CFSlPjnIaxL2d6Z6mdyXD/H93bAoWwD5NhwKzVdguxkXW6or8GT/JOUWp9SO3PGHBibKpP2+304M
vE/DKF2WlGfZnNlCLKUHkLXR2p2MidJTTx1jT2+ozq8XjNulUrOTaJjXeclz0dJ2DsjnGWo4Ehyl
VkLG+3NxcMpWAjZGFU8YnHPJ2uF/X9Dl6ppORe4VSc+mQRUHixVBY2bzD6L0fVj40A5AG/ftperl
YeOH6JHfxNmvxg1Vy10EpNR3lDBlEf2/mYopFCQjkhlQJPBAUf0KnBGCUZnD2xNoyiTQLo97xQwz
ESlaP7x5CCP/tekyd8MITuCy1PB/u8CLtj7Am4NR9aDtl+/Yy0r74Ohfn2zXk3Nxnu0cfy7VHMWQ
jG+837ausKpAjE1JrsMTi4/tbjsSITPpnv+6XjK/QTwrgHg6rY48wob4m6Ae8di1LVtmyEqEqYeU
X245Wcm5J5tK7Ia7MDN9xzUEueX93mM7fd8Qm50EHTRngyjFX392qSmEb43Kd/Z7cHKJbcSEKBiy
/iVhgTOruP5Y6m/lNY6vlObgcZvzKoLPuecF7u7qJEZVcEDd8lMrSoBwUk2KWupEJ19sGRV/ZE7E
88rzLWQdujOiznjBXTEsUDYnhmGPNdiusAjMZr6MPJJ19kqVUA/c+eiaAHvzwypnbXpfov9TOQfT
rIvsRmU3BQa1tpbGZ1zpiyB2+I+Cyy3TR6UoShdxGI/iZd6852bXuHpjn4yoxX5KDBV50EJsvHlZ
eYxCVXQ9mr4ODHeYCfIFS48oS9Ln4UuINtsiU2Tr2pBe0L10Zr857rbegEyKQ8AylisLQV/N+mJT
939PvD4b4CnZYhcyVQMavhbgvXljz9gtvdXluYF12qEwUxF6UxXOBArmMVYnlk83TCEhImT/YmyC
5NZJeXf0xv05bNuHSYPwRdG2IGGXw2tICrH69ZBTaLLzoEmQyk2uBS+wVgSgAo8pcmkTqusoWOAe
mDQNiu9RZesKmtpq202FvB34C7lqh0o45GvzbUqVRwSyGdzKQ6UQhh4q4iWAbscBHF6QWlk8wjrn
53r+HfM9f1XEHAswAUzhT5CG4nfIFaovZpMQMqdyr2lhdsO19AyYJMQBIIwaCYHweH4oJthVDfR0
VmtK14O2NoRtOhqEERXQ4vreB1WjbjIU3wm2ShHVoHJs3F0V/4/SXwEkBLEz3H9roZ/akukWjFJA
xprez6LsJmZLOizReAo3qATCARQTRu4s+o58/JN8GFebiqWsnEoRRi5q8dXtBOGTncCgDQMWnp/z
6IGS7n0hJh5hj3IqF5lT76Lc//ZuPLjJTa3s24wCsRpiFajQeW6Bu45iMxEwLfiTuemNMMP4uREM
N8+IzGBp9tFJBNPXNs9XKLlKyIS1VR570Kk9Nby2bWYI6m8PotwbSYQrOlj+z6/5eRMNCudHns+F
ladgAmvn1jJWwRk1CpyVXZEFDNvbs76QKH07ghx2Wpk1naGYAj+l3h6mPmeztWqgBKCIlljLqGg2
TaAP/bioyel9NUB0PrEK9BJW6Pfp+tRJJwg6vhJUJQ+P6iobXyJczH79r09K+JPUf+SBPYxIOcLJ
TVUHL0dJ06I8U8m+FikV/+EUyHx7EXnh3BR3lExgxN+I2d46K9mtz/CH/1Teb3z8yohv4tqmK4pw
e5A5z4FoCuO78fUqgIx4YnbekDxYNRe0V3xZAKOzAhj7hdqTnJ+QKeY/3OCXoZCklwGIoUmgbPJG
7kimKQ/104mYImFIcsN+HsNgawVKxYhHxIPjFGA0I2gQXOSrYqroJPgYJj8bpmkHc/kMciS+qyu+
gq6M+oAZdslb7KxU8uDhyxPD0JqdrUf4dzt+zC8MK932PIx70kE26EUlra5+FFsXlp+PP7w5gPCM
bCkH/YcJ9PTbiEZ987NxxXdbyJJLP0xj7iPWghnfXrOQ5/TT+sEL0RIbuVIu0jGDdNkfb6QmY/Po
r5ED+tO5aQSqGdTHQl2RU10O1PoG0tuQRG9/UkLJUChNfGyEjPv1QA/Muu2Sd7+yUGzhsZcIgJmZ
2bWH95NquzXN1ge1FvaJyEIDxsJm5XRMoueRKZ+Llo/r8rFiioqE0Q75HFQk+ok50obD4qxWFqxd
2tlZ2trIBU8XQqczhRizWv1eFGs5Rb2g+XDzxy1BxYfzosqAF3f2HwsEQfgb3/L7k4XkqZ3N+aNj
2VsOWvvwRCz8f4zfJtYhit2cZbFoKzowfLC/vpYwGThX0VAIzsP/DI7j/DF17MEP7p4hk3OHqiIm
HApYi1VnW7rNcUvKV3gROibZJchffk6u5rYh9Va/q2GOE8E9JcDn23l/pTvv0MYKvWSLmPILPOp9
CNVkxRxgvlj5noERiWf2cG+NThIkqNrER4EuRQfwLM25MHghv69O/qYb+9pwUhdXyEQb3kQB0Uhr
kn/DlXFN0YhAh7La0Pnwf6IBkfqFdUsR1G1CdeptA7m4TqTtZmLlSYFIk25iQNhL6Bhyvo7eDMp2
hEXq7u3Xk3qsJ5+UEQA2EFTtKyJDzyVe/ILk+k5U7rFCQQpLpvgl0kafRSZPOG41sdlsKVe6VkBL
Pjs7DDpHCKGxx7OijuW549unotA69H1eP5tLMQ+gl5UGW9+jBbew/Jm0USUDSRqToCcDEdth7VJw
ccLaHiIRTko3TYULLRhHSJB8SRtOu362ZLHIe7Q21tMbqXiVxin7wvACxv47jroOK/he89j4CHMo
ymkkfuohHu92CEWUtenJ+3RMefDA+lCEXc53hGlLLLP5DkemtirVbyk721icKFVpGDDa7C/y7yl2
6VK2pegDZkIwLcBw+Kb2ThZaMLcV748RG1jZqzYQ9V0OHSJ+BJZv4MbbF0WqNjII9CczlHiZc8XC
BKDvckUDX7UQOAbPLjxB251/rSYjFXsLeETeWTqi8nnd1wzkn9BSh5PIz/pLiSYjMQp+C1sfFnU0
Si250S2fs1BQ/qFDHdwyoAL6FOGWAFooyPdBe3Ho+4VAkqoJgI2M+SPWLdu0ZiBhVqe8idZmzaPC
gvu+PPvyk8ebJ72SUMdlhZ/y7lRpubuP9PsOrm2Nm9bIpLBn4NsqrNsE9TYVPa+eUXUmHKu7CHzy
k1KsnQmuc3ocbf4+63MbdyFsN7VNyEyZpZmrO8soEvfQaT7hJT7MN9CgrWrdXIrMoXCW/2OmYaIM
QtiBuXK66bsNG6k4kN2V0XObem7sIc5+X+juVdpES03SGIoYEMoLbW0R0L1erLM55dTYqPyzQxGP
xxodZ/fKRh15DgYhNeJpF6BDtK+S0FsZ6epLA5I2/DmIcsSoVo1a4bQ+I0xAFR3l3VChSWAmSzjB
CJfhb/bMNlp/HSt18YlK+tp36hI12hBcuvE3XQvbcUBUTyGm6vKtLa6vaJnnuYeZqj0pK17Y5KmB
UlYwNcbozmfWXxuRaseiEG7p30qB9uU3tabAHLiwO4Pz6SZ01t5+b9zNCCeM3Be9tdMtn3My+ak1
q8rJfNACBC7dcUkMmFpPerXY9g0VgqjHg6S2ZMQgZv3OCiEgUHdPilVH1lGNFc1yF1oeMvxfz6PL
WKizLqmMTzsw5WsVjEP+8ti8w3KKjnIdJbBf1qnNaiyVgrXvaWOiJ0lBADaUfzTroDQ4JBYhXzu0
zIIzN+Qcbm8O3DJCk9ynsLYRxYPc2piJ4VJ9wsQctBpvbnPLtbo+7e8ZvvKhtzksKx3rU5NlT0aU
0Jia0GarFjgPYskfnX9SXEUD2qgegELpThVwUMp2BMw04wXl4nSyMv4O87QNax4mA3brUqDtZw8R
7LVOic1sZYFVqipXO510fH2nMuDUkLnoW6TX0Z0HW0vQEwVkrwrPxzrD+eucPmSr+WztNlU7nuPA
ITlaOHJW6ehmPEjc/BNDBY/9yrHkJJug3ekIttmwJ9lVscjRfkaQhbFNZKv4EnyyYgkgRBI4NXRm
n5KLZMML/Z74/hbyq3arzPo17Ykb/FePkb7FuZuvQX0Sihzx7Q/JLGZ3kY5x31V51UwK5OQxfHDY
tJGkBf8IuoSHzIXUyxLohjBJydWPyMM3BvWlgfOd7LR/ntuRT2pZQz4zZAPVtURL9q0X909iKHwx
mnzc922g1jqF1R/GSLEA/GTNiT2emMMwxJ+WANmNSxG0FqEwO3PEe0xeMxeLcQ4267s/G82BX1sD
bChUzxJCh5qDjKf3P3BXN10hT9zhhPfLkPvuY6Au7w7t+wQTMMldgBCGmejPm6Vva0IZZUmg4N4h
c92gnpb/fzkOudaexe4yk6PmubmN+ZsdS8n8FfbGg9CHw0OC2VVVh1y9EbZ7ttZBnMW3gFEcqos7
6sJVATFRiPONHXh/FzCKXL6j9lvJ2Ga5GnWYcA33ZA+JzU+SYL0MuqymAu3SJQsit5GWx2FYhERZ
/lamuPyyc76/4Lw2rdgas3P42MncqqWR3yUvrHoiUCPXWfY/LpaljiuoACqJ1V0MTXCSMSr9T7Se
VJVL0ehILgdEl60pCfDoiSYdd11rU/fftgz/rA+h+kwu4v6q1utbjcDcN4Y6w8+vcLdjwy9XuSSL
NbcknGh8CmIOWLiSJaNe4ZiYqUXKwTpAtzNYTFrkPB9gJ+4PleqqB32MBv+wxaZjhQ6hdCxT2XiD
cz+8BVGW1PExh86kjZg4ZcDS8jKDlaOdFO1fX+RUgDzN/zlbEVEniob2eVcN7TR/FdllUYGi3gwU
KLJJn9XNbJzKM6vvLZoCC1+PXVDL+Zbf3D3FQnJTlJwERBYrgpR4KLoUV4Btdk5JVbWX7Hp6Lsyo
0ARjWNgYuhu7I8JbxZhCKPTL1/Cc/6c0DRABbaS//BO9A2RhNAIQ+Q8hIXRRE//+GJ+GK3cS8/u/
e44nDqhM1y/P88fsCmqrqLM0rQHcEsL0WpqRllDAGy/tPv3W1AXRm4IvelfG6YwyCWMmmAjwLCuS
Z9vF8PavokNmplihA1CvSG5hqMoD/sXaFn/iOmvpNk0E/RPDuS48aEFDLtjEkt6bhe83lyi6pY7d
pwZgJZzgwbluLLLWAAh7EfxINQK3/sQ1I4JzumMBVN9hWjLQuVfYTy768yl32WP9uoe2LvjUycdm
vENDk2NU9og8WRD1l8SyWyXutnQN48ItbtdGQxPDpb8WJVTAMlDTGLDZfv+bVOrlXzz3vyqO/Dul
ebdws3lpGpxQ3XbrZsSuJkhICMiFtbuDU7IaYqRZOWiI3P29J+O713F48Q93NAIeV/MI/Vo52Rrj
1mBvdPBYEIUvbMTu3wxdrEITGM2WTrByUnBWV2SbbpUMd9Krub7gkCvOO6ARXszcOt11T6FkwRjb
+r0kNyWZ9Ui+OETrRA9vHi9cnn3NS3TCk/Un7hlh998C+qugSJymFVUdn8lcbYTWcHi0ITrO/hnn
/t8qh4GhdssBObGL+U+UI8ND37Hn6QOgkV31SpraHcA41O0FYKRC159qeiLPVdxteH70tLLv7Zy6
80AaSkaeFrR0z2fvA8oVC/StfOO5fuejPnBVUEtfjk/kEXJj1nIpf7e5S5cqr71dUPkHFbGiHPnU
sCqJvcBZ5as3Uq+ODmm9hjU/4kjaOlowR2xRaP9kXjskIxG87wyIxrh9hdjCQGOl1CZwgYoURIfD
W1uxP7KR5H9qOGuX1dM4YIvdNDoVIACDLqjbfF54BPUActqPuyC15e28hJ4YrzuKsmOl2pdMW2CJ
92+EyIQwD6O+D0u41Xwobh8+L6tCgpsL5EJJyTMKL71oHqZ1B4YIoCgMdVb43yImNyU/uFY2jH/R
EkLTdjVUnsAUns/uc4DHqyvrDiQ6UOGJRgVX6rj8X/0Es6lK31O0NjJxNal3kxrQn2QGibf1VBIS
/STfeR6n3UcE3+fkIzf2AHO31x7rIIYU7/Endeajg2jzc/S3vrVXbY1PxOY+C39/FW+02X5PIOhV
fcUpqiaN+In54osTRVsMrg3lwnci7YOj7J51iqemsbymvcGWeG3HgULVYyMeQmSk0+LfgyXKHcf7
bVjKP982UXeVgB04Xo6Y8nMjIXKpXG3IXZKyPs+Sp3ohyQIN0TtHvT0AHXZjwB3HmqqpPM9M0vLc
simIcmTypSMbnXVErET0TI30MvkYqtJZ+WbT477doM7uCkSi4wNDOv9CId1NcrHZODQyHP/inJjT
BD/9SdXjHS+5Mwf5RAMFgV/DBjTCxhAOT3dZxNOYxfQvJ/oUzba4o5CPwn5bzsaPfO6DYh0bkr0e
kgMoo3sNabCk3jMAT2c9/jKX4rPdEkJ8t2LRlO2LFsqbc1x+Ui5pzboa01c6tBX2DZ+PNvgxwgCu
RtmqA527/nKhmR6eIg7cWUt4wfwkLFpxTWpRWPSDJKJ8Jn+uwqw4L385/AdQmYfmnCIGC41tSc5E
Uj1S013Yiw11SWbd6kwK9p9RuM3BCg0cOT6PzJZP9UlGciE+6H3hq+wQD/EtxANbYFJY52ea5ZPQ
zSzPzDl4KrW/Kwy09fzz3I+t6bWlIRBL7mE2L4tAXaLN091lmVkOUfINmahVK0U7Q89m1mFWBSUC
hE//98xV97Q/ribkknzu53mabruoGPcGNytnaRc78zLbVWviqgviZdWZuscPaPNVINeeNj8FMYuJ
K0BZtYDvK/ly6U5VUWiTkOFkqJf1T7JlqM2ItVKCbUpRp9KrUXn9WYHXLjcx9BvfTwegCrrdtMap
RNo/Xa1pUYi0UvBRKgO59+15v8bNPnACfCi0FlfTTw7N4aS0J11e1yVq4LmoC9HhQwBM0AUdZTF/
7LokVlhQ99zxPkzGBZyz5Xa/D8EOZ9uqg6E7IO00pidMXEeCOIt4JP8zY/knnl/xbiMjrc9ljAnX
R0G5iM767FgI2wmSrsiuUf53jF9totqCcxaTCbK4RphidgBphxMIRveOKpqp/h847IikwvmBSVRR
nLoRbeUisbzAgHQEeFXIuxTEdiTNVYhLAA0TKCOUjJ+ezZ1giDH266Tdtm/P7gyO8jxJlmtNWxZE
BM7mTH40A8r1HkUbtw+eesAf4Dv6lONzEH1qC1OREdpZwVilGUxO1hV54hcSuOv6wZYBbf6d2dbk
BnZofQodR/JmzGT0ZZQsWKR5ZlyINaAM/j+Lq80PDcFzWSu0ytipUNvhbm36egXlATeH0ipE4nj4
qFt4CVBmKvTfF53NxZegxjgZYgjRd0NzmSqRTQwl3jG+HXJl7HqhUfIJfe3V2t429cC1A0Ol/Gep
LrQmGzWUew7svQhrneNjoGw0/eRNehAF/dKdnVHcL6W1zo9PEITJBC+VKMLEJVTHjHmHSYG0tV/5
pexMFk2gr7mxuFZjkWHcLWU6FrYsIP/4MC2s0ZOV7caFDRUmxWyiB/PzDwia6vlxcefrPnNonfbw
aU9uSLOcT4MAU3PwGth5NkLpWsanFhewtvNYfqUyB3uI51KSWL1riQZliWSE2lsr7Zmqb2vazzXP
8juylZJwZh9PmM68Kx0EdlthjusoyIV9GHHXexRjqmdCqbgZjax6yFrj/ys8YzWzHffNTwTCr6sr
KlpVIJNHckalqXbfGEz4i2o9xIfiAnuhXPqc210bNFcCQJTVUj8Y/iib/fQ+Hfdwk8ZASyTJeDKZ
JFjAVeRrhCAIanxLt3Sis+TioRWWPxERFLEgEOup+WGLQgAS5NhliypZZoiHRemseJktQ1FxFIW0
IBvJqErfIRacw1l140VYIasV2jez28R9f/PtHq9r0eHnEtLZTq6XXnQEnbX12qF5+gbomX7tjRcJ
KMLYsSr6MzWRgMOXPUYryLGxmCa0fIy+d3CYooZPXkEOJyTjmrAuj/NTpzBu7vv8ushV3/Tb8F4d
R0LsrWeFSLHfL0iW8OfWDKjTRdvFQJzUgNQtBWFyvlbLDV6gm+q7K8pDa7/aIYVKNWKy0CtwZB/H
M2KYTENEET6TS5cg0I7xBtFDItgR3R56JupIMaRwKgYg1iPh6Dew9WL0BvFgL7yDi0cvdbcaWgVc
QWhWv39t85PZDm/HTuE8j59mi5JU0lcH4cs/JVl5laRC1LVkv82DI7OV2H+sZHmjhtsi+c3lzl/1
qTJdQMZhw57iWZuIbpTDrgwGhM4cra5QYX8wuzpgT94zuAhbt06bTG+USOkswRvUesGpC1nwejrB
K179DTSlXj2pWF7CAPk9+ZiCNuYQYRXz8LO5U7bCZgwiKDokcPyRNe6453Fim4nFeDXNRx+FrUBs
BYWCiUXjEoSlsh8L2TXRuZd7aX2stEHzHrX0rrsj+G2yddrCTKXpGFyGLgdU8MFP5RUkISDqlLQO
a4gbw1fXRKqU7t4Hrr+j6qgFN0HSu4h7gigdQKB/xw2G4LwejuMEwX3AgGbTzNEiFLUIGeE2heEy
zSb8nJyzW4Qtb18I1S9k348oefEcS6fA7w009e15UgumFvdh4NuUguIdQJZvDXhWFOroKASxMvoR
SsX2NepIxH5aiglPGtbxrgDb0+e5Rk4K5g0MsMAVXcUPiXO5IIgnWdGPps6iWRLWHXdR9XByCfT0
J1hHa7+JQC3hlX9M4o5WqYDQ5KvIqs0ScG9CHfXfptetOHqn6cKJVNRJ75djlIe+t59z1g9zmM75
06cyYcJ69FY88q9ZXnoRFwfSOPg9qThM5LG2Rtf2rsLAwpK2K6XAjYKvahxGww8EEno/1JLDxKyI
0+RfTXg0m4Y1rKLeWFZ6oPYjvI9fW3lemwRHtdaDGTfPoMzrINpF+fwcT0zK9Lts4OQjrYSa04Of
Etr3+Paf5nNnDV7OVFSeSDQ5UE9140az+1PsWIb/idakcgNN2LGMDwqKg1LxiE5fFGU7S4L7YkgB
EMh3oUOCB/iddGQlMRyYYxTTMxRCPbUD9Y4AyG+jMNZxQzpG+1OK5nWPOAT8DyO1R7r7T1xjgUYB
ZBYb0TLn/VlPzy+98pVuUvW324FfvpJd4BdtTLpiRDx69Wewjb5OfHPSKEUnoa7849/bZh394djr
tIlocIO/8UkjAKoafNTcD2FI228hYIofr3Gg3GZGN4SqFhpenGV1Z4hQsS7g4SUpflwVOeRUMPcE
c5MxWBtH4arZkTmtFJ4aFV8CuGVUVHQwmoZtAVSprzzaGaIo51QXHihDmnPLdWGCmVRsXmGHmNY3
ehtvele3KGsh2PVoe6bnulVv3jlHyxaIO6o7eUfMw4YOUL6NZ+Fz7KgFvZe3xPRCEgWdayTziLDm
eGObyGXwOP8NOggHh+W+Jxl1iHXa6TxOhBxtubzQdZodSVNmgeO/iOnJ8b+BdWuS7v5Pjk/R33hf
2Kfn581moBl29Kvgg4UPRJaI+PcvAK86ml+SP0jFWDA5abEnaSLziT7RXI34C4FkJbwU5HeHbq7/
50X4sHRjXtkmxZaJau5ZUZ+AKAlGt8JRdooQCZcnhKNu1D+TyDrDgBQdgGqc6diHjUTCatKdl2GF
G18gN1NUJ3TzSb9lb96IexApvvHnWF2QD0Ltb5wC5CSW4hGAMIYjI8PZXpM9IjiB3UjM/RHAcET4
Na40Oh8eQaOZC0QDKGz4gNhYkRpkWEKComLjXBUk3+YbFyEqt/8HrEqAAsvZTvp2Zy7gLy+sCVTm
qYN/YFSUc3R4NOOwvk9lKna7V0Rz5Ozt+oq2o3cVAvdx6zq9S6LtIkYc6KbWLqk2xUeVDcZFSVr1
Lv8uvf+VkJgYpZNzp9t1u2GF240PYwIvvl6zltKxcmKYs4f8UZv7SwMDa/auMBJ8K7oGjfeZ0BCH
C94HLVfnNMmIt2f32XM9//Gu2SN+9UTs4UJJSWh4Nk3M58UL7z2UME/CsFSsUroj6h/HOqS7I1OI
oM6yzW+dnk2oZkflKkqc280K+tqJ0C0SR+7x8WS5IQ638I5cPgBo0u684AED40IowOtl1l3DJb/E
gThs/3aSdEmFkyoSJRrJPqJzBctaFCe6Xdd5akOG4gugYxQNnMgxxNz5twKBI4pla6vGbt9js4t/
/jTFjQ9DKn7wL03A+DqBLozd4JtTs/NKZyOIBIkfYL8+hQbvAvnbt0dgOqL7WaFOdou6hYbz3dlH
jSunGZev7q13/HQeqmohhN2GIkBOWpNMUzOdEABNwp1/nrR0yxdqSqPjYcVs1ENgwzijlaFwphOc
V5Shx6HlNtfzlSu1NwzhCMXS0X/aQ+kl60p+fheBOpq2cHR1Jh2ypEnhsJ8NFGkOQhYlG1AjXJez
kN+RSV9dJcQld7xNzuWJwy7Gccd0a+W7ayFe0PibXtQ8A8qR2tE+oKNSq6KAPOmpIQ76zWgVxnP+
mzpGeAKPzgE7eo30nrSoZfAZe6nd/JAMH73HfyFX3NlgRszS7tyLZF1sREqmVVCLRIdigSWlsTdh
v3bkOV4XZbfW50Rr9U4pNdpeI28bDJAE2Ry0NnZBLZ4jNIe8CuCGZskYYgYAbX+6LGLkMW9gglZu
yeDnXta7TTGXI5Eh5UDzowlxUAdmAwSSnGRpQUcjX5v7gddUNv7txgpcTdqhYmyi/XccSWYwGdFq
UpyP8Pqb5GFWsDgcUKea1gou1rZzDiNLNZ8gAzXf7dpkHTHrxV84Bi96dlu0DfrthMWtq4LiSlAp
nFl1O/alOg87X/rK7yXDwU+hlCyAtP82N9X6FR0y/pmO5u+eITYBOT0QaDF5sXFVmTKaa/UW+DtX
nP1fl4WtYEhtKPOgk3oL4fFqNNs000I0HRMnIanBCe3BoV94aEPvoDttW+aeK0b08iTFgkHpi3iV
AR6+/C4v+DcjBFSvb1x08wbRupmU90Mj2cpoNnvzgFTW2RSvuVb138PSe+0sRGzWwUBji0CpPSMc
D3HOeDjP/KVRMxP1kZEDnkO+XTqiUFAqdfQ3mrWYKRz8xq+k9MOjjMp0iuB36422QXp+J3XOjMnV
mdYUXiPFrGPYvgP4AvlabCg+RlyciDqruLPtJuBy+r5VlvO9FWArCRBnqiYCA8AeL7gqkd4VkkIn
0BouLS3BLOFE9JyOM4Rry4+wn3UtbplkLE9LOxtErXqx5UIwvGjneWZE4372bMt+Dd4a43ZDA2Nm
B1DA5gyCEB1HmdvBSxP5iu0dg+MNgO67Kligrw6nIOmD/7MjbHFLLHWf7kPIz2uPG9+E/bTDijYM
zxhf8rU/82wAprmDwa/ogS7JldI/ODuz8IsZPc9DsmwRXNeh5gOWVF64BXxbbEKWVjjIygf+RWCy
fQabn4qw1Dca0YlhTlSHfEGGJod2qVTOaNelJd7BjKLbyI+GelQhuN9M/TCt/i3x5n9/Jxce1Oel
jen3wo+LInWVU+KeRs6FuAAjbaJinreMsIeq1IB6MFkEaI0PeXFPKpXdJM+gvWhgj8rD1YDd3Y7u
D1oWrFYal3oWhk0Yk5U3o8FshJM2CgguBLChsOzxQbCz6e+J7CE0UUgB8yw0eWoCaaaq9oLtNcrw
JbDOH0sGyc8/cw+dyYCiyB54DZhErWEfGhblE1xPratZO2J1aeTfZI/8EfHKVsb0xyugeaiBtA3n
beP7/agVePB78sU7f68Mrfnc3CtbadQmXnWbmJhQ2kH9at2sZYak5KkDDkBRd4Gvb5ErKIV6l+Y4
iKxNPa2lnPsxALloo5c9xABsRwCIspFmPWfgwNOJ/Tgkagk3VWoDdOZw8RSFOLFP3ZfllxSGAPEw
axwgR/38uaLlvqyZ4BFuSVfu1/NcljN71pdHzCT2u0Rf1IiX32VaTsx8ncML7DNMVo44urjWhknD
8Ni1p+5Own5nFR9QpxwkQZqweWVJHoD7+U4c/C8Y+/9Rvu6j8Wf0NrtE1jC5cVTJI+lTYK7IODrm
fD5kI8Abz88bRlgNUYESAgU2Oumk0VK0ZqcR8axmC5NON2HmtdKArfsnA0LuggH6UfalcGcmHd4P
3iCLSWoxbV9x08PvC9tBgg2f30VIXCVjudS2gkeso0/We+i7xsYky+WD5h+SSiCwR2eD+SLAiZVq
B8sEcfu3Tea/ArvfzoTzMpkDOftqXYoiP091QgqGLgZZz8oRcnmvWi14I//3zE9nla82mkmkKpkd
A8Tvo8QncpdRJYZc1fJ2AZ/gdOFS2Jka3HeT+LtYWyZdHQZFXom3g3QdhRmp68A2tCLd4dat0M8g
a15n2XCpZqXMFW7ruvaDrHgVw0KQmT0kdnVIyrA3dWcFO8bquNJz2rteXWw/EDpHjH2PWXKUGOJC
C64hx+8drQSDU0+kPyRMiJVeXbXxiGS6sb1N4h+02hYoBIxExlZ8yfIydnBDqyolfJsYkDBo/Ooe
8qh831M88CAsobp4yINpvTSw+3X66ve09XvCrAtuqk/x+k0sHiipFjscfnGcvL8GFgc/0wMjPlRl
CGX9jRPMdUvSG3UHx5iOBZ+iPDGQ7vv5bTGvqjAvkISw2ETJT8Famk6PUcP4QIuEkJjOu9G47+oR
492WBAgUlgRyOL7rdWpKoSwMWgn+ZdlExNYPrWNMf0J8ASgj59hw658WQp8PJC3mUFflzIosBphm
DPyzgCN+mER7XrPCL+/WS3o8S8StY9CMbsSh0njG/n/rvff8iZiCMIUGW/F7trqnLUM0rYk8Y20u
9JX2N5A3Fy5Tb8f87QRdGb/Z4J3lgbIif+LJKwTJzFqfKZkxv68UtVoz9AnhUrqGIkL0quu/XP/w
HwA85sZFEIO8lGJKqAksCg0hYy3L2SXPRx0VqUKD2u09JFcUDCdJ2tDP76DmgsncT/5aMIdVFeey
KCNS/8xlABEsacujj6plPjS+Vv5IYnLSe0o+CQ74HGxuxE11pjYR1/a6TucGShQ6GE4/LnAodHG5
dxCIk2MO8MJ+W+HhZdfP+HngPx+9JLrNDOcYCMaxBUHdmm0GsgaHyBuxfTOMfynmM71GRdKjsdOC
+aroIHAEZ77/e9i/6B/5xksr+yLIEpfNLMf5x415gn51ufKdtqZFKShBXQ4uQ28W9vcTBuDeyeUo
ao0Tlzr+YbvmcCctZE/gj7cbVMxWVcL68I4L8wSgmlm8Q5a5PN4j0E52ww2O70Us026bFRC7efAq
T5PlnBuLi7Li7ffplUfBPls4f9HKRFrWXdd3bOVLfFIsegHOaoqCNMrFhArCl10mX17nBvrheniH
QdwNdyHf9Ng8bIHcuP6FyClf64q8bUv1/nSSwK4LBlPIwANPuB8cLiYG1v20jaJ7OBFY6f6hD34X
hXt3Nw6SkNdTSAYuua8r+zBuvI5n5xoZrs+N9dptwXzjd/Z7Xs18WXYiGI8+3wlG5aOchWVSmKOe
isoHUTADrmjKyzqHIsiKte+gn/uPeEf7sxKtO/xTEb7gR+6iaAYsMrszXftDPgfh1Qa6b3tAryxK
z7B45G1WfdgJepC8sdEsvCsL1XzGCnjfnBIznO0hZZJ9pcxu6BINZtODJGTX2xLln3AXW39tvuvQ
80bxVP366JDbOW1zO+XCew8w02Z9pJeGgwUDUCjh3SVQjO0lq2wVXvmMYduy9Of0llYpsYF2n4CA
krRax/qCVoa5a1fcZK4J98QsW1vALZ913Bs2rNQ9+iT7E0EFDvgiO4I8S+pqeXhXmcymf00E1mYo
28aakR/76QNHqTI4qtGpzPcVB2kB+UGgTa80uORbf0RKLhzWhMJgozF4/XKeZS6MC+7hAMc3IUVc
bO2MOAb2PjZikFmj7w3S7QmSEGaBEUsxUTXpHF72BDJGWSWAuge8oUEP/OI/YlvTKY0zghqHk7N8
Xqtfrbt5IXHqvLB/WZdg3C32IGwr3+M4oPqrTemuNXDDH4k/RpCMJaeisSmdidum11Lnq8UEQoOU
kuJOk3CHEnFPH0sV/Hn7W2TrHvfonvtTQI0bCq+XbjbThjmWWZt8bbpeHlkN8Qev2nQCREjWeZNo
kAICnKrPUBKRIu4Zl8vq0hR9t/IIObgdxOV07XVxdz6cb3SJtZmAAVqXHsIy+2KPgjQEQ6laQaze
gpAs9+/dEzkGM8XMWfNJ/HPVJ0rQ933+4AvOrsTOH6Xhzlc4ZeC94P+AfGnzisiU7bauEEGBuqpV
Qn3mDOwaef+dXHkbp5TOGeLlu+yGfZTfOWXrStEJF5NSMlYsGM50osqxyaC21thvVuxZpAwmxH5T
B7Q8J+lDARv5C4FQcohSBuoFT/pd+qfVaO8zqpati9AIep4aXgx/Qstaa/Ew0geIQa4XkUqTn/Hr
W+4lUKng7KHXv3CaTNvFtKmejLEuDDcUJTPyM/Sn/4WoWlJhL9qfrfYjMLcB6QjdZo2NUHalbUmi
4oFc7ns078DUAOn+1QASfVCwu3t0xRjWP0VgV97xVpHdzIRtlfVdODzQBM7hnxhOP3LX1YKpEpww
qSDI6wiLLtiU/6e8dLKZ8b7o/Pk1/ce8cqy45LNCaX9aXrJ+fc972vzqGfZcWsninLMO04JNRZoP
/EBx2gB543aphQJTcnvREkZdiiNlpt/uvNAso0AYcRhruYslNDvAHUYBWlNaWah7sywa9LZebwGP
vDLPr/sXAvr5KTfbXNPRiDXEImliguj2Wszhop+w9GnXzNSOwQ1Nc+3bJCzM6UIjSP1Gs2FSlClD
YAdYPCTKOEKTL3TBfgzxB3ijkdY/6/R95zUPjVDjHUXlJIbuf5PmIjXOxxlyoLF20f6G66I3w/00
op8Lpiy6k8QaCkBQNuwg63tiuzirqRHZdL2S4djFsnVNngdbBjws5weBcWv1g6J0oxiq336dp+yh
xV/x6F9/CkP4xbG5tapuNcga4EKBEefRcifQUttpDAvV2xkn3VdrSrkSUu2OXvIebsvUpRl8Qs+w
18po3AoWDZZ5kcrr6ODvV1/qOwCqwzr9h7vFPVkHdhymPhu4eQXCQ/jyiVnRHPtwssfc4HtxvdxE
g2nRFvyXQPPiM/NPOtz27JfOMD3nv/2s1YCKd2UqYcpQEJ+NbHZSO2vXV4KGxeALvE5T7gAmF4ym
WnMeYLufuPE+XcO6gdL3dyl4VsXIj8/4nLBJ0eo0rIAkzZLF0W3Ire0q2Z4V1s8+xyzr3OZcrnrV
vg4II7VTOa2m6EuyQbWY3fYJ0cF6RZYglaKJ/o64a7roiUuHuRNlGKhT7XCu+AEORa/mYQ79Xax6
PtVXK6DD0yOZAqBkm3C82o6KSdq3ru+7f3AWN5lCkJIuYZrHCz15EizEODmyBSrnTrglyWckPs08
eagR1qIHePuYi11PSpqO3COfbA3QvTy3M6XBZeIvpP2KxtxkWVSDR7tyzQTZDAgALim+dQYFsXs5
HV/tT/zqOlHWf6hFZZaPWeJcJcWfTkl5SWeepf103/c2ANfevdbKba+HXvmL0LZWcVuwFexdMmXm
uSMlaN5dI3rKWFThCL3qtgv0EVUr5pYiwEKqAAYct+ZLm5CN4WeR8HSnifgchLPhK3uzMQ41OCVs
qEuON4q0eq59muA2wNXLfxcxdRXX6jaPtI7zHCo/DG00OqRHqkFcgjevdPuOF0uP+dWFAhGmqaNv
+GSddsEh3HLuVKWWE6oA/+KAr8vk2qyDD60PLWMJOM2h7QIFQ5Zk4v6u2nbTWo1hvHSzODIFOv0G
jeDIwKZ9nBuVtqHOcM8XOnPrh7wgJREPKQoKaUywdL9Bh40bLYAkxUY7gd8ZGJoHg+RQV3bRZnAl
9/KNl/CSz8Jr1nm+MVGEKN+cKPP6GvL1voc50yOmbOAEDSVX76WDEi5AR1rYBDhX/AP7Ut2DDCxg
edIVEo1/XVEJwV0P3DjgHB9c+33Q7tmNKQTlFbE0VYezinYnAZ+vXQyL2qhNu61GSzILazUxCzlR
/ZGczWWz3vswtJS4s4vLrm0G8S1mEq3SHAcyJCe4BTSAZsyjfBDxRLFognl8IzYZ9xQj0Yik7w7E
T0DPUfAwonzL0C42b+B8fPxxMmkkUmuYINDlyMoPc+PNSZYRiGwzOa7j6A6AE1iY3BX3LeO/UduV
hqz9b2DqpSoRQ9pmmidfxQI6lsI7Zsa9DX17W0HXpg89WAxD8YA0Gorw9uPqpkFCmPBYuEmXAkLh
AFXaItwuQ2e9gYTxURVpmnIU+she4HHo8DKBDtHXGmIrUF/z72nnpK/kB87XJvMnRjhyxirgHnkz
wnOCBfQ+5KAx6cl+bQqggUI3geJW/rGMKVJ4PzuiuCOyjjwPoWPjxzj+iipcVYRvDHbZwG9zvZ9+
jZw+E9NhgevuMHJ/zeyXP2CRj3k69B5DFOw14RosSs2VYJeyaI/QE5KoKzKx44Wv1JtcctxDi//f
2vwZBe89mBH2eEIBIt9Y2+6xh843k9ZB7pT0lMHbybIQKVWVylpK9zfK9Ldly7BksAi7TVStYflO
yyE47aIZBqwKsIaXeQ/Lre/gjV19qqHjhU86++4FknDUy3iCTHMu+W5armwXPQtUz8ggDsdOLX43
GFLs7iu/Tb8O+7Fi7cNj+MzlmcD5EQHTNF7Lx7FBD2IZ6QjLnqnD+1CTlVubv8RwVtcNnv/BbdNZ
uencqr2jloYbmF/4rt2HO3Z6EofdWtotn3fTCpn9exgZj+MO1MZbO12otZt1/BQggUoixWUbWSFM
8WZtLgWKQ92S8bT0ajRPwerBKncN/55raz78++pKWPTMgtmgvWtTVBt3fgUGMrQu9k3ePrAJRAI7
N3dYVfRSy6YK4aYnUrFURkN27hgsg6e8ohhxgfKTH81hl2AxVLVcqZnfi99YSFEzvIdBA8d36IFw
ObA9K6PkxuHfjF1O7CEveiezr2z5iPNw0lKMDUTwrDiOpxUE6EBmLN5Yj8KTo5RZAeuewb8EnaJt
M8gI7ixPO9cCBsB1iJNuujvUusTi/6f4FwF7lfeclEBJH1NKg0a4t2Z+T+4UKjBrsqH6X18NAFgu
IUloF9n9sfVQoutZKM1Vhn3ZCzuXRA6RQuLuzmHMGDAM0d+U3nnr44eXU0qZwoLe9gpvjSAyuciY
4EuayF7ag+9MUR5D7z63NM2X6sbrtVTQJh39ufz5hu8s+oNr8M0cAXlRFkoF+IZCS9R1AeM+KucP
y337PASoUht+RV5ex5a75G2WxiM8hdoEenrhRFEwG2qvKGNlFTZtWH8sUTN4MatQ318n1wCy3cLf
3WxczXt3e30rLCMlLgzs/czQ3zx6369lbpKj6T6ygQ/xMXc/dojmdOD4IuRz05M9Hxfu2h6OxVj5
R3mmX9kD5KMptKx3b3rkbL3AzbjJuDloaqlQXbZYjE0prB4CqxC7uYrMZYuTxyb6RgT64kctIEGi
h7sy1NnLHqya+kmoRto5P9YBOjlLlq8B94sppT9IqAkiMk3byaIW2q0W3eHEWjhmoubrNTV/QWEe
exF/qOFfXc6pTr6Ir5KJU51/yClFLup1dPcIg2BtV2cVGjQpN6D5k9lTuJgXxbEIJBPu2+r8iTLe
8O2GFXVUjND3+B4Huy04SDg2k7+KIniM/ZVsW1dyjLlXujoWsypvpe26PCUcfyExFdPsReoN+BOc
8TAVdHcrds0xQOsgm/1h+N0DDHrP4dnZCpsQYXw+CxczpqAPYtWXoxgpkCRhGS7CeP5kHgoqreg2
YU/gcZdkbBgyoUwBaH7yPOoDax1zbHwsqSbMJqQak1kMkH3XGs7mNJT/Ujhht+GBcm/giFMIbU4A
h9Jc33HOuWeR3woWbBlOfSI5ylR6o3Yo32oU3a4bbN9U60xl3z85TURtVGTpuQ+X/d65rLCMDAUC
iSRA8xE60n8jEeCmZsQiVi/q47FJwHKUCxtyIXoohmPa7rq7JySnQt2xfC7j2iITukEDmZDvVMK4
3NSZN50pKpyRDTOWy3VButcX0MK3jueOtOtE4tFYYbBRjQa9C5tV+GJB1dP3Sw6jwPzrI5gFfkgX
sV8mRru3zt2zpnq7rwmKT8hD1dhLqCVOqTEJF/ZYA90jGw8vtS6vY+QSffCDm5TeDgMINet2WeRT
1nI1qeKtgtZYCkVp+oSV/KS0rFSnK7GL8lYAJN84mHMu9v3FEj56YQFklRn0p4AOWiWfb+daml41
ghsPjnGLDbuK9QkPeDP//nSRZDdO2C1b2jXu9rmIJYAIW/xrVr4+hTb6X5JB4wNvh/VL9JVcQ+bw
FfXg0Xk4jLGg/vfwarMFNffc6AzwTzADMKQNqgr78hLUGF6YPzcqcMC4Y7nyGNLg3mWKEDsFyoC5
YMqCgro8CtUbfGYQBXp8Y4yW8q8W7amVWVLbKiZA8fyqqS/+1MPCGiKP6QGx8Oi18pCpY5wUAFE0
p6gB4NKa7HYrWkRW26ERln9GMNpUcobV58laBXf0hpjdgcLouHpM2Kl7ppqcrCRtd5aRYCl5BHG2
9ZlTryvmgyRSNBkIKsf/UUq72mQDh7P3dn2nZcxOuceoE3xnDCq5L3OSNvoq4SXr0KkNDN2XbI+5
xhzqzi5Nx8wXcQw/0HBbOrY7Tq3k5GFST1kUAxRHnZ3jH3zX6/5Zxz0vMtp2SsD55PAhJYEeb/qk
T5ETxUJekdF0zxdXr4deN595Qn0zqQRv79OfV51gk4VPA8H/pHT16UXhJ3uLJzNB+duI2WngysQW
EPH1cPmw6tqx7hZn2xFSraroU25Gc3gJJ28u0kwXE70/K1n0J9Z4ErFrrDptrwKUApHntnn5XwlP
rXsxSYnbiOrGDVuWjczUS1HOHyyrUT2bZNfAYime/SqSh11vExKiAb/8KlUFINu5HHmCZTa2WkZD
9+nRkQODUV6RMdiUH3yJ/zeF/psYH42y4StGCoplw8A3mBpN5XnIA2r3dr7/lTWhnrzEUvsVUbwK
PCTR+HdKYntTEziMrSJ+gjSRKlXEjEYa+ECXxHN+gja9SkOeDoNozRZdkuBxyMmVaYpGPPMGQb2S
xsWbE0/PfGCUQvuW0uJzTHj92kHgzfulJ17/VTlPvyY+dweNmKhYDUcFxrvmkkFQtib3cAcedx59
GNJvo76WofPmdxiyo/hlxBDLkn1yjMbJdvOfAb+nkL2KHsmnljHHpFIWaCy9Lq7klkLA1UYOCwjb
Kw75RCoNYEqzA2Vv6CrZc4vHAuv/GwCgRTspbndzCNpQHXMAiUetAhmZDuBBGg6uAUBKm2lCMRVg
3AqgaGCx9XebYepNGJbtE/eceHev2nk7Qa7ZhSxldgpXZiiu2KVr/t4E6Brc4ysGJgQVTnreUvEg
MJKRzHD3uSw+/g6wKy24+bt2WSdr9ZQRp07LjmlxSIV6ygnSHAoJeKg9VnmG+VxkBJ2BCNpypOZt
YqlusjwGL/1358ejm4ucDJDRMmB2YA03I3Oe9Q3cbvoblbF3bylN3kutNc7LKBG3D29LCtoD1oaE
xcSajHrmwFWeOqKXw4zrZRlmZSNzsWHuAWGsdI7Unv/LdjK50STjNr0AvPQhA0+H8yFSUL0qBREF
SRjnkxVHKIGbmJn51CQpebpW0gJKJdaR+QDDPrqqVMD1EWwy8FlVlZl08uQ/WQGcixulaz4XA21s
o55jRI1fMVsmbSSxU0P29p1Sh3WMUjjVQ9v+J7MZj1sQRYr1vhdmcGt0OnMt4z24kKqyCUfMYydn
Y04RGtiS9FPrLP4V4Li7AkPaZiI9NQHrMutxx51zUfExSp4IUEhZlv9wmMBOwi3dmQjvvVA9gfQo
1ZvBz8DOPlOqKN8Snu/h8nyPcCCIt2rtBjGc3+1xA6E00XGrwHdnx21i1B4OShT7iN9IRl39h2gD
Boup1MtIl0n2DVUFH1KkcgHbyK7ke3UHEW2cz1z0i5Hyy8gZtgd3gEBfoJT+c7uTFE7I6jJ36DV7
5K9bUMFLanYdGdTEj737o3PLfEe1z7Y5VFWFzCf96bALJYyffWxrRiuVAeYDt66BzLvOAYq3ll9z
6n8NFf8daXrDo9UpurjsUscbHlUCln3rnC042R8Tc2VDR7D81tKV5+pwTwxUgHGmvXFiqbSUuRsv
XUUWkqnic69IN+HK/g+Pi5i50PfboEwqN+M7C0kVHBQjMMeuF/NQ7i3RI3L9DzDL/GfvYA5+gfk0
4Tm5C5gW8OQpjLyZ2Dg7wHCsOzPN1vjAT/RE/TM2zrQzUwYaMD0GvXyOxhFAA/8csofIcyqvftYF
QJyvSM5B4upse9CQ1Pc7zVInrA89KHmZ0Rl3RCojtCrGHNCeJyPlE3DhhHSMni8++T8Up+rpqtvh
W6Uxmd6UeRzDVhQWo+EZZLxJ1s1CAvliKpGYD+bZQRidI6p2qBmc7dLz/8GsmuPuOu+2nElFyvoq
L7qyIMD9MvjIte83iq/qG9Jk0lF3YYcWwmUtcd9LVyDJuEhhYuDSIy2bYRhNlPLvREeA36EX7Nsr
9ZqzVD7MjGXElxwYoTL0jo+Xr6ZKTHbRM58AHc9vibQsryji77cNXONf7Jrba0aqXY7HtQRfv3BW
0AxqZiXx1rRBJS6Yia21Lgd2LlUF3SYMPER/hieXJ3BNsHOk+/034bpI5bECo9z04D8P0r3F9mbU
XV2Dolnvjaqo7DA+zEx6kcJtHEcx8vcWYq6A8r+9eEuIqxbhDEQiLt0ZrRyRch1ZF17tf46o8jMV
X5A2ZmcaGeuSarZ6sgMY+POiCNICvvVmqzxaRx6vgQqzhhtXm4peqTDJ8qmXFUmcrcsceKLTPp/P
/lE0kTQk6UaxQmi+x4tMYov7Jlcm86gNJzWY6eFoZqQQXosPP/tux5vSxLunQnkD394dTKwUUGMd
m9uRRnXCkwyJg6o+6vYLuMfnwuscBQ6AM4oU8JCKSyZsKWWIogWKxEUSSdHOoP/GAMn/Seh2OY2m
WsFQ+HGj3BPbvgrXpn/iMY4raBHLXJsZJZdMWuScVcGPk1zuXrsjMjJhktP52qBMFGlCRZdm3ENS
gsyBfB56Pt+wdK8efjhbBQlROOq5JgpAIl/eTV67YXclDxuQEjHcq1ODzDlb239v1Qk86ug2PSmd
LF/7LmxcEauWcKKx8+/OwlfzrlpIMp1As+JwvbAS2kEcybvP2mQG5yRpTL1N9I7sL4lK2ouujdTz
2GocWF4hE/RFU7NsedLEN105BButrwsgrR2Pc8s87YtAKkcMB7Ui786SFBibfT0OOoBuZ1+SFx3s
BHMlOuG0HUbmvkK40cf8BFrYsDXAaU5Z5EgyLaBy89Uo22xfNecGBEjefTOCuYbWI5c0Uv58RZHK
kQjTsyg/5HT/Di52Hm8brmaGtXEWZWiP0RGcUUm5K4B7VkEG+C8paf+4nMyCkcFy8+ptAquRAYBO
JYQX9iFDZPyISrWf48tR6knO+R3aRk/q5aVSTHMmBPDpQJndRv8vxGJJbdlgJz8cdOEnsiiFV2DQ
Z/CBI605By3jyZA3OrI6b4aF0CfXojTKH41BHUENsDS59kH5agc5rQ3Mt/q24p0nbW1Z9vx9ZQbE
PnJTvm0hN5E0OXTDVA8DhkY/FXPFxlRI0kOqROPKYcdx4WZJ9n9ZCSmd0p4MqV1T4x+zOTE/Yw8v
V2UIcVX3sPUtwB9Lv0W4tc4Oij/gbFkB1PmnYUFdU1VKn8cAq5xF6VVjvDk6JjEQIdNeI9jZrJB4
GMHiiUNbi2JyUWJzBXRu0Rr2J4TyGFLsmQ3KbN+LKF0jYc3xgEfm0b4jEo6Jkfrr8o/TUKCtyYmf
zbOQDjAXYEWlvQToOnxL8ozj0wXPsDvywtgYOP52soZncoTq8SRiXWpvA4NCEkNSN+mmgz3dIjTn
yj1S66mtkAkYPHNPAGtXAYlxKT5DQ0nU5nhSoCVtyUMFPE06TjaHjpBesWwQcxan9NU2w8WQglDs
U0Gjf3RhKDzXwcDMM5KBWu7sZ3Hb2iUCGg/jr7lUQXELryu47OMXROhdZbVnQyUWSCscCjq9Pn4B
/0val6c0Aag5oqgKj12IQmP3D6EXxM6/sKM9iWQ8aIvGC4LfyNxMuegCT8HyTp9sziVhA3rLNCdE
lT3UcpntaDpqpuPMQpYl3ln3YLpawnW83raX8NRUmg21hQClhQEyNUWGV0dRIOQKvfod1z08CZ94
MkEsiDS7FTAwzWrU8YYdq2v92mcjIBtcLjYxdawhyPVMS6oe4WmU708oO+bv5EvWYSrIKmBBFq5K
Ct/docI3AOc2S+QkLq/dE5pSKJ5s4+tzmUWY8wWd6DzafuuwwravcsVdQpx5GL4dXSOARwtaD3US
/q8df1GaLpVQo7WQK8N+pnXXGNyrBHpqSMWR/ygKRGC9xHFLhZ0NLVZVVOSIcsqI0DSglKQgeIRt
ZKr4ALRZgdhUhHLBs5qRVC8nZTOCWhEM3C2YdxZ1r5FHIahUpdzlNvCIg8/d47Wt/j4unP0ZNqZ8
PZ105wdCy24e7vZHBTQygZkAhrbL0s85AOfS3z9fWUDhkeQuhuYPx65MD4GU3nzpkVwVpgAKZsIE
CILrjMwBcgZRN74NaPc7dpkoTT34KxvthHxjoPuOOIXZtSMwDSWJDs/Ma/7iEfFes5ArzxBFeFsD
xcV9EhFCBfvZvz5k9+BDP9tH5XxA/FpVxDg28rmX8BNmDwQ98LCCbG9FwNixTZ8hhAq0FV7aZOlv
m1zj7xYuND7j2oJ4/HwUip8Hgt+CHN6w2Iqu03OVnw7LcUbSKkUxFw4gyhCD3qNxQhyjfzCmyH3y
lwCz2xXyycwPu+VsEA617O/5NfLTpohfRaxLYaxqANRQJvZMEuJ5nQ9moj/3soR4WzglVmZzVwGh
c8yAg5WhQLcpthqu6SHU1Fbt1kbVSzGiImfbf2IOSdTHc2EK/5geZrPxoLZKMqfCOER7ApBMQrYw
UnRsWuSj1wMfCotrCnFVTYxpQNiNY2biio1eDunXNmZi9e7I837xdyc97rXS/PsVKnA2p/D1RKA4
uoyWzESoTqB1xf9Sbg0zQAAFcOXsNKwbr6BYnfHzR4FuRf+PvqZQWjkMSo6zARBylzy8LwJtPc1j
GOQFw3zC+kBByLYM+o5Dk7VSK7iuAN9l2OAtybM5dkQJkak56ggT4cBi73/ZhlkUBB09EjuVBNFn
s/Rhz3O5zZRpS9Kdczbypop1m2EfcnusIey9erA2dLDClYtZLaSwSpT5/e5YkPFmxNlQljPvgHDD
/okYKZZclVyAfh1e48pb2rj1g7gOI/aq8CcXDJQDNXLoSMGy0Qm2UKyav6gO84I1f/FEJSdcPfTI
bi3rpsvY4K+A2diCB/cNjAND354n2HbzBaOdWdmYvaKirWSUJh3/EbNSTtJaCI3qTxmaQymxcZ92
mklfRLQR1MP+Lq8DsbWO+tHI6fh7b+m5C3tYkNXsDNB35p4YxwzHvXkLaqzRBvVDeq2LY5NLIAqr
NsngIcfDDM0bJduqDxhUdc6MNAWC2OGZfMinu8UUhF+BrWuO94Tj5JLw98avhZfoCiZyf51qCxkl
hzSrnZpZPHUgGzz1omesQ7cnijDMqQUsMEujj+0/5QOS2cKGFU9iK+pkrLne4Fn2CZ7ZfZFiz85r
KVepn6ceIrOO1Qh82YIOfFI9vnUYRRGe5j1Q2rOwzFvC9A0sOFW1sylA/1CrHoX56AhBLKxLBVlT
kJ/HgXwxQwATneRWykHwpS3juRC8HI7C38PRr8/bjNVMjLUmIOmTtegy3gGXudvywfnxn3eatMwl
aB01obipWvK0ZtYvK6Ksnr4zdVy/+vwwYx98pF2a/3gwYrYMROfmxUT2kL/diAsZcKOHt6eiwQFj
eIgrl0dqZQab4Sw49Q1tH5PX9R8VvrFQHUatviBwHW6UlqbBoFB8BKpzovgoDJsFj47TpTQ93SLn
vULOE/VnqVyemoTaszrpQ+ZkjiynvUj1rJhNKHSgODDdH10rjjAoAHIkuuTYwc/OXxVbxcouDTlU
TFUCNAY5CFBNy2WMhC5XENlNC/SuKwcMacRZETMzKrch6nIlWdZvvO92RaaQ7VWDmBrELSLrrTBy
HRVUfa+k3z/kSLW9JlRZotIdmBzXiW9t7r1xtRgs2TngkQqJ8mAKnL1srAqFnZA7RxNnYrkfGuik
vrInlcfdxRift0kk35CryRZ8NqmnTojAkQ+9cX9YFi05cWOzfjtb2nMg5ggXz+KiYtr0uZ6dOCdr
iluxLGBxcJrfJLeoAkFWgCcUCTyg3enUQ8+xLI7VYqXRgCdn/qMK6j5ze8Q3DqRasImoYEgWJ6Hm
c+989oxP/aZFdD9dtYLNn8qFGEbFXab8WUx3PjgoDC7nzocWs+H+xlJWMF2pMX5YALp3RO4auE/c
wzsNqu23i+Ii8idmz2g0qS0mJlSeUyNEvCNvli1AFeFQF7TkG0h8Zm3OQDqPBmG2NwrRO7cFQ5Oz
ye7Nr8+SxGciV7DZZzKPRWpyFMjLb4MogFzWhmk/EWek0zn7zmACZc+qBNyVrWfOmoVDgpELTGLZ
g9/0rXHhJsQEOuDro8TyQ/KTylG6EahgALgNZ2657K4dVXHW4Mn4bqgv2zYUhpVskatGzeqE2lQt
l0Op0opgetjFnOoBlyUhgNiOCJAjLTTfq8eYyyZRIJx4PfqdkkSkzlDAS9pwcrUc2ejShKgor4/P
ZUitp1wvAlxihGC0knouOqVM476uU799RwwEI1RsGNdD7X9qav9dv8Oni88jFZ8F8StjHmkFu4Mm
4JEfQ5khvXQXuiLCmr2rIdHRQuQRNrK710f2RlOynLYyaWKARdnw+HqTtlQ6Ho6k6wLJkUWURSMx
B/0o8je9Vg+mCVQCYY863yDJttVPDXxPi0lsgMDhFl3XA2/fKCBLqo8QgAXcUiARGegsnVdUCtSk
lSvnlFDbmIZymdc54Cz1rIBEzZAcUV11yy8G9bXKKIgEA4ZCcAi4BR4wKAF17zIYcEsaa9mEIrbA
SdUpjAiNuTi4tHPZ/lDbP0tSGv6ROWAuHdi1GppZ3fLpihMZPox3YzOZudlekarKDfZdERZWyzOj
BoErXJvjhpMgTdWtqqOISqulyCH3i/LEZEE0c7E5/a3co2LAhzTSaOnuLimhzZos/q8XWesVk2Yo
1sOWAvLZcfUDA/XKDYPa7/xItB4fSkP/HO+olGFj6KPvo+HYehWaZjUw5gfhZg6hZ2I5ITu3zYzj
7STbbmjshx+tOYE4jLdhTfCiZceRpWT9Nnrf9zVoj7WtbLyOLbJ007UjsA75NH1HU+x/lfwB43Hp
5zAtQys+4FcKiy7r6TbC8kHZDwuTUG4SyGkh96W5JMosiDvXb2yI0Sr8VfEoTdeAkWy8/Agm0+VH
2Y6Zzv1IExIqMUBMxW6VfnZ3zhTQXrbr4td3hKkewUL+edaJWqG7czuqMqd184V/OtqiTM/GztTy
hXsSCyFxSL37hKhDhemSHlILMbE4vFYnYsieNulj4GyJVuJmwJEA36xzQ9VkSND9vPpmb0jpwK0P
TdIvIA3mROR6urbAM1+t5MjnDuM1lDjN3LpIiiJ3Bnk5XCK6GCYC+hs1emDhm0C8/E9jWwAm/WHJ
v+mKUxGZacRpkrPjM/k/xKafer0zVHld08jtXe1IZHgvF38ta9TNI8JoLW4To2+MzHAU1BT/3gCd
e6jIVc51IXYmftB6zyo7SwlOpxQ/1teTgHazCUntLa82iwTLmLhCgWuqo6o+BmX22EHJEmda/u5L
cHMqQGAz2l9HY8Glnnk2vMG46KQ/i1WDJhFpce/F6eYXOzY6w7S2s+bkdk3VRbTqAdsqUBSCf94B
0ISzmZNguPhkH7LwowhjvNd0UOYraFPVM1nzlcBY6KIv6r2hMdT4JI2YZg4J5Vk5MH+cMiOc+ies
mq3Sj6InI4/Tu5kBwsJ7tnA5Wi0Hx5KZ551cf5ncpLYB4YI4Kt29hT9ZCNr9fw6BCAWr8ux6PnAr
A3SFV/LCYEKZQKP7OSpSLfbf35qyscc3ukwOLHGT9s7nIqdhp0VDWvtVo9VhFTHpjSTAqzL1EIV6
hkGFpQjdxw8ZorXRvjZY5Z5ZyXHB7V5DvT+LSlEsRajcbuk8qZxNSe6TxjcD9kvLlfCQ1JNBviXu
GtVlpxGzWVzwoxjw2P2P+txsTi2d0F6d36QyX0L5rRtKz2egMTypLx9muXGqXWR3Ft1NPiS/YaVE
aCUD7uZZ5aTOpEirL//RwfRZIyInOyLM2EsP30t09eKA0TpfB3ucSWak/jVvriWV+b0pkXvZLUao
raGpiPvq6p6dGRjPoCbuGXIqmOoa6soHFp94bunBYFWNicUCvBbXnkqswMSnaTbkpOlNYnRwiHAo
LfLkejA2unWkcRTBOZBg9B4m2kwkX4Sqav1YA+dwhw3oXzE+ZLQHylo6K7WOeQL5e0OucTLH4Ru3
/i+VgJYPAqqqb+VYzuWay8avrvXE02VPoN2l0utaffjmNdg4DHLWqx3ZT6Hs/PPww3Qscze9b0kN
ygq3cfWJ/LSwxnhE7g8t1ljDhDdqovRilqFYyzko3bBF1BkHJ6zCOwEut4Uc1ou7YzBRSmGzlmHr
dpGgDdq5B0bpJfXQz3gwB3dTWH+IYfZNg/vXjmyQ2Vlz8Wj4mbZZYw+pxfc+suhnBIjx70ggs6/X
nC3MCIheAZLI5rXFLGK69TinSrd1rMY6cQlkTh3c/pxjPf1hNU+qzbOsNTAY4Y1HckAhXeySlED7
hNJxefXglKwSm1p2IYv4NfhiIc36MLH5Jx8blbwRCdtdeU0Wh0RgN9ytoA8A/4tUEC3oS5CJAuKo
Wf162FywSpCMmewEeRPieHEtqFUOEyh5GENIZ8me5saqDP2rMM9tcmPNxYjDdIjU2472l3TDK8hS
40+vJcvFn5yhnlY1moNoBCVbIvE0rft8XFMGcBaokRiZBxsGW5UUqsF9MnF0mllrNbzD0tKIjl60
QRVejz3guAS3pMpsLfe89CevWr+0A15cZRzVVTROwBky2k+FcTydJUKovlOJn1Nm4L14HjePfJJv
INnt/Ug1Ub6Juf/8IPJKG7/SGQcX/H5OndD7Wa/KKn77MtQMxmwv01T99ZIZNKQRGspwOioYee7E
z615PoTrXBTXzt+9LWFhUFX8R2VpbyGQHykHiXrJ02ngc0mN+dU89X9K5xTqZfxFvKkGj/y2g0p0
Oh8rvkBiorb40PQa+MOWVnRCdYKe7kHeMsyk8tDyAPPZFxZMO+ooMlmThgWdQlcHQKXhRBWNkhQT
jhPGQP3N+exqw8ljzklTwmxGnczXTgY616SUiOmNq6tt3qZRcDybjMj+nYxlU6Znj0Kw+LSjd1Xb
1TazwMgybeZevGmmO12xl8rdVLelxj5PXCN4K3cyc+A51QeJvW/mC8iSCWLxkDJuc8c/e4DI9ycx
Mey+YDdWZtE/77lajd5O1WmDfiNdoWZABGM4NdIlEdi9EgBS+JmnEPTgwUOUMqBANxO3EubVz6g+
f9uCJoZ8xntbN5KlvkikBJg9jdeM0C0CIJ1AJXbwVwpEaZ6SsOeheGzfPD25P9SqoXenNg2LueYB
WluCTzK0zX5dWDoCarqC67IKO0tmHBKc8Jxm8ndMVp7grfUfF/2BauLB5FoTszrDoBfobTdpHFGf
77/7e8nqR3S91AsKRV0PTiElje3moqtuichzeV6FUsgo0Czv6x/spHI8Q8gT5laLRk1OKBrCz90M
mHtoo2QtkmTYoFpOb4oWZ45STGNu7LGV0P4n8yiTeT/xelMNS5IjGytaKIWrjPqfaykAqUqs6OQB
PkF4r6i+Q+XadMVLyE0aStNW8prW3AwyC/WYKLunjdi+ZOhkQ2iB8vPib6FVSnEWtDhuOHqq+OAp
WCzR9BND3iSsFgmU+COebQNc6SMZkBxggZmiWgFMZYxCZ5GqU4b+f7YDuxZLo29DOXfeelWDSMe3
2yjKNdNiLo/7marHsVa95qPjDbNTKBdjD7xLUh4Cf6xbPUKK6lehv9JFTj7Vea/kIUhs1aUwdctJ
0xsPE+5XNt4s61G77s8a2l8CddkVlriMBfF1jmM3jfmXmhFZpYwz/iGgQxWmZdu3sY2ULffE0Uds
S9KsLecnI1S0csWi3rutjJSkmGW8DxOp6DV6eOlarjpPwcdcA5IVPrEiEKg1V5fTrX+IxKzsAM5l
RLC/Xbw0LRGk+Zu7Tp62CoOq7IO05u0hecNCifv8cPulsZeeevxSGOk40n594QVyd76MtJhS2jpR
5ESj0RAQ55LywAwxk0T/P1DDXCLrGDrIeqpxOUubR3YCA6s2NogEcYAT8l74Zj926i2LmiuNbR0x
kA3Sq3mVV8AcMB5TsWpLlYe1aBku6vMlC1xK6OufmArR4I8j35HZ4p+sa1lnI/ylVU2jMDOTIYy7
N1LeuJLWRQQjjgey0NR24eLVw+ayCG2QqrIJjtgzUORlHbDBhVL+hLB39rtcmJ1CMU11LH+4mZ7m
UTR4Z85+sR/UWjnT7joqMUaeBRix3sIcEyKqk9rKIsVJKYHwyMLqK4T8o+lYJcH1MIuJMpEwUJot
WHEgvA1flz8XRbaaBq5qdKFVbj+AjY3Mlu1XTYYOji+hij7aH76SYlmp+TyoBwcoxyLELrg7pzG4
OFnu9qYIoSEvZ4iNMEG9rwjnR5tenNORATJ8Nj9IQKx6+iX0UK+/X97V414J3a3DFZMhANAyAlNs
SkLKe2x2D8+CDaIBrvhde+7uUsMrPNHwENltoZ7KHIWjmZroFtczwlB/WkaBNvjfiwvywPLJhlfc
bc7Wct9D0FZdkte0RZJp03XUmhJatbNlXtpswqEYQUzxgrg5S6wk+nj7UXRo0IPZ1SXGjh4w117s
v4hZDhhAGw9XSW8G7R3bg5taaOPp+iUux5eMTBuVqS1+cdqq0NHXRYh4VnrXS1m5Mj7lS9uG5AuY
QPLjQ1zlLzC8QQdFwLyyKjvfw8OavSkZIi97zqn/+OrdLkWdP86QFoe6OU507xjfRGnteASBZ2EX
+Bv5XGxfLooyb0ImjHPHS6+pET+Hyre9gVfegk+k+XEEk6iWTBkekqWJPcFBdZfT52Uuo6slShbr
irpDB8NKWMAuDUo+qre23U5jChhCEoR0ovOtBIYXMrkDcgxdGMQKMpZu7VoY9Mgll+FThHr+wNFS
mG/yBVKraKavT3oQnresPpNmGy+B+CJ36Cl6qxKtptsveds8Q/8buKM3xmBAVZYfz0aNtZbvYI4n
aFODydCDFXNEbG908dk/LG5EkQrAYHyrGJwFU8Pn5DMUJHl44Qc7e/KJksQToTtKXHFZIbEDlY38
JAfgI8ffKaofywGBt9XAhMH7b1WDjHTODM0HOAWxrWOzy03DIMcQHwC0tYVnUKfc+M0AQGTB68Ze
dN4qgUYwytXfFtQPV/FmCrKYD2YYl+TzANLZOXCsTbduP6T2Ngwb+L2vrgG9FtAqf9tugtl4l1XP
wW0VrCqn2pvgmkapUwwQWhXpQGnch0u1SdcX9GXHoqDtm2WK90uiwFOzEafNwm5hfKSfpIPpnNh4
FtqHyTz3paLn+4ImB5UhQDDgnXutSJ+NVy8i0nLwRRoA4XvGET63e270dG/NLY63QehcBeQ+FIna
fNAZ6PxVMpVE5C9X5EorGAzMeaAhoL1xunxhO3EKmbf6eEsegp+5tG8f3+lueJgDSTXmfvH2OVnt
AIby2wdnLmA6tvCekJQIotp9eBsmIPVyM8XsWwmndW+HPGhau1H6taYKGW2K1ArZN/4YX6gssDPQ
vQslQjGaoEyi/e73Qb7ixsX6VMxY3nkb4Pf+2kqvwjlNfTHShrezwv4RwFKiZ8ruu5fr6262ATZQ
/r5xnv0bymbwcQ51vxBu/w9ejPzzzxGg+iGafJk8YXm0oXbezdgyjB0+imPYvb0ZG+H92950X2mv
Zj9/OxNvOK7mLEPc/DzAKAN+HpJq6NznmbQdFNWGLmn9mQrJi8H/GKa+nDeL7Fcta+wMryfhpVsX
/t8pFjsE60dSVsbMYGpwuT1o2m8TsHkOlLStZxAdVPl2jtpdYLOxoRvnIMRmgFhkp/Gb7emCBF/a
fUTKaZV2Xovb/ns/I2C8EN+dr994a3+c/t/YfCYchyQWYedHrRjSOzR6lS+Is8EZ51lxtnhb6zup
IRMYVhyZzRGlD5DTOHxLQp+WuJm9aToOeKTt81WdNUNLyVrNP7OZGGMfhreEQpHaUfYhCETpoz4R
BRbtld8ek0WbX/POzO7QbAbW9AifNmIQ/jcg2U9WVHy5sshhORHHJilq+OYAyKv7q3+ZLCJxkzGC
xaBjS0dM7dOICA6rpYLLvPaBycP7oOGhEnXwzxLsvjychCmUebN+HFtiHk7YLRpNPqowAcnYXSgL
YPsNiNtEnXMxCL+B0CoIGTofrMGyteoVBJyy7eTYSC6MrKII+W3824baGdhlxzCl2Sd+Nq91XUdO
DkfDKa5yh6tNbnSw2pmNHqtBest7SGZ++MiELYXqRq5nY46eNRt4PSIvw9uJhG7BAHql2ZGxQITa
H0SOA0Hfgw7hY+U2SreKbPD+Lajoo9z3oVE4a4Yj1UBHJRshbOCnXe4iGXvgKl8k2NEOt/Iv1bCf
k+pnnKrS29nhwWqKtIMN1jaITd7kbmXn91kezn5GxlAiRRLObUsh1Fh3g5+mci00MH51MLPd+qkl
mpCn3ypoxNF4kIdZ9gHZ+CYKr+Pp0y9avsvvvp97FsFvF5CxPzd+EeyJYFbp8nbW3eS53DRZdnWf
Ie/Pd0+rATqJxysqFAOITA9SLXRlFaTHg1C6gfaLoqjjcXlWc77MwFXsGWDnAB6BgHOjaLNoM7TO
Lo/9/Nt2fmKUu4ufDE1mXcsasmi91La6JOJbT9ZuP1Y+S2d7QN9mPU0GVGTd9YDJENBrYAVQfAuj
ahws0WV1Ly04/Fks+WdYPdY4nKI71mFP3i0e4umKAji7oxrZMI1mbm2fIGndiUpfA4h9ZJmoURGF
++3U71nsMSFb3GA4SCR370hesCsg5xv/PRl3IfMjgSdQnqKCJ0Ywjuvx5sU1NLORSLvfx4ljrjOX
gRSV9ejfjHP7sV/k9T84peP3jo8N29D7XAQ1ivVnSQMEHY0KeRXiT8jnzsZZe1vFw5tGIPOKPbHJ
tkmtOiM6G0m/CDygEwhxmJ34iQzBktns/cgjoRW7W0/qx2f7NA/zJvB4tbGuOJMUmeXrqTvCVjtz
++oTynyHqfXdhfnFlNN4yAIQAKqgO/3qAQPx/CBMJFdL2lSd3CXtNrcQBUhoOOI+IO600ML5E6dP
1DeyZ0gH8+7AQCoyfm3hTgp98a7fGTw5P/2q0Y7dMZvrPzpCLUtkCNKGK76+arGZuHruwD9j1e4u
wT3gk07pQYmSsIPKmN563C6cpOkxAMUieQ7qidjLVOp0Ha3jsunj3IX4HTAniKMZYOse3fnqqsDy
g3bomE5jecFcZypdL3f15cccoHDI3djnFhpHdqXONwbhDylVA+Amv/KNh9uSxHQ4jvjoFilND//E
kfTsdR6fLDcmWcO32xlLg+W2j0GruiSAMdkYyFoaiKYy+b/ALF5JmMlrxPEwOR8gH5tcffJo1YXM
P6V24/AwZVhp8r2LALC5UttoEdXUGqRAAIHv8FQdjDl9Knm9ZqW+VU4IkmlBir8pst57tIRQbER/
f4VJ5iiAWiy/wdUFLEKSd15+Z6K3aUMG+mswcJH0HInrqR2Q1NZccw0yrGnayf4S6FuvjMRlbl4K
LQuZYDpB+1lxgjJYFCkkQuTk1wTmFQRqx5/v02fc+4JsqV4taZ7nR8bXJLvebtJY8cSh4YKsGeSn
bNYVKEvWb8XQumZmwYlQDwYDXRbcn/osek9qSRYYLSpClgnNNA6OhyQdki676i1DlzH21+Jtkpza
MT1iwxSD2HtYMa9xnE7SkShFUMz8PbZ4Kg9j43/TGiKfzWnwtl1uymJzmeMA1OIH8mpNF3Bzge4M
tkj+RE8r6lI5O8tiu0uhd8Rfu92LwpT5iNRlOL/euz3EBnqkKu9NeCweBKDYeTObSbUmgZG5KvYm
V4gBauyNkm2eiggJkOXys2r+zkGNscBPgeIitXlq4NPfgx4FqYqBlT2aEk1YL/o02fw63EEMOoie
lG/Dyq8moGYFlC1K17Nj/NWOCN2sg/2NU1lt3SaifD9J2NEVnk9yx7nMdQbjE0ArcZXQ8HwZhh2W
rZpZkHP3A4RIyQfi54gHvuRabf5V8zvtmmpJt8XtCDKTiYJUo5ikBcm2tWaoxdJ4tluGoi5uW+Uy
q2KDTjbVq+1FVLzhjI6sQ+6d4puPE2P5I1Ydlk7X441yPaMR7jFM9SK1H+9fHkBhHR4k4JG8zqhj
86mmSCdwlT9p5ENxXmlgkzOS6O34Msik27pM+pfLPuF3IFBVNi5ElnQw6s9xrxrF2FIhV6HfH/nW
6cIMUUlf1lGkYLhrhTaFdaHR+8TvRj1PioDstO+kLlp1YEDTzj84OrTpCKvNsk629dVp6nM+magv
mW+8Bs7xSx9vazxPh6uKE2/fTgnl00tEK5unicHQ1oSqq73YqvKtpM5rIInfT4Rg0YZ8gVpYNLca
Rucf4XIkTXe7wM/ufuNq70+53ZExRpIEUGR61n+aZybyJVNZW0Kq0h9GP5D1iziHQ7C8WHAf+PoG
9/H1NphEzdKhrs5Bdsz/H+VMSy/yZVCNNkIa46BHlnswvEFKh1zCoLVAgBAppJyXkg0DKQAJmCBk
wguWpqp+nRjzsPKgetqX8AoWEFgSXdeh1uLfjHCG9vWGM5xaVnQMW3lBx/JFLzh316SLnAHL1qjn
w4hEEuR8S7fv5+qOyw+xDzVMn+/5oUpksIeS/OiNwd0TPJfgj44+kJavimEoGxlROhP9DmQwiDQv
Gj7wZoubVO0KUrymtSOPA7dkTlf7cJOgIge2Ep1waTwQlIdU89j6wa6Y/0NC3T8oFsztVadXhxXj
JJN26NwtZuYmXf12RXjuW/6slzzV8peFrGX2TMqWBx5hhQk3NlxVkkxgOquoKlxS0Y63vclpbURC
KSfzXI+0Uk5f1NKwjld62Awk4b7xBR0Mxns4zbHPYjRNwIvYSsm/SndaNMY/uqXQgz4oOcrtDCI2
unH6x62rpW51yIvfKTmG6caBXJZVaKg9Xl1YmCM8ofeMacHybztlXjk+k3ebrKm/CmOAX8Qpt8ii
QTROj+X3+3E2SyxpYVggJ6XlY2YpoplKMxtFlpcgCuY89YiRBH3YCEMALDcIOa56i2gg+vcdfCt3
AHhJ9Ffr2uYUsswEnaYaYUPVMuPDk1kXOZS8dJfOp8cn6bzKMN8Sck3PbF1KLGm0MjIg7chkMzH7
CROTLOvc+qd6k6WNpCUNQ4PYsqijHSoHiEXHTeGlGZyySunQ2kkZe6znRjIn1+2qX6NnjsndYiUv
RRZV4Z4rqhohKVUaBGhjKA2y0qBehVpsoVRietJiXB6A1QfOVquoy0c7Lj0+QMRz82B3plDJUdb8
h22nmYu70C2lqk77+skKvw8Y5dkS+YWFau4LiXAFB8/FHUT8F7/iS5NbhEJ6oaEiRlkGF+cZd6T3
YqemyW2MYQFIr7n+qJHq/ikzd9w/P0YOlLkGwhNpldqCMlTFT8X4BM+S8HCcHVE8nb5Z5rLGi/OA
dwSVTHSbKCnxVpC4A7rS0d+Gg3+jPEwt2Z+tPTA4UPbe2xjEbAI5HELdWPJWlg1CfkREj115vcFF
SuHjAnPlA1H0HrDDbs2s7VbJiwwzgsimKeJBT3NUHXyrsoLzhzqjati0W6cHsZ6jjsvXD38ahW+s
+lVG2aIybzfVyE9bd1sbMIEPdJNZk97YVCATWg03O7ZECZbUCh1PJYqU+bUn7kFl+tiTNWQssgtm
bMv01WTfFiLjhn0JS3sfldBme9XfZVJOiQovLTG4S7TfoEWe6UXFm+EWuQZ6koD25m2JH8ADD/zr
QClUfp9/Zu4fIY1g4PfDPvD0lq573pcpyKxXw+hUDPn9lniZLZf47usLImZeV8IN7inck/xxYMYv
22Vu9j6l+cueNr/QtcrA87976fBFlp6PVc53RG8E5kOhfdKS7L8LpV7rujDkVol3LJgB6REpjNgm
W+tULavP2uc3RGTGh3oLlfiJrsd2Cc3d2XjGT588AU4Bbvmq9q48MS9bsLh0hVZj6fzQ/RBDQltp
tnHOs6Y4hctjUxEr12cLOE/9a5WL0OjTiIBkHbNQJPC1b4sQ2B9y9N8409XpeBGAf1xTBzJCouCl
yeiD2hvfia3taG/4gvPto751fcPGI8FYTMB/XedXUsNroWcsBkXJ2fe/Mx3nogUb1aoAL8s5zKDq
WPSz5ERe29FP39tImwF9YbnUeSBuxWnyQXuKzRq8EQrhX/n72xFglIU0kst6PxEVQU8ezVuOMwAC
6lWGbZ6l6jUTvNlmC6lgngsib2AVdMhDquR9+ec25v9mbbQW/gv4ZIAGgzdFSXGqYRROcUk8kQrJ
ayJVMc1Wvc/FSeCSgJ1jc2azhbmzlVpFuxjse07GFaPj377SFMlzTRWFNk2Eo9zoHntgjIkw1Wf/
MBMlGCP2g5XuGA07nWZDsjkHkqfa9plb6eKrlqu0eb5f+M1C8l8Sm+1uYDrO6NaV+N892ZtYmVw+
h+CyjPzg8dacGPeBvd9bmDC/sfcHJMvqRmpygDQ3TNe/6ORUCmVAtJIcy6dkRwK2/hngTBm+soKY
ma4dPCS0kgmWhzFZJ/NZ/Tt+gzyOXCkQUN0/8WFbu8VgnmKd/t7QHLEmUTadJWlMaEnFNokM9Q4B
yHnf0gK2UME+fWv50cto+8AGWwswgck0vffJDORPZrSklSubzTA1Z95rhrCqtsA4Cl0LKj93EUHG
Lv2gjSyOoNOcer+TU2AZaWWhHVzbF4++kqe5pdQsK/Y84WjAWY8vqk+f9lGGym+EgeS87zP4a4DJ
A25xqEAv6oT8tYgQW6juEnyRUL7K+QGhhxsBTdoIugXiHcOZ32jpwSUdmeQ17tH4K0HrVtIRDy4P
5Q/x8bcN+jPN1LbhzHpku+eTmS/if0h6R+RMjSI3euWWxCO6U4/hnqm3EfhTMTqqaa1vIwjwA6bK
AMCaFpBwl3iHQ9Cf3G7dUuyyQidrdUpKS/uQi+Cftuk09Uokcwg1t+XRVKZp7SVK7lxxXFrCL7j0
CfpvJ/rUJV7vzvCZStsVkk7+3FXOKggvxx7zO+rmGhdkAZpsv57FI1l4k2Y1OqH1gEBcYDp6Gz4T
mT0YRyJJH1mt9Eq0EM6bptjaG8RmxdCAEFktFv6N6ynNiNre+7uZj6fYD+LWlLVhXf0PjOiooJQr
ZLufA7TZ076xl0FFcT5yqL8cqiOdztOOSudWNDOQkbw4ngV6X+wecyC1LxRTuCKgpkeWgvgF1NH+
5Ukc5PPdiYmbNs1/lZAenWqijlLJkwBEMiDoJu+f7dkMqiU5ScjlxYaZ4ID5V4W1gsYTOpmQm/jH
P/Y19CKmR4CslzXhYhQ7LpX5fR4Z7T0vxoK9KrT9lFX19P9VnBG1tX0ak68hNGonzzTiLhe2kAFi
NDXx0a2lRb9lrjnYrodpJhYHdURcF7zVAG41ZGFqNgwaj5lkLMjq8oOdEfhFfaKObbjTgNCudVeJ
cssOlny7t+ALn+UPHPDYsOChNHSU4zCPoDGnYgiZTQQ2R8lTEE9FUKesWqOsf9ZyW60YoMfk2zqH
7LtQiCBHijbW/ayNBjr831IS7iI6ORqf2G8hrxRNP9ya5W/ugizWtTEpAM9EUDkQ/oipN5SmpO48
bSPkNGHpjClwPQe1GUIWMbqqnWWHdwYraGrlTw7kUavWW9MCX1ZJNi9xtE+QAxzCcq5qwvPCfSi3
khuivFkv9T9oN05nrFHlVX9bu58W29MkD22CY7Wcxe//ZX0AVKLKTsd+RU8/J2w1VpZRBy+eEVYJ
/jG760/OQ5dkEmNAAUbFZ31aed5sxrSGydchbXNQaiBdSBi0z4u1szatzvbNrroZuvNWTDloyvWB
d4/UMoMj4dU+DMn7mMO8v7H0xOqUSsirihMTNoUcXazQJpKvbshpN8Z013Vz0+7+ilzWYlqYdoDW
JpKocAVuYt04ksclE6jutgO+WPO6FgDJ0ysbHE+7KIyfUznwdctYzuvvrmOfmYnY1EkFphxN4tia
LycDNO5ZFWu6umbXqJrDBE0uxiov6RAj5lIC5b3DvCpip6/2f+v5Y1yXEB+Z72qVz/xwuG2YoK6c
EJBd65OBq6qvR5WGlWHeOmDDOVJOmlVNFFt7gNLuoTdPvIjDZkzuZDmsdTJrf8d0RDuy1Kb4qhqc
Cebl5Eb+BiR8QeuLM/ux9Jz8c7uCXkYidctZn3qqL1Uhlw0eVkrSbykQD9bjJAJ9RuVYdDILnrrv
SCzuzWTsw3/qhRDMRy7+61GvpJqyne0lOdQ55thuP6G3JVlWKG7/24BqnXGgKH7ZmdoAm0aSM2lS
bSDqj84kaFaeTpcVDxCd1firHE360YnazQFxlAZBl9OCG35ivYdR1uJaCHD8593iN1TTettus6cA
KtM8DeApgHF1D8PSeXzZ8XAZolacFgxhMGkeMUx7PRYouSvKS2KLyKn/BUFIEtJ7W6NdVjBSZjhA
TeRo+41bcr7GqteHjh8gy49bJezi5ApXo1oIHMAgsHgHar7Jhj/lfrNums8J93EgnZqigbKsdf55
kYCzZEMijbNJv5fSfrorVzbN4GJWelF9wgPcxamhrbkDpLRzv8SKRdKS8J4xtcUPzDc/56/Eb/r7
iUXZo51Nn5BR7EOuDgWi5/RpacZjW4ITUxOcxggo5xprRoxCnanbIEAOa/+n1+vE3KLAU5WcK1X7
+zUV8/SytB+d8jxJZikcxAYpNq47giV/PuBCuWF/cQb9024bWm8f78hS2cZZjHQdggn37Vm2hM4d
zz8ieJdvdpa68FqDLU8ewZpwApsPfb7AmnSdwLssiTwBtFjstcjm9DGubjZ3dVjxTDJL/NKeUhJN
+zlFt8UNx0/Az4L2WrV6aSW0M8uVsBKncFog5J6Ei+nMFopUzIoLnWExS9BqscJRnFkqZvh8qomZ
KCMS7YxWliyrRu02gCX1L+JGbGG7JYBRFkO6xevjsjnWUxYsNLfCDTiCzg+lJdIr5JiLLUegzlWD
QJqb9WkfL8A/Xyeq0CJ3g5qUMgTOXW94x5Ymk4tlSWm5JtKMztHVRo69MROVtrxyVwzw8Y+aChkN
U2ilEw9CDhwXFEMVKSsUNkCChAL1rs7jL0XKLMeTA37uQOkfQRZD79JD0Mfs0lJpWNbuqiQSUNnt
tCyrexWpgj3VucCR6k/3nFPcR/faW4e6hmsMQHzy4gFo8Bg2hbr3UqAbj8k67r90gCZfDOSz1e5S
rT89+WuR+He1urhbNJnuiIPNofN9z0m2Z2ST/xgR+NKf3gia+qWhKPVH21MtaHPCqCR4fpa5OyEi
kkAaJihSntVCDyNDTUFZ8dgp4YuBQWTR4rut7weiS2qWPtC63a60fSOzXDzIALtSna/8XBu++Qnm
NudNo3Tyv+5CncMV/a3NOaybrn2EXG1z2KrvbBUvTc+uaBEUoZv1JoKLUxzcq8DkmW3gnSZDCTYm
2DhxvylKmKwnx3FbRpZ8yabpwGOmI5X6okgCDxqujhX9+w5AB0l5tfz02vMxwbiXzuoxWiZGTd2Z
SxStfH59I8mHO3lFbEUEQDicg8D58O71dbJX/vMaScAPXN6SMku39OY8PDXvwF1Y5L8EjYLcf1r4
aBpXfJHx63Py90qkBJqp6xAufSyeBUlKYYDdVCylvlSNgt3kZuGtZb4Gtn29IJqUPxqtpg0G7Lf+
l6g1D5XLLnBnXtZETTaTcrnTrBagp+ADeX8SyHicTckzaLDIjupP9JoutHkf3e/g5jFE6GnmeTkL
jbNNG1Rl5I49Gm9U8D8r+a9AIj/Nhc/eXK0aUpBtJ6ZMSt+PFxOl1jLvkgUnU1SQ9m4q7cgbVTwg
6AqceEUc/h+ee4G3H++jknOK+LBjOoWAaA4k6ldzlxfrW7/LjKpbfhtooidCrcUygdoHyyJC8XR/
Pc907WwaAa+aUd/g0b4iWS7giodoYnvuwxKwVybKmUauXQofik0N7tt5zLcJDeJnsnLQCFfXEww3
jOIMa+DHxfPzNrPGHikLTODV5+YEhVQUMxdZpplXZtcK0DRgMGV+m0y9zuwUpLCfDD/cwG1LpH2X
s53t2hu183G7XKeTkInTnRus1mUbajDJHuTw6h5vVY8+8jFWKoEw+YVlrpxjY2PCPWg5Lqq5f5dh
SJgY8TaoLUQ3uggiNVpp7pcCFPjce9M+pFucZG4Xj3Z+sn3i2cvd0ncp1h+aVNEdvLTel9jAg43Y
vEKuFBep2ARk97k6NdjA4eZnm3V+hBhu8hNNX/AYOWVxamP76wDhgRCOoq21qJT4KtQoy3sddpXk
+2uHXVxGQmp8KAcpvxZXwNuecKlabXn8voxT2M92/K3H9/m7blrkwisX9wNJItU7ZdUFtgcWoX6Z
AUa/vVg8ahlBxmaBFkg2wMU7f/sLc2mu6fmB8KFy1lUxkv8bCUHYhtIGOHYCJFjEysgqtH66oCNs
djm919uKRF1aYt9Os7N/XDNVeJldmQ20pyUVR16CItjPhF84zFJPBL930+beAtQnKOO8zTcxFTQB
8POXvSkl7y2kNIYgCeuZcwAjJOLEXAGcX4NHyyuNhugG0mQ4LtVH/yc5ZU6tak7/n1r5YA/LkXMi
SwrokiSJTe9j/w2E7i+mDCIVsOiL96lPJvImKwI5d5N1A3xzMB19KyzSAgZsy9H2YOVnhdR7g/Le
YewF1JOpvOAAkH/DKzEbqFXmF71axSEOuoZAjdhWspJbfJ4utyzVpiFlfSvK/C+NtRVkgVfNY7Fw
BxXb8k9T2dT5FyrsYUEUD5pS3p1XBP5GiC3OYjxebVdicASuvyS05S7YYMhQv0GiMiSyopbJ9HN9
aHFTZGA3r5KZ/ecXCPGqPL3zQ6dnLHYR87svtbc+iEtGa6NShYo9KE9tSSpQjWcH+v74igIOPgr4
297iP3ZGxpDFcy0v56Dm4YPTQOqsN96u4zTO3lVK2MPr49lL5Z1cW5PxUunztYhZbkcng9AxMHO3
GD59POfmUQMCp9JMsWMbZIAMEypz6+kfSWSxqRwoozRR6W8w6c6gj6lxI18bEaq7nA4s04FtQTri
BXlKQ8MAi5TbMeDqwizDy1YDGExlMfnVoDRV4jbGn5DzsBns7HfS3VmM0U+57TMwW0DYePa/e0fh
D7oF2p8uT/1ChAQoDwyFPDgFOJ16v196NB9NVLvMty9EZzS2ZxmkV/RuTcai9v2FIgOA+UV+Kb8v
vpLFLGMAV152pz/GOgGtCIKgt62EaVH1yP5jFI4S7qGHqF7NPVeWis1xpN+dp0Yo2lxs11ctyPEj
mTt+gV2GiNCOLI9ZJvxuQ7OOPpYy/SPgznT7C+Uoq4QOSxYmsn8OIYW98ZIfD+mtt6O4TSXkfWPS
qomRigNMOrII/lE8eZ+OmhCJVVbE4/eZZ/NRU+XEVQMKA8Q/GVpH2/gp/IHrdgX6RBgP0dEHx+l7
SqzI9R4qTRhPQvEtj7kl7rwY0kXKjYrI/Rw6AYJeNVGiX3KvY9FWTD/m6CWL/q9UbMPTlAqFjzUG
NmARS/W72z2JofLoDgE113VMUKAsHe7fTeyAsQ5Ii9d9nfUousHoLKGstpk20AdRNLbdXm1krWlP
uWmF4jNAnY7bkZqxXay0fpQqoNu7eFbMkStyFZCfVFPKlBi3zVgUBesIC4z2Q7X7WgzRW3xXN8/N
lPDlGOCi6hqWYAjRZQeQ4ColCGir+SLdtU2BiMre1ktd7bQ1FeNE32sesUbWTeOSPbpASmAcXTUo
2w7XI/EQEdvM2s4fgb9myKkl/oUnKVfE8LB9GKV+skvfHww+HQ1i8Pk0WzocEKtR8GV2BbIDfcYb
LG96Qa7ysNV+uwBhuyY/uIHZ83m2TQ5OagFxXZnt0/AV8YE4WZR2xpVe/eymgWglcXQfBmt788FZ
7dVOnGzz4nxUOtNcr8buq0XxtyWk0qLx16aDq6NxGNYv+FyxT8kWZqRWC/pSxaWkhhJ7IfQxCL8n
ay8gYKQKnsjnIGA1ZsxHzkmxL+rN55cajSNMqzF3dEwmcx+kHcU0qJG7dnsh+UUDLsYKg3QTWKQG
3DgrZwe01GpK5nRPY+l5nWWdDFi5wECflhLSYTnbCP6Jwbz3i4OgR1Tf5OE2X2ZkBW6jHH/auMxW
cHok9VrRJ+doD9+RFxN6z+NCNyxVGkMX087aeN8oYkiICi4J0EBJdF98BpAVILd/S0Exn36duKyk
BEJ7Dgo8ZHrIT/hFk8rohyxROXzNbqYusfDNMNQ+8Iyp2V5ZvW6ZnvqFyRmr15nyznWxP4DkXWuZ
DVy9E0Mefa1lzDpMpcG3aUAlDJBifoGkE0lA+kfYOzTonG4Ki8UcTT5gN2lwnkpt7GjAyCTnVwME
fIvpYBqHo505qsnqh94beHaCEK/TianQ0R0ePgSOQjjpKl1bbljg6EzDyEFlSBJ5gycds1mzdNu+
pe+pe54/LEUiPFZWl1q97MgBYknAAJ9zmjl6Tv+dFjAYKeqtYVHfIZLRyuWNCXJFcitNMcyUYOM0
N4z3jWISw1gARO+qw49upI3/a5JiCQpf1aXSlbjMMh6tXP+BD7EDdWjFvxGsud8ifCEKzITLRayW
xbgUsGfP5jboiSHvez6mWwW98nWG7dBzEPlkBw57ofZDdlpTY9QT8fq/OeW+33XXP3E78AfSZ1in
1STMBrTFEzlJn2v/oPzNbsmys0ff3PPs2i7srF4Z8V9juvWnxROqfx+gkxZ3BaYB+F9XS6kzdj0U
SQuSPyR0iocu7U+uyZ/MHBM6OOUxNSzZp4cPcBo/XLi3Rl3noQR32aADiX0otugnHXxVRc6FMXBw
fTroHUMGLKNzIjxPwEPFlb+pk2dNS8vaq+Ics3cEBb496Rd7Hf5zoZ44WIPN+veU+5c5zEGClwsf
RJszrHjd52qk9y7LCaD5U84M6JBjoyeA4590frdfIxdTwDn+T9mQchzk5GcgoC9CGRpuk3T4IcQz
on4OGsnPr66M/RX1dOK0RY3HayUYH9EjNPzNJmd7pNvpiA1yj2HFXWhRVffT2y8Ztc5hhNgzjYQj
Ine71F1DBZQ5iGHR76Qf9WRKOHGtxqoFGx6pdRVaZspz29kK49j7dnz3wiGpaJuyqtZTmUimh/5G
DlwAdZIpnOrcTM3KWkiQm0fA2qaEXFGuyqzHpQv6cXpqpYQTeFBlTZaeibR5vSd+VxCvfkqkR8kn
ZaEnh/jVI/U/3bUFLQ5SoqAXOOfKoTcsvvwcASYQ2p68yvwX2db9qZk+DrIp3Rimy6xqdYhX+MxQ
ellcS8iGFPj3Mz2Pe46Txm1I45WZf3wQDuaGw823YmUS3Vi+/FcI+eolqFQmolgRj3JZ481CHhNU
SFOXo39s4svB77ehBLM6PsaP36695dcTXxN8Si6C40jdzMVQL972APm6/7RS+UkvmnF9uwD/NqS4
RPUW8drZ+aTyL4VfvmYF6oK8rmWfqhHr7HDQAWnrt2SQv+dGsXdto4RvB91j+CyiYC9TfjnrPE9/
L+TFPmLJQ631/4UV/Iu9i0O3I4qaq8FKbZCb4SDo7brviBWP8NC+UGZAgIoECsrm+PxK3mSMGTMs
HWbj8t5U4apsXoyueO8jq1+90f6fQZhafsU2oMHmtQ2si1lVhC06HQPsZAziMa1i+WXLBj4q7hav
TCQHwzhpMEMKkRhQXh+j8grtK0EBhMGgebEvQ+IJ9hKyCBymYbTN6pxK4cYxKArk2GpZ5PoZ7xgm
sNObrFx7vSEc9wMCG6RuMJ2vbyQmbMnCUZMobsgWVX+sLDE93r/3PcM58NURa5wpDTboOnRIf9eg
dl7ViNcH0e39Igtmybyri8vS3TxukxYYGolvmJhQl76kST0N3PXCIPImIKCQ2heKMXMHFptzeF15
CKFGQPkvQwGKSa7JX1BaBkZ1ZfmrOSsfd/YF0FeIKRrqr4ZYMN86vp/8cFSuVG2+DKyPsSM922Ya
f90m1UMdHcBdZa/7w+Isn/0kSe+JbpeiMkiwgzSg9JJoANSJ9x5xL6CYwyNbD8XKkJGqh1iN2Hb+
lWA0TXBAmr3eJyy/ELMGL/6tEmvQMxmUIjJELQjeWMwL0IdqcGnwf+ADiLv7OFxih3isVADj1Buk
qValxg7mDFOWheWt7wm3/cv7Sn/xMC0sRlDDZDSIry2ZnI0tZ8Yd74iG3XkZx97m68ObfeyRPSeh
UI6hE7BaQwnpBBv+nuM4DmknGlvpi4vx2q9OTogzQ9g6gvfNBqAphyLkunXiXv5PU2n2df2SuSba
ZnKom/0Gmn1svvc8Vtdc/lOpuFwzhbQ9xcPbsNJGNNBrCTeVIKplnjTJo3AOzEj/B2xTbHJySivF
0OJEE+5NAgqg7pIRxPxcFPmJuq9OCe62fGElh2BlQmEGOC8zO5lhisIgn2pTqRisHTlQhsoGhdM6
34bGHje0HBOcN2Hf119KxxErqQl9mZrNA4oNOtD1LcXdl/iIU8stYucto7hhVgNjEJWoyw7e5h1m
pRSOhZQWK99Ak8z5YHq7O7jXUpqQGjxEeLEGksZwh+frr8L1/RGo8E0VNmpwtmL8Dd/eh8P9Iagi
a/f57Q0CF7ZTyCfENEJJ1JY0PsiSqwfsvoUtjPKry2UcxIt+HXnDVbrEx8AhxpGEax2Z5YaD9Uvg
QoSGlc1X9jkBLBBhXgTIpyek6iXImPg8COW5fIYoj0Bxp/XRWZNnqb663uJLh86T2Adl02tdT5c+
UDS4We1I+o5ySEjZzB0lcgaWLiYgrWvCFwpSPsnR7CNlOpXTUThOJjwos5NXUzDg806IVeDaK8mr
84dMMr0kRR4807Xd7Yqiwcsi59PK6kGLKOkd6Htt543T1wH7QWOkZ9LfnsC6+Ii1l19T9PGuhaI+
2w3LGTCPkUuVQD+eQLwK7yl/ijSSwJQaAAZZFap6RaQLEPq6ySJtSJddfzEcCmikWBNUt4TMTspV
dk6iQo9W0FVSGSg2//dMgWnylabk95QAqK6FHqvBDJ+SDtQF+dZ1KbQQaGdC4vysZ6FlgDhRermk
Qn2yALZMEEIbVdB6KjQrA4Ia4zb/CA/G/jqL0w5c//Yeie/j5235/56KcWV83a62wMqFAA7xFjhB
k/AMmFJ2njToIX8IxrnRJK7SPxADmpkqkSRov89nDHu0cldw0NnutAJRvMS5d91iWFGY5y+Be/AP
037mKWrMCy1yy5uzhsjUufaWOI72N+i95uaK0ZQCSVNIdiCcItVH/X8qWESHrjxhqT9nNq0uywxT
wYseLdG9Q7g/4bIGvm077oWBQFZcTSV1zP7a9zLq8XLyYcUvpUtz/PABGuxBznqYMJzUePC9231N
L50smqIHGbz3EbrrZk8BD6nw4FR04YQb0OxKz5NdDnpcF199HadFrxBs2xxEH8zPo0wE5d7u+lEC
WbYNdlesXGDdtoZsI557v2QhxA+9mkPTXxoljZcWIfkwAQNomv41ybUfUGDvhXWoggEazVoyw3gt
0qUeZQVq2s5otJBlSfrtqWH5FuZH+8qDuRR2Bs4ZpibWky4isjahYZCVbks5eywgwpellXfZ/o2l
EgOW2VNVp609AKKvmZjY4AslX4To2jowVs/0tkUX1EtyXxqWk+dWGscGB3XLTbBcUqm0JmZsHimH
Aq66sgKBVQ7OZkDo6Yp2+3GOquXDhmCLJa9XblVAnlU+V7nn+3YRsZt2hPf1c45PiNRrPrZsKWhe
H+SY1ZcLVgS7ZUp7NjZyT9CbVVKgx8xyx5DHgLiyv0HqO3OiVH2ovM/71aYva8XjZnmlIRhknwc9
xQ75A7MTgz7dDuFo3NwayETyjyE9D8HnL8slw06Oq1tP7vdvh22/oDBuSdbFpicocLMfFiz8Pa9Z
OsEF+MLO1X9j4IxHS9RcTJvXIE04WI/hzGbJkFPGbTDvTIDSqsfiUDLlbzNT+yrg0nWxiCe9jmwt
qua5fU7Bhu8bbsacVh9LHRYY6tj3eZN/2Rp+rozOgrVE/Wfy4AUufs/7wuIEVmgIBvnTUDBCAtE6
GTwtDxerf+9WlDLypVPERS2c/3GvTZhwChJAI97J69tJqegrfxZt4Xbvqmo/U4uuxvbC7FeREDyp
nRwHVF7CMAQWjtQrYqIxs4Q46ds573QAAU/+dG4ZJL/1HwI0+bBNGa8zRNq4DY+wEgMwN0PKMsVq
VWkjUpdh/vuvoO1smtp7IHZNAXnckRGMiXtuLT4iYcL9VTeSVYViXQH51ddBzCbApeT1fnOADjmU
9Bw3bcF0DoAHzd8Ezy8DOFstCbk9EIlvb9pSXKFnKOaDBrTbHi9GSCxp3nvPhXF7adkumjv6UYDi
RLOvvH4wTP/LWCa0C7fclzJ8sG277urywj5PLji0GUrYRQa6Umqjs6ZVkofOmRSJg2a1oqHWJQZa
7Lo3+8Txe8ysnn4hj1M4PgYRlws6iep0P4bwYXFTJvdl6KynkKvbfJ3rXr8tfE7TH/dleifpohyZ
mt7N9zlQeE0ZCpaHyPE/5MCmdqWTrNn860ve4/88tvqnORAcSGQy7syGhLzrXWW97QPOOSN3D23F
zhpJhkeeGnqiZFm55Odisi5R6hf+mx71PewRsgr0zE+E9A6UGNCy/tfihsag9ulQIxg6c7sLpvVz
w0jYI765+BbQePMGgTgqovZ0JmrDNXyOhOBzAQ8mMW15ueZwpBQd8wyYfnYjluwpfhU3OnZRVrIQ
nbzBm8n8UIaRfQ/sBrvR3IFjZpZ1f041zq883/b5R7j0kJ7phZGFA8M1n61gvOwgYLwnunCjqoQQ
Uw4rML4Gpsu+7Kgnpvz31kOw0a/KQ7A+15rN4Z03M2Ao6QPnbE1V8Z5ErveIjTHo32bkgYd4Q3jt
77hm/4dIc9HU09/HoHWMISTcpVt/OcRMSJ1p5t9JPuO/+SakUuKAcauIRdRhWSB+rxxwggezJ7vy
IjGlURSw8xYUXKlo5K1xFFUUtRpJEZJtEwnuvj/mSgrWPfHyuF634CI2ibsJ5U+CssP9x9qT0qT8
qAskG6gSchSAfbsC+2CM1BmIE3yg8QOJcDwC4Mt3Szbi8JhCFl7GZz0oXRpSR8Eo2zq8aGBlhZC0
p1NQ61RW9h2LUmqYq7Zg1qcot3ZHLl+KovAxAUZRYuHvp48qZG0PJoHWhLUSXLP16ErhDU4B+dJY
CRM5X3ES9YBxUr/ICAoFbN5y2F2xwhRjShB4JvC61O1wvhPs0LpGnMk/nDqFGKwsPcUj/tBq9sTp
IKn5khqM/x3vHsm+dm+57eMYCqOh0z1mDPmPRw4I5xBd+nDnQP+s1GXG9qjrhc8p8BH79deHQIOY
YZeMrshKZd6Dj/o0B/7uLvMeo94HcoffQQgmO36aq6A7qx/lS9rHvK5F7gpjCIs3LBQSZ9CV0E95
6tqktAgnygoEz9wQq6zy57otXj/4gasAXQpvQy2t6NqkO37k7ixqq1+y8Y1PyJK2pAkiFcY1lBQn
rJULfjjnSptpupiFvgen0LSXSVCR0eha4w+FA665yYNoJc8KnyLgtpcKktsEKVGlXNmqQr0Sto32
pDVA3u8wUSsd1BU172Lyq+9irJRjZYOoQ0VXDDsuTdo78ISgneMN9CodeY1FZp6gMMZalCrIoGIC
/ZaACL7H94m0s1jfPm6AU44/behFN4xz0B5tFKCaDjf0vJfmZdHTbMVJJiL7f0bUbV4NqzFnrDxq
ooVPB72vGr5HBPk4xjhMv/2lMyqM5kbou6plTF3VGZsUAUt7JXfs+rUgs2qDIipMRotM0YCL8YCT
lcvM1V4ccEiLPvbtxleKr+JmHmsTK3zJif61QPJwaFHJHcYnUrSOXtewoU1XmyPoEXV1vGcVsL4d
KH0vDQB4hC4w4H4+J5mdxlsu8vq5luA1dJ49sqq9hUDGnGRteWJYY/+L8xP2Jvfgk49qRPR6Ly3T
oSUbjBQiSvGVK/BVDCUeZnn6pO2JLG1S62dur/aLE7fTA6mjbLlg5F8Wpej+0izfpen3llkGL6lo
9mclROXA9VYMVElLVy4iCMDLWoiJBzrB7fE6vZWb+ePMZNCjihVRCg+51eqQMbx6lJeVXC4yllIZ
XeMElvBHpaJvNtrS6jQupG5iL0Dnu7v0W+QsKF1hxCt8O/8G7ryp+fHWzvL1DNJidjQ64yWy7bWC
wdotrDaWcrqMgf4gQ8Hny+9qh0eKMxMSi7BDpBqvfRZTfqrEsOdvNWhFXFyqn2viyt0CmN9OTmGV
JFLCaiG48nX7Fs/+jMc/5VfZuGXpZJ4UjUaronJVX0Jv68I/zAlbFD9j1nPmRgufZgPgMu430HOt
7DFkz7ShutG9ULbi6UfqdRZy9A7ZPVSk1SF9ENM1C+HlslRuIExOUwS+/OmyBZQyvmXValTT4+Xs
jD08IEuhVuGu/iRKKXhcDUlxoGObVIABUcfbga1jhifGA9GtIPxxb7ziNnm18zRXuJSBgtRwzKzQ
Epau1/i8+/jWUdsKK+duwxp63GucyKLFHMo5HxkRvzgjiGMTU7wRZzl1eCJyM6Q3DcrAuY8LFa1r
TeuSO8RuwwcUHyr8hi5eEo/dKEVFvr2cmtSn9FHYm+E2D6bdseMB48T0dUJNLaOIEW/yHDc5tFCq
Io5Tw6DqHWAnQJAlzW1q8G4A/EG6mURYX9bhvQi6EF7+festo6ZhbLp/Yg6HbzpBWhAiACZzFIUp
EwpzXsMun9YBGIMs77yQXtljn8ZK6TITnx3Ed5c5iZ+GOThxza3mZIdobyD+BymYoXapgB/gX3KV
yU+SOI1AXeZNhDipMegHEnCm3MrP6PF+rU4l6NMqScM+96PA2W9kmz2gOjGwA247m5gRZz3mZWRP
4lKPgOcEtfJxE/e3ph3XUVn1fQ6SSFmyaO2lXkBLfTSP9YXa9gveK0Dy29D7k0RGra31hlsvwKct
bBKXWBmUPpBRXA3DekvJ93cv3DzyQERsb8XU2PUhFV12z9hfrk2NbZrqWIyPh9vYyRUEIJl4MH2c
ULicJVMe8iqQhUunJ8Qi6omdj1vaM73fXmYeeap3GcQHFPI90o4BXBj+wCG2uaYE1igHQ+1GH8ob
assX7JdjmxNHye/OlvMqMMP81av+kD0Ogl9UqhqpG6CrMM4Myie/8s28LvjiKOjB6d+M4dhMef0d
Z6oUZfIzEjyLC4at9SfU8Dgeg/Ns2JakBkmsqUCV1cYuXhI5VKB4jp+IclXqOJuy7oNj3nIQtdWQ
85AnIzhehBNLaPXb5J/ESr5zKftkwlyb5W8UWhvlsy6KOrtNmKiBy4vayOThQrzZVPyL3buMU7Uc
ht/y5ymaMFuuIPsCbFelc50FwGXwqrrsjM4UGV+b7QfRRFIhl7BMq9CtSqyAsDeHldPz5NwT8c2c
htEHSd2MqeYrP3BDDCdGo5ji0amUX4hGth4K2wQd5gm9I3L1QaHDwcgtpm/wjLcdS0GWN8iySO39
6aS+2/YLkyTMIYwvG15W9lL16u42HnNH73dVfuOCKxVgu49wmbgx3BGa5oEGkVbIUkesKhuIT7Bt
KFip9jjvsZP0+8rye3YmFZSMa2tYBwLHK07IacqJaSpsf7F5eNOSjaBZ2p0Z6BW1Muz8wVaS6oIL
L/aNXGPvWM1sNiuLGyn4PDx0H1aCIK+rkuST6Pbd91RWlSPCOxDqn8Ys4a1/PSMH21qNzsoP3fws
n6npJ0UUZHv80ZhPnzUiK+dRK3oqPdzFQ1GdyFaM0SzUN2CUH5hOEHYAp9EwWNx5aaoXlFLracMk
ZIrbmqhMX4Y8ZxXEd/8JkZIe+SmrBGq9+wG3hl8S6oZpW/LvoSS6GnujjSHoAD7LhqPt7aOm96Sz
V+3opuk0gne+nwrPJR8/U946iHR9Vrjn5X3JfsgumVzBPv1QgIMksO+MLtjWku2Fmm8Sjb2aVOLM
l+tNUVbCT0cmYBePNJVyCtfRPQFl+1Um8fmCsjgYFeS16+orx81Cm6nZoam86WpSGdPlPthswWGN
mWAd48l/tIB/JfCDlPsk+4EiKDo8e7H1WlJfkOeIpkZ7Q3RzVTgfbQZv25Q+UgSVmq4eN3km70VN
hoCDrDhzSVDIoK3lyb8w5RH9UcE/Zl6AewVATfvE89yPEMsuOMs3PaqZ2szGTmF4kaRSoXs3850B
UZPtqAktUpWKiQA/qBhzZJhCTnL0lOu98g83SiBW4/a65M4FLw826oUQ9un4D41VvQRw+hVOQVEZ
XxCu02bqlLgBa6K0s9TBYaaUuILh3IkxBPxothQj/LeXsLLD299KcvhxFLR6CKtwhlpitA24csBX
i64RCk3vgwQwC+iV4Dtg2fySEcnnaiUklj36vi5/OVrq+g2yNJTRLB21oCsxp9HdDPDYKNeaFipe
diXlIXtf9YwSQhb8IFh7fRZDQ6f9ab7hxWzSfsoEb/nGPJopw+HPYPxcHoFfsOWB3mEiM9HnfFvd
FyCAW8YLHsjrOhxTneRzHhoe6mHTUNh7Ai9df3BoGI+uzHz4xQ+lCvqTK6tP1V4csdt49kXcHGPK
Z1dUjwDJRejg15RYT0sLBZLNXKJnWnKb59aOHaozyMhPBJ4uTV92MwVLolEs1lsNVWLsCvV2H2hi
WRtbmSAds/dd221k1q3a9DGdlRMS+DnwIyozAjTrVxmImkJBu3At6ftzcltFGFw8ggyLxOV4poCi
DY2MT61XiBudAeC8zrQDHQo68ZYleDi9Zb/vb5P6RGxV/y7H68OANQcTBepqMspLyzmCnZo3NpSw
D2REkCNYn8e8HSVr2/UoDsadmbUW4QsXF0OtxVbL+k93Sz2kf918VQP8DC2l6p8DS1dcEpqEabjk
dT/RwzLhG0S57YcLnV5DgatG/hSsi5VIWK0/q9uo8eupA8ShaD8NEq119KP0m2dKe6z7i14Yr9rk
HluookWwH22XQ5syNfK0skD1AVNfCLpXLuVoeQA2DPvR5wgR+JqlWhrCIOUK1FWkkIxQ3jgKk3gu
qFDnGbOdIYP/LF+CxBQTRwuQgy/JybAXSfIDPi6UqSuAVN8oDSxwszEg+B2HIpsOmAWot0aYZomh
cZiePfD1yDzTMfTjr7unOK6gaWvgyu1UxT3wcE8WAkhyFRGzoTyOhDHYYk1nj3b3+srokWUUlGSa
n81upgoY+qc+22I390L7jq6KfvoaBzH1/nkxxkD1Xg/gbC/Y7NcBaV36gAx5nq15amnbKMGZkob7
gcjmmwl+xqdrAymqIUv26h1v1TGHQBzX9mrI6ObveKWzBAcr2U8yY0C/YBUyIGv/rQHkRBwN6mr+
CeURZ7L4pJA10EzyeJmxxrDKUTqQQnMF3l0+RtUIMh9/oec1vA37J1IRKfDKzRoMbHM0rQ+1vMo7
/Pokjr5hM6jY0yUsJ5NlsjR2Snve+8PZwuhxWd9lbhz78m2TgnzZ1/oAOEGLVi7r/J/c4F6KwAb5
Bhy+Vls7V/dCehRrgzXMqJnmKpH4UPYI186UajOlcPLeXLnVmJBcwZtmPBT/XEqidR9eBfuXZPVq
0EkqIq9MHgyzHII+5jGc2Fg7h6YvixN+GrvOAkzI6Pt1MBwerlAjeGsMHHIvglO8JazE3RW2NIAX
rGl+6dlk14BHP6EWFnMHyGCMZF0iC5jPHImFW+6TJszsKczjuKi/n/OGdLyXCyqcERYUGRLdNYeC
fmgJOyFagd/8Q/MKHn/3Yn1Mj44xR28N8fyBVfkJYW+PzB+VMfeJMpGZBZqp8+F6CP00s3sE+6/O
WQjRR8Z2862Tdd0JRsdh1sC2s0QS8E6upSYe4mPB5QvHaC1Iv1+BwWKSvjxN8uWYP3kgAnWqYGv6
+bO2nqpUGi/usV5KIGC9yEIonU4u6vZHQuhtbjkOIbD1rWi7D2ysFQYJgm5lIsUq2Jp1+AZka632
aO0ApKD0VkPhArXgsYWsBqeFf4tqCfo+OwBAKBzG3SdY+KO9C/udshWhx9HqU0I6PxlfkI0C1HbT
3r/XgkKSsUwcxziap5ere1eAiNY4sILEpo0NjwhZ2T1IOIoFOK0wN9ZQ/JtDV6fS3z5KDxoIaAqq
NTgUlj1G1ZWbm8nBQc1Vhc9gGKOnuAcKYrBykGfpMr74/i3T5IaCNfcqJzQsXMAaq82YlsY5P1SU
lH9KYMyBqIwVqm38wm6NxLm47IcQociCbXfRRxi8nvWU0yEzRlzTbNE8oD9EoMqO4uetDhYFyPv2
lLdWPsIqHN2MZAPJ1CMojusfk6mA2xo5qkTxIFxxAKp4I24QCmUwU0D1f1ndS8x/+Aa1EGH+DJed
petS2XXZwht5IA5vd6IyyZ8JVUDtPuqJ6X/9kv+sRM7mXRRej1oZhku5n+oIkRGh1c0BGvKVNwQR
/XyYMqdnoTmSNRgLKwJBm2N9sKwqOIDe6HU71e9xpDx7d49yxzaLBEYedojgVzH8gpPETCHJjyrv
bJSgVrffVZSgE3pJrMgtJtiDL8JhpgLKYnMIbkLSN42AXjZxV2vEzRIDNsqV4iLuJOAutLcNRpCp
tEqgnUDGI5iuU8dj/hAuV+Zq/IWuJVyT2ebuJdVH/0RqyYOY7IU11kPUH/HOaOvAsQgiEesa0ftS
kWOE7Djo3PT/gcoZ02/inIFpSTjRlldJBcb7gocSqO4EOjCZTn9PTVMMUeElWJ9vWoNXTqQTWWbN
+tNgCe5iy5OEVRRfjz4uZTehKJcOKdkueFcdTalVvAG3Ee3Z+lF6z72oThHSIbScPqCw1l0cxaNA
/COQfS2aAn87dsFiU1TrFtdZ62qrE0NEvoErRu/ZJLj/27clk1FGO3g7NlqKU+aY55TjLgMSB2TI
taZJr4J/cYyFbDRCeRdD2M+XBnozD+nrcgcHzllLBb2lafqaj4RN3nAFTHZjFozGIl3n2aAPL4G2
QfT9bu7X+xIDpHYsW6FU/AYee8KJ3TYj89xWACJ7o4lw5DlAZDbuTLC3MzCgaIje3qCM8n35JK63
lV54w58FuK7AV/nEaUUWdQYIgKUFNPKoBN6wbHjIdHRkq2/Ko2QWkJwx7EK9Z/6+rDqhZNdVZ24x
RW1KUm4TJ14qWjvYMh4/RRkESWOz4OMo4HSKBNk6FuHP1+T9pYUy9ctpCAPdQCudpUEEsPntjA3a
k015i69yJkBgSiCmQvLWLzdLKk1or2IZmFBwokXulHQHkZcTj7GHWhAn9mSXrvtdKax4GylfHRPZ
YmRpj0znVxALnCjm6aCCqhiSE0HjwXCQ9zdS6FsZvVExhuXoha8hzAPmpePuCu80pWnk4PdqHgjm
QT2uJfWVsx7j5aDq7Arbp30TEmLd/vqfUTCSApdx23tRj4qFM1rVxLXg8nLxHCabWJ8W9K++HRfI
zLTh8LFti+Z21E2QQIEyoOe+EXlu+gO9KKNvI0If//cAsOVgyJsihDmsv3gD7ei+pQjWbOp21a3n
za/ELzsJbRVtjj/BCWdzxSxyKgtI8E4PzL+xu9WQcROuFAn8awLzHt0kYKpGTPCR1V46jmCczVd+
U1DL1yPzVXCVYFe0Snz9H5Fcf6yEtgyXnrgUNA7JSZOgPwQeDnZz2IaFpNYFBlQJQ8F01cTrsO4t
j8KwVySNZoI/1rRUwjPsTfAst0q/ybCer1CqkrWSgE/JxyhSH6UZHQHHviGUs2IyvyxAN81bl1jP
sJz4S+olJYu7tSkHeY1gLulXlOz7R6LMinGPFJ0mITT8sBsFIBJO8LJ1bTS/GAEQDXcPYJ1V0VEf
pop3A825ytibrLJQjno6JrEa8HTg+3eNjK8e3y/+gPmkRdU9vvpQhReeF2ah/Owu3OUaBRNphcFN
WQWKaCtvVatsbUfNsnoEyVd0VM9ch5GFrd4ggmsXHTmi6DHo+qCJgEDjm4F+juzSuLPD4oxVzSSG
Jq3Cbn89btfnxCOPPjFKeyXim+YOwq1uuBuD3Kf7d4OU1lQ2mxfLTdL6gT6FN0Pj0UrWG++N3tIt
2Pg6vWvci8Zi9PXxdaCA1XeSGuf5ZRk0QrXIdw57HRtoRH56pcNEL8KAz3EHOv3MkNnCXqQq4kLg
FKhGNJ58/k36AHsHZYAdwNOEhqKClRHyZvoOFbleKvPJMa+poQEKg5zRz+OW/mUXxk5MlbFVEwGi
j5jcCTVyz02ZSx3aSVeckMbfUmSKPJPoOPxJZHiX87E7l2Zf/XGZCS7KrgCVVG3fbmHFFDXe9L/n
lgaGZb+LegCI6YCjkUoeHSsJ2IUTb/ga8xRorr6AYXjR7Kladsov+GZLxh7yp7pPqgEIsE9b7J9a
MtEhkpHKTsfW9ge0Vfelryv/uwz7R9YdcMgE8VUik0Bwzh69DJwLYCR+bHJvHNcXo6a6IKkAHyqI
18cMbM8V1m+JWbarXP7+9d3UmWmqJJXCnetjHgbHJ5i3GPeFFhB4+Ic04FkBQgNzUsPhpdDPXMcL
F/jCh/3X5WCctFBSAT9JsN5FnKiZ1VPshsnOSFdSPlGfHycOUvfh0f4LnhwOhYAUqJ9RpCX1tZ08
ts8tExJRsWrT/KA8qpvfsBDEw+j1Ew0R25w9FBlgFN+2CQMGVnCrK1OnNj0RY2j6VU3Xe5cs0xla
2Yofi+EKv4jEDvzeUnG7xmLwH1oUo7w0T2hXuzj8f1Q6GpZK5C3VCZrQ3C4Hd6yq6nbSQSN0nO0E
417HT3LkC4vQBUksvjS2tvArCp98I218N3iH+74JU+b7B6TitKNCz5jQE6SZD8mykXr+FchU8p79
QGCGXTc/r7LIrACerd9YePDQSxkGza+oHbg9a1pv8tif1IXe1JT4JThXoFmnpnjXKCHNKy+Tsjge
lYi9zFhd9VCyaU0+rgzC5NsywJJfQYHZw1IYFIwBlfjhOvlgdFzEu9T02Z11BAT/6l3w1lK4znvt
ZPEauoNXyh/j5It70o3GcGfjdh789nL/NQfai5ARjpuX5zlaYFM/OYCCymk+6smvjwfbXRagMhsS
pcr7WWY1lbWd6Pw8UubGaZq/ltc3S22puDrPpsMr9qtvLIUt4qkpSq4YfX4qs+9j7R7gXhdrXncZ
8T/c5JOQjzArPQYR/RUmIvam9na7wp92or+DOIJvk5TEWxvidXip1zeJBmIFFguWhqgtQ5cxSrxm
K0eksq+5khr3ucYcpborfyEPMLXH0n6CHRuwgxfm6oQ6a6HOh7EdAjT9ioAIl3nW+Yhwt9GTrdFx
Mhr1gBN/LlRtjQ7UwG5c21f2na9YwM830GHzKIPK1QA8cjOGlDQsvdjAMXifBe5DkFSd1i3iq1Ct
R8RGvQuosEj+U3QcWKN986dP4VjB7vofB0zmXxE760qNClvTJXrQUSAjTVE2mjMnAnF3VmVv/3Mi
lKglHf6oTbKBNbYg7juWOyr3PLoat8jh0hvJB/1gbq8EHvfjPAFGcgWomyXGXlnDm7v8JL3k5OIl
bgnstj0E68q6lPGmrZyrIEVXU6faIjADdIXc65qxmkKaSwgHsM12P+GhhZ1oL7TeLbQ566H5LAPC
n15RJixu2E6coh8kx/TmZLyBye5oTkcFkQUvpb/OXthUAbbdcNqWYxqPmgt8jHphfCAIE294N3oj
vh8gCipwSRwj0AfEMywwy8F+Nhwane9ZasRW9vYpA38xAIO5fMTU80cuJ28C4RjC3HT6c2Ws0B0w
b9tinvdBxdsleoc8clr1LK/0MmGX6A0IDtXijJa7h7//K+NefejN7NHI0JtEG+Y2oVVRqyuv9/Hw
CPM+f07mwPktBIj5X5oQqA6WhQU+z4964E2YbjTgyiSYY9t3j8MnAkSF4UfggV3qFX5fQ9h2p0dT
juxSBDV6rczc+VWbUSkPYteerZTKcN+7thIrzWur7DID2rCpesWUo8LHwrSyJ6fnx4brEd88FImA
ZRGbQ/W4ISczUdXkNStPqoQ/5rD/Hu+VqzTuX65iNyFn4SS4gUylstkggYbhhLoVVfr9QkDwmNmO
SBW/WwjovMVpymK+As/PMULTu+dLadt2qHiuN2P4bL0vQqh5Va7gBSt3V83BesEigIIzV7iE8JLk
eZ86DeeC/fjCZChYRFY7VLif4DVXwxT9dvLpkLyIaqWtOFQlCfPefzB4LICeVbfH3oZF22fpZVbH
OoP/vF61HFN6LYa+w89mCjq1sPqKbGFY2Hec4EICtWWEUrC7HPnGP5GU7rWbXWmDaytkLlipKcU1
tJx+BaJ8mdLO0qCdeRx0bx4IB72s/st7DzmAVuIFmAV5LIbE3SX44UVrC/I9nR1t2Cqd1RRXVMDS
MNliRhkhbxsTDxY7TLZh/Jdlc8W4wtWCPlZwQ3rkY0+f+kHDObJ626TBfMd/jxP77uOtd6J8kAuX
w1P9tRYDbzvSHBcfY67e8sYxY+QsjPbQQFmR9ENFa9CY2JK5ywr+zZUhaUJy0KntD0fx3fMKKCku
Roq4wCnoq0P0JlDOYiJpRi4sxHn6RCD4Q/vjmTB+/DvcFpVDB9lmypfICQoyt8Nrd/dSkAuHnDee
Ib315s4+QuiLV6V7+BpZp8TSa0aQTuMQGa8Cz7akLcXwwW2S/EPd2GKFNSJcIzxmYyKPRoNeigqx
n/MvX3UzknkQaARJ1TDeZozf/b0VNcz8KdqYwXmyts8GRtiqqwlA//vgSaNjmC0tCQxe6CmAqu5w
dvQcxdNbyFeQK1NFrUuGZ6jVyX6yOZw888qEv9lPQStA4zVZkG6qUgPGoxDZXpPqve2AEXJp+60z
pvOHkcVwm8vC00c62m/mux5i+trr8Vn2W56tZK+aD723sHNbYjmf0nCL6rSBOWNZYfIdufCbO07D
R/FLvUKWhJZqeD0Adx42349usnLh/WhW6cntZDuCbJujoNXnr/qLgPaqT4p1bpP+YXvgd3GOI5wy
2+t7yM065n1go/K9F4Ug7aV8caN4zFTgbGmz8MPJrQOrbUndOWLg6V6UhYVZJwuQnWIQAWmySwip
5z/H8ABYBRTOR1DvSuKfuTMgYNAAqR/CJ6lcCI2E160vxv2RBfgMqkp9bej57Y3ctNvjmYRXL+rw
1aU0fnfg0/rzivwPWNP6aREHxkaB34miglPm5UMyPnmxJDVhpWXYAqINTz6pbQ5J2lP/d8v9Hb9l
aVQzDZjei67Eyd+AS8LzMyMOUCTufyNP3MfyaavmyhVIE1GMbqSJd1H08Kw7mQD/AjohrNwNxLU4
+HJ+sDBkeu5o2AHLUFRgACZBUhJ6V4Vr/xkolp76OY1g3E1KC2gkR/MKNl2r8uVRqbuS9Zsi/Hn9
zzDS47R/SqZEUjZ8VjV5ilZxrccZhEyjXBff378bXqaHQGi4Io0PBsrUcd2qQ6I2k2H6uWlk6sHm
vNi60sJU+hpp99aWmejhg2HZ6/g/sW6HhZOfxWJ+nfblgu7CUV9qCR7srtjiDI3NDxvayGcWP/Yv
9gYTtEosrTCwLeDHlylc9GDYxThmygN1Qvj3sCPP0R8dJpyJEKvCv6SnFUsRh72JTJ8b6FBOJoQ3
vxN3CIrE7kkRLL9hwE6io5vUSZsA30J2la/laH6Et08rG6D4RolZcQUobXbEeE86R+ySqo2NaHC/
96RsSMn4UqBMRrUUV1PjPd1KNl1STIbd14GOuz+8HYKZigAk+JWNmBgSwXnNrOYj9FGxYr9diV+N
nMkRvOiaJsW+VIQA4kUTZXS0SQlWk4a/emZVj8a0ZCZWcYof7C5dIMWDtNzm7Xprfy72NBqabfc9
BrnEf/pSeuMAIiJiplYxhv3lTLN0wd0N/exdPD4MzCMF+90bx9hdvVSo6sl1e/LUmIMfmBMu27J6
UvhPiAJ1wLb0L71FwZvGnKe6kxooqZri49pg9KnxuGBZM4Ii1nt38zGgHGKR/IzxTp8CcHsrG2BW
hug6uWxBVYzQst6FzZvXFFDROIFkO3m+ppZlDNRvop1pzImZtfZD6Ilgf8TuGDffc2btWYryVJ3p
GoTBoomN6wIGI9SdqSNIhszNqY7OgvfUsVSTCq/g5Lj11Eagg6C6Gyjg97bLouIPR2hEMTnWeZAY
ECCgrYyRekCOZJytBONWHP5g5OYNf/3E3rVaspF1oP1AZxRenx/ouk90/V/Zwm3MKxH4jWthmpfd
SlWIJPMWv4PlliAPA/MGJ0j8V+XoustdDfzpisBJGMNDp5fpzdcTkTsXvhK0/yZcsjn9366WEokg
x3piwidD9xYJvzTrgXTaKl29ExTriqXorr5IIFoyUy7Cb7lkqqdqomByWSXgjQtac/qy+YmTxOHo
Td2hUhObPNjqaoJAineVxx5BRMC3VDn3d2MyRcSrveSVgr18DW368GJIJ11Crwr3WeoK8sTjwwJr
rtSh3Udjb14YRhMtFqMmtptCWMofMYWWueiVJcmj6BguM7yKB19cRHj4tCX7J+xkFfJrBB184j1H
GetOerywbt7wZ3WUO01Oy/nX1cMbdfrG7kasqtOWKyQ0LofBGorqr7uYogrV2xbB9m0mrn8O0uYZ
fWYH3uS6vK3KUijNLoeQf/6CK2zHREIJ8kI9jp6TfPjGNfRM2BOsROuZpy8lVQe2Lg8BW8HjTBBH
JR66XfAPiDpTcWY8CiR1I+0joVfF00icKZYQgkiqkCsFNnNBFOpI+fQqzEKnl+xmwlycpyZkPi+D
+fq8zB7Ors9//5Zi2/zq66py32P2HYi//bGqCUbP77xBy1d05keiEBaZhQzCjoEbr5Z9bVR7ZEnS
NwsP2QTyuDV+HthNIjhVjPL4tKQ4gNhJbmqxGQWruc0Gc/fBp58S2ga4DVvheGgRe7mQpwa2dGxy
wg+Pdk7IptyvQ6QVDKAGszm9ivWs0f7EomK8w86Akwl65pn6aWLVeQZmnBd4Te3kcYwJ5aEZmJZZ
3NTkHWcQqQJr93cjJuwq0SCYgV0uoAhPIl+uBtxvfjRyP8OihRmSUMkfWBh7LTHkMkeBqSNxX8gk
bhZV/k3uARr1EnE3x/U1qj1Nm87yQNMcTRCXHSYh/jK3wHChriJvHznPcQZj6BF10MhxOjzrGyeH
8rcyRqS9M6/IR0Wv9ZwqZ3UindiSVtko4QysLUnbI7ci4qAJnqrjDu7xY00FotR/IGycx41i8Bx2
SPpC8IVtptqD/YBOatxy3eNaFgWfDiCnlrFue1qhInIxmIfrab3tLmMAnUY+QbIhpRzO0e9504wS
Ux91zKc3DefWAEhgtKosK3FmTwGb3nbzMA3BBmRrgB/ow9k3dOmxQplRPvNRWKS1kdJ9MGPF9W6e
Kz3HQ/+QRqwJdGiyzjFL5UzLhiT7HB3H3tGqVme/VJWrl/pQJt5XT+glEzVVQ6hj5Om1hpW0z4tk
Oyz6HzN5KwXreulAoNxkJ7dGfttbQrMLpkDJ+8AW7Kkl8NQXYTHc17U+j+gL/3get8pFEV7Qzic7
P84/cWgC0VyHDEwAFUVwViW1Aioa80hHXrEorKQEChAh+Tgn1kk9C9QcAnApNPiz7Sm5+9SBKQr/
EVgUBPjGefx53uE2Ydqaa3iDNGxbC8kjItG0ilqVd7i1mDimerOyz4cibTQasLhgJsfyZF54Zw8D
HmuuX6ctOzOp3YK/jVUD06vIhLnc4VEVdaKUR0Xvm4ceIA1+xyWU3lQGeBNHboX5mGdoJ8kJ3zSm
UwCW7wvbuc4srLUqLVp2cijd5o3psSsbhpjxO6TM009EU8fKnTMehGUs28TUBK5D5KqEaF3IaWQy
UWn4eXErXP+Q7ZS/kT2fsate5fuuSnklmW47/h9CFS3vnAZkv+wk5tw6xIDzXq6N4ND6Y8NAdEEC
tw5iVQVmqDqE8NGu48LlyZ+KJCXdi3UlvG0Z7hlYKsRpFQ92n4IM0tw69q/uXYE2ZIzJ1M6LvTgh
b8h7AJAy/Se/QTrTqlIt8lksosS8wy4rYyVW/lJm81Btpy8JDCxv2Qo2nUSld94uqGIcS5H7M4Ry
cwmEPWl2LpzjuFhqt5nr7xcuktwsW0kN0wJAYK20wTh1K0/OQi9ekdYWXW7JeEqRBfWlEkK0dl6e
QpO+ItVegDOy3HOHJMufwWqVZrpQwAyUp0PIS+Bwf5C5IB/Pv2ymrc019zpI5FWuxI6NBy4kBvZu
gJFzCnv0cZ5oFKTH6cs4aP0we7aE+UYNZ1IW847Qw7RGsAMQTeij0YS0CQCGRcUpALcywuMVbJEC
zrAM9u/1/NofrTEbOJIKGRtyej6tqE52n31GfYC010BSVpyq82x363EqX2gQfTSGR/7KzJuwRiF8
WuZsCUm7mrJlreSKVdi9o5kCC3YvARTaKTXivP9p63nkycRHulqeuosBmjkon6s8TbOpdXl3E65a
jmnsbGkqx21NbSzikurytxArk74Pian7gzIF/PUEAmBO5NdadwowNA2ixW5hnoLJAipN/xEj/pz/
kd0MJGovas0h2VB7rzHeNzTWKnB3xs15MuGKKsxmxSIhhGbE6uBbpXXUTb8/ZIYIHxBQ+BPDRqWH
bSXEHdhXrfc+f1sJ6esFOEEZIsA0v/MapbqX6PlyETWDvH/65ZcLT9PXgCEHBaiLOhi6jClGz1KU
ZZWW6H1KPoxl5+7ASv78hwYzyduCyJRLnDXjO/Ri/MzFBmmRrEpKWyo6ZH3z9OVaaUMXoaK/Cq4s
dbf6P5aEb1BCkb1xaaPNm0LfRrf9UoqHF0IunIoB2lXudHCIGOz+3gBX+PoumiJtxh4lIctRNqUp
+UNGgS20el8+qxeQKg0i8IxdKqYRoLD9EymY1VNe00WP1OyFPtrGcxd5dOYNHEOoGY2wl7wofwMN
fRNHbAcOIj82Z9yAoumMwIkH9eiqvK6g5sh30OimEvdIFRGG12+UD1inxqZ2DNgSq8hobFsEWhVy
cgMdMS5WMoCxXJYVzfF5eWOvBRFUaiUgMmJB8tkVjkvuYMFUlX4ih8w56dW7x5R0Y+WiSRWMSShv
9CBXLe1x+VgRtfgoYJP+veh4RphGhrWlGFB4VWaF/MxQUSn+NpDy80p+aIIqKwzVwXIM3dDCGAHE
0/tPPaxANKii3vCIX1eCBZQ2IEbIzwDfy7xS8qZkcMvlrPzoPbJldMirXGTk5ZwdHIxp7jwzyHkc
AOLTtDX0rkEiyMyJnqrp78irt4OpI6L6R58IKX8nxCW3GESilGNpfPxzlMY+J6VZkEtOq78CQ9Z7
JZ4V1h9SH/9wEOICBPVQJRoMAmY0FkvpkX636m7q6iFG4DJ6kHkBMY+jmItoKExn/yDVb8yDPy9A
XMzl19MQkWe/HsKrV7ojn+bnLwouFkyTzeNytYH2PImHAC0c/NG+eUEjUISy1h6SzZaQe2NiSBoX
thj55R6PFERxY+Xj8HAVBrn6DqBFBTP7+/WUBa4jUWajQ7OlGQYlRaxDjoWiKOf2TagIZwqj95uS
b39bIBjDfP4bGzlJj/3rO6mC6JleR8n5bp03rwV3Z+Tq0jKWsFHcCs5rMPGXdfqific01U3M+AQZ
TqZDgKuRdq8ZTKp0NL60hz4aNoRGTI1Ir8qga2aomJOnAPSTi96rpj8pEOgRiZ2JWowQ7cCC4kXI
V9Zxon9koljjZUwXylcTfgta5hnL7TWqJPKOsDF6c92CFHjowbPNlm/EcBR1Spx1YrVNKcH5HSu4
6FkP9F0pLkOek7V6/Ns9yd5al+JN7NXAUY53kbR8tLlTbbvcE2BUjpAFd3W0eP0an7UFcu0Dfcdm
CaxIyolAsFd042aXKyhPa7DmmX8f2woyNpz+LPFO1vcCg9g2nH+tuHEyJM4Qr397X+AnGl2qwzx7
7lDdf7JfpZKh/LMCovHNg246pFD77Mc9CuE6f9A6+CUBMhVzQwzc4N2eMaTbKup5eHY8vSou5rAZ
ECuW6cHegDRLfI97j+rQOZA19OQsAE2M3YujXnkdQdTZRNP2wOMXrfsFHWApMYamcWjxuIfu4hDb
Ky7EyvUs3y5SG0CvfcpqkePlkNmMX+QFl4Q5VTR6rTIhzYp6YP3M8BvcGBFwiJh43E9kANuhRDw9
HzGj/3n0auSTixMKgmxhP5xvphBMxi33uNki+dv9BiD5kNTTq+ezNL3CMQhKZJ6RyFdX/Np+YPqf
+2bCET46UB8kwFOqtAxPY8gZlVBWAlO29C/inpdBu848upA3DAOZmsU9hUoB5iD8ySn1a/ZolRbz
4YAYcsCqJABipYNCMlKM+OwosRJLpltHPUwIugb4DfWTN3AxBMTP8rrL7N1ueU5h9XpZ2odrwVDK
VZyzMoBhgRC8++uPYqyxC5DocsQK/jmKVxAWFfHzun8z4ij00nOsOzEn+MrT3yaXupC/i14V6qYm
lgYTLvbwIasnaC2pPBXjqYpwTG6hAVIxpZgytSHkHpaqa+g8v8kXYSwmA6g8+aiZXQAn44YEd1jj
GtWGTuAXy1ywM4+IoR5N/Ku/+kD8fOJmZbRsjzdWwxhr5kS/eY/RyVcbux/5X+9JNf6P5ULVXpWP
y7azjqdS/n7xfmTuaZ13Wpe2+wmGVw0Bn8ZefS0Mq8lKRQQM0aWeSWKCzO2EnIWhIY9dZ24KnCR0
eQrkvtOPjxXaxPGoZGvj7mihZB7vj4q8Hs5CBTej9FxtmKeJFSPD+BzNs7BBKh6oCfXNompO5odQ
GR0z5JiZdgZv98VJrIkV51I6NE0z+uF0mUHjJwp4m5bSl1679xppTK7FLqHPXlVmTkzywoGwe0nh
CGTr6FeQawVWh++CQMKEg3hoHeYXvb2ssqHhmbLhJFwuIo/mfx/MODZSaCqz7dkDUEWGMpRcNn0E
z1uFIBIyt8VO7hzAc5zvZOSk6MM19cQn4pASF7NBdrTDUjfvgxecPjmy1bM58A5k3mXCnnq+s31p
FO6l6aYMkUm71vKaUIJAphHkBkllyZVWkrg70TkQsToW9XE6hYxbIXCws7e38wHQRLOnuQLwpvbX
2dtlCeANwTDkVx9qYfWuvWc21uVFYTWE4Y9j0eI6vsPwW842IxJN1dY9xmCjNKQ5qg90PNyO6ytk
W/OLKbRosBS0uErBX7JboIfCW8BUI+hgM5PsdolfyQmg9iq3hKAjMiAD2hy5vzvOUJAJZ5uUOChx
EhrQ7MNxq6PUon9bstZMPRJwPqcxKiFyvDH6g667kkNs7lH6XpWOloms4fi+Kw+Pkkdyq5i/Qr2Q
oKYPpZ5XsM3L/Hlx7fdTp1MPDhRT3hzc/UVONh/rj2CIuLM7hVgZhrPag1GrDtDPE6XeIf4yyWjQ
HVl6MThPKnq2oOrJnkRA2sed4M6MEKs7eMmpTTH4sVbIhPlrs7NLSF3uE8kLzGTzWITIo7dA3hVm
yM10XxycI7TxfB7i3QaGiIkTej/QQ3/M0Mnn4nMEE66pRLTMOe597A+28lqKi1gLWjYBc39Ts45Z
hDvaFsgeAN7hRZhiZsE236o+2W7xZxRqdiPKGOH0WEv3fN0khBKTRopFt/d6YlDevOE3cumPp6OH
nWAGXzrwd0OFkIHV8qScee1DxZ0xPd1ihC8Ziw1F2BkMDQHIvWJTznigIVa/UYPLm8+IwPOa+OrV
ob3B/yCF3KjGL5YbROh1sLEoeB4CFEYdoc4YSmVwousnFFL1sl5eG6hojWYjzvw4SRvRexo8e67t
6jR9vIG2q2G4nWq1TB2xmC9KQVutPsytbFv819z3LBTA1qr2p/c0sj614ltKqoZwB8Tk8JnrBR2c
SYCbOxmB+7ap7ana9eKMPOZ6KMDmcPexjT5sq8klX0weZRDHnrSarZ40jKYptLns9jq6EbHHRlza
P0rgw4WGk+evAT0HgUNvVw75tF4zQRrWQvqewkiW3DUwOM35hTXQB6efErHdDuYl3ELUZzP4s3NM
9cGSukiE56V1cJaCmxQD3S0Ac9gIPMfmmp581u5/UcJ5u4xroQJPqupTjOsD1PoEXreuimecMJS+
UMynMsYKpPdcUXnCxfGdn3cQfUsNpCDSFiNENJd58J8UjTW38S36s6f3a9TYTcxR4aHAHvafE9j4
H5PWCQ2Wxjlen2/GQb5WyfSEZodaTPMzgObkRIXi/qhohwWs6vKmPnlrU9nBi49hWo9Tx2eKdvUL
za4Qkjg9JyWzNvZKy8Eotg3gZcIaAmvNNRp8CEtzJafrsaoSq+BlqEdQUgdDi5qm6iUe9dRpWCJs
m4YKf1KXHOidiA2jU6i0poeg5xS35FKqkRFFwa91yqVzPVd4gk8r4barYyWzoVuygC6gOpxmA4Gc
qgd7dYAwlWNGf58DEp1SQjRbtI/V/VSNupzovASqSjQ/gDw8Hq3+GlGyA7f3QUKqfVSxlJ46nDrx
jhIXd7gpsOs+4bTbl095EJJuXr+6fSbMO6j0VIYQvaB1wwM+msWNoazKU5zmC136v/A+a8mKlgYc
mQEa4F/gJxeO5yh0SvX7Te7gAwP5K3HW33qiHGc4Q5m8gYAy6x2/tEIkatdIXLkbFT6HZc/rFuSO
13nW1gxGWOaYYGfNi3d025mxyawKbB27GPJESWGRGYQSSF9LVhkdFeoSqBcTsSvSc8v2n1+0TL2w
VCKc+xZFPqY2tloGzU440542EPvtSBoFY10fYQW572ceDHQHoq9BosxlT7LiEVtPLHba/uLH7xo0
8au4dNb201VwAZ2H1lfTI2aCGlHQgItX1alwqCzJ5IHfLFzpgQ8GH0YOpdloGnVcy7A72qtiIH5J
mySIH9oQFO+XpWqJoBWS0Bj5mFnAGZHz+bksAcfyHznmA09vv0kNaM2+yvI2TGPnKfAVTeEvrlor
12I4U1qI/soCAoP4SQUh7WdIzTEOBqnpdOpms1vGz/jvzXD32hhAAdKsWqoi+ONgLuOtgoj26+E2
zaHGBYi4YaWyudsFaRWHHaxGYWhucWc0eQSYEvMWB1GT59wWEQKy5I+9rCfnzhJ27G1Y9Bl8gj4c
10N2qLQu5OzAUe76bh05GOzzdPDKX9thPYQa5uavprdeChggzdpCbkwZCrMW7ZAP8eG2oT6X1Z0b
nxqdKx26FNZTHGfXed5mckGIHNa07o+M0VueRbONsEpiMTDYH45KgDFy52f7mEI3IxeVPO0fMVUK
ymlIAU58R8AUUg0pc0MnfeQmomh8mLMDw0ac8Ifpr/wn3a0fgZayqfSgU12RA/kiEfh0aBPYHa89
+AqphgwAggWBFNhP9TFLiBO5DKd1GkmX+GX224wiaDLsvxHWBuPSwK+pOiwE0wsE0IRikOWyzvy1
0trvF18VRFm2+aAn/4EPk9Jj617Jfb/V8MS2NKKZS94EZSX7FQyAv4E/voOp98OWKcIp984uryrM
ZWV03/V4oGYfptg8lhlHhulCsmhlzttO4OvFm5cuHBtEBeEZx7XLGJK4p+0lpmxx4uUAAJvU/GSO
CBGW2Y5UXAp1m+xOUsHVFn3cpD8YvTLjNM194K4wQKp2Hdyb8/AigNm19u4IJ+IARm8WM+hE0GoB
rOHY2A2Aa9W2d/BOMBe6TK/ua+D0YFB/9lTxhdi82t9XKcaGbwmzHEr8x5+/vGG1r3kSxyy9Gcqk
b8HnMFnt2sqH/GS44VVk5u0in+gW8kGsguuj6OuPpZyRM6ki6yihRtgPwAR8KVxqm8gcmPDeI907
PwbfRTw0SNRBJzQDtgJVIwQoyQdd5yi4abKwpKYGPWn5iZtn5IoKlJwCLsuNH0Xjs+Gz2VW9RZzj
uJB5YP+qYdsttLavJbRYCagQui7shw2Gg9YXLSIFR2NtK48UDFA1aLu0pVDZxkvZbJCT7uwOnNsn
Dxvn+9UHXGjfazC7TZ4UfpK32+S9BA+hWrkCLd0QBinXzxM7Qky3zWGVNYouBia7cncmkuaeWaaW
Q5ozMvAj4Q5Q35qfg4elbFB0ejz3PKoUOh7F1auR5G4y/XUrXCxUKa+saAsn193aKasUr5FmIq9A
8t7jcQnUbSqnHRlnMvaKb7KEUkuJ3NohA6gZrIgRN9jLjJ4nh89fWTBJtUP05zVx0yC8JNsMH+G5
DgPIFThPXor5gTBApdjtKnwU6M1sEokuA65+rtNWsh1uIX5yeg3mrZinN1ZIU+yaynZCqRU6+yeD
ITVWUIxQ7U2eh7np2RDQoo99is76AClnLZxbm/kFBXmuDtBtvJ9dsMWltJA1Jlk+ojwfa3/3PKiu
8xDBUB/gcbsmb+Ykexl11myEWZq3UoN8Mb44GPc47a2y4xfLMWbGP+qAeH4GxoOs+Pn2icmAz9Bz
e3T4NjpR2yJZ3Yow2EVQGhmOhNjFdzxlAXe01aFGlx0aAOX5yNnBUAQDc6I/ifEMs1lnCkA1xtyy
hpMlj2mMUlKfGTH2vgf/norLyFwgOVuhQpcn6mdKRdjsdqsAlREUZgXGC2W60d/IOqQ0wXUCRPmf
99EbmSNbI8HF9VTQsVHyrWNDRgWnE825tBUQjILtigY8z0um2w/QWhVCVA/MmsorcLa4DKywwlzI
cUrWa+7ACSioxmMune1kAIoRvzMhya33HFMLEofTOzMzrs5XMPUN/2wn6Fy3t2xyN6qFL2WR08VC
tMwH7B9wkvpAkEg3mMLTgmaeel7TTBgsTnowGP6q3GowUnrXa1KBPsDC+y0cI1ZSVWyroNl+mU0e
y3uWrVgFI8y0ksYqPi2FY+H78IW9sjBpMBownQ8UAmN/nwlpr0Beq39AoEYpDuPrHe7rgRf0aIXu
mXzKRGJFJOCrMTzirrI68VYXt8WsBiR8SaliFXKtNf8QA97zrrpA+85FE7FcT2FOhpMKO9b7xaaF
g3cqztRFL5orqHybOg4Uga/Zq0PfYNsmD0hUzXAyCmqekoTcEj9Kg6a3Jrx3hCaL1UGHLgbVvxXj
FQAbtqmENd5mWtDCbQnDDo8OtzqzZ7lM9Ipw6aIsTtsK61k2xJW82/9TsGzoaDhXLF3PEP1kRsz4
hZZZmW4kP91jJIV9ikRDSY/cjI5mQO4RgNos1wYrokM8K3G1HuL1fetOVFZY7Eyf5rDh3fpnZ1OW
OcHk1nqp0PA6BR6BB9PWy3usFge/PXc6ktLxQNgYqPfVdJg0Ijim4sQZ7BDYUAvUqZKSzpwlZLho
UtDIuY1z4D4OTZbTL4lJI0HwSekMhQ40+n7zgtbBP2IWbqPnpffIJrgBbUTNzfEPPNkt+9jjscwH
11YvpCfVgNYArG+Qzs6sGjV9e+5AcOd8n4E1ZFnhcV4ZXa7QNW4mwXosEP1aAAlawG4z7/Bi63h0
PhADsFPc7Wxn5Oa7smDpxB+yj+cZL+gF26/OczRZ3Ip+r7NkGSAAsb/Ao6xB97vLRFqvx6eWmIC1
g/+xfS8u/clT9veC/Gpm9L3/yif2WYgRyquG9eZ+BvA+yWH4t5IqLCoJwRWoYQZNGtKs/4U7hhCn
2+zDxPz+Xz9O+KxOJf97RgfWYgJUA1vG81alSPjVVQbYMOuYWX6uAP4xD1SqaRMl+9oQvmPlHQwL
mVuC+ARyQQXPisUo+ipkytaQhYoJDX1bJmac+ldkXeFX156tuwbPaUCfeu6hmSvDBEVsxQ0vZtS7
WyRwLsKJRZyms5L3bTtOM0/Nc03P3l8hx97HOfdrd+EZl04JJ02lNCYlala2VkdoRYk3uJwoqj3h
WCE8EcJVmblDYjKzMSu6bhwC/zpVjVdb/vyWAC/rXzbNDE16NiEez/1p4eoEunMO0/Yrd5A2xxQz
QKsaWp39Yloy1YM3LF1T8AkduEPQGPb1Mjf1Alq6713zHHtCEKOcv8bbviumHWpZIHTVGueU/aYb
VDdfyweX6IVsbe0L/DMLE13SKVQPYuWPdOz8TXr65B4eT/NNZLBXX9jyzhkLNERPicHXT703LIBd
lewZQsI6ZSEvXdxm/A9wrRou7Hmxqa8PyDoVT7Mpb2mgNjPos/EJobVGFMtTWjP5wLLtkQHNa6iA
s4f5E/fhE5q3YE/XrpRsTLkobkwne8KKIkM+pjZdErq2yor8+s1eu29Bh+AWQbuXrfpZkG9QhVD/
l9qiH8DuwlSBfynvUyQrCdP1F+pICxQa3/5nKQqLjg0NZVyj5TDnnEfFScZOHExwI9NcsfCacM5S
nBXZbcStH22jQWoFeKyBaPLLTVXR+BWteohgWyt+O/a+AfS1MV2bncd2NM8wZsy06VFzBf6/4qfH
eHNS6Go3q0i7AiuXEX920NaOoVcmLEI+xUWQ9KupPixkwo2f6nEquwjgAWjJSH2Ks0BDgw73hs04
PSbuIMpgn2LjOiL0/6iDCwLHgO2cIXe30lJ+0ZaGorCSwmA+TAI/3j3od+u9FmUDcNC+QQFEO+3r
I+f8gujseqCyUef/WrmhgonEdUCUnX5LbC+e6M1fJ74psZJY42sKvmkMf6XMoU+dkt/IuCyKlPAx
RsVj7glnwY8A9DtghKwjQJ6RIgsk6mwEd96lU47SiXYrp8sYU3CL6sg19gXFs3rz5tuYiLGjqhja
ja6OYA2B5ECvvB1tSjavtP8zBy3g4PQKBKCUxHQ3rIo7elynro5H2XAUyWDdmRnJLTDYUW2uXzhf
zloczkPt2DcrHJPbZ2jVNSYfqn/oquX80aLZranegI3LqxNGYQhWIcHSobUqqAK5D8dzoGFGLgFv
605Z/JPuaNmJTcZ5jJq8qF43CQEqZe8mhjsIqt2BMBpfv9gPXZVrK35tSPVXKVh73BdM3TnWP3jn
9GI0zp5d4Q2CEja/dL6JfVfaXqOpFhIq5Ie2nhorRSLy8lmZv4elWBuoT9pLXnpxfpDiCMHaZLtD
Q3kOrHfoGGJf1Rukc9Im3fskLlP7uTxabUmksUaHZ+FoWOjXeZ8myY//HMhWwYE5IfqsLhQpDHrY
XHiyRWZRrxbeSJG1HrVaw9t9bSRt8VHGJddXmKSz0c/gEcH2n2Ngvny3gRfQeo2r6xsvU+aDt1oX
nWuegaeSKsUzQCeQiZ8lZo8hhjskbVPGDf0x4vPGx17hJ6WH2+hO8P8GiH2fW8b9nDxpc21Oer/u
jdAlhvpA+ZQd/YnS380rolG0od1MWzAdLffNRMbuWrGlxanrdeTGu0Fp0aAIWzlR/P1Q5fdUPW39
MIuOqYm4fyysG8AVonCjaa3LeoH/TJ2RhII9Jg0wB0OCMVkrRBI7fUwJ4GfB065j+NASUfcZGLqI
a/s4nMOu/YMliD+mppNwoy6ebcvbgusFq2wNHt8DBkgFMt9z5BmYdHKMqujCJzaRZyeiVKE8wzZs
q6gSD82xn0WPDrzFa8+ynB4AgT+t8bYHJJxNLoqbS5qBkirYrdiazdWqZ0nmqqbTvsvj3jy1lNEN
GN3am042h+JYxnDzs5FQuIpPFuZxS52+TrYvX0Ltj6uqVjQDxSBb+eFCc30cGW087ByBLQlPG7Ry
08P9LuOGL7j7DpRt7DxKVr21RJQ0K0XLp0wIakO2ag2izs/e1dxbeqoaYvmiXIPnbParZ9DHBioh
8Zlpz5mptY4i2XzM0CrvAIofbNra61md/8CSmUW+RNtd38lyLl1XMobqZyDOSrr2WEFYGlEndvi3
CnVYN2w5WyB8XRO4dr5Q5Q8M6VAT/a791xN0OJXbZzJEYhDQsQlvQhcXfDu5/sGhpZ8dR4qswhaB
+rLcoXCSUNWgtviRICfJ73ymUX+XUzGcocSRR+a5kiKhLW7LSSF3Lix6FljVffwOO7IZ/KNYSl4A
kvmTIeKo/kyUrRbkap7TpKIOZMRqAzbPm2RLk33ioOHGYH7rBKeIaso/3a50gx2pzkgP1hIrA5HZ
lnbG0KM0RqGNhtgfht8co7dpu8w7C8TCsq6QslicfK45z6HQumbdlrJ3xEsxiKNgTIbnrcUhkXLh
FQpECHVNcLB4+7PY3L8OPA3CdMm2QktfP3EijHm93csnUcO/1Y0YKCDu0I/fYI7XCx9jU/pRCcVg
RWe5aZeBLt/irfvoAvxOrpGhuzf6nAk2kO2JyvWEWMWE3bn71S/YGGRGJHMt8Yj0EGJ+ABwakQbR
lIOFRh0l2l9bkr6CcWzSwZcwIoGfl6BWGgT+uyqvEeinl0p6wd6l9UVj/ec6pMsQlwpCrjXZNpYf
w90Cu7/fYK41F9xkj2KUl2S6F8e/QWiqwtzMJaoyWLOwZSfBYvCxhqmkIPJ+uE48A3InZJ4HaJRd
SfoM1alXjCWsyyyJtngnIWrwt5w2KDLq/8nY40PjPk+9Kah9o8uyPaATt2W/uXRJW8zlyPPBNnYX
Z28Qoa1isxSPMddv9FfC9W2S5fRoLti7405M25CvjB/74vhEvXHUS8YxV3pQmMzwqpyzatqOBzUe
KE8U/pkPk/VHx77FNoLIkh8xh4Q2zQPE2jDhNvD6H4LLsKEK+WFC+At0DFgGC9+ATC2TnP0GVecT
GvjdWhUPb4/QH9HauR+pUm+88M26cMNmq1eSouPuqCJmDYd9PEPwcYE3a5j3lb0+lQZbBomj9AWb
yVkE4NAiliHoS4UCN1111XgmHYl5aS9OQ+8fDaldXN9ojuSCYOvUbMunYqOiyDx/8KPYF8RJr+i+
ItIhoOwMi5Herati1vSqBgjv4TT9cl576T8hY2hCjb7Nn99ew2E97he5Lpta6QfRMePbv4FYmDTj
4DpLCk1VGAxxVVkrsoYIhxdNUn3ztdIYNdUTCmll9q3a5mZ1+zzizeGS/RhEu3B3/d89Wu22BGrm
g4Q4SQ/jjYPZzdD9n3rCRJe9/MD2CsB5qaamRhhhyAADWHh1ExCMrMZ0Wa9WbYcpojhwEEx52OGB
TCHku7oSc3DqQgKtcY0Pq+liA4CLpRg2Vle1GaDpguI/mWdu17oDSfUJrVbbeezeYrig5XuitEPZ
iuAUbOkJIoEN2OcnEC40gep2jcUIpHtXqUfEOlvBQ5fWSpRn1xcjcB4vKNhnEiERjBAe6bBBQ3n4
qx9P1lU7JTbgRnH9kIiUyUfRJB5gd7ObUr/+3A7QvKPQKD/LjhRsu6NhFNBgMcXxn6GszYf2KO3u
ISK09RMOqRT+ew2jWXyCAbT3F+X0/vF3pxNYbKMKE3KklENDkhgGl2BNnBVvorW8UnYTTSPFDzsC
ri0VWGgPwHV8ocGWJxsuzwyfXCj1SbW5iR1ziqQMsQ6BHgY1qxBCiI8CTDoHghkjlMP01Oyoyn0/
xIvGt9/fnCudwTcT9QFVl0zIDpoHJ8dtDbkT3zPEVOJ5t1MKCq+4k4At/ea4v6RkRP/rZrixoKfV
ls7SsHW5qH3jg1MTgN0UI9v3Xm4JHT/4hvhj+TkSz6Rbw/tud3celbB3yYv+82qpOChIn/HYwjvW
gXHW6//U/uBXX4MC/3bCBLWljeAbrh2NNBs8UpkO+MPDu8AicUPtW3MkvGydqbzJSHBzAjKNh/qQ
WSuAG7JCGP0GdkJPpSbvdiuUPdu8x8qrV6Nyn+xZgshoN70idvFMQYn/rVVMzHur9HP90fD5xQQk
6/I/5/UO1TA97GdHWbVtv+7Zu4Jz+Qv4hEbL+Cfn8b0lah/DlVBc3Hr7OTZFYvi/YkahLgfxvP64
AntUp/zTP3W/VtXeZmCSGVEoLiISkg8ZJRKQYH67aKuuYlcnhgdniQB+dIHoI8SeFZD6xxxCk0c8
rIZY48pJSTpn1oUlJyv29m6Th2VjjyoSpOD2tCKE2YPk20h+x/pM+hiB7tH4Mg4D1ZxV/b8ajYSt
xnIsNuNKMZIBMKlgilqj7SROphtqVkkSpM9TcoTIJD5/QcOKZK55H7SWkOCuYb4dUA3MXeLkwMMI
S7PfA/MWwis7N/GJKp9IVrxEwZncscRxduZYCLexhhAKfXeBHzb9tuYo4YM3+AlsegkSHLIxNh1J
2GP4FysGQnw6ykIutIuEvFz63NDc2O7vC1HGN5mY9fiO/54lwYfBrAw2daM3z585IxvK7dw0f9Sq
hmSZXUNHXZgQyZctm7v58duYmDjiQYp31w2oZkAfFzvu2x1ICYRMAlRZ5pf8HmuycB+KZUCZlsmW
VLlH4taYPFcARtaa9TirwLWEfr8Gd4KSm+m/LFMRqvVd6n/p3FkSC4LZxtiUzxlvwQL3fYoYXYwx
9hb7GmeV6oqmBA2D2S8I7t0IPL0BEP5uHKAqqlPmbR6KbIwud4IUYaWxTaeuhmNhBsBcmiVyG58s
9B98aENpaAXuyhnhDHYC1HF876oA1hv03bVUxMscTABUt/LM4WYI3VfFA0XWUa6Rqg2rQsj405rB
UnqDtEgXIxzXbEFICwsFZsuUeGdo8W4b4wmIVQMiAbS7BM4+jZWaJhJrL3CSSRlQV8Sb89CcLoEi
QwYj6hA7PvyFyNluV8EcF+qzTmttioNb5ymfna/a+yh3+jrxWPJYU3TZdG1ImeRtykS/u9dyWeO+
jxrb2CoCr1kAqCtLLlbGeA32vWTGYWRyRAjf6M9LNBCYArydtZcqdfzOBrXWauUTZDvmtqdU/yB+
q4PzBoIfHPPPi4XHo2dkjPwuep5l98jZyEMjNCtF+bAl6Hg6cQh7jsevp3QL13b0u1vrnnP8aGdn
QIu4JJXTJbUMxCoUo6j4hQeEZZAIfgC3aNXES7K4dqUz6A4homNFFjrOYbN7mjqTZUWoTp8QLv/H
xQnQkrehBkjNLYl+unAXE1Rqfu192MA5MypELDKTnAJG+max2dY5PYq/2JwD91wDyEJf31imndVC
pzyWZuTqEQAsmtddh76UukbKmiSEcphSHfd82rFwT61NKeZR0NQ3eG5H9PYXDeL1uw3OoceiKp+R
kRLbSQokSlpNnAOQhlaEJ1qPacZeUghz/fuwdkKqPlRwq+lBOa3ztgztHf/yjfv8Fa44V2rli/0Z
r7GS0KE3juPLIM3ELeMAK35friw9nRCZ2kKKd0icdmmNOdOxXFsuvvzGp6VfAEtFE4OX9VMHQkXL
Rg8vURag/sECXmLpsULEhwggu0YeTXVM8RZRHJAIeR2ntjSWG1LB7ZCt5b4kRsDVQVac2eJpMIkF
h5eei4hABZ6tWBAlBvJwjgqLxZEca4j1MT8RdalFP7+wjGuWNWwQh1f+6uMpRkPUo0e37sER35z6
trKpT8+CaeD1LZQ2UVJ693Dr8YlosMuBOze4c1OGAIC5D3JHmR9henuWN2N3DbkdUzwovUw5dvPs
MxO4H60NAvBv0d2E97VrxtN72Do0+qLOLit0GhWE0fpSUQgAGx3ehyca0BxfdU+VXn7JAxpz3mFM
YQz9Au+5WboDIQlLl6H6X80JL/58sVJkyOUjPZdLzxrGxaQ123F2I2VigEeIgSsarjuYO+jjyc9E
G1mTHztlFhmfp+33/CJHPmn4IIuG/LuWd2av2S7x7WMrS/6Yjqf1moSXazVf7fsgexLMNZXdhW/P
z3s9gE5J2ZARGCNO3OeLZpwELZoEiLwSYp05ZRvn+QTrod7m3+ZF9ttBh3JQ4ITs0Fu5SVCnvpPX
/YA4s39xcBUWz+UmXTxej+HmeTzJtACYSBWWg/+aTr71V8niR8c1BCaV95nCvSKIPl9M7ggJ8jO2
HQ8yg63p4KfmqLSuwU/maA7f4tEHEHo2X2jYHK4hQ5bJXXPBqFksOef8KC8R7GcHeR8P9mzKXxST
jBxX88vQAHWwl138qBamxcFH78gwuG0B7Ue/3yNfE4S3RMwx+if7i21Q2OREH0rqc3+u0N17Dg7h
PxuTFWUwuTHVhMRJ0ruAmUSBvQEWMPdOUcXJNZyUyUCtOWdYn42ZAcgWrgpIEvEsJRrsdPNkvXVy
aLmxT6JmAgSzFD71vrFcJ1ct9J0UxgM3LMDVYWlXnL7MN3YpA04OFhZMPAb9+pvEhQyL39R0jUbo
OISPvOQSAYyV7xBJ9MkJ0YF82zDz5g36QR0ZJ7cxbzqg5EfilIQ7crNv6iuiBpNKI46fYY9lyuRd
Q2kN6ThTOo0SPL8wgBRh2O4KVYdfyMfKpiXvLbIFUm1lcjc2LsdDa6yngA5MbQuxRowL4UHpnkJM
q7NMvaeRHcV6Qv+Zyuv8FrieEbVvp7vJUCxQphfbh2j5wbhjIVeOH+4nWV43l+8k5L/RvkN2+F8U
PlpSBSlrVxTRyHLkklnL+27sI4VcCE89DGu20JG8h4FZkDLu4dOQH5d+O/VSSpflQkwxpv0T8MGw
Wn9NqQpC8xUsp2VNEKwxzAA6UMr0t6/fB/qgjA9QbkTBNLV5wVoBtZVa7Zaw3ykuOfEf0IZBU+zx
jvV+7v4N33R8LALm0tTKJTgByq3ZEV2d0YK0uUtqqu374Je8oGjesF7+W0/JMBCzGrKNhc/UqWPd
sRU8T18H7X7JeeTUO3AE45z4/xeKIwAkbCyEUqexuZszeJti2JlmDnrpNcuBmJ/35Vo1MB6BGxWk
mhmgW3WaxnmBp4/wHMhfzkn8gfviMPmKhVfl/tUF0pJXGeqm7TKC2ojlvXTBXW42o+HIvjpiF2Fx
Q/uKx+rBwAUr0kujB/j55o19n+MtmlcuEohBQaRF93Pm0Dm1cFefWczbzdpKZZpn22T6MzrI8mcU
SsdAV7qY537df3OOTCa8LNnS69C8VjMGJN2nBEuZtfgw/cdqHS8PzMB9AMMqgNruz9cQDhKNZAqV
BHTiSZeada2TfFhHX2RvIx/Fs/IsAPzmAmApgsF3Bc+0Dtn4rZO92SR7X2MrCs8KWLX1AlgFIOTW
XAaGLJvo5HKCvMnu9UZNtIPEEddjIFcmOzGiFuPxldkjGBVelyDn/DZXB4r3TfI/ZtcRnHahy9v9
VX4iDcK4qb71/cHy8xPkYL0fVq6LIAxX2f8ONQz+MrKcQo3G4UUuVmN0H7GYECyhsnV/r0r+Gxxj
XSDE5n2pNUiUxgGXj5SNpp2uTHHjLGImFmiQBGXnaPmH7OBXSqsQMfJ+8H0vt9jt3B3YA9YP+BXE
uarXGxIyN+YiSKuWAJKc/rYfX5q6Qp1XgLbt3ey92HUPqzD0bBhKRuANVi+6W6+VLMJ1SLGW+qbg
7lPRJcowQpyxz/WovERlSxqQX5aWxagk81nENjC64Rzp+8mcXsttlOFSUKyo6kyPn/WrmMidFuzu
SC/PYc3nVMqr9dD5g/eIc2FogfYrwr6gocDlk7rZTFvmw92+d1pAnciNOp08mEnyYh5Nn9pDciuL
4BIEC5lKbdA7FDTEQpl82YaRaevAkLgih/h46K+J0ogUmaJp39/3zZmu7CfflaJ67/syaIR6sbvJ
uW6ouF9GnMhQYiWmll0hJT4TncD4E9pH6gIo9WeBI46OTZZHBXjp5ilhlAHNX0c6wYVdz594L6Ja
tR4we+Z1ap1kAg43vKd/1FVaSb3kNgjkmEbE6/lkjj5INpe/no7dN7btisyCa5tsSGLxZSDkySm9
633lRxsaW8FnHcI5MS44+UNRhSl28AUJkCRvIJYZPWjFfobQ+pk7730zevSEBG3srgdoHr5fbB87
wQjNbOI1QHZWmFlXwVviEf65h21GjXwn2uD9Mxn4lLQiz43i7NmoFTAgMNKZumClO+Uvh9R9GdaZ
ZFusTKbImRjxZiM2SZnl6lP6nKcFOtv8c1OYgskCr+nA0PjXMhGDNtEWST+j+b+/6jCdAAdbuVPi
JeP4ZxYZwQ10pmzX9iAsbH/J5x0Snw/dAkmXdhWAmoHzQWEa7BOAolXUp9+mtiOc4QklpjxIfgZG
eEvkDtyjQP2jBQOBNTsZP2HGB9+jpIQqab9hmaKo6aL82otZLJfzExpFjjlPtZ/HAP7QmLaReBUJ
te2FZ/vfggxszm9VPlJkeFJQtbXF2uydtiv59vlArXMe5woOrLOac5LeIy0TT9XOTqXqvPf7EgIA
VI73rARJueFbi7hzWnRMzLyx31RR7o3acTaETF2ShihRKCcIGqCFfm7Rh2rPPXpFmpoJJJvb1hBv
DhdFWIqUEgqZoZFy7ZRt8LXggjC6kdSgqeI0029SIsvYC3wxXMyWfJ7x86IF9cUWHeAtZ7OPYfir
bjvn+2LpEyDJamkyOCD5SjjFvFZ0yM5hDReprZpDRYsLroKFvWydGeslxdPgjjlTbNQr7JewwqoT
E0ppLaktZq/EkjQ5sy/fdQgIHXRluEQiGOyxYrRiwcLjd4GuvaJAyqGRtr772hvq19WGSvNvigxg
WPNIw6JMxA9AqkF7jDDxU3T2fkAqs77rpN9MtzfgWR1+B+UwZU5qxDdqSn/dThqj40nWtFMgN/5O
VxrXx+XH/Ot/W0mjcjlHK5I7jUYutxf6d1eyx0d6mYHlIvfkvDyhexA9LoOYJZ0hxa6GxnmUd27I
orPDDP69LbXfJj5Q2jjPsfORrY1qzRRysBVC4wzkSNDqxmkQi1BXN3N1V3VzVJbAuPWnmFMdnBQV
ZAyBZGQQeFmjaj1o6C/ukdSBhK1RmimejmI7FeXLLAIAJsYl9saeOHWvGsVCHX5MGKR+HZ2X06mo
VqEYlWK3UpT0h4mwEKacLcPKqR26dKLhQx0+f9JTQL970B7NAYxdfgOwIb4KWGNsxZbXUeNhnQNq
Vt9lU1eYJwqHIsdpv+QzK30G+hA7+EQ6GpRA5UVIUPw8iDBNhGttTgGgSJH45fnV9haA9Lfu9qy8
gJ3XdGmCzu0mVU2v1iGNLrv3dSXog+g5FmS/PCsXO/Qlcm25nEZUBpydvWu6i6z0mUtIoq167ggo
E0nnmDCq61qYz+oGT7Qf6z4nmpDeosXzgVX21+ZsyCM7HARFKfBE8sQ8rxIXeK35+NxhBmQEj9FV
hw/N5kFhYYj1vTDS0SpfuM3UFfoC6idIgGmqo6GYIrOGrk7Cq3LlFXmvHgh0pU1MWnVefwjBgGu8
JCGhNpEqqmW/iZIjdbjBjGoJqeu1JGhkBTVe1JlKVCT2H4+AgmkhOGwwTxYrgHCirzIGtjRo8O0g
c3xebG3xIU8EYtBuDKy/mCpOdkauJhWFXJ6Kg/q0ju7tUlR1a8ocq/v0keyWfW4ddfs2G25kjySQ
nZhevVcbteKumJ6U3QHpLHbQw6lfExyy195NsydgSmO6v8f+Za9sW8J+R24dLCUXgn+dwHEezXSj
ExILgfjq96tPwvC0P+AQHT9uM7F+s3XeT2QRwBoY/XO3uF7ac5PYzi9r/3t0AtEKRDHUZnYPid4j
CozKZLA/CCRbxVVo1lOcgB+HuWcOTX+u5dw8zWwVAOTfIcRFBXKV4j43NongDi6oXnFs2W6QeVS6
1Y+9UMaSBVkBu+gJbHFUXSq4Sh/WX2nrp6U6M9x6wYrZV1UmWF9tQITx/VVatb6amQM724ajm6Jv
qDiMhLxRhTZ8P46cGlJqxs6B9HQoIgkHCPsL+Dz7U+NDhHvDWwT+lEEX+9i3SKL2/21vG02w0rac
lFW15047AqsY+zGpCsr1MbbfBpt958/6o1UcXwlwkYBd92VGKjP7W9Mxl3KIYnTIL0uJNOUR93vL
qU9B9idBE2+xC0bPLPkly4UN32BwwRb9nPs2d//YlUkZkVbj9Znz6+f6lGJyMw/wzcZ15uWwtumy
uMPmiR2Xxt2S7jtbbD6HtXHiIa9sOQQQId5SH8I609lO40YtD07OgapyMIMkIt+YAxfG19bKMjco
aG8X2Rl/o/rlQL2cklBLNrC5bY9dL83CxypmEphYX2A4I32G+3FA38JvsADLmVUR4pc9Xj+o5kYn
vdxvfb7oubJ03uHnSwR5yBaJrkWeNlGuW0+Yyy5qFtkfI95ZwWecegcY20myxE8Y9f7X3JL8sejb
Wxm/MR1Rz/vyxKYjvXRREHWhHlRy/cIq5RIkHmdR9TBUJEOJJDvgQgqv4ElKbX91m2PXFz2d7CzU
p8hYB8YymZOHnuBP6bMJOPkEhG9bi7TlqS5xPtUebyH60PF+EmtSFeshP6ZGnSgRTxr7A7WqFLZG
afQ90NQA+yjblivKgTQ7xdomk+4+ToGH4+kn/PlXQnzaNVbm4cc64dbvCmJn8YowZ9NGONvn5DqO
BVrmuUfGieACdlT4JQ2qiGlwcZuGUW1kH/lrjz6DzDO582ZS2pO/PJp9LxzZbDvX66WwpuOd3ls7
HA7E8xJuAwoNAUsFOw5ZjYZMkalaFTlQd6CvsbTht3NG5GPlB1fYDODoNlfivJ5pM8SOkh8apbBW
S2nFXto+WX3RTlBzvB9O5XAaTNbsZPm2RK1dpji3B7hJBVtyskl7AEeNfk5X3I6qpB4EHJzQzPzy
H4RcaV+WsLy5AjGzAjKSnoQ+AT7NjrI6AguxpNCSfaShfvbrcA7M+LdgJ33JY8MB49/UmSmGa7Ee
KLbxRxyUtbbQVjueYr5FCQ+SXx6rzCofG9uIf5CvoWi7mQ4Sc7U+5A8o/KcNRMawqjTHxeR3scGg
oXFHkmKgdGyKU6Pd2bOgjcwDKBmk4UgFcABqBe9QoAdxIvOlVBJlZIOEiZSpCMY78GxXMb0e6JMG
5LB0nsnD6yhOFDGpi5oMNqyPPlf+hyuI0JWbnZny2wRzxPd3MfIIl25kcDLPZon874+3dT1fvAIR
VFXuALCTGdaCzB2QDClsHG0Cqbhm8O2he1024f3dLwl55SwpscK5YGYx9+46jGdAczDecqLvc/5v
tv6yGXuEAhPw352g3nQswJMS2I/ombkGHx1Z0H7zQhBw6lzAhMJKIGi6cFp9NhBSC9yYefwl9IuR
Cy25Mn17FAjlCuZQ9YF/GpEHgLW6b8rGqxOV8lGdl1qPXqC9uDw04hNhCpJjMS6bieWFa3xtmt6L
B54pBzETwOzM1ftpQGFtx/n8mxN9Qoml25b8K6ZUKOnHzv0HbnRJ1/SWIz+ewB2N9yNwIWtHKkKl
kLthh7Y4jCYnkPyIiwuobQiNRnP78mPWuMWKaLe41/5Kv5JiiKhqXxiLAyCKuEoSRJSmtLjkM0K6
eTIrYkCvSDWOSKrODR3b8QyLs0X6ae3lcMNkiJu1MSrvQZSID9NDZiop8gUTdAFZC8GtawQlSvM/
ddSHIU5WjNYuLj7TIzpEYQ26WGxvde/2akBgKheauJPMBQLjErjWBpuHPzeM37fdhZ+bHDDreQGY
I58h2gAV4HiXX+H5K3doQGm5KyxburcOGLYmzJ/o+rbrfCH/u9+sE+yjzWyhZBB/Ex6NNdUIO9qE
qEu1wr0VYGVMOg9Vg96fBNSlm1+y+Cf1DKVFSpTGk/R6mCS8GFaGIVTR0VefsBnFR3PrnbyoNhG1
4unShErhPWtaPZ7KKHeUpvNXqwB76bprGSfgZB7gEqtdHsJYMXqa9kqhCPy2Lul947aPg6PQ7GM4
z/c5CwhJpuXlQO8mHz3YV9Ei7rhSsY1SAyMqmgKnUd+F+EWVExdmYxHZkys1nBI4pZNF8hvXByaF
NkaQMXvVGT2O7XGdDzeNAqRFnb1MEDOsrxob4ezMJbDJcRJx+MAxKMy/xuurxQfWTmepq3K3JiBQ
kvqu9UxZ6XwnEhz4uiGkcrC3nwEMWzpEKYlRxHu6s3OSv7fuoQ6718QtNqPei3VN671UNAZ6bUEV
e/2e9zaX8mpK8Op5yy0M0qf4gGrBS8yMvbIFXsv41QBiUu8c0cO66C03md3Pn+/BygwjHGTnIel0
I42OaXzqMrnonQPTRbSgtlHHr12XPUgVShzq/rRqf+bapmp3nuRXvIN6nTDjgeXAezCbEU7vFlE+
ColrKZeklJC/S/zE0ig2f18GE0ikFoV1cBJZbKT255bRJLlTjvyYPhncmG5G4yCKpJDgRPnJka2A
6MUCX+ZMv6qcwbkRPjmUInpeGSTki4qLvHfrM5JDEudlYArl5mchjJuyY/j0a4H0DbO/FZh7uXY+
K3iEBOFHblSrPqqughgh/I4h5x0KQtpFB3wa4ZT28knKDdIwOJpsivQl/BQGwExvByabZxYg0zJm
sNJzQtpbqEIcICu3ls73qOB414kYAIJv/zBv8YROLyoOiJi57r/PHiEgclMRSPGXLILqcqKCCthI
rb4OTMU7VvGRoxWcWUC3gdkffwrMhwoS1TJLflAACc2xC2rZBEzTwCYZErv3TlLwUDcUc1Ku6uaB
4Dcov+D9DgtXJ5xhIXY3J+LaMGsDxVcD9kAldeE5bLHaJaoN+k0o9W6ZeqNhi+Xgtqq7fZIJskdg
r5E0r0F4nLG1KO9mMg+lUFC3VBl72OsmHYl62E8IKiVwPyJE28isLXNpTaclQwu0fa5R/mWJlJ6P
sfwy9Ga/5xMofS+k2J4oLXmhTi6SHwxYeJKBl+AYkR0nc6zZZk4V2KanVF6BM2yss1AYovRSmA+N
q7kREuE+v+clF4mtQQC3rZkRikvH4eHV46bpAR5KcG9/shUcKhhGYl0wocN+LK3DoDnRWwSz0eze
Kxz9SSo8zKYd/SZFVn/ekSPBflUjdyk6T/MMq86AkLXnRX6FigLdbmnHIWvFXA1iiflyl31SBe4W
KIXAaDClwp6i+ZRnIE+gTTcN8qLNOZCXEBCJP3xjsNWjRnPU9OotrorYH/HU5ILTjBOWw1mc9itx
ZKvV75EB0FhlDmdd02wXP1aQHQJJWX9/JUZ2zm6FIMAU798hH0cAQV/pilMvKOGSuQZz8SaPIuw9
5237kflwLdGRAg/yiRibwGrBgR9RHaCm9n88xCVMocpc3qGgE7bE5sNT0FGMS/gyRI4l0Cfe46hu
U12c2eUX4v5OLqCvHnz8e6sIqcyrKHZEWS5fECWhw0WHe2Gnb8vwb49SXpitshOR5oMvq+ttP2NF
Chl6+8iTvM82L0GP+rN+zR5AbAsXboVuPumWBuNqA30O0GC5XvU2SJs9DCuK62RX2pw0bAw49e8B
A9YwA7huUeIjqVyMa7E6aRuzOdIHWuo/dHDHcJhCSi4iSxxUvtbzIOv23dNcD4WvdXXl1Ahp48lm
Js5EV588n0tKVa9AK+qVThLtB5HKb2Ix5L2MFCC3av1ICa8oYRb3edWoXnRaiNiOyAOMBHMb/Lb0
SOqLcDZKGxYMICxzuTVJ1/eCMATnQOG1dNTy2Ynf2XKv6Z21t0jb6jSjtE+s5e9gTGpxuUSm7Dy1
YUZaeOOT3rnkPkHrcebMD7LByY3HSLWnBpgM/2wGVYdKWcrMyLsXxCMVHX+orDhqC8umj2lAOFNg
XWdjs7s4yFztMNNCS+ZmUE2pZfevzj9A2mLARrxcKqrJaWIicSKVQg/ZWkrlbjhq7j0S5uKpfc3J
G/SlmhB3oO7QER00sgpaltD1QXG9eICUsV+0+KtPiOys2NCAl/AUBpU69ipPDMP1eYQncMOIBUVk
iY9IPHGhSw5XsIqLYS0Zsuai8KJ4EZ2P0LCQcxb4/EGGVbYb/UJ2lvf1FufdUC35GfEjPOCwTeXe
NKLXfgK7rqMfAyN1xGOFd/rvv14z3TIC++yKrs8g+j39ooCHG6OAKfN24F8slQvlAwHPaBZw4cj0
XyI+OuDbZXWd3w7tNeuYYJ/KsKQ0v5bLczrLZ/qhUntVy+7J5sXy6Qz9pfZ1SaF6FMczxa8G3ouj
sbfQZDzcwrW7WtmaSGzL8kR/xjcgb/LKOPfHscaBpxOOgZBxx+n73bkdpZT++KTKb4UoT91ncXg3
NYRDEKaymI9gSpyggEtu5+c+W2f4f4GmQsqacosg1HtMahGBlmTzT+0QdEBexYhG7i2NUQLJ1jPS
YmE30BsofTGRj31BqmD6EFqZgnIeAzG5iBU4xTgUVFy98irWdfuAaqswWF7pYTKMCqZhrbgwuXr0
97pjZMqndZPaBxhtrJdTarj6MKYBNje6nnKkY3Z9hWQCG3hzYqKiQfaMoAnMcPD3W3JDIXEx2WHa
g7nUyWa/XKgG/QXRm5mYVfMdlZ1VOF7VZx268NjoQn2XLiZyCCW//uF+r8fmGh9oAsIhvJTrNqs+
lj3qLxlNHAAyLfjZfc4l079XOgK+uD4zMa/LrCIpqroN4I1OJoJbmbS4kN/fRnpTupNzTBYUPXsB
C6jKaMojHY0HubV8mbEH7yBeBwk0XP1e5qVhK2hJhrhaGpxCifQH/KULL9xHGp0U1pbeiNyGgX45
153nw4JpGpVP2BHjo3zoM8peHYSpqKQFuxzbwCqtfnf3qDleDAEwVnDW4C1fFsFNBCU0deTXS9Om
UjhRVi54+IgeC6z1/n1aIbkl8VYziiivVkkMpqRui5kZOaUBD9PZJ4v6LYvEYOac62GGVpwLLoDo
ZjUs2fuvpr+1Ab6vWvdQ432agsPuud0OqI3qHa0M2k8i5+HRaoyb8qmoG58bVNzHAhepQ8PNr0sW
Y3PCRwVibMLcGZz5L0wav8DYDHbVudi4jr1tHXJUjzuGAJ0nQ7s67Ld0sqalwuSRPGcMScFhIKFn
LOLPbHN5iQ8pH//I5u/gb54Af9pnk6c6EEx1uKo4s81orGv8E0pY8QrBBsbIFhvJNYSVk6PqoRyI
75CymKjU7CZb11PhQUbb1o01zTiSlqb+oFnTrIwvNGI1+OsKS5dRrQoCgbmh9oDUUZRjSUp5Mgvt
KRLXvzKrC2hIXvPBp+O4ZogdTQcdpaY0vpd7UjxiroWUaCV9Yj/gfQqdMDQQ0q61lpmZLgW1Q7p9
yjLWzTfjLvOdob4ZXdnBdguhZhNFoA3weq+hZu+c2aOqgcLQnPfaRAvP5JhnSPPesqcZKRZAWBUx
mP62z+MdRwp/xkuTFivJhjJ+4rPYwBPLlXt2AngLidvMkdHWluBXf8d+UzSvyIhPBKGWt8rLJ9Bk
D9SXG9PXXBDtrrY4T3kFu0wU+unmhjLVi1qnApp6Kc+veZj19JfhIxFa4R9uAXoPHDixg9/vobc9
Ph/v4+safSFCZJrzr4A0LQ2zZ0laTlGsQzWiAzobLBcNK3KehlIiSH3WRamZwlQ/uL2+6NT1dCDm
XjrDxmXFNHLoZLyZ2BDoSYn47zwEl2IHuUWe0JsMcMBVR/4DdqbBHn+cZF/vBt87xlQW07A/Ud2s
KuzjEyhVZe89O1yKm7s6upp5KGqRIkFNRzWeZF1jabAiBxz8hFEuZyjXMnLY/MUXFvrCI1KPsjkN
83akffRzsVcak1f+adwzQKqMDLU8LqoHNN4h1ohEIAWdGnowxUqQ4Bno/r4a5tSdIRU7wGEDz54Q
VfcvypcgzcI3LbhNjbbVOKijQAoHL00fyFmqMMYWnvdnXboqreJiWdazKMxALwtL3cizLkMSevBA
W60mM8ngHQtU0cMRWSzu6ix1LaxGueRY9NQ4/chKTWL3rigQIg8C3HbGGgT/7FEojKP9eYj4+lxS
mrFBIBTt7a8xvKHg9oHmmkYEwLbB+/Xwl5cHzPQ+3cmvpVBwP89nRsl010G0kexA9JxcgHejE9Q1
PvhWd8QUdMz/cjWknWwGsyVdqVzba4tD68Enrdqc7lFV06K6VJPiX2CPpgBrVlXvT55UfhsLYsHX
Rckorn0UXCtgQOoI3QRkEzVukLO7SDTqZ+Q3gRLwyETv2i55KT6xjh2FhtZiAEkcalgxpnxJ42oI
Zf31OSVsefZMUaUp1YphqXpzKMw2JLGL1/RlmYgoJ0DUlNnmEZ7KWzk4BXRqU2S36mL3aMBET4Yb
iHpb3sNq5f1y0OHXrSaa9V9ib5kdspJxo1lYop1EX1dDJcA7g6C+yiNawPS2anqsIwTcRfHaMFMz
KoDWyY35PmSVtQfzQDSl/IYunGYEOTZCv1ZzvcEpe/zV7Qy/ECj13VwZ4wkQLMxOmvpM+5SFhvrR
SAVcgC3yk3JNEnUj82POSffKFD3hPU6M5VO6Y4QYKmG1XYPXRq4DNTY246O5JMt5jiK9MVExRMjm
oBzJOczqlauyJqpavcGCnN0n3Kkd+w915KhUxePAQ49MB/0dX5RpvxszGZ22M2zLGt6lZTo0GE5B
Biz2I8E4BtoOpsgBchq0kgid9zD9YCf46pDGB8uLaW8PMOUyJmxohOS0OnRJI5UeZLsEBLtdRQnM
W5McwTBtxTXeyalT9f4wtTFZvEOlKj8ew8GHQNdy2p8RnExK2yRHEcbH9dahjPb+ESOJDQlCWsRq
xnUqshvegQ3EEkh3Ut40+pQpSR+Ne18d/4y9VNuusZKFSW0b2HsBu41r4X+HLGDhWI3EshgPVWMY
d+fLK8hDuXuh/Rjc1Eqt9Z6Bhlylcp7RpBhoJdZvTfzzEsYvP9WjM3vLNsvsPWF1n08y5n3YcgRJ
nI9HdKD0+xvQaacTP+CaQ2o25GZ+KfHvEicDWMlvgY5KzCbmZxrul9nMOq1piYT9jPmzKHHSqMIJ
yBIw/XcrdXqqmF3SnFlfH3zgOrEWQEpHDFhzNPIHp39k8V8vfbsCEhj2qNJYQ/I5Ip0wokRgC0qB
8jp5HonFFRq5o0dpcFzBpTzIAv/vZkugSzkIL1Z1MQn+e2w63KommA8gtiFzMjRRTGDBVXUuXG/5
t15xNw06IMxN4S8NO9A3AvsImBEBzrV0yLKFoMb9OksiIQIH0Ut+5wUH1LRSe8fROMIbzIwK9uXv
CAM3pWZwzjytuQmaBZtN+VIQmTtj9fSEkzyHJpPfRI8R01/jLVEgJpYCbRXfYOs5Aj0ottgimRPA
B2krrcQDWypUD8whnuydzuGVPZZvksFbIUkgFdOMZbWx2U4JifUOqhj+Mbz5/8Kca1N6ez9+AATN
gqpRKr0NxBIIQKB8CjWuiCGsEM+RiJiOZXRA4l4Fr6nJvXQwtlrc1E9OHmJMbojGqgGqt00kfI4i
T+63atvlTdCuSBf7AlUn/DU1C6eX7yJMnMikKi+6TQkyCsM7CklthyvdZbU6Wdt/b4gitOeL+jHF
1uIDEINZH/vKKGo9aiGOirVUZ51u0jI2+BpqRZGmvrUj4zBbhZhXFfeXn1rmaQZ1qAVmu4Qtvpz4
nNYiEKgPAm86NJ3L1sg5MDcR3Vu/RGXhUNZDr3+7QSxIGryiy4nWhCKVtVJPtNo2WOVLh3EPELrm
qIXoYunVreawaEwziND+dVhrS30FAONmwseVHhn8kcoz6BPDrypjtW4RDKVRqiDcW+bsgcgD3O9O
HNX5EyaRmt2gmc6m1uq2A8zawRidVseucj1avf93hRQ0/RVIkFKKw1DnIG169yRuwA4aFQjoKSNV
MCZS/cpg91kI4RFU0sNz3kdPAnfMS3K+WMNfbfdyFykmLZYI3IOExxqkUAIXkrZXfYS3xVobZQlr
Idj9eun8y3M+y4lvmMOfyTpGhfn4X11/+YVCb4OuMvEkiIXARAPfOldW8TmfolVqrBKdHX4HS1gB
3RuDuTPVbZJCSC33gU69aebaFFA9qlF469oiptm7wTo0TcghbDmS5+1DOqs4fok4F1JQypDc/Ils
MJj58IHUX122GhHAdhFcJwj9V49bhSsa6/b8ogWTnN04WiTL9stB1CnF+pF9d7+mNRPgtirxlzz3
Gn4C3eFHlH3nCGtbFYxXFbFogGUrVVZEKSPRAA6NPuuUuW2QxNA24dua+K5RXFtzh5YSwzDs/+gV
fN+Hb+aTrmyBuGKRcBRfkOwgFbMyArSEblyU8GJQHiqxFvMEJfx3sErM+rodTEWr1KhrySdEsbKT
jiDRVbJuhsOwOwPz5YVgEnxeY6jhJSYNn3Pf5jlkQ7CIHqW+yGdErjT+JDlzGjD4JrxfaoLrooTe
xnTTgqdq1tWwyPifb3Dop+w61zJ9FpavtNh+oWInAwagHZPteniou1PErZsAZ3zi5ouVVmcnjNZg
ovXnA1GfCMbr4js8jCoc0D76W88OP+k06/s3+VIrWPrCO4/o/uPiN7aPdNHeCR/6ixoVZn8UdD9o
S0/tWWKOnK/YQ0d8s+1Az/fZo4xbSrpsQndgPBBDClynqP3J4zAeWyJW2Y2tQjgKi+1hj8ZvWMvs
HXapx7XEuI8WMTEktTwt+AzVQI3VDC8J6Sv4QcPtN+69DKqsOL4X3kpavga5Q9Vfrdv3RhL5mNES
3BTWnPx1r5RvrnVwS8JyBvX6vEjKi6+hnM4ZS4dJ59Mo6qU5ZeTA6psUdjQQzPbqv+T6rV4nE0oh
0ZAg+PMqWNFmvuQeqoDPK+1Pv8THt8dnYvO/gWIiUu+vQ5IAsSzyfZx414ZRQY7MBQE5F4Jvtiv5
EQgIwWArYccWs3UiUfSRLt28ip5x/wkEEmp//qatPKgmb4AHvIhSAbVjjR3dHtOWMd9xo7npn38q
DT9qBN0oVwRqPrs/f/9MtAsqKWmb6CwnYSbXQwjobzMzUklogWX7fbtDsdEQu/GngPWusXKi0E1/
Vi7G7Rp9A2hPj5t460NacCgdqeYzWzqOrYWpCaHiD1lVSEt/+XfgWu4mVxv3m3pt7RFa6kOjJgZ+
xHa1NeZjyLvW5jgdDZ3d3PTvg9/khe0LH53a6u+PIQdH9eSSJ01B1VJ6jIiiYoWcgW7o3MXBh0D4
Ns9fRQGGpIQWE6aB8HWZ3gAm0yJBQrkVcbcFGOqfqSPVQOOS2lJ/h5Nsf4lsBmLGzG7rtDRf7Cpf
MrscdWOczIglxfWtoOxVIR0zifZFQOg2DwMvzrSEigMwGy/EvsK3JVBsAO8CF852LBzBC+LpBaSd
Ud08acRfjmcy+Rb0rMh/tH8c24OA1eALJo/Ub2Y5QF5erd0DApOl9rE+PWVKlQvSehpY9geUWCnD
A26VaYsK5W67sEzAJMIo2wFmDAGajAs1L+vnuuoWoHeD7XRC7i5dgmjNnT65/3uC9RYAwoAEpc+i
lHj8luwITE9EZsHhK+5vy4jiv3qIlX5R+LJKW39bKF/Vd2mWvgAdGbOn+D1SoZAD7Lz+VbTkEtW/
z5P60Tksri8syOPEcEdnNwiT2Jqm01aBta6LaXB22ToUcIzLv9JdvDvTDzyMr+O6jHB5hLAq50/w
dTenkDuj/xH3kANDlEy4NFaqOifK3WpGRVXV4lGXxAxovDTpJKkc/ALYPiwyZze7x3Iwfek8IEne
Uf4rL7G8lsd1eLgm67x5RmYy9V5FLQgZ7lKc4Xd14MaC4wfMZ6BH4UXuleey6r9vOauG8rDd/1YT
j95PDE39Et9YpQeMApZKWHB3eSJz4tfwFqkMZHAysqRUdiRQ+qj0+uLb1F7rq2MVVOeHx+uAz/kl
0GcZ6poDRGMTCovY3q98TII1hOAh5x3V5/1EVGEIR/IUveyyrEumWrObuFlR/aBIJ0WCsn/n+rYA
Dv9EOcMpTrntKfJtDjWQaPCTrm2ZJEMUntkOtU25/LFcvUOUJY6uLPg+jj//jaxyDGx73G8tH5SB
JYON3dnFI8nVErWTx6kydoilaxsN2RhtoR1B34oY68YcVf+vScYnFAuRftM3ritxcvOJcizOA4yE
K3B1y4SCtOEcUH3ciJyprovyLjS55xb2cZRt1Vuw6C6PyVvFf4m+EQiB8n2BD09K5QMG7bScB2+m
H+VCWvJWMC11RD20T5yHeYF/mfyY+v0Mc0mgh4G7Q0vZR7E3rhv37j2jKGtzagzgZyZjc9YZYs3C
DLBaFYqyLi+ymVGRg/avUdo6WUzg5FeRW+UtfA0bf7+NXWCz0F+YYuWT4pICJRuhcs5dVlWNTzhE
kqT0hVXlO6jB3gx4HRsKLdK4wSoKkdrjs1B+huOxjWvO+3essyPF81gtXudjPdi69v4bZMronmWO
MAxsTozSXXyzmZBtC+XXy0FLSIX3rFiDMJfVHf6coFmmP42CffJtg07BaHSNvzW0AVQozHzKGSVV
Tod9QE4TQCqkvNUTVpBbyYYGHKNudbrWY/OOKHIg/yn62oErcPHwy+qpRLuP7jPL4sXyOLsSJVQd
VMRDCsTtQ84kJ6tFeD6jJQOVqf2DJcEgw66bisWsUB3sC9ZQPRZkK2XKeGTmiuXg1kIrfui6YS7B
vxaAqO+06LWiQslGIYySIx+9DopcVDUOyEL4t39JXa9xhPS8Jf9b8HVVnMPWZgvropjwWfMsfB1K
0z9DuwGmCnBP1+b/fWT3UOt1C24VPpzhiXpG5zF30z8PKMLPcHCjnkCbweusDBthd7Y0XPHFg7XV
rxkBZxwt9Nq8kRC+BQ2jZeIEABp26kSPP8yV4EkdC+ljbIykyB5ZGIItwAquL7gvxP7pW7bWKgVH
JGXMtmmbBmWKnOMHc4FKhyWihrHNZ2HyZsyAnLQmyVjFJBDfSN2U4gNB+mm2l5f8UY0l5l593wEr
T38y/T1Al90IqgVLyICVQxQlyReRwntPuQ/qOpRHv4KKNEfnedhWiNi8qJFIszK64p15EK/NTYyJ
sa0QLoxGxhFthLRJr2uzjQcxfK+3ElOXmk1i0UzURyYZNDOvSGJ4SP0AnxfvLaHEROB4hAnrYDij
ttdQmbBen1l23zh1OZhMdFdTQZqTcJumvImoSLCTzzdcfDJV6oKUt34/+MzXxESJQO7utFGg020C
QIoa0IXKHvrSLrwEfxQFkRelsi1Czun1c1trIhf+boWMEJWCnuHX1cbZ2Hj5vp6kYYbimP+A+Cp6
pFv6JhrjbXFzm1EWyQPfFQuf76pxbl1tdqhjeS5uGCRBDadI5cxjV0tKXqrifyt4eON5wqWVvGfz
ME8G8OxMaQw+df5DWHEiGX6AwlUfBbpIMNCt59wIfPTb6XfFnV1Eul9DfBQ+3Gb23nBOwP2/tWAq
WvkKyx1lDNem1Ya47b1W0T6iO2Qa52bD+MrekWPj8vY0ITbzP+4n0TvGqDrtZY98KTfh+V6gU4oI
gTu7xXFARfdy4tdOV+t2GZUhxehmsekVuKI8I6gWAYtHsuAsAnuyXlnpvVBeyql4cEenQ0xAZg8+
k/A4Shb1Pg72O0OYAVmyFrQafD+b8Woum4KQ04kRHI5B2SJI19vQRETILcR4wB0B7BonU9VjYt1L
1WMkeSE6fPA9OaDvvOdNuETvUrUoaRRhnzqrgwPLxiRHMLhVPGDwpHv4fejPYfDyytzzMvK2p8Sk
b30NsQl0WjQCEXsmMat9ra2cILbKy+tCMeFNs+ZCmK7vsFe83k8Qs0aLQrndo0N8cWEKENpcozZd
RL637/o9Kzp/iMVaWf7labpeSZ9EdDR0XVbkQifQhR9mfcArY+RteRvfv5aP/UD0TqvO+po/ZQ89
8MI7Qphib86nFUcBtQAV0OJNR+MXDTiV96TT2nZJicIzQ7qXbsPQjYwGHQ7Nkda/qNV3WbScc3yD
AJniv3UdXv0RSlRzEtvK3n9G7gcrQ2520wIrwRXXvP8V5RDeWy5se5yoqOrd8mVrb9H1VByHNrzk
PzOqUfPMI5HHvNcLV7CTCMHazl3HVlby23xaQyKeLsrBG8BKfv9idHN6ScmvMBrcUZHEPFsynTrg
Q0ia3nvWepXMsVBfeRoj84JEVy8sEwbSE6RC6hmbTAEAHP7cjlsKPdT+wV09WcjLCj4n3KQogtQI
HJWpjBx+jScwRZaS5BLJ0vmIA7wMnZT/qK5c68kpcbIBDNoTFN5FCNJxXt/+9SVKUdyJilJvjPoV
JUa15T1JrznA2Kl+GF9M1gjCYf3drF6eQ9eJP6IJTWtT3XehMtPsHnszwPCtXCsaSvFWqUjYn2pk
D5L4T1vi/L9YUaqfyu96qSNIIqK9Hkv8CQCC/+NbmYf4Z4h402Pz0Sj/m8EKHLYWdbk36e5QecAC
8m57N/ign2cdyelXcYOWbboYXDWB9WDQW/gIpkxkVuq5wdY8/t8+8UyyA2+hp6cXqANSIR32DJYG
uDozwEjNR3cMfvV4RtUYrRa0HpXEI2pVenu2ZaUNJTV4yGfq8i2PT0B37TRKZX52wR98YAnniXwG
e51PxBCy3a6V9vGzofkuXxCxodDca+MZEgCbrgN3/ZNx9SPE+c5ksX2aQpJSWDU6giqNhS2MumAP
3b/kKPDzuL3xPJgaKiwBqdYlYDdtqvUFCj0o2uK1KLFMckOuhQ337HzcH5fFy2tkpHmlt0Fq/q7K
yYsOGtXHjh0dqOXlTErN2HtifGrGgrt1qPfgbO6xV7+FSBib4Xc4AFPPSVl569nxgqqv9/mU3Vx0
zcBgAti9jndTVpKoAL/uEGAq70UpNv4oU7LqJI81TiCDrzBwuxEQxhNJg6POq4xgylPk8sy+HOB7
ZZtCFIB7yfcbzdWl1/M+0oaz4+qBDIl3t+kkmmSAlC9FzAnDyL0lEiTTBXPAKlFjKLQy1S14Xjg/
b64q0LFBc1xueC2ADrH/XTmNXNErywo4DgrrWUvSPgW+UcHL6w0QE9jN2PldIXGLvGMKx++dH/QK
/QNvJDXQXg0qz6umQRZfUpp1yegd80ugdi08QKCGYyIgVI32MGvVSfBmAD52T7djimP7Ti1e4sdR
tkPLNF6lqwalnBz+Is8mGDPhf8XKKBwJvTx1PnievF2yn0ZcLoZS9kyEKuOapHBAS3yNA3aylp1V
WuoU9Sy35vTtHY8Hq72MHxO0vJX9wVNAzB+Hj7t15bO5vuRBujs8vtt2IPW/pTAIj9wVF/XZ3Yus
wGSMDj7OzaPL8ceaXq//95RtRZ6a47C6OW/7Pi5DGUajwpozLOmDBFqBsP6J1FnASFXoxFp728Cy
XzlidErMhNInUSF0kt0iUQi1arRDONvuADuo2man3TcN9Tglmr4BR8WmUQ2NDp3XrOkeEL5P/bnq
Gk3+ljkA5smm0OV7ROkal+hlFups3gbRBSr6yB/cOCk3OXUMN2aWvslZlzUVz6yi7v9umryHTbVR
/M7VERPtJxQULo3myRamOWhWvfOFThmW2vOOk6km8aoK43C1QO6QMFcKFfWhF1TwXYEVMGcIZr/E
iAI2TXW09xOPowKkbxaGMCc9WH0anHW7W4Ch61ZJ2cJAm3oRxVnchdaeBu6SbrThX4rIaD4L4iaX
esqv2pNbo7i3lhQ8jJubo00+wAGTeECMJZiTFolSo4CQHRBfdve5jd3d0bzljF6A29eJVWzJq/82
r99yIQ8vC7xfsQ4LPLKh/oyNokcZBDTaRFbKZn0oIqRqAFnoUOdS9EnSXEBzNw8odgXzbCavzI3X
BrxUx6USaApFTmjElRqugTMHWAc1SYPnNmwQmDjmsoJrvLiLCPFsY8wv1MUb2BFPQhrrmcTwr1YK
07TIRLE2ILTaSLxYnbVLvroY6R6TfgthZ3N6CJuLtwQPG+1Ti2fYhKiww1flFzURn3ZkLHDj3m68
rQMqhbEEKYinopjKbn53rg6WhtlBVxDq+J9t99SMqRllVmqJ17A+kmOxAMN/qGubGJf0ypmcCG1u
QnxFu8hjjGZxlMC2XsKwMqNslLiM7KDfS4udUiPD7dR7FrZmT6Qq18KLuT9qzlz9K5R81vZFdYCm
/4PVTDVAvSSbh81gRNMdm+c0xJS34h5qynEg/3RI/1147KcRXrXKIjLOJ7xhJzwg6fXBtFeb+9sX
IBSdqYtyYeAZwHPHk6NVsZu5p1gk7LA8BuVFBY2ZEOMh5BUK3nx3NHgEPz0GQHoyyo2OYU4b1v+M
A4qOwwxuRuqJ8+aeOEAgXM8yUjPGdYof6aHgENg8PPrImW8JEjtfasU0EcJpk4+uuiccZ7SkBkgA
XnXlhhyib9tiiMBVwviJH0EP2SKSMLGYwVThjRd2lENJDutCyhZENSr786gGdZ+VmU1amZv+JjM5
u2mRSqIsi7agG942NR15tXS4OtTGgl/x5/mkOjF463kRcLJ3ELk31JA2i4IpabPwP4/hE3EC6Td5
riRNtFMcVXK4kCkZuzi44NL3ulNroAmB6LQPiZpUe8wkWyF0vsGtzCTH11zTLpSXU9RXmgLy77Ya
tomz5DQgIkEjKGvmQosYVEKMwy4Sm7akbbbHs+l2N9LJUEMqyYMyw2uRJ1hfYOBQs2oLHfNDbslg
ETaLGaSY66wch+Qqc//6wMcp6ivPj/iYafuWBV0d1uRZ6xjQbcMubeJETg0KXu9u9TaqrGHawV/q
m4aY5KM6T5S1MWpbwp35kTIvS8P46MD0EHUg/g3U+R53dQShKbWby+wyGjyi+FrtRWRg6oyyuIQZ
JjM4dl7a1lOQ1RdMYUF1MuhO+3CBh0J0ICbMtedWgOjvcHd4jV2ysi4KVIqkMOT/D8qKXgcG2KnW
vtna3xg/XJVkPDDk2NwUviJmKD8mpGC8CL4dTYktjqP79VU+u2EP6AUfo+swdEzjviFKRyClXrv3
BVkNNDaPxI5CpbJDTF6Jz/9AyXKUbQ0QHR2uboFi+EgENOBFacxHEJocXm3EVwM5bPEFX/mY8l1Z
T1nNoBZbXt1ort7plEiUNMRt4RntFBgpLiPeeJzEqpy4znRx56REJKW+eI3SSb8C48dH+9eBVEaz
x5KrYIzyDc67T1a85N7kN3WTIC4ALxJDJG7yT8yRv55gsx6By0RMCcwbVc9NkZ6YiTtS/HPteI88
O1NFY6S1CwkdDGsbWhgximUoggAyOy4KvCiM3AypPySZggNnYw+mAbWBkqYrsOHMa2v+aN3WlzCv
uS6+yKX4jzlm0RphQg8+xDE/Vc/fJzNezzpT9HEhdmGFt4pZ4Eq640AtFZ7YlvnqjutGZqrp2G5K
3tIrkN7LiYs2ocKH7+eu1pJluG7WhCe/yrhrK4NIHV4SwCqHkXjEznRlFBDf/RrlLjNKBWoNm40/
mQoLOTg+dIkxLbr/GSsRpDd8AdnKpAuyO3lHAz5hNRJxkoK4MzM90t3LxlJMAmctP2rRDWd+ve0w
hPepEiPLNfslUp6mlhDk/IjiAIWrdbPw2Uf4AC6/VOe1elRIRBGETckt/RvvntVMj+w+zrXFsUM3
LKvMjF08UyuWNCpsWPA+h0sGHkuAiw3ykJmy0tP/pdNzXEL13dgrQenGa2hlFrANfaW2GuDrYdqY
OKnZylel0GIV2EnU4zWdWMuEcglugolmuoh3Qsd/OuyQAXOvuoytFLc2/io7+P8ohvx6jN/Kkh4i
+D2d+ktwGCzdKoWajIo84HdWXU+3inTdjjnQAkC2QgaZ8Q516CsKUyflHi7O248hzOLzmLsHVFRz
xK1/KaFllZ2hcphQjW4a8rAd9qJyZCWfLcNQq/hibNeH0ueoCidDMGD7sb34rwmImxNL0Hkn2j+i
LbnuMVjRuGfXKughwlj4CX4RLgP4icMVsyK+Bg93umLXwTdue0IPhkQ3BK94szwSZXBHPn8S37iB
FT1d21Pghtfa+7bh0wkGU/BP8A4wpOQtuK97Tmav3I5M+wZDyYO8+aa85ms0nQKAbP5SZZtoQOcf
JBIoKrVST8jJahff1smtvm5E0OxvmQvjtXN9TY7rtJ1kir8uIkT4rCAgA78P19Nsr0NzKB9/BJmY
M+JpjS0O1geA1X/vrxYyW7CaTqQVRHcO8f5OCGc0fM2WSqRlzDNpFfnqi3TJuhLktLxlit/XRqxw
PqeRT+hXWkYGcDlnt84riQa5yUlWX2rbiZ3GoovesMp2R2bPh2/cNKLtwYHrxbJPgZeZxPp7ATo5
pNWfFPUcid6fDuXU+YY7XBGHnAFbvQr6QLb1QiQoldS8wvqyMMnsluOyEflQDEyjRqBxts+QFmYI
3sesu8fVB8mGeif1FT/vo25ixT9IxSjdMahopbTMRcYChhTMT0q7zDSB8R1ym2H2KJ4TA0glU5dy
U8QhNeWt+OmHz/ToKaSXwM4bqF5l3IJWcW++ZP9pF+uNNPcNkpUzR798T03w7xcYvSDZU4g1QIXA
O2C++KY1Q82Ec/+BdnwNYIhxqPZot3UOK8j7ZJo1U8wrQN7hx6LJCiRE+jnuLbC2it5Mlrrrkvif
d+UEN0zZfgCivAr/ZYT4jF4Lg1r8bWXNquaO2/zGqAG1+bt8rHtkhHv1Rh/jwQ3Qn4d7aXEJ5oep
bXk+iM2zCtynIqHyV7end+Rk7H3Nb8FuZXbU5uLxVu968MwGubs6Jf4poWbmN3yu/VTnMf9zIcEL
hcH3J6yOlRyOKrf5/0SzS/tnfzRw0Kl3KabhRlOoReVKlxlSn6KHTy551DV9WprUbCOi10Ww4Znc
N1SGvwR/DESdG5a+X1nwoW0vQW9/mMI5TLY2w2sWVexaHCV/W8DXkBzZxtTtL4yXkXFyEbMa0TJ3
JtObWgRbgXVoYiIn2CG/7gsqRCY0/rIuZRce9XMBsdAeqBYm0dgMw3oB/7oAkGV95md1PU/K+GFP
au8DLHJemOFFceM8HbQlY+p1VvtBdjiyltwLQwUAJUK4KakgDrBXhGeUdZLzh/ZVr5WgtU3XtAAh
U2gsEtim0lqIMc/92FjwlT7Ozkqa6wd92jK3aFZZnfzRH24yAnUaoTje1faoqHhP8XW2TzFRo3cI
7r9uUIMs4osRtq87SsjDdBlosyPATmXqBdqlogHgM4AJ8ezcMsQCbBpyj+nmPC4HT8hgIBZtbI5w
Satok+bQCMz9ZqKtvjGGRPb3ms2Q7qnJZAaqRHMdAcEwRRboE7v+CROOWetN/r+oVqApgGOrJqPD
aE/VAc67J9i+dBtpMlERyBGMkiOgCdMtoBpsKTo6YOqV4viGsDkBAQL8DaTgqIJ8M7AMxcIO3/WP
ToW2Swi2oovuSyfNXYH/JrRM9EZ4PG8uGvYzv4dZ9uOIUsFOkyLZKk+tO9t40SkbK8dGkIOm2bRM
msti1mQ074pSyj3VrkSPfMVBzIwm/ZnzT9v//IkmOtl1e8QyCLpEG6D9F2DBDxgGDE+HxDvKV/hQ
p6KkJS9ARLQlFpMidMfgTN6FpkufQkIYFdN455ZjlIVMAyCG9GSDq0PXPEr6hz4UYL/xKI0/M1EL
ntRHGSonVlIngyTdq+UL7hHyUeHYv4m21Sij8o+lne+NtmASTnI/qxwzMnPlkU3RxoDqJEFKfMp8
dfPtFlQ+QGQUAS3rMFNSE+SmUKZOBmUs2KZ1EhyKrntPn8n66JTiiNzXxVK5doqWY3ScvEX0h8iY
686RStk2CJuyGNaYRgZbLiD+Axad60Ky6nAtN0pUG589JoMteVJfdQhOMhN0ETYyCpLDtewMLRJL
LF+P5Nx1ef2zIDkspVA7l4RPLyD7GyucZTT2/cxnn6KN22azLjEatCEJw8Zl7dKoi+wyD27FT0fe
tqHMO+OXHazcN6m865rq4N4G/5w+SsXH4fQ1oBO5XfDW+Y9NYtogWVX1yXG18C9En6sdUpE0QloF
iqM2ZVMpfyDUAnNNwVgYOYVq4OMBRqjYiNbuvcEU66zVxevEN+u6to3mnnNJHnj6Ga8TTZUehi3c
1h2yS6f4YqlsJ7X1QErtkCjugNttVtUC2fyWEkFxjmME89GCys2czQXQqulEflr7T5oH+8fh+kvD
sNJIUWuZR64UwEWgBxsCS9pAq6cpqtL7dxg5AaADD8gKzwop88Is6doPqx3wnTJkNXQUJBWypC6V
UukqDk2TaIBEo5FX8sfJ/BHmjwbQU2fqGc74BUjHExLwpc39u3GaBIzIbfJPo4bJnyenGF4UIc61
fKolatVn4WUh2dTfDidi57WFQ+hpSdFSP3zvWOcsgH+S4yyTS3u4rsW4Lth10Wgf9nC5KyAxvz2/
glftmHEH0Kws7WbO7lIZIUTn9hnN4uIyJPUEJDL0g6Rjsba9bNGLsjWK2eVgrxeRGNs5mFS20ThB
mfquCPL7R7pXzL46zcSuIvr+NJJ9P2hr0Wd83YR0sSFV20JwJIz8SY6A5MTfaNJuV+rYvRzijelQ
clGslsPXvDeIM5665g5bMaKyZHbtiul1yYOfg8lIlOHYrUpZ0b+n4ETkhJF9aaNF+TWWrRy0AMAR
U2cA31EQ6Z0ZuzNqcprfZUxmoBY+HBMgJR1s+IaSLpJlDim1qW3QuuTEhIrLrSkLFMksfcrK04rD
7uo6W3JBxzxpR2YOokFUWSPKuyUBWmnHjP6vUJIqJNHMfeFSrhI0RSof8XXwfEGnsv5skSbxV+vi
rG0k5PMH9+piM3lCBGkCv7astsQtGlEjd61UQPlR2Ay48MK7XeBeHsnI6V2F6KlY+QRQpPakm4tO
B/ZDnEfPF5U2nQvni31e34NVXkVcQZQ97UljQk7K66kT6mpHncSE/YfXvF2u+3l8sV5Wwp14Y5dc
gVDk3pWG05OZ7jlJxBKT+OEW6brxp/Gm4zPektzS4zcL1B1aGm+S/nNpgjX2RKDqjtwsyWDJdgGt
Dt7mreaTswzNfl4nGEJayf6SZY8K8on7jwFL4gDePakq+j5S5H5ExzTp0+fmFMrGmHm0MAnRnMGv
+tVRAv2l3eQLpSTuNzXTUGVNtvfxq8hnk/ZROSxfGSHc7bHJdQU8qHuDIN7KrLdT+VyasDmtn3UJ
fKo5T1HIrWwadSpUaQrvmBw29x+rUbzC/E7uhnZgdIYtuXTZD4g0KbEgxcXhdWymJEP8K/J9UBuz
5wHCG+kyZ/OgDbXsYgf0hR1dbfRa9Lg56T2fmezHMDk2GK7L7OmhJPna7UTJd4msHpB+0wfqGeo6
i/lkigJuetygHxgpXh/hoytS7ZeSlNxknQl20CQmUFTF+zD+4zTWf5+afyyaOZ8+yPoAK+hhQKdy
3OmVV0RypwpJ2csDcxYh20YYyBPdFCqZdIetdwhW1SLNOZ85Xxxt8amDCeUBhhA3heTp0d/KVAwh
UOrczkTFomNOX+AubSYRn3YLXFn0jtHTD9A5erSk7PVaJI/ZbW+c68MgS40EwtR6Nt81k1BEYJSO
56mYmU6E34cGGrB48BcyuBSbUNqN15U3NVsKftG0C22Y6ji2ew1+EibYdSMbKhitAsV6+8OFjXLM
Y7KE5KSimvxl1KGkvQjnqD0kHOZmESQ2Kbo2VjfwCvVZUMMs6wiJtVM74IkvtJRYheIjehAkkEQi
2fqYIlRldOUvfgNLwqO++qUtEXdf8x3+H6OgK6nDJQwJvbWLBZW42G7gsE9QRCaHiL/D30iSDXDr
nDsGimuuOqcE3IRS0v0ILDYF7NxpJpnDZ72p+NWWucwh7V16v4EO/qn0mwYl6RX9eR/70h3jJpXK
uWKrQdDC9ynRnWdqBzwvw77hq42y36FulKpNh/EYKppTa3DGdvZuZH9IhcQBLCPGhLtZHqRruNok
jv5Xayhs0Er+ljlLgksztT9TRYBGd19X8n5gsaEUbMk56M6+wprGpWZs0x+2xGqICbAL6Jxm8hVn
Jl5RoA/B2xjLfVuIZPEdjc75YK8TJd8YbaZ5Hxx5ICFItBeglvoat9VJbyzzc2GAO3td+Nz8TbPh
edSalrC77jUNm5iO5o8RG275P9ErHPI6okjUFQzcGW76PeHrfS1Gw61Vs/3o3D53A8nHD6wGSrgX
LDen8kimCUaJcwWkVpxhSAgU2FV6XwTIcYTfPtK0F3EcmNBRcu2L8NZd1ctvlBuJ0IhCEEz95W7d
g3YHFfsLo7ANW4fks50ItK0g2b4kvGF/KodMz2cHWKuW3nkShPlvIkIE2q8b2Vnv5fG8slCKTnbs
yPdH4Tvsrbl2lMIBobz9IEbC+SWQOH6LK0VNmXMXmhBR4vL7LVJWdTO/X0thVdcLxXbUWyYOHm8o
zMySVxI+Dntr/Hw5HlNCMVRRFU3nFWgqS2R1Kp1IKtxulobmlEk1ftSPwO0ZqkdbENF3HnU8kqYS
ACN5iKm0yTDA2bdQAUgZwNSjusb3JeIMs7SFWpAJNzCMr51wjqKEOhPjuHrzeWhhPLCg9yNjt7KG
URMkEK7REq0cRGI/WN3y8hdtO03hMBAqgrVdRLdVh0aZNuexNaKJ+da2XHiKR3Q2dzr/Yu01OoPT
2imhF7lrrI7QZIde0/t7j0pRjcPaDIds8OgR3C5BpMiRUlmDmwuvChb8fh2GrKKecmunVbwWrOnP
n3gQTqbbhhqA3IY7+4PUyseMlspVlyAm+Eb59kc7Sv9Q78MI1f90NSwvzzlx7TwZ7id37tO8/4pv
d0o/BtLPp/RjJTsYO9EoNL4XNwy4twpsoCYRx+8vC03/IVPgEuo4SS6/7aL25VQJ8kax9Jahbze9
kzvNlnX2d9LoI2cBXCvQi1FhgabvHCiF1qh3zDnxCFcG05bCXEuhKP3FXWw9od6VJw7xwiHOrZn7
8b9wu653y0xswJylQ/IcTIsIXf6X4E0DhTQJyJb8Sgpxb8oixS1RlSmMZEB/5XhkAR5Lc81NOEMS
wpMPRnQfJ6PR6HVYtPAYsd9iiixfSq9TcuT8LyNBR4NzFEEXfe9k5bXp00rT0fIEVlmBRo5L0zbD
uEbGcAjJ3l+xmf8pzlhwNxc3lhIZAzjpKgBY2p/aXPA5XCES+xN+Ursh1gpUXHzbNGhYjzB+gVJf
BAJtRwwNhjMJW1NtHVXPPtAZseXZwnpjDrMcIHBwzNSM/Bq6ZF1Jn55CBfdtWkatvmOC4NjVb6lG
brpCIiuElfAUWbV08qxuJdtOBABrrLYKb2UD2GlVOhtfaNLMkUNqnYc3Pvi39lTk7pKDMdTmcwZM
Mr8iEcuuhlu5WYOGQflQ3f29L97k4MRLB8N4YDFkohD8y16vT9kbmhh7Qk/iX5jR1stdvG9C5oBb
pTMVCqojJBxMSXd+6rymVJR/KyGFfMcoe+X7ce6YcvwL/gPtMLHyY0lGnWkSW8mz6XxiDIXM0RHO
UI3YJB1kwLTfvMcrc84fitILLHHvTfd3vi8Xrp51GLMk0tmM1a8Snjk0hI6KUvbha4pvCRBhYAtf
zEG/+JGYRp/MxmRzZMwtDsZh7BfADDnsDkYZRDMaoRTq5WPyjTWHrqh2GbtT2CSuBNhmYjHxOpn0
sMvfjucs6ytK7wm/SYNA9Lm/XfWQvqBKEwB0uiJYwBozXdfySyjFG9fgp/ht7GGwD4kokJkaVNaV
3DM8lmlQAvuVJJbO2i14fNU2MKMaO0pDeCEAXuNU3oWzwX7LZeoHhAbeBfAc3uhb6FBrKzhujcSm
zXP/fXqbrOYrjWe7QFwkSRcoTxj4Un+HePWk4WC9/eLuy08mUyeSosXQCiKHBnjFlBusiQpdkpnp
Y3cY6qZvgOMUHMN93+lDsU4MKxOvdREtlH0HNJl5imtf0zMtq/O8YZAE61NhFP97Qz7YxusmjmqH
nhpPzfQlM8s9eVymF8ZsN2AOvKRD92Z6nlyZai+0GxpftDNWvAcNz+vjNZwg+yOchUGVoSjqiqIp
jKuoN35CEYKX5wZoygPc7D3nWrmQuB0iqS/EdyDW6RKVJAkSnhltUkH3TKXS4JMkRNTAeesYK555
oBfXlYfP/7nxXRkDOq+DM3B+nOZJcGqZpivO7YBIErwUtHQDU8Q/mwcjKl3yqdzgQPjAvJOQMnTe
f5q/Xqp1ZvLl2dVtT/6OIbhsmBfnrv9Us8V0CfwocotjdwksDS6WIj9Zzr+We/eM9Bfs2m7RO7nY
qVX3Dz2+2PEMCu1Y++XIWN1dizBjvaijFA3Xo9Ln7Pl32B2IARwlSf3ojVYd2SW8W5WPu38VCOhQ
/KJIj3xxjboc/FgUseJJf+CgIv6YRlFlM70D+T2lsQ5PdJZC87X+KExZqv8d75J/lLtFioiK1EGs
jLTKMYX49eb68wenuNzUHyBTtGgwF0e8a22YvQacR5/cIvvSafmAoT7D25YweznfKU1VXzE61j7+
6jSDJGekIXysiWMUkZD5E/DBQElGRzPVS5ucAJR1v3hT0JREjVVQPtkO7JZ/ra2TEG8oXEaqRWV8
lZd763XpY+P+rSwW3LtlUJnJUxJZ/RYWm0B+Cyv52susjhcp6JL/IowzCYy+GhpxdogysidHJ82M
z/IRsEVDG4nrx1soPt69wCVhWPBJ+sTFI8M4ZNbTvKfS32CqupJQMzdobZgVNzBD9ZSQcTdGPji+
M0YzKoY/sFvk25iciqKJOYpUS9gb6MS9H2ssCk6suI1f/4UFxxwBLQ02j4UnMJ8g7LuLUu3zg2XO
FvxneTp1bxnzhqkznDuw+Ux+BpXcJnLBdGO25KStNfUCBVieslonZ0jnIaFZcQhEdBInWQbRCmLA
JIji7eTukSvykqK3wJTAeHnrgVnCt8TvEW+s2Oz+PXHpMTBAXjz50GypV7v99QEIM5CWaKk8YUAg
acZb/JzF2EgxL8SX6uuJQf49fEokVtz7cMo7/oPYh2Yhljq0WbhqwPDR5zMILguMY+3IV08JQvf2
xfFeXhoO6eH9RCAvzHk1Gh9Zy5egmNCskxiW2wlAb/Et8YBt++9e82jNBbVrK0TJeyCOmgA8Tvgq
MjH+awSVBXA9n4R7EvhBzRkNte+oZzvaZhOziiHau7P65DoUE4wpXPADUM7p0a3nQGqCYuwPWcrl
PpQuwoUjnlg11b9a4WCc+C/6p7xlvRj8nZ6Gp80D2HtqgQhnJx1Rji2SC3nXRmAwcOaeHGCWnd+l
C5dhP2TmU8J9Ry3EnrGztlfblvFzs5IN2xdX1/dMlEczDgYYXXvPoBxnxn8zTJdzTUkbgcuuNN8i
DXa+jNSZqyICvh9ssMTbsfpJbVb5PA+ryzBwZVTYKnHeSOYVV+YqLANo2gMRSmh4sfkA9VhLZHIM
bqlv/vG4cfmpI8sHfp3IWxWqVQpAuAPTo8NiTHmgZNe646r2ilE2EnRLQ2/LQzlEXRGq9AaoiNCo
K4I1MgchDBSC33lifxhukCeI/mtcDmUfHo/5FYEBafYx/FgbyJjNeGSCG9iJaWcFpgZj5cOV/KO4
+nuNCdwAk+kljzoxsEO1XmRaJ4VNM2vPlz6j9f7OnOOeTvw5PuOd4mf2w2QNrYqADI53PYduLc1x
uN4Kz8hZPPOhaXWknZzl8gXqYKci/eMJSh6q3MFeBQAuw20lduy7TMZh9FBfVAneOvfxKrBeR6qR
eNCPNqFg1FZzr5+AX2lwN5eanPnF6oW3DUApcVxLth78RXKda0MPpBjhADSn2E0lLu9FtOLd3+f7
ncQGLn1Msf1S40tVH+PjMMUgo4pI5mzEVGq2NoylUkhS3C6oxlKBAzUd3hqzkbXMRhFa7qEVE7Od
ZHIsay5++vraJbgDPKR5Hlqn1e5l/hbmKBlthyGT5bHF9+Lcju/P+HzW4IwMAV5AxrRLExRWKkY4
7uVX7b/ymUMMyt+uwPOSFQEDHt/hZaGe4K9hPFNISMG41xwgcN6Lo7aoJVjz9HlBFnywLLbpMmY3
DNlkZ8NmblPuTZnhiTjKscDw34H1Aa4/CwSeYkjrDW3OgIcIl+i/H6XQJyDmFXcn5P8mOJnSyUJJ
sTH5tfheVGzYV2A1nbUeHrechu5cKdP15PSroqB+YFB661JhNkyIPzkLpUyZQF3CoR3i/dJX0fqc
ku3ycAdxGivJLeWMXPCOO/VsxwWmR8HNjgPJn+urAsqtM+MsB5bfF5Y+7DMp6aHGcN38nJvEpbTi
rn1GYfBYSpusfq+kFCg6g4sMMxc/B9bPZf4ETGO9cJnwAGwe4n+PoN0JTBdxLn7tBHfT6aFHOM8m
yt3MkGK+wa3Z659qN0uU8Yl9Ic4ObzA7bVSVoe/yK2zoBcQI/Ix4hmxp1Xz5cR/iU+8Tk6Ef9IEV
V0bwmt/ERMnTKcMDEALnq2MuHOIn9a55qjvkrzY0jKcCsR6N6o4CHc8BOIQLWVFLguZRCZ7cTYUd
Igq3UrkegEMwmsHs4wPQBCc2nfyndU+3Sg+QSxIXB048y7c1IYcvv0GofGBfP4AUHYoDk8I/wWv0
2aaBTjuw/e5Y9RNEAiFBwRT9yjiu0VXWZx0U3ZEeeEZR6sYgdiU2/VpFjzzorWMbzbOliyAeIXCN
qWLwWZbEvIAuT2b7+tyvF09fdtvOeHhuT/roUEiFpMh+o1dDnxEQlBOofOfGP2qwmK5Uq1m6/NPS
bN0X+qsrBDJ+hiwcaFX+YGGwgi1KADHwr05u9C2HWUysvp+b+6FUrKybWl39ryl7iVvOA3Cxq9Zw
A6CDU15OAka7NhbfpLSkwrRoRM9n9e9b/Ac8uf8CgpU0Qjt2lo9gIwwnDitlZ6BJqBYgXtFhmDjl
DYkR862XXVA0dD2gjp7mPZztSZzF8f4tdcX7tGdyNOTBXUvgxV90SQO26g1ChlUdTj7Dp7kYEpAB
b/c0uIH/FRUO1BN5ljKaUuYlGmInShJPCLwOMMYpjjwP+EYUyoodhxW0hXh/tWKujnjE4IASYBhO
/XL3oJP0vkXVYwyXG28cdQbXg8PN8mOS7oAZbZou0Po8zceS0ugbFq1YtNfbo2KzQZwRt2LIiCJe
pjEi5tzN1z6aXSr8heUHgo0GPk7JoULUL04VBmFDx0Uyj+1fM+tXC72pSZEPdpvQctAjc1M1cV/D
cUAaeg/UKxEli2PsAeiS6wtyncM8isevsi1msZp5VdQ4pQhLmodtRKNvTu7uahcfL8qbfg9rCWXU
pibOW9S2FCaRjTixWGwac+hpeeGTMIvQ2HqbZMPmTadCPx5/EobKqYD5PsWYcNa4/NiK0P0WYf/V
vb+jcnQ9VqOx6u4kl7kOODWQ3dceCnT+KzKNdLfZ4DbSTbHviWf42c+Y7wDfAc3l/I/0xCnByLLl
3WD6+a4VpRdCJ/mq3I0Vzc3UTNm6qeQ0C1A6wAO/GlIPg6lElSbG33Y9/ga3O3fxwbrmJIha22gF
0CJuKEQsgtZndKA7ZO7OC1ju3ouBHwaTp85p5YyMc1EqnzdD8sjDix4DukWyPbW9lTrf/+j4qA9A
v5EoInobBxCrrM63IUhhWG6s6Dzhn9sgJlGqMi2ud/BOjpSSbSmaufXwOtYhb9ENzpbMSHs2eOhF
Xjyw9l1LPB8QSarsjofWkLTMCJjQ3UkJ7+gWlXFHyszz3qfB29LIw6P/EBMALu5fOW7kYSOIQXJr
Zn0QArtLP0S8BlVx07gqz6HSa6rUwduxueIf8hCaasN5Acu8nEaIqs2TfNBLTr6gv8/XamdVqxH/
6V0rXNGkEOn6jSY4DTNV1urm//FttRNMOwjPc/vyEE/hFL/wlQXtbSe70wEQrDyauqdsI7bjan4w
E0zFwsm2vZrih6qN4evzfNvBclp9fp32+jXO9UCLWh91gRX4HH0gzreohTgq6ePDWM9GGQo7hW5o
2louZJ6hIrfc4436Ev7FYnaqwFaqC6UOpXm1DzdQM5RP7uR7HC7egSft2gyEpStePw0nQMlhndl3
TQHB5n5S1AyfT9KBGTbuRhTizMa5F+ADzSlbSJb5+gFiB0hmnW/Zgg5NfW243MQ+fL28wEWJbmHu
VpI9vQ6nAW07KAeAiOtpDpMU1CdAa4v8dKJYwVCb55nQ4I6ohqqCJPXU+nR9qkn5Nn2GEhK/jeK8
G2EdXDKdWqp4h1DZDw5E4NiQG00OE+2GSvp+wW1nwAGq1k9qhicJAiNOQVza19yfsHaZUDRUjmvb
K91aojLQDHJrcLY1DLlf5umzOKovkz70BB0pwEf2t1Td0Xo/BuPykP5292L/IYNJnmEC01sbaeBd
XnJh/xDgQ53yHZhjMrxMihXiovDZinCgmrJ082pd/BaEUi4rLN9uZoj9XyeZDRa0NZ+R6HzTUhxK
B+esB/900d+fKIC3Typ6dYU8NYuB4+bUFck+SxaXRks5ZBMw6k8q4NG6DgKCyBcqho0CyK+LL6yC
qBqYgw4SENmvtEIyrEdwYM4VA0xBEIMd7ayBq5hpxoHZYhpIy+I2aYXYmmjUlytZ2r47knetHRbM
ePf8OSEm/Y+KMD4izMnOXCVK8UBdHFXSeDHOk4MHjaeoVpHDp5+8A0vNJTDMLDpLaJ6sCKyggtTu
HazqUKca3g40M0drCMTLVCq2cKfFP6PhdcafAzrt9QI5cJ1ATkES7BtjUaPjOrql0BT2v5L7xFan
i7kvOd+WA2MI0e0ub9CPDKEkSd36vNDUF+gJtho0T1v5e9gCZlNFH7f5vCr5qe9CQqh/wEAgnVG4
qdPCmDPIKvBzlLYdbNQ6CEN2F0UB4cArOqjoUKK28/rCv4OxK7KOkGydk4vYXnzPVNr3+pR0+kRV
ysSwDCEc9uV2T3ik/RLWIh2To/ANUJI1Xks7rcDAtIVN4BwkpM8E9oQqMQy4gtNWAxQFHyoIYF8D
+T8uyYHDXVubqN3POrzzjqnAM+vZWk73XMsjuTThgkYPT9jIex3pxLwFggM128iAuN6kY/tN7w3H
0i4MpNFwQf1eXnDZPsPSsEL41iQrZ74WIiy4RujwnBAapB+7JK7UDzANKz22ugETaGFDHU8lklik
HRF8WmpuHbZb3g74rficJjXNxKNNjZUwG5z0pUHA/T/tLeP2MRbnMyiHw8jTGAlGszLhyzd0NXcA
8shx9JjReSvqFLGUBp0VeSFPCTh1yIrt3CAN1cE+EdBT2bI0UV7bDsQydq2P6x3YYPtGIr+AI/V7
nlZyA9rpXgEshulh5cQug4lNDzE87WDl+wthvoVr/QyXrtDRYgq9RyES4EUsQBMTEi/7kijx6XKU
r0bZ5BXkhJ0LL3xIicniUtFJuzRwFbZzAfAv0gEW9VeAhfxmXDA3fTYIg1MIwOAUldcHC9TE2p6r
nlwdeVaYOGPHEeBH3smBke7SYEKiRrbjbuhwp2kjZJlN730S+qEZbyZ7UcQ2wkci4QDipMIiXjGK
lWdb5wtlfjoptbnJZom2oG8AcRT6X/twxnNePNU/KJ6rGca2eHQqMMhNrCAs33EF58JhlaotFJNW
qfuzJZsjMO6WUtKT3NfFV7axC+L65FFi36ZZL8QTHS8x1z513OHqnyhlKcjPnfYtJMY5SKBtNury
QyeOYRsERoW9cQs7LAjg+D373yudvm/646qjA1+mo6pwBYN/4kT/ZJW89TlyqrZ2rhbMB0CHU7mn
gzgUmCTdapJBm5GQeHuxv9JgOeQRiML6SjtGa2rXBFuhkgnQFF4pPtPs+Jls3Fq/s3PLVwK1Flv+
BTE55MnmMzshG0qcKYWMXDZ7GJ9uskIVx15jfWUGhPUiy0opF6MK98Tys0hdVK8kwcihN3GctVkp
hFyy4WznFtiFv13dNSSO211iWk6rtwi8MZRahzcXogjd5jqmZk13+pa3Uv2qxJUEX4cMTqwUptaP
5a0qQAPUM2iFSeIFdECUcKfCCLwOXAhsMBXaSJ2Rg7ohe9Bo6y/aF8pVkg18pt3YGZjj1ZfLQL0W
/GSq3iMJ7NEd5LMKVLoiIR30oRE2vPkoEJ5gStb6VxIWAr0P4VwSp5iEg4sT/NQhKWO+W0eLOK1d
3hBNyRWSBZZq0Ag4L8EKoqwZEErMO7+EcNtE1XVoFRG7sE40gPiubPrOr/rluTittcam3YFFtnNQ
AcNZa/KKYeTBKl4VyUmij5jerKypFVadcUPr7c9jh5a1MKvpLiRpnZW+wpRbC19V6haMtb9PNHKX
fZml68HkGavR1VFHei2/FkgL8kSzrnppJyABbnRt6O8yOOGJvcbI+TNklv9GsHNdgIoUnvtR6iZi
PJobcMp8NfF+OYNFB+CZvy2o9klRIf0ncIxntRz+ab8wjFWMhqAxXPkMpW8oq2ivyjR3FgL2Bq3m
RQmszK9WN53fFHLrUMCpftS92apsYXwAZ5sfmwGeRdGUkfK6u2wtq5lwJXjGdw0Z3t7lTEbgosWv
3NPawmcsknZD0iSH5HWWA90lsiRVyjCI2X3aOr/NGLkQv55cNhN8bUCFUFsafDw26D2jwz5y0DKk
1rMOhUiZSbRZFRJGW4GEBKJIlolByECN+b6DCj3pUQoR8EiUDf2yXIk3Hx/WHRtEJN+YP0QdwBud
PZO0JRobCO1VHS0fH4o8kgPp32FteMEuuCPYuzEpqjke3NyUxOuKGu+zEv2KYfQaccKvQC2L4ylb
IE0aVxHxgdtxJ7DcKFE+f05bMZkPsBn884yccz5rub+uNWSLR7BXmxpsTv6Ovf2qpE5C/LzfFIps
icdcyf7/nCdNSRm2VETcZGqF4mV9CFihPWRExLkj/DRGXxQ1SWlgubcsMj37uFNuAQOiP1MqOJCr
H26zD4UdHq5XREf09K/8UckCiiKcoGMLsxj7EDNRuzsWyOn5vvThGnuRKEgyb7VZTXOC8FW55Sow
qW/EF8iyKKBUEV4QYE7fzGEHXa3l4y9z+er0So7uFYi8eJjTEHVWJeoJQlL2ofjCDsnThEXOVkMw
UQl3w4eAyXjRnyJupcVmkwQQ4sqh8ytt7eVQx3aLPghQb0Tb5CUMGssftUIImqfOwxkwLGOAcaus
RoBx0Eaokve2P5j0tAj9NrrbkCc2AX+2eqfKUvkiQNmwIgXSdDRw+JFK/QkaY0omNa4a8R7i7U1y
ZOok8/iZQYVt2TbEfTLJ5tMOh0N/qHYQ2gyFA95aEeF2PeEDA2M+NYAT7e2pyoZcpY79Np6m6SHH
mQJillNWZUnHVGX/cxz5faqRx1D0SR88uhQChbgDzBgLf0lfD47dJFbZV+SHBw8aPYjALFc0bicL
eY1P9JzOXQaXGUaFteHs3fuPZ2LtWW9T5+k5v9G2KOAMI1SIWJrZupQjvQc76a2tjJCkAhriSpZ8
ousSj5ytjxti+rPlIEyQNaBhHF/KwZesqoRNtG1RiRMq963x29NpG/9AtpVDx5Bp1n5CI9RQDRIh
euNGoWMRywQTt8NZxD14ik3RJE9wB4Y0e519h8Upk3izYt3LaTotlhLKqKflCRcjqSMkBlVDEOyt
LOKkjGlr29GhYlh/klvUHi0cm/H3Tu2DJtP+PTanCAUb0RzkARcNLC9nZMZjiHORgmMr+1vSseD3
JGvXfb2Br3iJIwJr8EYPPNQm8Nqltu1ZnYnQPqQcTOYxVUsAuK9eysLCKlG/BgigYDUjWyDIqWfP
1Ou3ThYufudhHrVMx6raozi8lhEMTbPj5P8sfVIQw7rYa+CFkAjO6PCGw9W15YZuq5NsVupDL5bx
dxHHbRk2Y4hZ9YQ3c2wTdRGrUtqihAWTxHUZFpPS8xyXgk8/kXY/uE2O/21Em6/zDkBE7ZPE3DIw
BW6V2cz76IWubWuyWK7TwmQzzHqS+zemzTO1EN8mCzyXa3ZM7X3YE3fua7Tf0CBkdHt4Mfb0mrCG
rl9AI8bdSpVYV/QKnMpscSN05eNKJ0oHPx/zx9FqKwkWKgCCcy9qG1uNl3BjTgdAly31lO4kE8l/
WEtFxdvzSHm6K019zOOiiHXEqZVkC/nAxfo4DGWhrEH2FIW34PpFlLyvmjDR18RXhNpUnCzyxCeE
rFUGIT8NlbCU1Jx8HSkyEq2sh7nKMpRizmfxBpdqjxTz6RZfDa3UWsW7Yu3+zcUEcFo9UpFRXhPL
qVgNanKekq+vz2bLFgeM4LIn8s5GfwYRBMraekSvVfs37DJCBHZ19xJUq6YoOjQkltnkKdjmbsDd
XByESzyk62sOYkjkr3P3yuuZ2LJtOktZdt1EJGUZY9+Q4kqItEpBWWjk4Vu1PAB/T8QDQ8A6k3EW
4NOwhqijhg8Xkw4Zot9rqm0gpaKYtl6DMDMeeP1VQdgPprw4WerHGXAzTxnAV7JiQa0/GG967+h3
the4nhsf3BJGIlTewunZ+NJ7Zg9taTKlbMvVe5ZKC3bl1WbNeZ7PZ0PTm8r79mX6+Pxp2cwKA94s
qnMOkq+R5SN+ZLC5L8O/krRQS1/gnSmm/kiXgQTFI2jJj4r5lFg/9XHWHQEXIUhpgNDHMEZ7SjbU
tZZpxck8GeGJBEX4OZLVyYXrCQ0CdGzvo0IV1xFxEA+Ass6W46fK1i8+Y2zrS3wsuzPV38wvs8Mc
2yXqOVTGKcTqfO7cMkPle3+/cQywkVBlB8CI5ZqYSjjI1cueA8ZdmHq453Mec3pGYBvaKj7nLocH
mijH6RVMhtGat0nWDr1+nQxH1X0TbTLQ6fVy51cS8Nu3KDjhzlEZOwqQh0TB4ggFvcmqJLLAknxl
WxCoiS/n56jnZPcuhv2T+jmVbYXa1TW2csh3yxqStmyxSurKGu5pkVHHx+PspE/CGwV5u4hJRjW+
1CjCY53ysw1TOjTzf152VYz+dE3B5nHRMBk6lk7rypMyCEYnP99eItZQolQqqwd27QIkzDcCwUa/
Lh4V6Z/NnBdOs/Xgw4/gU7i7s8dYbbd7c9hhK4HtKtVNjm/QlATfDy9d3nM/vtAbosbCB4mms98/
b60zdF9iTzI7gjTPYKQ77bFOyw/F6qXzAO6U6SG/UnR7W7rmrZVNT+/p8tbBhvywBATIu5T+BM/p
VK2Je+HqUajX3NLR8QVU8VrowxahEcVxzsfoxCP2JJOWEcLRaWNewMpNvDYM40eBLPHbPe5gUpD8
4xPk9pTs3fWQDvab7wgt89MxirWubURGeQSfBGTmZGhwR3FlS9bzmWj169tVSYgHILX3DgzHwB/q
xgssC/rOs5p8sOzHCHfdTcOLVJaR6A28JG4VmoJVuL7B89DXj35M0tqC1b1R0nhb4g4HVwfVcTEa
4zsGaF3TOFbz/0XXgLsEMTb61eYXjPiznGiKemENtLfvL8S/Sx2klXS8V7Wht6Q/BYGNkfHomwyY
0+dzl/k8UpYzf0OOeqTdMthwHRDg0uaSit00zGgB/3t/iBQvLezPphbTHT3ibZFRLz/RgsQlEqkG
0BhJmBzlIibeQMkzhkNYndwp7shKid4QbkbHFovgZ68cvIqdKZpY86Dwa7uRi2JpS5puphkhUlOI
6/a+8x/didJvg2O3zmzpq9AdjS0iWtUWDej1/TDIZeDUMoubitvcRYVU4JQVUmvleOykZnwOWA3s
ddtCe4XzbkR5TFLVQMxuctgi73tV/cte8L1Q0bLYSF2ZnIE81saqontJjaili0uHRzqrtyiWxH7C
PhZC6JB3E0SEepyeLM/CbOo0P3XoLAFmYwtcKqN2gt2iw1UGCX7gLx3zkkBNli/N5i6puHu6t2S0
BTCtnYaxdtyPBnYL/vu3SkzypKTP9fbvWdZ3bs7puv2Ps4oF+fLCnhOn/gxuPifvVsLOU7KeApNl
kT+1pGKICLFJY2zAw1Dlibph4340e+gOH6l/1oi9gHwzz6/FIqtelQwMqF5OA/qQDw2n3qUtEn4I
gt00ZNcPeFSHx7rILsyXZp4ZjH4KmtZVJGODgEdvdEBPADpcAL9nBghN/05nZHHqbxBzPxXHZpCF
7dUgGT2sc5Snz4s6GC+pVhj0ZRrvUA+2VqVQV5rkwQYdk4cri92t00nZClSf8oc5IF4IDAPLEQM5
MPIUe+3rAPVWRDDB/MHX4ItPAqOZeffO9kv/VkCikqgNgfwhFfuVhpnvDYdV1lD14WSHR68yyWjG
sCmj5HbPw+SYTRQwzwyHIPuEUijlTNzExZd9wfCxn8okVsqsA0BER3XaymgPqFjHnqIBcEMCoP77
lrz5CMM2ZRWCtX32YP4oz54woixfSX4YSK5rYTAT4OHgYZGAGC4sNGmgH+Tm80hboMAC/mccLaGq
0gtZ2T5WNSl1QNUbK4YvTK3lNf9d2ep6LLoyF3a31BrviJKkLT+2eP7S+A6jDxFxK7ad/dx34dun
wYfy7vTSmz+7ZI6GPBTAS1o6S8X2Vn1JkWVydeOBTjIBk7cY/N+BoxIMKpRuc24tdnO5fPCFRMbv
vHRSD6D4L3l2PMWp1NTu3yOhY8nk685+JxjCRxWUV1pvO8Aw3QYYEbIwzvlZhhvguz8Q4EnxYgwq
5r+t9SOfy9WOhnk8Z85jlHHyLGo/6unvGF4czT946gXFASX7h5udNX1ZJo1ASxfYETL8oYyBZWWN
xY5JuIfL02ubLce0utmKQF3eVPROBMBXTxlU/ZiofxOZ/DPoWdrgWqiZPcT0Glh8FzUWJjNoZt3m
q8atcPkeJaXgTVHhW3X50W6XAgEMYqkXnemHox1vPqiVh82Jq+zmQHPSnmqdCay7jhi7kROIfjiF
vcxhZXGLMl4FLv7IewNWfHRddrrkxCM9YRWtg/RqvQsTrJGETtS7X1r+keP5IWZ0DHC5fUDbETuJ
1i8PtnTXknlYLZOUgkdhIAuN3zQQfotZcQBJRnUVCAkj+TDYn4YsyysramErE61YL+E3ZlBJV8wU
sw/KRvCJuiRAoc+jbrqacadU1+c7Bd4IV/6n8j+ohK0QbUYxx7tiGjZvBYt9Dt5jwHDwyEh4RzlP
LDoNS06Amxz8YdLFD5NzRX6UDvL3NA9Cw/28n8+j4pi/+plehbHjkSK9XmPX/NA5hcC1g7+AgcuL
FNTVP51BPNIM1oMpmu/DHhtxT1Lwvh7zXR2iee+83g5H10d2odCdQfiDc8utHGsoGxtGdI7lIPx/
b+YpipucLh3BgOr8K3LcxRS6LYdfwTMdCsgeEQtvwVCN8SYaJtPzzjljoLBVquPQ+eTPhl2+knbS
5bh826o4ghRklJOQLeJ++/LKVxjCIbheIGHsLvUKrLwwyqA/eHFr5Yi1kGVqXQsys03BwUgUsXx/
XWWLT4M6kcuY3SY4RFZa2QgCay/jt7uZPIQEImtdOTiSv5/4izpp8QsoxOktvf5xSe+l2316Oqzr
4FUYWmRfv86tep6QSrGaL30c6G27mkSDwImM22W/RQOasxxqqDxN8usEHFgN0INeA59FSkbny235
Ij3xQW9ZeE4B/IIlasJnAlUNf6QEUkLr1yqS6EY+6hJN0B8/5UbMJDBPIAorUU+pqM1PSStAmIR4
NCYi0PCWfLef1i8mau7VfgVTKIbe6SC1JsOPhAet0Zeu5N5FW/IQUE/+t6vct99MkGcPS/WsqZfh
E3Vpf2lTycAVP6LcSqFwNjg3xt7GA6SkAG/YkoXOdTGkj3qWnikqgTnOyafBFFhilyN4YBEPj3yD
G3fYtvsSshkP5MqziAlnvX6aP6fc5FF2hi0sdljENdOYmKRrIQChwWKspo+bb6yey0Sfiheg5V/Z
vRKSEPKcl5aReLFH7mkqpZxFyj1bObXZZPevBWYNlxstlwcz4OrChjSKGYO2i19CCRgAFoF081ei
FLIIEJN/ehk3/DZzr7hVvjC+PqjydwA+gwqeoeP2FqB2tODvNPas0T+5QCgUIUxAII+O4kmjfUu1
nkzhTjDqmis0hTYTBczxSvITNZEemgVp/gDFW+p8GmPA9u2WwXNieOoDR5pvgFZZcaip1hxvv9l8
D6EGEbVQlu8f/69pvk3vspXn7KX1+Ss7z2O1ZzTZjUCqoSb7EJU+GWv9+Rs97qI5T6YTsv0NVBUg
sCAHVaDod7oRHY0PUg1OgLhlCGrlzcu5zy957rbZcD7F6tq2riciNG5FeBExcTBFufl6Ge1sc7wy
o9i1qzv8kxnhdnmFFTRni6GYTaEiFCe2hfkNkFnpegUM9AZt/BW4cHnuckPOaLW+qaF68VNBsdPF
r64YowVJridZmdOXwqDTV94oAtN1vl4wsFSxGgTu128OezDEB8lpTBzD9WMDA27fyILf7/ak4xqL
FniOorOtSWXB9jJLh2q6tWs7X22I0aT0zhLb3mCKxUpvJ4S0TpisUThAwjj/Cag/5J3ek1hMMDyj
qtBr6wRTLUedoLM8ESNzChVH+KIkiUjNnlIqelj7EXY9Nxsr/+x7yZQIfT19FXeQBt9eDP5ocZ0i
2wcz9rbCq+gJs87XnYgy+LIS0d2cqVFiAzxnG+viMO3A0juoo4UDAhMB38BypBBI5hgP0/snxKYc
Gqf8bPm+sBNas/PXLoX1J5B82SYA0xaqJsHmYPVqoGVlvA22tL0qwEXgNVxuT9V15glwkIepE3XO
o0eM9Py/3qAai8hgxZy12YSzrrzUs2znwIn3xtnfyebU1bAOhOgeaytzHU+8LEmxKs5Ug49Faygp
hjp9uCe9ivnMzTgpHW17zbXNeEORPw9llIY++SVe4OITYnlVgTb7+pFpmf8JHleZmLiIq4mh3o9b
t/e8ZbrPyIXgBZ+jEIecBfZzbxtsuR+m527JVzSkEmjYIymOAG5vXwJH0QfaC/4Mh4TPM1z/WgC0
MtVW8aS4rg066oR7sxBxeLqITX4BzuONc5oaEYbPxGt9SLDHi/Qe1SNoHqlw6pjJPgA+LV2Eehi0
T7Eo2NqLFYiuzLtkHerIJzhZuWTutjECj6FswbawFbvuDH4H7Uim7MlSfhb/iwaug6TblxaOhffr
Vcpho7NYbOzy41OCaZ+cX3E/Mk/+t6deson2MFDD2PoZ9uJhODDo9eVJnDNP73p15Baqdy8VamOh
sEoZC05a8W5NRGnFsje7DyZg1K5eEzKsTRGygbPew/RB+F11JPpNFyTXwii2gElKUEryd/rZ7FOL
iItm9mZLWnimPQTYZODpuu70cEw8FbSAqxW8LKzEy2yTZDeWit9iks6bKK472vR/3/WsnY6sm0gc
RwIQ/Nb1DAvgqrWay/vxkNafOWtf+5C47Tr517dCRjUnQ2Km63FvqW9hHoRstAELIoiPS/YLNHGV
KTb/OauiGfGeGlk+8GjZsdP1HnSYOYWsGwbPOy/CURO+WbmRqTVmD8VtcHbXasBSwwiCwnUgy1Rr
lXvS1X5WpGN9oHtFG5LkY1ptVfKxKisx/XCVuV6IThlUhWxtky+Q+63k8GFPQr/ekjmo3BRUFSQ2
yXSIOQ9/A6Fk1LGpYwVp4S9xdGIFNEFi7NomO/Z/n7FmBp0pIJb5rEn6Xywz6rgkNLDpndc8mx79
7OS1A/V0P6sS+PbKobGYwPs7TGAEG7wdCb+qEHn4qAekBC8Nw5Luc2Q0pv1ijPdOzzFEEJAPqDlP
U/RsqRplEG7A6ZA/6SdXkFIC0YjIE6HN6K5SV2jzOOjJFSORTeAXS6tNkvWzJgBxaFg+67i13eSh
JGiO76onOrrH0MlxhylF7VYS3/dc4q5URaO8klOfZXZ4DLs9MeIil0wNNVxa+8bn7T9L8C979koA
MTUXQSxKb21/WtlthvlZMtezIL+C40rj/0iXnsuxEk8zzknBwWnCrhmqKFLt4qLWf+7wvI6vtKGA
GJSjxQcZrxF+K8a3fBnXR6HYkZEE4FJUBNvwRtveSmNKf9C6/VJuD0dLAn8ZVnVfUc+0xk1++kVt
oUUN1+jNZRmVtEZTPagCinjPST8uzQ0l3F9CVJWqkWGKAW8G18FQJt+9DvNRdfS5avpNFzf1zY/Y
AB1OWvZvFKcK1B6ca1e8fvQOZiiTJFf2wD2yvHn7X234BKlv43qSygcpZ+nbJnGkud2paH2zF82/
S+KAzSV0eqt3/tQKB4q/UXlLhCFWAhwx6Gr7fuMeVZAXjORlEDp6Rh32wG2nUIm9z3f5XvgWkshf
V5GReyAIE5/8n406h1dCsTrt+D2J42rPh69QNCSjHsBG+pJ7XhuQViPQcsiQ53GYhSSN/HRxD6GE
qoTXe5jYLUL3sxilj3G0ie91a0CzAC5AnNduzQ6XdwxjmczUP2ueTPnyRhV7t9QPlwkhlVB8J8cU
gmqmNUlA90+AVvjb6a7Q+ieWkAqbG6qykGfKBP60GsmEc4E4T3/+2ENVA96hk4uwFI8GqLpyFHRv
I53pMgd/rI+I8J52f6thVvxjxDUTA7O0Th7XU40TbrX+IiVKKR9qKN/X5KKtLi+YbBM6/xklqP51
NaiLYuFO3Kpid9PbCdgXn1ANeHFaOiEvNEyfRW5e2wuuIffX2NaQLVwmAB2C1nKl13nGOGi68ttp
alrKeSRW/qx3kCzhNR2O74TSH3suGHGqmoFyBN2cUsKqFunngSs5aROFvSh1XRFYTzAeh40H7oEJ
Ek6mpe3PqpQ1liDw8y4/+ss2H21PMMTnlDfm+bWyZqs5gDfJ5cNTzG6MsdbfsoOPeP5IpsPG1gQu
OZ+kqRNb0iMSwhNLoetUxVWJ0Dq6Sr12Y0hits0Ov19Z+b5bA3fnQP9xsNysGf9Oov3LATDYQq+7
XZTeD3ni/HASaIgRYLyoSTqBXdL+5v9LQFNx4I7vj2gHIY57I1NLpdoGfn01PfDBkaY6FQcdVvUF
6IJQtiAVF5Pwhx1LbiLNV6zvkj4h2xN0qjSc9pj3u44ASlC5rSgHtEtgDibHJ+qtiTwJ9WrvaV/f
f9DLwrz2CwqwVBZmS5pMsYoIMs+626v2YeYVeIkkrS5s8g7CPsZll5jG9Ho98i0PbUpHWKAjmWoE
lwk2jYwkfWDeB4bbOBaE9ZvjW3yIElNsjWV+P59cT3TGOx9gPCdaHQfyRi402i9twgXjuPBepPUL
/Z21YSNqIexo40H3nsDVd3c7aosqdujRd678Ufd5YMqEACfCFjqTBznq5sQCR+BpmadtuKH30Fd2
pzvAVsxWcfLb4lDE8f1YwKgjy0vcZwSu8bcnhzIJBR96xSNQuLQw09mFXqWSq2olIEeURu6jXMsB
Tke6B4/ROT+SemxOjEjO9M/D6CIYByevlsERwdRDYu9+JtzbkXVhqR764E6Yl0yN682KzEVEUNnR
I+9btix/p8Nva77E8NPsetZXHpHr2Bjtgl91KlPzAVed3jxtod2FT1TVvgP5fwyQncJMqFrEa/c6
7Tu1kOYyUTpQ1n9mSw/bTKSHyLCMvaXamiHQJsSJuRgWk7KBQ1EfVd+GEgYquFXRNvk0s2a5J7HH
QNik+1mGEltuWSGXtDjMpZ49BReYALHIbPMrlwYnbscB8Cdl454/S9Y9jKi32ikRln657sSfZLAy
j4AwbA35UFB6p+Ij9BDf9VYoMuKSO2T0z2SbkBIOoiG4hFZJTejWA9nRb7GnDBaynMLjqXSE32iW
vvRhX2Zq/vQC+LhPtoke2zmX/MSP3VdFVAC1DMEAcQwoy6NtXjDmMSjVOPPZPNtp3eJnGTnFU2xT
HhXssUaW5MGfastDBtpkE+Zei6PJgcQYOaAwqWifFX6WVQSa/5GTtRVW+9agF+bpYkqAeZFmesyo
urTHnI67YS8QRgxmwkGADYZbNN6Zmhm7yWBYm80zbPd11jbuDCHOdKMDh6RRc7XfHvaDu3VHtokj
+n9u9AtaiYMceROuxwITClqyArQQOokTQ7/sOelXBzzuAbTYnJyhhgmNl+JyS2unq2tnhONew9gT
LCzhiCmug+5RFWBfXoLD74Y9rDoCR6/hjtQmULTP3OZ/zw1CU5NoeyBGLX41GugfUYVtzT87iJP/
Y3+uHO53KK+qRVKl89hCOL2/Ow0nyCv+LqUN+B7YlWJPI/uqB8Wfdmy21jkgjFTwX54X69hxN1cO
Ku1Yz24ycWO6fO1uVZcDRytWQiPddMxRHhPhi8WlOHhXgDZKT01X6pyw/5l/yjRLf/ML+91dIgoR
msogxuTUTHrR3/PI18Ts3kSncJFIKhwNtB7zI3af+IUh8KWRUiB6enBl4XcBvNskHX1eEJei9b0P
Twe8yU8EI3H+yEMO0oLPY3VY7BuRd/l45WIpRDvJmECmzZy4wrtiAxJs2a/IwAHKonyLdaHugLC8
n88bMxNqV4VohhtBc3g7Lj7jxJnno2bPQkbGmYvWqiK8MIFHJU2rP2O3GnEqYMHcPB/a/3+mLl5R
7j0HL0KKkNPUwOF0PagRZGBe9mTPLs0OqHwD2wIbpeyEn1VU51S8e69VVPbczN0bYLRcI9hW2Cj0
f+87jEd8DFGti2jytGSmZ/pP1MPNtTZ7JOAG2xms1viZg5fYrkE2+dVs3GRch5pBeDg5z0jIfhLK
3ylLIiTmEGbcrkYgiqimdd0e+2RgLnbxsGC+3AaVTVZjNk3OYXuTcdWHdsKTV7tX5Vjn7uvVPf83
qMnUKdGqJ2VJho4QPmGfS0jsvAS8RRSvTDJxPZp5F+QHSu4Lo0zJmu8Tl6cugDM4RdSy8320x2Ce
w8wv2C1DsyWXgHRSyUZFQN3i55/EXc/LjkdLxiLRgDBHcJniSEwxullniTNkq/1zqu7s1euCxCD9
vJHqWva5cX1+PVU7L/KzzvjoMCnHc+sVMzK+ghq8RtVf4anndV3OTPH8LsjSj2L+rs/8xOBaoiZX
e0aep1v3MIV4hCWlTr5K+Wx5ovNDfZpjvfwAf0yJaz+nosPyWOZZ8HO8L5JVufEIUNCjpDIs6sz1
J4KzxT6JpXN5DWmVSIpadvhZW6/wnZTzdtqhx2yxM5ftiO+S7na/sohd0bfT+/WzYqHuNHM6XyrD
cx/JXGnDbt8XOyL6nMtXf7KLpEitxUJX3NPjoho84xcydgqqye1oh0iJmR0p9jpnHCqGSFgVcSLe
TkbyO1OoouJuVRrQv0fqO9Iz9fORg+eDwWWcg/bK5HSmDEbuA/+WrcV14kPYIxTsaUsH7g1ywplM
ZWnV6Hp1+vvpPTMidEO3PrjUNG5UnuFXDM9EtXCMLUAjbytoL7e6nkrHoM4foAiFY8pCJTX5PUX3
gXM4UbEOhjV+uW+qeG/z+4AXeoRu8yJ6bfuCCPc9ggq6CK5XdwGfXtrq+0qJb2lk9B4GEU15W4Y5
rdwnpiOLTiJcxTTZaQ4qkoDTmiCjfx/DKumNC6A9BUSVA1RRO+0HXzOTLTKUNPaFJAdVKdqFmihf
eHX9Z6puxiv2Hdgng0RRInULTozzP4GUscLxuOUc4DrdGjpD388QCS1/4f5L527gcpcAJ/lodMmj
1XRy6ReAeoZHRm7gDkmsYJY+89D8087CCb15IXUw9oEgk+UjrDRkhMiRWFb/+ERQoPZV4R/sMiLO
phlaM9WhLhUBVu1ti5dLHwan0kKHvFM8mmR5CMywKB+2dQJlXLYgXkasXViCDUy6z+7o6iT47G25
yJGmEvnSc88gTaM7VS3Y02KDxf3Lj6qs4wIiMhtp/Ag7FgSpskxoF43naq70+umv95Xg3OanY6Li
X8pFC4qIqfbNvlQHFuyv0AH9q8ZWzh0ZRKDW6YZSSVdN4TkD2hr8QEih3Gg0rKsl56gDTZqTue8Q
YI7RQk4Pku4zJMv7ac7GdzBezo5qeMX9dhW9/+gdfV3zfoeL9S7AwUrUWPJG1bb8cLi1cu63eMp3
AxjrF4JmQNXyQwvmc/FjvNucXIfmyd29xjT9GYPtxAokU9ilTCaa1Eo5u31YW7knv3KzuIX3zvGs
vJJZ8JfVWANnU5S5ECjiXk3Rsx3Jiu8iAVwd2SHS9/lHzjoq4+GNHycXu/yQQ/6pot2/1O0n6t/t
XA/nD2JRDeKklfErjYXpFgyqEJtaZAOSnFkhgcL8mbwqRYBp5JYKGpJf3z5PMZzbNEXjE4qZubwP
2Q3VpyA+M0IlcLOVpFT8Cv2SUU9R5EYB50m+v2qy8KKYhEK6V3pkVoy5jiz7udSV0a7XgcXIJnj6
C5onJ+3G98fLG48+KpeL8vQ6P1PZqIbVyiZYqyznzBwmUinUJ6pSc+oje3r6iYHWkCAcTN7MqlGa
z+IEigWIVj+sydyJHiSt+QZ9zdkpS6oyIECuYwQDsBaN0XFHUNltAo/j73WDSWYj6FRl3W1yV1Wq
ot/nuPFxcjtnnLnvi49xRnJJNnfUs+4Y4JPL/F/rMiL+dGxJnCRNYre0/H0yNzndAdURMVHm90Vu
22pX+XjV/zRTAApf0shz54Gzw8yv6cZpDk8keaSwadAAPsLufhK2r/w/+dw1gxSzIw2ScP4SUKlr
sI3BIAGlGMO81Wa8PmrvtUMdUH+6wjMGzK7SE/ZgdV56g3TGnNDpqYY1vHZ4FZzWyj3h2lEk4Go7
ov6nBrpNNpSSXz0aMP48GgCzP0DHhKxHd5jvf59Up3/W/MzdrDDoClh5DrBSLQYMsJ6352whmLLJ
Ox/cMJedHsTaUqe7eAwmqJHJeAOvSAi1g1VsRjd+TRsg2B3ID5JSGjeohhPZdHaXBA3kb500BrNX
e/4IONObAAe04dnWkRo7psK3dVc96G70O6YX9zmYNTAoR5+gIqY07O/Xzwt74rt5J5ZM/Mq0ZuiD
nvbew6hcTmIOEU+Wp06MPSaAqmhqpoN9ijpmvCr5MYLY4bFahJztajvJ27YwNbynbllqwUnfGqcN
riGKGdOQ5qLIZBVPAwPMsbnHi4B3rV/4cpDcnTwzA4WNXIIDYaoer0C+P9J42Z1vcdbpAREmVMio
TKjODg6vYoLfA36N3M19U1hhFAMgSU4L8S1P2E5nPKrj2LqUZxRBYR8gcLehT+29cWx2InRXndlW
6R+M7cByDZsAcLatT+s/yPWsX5EU+OHTIao7dbTkwB4bZMLUJmj9Gw8LKo3v1KXGqX8iHXTvkK8f
UaJnzZw4NwuLe/Xj0yEkl370alkiTtae3z3vaTtrw2528Nlq10pffxECKQKU2KIPrqzfz/rh6plc
M53KJOFWF8u0x0JqRWMLx5Nn8Uv1ChzrDBzQ2q5WQ1xC7CPTrRXfkIX0OM/EWPmebYwVfNwR4FNf
EHYYohHmbZj91kkAwqgtYObXUX2K+rWBPY2x+2ndiVvMkBGiIBGnha+YJrbsPbnPBq0z04stdEuc
Q7F3Sb+/zWVXPW50OJUBUJvn09G9Rf2szqMMZJeyFyS5vuXaavBpxRQqeGwf1twQwGicoctFKwQD
9PKufZrJ4/57adXA8BEB0WyADj7Fh+A3/uEfeIqG1+/jeDHcOWNiNq4V838hiiLtDtx5ta05zP5t
uXg8iaWMQMgZt3NfWOyY/5VgjPwH/YW/3v8mqONVf8HizvmpAsbCuo9tCQOnw6wJEtiXuGSwVPTK
wkepJd69fBlnjcThNy4Q/gnRXKeJOZ4vZmEd2oWz5GAA19UouOjzSZ+jHq2BvUs1/ZGKku2oJHUk
+l7uvrPwiGy2UX1F9tE3tzi6PVyus0PvA9QUT6Jxv2VYqRoe1FOgMSjDVaRH0cqukxPwF6LzUsCL
yinQgvc0FizQ0HplSS2Xl/KbvqglE/uMZqw2fPYgh5IfbjBt/rLR+rxykc4iUhI8wcppGZiwr/P0
BOvvTuAykK7wbVZMuHVPIMQvKhrsR7vZN7Urit4CGxloriJUU3jSvYWPo1UTGjaKp3Iq4xAt2466
Qj0twyJnA7hMm1n2h8knBOAWLj7Ufjhzc4WXJBoZoWXPDrBNZ2cPFU72djZQjIBBqwomhwjUtHsH
xrVBRRufpPAOw2IBy8Sl0uIBvXZEO4lm1zbH7zC8/Lgqg3Y12yQYB6gTTOiyMWoPeH5rMmR2nxb5
2n0ZpxQG9iD2c9lZb/Rva0h8ivl3NqIhNFrBN2lAAHS3MElD8sdnXGo0P75z56SGjwgsObdR4DTu
YXTZuIrMSfwExTA7P8xiNCyqf6JK7ZCY6ckQhEiiPlVJ5Eq8t5mkSH8m7XpLS2j2W7LmUjX9t4gu
OLjAtJ2rhOCH84yK0ttgjE0suSQwJx7vXXGoRN3ysDDUZuHudNYWyfb3gIQfBAmRjstFKulbW+51
oBLMm+D1J8YNDIJZlSImTnLdnW7ol8NA42t82lqzm19hpsUCi4WdU/WwQui9CrPcOZ7mfOyVnWbe
kv4/O49CpUy67e4YKd5dnyO2wfe3+iiTF242aKMQ6NqV19z/TleyKLqZnHu3GSFk/AI6yLnqVGNX
M9fQ1KoD52Hs9Voh9rq9KFQyxABdzejawqlpqmqaseo4bqhyUY+J8PaOP3LOM/T2ZQJtKlWrEQx3
Cx79+zr2btX7XPovaNBUKV1N1cq7R6zG6Z4+0tADv4dJlApS22Cphuv9xo4L+4kn0tcMX2/PrO/q
VhVDSKLoTJ+YHwAj9vnT3+TFgA/brV0fRKFqOJPZJDHZl1uuqaUmGlYaYnQ1RcmgLCijsF9FcmPc
uD581G8lpeGBEyDHIgnvvh5U9uxiggvRjOj3UypIVpOAU8m4I96IUOoTRavgGj8k6b7Fgd6CAxhs
i2H15XCV0hLC9UfAo4qgL+XtUoLSC34pnDVonC31GplQJO8JejIMK58o8nFncgA77hDe1KxFO2Z9
G7ed4V9GJ/NF5COXIafvj/dpcbzyyYhARCIkBbMizdtTbiW0M/0EyWapmA4kxedXs/minbaBl4g1
vbBUHm3nA5QnXKfJauyA3GAQDkcEfr5+fyCJA9lRC5NTMPg17dKXi+geucQZheH5u9Zz928yPQTd
28tsxfb3fWYo1rNyRAIvhX6yUCowihIArmvdQzgyYL6d25yFHC3Ufwad9RKX79LeSD728idB1Myv
IAtS7ZIXJm488mw4WUdmUYewjaHkMgbwuNl8XsSgkdT/rf2Wkms1Q99HB6ieFB+Ao47RIOivOO+J
ObHGZ5X1qTuyGjShtHeRqP4nO+ZR6tadLG4opNkX8AKGAGM36NtoLC3jIT5tB8r4iOu8xfhEmjR0
x2s0thqVJDJlsMtOTdUgbMJS9XegO0xDXyUUn7f+6YbQ9pdymG+59A/BcYgiLXXWyfIly6CMAP1q
aQnkGKXWoFg7CK9DP2YowbnlktLB0sc/H3o4OJOGehrUYjseb2ic83otFoMOeBvWaecu938qhwI/
25n0Z898KFlT1jzJchDtt8a4mWPcostQ1Usrj4paUAZ/85KDLyPCNcMX4mHvhFuGC7w79hcK3Wlp
n19+QrxzYLTinr/xrmbB4IxT/wEpKairMxXZAT0RSm2LAK+u428Cd7sUpx2NlVTjTcoW9VEGTfcr
ccoYjjcDSKWnjdk6Gqm1Dci039UQOoMF+ZZ/eFEBWdJu7YEOwYLjq9k7ztKc5wIe99l/a71xWS9L
qeXdhsnSelylbR19aM8SUcoEsuaFk7NepksaE8j0WQ/F+GU8et/cMkgZ90PeD7gAgKMUIKx/NN6p
QTDyCIir8ZWjpS7w4Gl9Rl6bEUMpfyr1OV2x9F0regqVj+uyAzfAMG+1wDFMOw/iskUIpWfwTFPk
Tx3PxQvBJDKTLq1zfBxxjsvi3N+JbbLSpv7oXJKkyDByDxWsdt+BCMe/VN3kKUP4Wre5B8ILoEDN
2EQ2W4BgO9K7fQsH8VQ4QZdeJMt40K0RMnJyBIj7Qvht3FOsYGBbYq5NglJzyPvMORDyDkFpjBUj
MSzpG9t+aH3g71+Pf20kFUZkFXOeCfWivh3ueEQy9l2GkHA3rWZiX/qpjsycHluO75CKzU50zX8H
xOh1NQiraP1dLKUz15bVBFSOQkkBB9+kC4zgyrYLZtVMXe0PuEiNMrvrfJT8FuLPuvh+nQII2NOs
kp8N3WLIb+00oPeUV+1Z1hxX4RjkXqsVm8vCU/lhbZSOSddoQlk/emhR/EhJ0xSZiIetfrY6yJd2
srAIUZiKgU8vEYuCwDjPphUWBnZXfeZ+Rfm/j9DsyHqp6Q12gLRGyNJgZMdcIGRci6rQo2laReUc
cOOX/GSAqUtKfPjQ2TIl4XWc6a/1yjfgrFmBQlOp96RkdkVi1duRKrxns34o//oRVn6qx4jZnWXw
hDZsotRTMdt2Dqa5Vwmq5vBEYGeTW2k7mkaYS/kxk1B2VjPdcb8MgGY9YVdYamBWg0VlGjwJxepe
nO7CCeLXJkOnqHw/NkEx2X2SmBvwon0Es0+ARlMRtAXr7jWRboc9FVsSgPEDzzGYaPEKLL4IQGlU
lN5oy4NDH6q68ZTf3w5EGWpvqvWcBQ/H5PHcUaSb+u9s6XhfHbMF4TJFYnp8h4xRe9ybNYg8Ketd
jZGN1u3pxvLwtTsX/3mVKNMgIbUUeNfesO08fKS7kX/lMsuzp+YrzXGr3yv4vXyf+NDAKviJ4LTP
XrklHAF6pQPSEt9l61Jgu1DVmtqbgEMiCRb6c01ghYHtST4kV7GmB5c9EWV6nKRgY92ElF9mtUkW
F4Xyg2MR47FvlsdIPFFhONs1D5gmeCQbcAuuRut3zQadfDPEDadf2n9hgjNT3va/dHcgzIylGXaD
Z4dhoyF2cWLEQeO8c3dc7hxW4fEPJZYFZjDHRWjgDoSq82wMa1YyTxGNa5ojm7NMC5byNiGy1HXF
gbufp7djUDGVxYEAmkgw8tfpo9ppFrAQCWTwbJQs4PGy2MYWy65gv9uIF6FYn8fgFj5sZGsNB+zd
Ze+rX9a5aT5nSLVJfSz/5NTRT4VSB5N/3D4s9chKHtUoRCxzVs1jshWyUvtLsi8yCnokBagt3pdl
j1OP4FutZaF+9ZgQbgaLMN2tGPXQ1XecM74+6DA7ky8FewQAhdl942XzYzJEAzXTPAqS5wEv7N75
EnwsVHhvRjnnUvMLRADdqSH1sN0hVoESSFPs9N96ALvzzoH+M0vFeSGbbPSCXtuJ0pN1OXz94BWc
RVz5L7iq06T03GdUlZ/ISC3MAyu9fD7jFPIE8BYTRoDG31Ynsoqnc5QZ6isvHVaDmIAWOdF+RwDP
b4yCcwbD2mPy3oe4Vx/sya0Yz7zphIogP3ot3ER2LPILgWBzyG1t+Gfl+Z0HPuwiPK/We0mhkWFt
R9nSOXwrThttMjbyWmUXm4902wQoCDoNvnOtUftKU4H30gfjxXZyBnAzPJClmTAh6CF6beavsicp
HKfGKS/8WGAdX5OEUZctyc3Jx5FDv1sjr1SBvtBvikXEBQMaFgkalZlzkbtxLvM/ZlDNUdwb54Zg
tKD7I+ibZuy4CoOug4/NfmPH4hSMuPN5kHZaijczb/z9WBjVokMRhSd/nRyWF5CJC1vF1Pnl+ynz
uMn8YUNJXdKpKysAkBzirSChv/QWROHbcls9MRR/fig1gz+Fu0TlBH0yOohab1gWqLlglnwQ3Xlh
vxORZ4A7aAm6G7e1Oq3NeWG/pSwDRcuS4d0rNvL++hCdWsivbIYLcbQMYeCe9mOby4uxAfH1bOAM
Q0R7vrxJtiB1brzzy9yrxIw8/djkUzHv1CxH9dDx0C734LpmQVY8L+cXSnIX/RlAVvuTBSiQsGaK
LIp/PyU72PJ4/+dU6ghMN9nZlDNp+In/lB9YOJLlA32MO7fXICpIbiaxWNcWfaQA3IvzG42G4g3A
qlfBINutzhVxs0zgsMfYC+R5J2OWaYcXmNFAY0uxpilXpM4ZohTR+TUwWxrUF3rtriiVBhEUstij
LLCTN9ntFcQ8FPvzeTsGCubf7j8CwQHvHKhvCat0l/iByh2O5oD6bA3XZPkG8oc8vJJa8ABhsjl7
GQEUjH0Zy5n/jM3KHZTAqbIzG6pG01b6KlfkRS9rcdLKXYApNNF76ARGKnVfHE6EU9W7x+c93E25
tkMiTDzlg4RV4jGFBCA8bf1GfwK0/bwPy/4wZrG5iAsNl5azET3JQFD3aU31L7netEsIIhYyZKgO
naUIFlviW8pbLqAqqLHP4N6qCucOOJNEthOxlmpaHOwra2/NXLyGA1ggiCnopNqojTUQQpXhMBZZ
flhcZDFvWcfsT94AAAgN/x5wyd7A5gH01+gLnuEuXVirsZH2pTnB6WfhZrD4P40aOx9TN2uxDMEF
GqIcXQHrs3ZpztiSjYrHkviUsZW3XdEAEWFl9a4Vl2a6n2l8UbEKBl2CLDkSTkRDoo4aWLerfi4E
sOp2PjGh5850wHkCrkl9U9/4VoPuzexi8aDzhl0UEJvsIKsdLZrp1v5FVEviBBsQjoSgRdGgD4PI
aoYosyGkawDjcNgP/I5YTIh/YoZ42KZIuivhdyYfyuPg9fKiseoKy5yb4TJ15C8PUHbP2lULYx3U
vYmsPAPgC/CdGMLOQgF+8zjtk5HtJ/VosPmoLKxQEekLqMSaDECiqfhrVvajWniiGzQ8rtPQeJc6
f9uOn6iRSwYmWWptCJSvXWNtri4klsZQDt74Nxhu7b/WpOemEBFtLVb//wv9Qr0QGG6MHPWsL6Ud
RqoZefxV/Hls6a/F2pS0CzJt2kh0OmKJrBL5Lc1XbctpkCfEkORTaDtRPXIGBcusJj5sPpgbBOQU
aZ1eqp/TfEfMx7DjtVyAIRmJ4Yfzbqv6sbAOSEXFYp/v5g8Gtp8cxMu2C1IsJ3bIivzUIv3lRSl4
WTHvcG1OjY8FfLuC+u8ytEEcH/Zi0ppxE0UDXjTcNlJ/ciQvDE5GIv4TPEo4rkdFbJeQ2x7uee0w
GvG869rqGyopCjgv8KpzEa4tRPnIndQE/JEyfrCiM1xPXhfk3lqgeo/y/OQ8T5OQW9jCzqPMAl40
ZXX2j8EpB60UMQWnvkvBBijKkngZRQsLRTHuq3AUe+zFyvjkBm3F+qth/kfIjRAPO0zg4u5aT2gy
pepiIW0YHiOpVSPpt7z9N1KSkG489Gw4xrpG70/dOpr7a8NrClKwT+yBCcS7JM+kWf1Kv/NOApbP
YxGE9agH1ysKqhANNKcAx9KlcaEq42MAPEhkXqFmaOMTWJcmKwQLJOltXC+d7jo3l0c3wduHMeMC
2R5DX7AgX/RBAMV7qpwBgdJCJZXI7Dh/mFerjp/aBbr8Xair5NQA7bDbXzdnhmDqV+YRc2cyzMqp
D7GGqmmoxuJwbjznnUua8eRuW0nd2x0sTU+fgnb20OhNkC0Ct0aEhFTv1tOUehKz6kHyaohPQGvg
35PJY9lD3w1c6EMr/2U7brNmu1UDPK8jjYrhI0HY9N4DrGITmZ+lx2SdWoqc3KfXuw9Q102N4TJB
YKL1xPH7sdTxKbzolNS29EfSOPz/2bE6HRg4tdJvVA3+cwIhBVicpYll6CUkxpklN7CtUPTsDYiX
NaEjNCZzW9uj2DYCWU2eGTRXTj0SdTgSTErNWptfdV36JLXvL6zsk86hHAX5YlnPJFWpo/X+axbI
Ou1mLiiAPwcIOyXhjwdf+4dWQ+Zdxy62jtagIiFsi5y5YPZqhz6vd7jcegDESPT4X7w4NFZPcA5Y
0grIEm2/kDY0ObgP2mbgnJQDZmnMgPOHQ5k3ieDCL3/2GUjiWFMRe8sGacjgi+hj9cKE+AXRyqyu
UnEL+Cd8suJjWzQdfvSRPAqn1MDF0OngEqOVxjkFX0jfBylrY5YzGp1fVppWATMhf0fEsTk8+5+Q
foFj8+CcOX+4E6s3vSwrp5apoprIbs/CfJYDbXTyHlUJOXN2VE/2otRjGOIxG+usmnZcsn1o6mOi
U9B0B5kUrSUvuyDidVdXevpFKQDIjYqmUqLh352HPaslwMM00nfehKUT92CgoKP0cgzLnIjn9REm
oGHt2t39yrhpkog4XjqIf0jwzPC69lD69ORp+1N11G+0c7pnEMwjiFB2VKrkTqWgLRk2R22MYGXa
c4cXnW9hRk8/TeouDa35L2F93P/brTr0FNCwJjt9qYug7dlaDulGeZCWR2BxVq3SmwL/OjIqTUVf
hQ9B2809EG9PTuifhQlIaDyQQ36SDhUfekBuSd8hWtq+lW/QX1G14Osv+IZLyR/Jr13kDFEcw44g
kKPX1d7g2wqbsNvluN4DLi8kaohMXKx8emI4RArAJzahOrrq8C7g/Ry7QNGXupbqpU7eMQvNkEyT
QW14Q0Y7aIMyMRJnKXRmVfguu6E+BtwdHPV78PJBxiyHPjfrE4NJ+A4qwWrfyBd3m5Ln9tYzPeIO
JiyR34aDEMH4LLLQuCjgWq878rdk4o0VdQzTcy5zEHOtevtKyNL4XfP8w8IuYGpoB+cYW5PCU7aX
ZbAIbD1e2BNchXUUPYEKQlGYBGGxg7e+KoMfhZii0g+QycYh/LW4m/rsJxSoxtywcgNuINPyR8ye
dXZ9TMt+rQ6pHIyvbd8Ka60xuOMPXhdRXwYvFSfnsGdmaAa0yhgpFOXOasL5Y3jLqXcX9bWcRv+u
LY7dpX27BfkUIDxOk8epNWLiW6HVn0j6CjZfd9ERLAdOqPSlAZN6MbsiGwtH4StDX4WmWn9plFw9
XOliKIU7daEgo/JUqG0UlRsGXx+gOjNsCXocp9znf1735/QL3Qhk6JF3VCzuOQGeF4TEEt+MkKek
FzvslV9GDDwNwvXA20P/+/tolOhuzVabk8oODyHFcr5oiXGAISlvIMHZn6jrsL9DHO8eAO9RTT5Y
mqxtebTkwB3RJK6zedROqN9zD4aoYrQKYfbHswKMVtKViXbadChBVrMeMLoxlfIqRkeFtC3Y6+J5
MOeQ3fwXzeE5zd2wePFgEgfOfyIgVtO1vvQJFTRPOir2Rr9qxD4lHy17Nt+ZNrsfvfw9b2CwjV4Q
ENHGOW6qaCycIigqJitwrwgFV4Eow/RE4ZLlZTjcCtxErQcYNWRsvgoN60SmoyrIEhyO8pGxKS5b
HtGyAnPEJX4b7xmEhsnuBI4bbU92uDWTvmX+GrGcbPhLlDYQwRn0dss3NpUX/+8eZF4MysrhbZtY
ggDrv+d7ZDuyck6LEUZeoBdQP1a2mIZPYAodRpGF8LgFOkqXByce7ChoZDlAlLgCf3MjllaZL0S1
eXWJoT9NeyfN1GBDuKgOF6t+zIrpibuiOhT92LwPWtME37CXn/yPhTCSgfmtMnT/YQ4DkaWhg3gZ
TCKseHQT45dEi6SuoR+Ih3UFhe0hK3r5J+T4escvn6wKcxw/EP5TQKfvMI3fq/9DK7a8IOchQnKy
9sD7OyKQ6/K39oIt19k8clpkdbSmJqrtYeqA02wFRfo2Ml1H36hw4ogytj78vqvUNgXtDtCR/oXY
BVSkpmUl+BxHp5AZb5zEm/1NzhlyDdm9UoilRkwdNOiT2yLk4/HDeZHOIqNazMPqvuWNqPotzVaD
jjemNIB+lqV1dqXbNUWe4XcKl6Ymp0DIzv3NZyf3Gi136mbhTu1veqLfe08KgA2y+ZhUyRUgZE1E
xJjjy5FyLmPWvA/an3gsUv7tEe/IOx26tv1Eg07Ue8WgylqDVZzygDLx2msPUGXnVRfvt7pzmJGt
tvUcIWhryQESRTDHuLsmpW3x57PRsd/KhYuubI9KdyGCc15TzBnKq+bfnSzH2W2TID39z5qvGLk8
9IwsCMtl9i2vIjODIcHMWQ8QXA/T1wHi1ky4raCuLp9DBphK0sqjH85g4SJWJ54E7OHPtrYOyVxD
zrGQWBq5T7GnW0w1VcJZns/dRYd3/niEdIYiHeleJ4lE2/lY8oaha6Cd5fnJJtbHUeVZKXvUJc22
HCdXGeXzorDb3o3aP5j4l9uu0F6bUQCt6e5/Dd39IIU1nC/9NI/P6N51HuZMyqKDWD69xuBa5Uwr
lWkSvPQAZjTewY6EzxZUDgf6JSoa1Al7RBJlHrK1ialq66UmZiYpigfIGHD32suytgvsIXXFiQmZ
gKqk8IGZ+CFM8Kzm7egA6yMl/5MVTvlinF0KzicZzfeGRrFrC8nGvDWMuGPYcH3doX2gdfyh3cJj
N55OZeMAN7iuSx3sHUEg1hiNr8jR+PecWE3bZMAL6nmXQR8gH3bvRVgQnCD1rnJLa4IREw/mvMag
wTnxvq1+swEIgBj8NXj5CNOYwKTCW6BjWjoAoCrTy7SPZccBj9RWQ42iQwkrj+h0xfJJMW3Wng9G
MxM/A0BdX75vE5Q/b52fRjwG2F57ahTVwOiHfaYOYNvIhxDTMssDIyuHA9EDmlRXl9ZZhLVuW06H
5boljJGpPi3vAGm+XrFdOnNgDfj8Yx+w2JU9e/2F4Z66jrYbgqW77Nz7dR7zm6NLnVmr3BNXKRK8
LnsY/TMWyC41gIpuyOxYallKlifXVQvA7hwOZ60VekpBPD4MuUJ4yNy2fJqCLEGzboG0onO/pnS3
mPZv5cNwoTMam7dkQkcBuBv8JKLRJ3tn0GJfnh2QxIt8M9eEprUTExLG+9TvwPz/e5VZYz2g5psB
G2k4oePesfZD6LmmJsO46wZf/Yjmq/2/VEKR4rcioK4ftP3dsDUl8j6UmjuNrt0dme6BzQ3hA+p4
WUgVWh4HEDiXGYWcKxF3CalaHFEmTbzt6VNgzO/EHDQE9A7u16Qll7gm8AkTIPVFnx4b6cwR3HDX
mMsX6CtkQfsygxcIW8c3qq0PS5Lu8N0dgGjwtofNj7P3Ue3KjCZopaX0FySNJJEXh2p15vYl/w4d
Bnobcl3stt5zVo4g9bRGCEWvHlUGu5fHzPTetqb7p1AbvwTmKSZEeTW0HMCPqhoqsJDAoxVHj4um
97h757QB1PiyCDHeZacMf0wCVKOI9E284GnKIYTE6J/gf7GxXxqxoRN2gR0hjcXQFtSVXTI1VCSh
iib2H2ty19cbg7fied4zwmZd8fXKY6cbgRXTliwiswbxsZaRX93uNYqdrBuF+f7wMAIwo6UjSYm6
XybPGaMrdKnJ/uA9O2KmbL6zyXFP1wJo1tOacI/ReLeWvKuIiz8v79GriKrdlRl1ICgjuW+VWZo4
H5P61u/s/nPBN59zADSvyxDT5CC5YFQdYaNZ6nniThzJc2xlgftUE+nf4mGUAEn88cx7amUl88z+
IirodyHqsyIkKDDZHT7f0Ed5QLvFfPtbLL8Lh2EIgyzVnVCP14tW0pdufclNSkPXApWqefZRbpyF
ispO+WbS+6tOM4z0UAP41FVXVtdNM93VShnILDN92+znVW6ib5T4po/5x700jyQPlEqmB0vFpQoy
pxE03RFPBDo43SbFEFUzldf0AvvhLXu+uDl8AAJxetEVue1Dr7YINkmy1Zz7eOVFWcZSvd/X22Qd
y//tU5vB/3IizKlCSp0fObSNxntXwiyQV5QfqQYpwpa0Ax55lLTdR/WYbb6XHZS0tJgdcEdwS6la
VGyk9EHpKeA0mazRdWUwDXdR/Ev92qbs00eA4v16v76kCYo0E13JAzQxkY4R57xIj2Dj1Fjdqj1T
KWZ3bXbkffFUjQeT5lntSmi0xOrgWc8TFyzCXVv8X60gSajbOkIG+w8ZnW52ZDX6qlnJ7raCodoN
BdjaW3/3erbAhZDyS7aQj7U8BHkCSfZqyjAGybopzUeRDJAEZyfXRFVmTxZTAuMa2XtDcTjmTJT8
oIMdD23UOU/kvoQGPNlhn+OLsGG4cBdURUbkUbnEYmIvZ/AFy8yJ1V6zhPZAxAQqcZAZzzuMZ2ZC
NBDhUIiDHhpE3h8Iu85yEe3IZBWR8EiuyFgrC4+9CAgSxyKFntB2aM0SIrEFZ1tLfGUPPi9Lm+AE
E+JiQeEK9I7hdopdYYKSxqZkAF/uEC0MwoxmoKKIUgw4Bdb3+MewQQBFJekeI9M3VJQZLoMBDTFk
4HAFS/gYlDtbsw/vkbJbBG8JYqagPQN9rXCXJRJUxOk6rREGVfVqzGCRHl+8JTfGbrCq8b02vERh
mswg1IsoTwfncs/Qel2Mu32+LyZ9G/tyC4qm3iXEskcUN4raDFiSzz5t0vvEvRTQKREanGUI/oea
2ErHHCx0pT+5rlG1UsyRno+kaj1defz2DAvL45LgzgmSIHj+B9z6IkOtvZMKch3Gl/ywaiUoW0W2
8g7XcJ9IVftS9VfHwNV8gB9L8RY8PqV+9IOR2QV85UVB8D5j7c4fc9Mf2WR7+Z2D5QnrStR3Y4Od
Sc7tc6QtN6t1uOxxxPQD2GyYAUhndOZX9yMXjJgvR6nr5WgIwLLKkKtBCLXQmi/d22I3yxOpO8wg
KBuvs0ZJf9nflGH3UUh3PJpOuQxISgAE/adQdLnXNnpc2O6D80OywdSmc7AwkWDckLcDgPZlD7Ft
PyATJO5JcjCw9O99Ek7OBcG+eieCJb7Ghr2NCNiCy9lu+KhfDLptimU6CyQWXN8F4npryt8ZJpia
RKzhWqlgvyFtQtvniZYtfdm5v383SyDZqPZ0XRqYPiHaL6QXCU47qtBszGnSywLuDaDmvFqh0m/r
/kIJryGR2947ZgXD6Lf6oYxgGwgZQmTogI3bHbkqPwdVEJkZsBcJL/rWZ3yDIbX6R8AaLcFA/4VA
LM8pjgSMUgxBGdhydBLZMMeTk/9ko5zSCU38rWqTmMYZ/geJALkkH8RH4W+TvsaQOlf9O/wSp1iw
sY/vJEr2bvKKMWgm4ryvAKYWN7nZ3dXGBqglz16GDajpqdjPO8lzmkHAD4VJlY5sBJG9R1CUxCgt
bfzurCGkGrD9CC1b+YlDQCpdTWPp8/NMvcrfjeZO8W+Gr4HlZiku5QcuLV81xqH/BIpxAyIBA+wM
KOmFLxX3cYi3VqvuOH9BN0kuRJQEmgvSjCWXNsetubqwLJrm8bWeG/UquMexVS5i7XcJ889edrlH
XRGJRbPws6BR7l11IlbfUYFkehmG//Ft95gpZTrswYfeZ1xdmJP0lQ7Mj3SOl9ESV9bjUJ90luLn
+uDq+jewkR3H0ZFnULv2uB3KdWr/J0FwBWRzR6TB8oCWSTgoS5TyhcPDXI6K6AtvpXPwlt26SsBJ
2P62GIGaRSPJKWESuuuJPnIFRVBRusxwjPQnEIo9I3k6xKjaVrwxLCeFBdfWkga+d2FhqmkLiQOL
7rTafC2qOFtKyZdChT8U2BJyjz/ofyUYkpAwT+B8D3gzm76k2O4iPvWrtMfnoL4EvWMugtdf1bb7
2DEErRCrhDvctUZQ4+ssHYwKnNKWgCuoSJMZTaf9i1GG0ow15O1jTYjnRx36k5eDS2V0G1wvDbv3
FME2WTafEbDhAz2w2w6iPzpkhisVnB4HwDJRp2r0fVr7aX6hwWFb2DVoUTBzzX5uFBDaatUJQDpS
XaMrqp6tsaCVK2HpYOXPcRr+VjqBMtjQEx/vq7c3+7kx1BKsqJ5GRSgRB95MJF6ltS2xtO0q/Vyd
Xy7yKnCMRFHcqshf6qzpwSU+4B+vI/dkbeGU4Hexw2VHVjE6Yt1AiUX1CBJF2ZZl4k6YtHbpDFD8
lHT7/i74EoVBUJQ5cmIfjS685fyJonq050rDjk54imK76X7zUCX2ePrwgoiuziat69ME0BGMthKU
clmP50SsPBmQavtd8qBWxWLfjgGazdGvsTJTILTM10x7b/R7KRsL8zgpc0skvs6SYDMdhjxBJYW7
9+/dZzmFR79rVSsl8NqjFv5f4To8GZ3u/ga7FDRQ2WIN+I0ELRIKQmhy6m90HvVVvUuga5XNqlWp
n+MJWYZLjRkHuy2MTpZQWnoaMQLyFCUvC4K0psKSAT/CX/B7NBEcNH72bZklhiZ7EPa/0f3rvjFV
gQkSQnDmI320SIKH8mKhb+CnYAgWRyHpCIv7xT7ekKJ0mEZtMqPRRW7fPkrTxM/D6fy/jzDtoeZY
FD7wNKw2W5IC1fZ551l0YObv1n0o+BkC4xdwRTogtU7RaO6d4mwDxemDVkPrh0bfihmBZVjtwG2l
E4CaqgUt3+gfYLly1L2lObKcsmIMsRuIyJLy319EAPIw5IJj6WvSQZmzAkk4LlIB9TLMY6nOze9C
uUrTObYRmPf9PtDJuXxGzxKnY9aGKiisdeAltiPm3vu+oI2+mL84kmO0ueqkB06O3M/+d+gDKVXy
z5exq0fqYKHgEpa0V6KLoOIz5mx3rUXXGB3zXzt1W03h1/q9DXNUzeKuh0J3ZjJkPqVyZT3AR6nb
EbJwKcBJSFO5Y2G91li1dk2CQfl0HQ8eCfypPPcDZcFisSBcE3KSood8vgdeqAy60FSZbxWlDixD
Akx13osCpO/lrHmdP/eK2mzPe5m+BGU0gptPR9f+9L7ZyCBhoB2HWndQUhbjmetc4z51e0haBBYz
4wxKzH/SoqdAaOu2LKcZss0nLGsj1v+0XwumF4/OhtWTVaaXEHXS6Q7h1h0VmEqopctAHHIl0kDR
xO9DZ+G1kkL3Jf7P7CGIFN5y2BWir5O7um5Z2m3q2fvaUBQ67WgDED4RVc+VaA12YSnq7ibM3y7e
wo/FLGnnP/ZJxrfghw1MWSsDgO9lxYKsi4uGxluot6UozmVOf92Ft8UzS4YrBkCXz4stAtM/zm4R
edCEQ8acj8SJxnQKDfyHKv35u8/XuOdLn3t+TEOXugfy9UypF5JNMKL+KVbmbqyScUJivaUs9zlj
QKeMMGuatU5tfroWNoF6W/DeMUS9RPzRkjFm2mA2xc9xWRbRMwuQhBqn1fChpUxOvukNqLeoS/mx
ppTnOmV209bA1NptlpOQVC/GcWU7exRrd1fHNzEeBDIoPtXPoeB07Yz0K5KF1de8n9wk7ItqMamz
ozbO4pJRMyuIQINabYWgDGH/Ry0wesBUqm3mdKLLyNlWU/BdeJSta147hnBHaAoh3qyFsym9Iq+J
STBbPqHZyMWFoUiBhpGgnudCwDLKEAkIQup81m9Wfg2xUO0K656EHQsSGrYRQJcR/Fn38+CvM7e4
MdOr0tL9+8MlM9Kwck+bYFEQdOC6YAjHpMlRKEOEIe5moCiObCgcCxQD3eos/9yO+nVUbFNCALLK
OOHpLI9uL6VH4bI8x4OOmWowphumql+LTjCQoxLsJaTbYh/S+EXV4HV+NZxBs77TOy5ZK4Hu+hnZ
rSCzv+Q5wGgKmYHbjqgaCUIx96lQnDg8yxPMJXqsDyec3NdOnMck81IWyi2nLfNdZvuEeIms8+b8
jJC5Wq+9cTAyqyHIu6kzMzEa8U6VwNR0ZWtYqoyt7kK6ziNSADCmlsjiO71BDapx0bUKNZXVICf+
d7q86/DQJEYr2qak/5antpnZbQj/5tEjmHy1OlUjLsdjsBL4PLbnRvWaMudbpmcy09dI5tRopM4G
3ji3BrzTZHilp7p9bF36DkmufYg0sN/gd74Ou3Q0zLqE2ZZhwv6rFzPmY5uUNeBTkJZi4jf2JFAw
psoeqmE/ZmYV7tHjljwngMzF3ZKN45F4eUJTf/G/usltbE2G2YBukR/vvdVNtmosUYbjM21pWqjk
KHd6jE2mxnfhLlT+raqoFDMi4v+9GFDuBsUr6BLs6LnjXCJjeKUGogMcF7V3RjR+nQIxYIBF7zfk
JKnZZDW6fC9mH3/jMZMmgVFw6exDEik/KRXtc+KCbZKttxcR5aa8UW11YPUh2sEamN0DCA+CSr4X
X+auRKDEFtb7hvN3Xf6QNb11FYEoxN0QoUw51AMvKgKKvN1QSXuA6fokGMtxNhcJ4KXGjIpgha36
xuGaJYEXXNZEyNuSVa4goJvs2Tyw1lsAwO8Y8SDME0cCfAvCEpN+E/2uZloT33ttMuA7hE8kpYtm
ChC29jWuyl2q8/VVwy5a6APnTd/S/TCSXftLIA7gsSBeCUhX99/Cu+AtupnCj6LIaOTDOV7PtX7g
Gc/fM57KG2fJRkRFMtGNRtoa70UnYzzWLMU/LZHTrcVRE67O+cprO7rvxl8vD+KKPqwlXZbWmSFB
kGLWq6Gxrqmsi9tc0ZGtalhnD1lwTl/3fhPDoHjm77hYxCp4KYZVh8wlcaFi1pKf2VdqO4i3lUaW
JRxajtVESgss0gxVhfRbQ/jqLJ8szdSQ5Ques4Bl0OXBl20FXTJQwxEmWmmmNc3DOxCMwUMtp3za
w87EEu8cM3KUo37hcb05BypHbXt+IIp/Y0+8Q8s3Yjm330VYQJkn39ZTmgtHlQ+WwZvAan/I9qAx
lAxzn35xOa2HGrBd9JVALrs9tZ54oVbnzv0eqYRvEE0TYRv882eoLPpwNh+o6BXK3XamN2eOSw17
UeQXIeMmTJDyvgoUGNfzn9Ol+rT4iZBwvpVJ21PMfIbYUPOQcWrhA0LxpbvXmYazld8aiXWcgT4t
0pYXq140S9zXzBl1gx497U+0Zk6P9VPL3ZDjIFkXs51q5ptd8fSI4cORO8sttEe6XYZHq0Rl5hxi
RGwPJkx2dmYeLNomIPKYtJyVwjK9TgibQqfEuN1OUez4z5uIDkSgH36x6mg4PiXxJRh6HkSrHg8L
DD1KSNBekAk5QHWaMdoObFNLIedvfhAx5R7D0xtnB7UAovSXt55Ez8ypFx+jVyQRzisHfojWJ4kG
0FoofaocANajmiFdzzR/F7YapRttNwM4oIqH0617Ew4jFYTvW6L/Ni5hSU7gPO86unPu5iNestS8
gucZUHSS5bgJoZZpiGukRP6Rn7uhbPyu351ZE6c9zYeva5SFl1eTmXTFqO4VOxx0v2kP9x0FeQ0u
/wkWJbc2FVry4hkB15/PYFCAACqvZzjezMDgOFQFyd+3x8+ezCE2YP72tRb/IcXk50myu53v4fLc
wmbHjr453wuBqwEOcnMQ3xEbb2xDnqyI/ItQE3tNlD0ehkmA2IQCtFQzl8sxyg0dd3s4Syk1iVEe
E7racbWUCkBtyiBzkhSS2tpBfGD1ZiqR7Gr0ofqvbVop+kFx2WOFCANZpgXV2TqyAl430k2LAAKy
auddW1UpF4B+qGal7QPCuq41HmqDsQYfJjh8Oijyqa0p27cbLWTRxB8V3B6S2BTSzaJYZRlIxanY
8AYt2hv7hWZ2zN9AQhYaD/cxekHSJ8IIVGirDFcRCJ0oMRzv0TZiu07bdFFFM9vRFRRIuYxjTdUf
hZF5IJaLHtyAhYqZqyGeZkEey3HzGphALCPgM61YpktZM64d8ROxTR1IkWfyJS/yArq89LL4jddE
b3vhRFN1YCe95Yy4GI2D39ruY6wq1jvaWONiLQMNuyxayorvJ1ddyv9veqko6JwVfsz57Lcg5u8x
v8y5/26RnP0c+ozVUCly92SBDsKyFqTTOox6+09xnlJQH1rpirgaf2wOzKaGRWXzHI8lUfmBDTkN
48mjwD9aPG/Et5WodDDeu67TGhUO5Oz9MTFjJu9QkgOW397FlgUcPYCloT+xUnfNyGS66g8xqkAH
4+wgyLMqDR+sarPD6T2S3h+1mSRyD+AL2St55jqJKwq5vfVjgsW888Mbugud4qPp/m2SbRd8CeOP
Gw5xUVkx2pLGTPS4PcCwxA1GZ8BrEjGnWmkH77dPghuOqKAbu+NWgg/QPsAeg8tYFJZtw0LfbtbS
c4xCjjKIrplaHZE0Fmv8+ZNENkb1bMoiox1aMFEZWaZsh6tBoQVos/vaniVWc7k7lhXbeKi3yJmb
fPiQICqf8B1yre6307xkH7q1rdA5w16xY/boU9aa5AGANLrNirS0XltD0cbeYP5btQ/8cqBOao+W
zEkuh/DaLsuDx1+k9HgbePkmz/MFr6eTFmztgp6dEyJG3vbAZL9ZCNJHed5hNfNg8SpkN6TAaF6M
f+LUZjBCS8PN6X41u3GrJumxekF15lnPSsL8JFxUY0a7bD9bCYFoL+D/mc/wxCdMSIbnr4h2rZWU
8Njt/as6MsbPn0XYAFXGsC4aoFLNj+mDft8+f+fQDFYgNuWq4I1azFTWfPGrfDaj36oKpEZReFlR
ytIdfJmz+TDYu6XRGQ8q73cZ+uy/g/BUXIRANqc+FgveeK+iSsBtsGWd3/4hCunNGjY9SWU7f6TT
NC2j6/q5kXqHgo5g6qcHo1QzAPNpfprjabBF9L/UrWI7hEUHaCrz12bcbVifq/jofJq9t/FZzrL2
nd/l7kGS0bFW5hK+Bd5amxZGD7BQCVgLBv5MYu8XRnH3df1bvYxkCHq9QMG4w54nYJngwGCKIdU2
y9fzWq3fqnOZwWNQb3zQ2LLessnnNo9DmGxMgJdZldSpXioCG3/XAQXQMxvW7kQMZ4LBGTNfh5Rh
GHsJIuuJfSZSkboqGKjPjwK+VaGhqxXO5FbbHzZm89CMWaH1+tXKzpBG1qTxxkwgxgiz+YJkp2QI
MAJO58jwHUAxCCMf4K32Mg+dbVLph83HyMCRt6PBnHkY+uwnL3Dp1L/uJ5mkoLCLdQ3alcGWqPIX
IJI6boMcN1Uhq+QKTxZX6VAoUYKTJx+x6ssTLe/2DhJMLeBgAjFGBfo9HvT1SVQ8+wiNFMLwl9tG
mY2zH3tHGVdAxgksI9dNenGE8DqzI6GS3/M9KF4SRbaCO0D8DAZyXNSnccg+g0Vhsov92CZEhLt9
d7y9f+QpqqxABa5pWf6stMduUvd1eC3UZcMTp9Wu0TUNMqZLsdj8RD0fyw+kR8tjhiR6uu/R3C6J
WUpj/I/fxGVvPAyF6TjzGCG4s9GL+FhBhJMfdgLRZAphTATiHPxQKMD/gdGVTPurkoEfTLUQIRXE
Y5tQmS9lLX087R8rwLwuwLrziBk+P4W4zQztIH7v/1+LgUmXR1Adhg7FRmCTzuZlX+Bn+Lexb5+8
Mp33D4co7+eSr4jLWlN8SC1vT8b6N0KW5IFvjhRJ9QL09ELRqSkrWsyEjx4Cfn5FHVcicKfprB6i
84NhSQx4SZJKjVbnAZrY3vxtIWduSkWis1PrjA9Wy7nGUbbclH8wluJK0VF9yo846UDKSA6Ht2ud
ULlMPY17IvU2+GJWQE+NYDOI8hEFfeMbyfWZL3D/X7DTvgMNgnphMNvwpWreiFnI5BN3Hj0RDZR0
Icm5Z6THg9w5MFUI7PtpMxpzV1rYtkBCOg7h6bUvv39MdskBWPG3rbsEk6fap8BvMTUKIBM9FSZW
rk5gC2mU2OuqW7oXaM2CcGwhoybDDED0dCEgQ603XesoZ5CafN+IHoXUvtFCtJkMiB9ipN9qiyGA
kNKET4V7/25NOMdrIIv2muHWVSX9h0jtEAYoBJXTxZ2/QnWbGwEbNEnHwkeD0oIUZ/Aj6KWEqDuC
EaCFRVQvkBlJwxzFwkPlR1mcSNHNKbVq59JqHtkCkSygaMN5bFqXKvdCW5XoDAxrl+FsoXq1rtbK
OZ0rzLZrwb/Zl4JAFdB4n7OTb/KaxXsr1WClman28jnbZV8UuDlNIaTdc9CXhGlcPH3/aJj1jzbf
8wD5EJ7Bsjlkr4MXEQYzWSrKJK08P329knSRDcOY7nuTBJzntnm1zVTpdh6dSFlZw0S8cf8gFqrM
/tjPAbjjhBYoEyhQ9n5lOATTIv29GOtw/0nZUcbg0VHBkUqRntLK393mOHaVX6peyYTMdRqvQ8qD
9vXDJhualeLFjgJ4nWyVmnrj0fz4I9M8plp9VyZig3f7Z6qahIt0vdb3mvEuqx78FRylL1tfW289
MmkSfRtCZAviRf6H0xpIsmy1zjPHIu6Ho6sq1msOb/z2LOWCoMnwmT6V+TLCBPbOCvY+TZIUFxy/
I83z7a4iwuQjIoqWmzA6uROFx1TgvE17IpbqCu740BUxl81aYyypaa30zV454ztFZ8Z4lv0gAFo6
ovuk4+ZVibcuPpncVUomqRPeoNtT1i5qvOgwhA6uZgmlaY28bKX1qZCUyvuInHzGlwfR1Fh1bTCl
2qOlKYNKLWvT0VFAZ00aBnA8A2O4EWjARFYG+vILKVTmC5ZcNes26EKiTWXHfFRJGkdWFXHTkowN
FMvZDY6LraaCdjdh8vDCsxrlQ5yrja/ycoCjFoUbCc8QVv8T4n9yMHas+JOygP9dPo3L+90/08Nr
YE6G82pC7F2iRD8kefAaOyXcGNoO9weAaBJuWfhIxrs/TXi71JnvxlzFY7iozeovgrL7CfnWKIvP
RiV+kvZqIQ9c2e158edGR/q6UUhBwmxt+eBv+fMCWHZ+Y+ASVJxHYgOZwm/8lHu00VHWjpzJ6HmI
8/o4x8V/PkYFqmArNOKwNL0WBlIP9es69L8Gza6uJ3Vtlj0npPugIq3+XNyhVcV4mdHCUppbmBqT
7YGn3CT/qWbIYv3izq4vVqUP7HDeOj/KoDOp8aQfIEuWjFQJWynQPHszu8GGjI6S4QlpL8Oy+Azk
EccMzUfAw9JXiZK/rxcV+/S8V4CVWFVjr5Ht5g9wU2HjsBvgpFnrzkfX7737j3U9gFWDEKdScdpj
rjlR3xkEpMISvKWpu5xNOC0wbqrh+x1wGjtBNN2XHlaKnOUx6HZt6zydQun+UyhH8E7NjyVcFNpq
hh+WPV9w/UgS7DdlAgjl1QNhTwlX3lr4t+r2vO+hRHPRKKrwU0tmN4MpafY3feIOzKoj1d8bNWfc
URIgPWoJLZMkoRmh+VQP1b5OaVWHJc7fbE1oBGH84IAFygkeArNVis5kuV+RHWT2raEvyGb2AUdN
QN8nOryWr1siykf/L0urhhMsoHc3sWnhJSKuwUq2/i03EX/flo/e4byIxr/LLD5SaTXiWC0Xf/dW
ZX5sgkONHsMk1JJBQwzzH0jE+VmY6HH8lQ4BgVvJZpkPgbUn5xdAqSnjr5xe1fNdyjlhliIitbnJ
ZnDj69lMNj23rk2uFCwbf2SfoWWhEW5VHP/AWqN+Yg9NjejvHh967IEbN/0s2q2IBRgH2c1CCb1q
U14m+Dk23JYrYI0xIqRgICAFvri5OMoK7NmDkn9Xu2EXSpzGY6TNr+WYVG7oPa/w0x8hxWcJqC85
7E3lr8/vRju/QpF0vXNv9wTm/u2quKStZMA6WovuK35DWfOLN4PK4SOSlMr23oPOENNpoDyOpBlJ
q8palRAHeMOY3c/KykI/H6ewv6aP/hutIDTLteRnJe26abnpbR/pob3dVYvRzWovoQnycvAJC1ut
pYN2f9dsReoUqrU3Utljwn+iZfacQwlKWJxb9xTXuXxIyEVSeKRMnWccqarpAPrp3obUOBSv5K0U
cmOTj+HZett03KviyeZoy7GAn7XlkBj0060YLRDPNAtIixl+NkW1LCgy2fShWmW4N/SsVk+0RV8I
tj6qiTusOHEoGY4KmnGDPEwUoxyeIUBaqZsiAj9k/+ZZlYIWLL9xZgYZz/vlDPvxwjLBgnoezAvN
XyV5LzVzkfaFUXYlvvKAKnzDLl9HMFQCjS5eiQo1PlXjOmi09vPJi05YZQXtSmZ5qKoRemg3csgG
8sD3gIzMyD/r92X3V3QOkRYvP2RzH0j6+Y8149SszefY/l50WlFXlR2kC0m83V9S9kmntC3NefLs
IgQ6XT4p92sSItImPj/SIF2QPwYyyqoAbuQjQQy9oz9T36D5UpDXr+R5re6EKNbm3RQr0RgjgeFI
9iPEP8LKmzkZbJFMduh1GZtUiVCrvmhCTt24axdd5yShe+aG6uo0E+c9KgGdklk0ZD//QbvlCQ+3
v4CzuUyg1A7I8tWxBEmAFNpimC5JffOcqY8O0H5PoHnAwmHvQ5pgGDBgNp+FVw1/tQI5jiZ6p5Xw
ZAjjD8j2L1Clze22QjHkj88npuMkbwIk9VImUH0VATf3sxZSeV3CU2/5o8XnSBCCky3119QdcWjV
iv5piPHtPb+uvTAXrbyqkN9Uq3DcSCuTJq4bVKZqik+CC8oS6Ev1q0TUXjGIZcmjk0/IFehIuQx+
pmQTC9eT35p0z38Cw6+mIV4xIpd19JvmxEQVDzO1LTbTDfN8VFY+QAfG7xfOKIdY3GIj6f9YyJ1e
j5EAHpDMSwXMv5gtFfwheZhCQRg7ojY0IOIimb4vXPmDJfenmg6W0grmzdQoDDcZNYJn5sDU/SOo
5M2LdkyBMeyjXqqaVaenT947qsQW3PDLBb+j7pKA9/ODoyOH+PA3nKlkCJI/LRvWQ285Zj8irAfr
1th6yZcYayoikf8veYSZ3ivc2eWgNeHQp6YsMZQJcOtA0XMCj0e49xOnyxerEhQR5ivWA1YrVnTi
qN3FS1LRRttVGp1K3pBhAW83b3qh2xtII9H5TjsoghvldRvwxAIcPalL54wICVRGgk5+HVR+eHKf
mmVWyTkKMPmgFTMoBhzV7esI5gTkiD1UMH/9sSG5XAoZmWAsXDAVp9ddmbMWg5jdQsiYv4to9BEH
Krrzsz7UTRqMomjOzeiJUwmqtpneI5KcttdXO2EEEJn/L5yEEtRMXcLqJDMc1Y+qhf9o+Juj7ZPJ
6WL3zwIGq58PdomVQnpnsfI97k9WAV15i7tiloFT5GgZGTnkplzG2A4dedwv6FBsgPfNduq+QCP3
ai1CnftfHZxQZdQNYJbJkkTgcWQQXi91nJ70t2kzdY7mQmq3k3EPzKYSIk4F/zLHKgMTC88CMej/
qwpy5lPbZA+fzs7GCHLM1bK71eQGz2druP5DqtIG/iOOSuypKUg7Tq17LhOoHBC3Oq7zTHDmk6+9
LEjEVDxMTLOKdJ6txxU+QR6sUsh/PeB1MVWdYGYokKxpGqjZ/NKxR4+pGyLWyi/R3n3eMPiWZd/J
5pxWoH7UEjKLj1+N+jTWgMGulC9HEZeR1cGG5piU9+6QiMSIxWARtKU4pKPIQu5qiiJF9B5b+7ka
ZXNaaTMvW7vD0dnppKJe3hrOdq0w5ySrB/T5e7yqby0jrciAPivzyIncJxtDDdNBL2hFGYXPFf5S
6PmL8gxxj75B6TPqYhCqx5yU6I/w0SQb6R/BnG4tLYApkMe0vNCtaPSFOsSqKEosJm+60F/jKyn5
L+1yhp7KwYmSxhdFBNXaRwa2qB5WUoEqeQDo05RMMIlfW4q524tnBr8rhaYQJdTm+uCDEAllQxDp
Cz15KSa0HJ5lRJkUVNAlLEqE+FZOk1IVhxfgb3qei3FzoR/699gWtm5BBtFwoQwxlmxhS3D7lGPJ
jO6yMcM3GPK98CFf2a9G7nOR2n7jLGRaP6NgessijuPIaQ5ZZ4kC6UpIkR1wm9NC36WXfZ6aotHF
daw7qGvJ2cIoWJGnR+gk9ADJJs9TuyKIeIthqIvNZ72VmuBqFIRwmREbXXVrwb+XNDu9OW9T2mPf
VYj+6hhGxanPj082Fb6FwqciWNz5JwtPRl6YktWOlofoy369B7BI3TIVb12X89FOxgvqW04NiOOl
3tyfD0BO+lcJmBc4JdJSSQfWI4SKoLr6w2FkfoMFeNN9vsx7004uPmHVEY+J5XJngqNMd+STkk/v
uZcujEMnAWqoBhgG75hfhubqVExoLO60l9n4XAKG4//7Y3KQPO9f96mqg5o1gwyPFY0gtiuSou2D
7g/U/PGHUMPDwU5IF7F7fdycsoDcnXG9Vh7zane96VjC8F7pY3UfGNjGA5uZRK5WEG/krDo2EQpD
qoOpdJ62JzPtIEMBZv5T5kQiqWytaTytGzdTL4IvSr1tLQS6l0eECv7M17KjUgjCAXCcJeJU20cS
0G2DX720WhnS/VbzpvihkdCr7WMJnGlKvRtdWc8TRwxv3/C2Oh7zqtTAbvBK32xDc0+vvoqHPWfm
4aGQmvAUqweGWXrRUHbEa+UdTAno+rDd9Vi1VerxsJ5eOBXrA0YoO9R9g5fI37pCBaiyqzRnwZTx
rBOTr4wM+zartu1uZSNWWIZSDVf1XTu/185NHS+fW5ZqCSNIdGEfd9mTwggw3NnVR60moG30DgOS
U5nJ+IsYi47n2VrpgGmnBRi3renU5DC85kCH2LXf0Gmfdjeg2RkylNjWvO/7FtNcVZ5lXTD5buCm
Rd6cEj98m/8aG9iCY+xWLIjpNuTMZi59nrZNGxkX53R8uBVRdSg2hW+GAAI64ypJrcXBZ7OqjmFi
0sjsmlIoD80QMnVOSmGDMcuSYX1TtxeMZHBYH4Y8RFA9ltCvd9lrzAi6882TB02yBI8d1nbV/3pd
+XptNW7GRh0vZNn4bZtjin5c2ILPXwKGiwwz2MUJNs6JyA20Y1Vsbbzcf9xqp5fXoVeEZgyC95ZR
ZxB7c4qnqotnn1QWRkQJOTaKkrwqRuZf9ZNPp0WTL0S+6gbDCot4E4CoUfX3dD4wJZItP079sdSw
E+I19v74FhkNJuTmRyEBmOTuQY5QY7ympuF47DYvXcF9Bcj4wgmOresYbK6Kup7YESN0rNqeaHkP
heut30B7gUgFkaJr+swDH+P6tWZqQJGMucsoaUelXzFV/DA4iSFO18pcBXXlu0HGDKTL50vrzdFm
qDtNfQXy6gJZnTlT/FrpbcJJJxnkcmWnT0W6In+oYbr5OuFi6ABgEcqU33MgRWdqu4WRboaJ7sTI
EaqIHjmeSNtfFGJX28YjDV/R94hcWERNBAKNFrHaq3GJBsF+7BfZyIEdn+BsG8GXDKP0gdUcMNWq
fr3wGlmuITMaV+CM08yfhtyPcLkUq2wccSM275X9V3H9CdWTfvnGS8DKFaJ0Bg/MnkMjQVc/+5ED
sZ4jEK7CxNq+lZ5Vdmz7KmVZl4rh++nCXckBMmf4DOG2HADWpzJSGludiHXsQ/Z2wiOqsRkcAvLN
tsRr6UPaQ5v3J8iJq5D4k15i4YJGDk5uegL8T27SM83utpw6O4U6CyiCsWWq+GwJvcz5z3eDsJkx
Q07es55sjcy+HCAfBrUhESx+5JC8lE/pr1CQ30P7Zo6tnVlhJGu7JSdMijg803pyQRgW9kcYGxRK
TUxpHIelTsaZWDIMLZ0GI4Tz9KmMqI7gc1ee9oQSuRvnA2FwLFCmIRyLzMOYCMjZbxYfux+dsOk1
TZnfYNQAxMAEwk3442j89iPs3pKJ3f/UOWRIvFMpmb5D8Tsm8g2THHyTNkv7lZB9Zj5ALxFUWRUv
1KEMsJ4XhhTgPUTbSIj9sNwHoX66CRy8tAVu9mDSa/Bc3s9MtnGq7XY3PwRer9mKfHzCqUy4b/7Z
Kic4XTP89A1A0ia3uQ4Q5T5aInnbr6L19QayflULY58gQBb7finCfGi3wm+gXubL2+jx7UVSa+AW
hTrmift//rlHfVB14XrtPcaZ80mXLsanVS9XcIpei60am7wkDf6u5/Oia4oW/tC0Ki6RbI3hU0/r
OsZW55tTBdsY/7sJEZJFth+kur3rAKKPxnM4WuFFsMr5MlgsPkkxclah19oqr/Ffi4OjZvadcRkD
ehipUu9IhcLjLsyBlWJVq5wiHFfOjlSL0JKcMRfRL7+2YPGhHdDX3/PdBE6d16D4A6v+lpkHt5sQ
g2LKp0URqK1OxZEQ2o+fD9ghUa3jAnDBBKQljEQIMbPETMP+DIaGuhfN4G71o0LauBKBKlWkeXdM
kuhW0vN3fqrRDBTBEyiL3QUquAcgrpN1k2/SdU4aG7nTaF4N7gb+jS5LodnqIiP7tdfd71ACDEl2
QfJC0LEcR3c4vqwrE4HrTOAfvjtIoU6DLE24A56beKOox2bSBLJrtY+qP50A/hDscz0PbcUZMxeb
nJUvXb+flqouzjx4Tl2jK27eDJPD6S3Fj9mcMejoHyBR62lRzR9EamZGAeAxEDqfpnT7VA6GW4F7
td60mW0WnMqaXY2uzorxMioxBNihnrWUkhcP1H6FyTnyRmKRFz6Pzmwj+5a3lsfv4s0caNsn7iM7
N+0WpsWVimZggefRF19DRODzM9p69lEmIxTs8dnPnfsgeXlV6uUAlc/RcyobQx2S6Xke3fyLuwyN
r174HxEQG2VTQUH95zrKESvKxEgdaPf8ALfTBql6CmTkU8J33wdQp9kaWJDJ7noCGHxeujMy5/MI
mmeDjey9QxKIOgnEGQ5Lv3vsGWcSZYxviBrVK0kIYwidZUaxbIg70YEttgMnjCp6wnlWvb032YOf
0I2vD8MtR+p4EF149o/b4F684w2yDCT+DHgzkD7mqzAvqbK0d1iG1oMcfUJHRxqW5hJ2uuifZdcC
c7D5Tk7Vfu8stIw8dToq6VeS6cDRppq8rapKLPpIoKvo54N0jK0VFHURMVTH/Yc4m3++dAMIFSaV
Ha0pjeN0rhdCc/h2hlVUVpEgpiBlr3gfv4ixdBWYqYJayX1Hxl9UTkCfYl+OgWdwur4JSKWrVR3B
/sA8+DsHbefz4jf08Ids4wc/6BAWmX5gZ+8wV4DAitUGh7v1IxC2AmhEIiUuBuiM4qGLDuxBozoE
c6ElubxKco4NCAQngBbP6l6oTNzVG3VSEq3eyA7tX4/qH6K9t2RJ3vi40UAfin/YSlm/ggkowP+R
egnMwNivWPh6XMoYMrmWkVq5AYcMgUk7nL3XGakZn+BpIjMjfs8P/blL6UDt09CRsBhpCiXyi8u8
wvkk1oQrjnEbzqZIENS7KmNqNHO43424m1HdoS4WmJiW0cAftI0KN7fqKIayru1koTiypPwixaTV
3TdiQ9XBVj5QnEqvwj2JwI99KnlZP0IPSXing9qa3K+KBafj0BQzfKX3jVx8wxJOiY6Y+JzOOrTZ
KI/Yg8wbYzDaXQA1o3INcp7PzQdqAnu+mWHp4h1/H1xgMgP4UaBw+Rvm2dcQ6eE6XslQ8uCp2grj
7xinChrulTET9dNzVbLyrdK485KpF3yu0fJPZzeT09DabR9/7fiEITuuN8ViFCdiaLGSOoG61sXh
nzD7yqqOW+dPawHpc6cXsgurjalpl2P5y3iodmv+bZ8meihsSSHkCbjlqLXp65EuZH6vugj8twE1
WjBCYD6F4fQcFqdA0EjdOAmgRDPP72oWa24gv5G9VdQ6UcvFA9wfhbGKIVSVu37GqhviMUx5ZALa
sT1374B5rfYGYVjs3RIHlgRumHXCAJ2lyc9FT5Wc8y1SSs8jihbG3xCu/5+5n6Ip0o9fTCt7ql38
URTS095oPZi6rfcTTFCoeooxAPznvatUNsjnB3XvueiIaxRea2ZMvrmiqJi0BlK2hAW/RocIbkif
9sWfhIORclWqm1A2kAweDkqdLi0eDI2pMWxn+8mraKN+heuQRSbgm/mufEa/qYzmzS+LYpoeOFVv
/WACbgzXxyAj4HJaoNXJEtgeOf16MW+/6PF9haHaFSlLfgtumPx78o9DKSR6JOEW3leJ90K7TvzC
VTu5wsBp+wUrbcDEstvyGOFJQMGZXPCn83EUKBj8fAb99Al7fvKGx3GqVRVc5MHyg8lfufednvZQ
Bl02MiEE6RWke9Wd7SFakKIPDONsiL2WuosoKXZpyxRZMa2UaeskVndKJ1OdW3kPoLpgUcE7zeQa
bH20Un8hm8gbfoFxVrJsDH94bYuIp2Y9LbeoxgPuGbW7oWn6Y2AgIEXWZFz1jCXcHuii0B3+tCIy
P0WiiJ39qUc6GgeoZru47nGS8/7vnALpUwkw/sQ8wLjpQcM+LlMm1L94HoRzXC76RAlGzw1UHq3A
d2d5gbLQwJ8pY5YWqhw/9aZBptCFk6WoA9lRqW6S12dD578Biv+yBTde7eG77W9NEGJE8eA+OacR
7BDv8BD8fHnR0ekKBwXajeu3RMcpw4VFQiqY2W7iObC36cVJmauk30DW14mnWSIB+CvNRab4Hf20
C3xIgGeBrrADoE8YiLABKkTZXz2BY0pH+CXl8hr9hvF5Xy/kurl5Sb/dFAw85TggSksoC6M6bPGz
ExRIlwenl+D7TO+YKVf9uuChA+vhb3JWF8HxHe3i3/0qpGKZRL3rACnmjmCSICA+bpgXc90rRf++
5G6UYiRG1jeTo8kTqR2WN+8uQ2F7/iFHlQ8ccnbMabw1XOF+dRNX86uo+9erPbPWRFKpaUgV5Qe5
U2o8L+y2I6SsmtZAsjlucncftS/ll4BoAPhM8ydbbsQmVDMbnEN3PsvRTb785XbB9XIpYCqHtUU0
djrVi6NMF32PGMDPOW5DA9uRu+x1FdgVO/TMQW0S1oGmzG30blQAYMtMxy204SXKvEz99HvDSaFZ
PhDc2r9V8OG6tza5mlyfk/f79OrWRr7sI+xk1qRuhYtzqkx4zsG/pT75bdZKbSnkEwUkGVS+5o7l
nCZNiGKALaUIc7WCrTYIk1Yh7ITkic8PJw8OOL4haxST1C/CKSUP+BwWwjSjnZACIpeU/OwKPOd9
IYgHEEEFPDqRLlrF0OsGVMJj5sjHzX3s3j9tIXhlOl2OE/T7B5JqpcOvJpeQRR3ysJ+o1h0S0z0V
7q6XZ+El4/xQ4erQo9tlZ8Jsh/bAC7QqUCbStqKTDT30ooO0ypAhht4Kyo9m6FME/IskRiepjOBN
eZls0ju5EKkselpC1w6/PQt8hj00T36aFJdbLht25KQz/1dKbm9i9JnKZbdKxljgjg5J74Cd1qg9
yiActSx8QEMq+VKUR6Z9MwVrImPmyn/ZOqCMjJSriN6lJInkyGw4DR3BR55iiGdXPTHid2glPh1y
SF82rS8TtCo8CRokSN1cqcQjsN0anLHlxkjFvax8ILC48whF8ZZEI7y4zLWZstUBvmn5A+2pKV2C
/Btx9ZPoAaLhRamDY5tc8ei3sI4Hoc0NQHezKjadAS13jItwE2K/NGJlQpAkCVr+f3lQQicuROyb
mx3WqLzdlJAOOWZ2idBjZ/bjgAd6TtQJRC9n9jvyjWWHd3wqyhKHPybwCggipffBZPged4VVaHug
5Lkgb3sNaKq4ThIER0VJ45mM5f9XVW4S721eJXMd9jLD5nX3TqhG4kY7yJlV2XQbD72JFyVvRKGu
NvSS1Bn4goVA4k0j4Q8LbBicTGjSdqDrbHac+/i9tFroDGuk1JlyPznpmFD/IFDzHRfKgDA8vLW/
sUA5cCpxebult5u/XBEtRki399Vu+BYaaO2Kdbr1HYtGtIMEJzMs3PMygYAss0IU9IgENXHfJXrg
itgRhaTyZ5kdBOTJfdgqPm6fVlHu3TRM46hf5njFAEybFcfqDh5MVlZ1WwjdrArjhyU2FZ1vP5u+
MXlOQi4KQCX20W3m/snjnHe/AN2VnsLJE1TbXY6B1K/ejHTF7yWPK5wNxbPjQgKEkdqzj7QbX0j2
6E8r7dw3TMqOGDiuRhViCm3smk04DorH0tnpdK7l1l/u9BsZL/GNjhEtZxYUbIBINil77ELUmKTn
xCHvpc65BzQd8IFvEnIqjFekIBEOsVjySvYudZOEcT2sDSu+7zf1b5KaHM9YV0cXzA88m/kI5Fl5
fbUOJThTqrsABgCYm5IHu++E5W0VNwSA+cXDFrDxVhJhSM8u/Ye876jKhBmRkzXudwSyzpa9B3X5
KklvJY1ZRYBTuL+oe1tPR4TpxrLjUxQAyjXNTSLdDZlX/K3u9WLvub8Dz4pa6zm105DdVfp5k3B0
cORiEGdEJjurL6xpVAmLf47s4SNKMGkcwluAo7bTG9kMf696WJ1mSlFgj/mIQvzsDLCQESTXmD98
YjCNKdeD/Rn8/LrnPszZsGz0MfvaW4kdsuAuW6aOH/QAhkkUoeP/wk7114AOM2hfdkGHkrHnz1zf
+DmVgHu71ypmTnk68n5u/UlXgWRfVlS2lYqUlB7ma9/fmGOFlOYDlfnNPSfNn8fMAar77bhghJ6b
Nuqr/kNgtdok67NK67hW/WNbok2ZsUHw3d60cpF3QuF4sPCH6LyyQ/pbT8vGGZGT/jz/sF+GfChM
Ym+xMGtzT99ogOPPhvqnBJPmxeza2J397Rk3htdmEX2lH/g3rNWKpAsoHQrnjcUfndjW/eJx2IjH
kWHNq/cuw9xPdv4f+2Akm3qdx4Z11th03rgSYYrfhVpbmxuSxvbi6DVjr+7fErsgi2P8qKWZt2Pe
TGGgWsfWdIJ8vHsVL9vChs2c5apEKaO7b0sF2VfPDgDlXowOVs62hqJGb5typgMbJRYSYktpMkQ+
1SoM8DVFP4/eNwVXT+agwCg+G7/Bto5xsNNYrTWMTYNEskOi5cXNra1/Vd8tyS+xtVgcWHWMq7hL
MAvmZfFfpiAj15DtFLCShhYcqIYKY0mYDBSZYqNl8M6MVFQOdBnY7QdNSK8yLUGrpT3rAkVvNC+R
SwtsfAbilu59Sh3tNpI4q6j91Cimsfk8tR9tG3rKwL9W8ZMwzNh4z1rJC+Dwk1v9Gxjab4eUqhGR
J9ISEt1R3r2PTuzkU2CXhR1uM/6n44vALQD+6xAjHqmMEgtPE10ziB4gyoyGrP819zEvZUk9Gd4z
APe31VjJcYzSH8QOPjMMWimXCn2hY9/sDrcrZBzmuNjO9MxgCOUi4Xp+Qdtz+ZTIW1O0D+h0CcYg
N6GpDHXxINx7xe5msiDO0AJ+jTvTjk13fthRmZgZ7sBAbANVTUwcltDzsKx95lsc/eO+sCE0ukKH
LXHobn4dsSvqnEW/yhxzjhw8Zag3R/87IZh0C0q6iG499IXi0KUAvNIt93Ryu71/tGtkx0PVFp5S
bQmJPtizomfyuVB+kOQlK+2pjIHc1bV65sbxXQGJwGMkP9LfHW8gCay1K1D3adu5Jnmeye1/2yn1
5Sma2ZKrHELGofIaYOD1uCUMxoHldVQMXFN9ptF593Toe3CrJlfYadzRv59HIN2x4gVuOP79pchi
HPUQ+XjdwA65o8tRUzsHerDeEfTNkfOtdGGxbfmdYG/NW5RRs2SabNmnhzVSWBk2iIiBrjcakoOd
BJICjGvGo4q58p10NzXThBZ2awBdjv2wLsqsc4YUv1d2OGkGrfQSx42w7C9S0VejDG0bPJSX4+Mo
PQ/fVuX/9roRN3tZ946RGyShh63aO31FyEtfeghRNYPvXAlfEOrJhLRwQl2wrOtxAc6VRmoToDiC
y4Htctb8CMPIUAOaBp9IDyrlXisog6rdkMt0ZAtkvnL4qp9yry+lAQlNL0argXIwOQ9uTv+AvcpZ
I2gC8scVkkl0VSjzCFhvGv3kU+M4agjOyTwreJSPvJI6qmKe36qZzJwngiMhcihc8EuZ9g9cIhvR
6a2Q87C86Pbhi+VGbjV//RPao5T5DNQDXSGLzw/8q+eXXCpIkIVWo1ouy5FxZ+7w8AtTetyXCOaX
KFm6n2SXfhWEUA4Y8So0mPd34QymN1x9Q/NHt8M4F3PpmniGo0w5aX9j2x9HK/hmc877rp07ilST
tQ1bDxj4ERgLIkp5DDbGVW7fWYcSaEq6Wr9QQeQmy92MNTRm31ZhBvfeGD+EylRfxFQ6pcoHGhMN
TngMhPFRSFDD+qlxGlW3qzRH6Sn+m2bD/S3EiDX8d1W9c+OFloRjEj73G1RxLGUx3ZfN7Z/NEHyM
AdXewhXsR5jiyFIdBHpsJH+byfBYuY/vNH31fQU7b+16iZLwlym6PLeILOQsN5K5bw7WzGgiTPui
FUkVJEZ8ITcVYQUEcYmCKPsfWOV7O3hQcNm2DfxJLPz/N4sKyQUGI87OCmEPQRr3OrDOKvQL1VrR
5pfbM4aOrQPhIlWcKdEcefe0GdRcR93d0iXJvjREpFq/Jh2j5cXxYKpJHF7pVnZGzmbccsOGrGAZ
+2br1Q6J7IahYZQGhtiTVuV0vfSQrnZnFAu9d7hotqmh5NZsaxz4DXFeNXSgz3GJndMwPgKzTmya
ckovOUg0yqHdng9u3iI9Lfor18h1OZ0s2TG/eudr7A18F43v05jSez0YXdWBcFWeOm8Lj5hgISmJ
2hLfkvbABaIUqEVve7QzXwm/UC/dpXvziGZodlh7m//x9UHXS7sCUkQUIPwOpDJMCqPdlH10+KIi
A2jU+RYy5iclyS48LJbEk3mQv9g/gGckqvpQ6ZIGBrC8XE9vEdwfyicxZ1UrozbLkmwsKdF3er3K
z3mJM5g6B0U4r7bCMlnJm+1qkEPFEPDFr/FO/ygzmx67u0+rcxHMqVvaLns3nEDZMiUB9yuGPAds
4Zlzyy3sAOIYL1zEbIFt376PeI0S5NGJ40hY6K3DKhJ4mtsXMPC3k4AQfw9rfxQ+CD6NridMENC6
fvgRd1SQXY8XjMGSbbWIoJMSSYsX3eC3wxMGld1oVMujgBw/4stzRElKhIGiiZ/9m1m3S2Drb4De
iGDVrFtRW3bPtG/3dU829a8EEo5It1WLNu8bsf/xyul5JhhZtJZtFlE5Qy9ZBKQZEdzMzsNYR4A3
qnK6E5lzGyBvutHVrQ84ULW20QD7P2Zyh1ITKXhchY9xCXZaCV302xGhSdpzzZ3MTYFfwAYOTokQ
SoZ9SLtR2OxV+1GnsVZ5/qF6RqChUDSzOUL6dmMTOSTMKaOBxX0C8omjKyIzkItv7BaTQ0QOn69R
21tQzHG2TnCAy3E3wyN2SqjR5Tmu08j2nY+TETNrSvqnrg1MPrBuoA7p/w5J3ieaYL6ZGE+DD+rH
JUEd4UxcXu73bME5/TTKihJEZ+nL3cpTeQaahheHqrBGB+n1o3/zXegt32nrBRHqQuuWBuI0VBss
5kRM7wEHlSYOTGecq+hRFaE2IU+rqcgzaNyAr/flofCdPpz0ZZ5h7/e4vf4h4biIGhxwgMmEcBBT
RWwpColVUbUb94+LjO9rSG+WwJkmEOyn+9LgkC0xrIUB60Fw5tE9n5SiUvHA0cqZhIya4xHu9faY
b8ZThySNdFtxSNwrvMYH8pGPfwnoiPxlweXfyCXOHdRQLR+qZ4f0FJPqHdOIje3ox/jkqdiFr78D
YovYIE4NNgN0eD2z/SqJS2vu9RfcnLFwS4XyvAyWQQLOwu5rLm07LgYQ9ZXs4ULZNKLXGhF1G3iw
u80NoaoGiXYYoZAXOzzDNTvMGgJKxwmHt6MQWB887gcSwr6ZL+RPz3Kd97F2jJI/3CAUQ+pHizy7
FSL550MPhR6vqO2SzEUWU4+jyale01omocBYDx7wVRUKHhmZ6ABpw8KeJTDyD/KeoxlKBbKoE0Jz
w6whD0CSSijdv/tj0rQ7sXZI15zp/vqthZ5cx67uPwv7AGUIyyPrzR1GxcG8j7Bn655qu5we6aYx
4gOFpjP6LG12UsqBoV08p/OzvOAUyzjAWBRthbmLPBULIq6BlyLQMCOpH7YYC0oCu/ua16yC02Hl
pSBTXC5FZ4oJkD4W3Ca5l2efT2exFNVdFPKeImdqNUO6FEvrE/9+9KwCXuptaJlSiG83GH5pZNPl
byAgzhBVdVBz9bt24ns0yiy758m1kbKC6rGKzYjPvl/j9hZ4QyE9YwEQdaAo0CKCRpAqdinHwIGg
mNABeTxsVX3k1XtymJkTICdgwEpSaNtgCpxxuDzdj4EZszZaYi2WvPfKRvxzo3WgYP8dZHiJRoD2
fAxuDQiYE3m8Cas9691hiZl9ml9XlXzrPBOjRWThCWPrMN9ScJGaU8tB/XQaSmG22DNrhJkANagv
paSI54Ep4qeSBwRqQB0B+5t4Zt2wcDiBRL+38a0KavNlxN/hB652m2OhxNQSo7WXlRMVcXMejq9W
jTGB2s+Jfh+XPBWHUZ9kbBCPCpDtzTl54v/eZCSI8UbHVpvB7VxKMs3sS2n7DRrXNg7SnFUAtmnx
g4NpVMTo9WkyIZzIVOkY1qMyjfqZMqSm6ku0o8oD+McpyPmFvkqpTy/4vUO9lXzXyDz3d/eguXt3
0vNOewk7x5f3OMMP4l6E90WeZTlib/AOI17n8utwjTdFww+ASktE30O87mVBHSUEiWRjAOcXQBvq
jdCepU6QmU6EQjhz6WjKxJxKh+dughSD2nCbfRJpm+rkk3HkqiFdk03Wjx5ujsKnE/qLOzZonPsG
gEIgL1ca9AvVHIPcxIG0NZmsTFqYr00hHjcRJFoRhVKg60wOoXtcu87GFOoAu1LYYj0p9ZjtuVTu
3BhVGhJCrJ8szCjYtVASwusonwKjL5r/vmoAAhlBAUFtJiQ6TViP5vVYoG+lBX0V1PrfPUO8Z+mG
WWnI8Ixd/jpzAy1XTIhOy7Qe2P7Z9EqCFtU3uycfymNNmhMQxXSaFizb7NgKwxjN1tY7K8mVUVsX
bf70oYulNeFU+yAOGmz/XUydj7P9PoyKDi4Y2qaRpqDCGr5duwZqMjDoLcmMX9becXq+T07epKEW
Tqjz1nJ56VhuK6nIejjgb+FJtc7Ny4V9nAgdn5NybKUIUbeFEOeARCHwTBMJKSNAcin49jietOQB
hLtHnxuvRs9BA4GoVtOxb844ZXKaC8fdVAlCA2q1KSGfz5uSE2XMAeCcbNx2F92qjKFB8wrDV9Ok
QNORBltqHNdwahg4qv8Q2C7JPlhf0vejElE5O2ptNTHbZC6UNKDlQcMp+Bec9SHW5MQPF8OcDvgF
sVdyq2co+U6wLdnKoyf8O0iZwEK3xIx9xfiHsnR3Amyl3kYlornIJPK74U4GNnHQNjV+ExCephZI
QmjGq/NM9FC6Z/pVcrZ9zt1H3mNAQ8bDgYjLtZNdGSHjpgWuKNVsmvubLIUqQBdT/Zq4/cEUlbwh
wryc/bTHeFdD4rfvMthuJDmff/IMFg8vIQ0y2Iq11x0lO+YPgSIQ2bYoO9IV38GALLtN1q0NjX31
E+UkAGO/lfd5/Jrokl0AvqPK4e1cRZgm9bgUIAS6DS8vRZ+JtR2hkrMsM+Wu+W1oMHix0txz7Zp1
wCdVTifZTBhNMiCHZ/t16c7IextGaQQ6rQ7DsSIraog93GPrRbAa1o42/X1fl4VCk0tmVY7NtxP/
jBH5te6bDYf3ktI/vMY9vQlzYIYXatrvYrC5y+mtAAZ0WhzBikRZUImCt77FSm0nQfxyfV9Cl9Dm
9gXjc/antwWUbq6Jm8Qgdvks5tOBZnEoHFADOFCqygv8NRojBoZXaDMI/xI092UP2b9HPiV5E5l1
SYgi6Ic5HjAPVC2hNXMtXxF7VRAMhsGB+pjUg0hu879amB+Mn+XDv+vwVu0K5cGUhOO75n+046yp
4GDkCfUqcF89l6ugZ4d2HySumipAz/ny5t3Q2jVQMHwIKvniu2Np4vTaSGabd2QblaKfoXQ6BJqh
7jLRFgnEGSHPDXcyNWhPwSrGX5VMUu5X3r0K+M3MT14ZPAgWV7L9gsJh6fshsDVmG7pOGLBjILY5
fZEuJnNgP1hw1joecQXUOattKTcSS8s5A8KFyVk8xtTUtN3U9XbKj8IudRkNHHImZdgxKlZb36ZP
GE2plbZD7UDm1Usmrn37zt0xufxk8oFMhwSHGHm5IfV64rXkiVaFwUY2DQEZ9DHx/CUmlOiAGlAL
RWHi6iO7xdtng6QnfNDz/K6NHjoloz4vy/sRWlFySdjwHzHKPgk4yFijClIiijG+QFUgYyQkXIwl
aiE3nV/ffiV4079yKy3c8+EPyUHDEe2K4i5Vzv8rt/H1xjOlvzkt09BlAG+5eGw9am1XnfMCSXx5
oWorgem1G14yoKnntMRkZN4EQ9MNBw2dJePVcPdBkrcEr8uGuk3ZxLCI/6nhMl7iHJYh5mMJP25h
qMMU8L3Iv39p7QVJVWzf/rkJTe3GwTRQzhxbpIjOaeyQGMbpAi2AZmtrr6xUN5aUGT5iuDrBti0j
F/GhuoqhCtC1D+0okNUO+/hHpXC+HixNoatx9taWLU7o1BBWousVVuUvqABFbsHJr27fN5vF/ycN
A1Fi4QBScoiDJECUlx174OjO0QtTNsYcrzXUwydk2VE4iQSbQmjx9FGpT00EBiK3q7MKutBfpveb
o8woq+gPML6EalW47NOLoyIC0JPpflAgZpXSoIZ+O7GcrLMG2xZn1VZtQ6RV/9oB/hjIkJ2Adxhe
dw1eC6yJaGBj6dwJJ+nFKGLMGDJjFgb/4gdSMbPLwYhOo7O+HynzTv6Im5zyItwislawW4l6zRx+
lPre3dWG8mxfQ19Zu6D+KL6j2GHeHPFgIHUA2mWR6uigubPE5JfPVEI+0fmhmCvVwY8fYPXzQpeR
UFBqPWpQJrvxAEqpxcANKYyNlcroK/lrD0PzE1kQYsmu7sjnnJYvYXcy+3sAwvFBZUVRqtYNK1gw
iOr9odNINy4U9eLjlQ6iRlt4LJKUHzrekWtGEKR4NsEwK5z7GVGZuaXn/cSDOx66XXKF8lfAvCaw
AyIxlXxJ3iLu8qp4caNXbBSkHHL0lpqZhBRFXirpGW1zXN70AulnxTBsuys5nZ/ghYOo+6z0CKZ4
HIPRARQf7LnVnlWyGR0JWvrtKdDTEw+LXemwZJZEYLAS7XgqSyzRhtYvoMHfYXWPcV9K8N2sq59D
cnvpBfNYV0bMdTPwUIJ0CM++xSQ3eQTy1OocstqeCf3EV/jAUL9JpnFCHtJ0vhXSJeSWdNq/RbVD
2J9Lppi2rOmvbIMtHMyC7shQMNPtfUti9S+r5bVIb4Mr21I+x0T0mKpKNh1LVE20tRjAVGuIjIvV
iLODSVP6A65qMjonfR066NmHC+QEsjEFrmQKRfZBh0lddPYb5YaNE6ezOvDScYI+SJiAzoaeNYdj
iQyAukvHahRPDyPGCI0rQmgdCSb4/+JPkAdhsmsoQbq0AbKLxtp03lYf5fJJrZdTK/WsE+Hh5IAX
8I7US/zTJb8Bt1+7yg3JyGgWA+tu0T7bEx2mHbkDBKGvyl0rP5aU4MMRSTnoQANXznDYdusJiM1O
HLJsRINPKqTce/v0Wmc3cFbYTdYV3dM0B8AfqpVrznUX1xKSdoLBGteJVTUcmsfV1cEJHZ7opXZt
d2L36ZXsUrXxiiU22as8Mm3uQJvZciGsIwCeJXHg6WCsSBNmODJfmhQPmHepbvfZe/7jTK4IIFNm
FrGNejl/epP2rU/HT2Qe0wKzBFHXNZhonF/M7ADhra4Qhj0ATfSmAFHv/vmArHL+NeuEJgYKf/JS
LxYTcaPOIUZkHbxyMXXGUqyvW3dZTXNXEfeBfZyjPZrQQYSXEhbYqLzB0007V0Rm/NKfDi7XI5Mm
Zdkpv1sVrIAKOTuyxJmlew4C35kDsnou9/Ay4Yx/0hd2LZu44dXYMbsxMInh/njCYxyHrPMSiLXM
oVQI4Fb5coB+DlnckPjYHTMbQXiXrF2XOL6XtrQDMg0ijeFwH5fe4JhFZ5EFnl1Hcn2Z9Fm5xR4r
/JdVBKHeuid/75Fd5e+eQxHGTTaNlFd0Uzx/LCgW3iuXxBzsjHuVtlAdlCit0cPtElghgk8JzOHS
wEFZUo6COC68tFvnoyZcGX+GtOLkr2iJrIFChTlIL3L/lKnpA5YJTu5RKQTuTK3dZBhHKH4b+QdQ
BZ+uLusAVBF9+EAJljqfZyeBApWmAPD45eNx+Gqsvmv4iZ5V/V37YoQMbavlThgwYvaI6uP49EAY
5wX8hCmGnBW358AJHa5Ue2TPR8ppu5mm752jIjK46iHuYmUiCfdeGpGf13Jbdxy4RWgmbz+rxUzN
y+qtVImC4WdJJKmDcmSeYcUN4CHK9mIO0UDBNHdy0qAnLLi+/yfeI1fOjPFxP3sjOi84R4eeNzEt
UgWmsA85CmA9wyNb4ZgtsLwVvYCF5yudySVQfpiH0lqdRz4OXi5ShNN1t4zyGLcRsqD5Eub2wJaD
LrNtLYu+COl8EuKECFgur+d1Lj+zKCGDtlrbV8auednqNxAta0Hm+T0u5mnWRFppUHgW84CtMH4z
CUW/WH07tiPNVA3ChFJCAmDv8Po/tpIIhsyJMD0hr1sl37YngBTy1bihxoN4vDX77r7t1O6LsbAm
pkkkl0rj7XnOJg4DvO/QsJbVw+RaK6GDVQLgMT5fZ1cqtAhJ6JwHm+VzYxIy7xbE5u+tBBdOTsCI
RHQLUcGCGKALumpicBqQ3GEaC52iVdCdbEgFSurNlJeGYMWQyOW3wToOGnl9FtxypFtRiXtHKW2f
AqKgpA1PbS5fNeak3Dj90sgrH3iGT5KQJX65rotqhJIS5xNSPRuR1DLiQcMytbWfXr8PTc/8sURy
q2Matx/438CsXYDTCv4BIsWV3gMi0zmuNSCq9SmXJbhasdU8UEvnnDbOMibi6mU7hcJ+eIt9X/t3
nBT4XMZWIxgnn8+MwAyD/fJcpJWUWfV0Qxg7Ele4L2ukIUp4L2VjzYZbuiKgnYB5Xnxn/Ok2LUj4
29pJNSzTHKa3BdtxRQzRmLooHc1YLV+m+qHVMzbXNV/Rs4QRY6hRB+MHYPzV7j+iSh8+b423MAwS
/5cMbD1XwYIV/Dz+oH3hxG1RbXeXbnR/Y359I3bXtywXskTgw1BXykPJS4yPLbZtib7YQWEyDS0Q
Ze8Li3sOQdICVRX+MwmOqCMtjmwgZv9j9LHMsh72IPB6h9dwf12yX7G6i0UWUOjLIBjZ+TC4L+Cl
h07NC46zZD4Ft7WaXz2xEcaDWBHVR69stJLZntnuAqIJ6vcuVV+MndDdcqypLijeqtd6O3xygreK
TivHbliHOwikkz6ve5FMTQv76B5R2ubQ4buWluIA5X08h6SdMAFrt3cE0ClLgpiGKgWkxMHRU6nb
fbIjCa6inaU1yXSMvGvbLPGIezSAs5y5cKKaPKQahaaQ5o8J2bBTK691UFIaSZeh3F0TmDXMjdyL
Tjj9+YdnaM3/+Hh4TmUVJ7hki1IvGLLnyVB36+LfGgxG3fYUrnRAvd/+8h1e1xXO05Ikxjwhj8pS
O1BT8G0S5q6GlH+Nup8ByOxBs5bz8BrPAL4tRS++WbckyY3MwSEES2PlZ2vSy8PmwN3COHvuyMSh
DqIKCxMpgRPx6dkm8NXyr71tDt34dvMvC4J6A4QrvsQhp1XEiByYDYctdaUNyX7OPNeFY9BUrqMr
oWwqDK7BsDcWAHYv9Mqv35E0QSC6WDK7+kKvA/0/XaC81MfyGpG37XeY/5SuyYFL2ZKUXbLlB8yX
gMVIJVkG5mp70qzFbDggMUJg99rLcvhzDX+7GZ0o5G7f2AwyIrwKCxPxC0q0GWwE8XKRYV41q9Jz
dFcVfVcZvyrwHHYvKIqLz3tT4fknIH8fjK9WIsUufnqRHf1CmG1qKoxVoOVxfEQ+zMYS3+fd+lNi
mojM94oALSHws0qdjptnZugonXf/iUsTKquROlbfAa7uIkbxasPusDVcbw+ohpJTjVpbsf9O2/q8
APlCYEjrLJFCDW+rn9KGNLnkM5ShsGrw5VX5b/5iE1EEHshgSfv3LpRjmBIhg1FvwthCfERsHEP2
7mURmsngjgm0qyo9XA8YVUdJ2Ez+p7QWNGbZCUV06OMXDLquCwAnPrFcz7aTy3gkldvst9QIePLp
qm0o9+ql+kuSG+x/pamazgO3au0wirsffBMzCR+qdMcHrHDBIpZhadx68h+t5IrOxo1Y3Zr/b3ND
nj/m5x7ZcHDkdGej9nAr3Se94OH+cJavZRskavaVSXB35gLMF8Fn2B22FHdlfwf16b460T/dT129
pg4RTyHD7snmC1YIEJCNrjJoUNpXa6eiJgS2mL1bzCxEJzvbJhtZj1oKBgbVpVg8MxSy/e456+3e
UekIbnw5Smpg127ZcG9LL3J9pKu500GdoqW9FkoKtEwJKPfwxYp45r8/YUjl+c8bDa2L3EKBiwCp
TyZBmW0E1GhAbz3Pl7mVidaed4IkcpwtRes3/5HykrSiYfrOy6VZnJiTQvKW4QCgoIuHJI4I3PUE
fbq8HkBVM2fjaUCXhfUxGBqc008Mni+YIMxAJ8JTuHdJ21mcEKI5LNnM5ZrzavZnZw66wEApxyVf
oc7G7dsXI78ZrTyzz+b9Xq+DF9n6GD2zeohDD3aLAx5tQQlPj6CGLrsEGPDn/j0vbZqPC8z+KqDq
N1zOixKnWONUtfZ9ai3/RlWbmXkVU71hzHryzS2sVSE9L2bcOwiDyHNerfILadUguWpd7nFGYrTk
hjZE6uB4KKM7sP4PCUK9cA1Q4EAqV605WDYM6GzR2BMusTjMYncI0mtXU/6rn25ozDjctdHzkuEG
QaiiWYAZAtS7pJhlG0j06tHTT1Cn6zY9MFsSapSnPghd+i3COMCETbLMT+JVV1zVo1YTpuavNlgw
Qft68lZ6CS7cB+UG/ce5aml/E1s9WWJ9P8QblrJnuj+XdckQVtGcSkVg8i44KbfjkMfRipd7tDYv
w1A6NbYmtkP9fYmgwU6ktTpVQnT6D23oA5Do+67YCjPHSbTgbIG9K3uH0m34QYxa+R0d5njaro3a
eMVA3hJD0etgyTSOQmP8x03KB5UzcSDRh6un13gvO3WmFXqbSwlTpALcls4hmLRP7NbewOCzOyrP
SOk/2Jfnbnd9D78BTaavhVRHqQCnqOwgPU9+bcU4K4gN7rYsCNjYo3nC/oqUvIvQi2gQZx3nr7ip
Ai7AKHIApJBAIQmalESt+Ziq+6TDbB6KSfwMmTYPAU+JDCepK6Gdo4Xa3OkbOpKoc7ne88vLcEmz
Sf8rTomuRurTIz3rsy3u5OvpzYbLwGAWL9NfZ0pTUEE4dqk1TSyPRvN+Ae2wqna1zHkLzO29ipbl
lHYM48A9d0+B8HxXGThR1HvANFyQ5IhmK7TNBQ28B9qvI17ufdBk+U93nZ2r+6I2krd0qKsAXEAC
LZJXPl8eNSM3+J7EqgdTs6Flw3fYt8ynPuBMBqZXbnil7j+URR5qlGlJa2OkZKvalu7UC6zK8ys5
aX2/rRgnMygwzyscZ0M5z2tTQA+ENHyDT7oGCkSxN78ByfrKowFmTAvT3QkqyL6AF9tmaAomLHX/
eQKSkByIMuHd2T9yXzHGsBQYhydnlw+Bwe0bFKOZuRPcD7f7Y/YykybUU+CPiG/KCK3nfLKV8hNk
ekPOAn3pqkc6d4TnzjtC26A+e17WI9yDqwuyZGqmet7A7IkwE+ISdnR0TKk1jvNeZ8mMqJF7h7vd
k5xzFgaP9f72CvOVi2sQXl+cb+mh5hqGyJA0gIbBKlsG7s89VYLDj4N6VeeQe0MinOSienX2zgTu
YCbRytKWjfywAbVgJRxyLZ5T7XrynkQujzudWB1Mp8RwhFuuGcqxjQz4jDIfgmqJh/Lk3aI1/ykg
43yFWomYAOkZaPEMAaBWLoFz4C8AGIu18xowJE5kYSix9ipE1IBjM8i485ovRY18BXfED1hdPCxI
bLf2vOcoZ8I1FPQpjDKbmaNPC1bDcptgLJkcsJZCGmEO2EOOotE/fDjgDRAmxfFOc5h9y0IsRq5D
J0ZC+XUoQFZhKkfafwfgbDijR+hbimHFVVUS94OasJmokDFjhqsttIfHkn/yk5PVQhJ3afz70Er6
HjkZFmXJTBnHKXEI6ABxx9UJyBZo1oreiYvyZb1PMSl5ug1RGx8j+L6u6/1S8ekWFGc33ESgWy88
uZm8rBP6065d8QCZckl3+WWwaW0Q3LMMd2DISsu6orMJHuogcBIeMMoSRhUC18Sh3edu/F1qxFCa
IRbDxRHZ6Y89l5BB/UwzAy5BUbGF0PErV0teBlq6YaIr0UHZ1TL314ngv4M4yXJEghy3N0j56cIS
XKkrWknbBtrQMkFbPGWQu4Ygk9i04VZosuOZzSx1xurA+Pb07aYQPE1wfKEZyCEUqzb/dQfQ4E3b
v2yHtmcqLQWjlp3mI31CPNTg4wDWOgHMh5AnUJQhOCOUaQzYt8zXy0F7WItqQxmFT10XwXyYMM7L
BykmmYtCXVa1c63/hGfDmLkRItLucSGfvLjwIBwHrJotyGNhqAlR0vYRC7SEHIMpUKRNv6H5FP/o
d6RLfys9h0jGSARw3+dGoqulZpenBq5k7qf+tWkx8jnNXY16VBFDYbPOvP339pyd2dW+n9kpYzke
X/LmrRVhESzlc2gTo7VJjbzHn/VWdYmmDjPOwpCWnkgJ5Zrg1aPLXFtN11eVuCqqJp3eH22UK/oh
1gAd5JyJxCMbrxixg9augLRgefHZJKYT1b0HCMwFpaTQ+OJ6Of7t9dwtErnTK1p1RBzVKd7ZpUcL
eMl8QBWruyw0+TyDiMbUyFGNI+SYpLVK+ZdtzJDQsidzv6fmIXOV9AFEA+Sjt82oDi6i2UbSXhLH
QoJT+IVyo96BCqSXpv/ZrfJIro2LU1YDCMQAUaQA4TQf6glyxyeRHd4qSZ5C5a3RjRkyF5OpBp8N
4G1ybH8ePKx8bIBXw17gOASYNmNz9i0kU2IRnKd8tazCSMsYrXOOqWEqzYQLTmkrIooKnHyX3VgX
WUfaPLvBtg0gKNbvh6+2QPUpoZJlV/q/In1cpXoJsXEZSFCKuBBYoJHrBnX7pBtYf2lavGQaVquQ
4V+XzzX53Sl79toDZchTWfrnBMuYexWoTF8iZeX7IXt5NaNeTEuW4HCaxuAjU+z2e2w8a78+RLug
J5V1qEkmjfwqR5muQkkAIuUfuOVBYlMZVhK1X/wdPZnaxMkGNEpxEe17rJMHZZcOK1ZfMt3L7q7r
bloVxw3ed1kfoYoi7fyo3mZDD9neUhjnSRlXIYXorQGkyAsm1uoVjs+0/GCTgEST7K/BJrU7Hls9
Fp/KkwWFz5xEexjZrwmXXtfczMwBUZjYqGmejSuyTeCKtiapWcUEP5sp60mL4nPeM4ubYl+vUm18
PwzDMetzwpfulOu6EtdGuC+vHZKCVn8pKyA4eZt/5IhVi4a9JO1W+GrzYBjkWm8gnzmtakfWxFd5
zY60yxwSSHBo/N4DA5FzzsZJpbtpbunP/0Ql0DO4UaS/SNpp18RFKoC3o4t/L56nWHEGCLWRGoqE
Hyhvsj8R2azR3Q/gN9Hn7VqYW7hUmt6oFg+tEWgAMIEg/l/p5ULhAmEC/Zdt9SPrqlV+W9yabwU2
Ikv8vJYZ+U9ZqJ9T7d26p0w2JNwOGg8qy4NEW8T4xEk3I4lkad6x2inlQ4EXPowXSL171WcSXjnP
rA8xJ/zcgVVbJpKAqVvKPFqP63WT8rRPPBHPdxpN9hgRcQmoUpfhFBRNtFo14HwuxIi0lUaINowQ
CHKBs+YfgceJNcxR9NyDqto9cI2CNCVKojWlyEU5HBnYBg5voCJmR0K3la7v4vgMgho749AMWkme
XtKPoHQqa9NOCZt+KOo9koICsH7wWJ5OV32QT6a8xpISPqy6T1yyC1TqcaPhl5+iYNmaVcWYwSUT
8Pi3YIr6+ZrAOC5UWn+ZubsTob+SstYtiVgGHV1yBQZNOJLK3cg5qf62BGksYy5ptzmI4OGpsKIn
femQCN0jhsxOLBt9YYFV94yoO+8Bk2iOoCTqOhUQAjXrd7FXZ6jIzM4lt35Oev6r5KttlhgQts0C
Dg9S+3NT/vGnXMKJo9cQVpQwY8GQXZNdmtgBzqhccD6nJjoYcQKkxn6Mhd4OJHhYFdymaVKV7KnE
+AI/teC206uy4Gb5kuMR3CAL2/jTR0WyA5G/BSnaa0FPQwAKF26IEfdXjaw+iJbT7IhPQtiTmjoY
ofwEvybaGClBNaFIlaqoiytyo31BHFcw32s/VOzSENEtGNNRt853LRCNLkY0snMky4A4xTZtwHVo
27VMJHM2ViZwuAOXXspFpmWHLBK1vpUQJsarad3P6MfzD5tMn4Cmt3SLT3atHKv543ezjiK+QqxK
KuMegDRg5han0goBL5Rr3/EOiJm7LJZlV58OrF17i9WMSsbby/oOL2lk61SqsKAV5bBuqajn/YWT
E0LqJA0iU6AkN2DE26sGKyLX5F0tfsu/vRfII6b49uPtaEkZ+rEoUXlLhjUwMRpN0CdMA7SzZOgf
V52JnFlryU5YMgnbuJY1WUXJDIGEqmpvzlLaVd55XMyQ8ncTPxQhhGZQam9Ne/IYCkukiRtrE405
T+YrBCyTlOK4BAUOgzQra50QO/bkaE0zF9o+z2mdKyNHGLHMIdCSEmP8mj5MuVdwh0w759kOXqNM
lG4HefGdCor7j/h6eyfnpwxaRI70T4BGUzeLvM9d+7rTrLkIdNpMY41IePrdXj99gazdisSXVn0h
IJtk3SEt/XMWqbgQWpfZjJ0c6ksQWiaWsv0dbx/6SkNo3MM29CsYCYDpplJx0x/Q3vTlccuKNwkN
8J7FLx8GTz/d+I+JHuJyo463DaRdOEH0jfnAkN88Div8qIkmWXdk8+xhEYkRGePsHiVRXW4Ot2lQ
qmi8Knw9OT9RFBKx+jeMNhdH9EDJRotrV5X9APIXiMxdqNK8nA4h2eG8VUonhwBpkJ7KltvUn2fV
FV93OpjD37cfIpVwrqmRp9bF+ukVAHD9YKI2R8ahmPZabgB1Uovg/fZ6gRpb21mDVfhvApkDNAvB
7vPTQLNOazotR7HBg2cFrpziHRH0Mf4OEWcsjrZk7sCZ+Wm3pqIJNQvaMsSYhIcSZBB8/BhI15pE
MLS5Klp1nuEWnK1O0Zx/yD6oaP6H4xod063YcxfyoNzXflPrDgeStySYy/Az6kSNXsscPeHCp54E
2AE3Lk1FzXLM7b3b0WeVVn1BD4R7vqH//5Q98xORZ9jmwogwUspNkeLkIfYDPexsUGeFjdyqcPC9
qk6ibgdFGWeV9k33erWu0V39mj5WVeeDDVjd9pHVpLvExi5CfWUuIPwF90GOlCxT1GACGgpsLPfD
m01I0J90LpDtZBhhZVn7PEjcjK3rlriAgURgZz4H9n/Rdxa6OgFnUa48B8RScyTCq0V3r+lRnl51
IF6MpU/qatULqjOr3zlWsaWmD5m7eiZ8PgghYScQz8+RLPYpnR0zkL8RlN/FRU286RNGJLa+vm+c
HaT9zvoKhHZeu5IV3I3NZ9rewPti+u/uqsADcpHbf3HiQHcgnPrtqw1iSSpujLHxI9qrU6K89fUl
3p7PVsskbQTH39VkmmoKauOeusEfzgUFELVy+3rTDadQzEIJapFhzj4C4brEugrGAGceGpfO88jc
i22mfKxTo9pHalRUDiG7vPMK/9xfn1rDOWdMYeqbYONCyDCF9UgcBoj/mbaj5XZyJg4r+RxijPqr
sQyCC7vrEdSZG9PXYrm/O9strtggCUn+TtiujfvlKeNcGdnS/70OnCeb3dG/oyUSyLh9bpM/8Sxi
rDQg7xU8K/fHy6gWXaQCjNhRQIC4Mh5W3Tjkn+LCNLWAFf+5xb13Blxoll1Sn1FahguMa5FvQjwU
da+ImCiXkgd+ceCfmy+azxMBoWhzfEQjcKmEbSNpEmeFOjDj6AVtGLB7aamVGfnNK+89rwuGAU0s
KpMy9BE3bhkzafNYZ/j5zdvSfB4fcsiY+qn2mhthEihcJ7lwnVAv4Uyo1HTlaRdRWK4TYlIvcsh2
DgC+N0v29WKfgxIIj4ZYyqLS94hsg84PnsvG7Fz3C9nfcd721GWc38TIVW4pKmfptn9HVl6QHYGr
6Isp3w13lD4tvV8tJ28a9ISXDkGA42aNBe7VOqRoETe27MAfn6riwq6PlC+2lPwvD+bLhhhrEk1z
Lqaa48ajmP4Zk9fqyle9Gxcph5B3Ge4FTDSmhXzUHJOa3zKPK3Eipm5X4nF+p8d5hu9LG9eTtVo3
9WXzVgo+mzMlE2UeKXixTLcBQKz+MLnjsnhMuj9F8R79Y8zse1J8XpFbIzZxQXtb4Wtu+DA0odDA
DYQTH+m2ovdtId4etxqum1P4j5YuCVDmhFWW/swXDj2X+FJ5++AzO2qDZ1yA1Xp4im1cGd88OuNV
cl/PI0OUcLa/O3lDTEbqyy0vtvqUJ1wNW8Viq8RkZIEe3XyOqWAVoNjbfSu3Mvk0e3CsZL7Nwwgu
uR5sgeTOnicOxV3FlBwgvDqtko1FGrO3uyYpRD3WZIZOXdjKcwTBHDq0VuU0tb4BEJRtOGyb2bau
P4f/PmeTZtWZzz4NlGc4pRxHUkcb913+gKIGc8xhhp96JntrSGxaOeSj76i2k8h4mvI41/0Z0j7p
l4Me5a86ZLO02hhXS/NLbkiy8axTv26bfKvhMgkY5DG/9zG9EX4zqlAtJjY81yswzXnWNUi5DSwD
Odc55MRlSJaFqIHj6v/1i1roZ8aBfz/Blodi/rLrozV1908arEmC2jUnwX3bLq1k3RMbTKu11xdJ
FS8YZVs9RFz7W+NcaHiMhOCRbSUyHlWTyazSpkYPOFe4oyKnvoQOhH0MtWh7oz1JTqaGaz7d04g2
o8yg5dEWFxpgKzo55jMh2avzV1q53e9XQfjGs6O17Kcnf47jngR3Qbv0fq1q6xaty+C+molWIkAT
tj9uol8eKpKzDmv6Rn8vUOuCn7X7nhYXQs+jMhZ842ZhYFWFqKr/Mdy7Cyaq4hZwfMGFpMnrxv4A
cyVNsJdnpTAQFiM/BLMjGlOyaDK/0I8/nDzLGLmXs5CGKaxVkEa/ff5t/sbd6050lxXA+5w/Etii
fv1L/HvMd/3L9ecfmkk7m9kLV300J04aX/9FfX2/m2lRMxJAHcCx7HiuA1KA66lBo4LONG6jpVOf
MUMmsUgFUVqnGZNtaniF02DmOj6Z3fFVD8g3XxtuB52+VyPxfrOmR/4CBpvRhnUsTO2T111rzHxr
zaGMA8SwLQQgIVEiAIDk0WEFaBiWTzhA72tOBZV11b0sIbN9f4iaL6LsV9TIeKfN/UevyWp9fGe9
3fNXnY5BwNp9ihR2X+ICvn7qHgeBhDTpWkLpmS/m6Jb6tIXOaN2Hr1RLdUPgRobH95pT0CtDSQvx
/tUlkrRPp7P4T2aQXFtW3TU2AipJ49CLpfjE+EjWmqqyg8IfoBTmSGIF5Be1R3I4HEl4tEGtLY4h
NMYhPe6jmiTBIofz3mS3juZFnLJjkiVe2RUONRxoLOiurvhj9R+Bqvezmlxh5XnG9sbdH6oI/JHV
cVuONa6jWbJlw+cB2Vs5DA9QNJgJQU6NmnlALnul2upeZkcSBrlrS/+gmyGXNHiH1VqBHyAgSyUb
4Tr5L6NhL6gtTpEBawazpg0xu8knFwIMcfDBV0QCBAbUI1jns0c8nSHDxU66HJlAjp4eqeTUlhgF
kbx8QN4zZ8CyMIW/zsUGqOiOLmf5L8uXNgPP/gGw3CwPFugRTcbk0USAVGlia1JIslK3QwpFog36
E3kYkVDzasCmp2i2R5Fc0tIP8xxG2vKxOWsQGOXwXd89OQ+20yvaOrzPsET7LxdrvZJhqTptkpPW
cJnuTOE1ZukjG2cRZ/jMs81z9Km/zTbXNtBRVHvrWoiJDDD/aAnNZFyYf2cMgBIb41ZDI8prnada
eXuTQGRlUnpxslMT4jps4KDULyau+mCyaS6mUfAZ1YZ7kwDyeqeg8OtaCNfdpvqNj0Qa38TDLURZ
VO5J5OVhcSqJ1daMBfE57/mjTeCHUul6hS9BgVR/SkKTFzJ6eDQhhu/vwtoeQHLmmIT5S0ccJroI
Jc3PAof4rfZd5J6XtZsNPHmVi3KoJD0m+jb6X3dxSSDkB3JE0U6qqMxf8JQPiwR33vKIf2TyXAKB
lxiUaIbMEPeeC0AVu6uaehVA9vGIGHzVkyZbnB3GpCVOFmomAcA9D0NkVt8NjoU6WBwtaNht3nq3
aKlgjpkaT//wrSwrrnxzyx4hO5cfIc2jJFRPw4yw4Au7HwvEWCOohGxVjE66g+EWQfgDiK5gzid3
BhIUfxESrN0XPfgNydaBAYRuE4AENKSYOx+PgyCOQ6WfRB8dgxkoCw+xIl/T6JBvI8n9kl92ysrP
7swQEtKMqcfPcGqHnuZdk4c1nrCzcGG/5fNYxx9ZtANBJPe4XqkA47Vsm8iX8EKAVJcPp9Xjpc1L
A1lCZV9ZA7Xxj93FY/8FIBiz491UPUvAnnfVhiCIYU1pG6BjXFB7P325DKjbkgdeaHOUe/YdvEOr
bqMqyRzCv/xJ8g2H7qPU17tO738KejPJ2yklC8K+ZXnOx5/Ag2kRj7IRrjnYgqUnZQscy85Y3dKO
EWsXIb4ngDiYrSuiEU/+ekZzm5mY1MHf/p+flpn8hR4CfE1/Htch5VbGjV/ik+V2UXwUZC5Wws4/
RsvdPI66i2khUB1xuR7JUhzx4YAj3vS2fryWJw8rVMUqe6Ksy7pUvP1k5do4whff7fTodwuTZcf3
R/xoccj8nHU6ilwO9ODK7TDr86QMBhLnlV7cfS1XMWdGAiPa69NrgUC/2lURDU0Fc6ERoZyJ3/aj
2rLXvo/rJ5SogkzAlVn7YZtHoMPd6e/yvJG0njqfG8nGyB1eooeivb2WjcWqw3esUvgLXlfxtNrR
qPtz8xokuPZplQIb07i5wpn/n4w8BXEniN/DWY0LuyMO1QNlGl8f+leSNtAaZjslqFwi5LI1Vg6m
hJo++GzwvgXEoeB4W3lIXklOKOwcPt3qJhFKpwRDDXiHVUjt6ulPPHxzw/UB5NBP5ef+OcgQMx1N
0KdCfigvomh7W601ogsmIbFkfKTx4JI0RMkhEf0rgGnSinNBU4lWiH52h9Y34rHL9gfuJ8ksM4/a
8FiiWkIZmJSCyBI0Ai8vV+PdPGIeTYwFlK0ShDQTsD1OkpRJrsjQBKtoRcoPxFk+fhl5vG0flQnj
XYMq1v3TqtvSvmAZtR1I/OXIHEAQDLiOg/V4UF+a6gEo0+TekdZFZSsHfgLfQUFSSg2eu7wulkMP
GqaxkBQabu4muUMM8tDC1/e4iAuS9Nz9llvcGl4XPuB/mRMUyWlEY5PHOytIu5DgTycJe6ooWc1L
GeIHIJCGsS+OgCGFSFjHFLhgtpqZ7NMnZZNaPwsJw68+gmPqUcanppEfOPwDaYIRVnXfEaWLj+Nh
bKM8gJlg5zI4yc10OTD4wrpQvAZLmLdpkUdH3SiJNp95v9Y+JnYizPXPKNlgwU1D14GUfYlBo82r
NgAfG5WJS09Q02wpum/MYJNe4x6GNXU+cxNNXwEzyGwyzm/Dc9iiOWLVNd6zAFkVoyglvpilKkgg
LXj2e8U/KExigOSQEaoGoUtcTrTqCJhOhyG6ZsbFIkwhPYwvJHvLFdu2AlgayZYQCsxFTyPI580N
pyOjDVHaQly3uOkkOF4+LnGjvXbVxUlUcz7Q6dcGEhQWWmnTzvrgLzzbzxYSIJR9ZPE6Ii3d6zcv
+Y37cbxKwmwcQgv8JatIiOfjebxQ3GDD0TgJe72ocllFs4vcEdqxE6aUuGV43QeUT8h/8kabFtI/
j9zBBwhIPWVHVTm2vv8NWGEtVGxzCwTsNFX/myQ4SlXbxkx1Up5+Ak1k8JLVsWkAFbBGS8fziGPv
N1tHQm9H2RbP2kWdfT0BMoYEUirOq9+Gb8O6K6rDV5eIV2Zzkoa3Q5BPl6y8sWuEgTQl8rOxDyKm
TvU1CuBV7P64FNI6EZlyDdA1FyfYwDqgQchTjfWyvoeiy3Hn9pJCvP4fjSgoU+b/JdDACCutxyIT
0dEwHsXD/deI9e4ju6i0s3dmJpLL8NohNGMgFJl+HFTrZnNzpMiZ/2Fd04hI1AhkafYYGNiCj9H4
qsup1gMT0dwF85gENQ58y93S+kmiZryqYRdXmPBRJlT+CSpAOP9qdOGsjqxWa9bFM37eqZGKN79X
8JRcPwwdX2hjHTmHRnvxxu+fPDI09D7doH6LTpbWKRzEeVVmkjzUfEfKN/+mNDinvSMylH1m+tmj
JnlrXw56EYy7H7A0VY1nHlYyGLj0CTwz+AR/bMZtF8W/WwLoECy/xv9drDcRTRu7HBwGAC9nbWW5
KQmvBU7+JemduHDVRqBB9SyO0eml1FMDRoKinAS1DSp3dqddSlymxcwiuMitF4x703gqLLhbBmTC
70GkgGcmOKh0vIhbcE1Cjp9o/ldaui8KivqC2syCJS5dAXtZ7Vpu97zutGTx0geyinjUHnNWlzFG
JbdBQqlqSmP7MXcztQZoN76VZA08w6c+JeqdVTpygKxjbpuEfgU/crnKMrxuuH+KTFiFqcF0lBL7
abj27DdsnB6yMsxTloLbNE8VIYxc1pVAdGju254t5WzT6aqtlsIdTZxBvdxN2RcHedZKI27854hL
1+Wa4B9wgAweDWtH2TsAENGxcqo+blhuMVxlyq0e1PrshvyxbiGcy83l7a9lYeBlbVoKbAsAS2Ff
umfW9Gx7oNZsfAps58P6zQWYJhy0vRxLBfAOLtnCqyiNPkPQQxtGInrzAFgquh1ktlSjM/gZgmue
b257xgY9nfRhChNCDmRcPT8U2B9AjLPaq4XuBCgYe3yuTecdGKAUcyxU/Tm5mjI2/tGkEk5O+zUR
mT2Yh2lBPmCgmUK5Z8r7rdq3mQ878DwZhi0QR441E7DD5r4iSJZ7hoED9T0uTGngYti2DjUoGegm
f2kq6iXUnKcAvRN/QDtYyuCyNAT4kn8nxUTm2cMsMnopOr1w+xuRD9rMz2RtUzpyVL95pXXEWoZT
30YhaToruCCODGD0mR0RM8+Ec9YOaBm11zLFV7xa+dRE9JCcAVyLTGQYdudVKMCT4IIPz5PrjCtI
TXM27DOFHJozDsIyRBXqX+8wG0BtYk6GHWOkYp0SB0Qqj7V/J+anDlzFiG/XR1PBlaPzbJ4D7Ili
MCnVhVOiPH7s3rL8WexJx7OelnOCIAg+o5D2rwg7QqWXgvKkzfwhR4NDGgEUKuCr6EY1vug13LfZ
dyE6pehCG0I54+Peichu5/2rBZPpaF45ZSfCdcOYZpmJ0iAZFeIPyqh4W3ba+/eHL9y2Mzx76pWM
MHufGRv9JKtCBfP0TYz3bDWMG49IVLLYs9nRFLBz53rn/J7Sy9/Te5V8RI9PQXbu2bXeGqCf4l6j
WY5EUAuxy6LfJaUCq/mZjDfhujfOKjKmvg9o/UVg1cyhUdIPofms/UA306miSIwyQstsFJvTK3xK
zVnh4Wyprw9gP8dWV4grqTJEHjfXFZaS8j1D48XLPOwRQ7IJsKAEMyiWeNGE9qb09jFIgAXDaxMg
UaLMebVMp5W6OwHEfWRkkQVT2bMISWaP/Q1xkqsUMEzmcIfaBUyHEwU+FiXXj/Tjh6aCyQnX2cy4
oAbI01lQ15HTBsQTE3VP6iQ7M5+gM5sEgQpMvfmbcsf5k1eE0Hxuv2DvVre+MTRdjFYfKbNqyW/l
o0BrFMPJAleQGUdQVn1vCC/4ZdYH3MCQ+5nX9REv9UnjLHl7lg3BExxhStQPQ1xjuJfdwT7JeYl3
qBdn9yXBwB2EhrTcmgfxlH46EBmJIoeieCpS7DCvVyPfZr95Fs209kjQO6NTHbhFYdPEk2NfqgrZ
7TvpRk5kXf/GeGerieTA4Q2FhJhbNdU2hCMyKj6HiYj74NBymPYceLnL/4+1tzI170E9L+OJne7t
Z+2AXyS/cVmPhmxbjod6pHTo15WVWkRyTNs6vkd1rZZiifIbsqSig+b+2CFgH5fGALblf9yObqa/
TyAcROBeIHuoYUnjKclQpGYJT4og43nSsfGi7HJWX8BKiwAJzohHyAHdds3wi34DSlPpH+bAwhpn
cnFKBBbR7fy3/wlq+rEGFFb1NaYvU1c4pXoBmOw5VR3XprJhgRduilQ/Xo7thrB1ZiIxUlyatI2U
QUTjP/AkXHyqwZdriplCA886dzKBINakGEgYBevvV/Jl3hz23xhZEyy6ts+lMSVs3fTblrn4/fSB
Ho2Oga4oR1bwnBPu/tGOFsTPB7QP5p+kGJf3ZwPiX/kp5UygcmMoPqbuIlu/VPo4eBMvKqWIIy9R
cIhLJrnlL3v2/vYzqv0DG3I9QBQNuypNsvJcJbvmNfQJppO1jqiWlZfIpwMa461lSRokNBjIeijQ
vvg3W7ynxisT2RuDlVQB+CPvTcq1XmwuREPhV1bRedxndmjr7y6fpOO3txniJDsllKDTv6aYSiIL
A4OBzeTDJnmT9AIZjvZ1foVGwJerltPlOZS39CcudrgSpm0eVAtzTFvuTC4DCw0x2U2LC42XgrOt
c+QWwbiNrL8+vZER2FNSR89rxFAOegh2wU1AUoj544KBMv/NW63qgvu1S4y0Y9NYKAY1nRpF985D
Z+9JtltQJDkfMsVed3WhfzmYtYRkNhQROqczQtqkPmv4ZpJt5i3ikXXlvzrwDP20dveNLQfntelu
V5k+9Al/GPYVTLYf6ZgXMP2530s8/E8mdDNT5N8e301yaDw+ZxeLI27H3c85CTrR23GWBN5wSwb3
O2l+60Y+9SvxVBjvw0gNvVG0m5YTDg1USOtrbxHbpi8iGMOyc3HNIm0PUslzqq9z3gAiOHjWeh92
Qd513vTDGTUDk/517fTf7WKQ6DZOlztvtHHiJSP59VRTCd/Vtfrm5ZfU9YyQ86t3fUKfSTusdUVW
kLLhf+WjyxeI+p3R0wnjRXbBIxmZxkNZ1AxTpBCfiDOHLjsxX5By8jznS9mbQp7MXcTG2ST5kiJB
T/shOkxIlDn435J33iGyDWSiEW/SHE5uPD7kLSNETQrk3i41m8znSTT2HvWNKQRUZCishb7PqAaV
bFKuEdB6ABtp4HFDZchLlcDsSoVr4gbbasrJMyjPuJQ4zoVyhMHbz6TLzHHf85l60k3bso8KIke8
kX0v6g454MSY66khf9CdyTm4WrQomvIbhigrCw3kOvSZe7lrh7+b/AklZGbDUSbp9+ujiV2FYSRI
QyXXQPfa9nFseLra7X2by6ulbRJDlgDZvmdJiKHoTlPhW+6aLMMwd8s3F556GHJpuL6ewUhRYt0m
8a4pzGos/zs+1n3+Ww83N4RDvKik+Z1Ymrap+kVzGfIWdlM5ZkNcH265XLAGrpmwc1nazuD1kQGl
SwEPEYiUPvnYXKGd9E1/gn+vCYBbYv77WOpPD+7GeovbWtvDWIM9lwwgl6T22kObrg3MBHz0MnxI
Dic/g5YXfnkwpFgtA3i6omXDJ9gxtwyx8+XLCLoe5Cll7jR8Im3EA0eEqz0e4rijoTRC4nQmBO/g
+/yvYLGaMYlThUHXsQCerQKeIvPA6INGa8aEPzm0yd+5WJ4CmW+xLrOEdTT5TAgSZX5tI97JkEyr
rDgFMF08/Hdt6kBgR7jiqZpVnm5AZkQDOK0J8pjuGXx/3hpnAMDiu3H0SBNKZTUweDpuJtazTXVA
0jCEMjuhfwyxis2TLm9MKLggKaDl1+8jR2Tv8M1Yh94skswNnRmSMLCOg0QujCIWEo2hLyTgdBp8
POWbDRRL0f7tJ3aLDdxX3mdQ3kaJggWyjg8HXaHQHDdDUwYtNMDJ7j8nsb85kWSnSUSsESfAZm5r
YzQp5/TE+GEW/kYplDU8jH2XTxC62F4HeSDZDbqPUx4sg3fkWfjvlWecRBnQ2gTTfVcjsHb5+bQF
duGt7ieAn4oypIFL+AX1VywvfSSwMUY0gpCey399zPY5qDCStfzbRghJtWBYKFXkeLQz6UNUWY5W
7IDVe/KDdXCxxnniSQy3OQhEEDyQRXhUkYKdoCFR0QaJHYfelnW1+FdcQk3VVBc4HxqxwBGOk2Ec
skoBZIQeOq1UoODH0NtfmoeTRU1Bq7T5nCT8tCKw42HURGcd8CjcYTFGUMTtz/4k6j2UBbmNwPsc
JQZDXcTtIOsypKwX6J57fUC8nH26oHYwKcJHA4Z4OS9sd2jbg67niBsEelOgyuUCxhto4YUXQw6W
+vT0zpQ3Jcai9QM6yxK+zP8qMZx+gPdrS7d2C17DL6bPCS/+ijmqPOwzpFpe/LvL8x0meBksF9gi
PYvemDf7Oiwqfja7Aw92Fr2k7Z4KZOLmUUQWkdrM1+to4kBCFUqvwDgrXEkKuoiy9uxiSzLVoqR9
hfLuTlOAOmC1pVCLouJJcv9WJ3wgOU7uS+5AFZCiKzHFHw88b8G4pAD1bNVni6dpFk2NNsZJ4g+m
taKxKlMb2kNS1FIl/GGUxfjQlOYk77qDCbdJZ+l2S9btZmLTPwWP6fTHonD93E00ve5SQYvXby8D
JW5d63a7XF7l+ucAGx+MCQxuGEK/WqJmbB3+tN7HORjX9r7zg1sdLZhR+vO8iTr5MJsIE4naTgYj
fj/AszIcuDGUa7d1UAsjfckLiXPuVhsqM5hEdvI9NXLQuK4cSPYNvRkmQK3SWB+7hZsQLlCvyzAC
NAH6gDiOFKgMTGx9YlCLKg1PMUwtwhA0y62Yv5g6N0YV5lHqDVUGV0kt+A/zg430Z7KR3v02jeBf
yTtMRYwvJfWYG+4sKuecIjINxGy+xKoESbCnuLMuDV9bNfTk9DBnTBgPoeHgKzbAQ5WeZrch93w2
L4gM6BL+IyeBpEMPcZph3M9OhH8RV02YdtgnZC9IRRly4o+aEJwnl1uzW4m20RBOu2qG7sNi+yFq
h94Anrg0u+DbbYcfM0/UA2qcLjEtNA5uR1xdjLLLz/pkPcP5LhjHnHhLJGhffhueD/QenRCBMZSy
hevZFMzLJgpgVqBJsdseB9UEJmZX6/KuZ9RK0rKMVtvh8MqYFB8M5YiAPFxTWfHD9fyjJDdYJglB
oMxA3K55YonNYb455biSF2mspbaaXj2mVMFM3SNQBSAsFqrPrHKKE6Ur315A7xCw8wkxsRKoeEoP
DwYtGBKOcIwCtmfDWcyEkHYgYRsY468X9g11855ugL1a53N6UHniAD57/tEIDOupFe80lbVmmfNC
VKA63Av7gDHQmSRdutsBYLgVR/UBKw0bbfIAv7LddxF/LJAppVVNlf7zwT0oZUZoTSYVwemkEm5p
4VbwuGjkISXON1REhFLkN4kwEwkFU6b6JKD7L9BhvUs7USeGsvbJc4lksjPEYpnMhp3vtDT3hIYW
O2oAFkFN4YRD/zlUyWOPGJbxfzp9AdCoGaFYWNAC8ueZjFDToyZi+RNhf+b5YvXw8QjNetSm+QKq
m2XVE+WUHPIxQ8W6gAuG+jlnV2lBC/JjOUP1eq297zTjqvwrFNdgLlWxKZekTDnckvZnjw/z/RLE
TmxL6KrzeYBXuQMduQYgLWwtnVtd7sNIXAzXWvmVDHmTicfswBszGjuLtrWjGnkl3xKHOjjPeUXd
UfXAFmAfk6HtHCHiCT3QiVHb3Ypjn+u6HquDG+dhgSOEY767bREgc/9l/+55qEPM4yghXyWmU/A/
vjiwoxpoJK6b8nJq7WFvaZS5omTGVpUoQHJ+xRtbuATRdtW3SCGXQPM2HCyP0AXQpiYtVkMZtx0n
qTL44B58zisF181X2PtZVgrOCnHaCZEaeB9oUOpfWMqPJNdQJkUWn9xHzO1FIFDHBYJfkTceUvtv
uxE2WUggaSY5uPPOIdux/Mpymj9Kr7vNSyunEhEZ7GTEQdZOlWOJyjepbDmeclxvtZGmWBWTkfMA
fns/ohR0XkTMktsYSShJVQm8JZdYnGEqbKAXxKld/o0dnCwqK4EFoDLVd4SsoXzm2XCarZh4QvX+
0oOjog7MFY11Ux3oOMnLZQ1xoO+bvJ5AgQbvAUxZdjgX3ynPE5K1NQs3AVRKmxDjJrXddAXT+++W
I+oG/NZazOg+kD+RpyFZ+20qdZv/zab1yJlleMEoU8g60UuyHu5fIUEejhL6/Rlhow8JhvEXzwrT
X042C+ySmwoaQJkgjI7EeecEcW9nwwt+QDZ21bKtkBmJzV7QLorSdflJfsdjGxfOX0bPQYOEHxq/
35McaqjGDV0GbZixSjK6w1WkcBHhNFj6S8490pPMnKuDdGTUY9eFqAosizkypYgc7Yn5SYAVifla
WpBdnmegHa8vICFwTVRHVZZwmkstoW/wZaWFtcoBPaMzg2cu7gk72gtbTFDNkULOpVvlk7XYB0gH
N7vWP8BGnRRxaXmMRZR1HQLojgFyClh48rZK2DuK0LfjgFAuAczxu3iZzI6t33gPiqgVyenScEvt
QCfryr40xvzuj5Bd+X6u6m4TEjeVibvM2SHTEfeuxRAjD33x/fe9BGeua2Iwvx5PyXADUUlfEKT8
VWRM/Nc38/pvdxEeGKjThoCzklmvao2NRFHfE3sZ3HoDUsKwGa2fRsi+5S9PuTgMGMCwbgMWaC8O
/oUZIRk12NvFo+ZVZhdb89VH3zOlrHg9O8Cr7i+CGzLbGB7xXEUjNX4VV78pv0iRZsGJSp92IBkQ
pHHubEbKcPy5ORQcWf/wq/CngqkkjTkfA/CjnO4oHqa030e/5l6S0oym3gbRYKkfIvs1zC9Z940r
4pG/R/qi9dDyUmEp3YcoYTF3+BrM/etoW5I8h3gBLp/lY9ZG2pWLDLcntxx1veegqXpaBBcvXU9k
laCIgbNNh4k2KnRWPqry9HiO93vTzq4R7w5ruAT+RFB2PiTT+wixL9zxrTywp5guqcWhcrfyaHKa
/nERT3Yw5pXCEDSMxNvoUPa0fZD6jbwAQKfgf8yy3jS1kTkyhx11ltvFqCuIfiyN8ifzhUM8nKF7
QOVZvooId53Zu2rGl6vw1GQplSOnc7d+hHrHiT0GfSStW7StdTBrEUF2QZ9bdVcEfSFEA9aPfsqn
rDvLmuGzhL8njUXTpGWe8/shyxdCPdoLLddHq9wfto2wmAUyoWTk+gPxGVol4NAPLDHJanaOhFZj
yiSk9mhr/IHeGvDJwgrmuwPPFxBYFo2sWOCwLjbUax/FuMm5NG65Xwc5NEEVVlJEs3F0lsDg3e8k
rR/aYeMhOlTA1TCIrRxnPtHaKhggj/DUoHMkCZdaXm8ojOdFh4+pycczBACLKDDxtIUB0Epp5x85
Am7VLgv85a6huLam8oU2hMwF/6k+aqo5mAZ4sId/0yqIJR17UuTHhYOBpFZz1LZpiHuxvYpNyzWp
gbEfHkpMPYVWowhogA4QgftD7xMnuA/zJe9KYOQtCoSrRTkpCJcKLp+hI6JyeMHFsXhWV5xDNggQ
FgMiHKAXcn/1JSK9z0VeR7PDYOvyjkVcvKP9DWLo8SPeuQeoD2xMUPv0uSp4aS9JzzvgAauSrMoJ
JCxUq2uvG0+OnlKcahQUYeZXjB+qkdprSOCNvqNeAJ9QOlJskrVL7YtVzXjUDZS0dprLRmvhjde6
IAuhCsHERCQKH5q/1NrGx6J1d2pcPSFfMYjiVtGQ4zvfPCEYDARUq3On3QPba8DyjLs5oJfqDKSi
Ir5bKFZeTkH4M93zaJTsQ52WRjxJVPOGs9ElnMDqVtG1Vl4lQpFwP0XETqfhMNfw2SJWzLUfpebS
MVSwHw9jMK2I1Ss8gCrmUs7RSwiiwtFTiK6BYBBwAzmlHVd04EpLeNHmH5l7y7vGaPlBSm1Z09+8
ZrWiZ+4Spu/VvjKGDpJYJZumUmCq8SG1v705CsGINqph33n9e/p6tpzIm6McaCV5UiSXx5Q2jKWt
D0py4TteXhXT5lmO7YbpiBH4Gf862GwZg3mCvb7PK/wB2MblgJ9xdMDiijrNcEg1k4t4cdxErjvx
PlDjG01Wff2GMwngX3ZwwoIFxZrEJa+81U7wmS0Q6k+KjZKpdaqv3kLYtk9Y//8XZ7Y2dSAP+ydW
wyBYtC6C57KsH82Lp47eAZEl8A+x9WOhrIg7UZbnp9y41kfekM2+v+fxOkHxt/J7RbA3Me2HH1yY
p+cEEExii1Ndb9m01e/qTS8Jg58VrAr+68NTXC4jFjf2R2OyY4UrpQEyfm2EKdcpL1BeXZgkrrUf
Q6cvz9tShD2+A2pjj2tslCmQ8HSzccsyuZxpxk8zEq0hjd6zVMYcdsrc8XoKxOLMalnj6/Vsr8dR
60uqgr/2lRBfb6fkL/oIszOcHIhuDtGMRNrjlc7JpbI2AtmjYk0BMT84EMuvye7G8fWDPYay2Vnm
CiNDwbqjKQMTxVs6pFgIkhiAPVcKu2tsmq8VYVfva6eE7uquXfo6/CPmmey8YWB/KsBUkf1w/Hsu
QBaJrW2YnFbz59PLUaVAzyHSxPQBR79jQZvrQTV9AEpKntCksaLGS+FrUwqzE8IbGRcwJZVokAoB
iGOZwyGImdPh+HLBwDzvTnFnbu8eu5TnFEujs+qFl/q0w9cJojoD6x8Lvzogrfb3FaMKya4I8ByM
bBEUQc0sAfDP7B7nFk4cjWaDITYYo52ceWmJhHby0pZXQmQbbBwLocPlEY4O0jClOz22/YfXLRjn
ACJBq8ybhEbAUJZLZPqmnbhPgNsz80YSYsPC5WKgniFCGEKpVY0S/qTXvjOx8FM9qezLG/95vR36
nVbaLtyJomt6HM9pN+Yh0v2rUPsmeGE5tj0iLNRAENBbwX1chVbap8W0nTbwUMFgo6k7QW0hgtvy
x14pyKLC1GcCfq4lJutpQK8stpLP51aYnEmPGQ8w7aJIIB4k/3wq+3zYvjXHBdYrEVnu62jCbWFR
b0qe4N2DkmqCWV+/pB+Kqn1TXTIAlzUBaFzGY2JtG/OnIo3V6C9PbtCwJl3Do3Y5DlPxlh+cV+6/
JtaTf6l7BImPkiuyBwHePhucrVVrssda0NrrrcU/ngp5mydEYDieRQvwDys3w8+TSjlENdwHFhPA
LrxqRNbjqK5eFMKKk92dUVeRs7LMLhBfJowUra3idQAL8QV2lWFMW19CfFb7wr/Oovp61JJuCycZ
wJ9DB0CccrBjXkK0SHoaZsP9wPV5aFA8tU4yz2+wshC95kUOhJgjGKVIlcL+eUgBFFyoJ9DRpuwj
6TT/hYbnGwP6hm5OVkk+3PdtQUO8yN8RchzyBCwWeZ3uLAYThBthRUbrOtcXjIyTSU4YbBktJnk8
NXHdcyEHxqaCLiDL4TPwynY/iqbF0xHC4drw06goMgWy0VxUL/SVYmcCixe+p0QdakJKC3rs/5Ln
unF6iqaeuqaSNeRWJnzuFyZxkM45AsO2tLolAFHO9spC5YaUe56AWuedr+3kixltLgCDen6NlAD1
p/9An7yNWj8gsF1VD3FwluvdGtWavqd/3xWyya24cCZSl4W0RRrpDXhwyvGH5AbA1LGGILZsUItU
0DpC2E0PcGoaP7o8rElL5lwKxfaHgQqvTEGIaq5h9GIduGj1g+j86rilnkvMXonPv2Sf458M9IkP
v9p+Y4hY2LnY31wucnIXQCzVwi6yoUy1OBX655UzuPx7H8kiF9dBNTc2YMickGG1fBuG2rMqxluu
0y/xogBbzkZY4IZ9pFnIxpiRAjO7ZEe3YmZ0Ns8r0B7gNCZ4ZXl5SwGmQu+JGlUx/HJAQCAfmFBC
pYUBWc9QbkySvqX5q949VtG1O3MKVeOIVBoSLvVGG1zaayn0gVaBNTjRPOTbxgcRrXfvmXZ4fgSE
25bzqLLzSH068qrv28cjZSfsN7+EgfGroKn9Aw5hE/0FlbXEGfrNuEPEihAWYZZYlHh03mZe6GBT
U68md5pHSzy67n07/a54f5U+FNv66kePKo6t4ujO6BihnMO4FnlP3VC81tuVUV+bc9lR59BR+We3
iSZ5my+RzFJIV4DWxM7w8T9L8N36xUMeLqubW8pG4dl/tUrKV3Bv/NYSBGGo7CBSBZoHdsTHDtAs
PrRpLxrTN7LsS6d7PgBlRA7+oI9hWpn1QxSZ+YgpYyopZjx4nm0gAKaNqfGExg903iGiojry82Tk
no/niNY/LN6cmlT852n1iaPU2VFhKg+4v3UAa8L7f7aJn0bU8CZrijvAZx+Kp4/r9bWNdLNmWMYI
VTah84GFaKvJa5U5tGZflG7IYrlFzj4FamhHvnlMp1HOxdbb12HqpbqXkx2cG/Is3DpcKV6+bZ5G
IYPs0eBsBQpPYSTAJjqxI9QVhSYlSbPnHdzKIYvTkX6CzmIS0Lu+6BykLqDIt1YATbgMvewg/D1t
WqzH5XAPU8hl37CZdSqe/CTZtYI4WCmEOJ2ewnR2wXfRS5pJOTf8UurTwyCY2YGX2iB0mzhIlFBR
CgnmTCoJMHy1I9kfqfgxFXjmuWH4Ca0Yrf4UKU5OQ9bm21SpYlhV5zPc0RhoTuwqx0j11baSCevG
3tqJvkFw4I8cuq7Zgt/0eXoj466kOF7YwbjoxxHG0WW7zkMGVESZU3ghMoz/6N2d4/P5KutQmM9M
wUnd5DKa7XYIC+EcUBz0teeGTxK63SHl8xkkmv1dtVneFLe3rpDhWIv2KhZ9oGyovrV8C7aYRA7J
PKiCFqsTgdNDgmlf0QuoRWSpI6rhQsx/1hfBEi1U0n1mfGJwDXMWTzcYHXyusUJTjNaGyTXIOkC9
SsNM4vzeEBH/zWDwrdZsyCSKGRwhNdjLUoxbxR+JZcQlu3ryuOW6NJXO/rtofJnG6WH+SNuh/y/X
efcRkGW0WdulUbnGM7lW6ZkftKy9gNpIxzmIf5Y5TY0e553z8NnGrlAPLICKlgac28AJ/jNOQoBJ
vHDIxDGAiVFJA0TWwlD5B/85WLcYwhGBBj8PIY2et6YfV0MesG3B7wTDcf0nCx5iH6jheBpLAWXY
M3jpKslZSaLdeux3wI5xmi3W3bwHHIxBifO/IEwPHGYlZ6pEcs+XmB9vcUARASpSDjnw5HqzKQdO
YEWDco+MNqjYBaSd1tP5K+ySAzfETsVYv56k3UALvgZunpXD5Geh3y2dhbl2EjdUhaFMU8K6ZvaW
dnf9tvugYou/GYqUAPwIhNCldjtr4p0tSLz3xLUUOgAFyUXi81rxST7OLoT1j0RbxdI6CapySmSs
NO/U4fy5NE876gfJpfPtSETuOyZ8EHHeZA4iWh/QNT4AfdLBt7cT5whyfivUG/uX7xPmA/2AzzbQ
36+s7PdQDCvLaWRPnud/pyD1fwyTyGUf7vYYwHV58i89nUXqHJyTbVL/cpRKlMvN64hiIYYfSrxX
ZV36uM5Owe+MhO2z0QAaD2RY68f+LRofcSGyzk50FxS7lDEaQwKF5qMtHsUvTmKaRcoia/Ysrir7
m0dozv15FkD6F9DO+iIJrIhtcTqobly90QwFvQbFRpDArSm0huxVswLWf+9avPD2wMZiL/Ct0ClP
HXbDN5y0QEJ+tbGnZxr44OpBbqAM3SM4szP1PCAlGUF53bhId5yrvQ6pp0db37GNnqAHKHBEuljz
ALo0O24ztSfQo1MsHIDk37rkMXPia/1W416gpKIROPSZbueninncN00MvPRD+j4WDdlXUMBm1ayQ
r+OUyDaiJ5ejd8R9NEIgk9ZrEcNs4MB8scjJJPx2NJR3S7RNWPtriJHin4mLKQ6LELNiUX8iaX55
Fl4Aqdrzjr5gQ4Lo0NRJYoK4mUwVvHr/XWjRJdKhKzOBHCwoO95cjr0S+oJHFoKipX/BvfDJggQJ
OC1+BtLAEngLkPDCxOqZkiGAg+P3QjrlSSKozuQ1/K40hn9GOfVC8dekmG5IjbFw+XSddTcUzmWS
G8SjRATEBmf0ngSMeET/glEu8hj+oBomH1fbAmqBp26qM81v1x1jG8FbwdcCIMHvJsenks8dmUzt
fJbh+W2JU387RR536z3nnW4ZFxYTERn9sttUWrEjWFO/FDGmYDyc0IvE3W2ayikXrEQp8NFX2/dw
XN6Qv5GNrVco2nkvWFoKUkTDbcNGaZuf+9guC0sM/lIP+QgnNEKWdr7Jrr+QcOG+Xno3zA1Ry2o+
ns6tjp0xwDuHybS1eqCwS4ruBj+AIvUvzDZDfOYi56ND8/mDiFU0nS3NYxWeYxKKPbhPhuCpub1t
sXW1aCZD26ykjH77zA7AUQ/zcTchmhU9V2tQ3CTrwyv6vnedQGS8mE5SGIgVgCNDSDaJx2yzbl+M
OtrBj5/G5gieHjzHTgh7hkNSRwEBzNEODIWSZRHymJYa9tWUTmUS4+d664EKv8opgNnCHuAsQHIc
LYikjefDzWr06TdNikTrwO7oqw4eZ6sSwFkGNT0N7KfG26X4RPDrxJEZw4C5k338wqwKKsrOjHb5
9um7qaGPwjpal/WOzdMwiFqkrZgzn2qtexTJM3y852LQBJwb9m+PfTw2ZEOzNVbwpv2qd5m6vs9c
RVtiKITA3r+FPpYHWrezzLrPum0uqKF2dXD4vOlcPd7+S3B0XlGMhwXMIJyAJzrNbkmE0ck12t3s
p7sgUXIInJUR6bTpTy0JLv75RuFe55xRa9FKXal0gYtASgkvBTSfpHK/Tv5LWCSJd8Jd4DPzW5Vi
vdU8xWQo84tdvMjaby17J6v8O1/KJ7sNdQb4rrbn5gDDNFE9KITRQkWHw+ZVyudqdTUAdCCMOCAK
UNJJriLN2EgfFNUN/YC71UygioWpwzp90z8lieDjY4cNoARS5FQsafSaWljZVjSnMKQgQKVyhCyx
bHYW7/6uTxd49mV0wv4w7AnHOoY3R0vldLInJpZOaY/uUxnDPSpVLD5/vqmsSH1FIpKnZJEXJTyP
ZKSg2Kv9M9e7yeHhXdsWD1PrC8gHmQj2np/l7E/co+35CeqOyLuu95+szGxUvt9QVoDJpuSSI0Qd
4NLx9j89qHkNbKJGruhfc3BNiB4IbBu5ed1/MIUPRPiXnJp+O6JdSn1WujfWK90vauXNoEgjfbRH
prfPj/1SrqTjSJ0q138P/e1Hrjn87EKQUG9L5fyXn7KFY97C9/uFZzfNnbIaS0vus86tXQfp9TYR
cW42Ju4+j0w/KtGFEm37ljrQbdCMkniSA3TMkVXjxogcFO5YR9tAug6sZLWMicudAwluH2jEu6DY
ecccxD2Q3Ap98iXFCyLjuZwY07dzas/8YbPIsDnDtE+edLkANT4qXHVSpDKECXTKkpBvT6zQKgRE
8kzqfFhVSI4hS5+ZUJ5j0g6QzeafUBCHI4i2O3an0xQ67iQqaadwzobPW0fGwL1wmrD3NNhqlvHX
HIiGLEhoeUYVjusM1zmC4PUgrpaENahU4gM3NllKndDj3VelS6bChDZQhZtB32ulT/iAMuVnux6F
oLnWNNwBxYRQRnjr3SaH5Uwh9Qo3uFbhoIRTgDSUrd+Yca/EY6PSaVgDJ789CeP3eJbDDqEI+iW1
E/S/Knq3P1YhiuXWbuoxt1VoL3xKVYAZ0PqHSpkDDZz69uuat46u7ldX12NjCwo2Pa2ipHrS6KEB
ly5C20g63MwmvUtotAL6i/m/6/RtYnlq9aAYqf7HLvjeLquY3LHHfn/oe3GJyx/6wccr4LgtdHPW
W4IdXWR3216SMray5ndf1VdAAo4Q9KEM5zX5IrpQTAaqStuTklOUGDc9sMZKMNCC156d6/yrXX21
gvgiW9dv8dcF9UAulBu6lcp9zjcrergC1WkGn0yEflxL+n0CvJUXcwVBdW/DW+EfJPooYi9+QpbU
asuyUT/5CM3Q6mYtBAxAnnc650ZE7vYoGnzftLMZ2NA4WtcgSWV0TBeizU03C1q666255IKbHfoK
58Wn5nb7hJynkPS7mgGWo1FMGOvZqt3rczuTzEWsFDjBZs1SPRSoe+0iVO3MOvDjvA7ZJLhet4cA
AQxlu7f+jJo4CZpkC6YYBORh8yPzLnes/pvkyQ7scdsqmP/TQbR5R28Du4Jz6kJaf832VO3BGWHE
tB94LYCroY62hdN1eM73IgrMZOTWeTQBZpy1DA+EcHaOSDUGxL7uw8GiVoDAtwlfDhLmCLjcTpdQ
NMhMfpJIDrNbIAewf1OKWMlnW77og9xlzy7lsueIpUmXZthSFjN4Av37i9I2FyMMLd/LKf+jwZBk
vomH0tZW2y73Ly4SaPbdFPgqjt5cx4TrrYPhTMDzAC8gb6rBdd6pKEyag95G6sRJXeGL/1v/pmLN
C5EiiipcheBx569c1W6Be690rk1s3HQCALpQPSFwZe8o/0BlVPHmP49DRqKht85PSSWLxyGkoF84
W7lGT21N83C8zwPZtv23NvLeWObWQKfxW9UABpbT+soPj1JH19mza0CsCKepl4/NdUuvMpdbHjpB
vi9/MTudAD2QfMJ2VHJjo2YKTVmHM35W9h3fVkYrN2eXf4j0MOwKb+Co19TAuujc6ZNNA+zJpBAc
l01XQ6KxDaN+0ic5y0LiN24ZrCI/Mrdn4+f4mwunqGerHVgkjJj8wiGOEOL4zPKhakf6lWoc/SBs
Ni8kz6oRmIgnUoj5CKb/+qRyONoV1S6RJsMvrSXTYOgYkxCo/VtFg2A+TWIegSGiosc5lDEACeIw
lt87PssdI7FxcxHoSc+Jl4X6Wu8HBtIgvh4sJgV0s+9Bbunpxl334KALnAqCgrdfFt4jv2zONkQR
3QOV4o8+ZeYyM1eM3X6lVxTomG3P1HjWh7wFzYiCtP0Q1cBVji6RQOGEW0fPqVOlL9TpTUe+kFd7
Zz7Fvmv7s0yi+LDv2TVy0fKu8EQqNPdEdf8njTrXIqFgF70KNwwgjMwoxFNDdyw8XlW+g2cy4Pho
xyS0e64+FiB2nxwC26LvbSGvBJTDGrALQ/PQVXenffw/MXXVvHNgrp6eZVVJyt/dtX2Qx70vAlwS
4cC837Oml/IrB14OHvso/tJQzzh3eLuUG2tAftFvB3py3+WdVJ705I0Vpd2f8VNc0k0WFvpos78q
nmwrEfCLUoCusTvorbtqnpf2rVHjjGv9lGRVFNS+9xV95M0yG3cvpDQZ4vGnD2vmHhDXIT+kwtU+
9RrFXMVQfkGNDZMyYrxQ4xKZaKJWy5eTikJC5sD9/CiiB5W/AOP4Krx3+N72hRkNmVajg2NieXjV
0w1AdCTUwfSNG6l/h/2Z5ed7a+bMvB4unpeOkw27NcXUW0Xi4sOjDaQEz0Eypjj/KLH42QazDdqi
gxfg4eMKyyBwFNrB0i5a+V/E3wsQho/mX9Scb42AyAlLSL9ozDawKseymPG38M11jZQbuNhxD+6b
IGwBAJ8bspys8tEjSa7mqqgfKFiBRUzFjctLCHjzweBilEiV65Rg8Mmnw/kzgMQPWqE1YrqpD4xM
qnB1j8aEmhMLQ2OsDfMDXNljqoZLRO6eGc0bcB6dgJI3reIgV5axbUm7W4nmc+CipqYgaSmVZLLZ
ISjGhIScuvrZooHHK5/EVLX7/ay81JxP29Th8Fz/ytC5+LQdaoU4sFJTBamrJi9/Hz954erazp7U
pY5n1ClgPBvMQo05SEhKqQuZ7XCuyJnBndvZmuTS0Eduv/pitEENs4ZF35IIMXYKnxGq0TAMIyLY
rSv6YOuQidvkxLM/CnkMdXHhxYk7zZkM23RUd28ayWx5LHeLRVM5WQLuUfEVzjJziDIgaGIdgw20
yyo1TfZeju/Mxps914rTw9zdDz5Ge00lWa1sGO4nzuK0rtz1wm8s7ewY1wiHe7/BCf4frSTm0Hiv
N6ctwAk6/Ur4I3g59gNgXotvafZ0WI2J1G28UBKJdQbnNImdrk605lJErdxZhm/C0OqUezekTE9D
m5QemSoRekUpMUHdgH84lTazK1gHDzaLrvDnat9gP+UZlR7tket82DdtEbb876K3VB8nFSVZTb2B
HAgdmQAMZHbH/81heGng3ZYEQ/liQo29dr+NofHbcR1hgFJ21roTm8iqGphlTfo5WaSU0vUeBctn
AT7yXELFWXZlBrL1IGWSlZQ4Bv7K+doPvjoxOPbhSQleKrapsr4QHKyG0csvyU0zqcUKBJjHQGXX
3ETYAgECPgL434BrStX16FrSKw+z0+O8PNJcTATk24Cj017yLqs4RWip0c8QCuuTIALsgj/k7eUO
G9QRvIj2BprGZAWgLUeE13qf5ktoz7S54KlRtirlhRM9LRoXJMfUlpD2arnFV1oZ1kTXou9h+QUg
/dycGMZ83GDPsV487vozXn9JjvrmFqIThtLfClrHsIZUoqfynZLEfZ/mcddAxy42uud/ZN/jm/Gc
VrpMIEVpDuz2gT5X7Cn0/IPFJg6i5yA75DNubsP0NFIUI652DH1F5OOhxkCsEe3h1/gV/WA2ItMz
yIC5PkCfNABAMwX0GM3bc1J3XCaovkDgAd7HMPfQV3hR1tGLJePCO7ZpDquerGa0hp24BvkGYrnj
ZfaAOTQ6BEL1Pd/gr05rMEhA0TNlWws8zm9IZsvajBokOVo/86oRfqyFFX4kJkqySnQRJUb7HX+k
zF3h6P/ZfpEYduOqMyiRgk3GNPQaRnrjUmkbk0xo8dGEo/AJYWC9l8H6FwrGMC/IDD88OZEh4U6z
JShHdikxb3LO/Fqkg6X5tspDkzoBoinlS7DC0i5xtPJBOZU0/lHn3GW6iSGzCE42o+v0XJqbUyif
UMsCj6Y8XMdNMTTZJqKZNTi9TZDwmGlkroC1kNISZMvEecAA7lcRjqBSudU6IO9tdskEiScC2LY1
HeSPq2rmFtnd1x5+V3dgUIMEiMwkylPXJyJfgAbjvDu5tDYLM5wqw6DDGETv9aQKr7jbnQny1zOM
sdMsLGLlKFCysU3Z2qMx7UC/5xDKv9q32YSUATzKE8uU73jv4zAP1r16M9qRLitjJyvOMrn3Ryhv
BDAAIrEF9p4hGORJm1FkL7BcgdEs/QO0xG08RE2ZyoeqgPe5PTJ0cP0cjOz+wz7LAKbqR72HfSal
ddCLqWgN6IjqNrkUgyRwUePk3WS23eOy9Gu09qdGtsQg6akW6HrSDbS15CSLOsPKgP+wVr4y3Euv
HIDfG5QTXemltduF7MX6+2BK8ia5Dsc9ipkhzWb8Hv702HgCbmT1BygjPMzBxQSCtg5p/+Hc7swd
qA3CSBNQ9JD5uhFmalwQfJtetTutLoW2SEHmZ9hBVOa/qy+xi9gHt9fXJbFZmpCHUjfd6fIZXNit
3QApMFHVWjwsbzn4RrvL4nV8oplDZqj52/zv4KUSJl3xUWRznHE9vNBhrRi0SFKwsV46DTZzHhZ6
oXukUj6WA4/BE3I7T1grc/VYRxtj5UnzsMJgYUJiYgMCXK1409cgknyG+xj1Ej8/0V01iiCWBCXr
1iov/WvOkFPUkK4Rs5EpIL6dYrrF5pcyQnXow3z3h8wTK2Z9/lKCi3FtoIKJGVt65rDFfIi53nlg
ir4MsLgIKztDfxXeQ7q0HVpXMjKn4hpa2K9F3Hb1j1unYpZGQhicHwyPT1HyjHHLOdxrgWbdzBGF
kFKuBfSE1QWJEs/i2lESdy3BVCe8H7rYRqP1x6k3r41fJiLN1EdYUNQKpqAy/lvu40kxcSEn4DxX
H3CgjwWdhu+0YnvOBPPvu9+hJiNvO7gXpcUH1N+ltwUdQFujKfLSVP8Co14i8RvL6ZgROQO5Fuj1
E1DAdtP4iWxPFOqEC/8BngcXPkXhsWwg5i2FCT1B0VuNJ3Gw+DLUFeOq+5f3fnAIcjNmmSSBR+11
IWYyFaOy11gI9W7C/XGXtrpLVEQTR9Y1j/YMwqm9SqDkDGHVBcDAJUuoVhVtLoynBs5YK2zzzqJH
12hKhGcE0qZy4rphr8tHHW/Z/m5hS18V0+jhYGlKBhHuX9nMqg1twehcCDCwCE2YGCvTL6ZQJ3xj
heQKsX7I8nxSJp7WSjwg1JYIcC4FTd8/DB1oyfKoShzbV7FYIonTBukrd1O2/YAHdAFPNWZSsxSl
b5hkM6797LuTJ+y3U9LNXOmIkv5SfmoDCrG3y/uQ9xImK6TDQaNlzkDGBiuTEbBEHsNL1/Lxv0Zv
khjYxzs9cscdk3YwpYaxH4OGNjoJ0KJOIN3sbSplmy6v5ohTe14L/4GHHv8g8IQnI6uUxgpwS5P8
GqWzZQTdKyAkIANRYVMjtbZo5jCV2EotPe3uESDST+BFh2bx3zJS0zhX1PvSgZInTbTkGdPm8nH8
Wi88pD6VaRp1qJZrIftkuq/wi8qmSDMs7hcSY85RNXjnGDcAOR509gtCUOL65ZjOD+rAKgMu2EW3
9vX1+wWsr43kVUG9gjinGutVAHXyZdN2UOpOZSBL6JxorFSK1ICSEWSzacwXoZkA5n9hPOy+oyR3
HSeIFX+7eplz+kKh/JT0G+v085WI2jg4AYJ3WfBft9izWRPLKf5/9JCSX49HB8mve+zr3zRASIuO
7MtKvNAdvPbFAJI/5MH9xXhxsNXzMzpLcxjg9ZOI1/PGTFKHHdxUc24DVYrk8nxbipraKrx++hse
GmDl4vXPBaR7chVByhdFoV/oPjT8lyX+unCFFwki6ExSby/71bOm0ED9ohdTdTGF/Fl5Xsw/3Dg5
U6cZYChlHxzqYkzHgM6TLAYktWUd8KBBpPQ8L3bQ5Rw5ttoloBKjDrYW8nu9j8eyuIParChCg6dD
wJTDuXX9M6FzhrDQVHHwjVQIoCjz57cfyd+TMcne0PVeenAOlrC3z/xASMvn2dUsvYTIVIcKzUh5
P9XCiQSMIaqkNK3n8dANKT9hNh9iK9YnzSwCz+Kp/Z9kMlDN9Z25ID+WhQ5VKYA1LseTJ+mYcQzu
9kyudMor42IR4R+6AgGGE6ubiDv0LV7cFEKkwGOzB753aexnJGV0lydCbOjTYAyCaE78DEMLCCAa
RSKEth7aSGn2ILPufX4RXOYiHWRjBlGAvYBA461bSxGNQGDzR+75CqcedIjNN62OESCelXZAwlA1
ouqTQCBsmnCVl95Z8BelCwut2n0enXe+NVs2z/bp+Q7wJVtmCQBklpsJC6uY/VdHaNM5wCaezvmg
FCTUJ4xZW0eXlzNdnYUZNCRwXvwcTneHGlAwVfHy0clUCOZVGbL0lTZHFlpVRi3SnGwOQxhX09Hs
QlXqreEQaBqBKcJnURI4jEM4uM5jkS1IWU283WwkSox1FQGFkG4NVAONnT4mf4iNYDAIWS4pEfxx
c2TkZJuorrFrMHLMbiizFNyST6Umejwv93D4MeR2A2KdmbJTSggldNrVKKjuomwqLvnPXMw4GOcv
xk+ZcZQM1CZBxjNrB4l1pMNd9Z9avJ2aTI2kD5sREbM3/pKrbEj9XNY8hMZwRk6pYVVoW7oRER+a
+exj2JkTBl+ZqiLY1gBBhwJhvoo1m/vBshm8HYMQ+qE6alh5cBCodIq+PgbbhbidmJG6YpwxLkhp
GCz0GWx278NuplVxXvmGm5dysNg1Rk/3uqaEwhiJ77lGJkgjNmalOhckEsF9AK6MPQ0UaR4JBIHG
tevez+xvBjBReDzsxHjmi95PS8kRZ5xIGtnFStw2J5WNSU9gRnomcQkYZ1H6J90cT4X9gXPY2Ix2
EU9kupoyEkRHwS+c8QRvPvB1uVI/hgWLXI4OAaVVBqfFMiybbQ5mVLy/Uq4WtsohUpCdtCFRLen2
jwcUeSeRkOyJVw2CfisOW+yLVshYq2MQBz7aujJbpJGd7nwlbo5WAn18aLr3kUItiSfNmy3cS+Lm
e35xQ9/GG9fMz8IPCp2Q+fev46TaVTYpj162E47MnhTsakqCV9KfsXpOtwsl77rw+3ofqri7iZwJ
LE36f7hmHjUXcfMaqDfXSAzHzYryrcgJ6P4VWIGb7EYM8VHh9Ei6YDwSBxbaWNwmpAdK9HToQWmf
WH+XAK4jZRdOCfyt5FPM84V0tpLJ0IJD9CGIXGteVKiQkDXs3SBczoSLBPDQMa3HrGyq36vhtLVj
BXJHJtYPBNI2NwQQCh1anTRtXsvYOdP/qPUvjel66zQrXweRM4zL7jaaMmPRHCGIGSR/OWh8trQE
3E6RtMRIf4qRSPWrSbbApY7S9Gc+YDUPdrVPqyQaaborbQVpR/mhL4oQCswkOVT60umBPsYEHyPu
bj43UwfBH3Ygp5I10TI9hDbks6CZ55xKX24BcnDAmzm+dp+wVh6t+ReIqwQkuJjsvSV9QLFv/1Iv
gHDhqLcqDaU3YN7gjpp5NVCpoavT2yTvLJMyNrSuXrHsoPlVCfq/OB7n4GjyzJ1tOcPnqKDMb9vR
DiN1V+WmTwEFCAG1fK4YMzu3GSnKuyGqCXcCrXWG7iVXX8gFE7IGb6fBXIj2uCPCPSR5RBM+REeL
K8dJhN9+P9SH4sY8l3Vwa0/RSO/5Rc4P+f0rCo/NqlwMx12xtbU+tm22wEqBz3IMCZHf1V/H7B0t
HsiAJvRHVOePWY+SHcxx7MTrCHtKrsc5n1QK67KrAcKUhZ8w4X7vRZuuYfUC0bNdvBEBWWivdW/c
bFRJXCto8pPfBoNdoYRCU0Vavazz81OQerXwTZg9EmfPJDbnGx7lC+/wqc90MNoHYY2zDE8X3Xyd
lwwczqO8xBbdQbo9dwltUnvNaAiQgZZabbQOObbJyCm9WcUXLKYAfV9ici6Yepyu2/599+r+3ZBg
E3a5K3HjmsUz6qulYCeq2lJ4GdbFEDEf+fUiFhvt/ONYHIcWYFzlJgjKfmW4CPY6ZBj4/m/tJVYF
gQA1L+2ZBrOgOQ0X1nLrvyltnXz/al/xOGCT0QMwwicJJ/JTHFag4N6nege1Gv1kDePqrwYoHktu
PiA5o/4leBqcQeSPf6bhUmgC6lgiPNtgUuLVzJh59Ey10U4FlhDPFTyOVZ5sZ3Nb3GpG3uaYMCFj
XUP0IfYlfL18FtREm4CunTXhcnfhgrChg4BZ2zLSQiM0343zxcVQlGl/qBE3TkO5rpRj4YwX32ih
LzAJ3Uf5detu4fhJ5yW0I9bFO+mpE7tbSLB9IyKtkvsCw4McpvuNzq0i5weKI5VbGypKtr0ITwdm
Er3DxynEAy8c3wl+grFvA4BX5KCPvui7+n8A2jYYvwu3nww3MBi0hWw0jgJMsG64F96+WsFe4wzz
PWDHi5YcezXsITfZw5FdvrEdZXIUOXZ/NmMhmXBugcOFalO15vIEcqpD/IksOmkcjc1Zsd3+nhUM
df541rre861H+5qKn007Jt7LdUdSGRjgYHItptZGTP2r/5iYOaC6PEZkjZW8zLR5+cVW6Sx1oyHz
l07bxIdGyHY1gjDw5pj4emzizTKuJLFJKvI1qiRva/XrHo9SiUWZaGcazP2g7lbStHbkXcxGb/nC
rbfbpza0GNI/pccvO7l0I/xFIBOTR4EMLr/9U5iegIVfOkGaSs1fIYYC3ELdVCEM/uRvCz/182/i
Z3eT3NE2kNJ3+75kg5Pg2QJWByfGyE+uvxQFNXupaoYWr3bdYmM/NbabOQocaT9LL1H/tipM/FZN
UtUq1/SAWwJOsRfBotz1z6xe7pQZ6L1uZYFNGk/5wo54vRKYxU/LShcXmQn8fSJ3yRYleBjdyAYf
APyQA8zv4RVzoP23UjmEzhZZw5kNSKGFQO69zjZQQ20Ksjxc4aWik/xh/+76CvA7cXTIEpZXZwkX
I2YPUctVMpn8wdxmP1GQ6Qew1YyD0ZvPGYvxCRlRBDYHZzYaisqg7bWj8JKkf3pmyy0q7iNm1bjF
nJOhXVfbOgWT5pb3R3QEQoLOwSVKfD7SoY4I9iJiECtKi1SExfHpPYb7Cs5OKdIiu9OyJo05zT58
awy2yVmFFm1r5sJn5DvKxqbm3U9ChIg5gan2DacHOAmRL0CmC5f2O6T7VPytP/ltNiBLtIo5aGfb
0t9+uFz1CWmNCIxgirdoLnz/EbRcXtXgV9eDu5V58aRyGNf8JUeo267INkNiafDD2gVHdHKPDsHo
k/EFGXh33EdcIH4+AGl6VF07DcJNs8e9dkOD0ZtvyrJEU4JFfjnGScxzi2EzKJxr48C45LucJAj5
FKwt2aphLJb5vKPAe8uw9W9Um4D7k200bsS6cKlJtJOz8jlaO/1k48cnjDqUuY43YR3XXae7wrma
iinnDNpKM+pmd72YEM1iBd1SxFAGTv44euLrYWhEos8sIRq5OZ8AAwUBmPloFNFeK5570xbZN2w8
aqHVk7ZiQ+qrLobK0P7Td3UQ4Kd4oUUM0wzNz/a+d+lugjTAQilHOTW9c0bLE99DyGSRSoeDHKnW
fJ+Eq0np1cWqxhelq6kTZA1Zfq2L7C+KSI3WEqof1UCgfe0Z81pfWhzFV/8vDRxf5gq+pCVQxKBo
ocD0jLzoFjGdVaFPmAIS+7EML/VEjN689K3i/Qq9XtblXsyPAniJ/FSrgQjVRk3cEy9EbVn3Z1z9
e8kLFIIzjHYAdgpRF6+16E6JjAz2sS6cyLYVyHrwuFADigwkgiGM3O5Ljv+A1APYXOcdMO7/+RA9
V8wT3mhTDR/Zg0IUzskYiKX5v+JDi3XUmM121ek4T8dLIuKd6b1eilolfwnbbt1MrsF/VvUgYB1V
4QpwS5AFEWxUDGyPuGHV6cvQVeZ+gYuWzQM+alX2kH6pzrCEGOS3M9Kg1khhRjNXyQaM3eKI9m+C
poBdULHGzBfLNOrjbu3C7VEEe3gnFElEdXcl1SDy2g81rS6YZbwK9MhOfEd5rjG2Ac57IZZ1ti6N
wyMv5GzGX5PqsYEFdqberuWlV7FzPIpqEddfRxDgfIsmKtU4PMw/BnbBsSH+3GeMVgcVZ3bAELuY
fV5TQHaXQGbhVJwXaOf/l2VxNcXF73MuFflqr9PGK3apTemDhJnU3wDBw0muvKsP4CU8FztDR3SG
LvO3PFo+AQPWcKj03w7GoqD0MFu8kIBXbQIrS6duBe+ktnBD0MVElmidQ0VkgqPJ3xQ8eVk49chY
mXgcozlk45JxN9Zfk98egYhkTxyi0UTScHvZt4iD7jDwStwXEqZfwpkwHLag5Spx/W6DP4pnaTz+
dT89FlpGXYa1v1rpoJleoaedpEmgycIvQH3RpdMtdJz2itOHrDhTb6y2+9Sjvv+QYI9zVXu+CwBq
VazzP/SbRFTK9nYK8858ArV4bG4XvHEK/HmfdQHpj64QvhPCnVWHwEz/CJgOUEj6N9TeNNh0sdE1
9PSfBHCzBbQzQz5SKCcVYnBRUH7VRGX8DX/Ihb9eIcKGQ4VoN8/GLeT4LargfAoNHozdEbauXYKZ
nVDJrpQNcLfTdq+zZDiRdda94g5zDcmeg95h0ALinyNEXlJEwVduMKwvPR1gAtP1LBoO2xvoWMJs
Lsoz0S3XSo/dDtQGf6iXUEpDD3gCgZT83R6AtaUPI75aPZN8MOVka8vDQslK62q8uVNmalnOFLWh
LokDtjN6IKiMWHEiNRHGZJmEfxF8kURPZNXgnEZZahMlCEfEH1VhrghxJd5iyqTFyXDKlKE+bpKk
Ahr4pQ0bcEyDnuBOTQmYoDMtHI49xmIzCUb/pCbTTKHwcnHja4eQtxf9pIqh9xwgASAkf/3aUmhx
+9UOJTU9JkINq9PXagwJWqtuI1rVhLXY7HyAXQmGyRDuOFpKL5l7P6WMwS84FhEga5jLimTvJZLV
b3f2eBFV3LoYVxQ3s28JUx7AC3DFU8xQ73nlWhKWOvI1A2uPjBSNC0OC4csTHcMgaji+C23mpb3e
Q4EArB2lLZr4zJsAdlj1olwjQXG8tMhvhzFIEkac6FUuNWBUFv/pw8hTdwaRZVwJ1/PFFiQw7xnW
P0SWxUiyG40IZqrLzXYga8PpJg0eqwJvZxqrLWUz4fniuq4YzikWUYerPuaCPXdT0IolDUUPz6Gs
owvNDLhsfzzO4J7KQYS/XEDl0a64cmsZPTwq331vuTRWGLD5cKnKmJMAvAP756Jg6yHfvgMbkUwW
8Psg6IL+Sd17S1Pj0W3fBapA9XQ89iSBZ5jqB3Ks7jZXH7LwXzqvDK8ths5nGa69x54uERccT9eJ
LUJzRRYxc2lxNR3tAr54p/T5QayO96qlgzKXNyNHIzOh6FukRVU1nkt6w/bBwSrWkaRk/Om4eL6g
/g7edVFrWaBhT6gPzTWGcZwGYSZqcp11vo9v66j/T9I0QCJpZHqHekwGw0pOOrWad/uQ0mb0zKLx
1XZ0rZgJ0jrRWwxLpdpCd3bcI+QeNDZrU5DYRRlMcMeBk3Fs3TEcqZZva5GLplFRqZn0dSOEYl4X
STRhCbHCUMD2u2AAy26IwqKTb99Qww04vflvnn+JwsHbxufqkj6oJB0as5n0U1GhaoWRLGG89dSj
naPG3kpfF6xelEIIK4In257NmDiG1C+udW9yA+KIKsU8qxs+zrZq+y2MWoL0yH9spmZPKRhkf/mR
EG1eXxgcR/pH1EMtPk3w2lhopQPOabSxZfPmzVf/uR72aNeuFNlDJXuKHb1FcgcNqPxXGSst7bb4
YRedM+kPUuHEs3VVsTva+X5AJDnmTuUyrz5OgLRBvzZU57/Rw5luuWTjpf+RmVygP1PyToDiHpil
X5QOKsOdqCRdjU6TpBG7QAK1s1OKxoL2payEvy7xptb9xUj3HL2QyqvQgozRcIUVYtg08uMvCUNA
VAXlxzxQMnzAw1LP6wDSAuGD7yeAGOuGKqt7CCpyUGWsD5xbDE/s/fQVOvbqW1EZ9VJhry8ebCaR
qSW73uDTe7VvmlgTnjUuvYxpXcZu6UfVxYp0Zt845VPC3TOq0CdQ6xeIRgQghZoL9AbehJxvZ+km
PrzDOeku9+SEHcCOq2IWhSuW4NYfUZ/5gi9bLW06AGpKsfjYc67UQ8VkXo5CDHj59AyCJKMRYPJI
ETVo4oQSP9vwsS4jIeBtEXCb+ncP6eNlbbo1Tvu9IdFBp0C696KjrD3OyrFTch2lSTW3+lWrNFBC
SvEo75NPE8ok09Tqgi2BUYG4CnVGXLCZebpPdsgAi3QH/DnF9YTvMcIip8+NnfCtYvCHKiuMDvyA
8xA0cSKVmU67qqLs8v+zNnByCCjSTlwj5smaBmf2wRYZyjOhuW0M1kLqKdhDEE9cbOC8EgJ+JF42
AKDu1496VV4paHmDx6Yl9iR+pTTOKPf6kNY0lUQ4YLILSLfgKEhv3FDPQnTT/e1uYfGyxLdmDM1h
H2MHb1nDwqpvc+oJ3qmbQaXUTKwto4V81sPRUULN6bh8lIbmWM6k7r9rzmQDDbjPp/S5IN5Dhl62
x3PJhK6dAh+G2YuXAKq+hbjaEgjk2LxmOltuT53h36kBLdJNJrciqRSR1xq8J2K2wxtQPFoxHPKa
CIFVND15Kp+C6QBhQcGkaP8c/O2WgIjjv1QkcE8ZOoIA0t4DhN++JKW1y1lKUBXU9BANcxyS5KiD
P9qpQSbkNKKHRGDMe75+GQ1ofQ1gIFEkj3xs6bztOZZj6EEDU5FmxSOMY2+T+3OThRp7939aarLR
EbpVg0MtqOtp6185WfT+K+aS189zot9oEvfJM9wANTYMe3AOhHKQJEDr78AlFEx+f9UTEuPn3iOU
aG8FMeuuiiumwk5mootTLl2wcAnLFX434JTwjFOS5kCUhVmcwr6uZBeIbp79+dv4gT91d+em8arO
/tVEjEOwDoUEGdruxCuLgfCuVFs7pIEHRrITz3lqiSPLfOCNuYHRTFy5rck1gD9JmBLIQy50hQea
0/nl6hDq8bdSzRKxOBz8KR7OkBdaapNA2JIqu+h4SxQOyoPL48GnvA9+knJiStijy/ec8MkkK+rL
Gmpkm8ApUtr115oSrh19+k2Nobc7XjKsBxWiwCpV6E/ujNhNcfM9G2Ngcn/Y1fqcxepRNFEygcRL
yRhJXQ7uTqSVVHH3vwFcWbUT51qyzkaHvZGJuXyyhzSSX7yl/A0ZrULQrK1jyfpvw5EUbiSeagC7
4FhuWFE7baiYZ8KESf2GR38ngHYGCFNq2z84WRF4v6/cT6SgWMCTk2/FyQis38BnTZXLp2t1rvx4
XshayXtFOhYm+Rfj2Cu5yzwOb7/hCiFMB7oKq5Im8cXOA9nC2F1rVGr5tErFMwsrQLkHiSjm7aVh
hagCdAkGaIWcKII4BzbXJrTcXy93DS4pqYrnpCOZVZB2xcObFasIm/yKzx3qDAuPCFRzaA57sk/N
091dauqY+sQPoTfwRDkMr4MIMnYZUJMbOWSoHTCbSJiM+/4UnGqZNGBLy4uKb+ZSfPZrhxzsxCRP
hoTw8Eu83DNjHhTbAnRyej1g1fNNNxA7N6vYOxlqhpB0BwWHpqc/u3RBbFq4jA+q6p5jzPIlEjxC
+S54GqB0ATiQTH1WD1k/oE1IjqoomL3uSB6YoX9FvhKRfQieTOOX5DHC5ut8Jx/+WQtKFDw0xLWq
0JiI352959MjV5Pj49cHg7DClhIMvMzOO8seMKmmT72Yf8EtctpAXoJHAqUifyY6rCrjolxZsUo3
bJtUh07Lu8CKre0D55lxvczGv5S8zSvKF/pyC+zBhzMCFj4q3bxLvHEzvCu8wES2OXSXR/L9XMTp
acklLkls3KbDtffJi2/DYp6pA0MmNJx4vVUmBPX8aa11Dw6Rc5oLgjASHzhnpksIWPNBveNvsFkR
Mtd9tEUBGpdU63N6VkHgm3JnQnvMNCUjnRgkCHRG0jB7z5GLYuIEWLGl/NKWrJtuo152ukBsB4zw
pXN8sSs+tLCt1ftnNqmb8U7GZFW+HDDsiO/b0tm1kUxmTzdA8RloTP6sz7APLmMEHrQSwmw6yG3f
jEZU0SOQRLRsHnMMM872IhbyfPsYPvR5wI+AWksvMzmW7u0lKQ3eSyYFueMWEbIkvFKH0IIN/3TO
8dBZjMKpDP0incu2JHJkdA0CovnX7cufaZ+lRBUxwd76YHkWoAMDogct6JxlYNWPyVxYTfaURFx3
X30eClXwQ4CIC151bKEJijS+LER78Ljt710f9vCYmE9VUie1j0usilEq/TOj14m1BgJoN59WidgN
cbA8BlymJg1s11WYVBkEpIO5uCqQH1lci9+NMFEYbX1gDsyzzbjXzkUq8EkWw4ev0cInfyXF8t88
YTGrZKQI1U5ApKb+uHGta7rHhUnH2LXb9KTnxwpaFXN8rcY/uW8fZabZp57wOyTqbMfpRo4a+aPt
dLvNkZ8wpxEbHJrVVIW1L2E7CMhpp2Rk5H7qe1jGR6hoVOjiV8tm1UMAb6Rc59cZriZqqnYDWogP
l53rpTPcCSp05DwkVy6yAjIXugZRtn+v0V+BluNCtdy4m+59RfEs9RAaNPHkcMNWggnvmRawl/Fx
Wy7S6P6xuIsL3/GGP6+7bFWTDeR2Clq09hNAHOD29iyHHwZetRz66mt/+hmdiateKDy7EPP5sQQ0
qXjdVSFsAuUTCPlLT6bKNpGx/R30tJp0xtuXHoi+RQCzlmy94yT+bMZs6H/1Z3BgxlsLiY1IgPo8
uRYxg4tCnn/mlF5gXMKqWTqNBUR75plp0G3oqsfyEDrwF5i8OTKUAcXGwlwMeMO++RdRiMdWw84B
OeQ26/czenwkWI6BB8BQ7JggXsPZf5882kDtKRe1FH5oXHFmJmpVV/qpwZsbjKASsOc+AUbOw4dh
4FG5CBFUUr6JlOkOvztlqkMAgZBGN1GCSxEK4xROAoTATEq4J1l4cIP1AIouX1qkgxDg9Q5l6nSG
+g0wDxuqpK85DMOimRJfnGa9h39aTBtyFSr6b6EE++VOL5aniWQoSmBPhu1ReexXSWnfJF4REtpX
hTpENCGzJU1yeFS8ElaQXvZHw34HpIff362fYDuZ+wibqM2VXouYPU2A2Rfv2Xzm3jBnWtMOGN/Q
J6V8IaZwIbbYslig0jIZc4zMg+iuVscebIcdJEVkheAkyk2+fMQT3IVtSLD+PHg0kf+PrOLKKxnu
Juiiuw3UJ4CcTo60Jxv8CWXowhHtHAoMn6peb2/Zp+F5wbCu1ZuNEZZiS7LecaCPsf5OIqkTvtEF
sINwOnGzve0OELZfkZNBPl+WhWugWt8w5RM++6dvW4NtY8DjQ4cxd3zxAweeNpD5myzIle/OGr1v
chZgEQC9j8PHE3GnPyRRxWaOgsNkFik8TZyf9DjSwtdq3Wlh9zyPQHCiVOpRZEOvTZ52wy3Xwjb1
lhLgWolFkUt///GWa9Kdjat5o/k/sXDD6aCIJUiFJxwCFeJwX1oCUUmSFWnZ6XP3pXbgaC2l6eVp
i/JuLsR75ArElTn/cm7SupaOG8l2nVsbw0njF6pXb5yHpUleQ8QhZX6Kq+G5OteBp8j2rxXX4MCp
hQ4/tHjXFgxw/AC7YsrDN02U9io7LLjsDODEVwK4pHvnEtTU/vKZEzBn1uudAIIEDwR1O7XLWcNu
TGgCAs3ws1zonSY2fUYsFcn4620IbPewHiZBndJyTHeo6WUR2GATPlgaPJGRyjXsDimMb0tOW2Iw
Iqc6zSslBYpjL7bAjLsslXuUJH8/SriIblU35+kPkIIt6ZgmMK8Y8iw33JfSaRsAILA3nk4tT/lW
GZiVbdqiyVCxOM6XVkVDOFDkE5d16V5r1BbE66FYvSY4L+wVDTML0SknUxoVELgiOrxdEzG4/cXY
ak2FZf7Tr2GhfJLR9KdW0D/E0nNRbbMWxl7Mf7gzifoswAfwmiRrz6F/aanzIVV+BGAqB8BG/+6f
PgH+PozO2o4rUSJlctJfUyP27B47ytr7rQq40Jmdl3EQJvkTXXKYiagiDH8PVOUqwsLjDCa398Np
n8mdKNW0Tm2s+KnhKmV7Yd5tn1qikF5updr/TVpNxgk7ZaM42tVseq6x1QtM34NZx5JLKecfzk9W
Vhb49qKVv52vEB4xEHGja129cYrOZRBWF+y1ovF9VTV761RFQD9gHLuBlmnrAmuPUk97jwjIapvd
ieGJFurZ8XL9hFnK+UQEywueALFRcrpxppL48Li2t5kRzu/04l7elVrcWYtBq1oiPBQB5N71h8Zm
pddcHjtsHZPp+RgCZRzymVVzFVRjIgDG1z8rt1R4XEl+T2geq1njdsZWJNht1JsfNkLrcP7kPmYh
hdo6PWWrPurJlmknkPTQ7OXeKxDe64OFyOH6qFLMqJFeSdX6cpRo5I6P9V/KvgQDAFsOVkrAcM1R
4/vDtQMktgv+MDUni+gDZg7+UjH74lSowI2jRtxE2WlQnvzRTabMQ1Ngq6XWZKN71vws5shB8SdU
U5vhSvvUfSvthOvTarmatCgIM8W0vXFpjf8SBrX4SIK2G/O32cuM0owCy6oaF6byMjW41KbHbGj3
1Qum0p28+byZVa3O8PJHMLArbzXYMsJyKnqh8B4Ah2rj1S8/Y8rXMR0IrWEvehWsS29zylR4dAPZ
u+CaSKa37bd7ddLZLmUD7sgQVVVE0iSbn9Utr5Ev+kIPbBHF1kTjJ4IHe9Q6thxiT+kvBnE8LOpT
UU753RikRZ8o3buqf4RxEZ2LwS6siI2dSTFtsb02mgwF27vh3iBLikqHmxs5KWTt3tSBtf/CeN3b
x7lodj1xq+s/XesnSpnXPxvGmJxxxsOMnFyIE5E9g2rfnK6VsOIvFLFbEb0rxjG65U1+felqlyYh
8mSg45Qmyiu2sXt9pIe70UMlrYPXNckoLSQYxgaCBtVTrfOOkDaFWzyXIibfrbdFrtXnMQnDe1ku
VDAtfNWIZx+iw1M4zCcljxpdCUGt8OKE10CU/RdnV7COm8bWB5XJnmt2xL+0r4Z1hW+ddIN6OgcQ
vCsD0AaepVzV9rQ/DNHO4WpPXFyhYDLZE/L5KWZW38MtBELRx0aZVLNuE2H5b1C78GRDPUyBb+TO
AE1ZcqXZDz911oTWDiN1pfxuahAURs3zeCJpSD0iaG5YjP6/5JZNzljlvDkhjgJ/gigRmLax6jyw
pqXFZsm8zzE51hNnxfONBkRzpOv6BuQfvpR2FzQxC5cafo7F+7Ln6ItpHBXkcwweThwbbVgqm1dZ
YDHwbh7hb4S1l+KcYASkiQRlOdDblnH/jUp23B9l4vgV3M34ci55wFRj2pPMlX6u9uqjo2/P8djq
B/qZ2XcspxaBHFG/OhwXELRJAt7G/fFYC4YQMD9ZDkRVL+XoNaJuqO+uZqwJGV9GfZO5nPfPurTz
adEfcOOvDghy2BdezaFfPwb6ec3A3dbhKNNvxDX4nL0m4yGZ/JPy7pelD8BU1NFid3DgxDDEKay6
oDmVbs3/uC0JD91gU0UnXrOLKZS/o80UdvZSwPgaE71QgYDUUiigAmyGSkU7LGggQRXtNBGoqLmU
Rp3ki0OLo3MtFLq6KObcJag7HABWUH8/78WhoZBFQuQk/8kTS5ZZ9HHwGzc4gkz0fzNj9tvJYOi2
/Jj6N5JyJyYzlOm+k6MqheB86rT7gQbjqPQmvBoiTOLev0R4GnBVmxILa3osp3orAtVNbi+jxZfX
DxS0HUxRa80hXythvC6IXuDBHTcC8vH9VmJn5RIxeGBvnezdHstBbuZ+xl+1c7fpD8+If079Xb8Y
+XwtajGVGhLDPA2rVlmZQDyxjQmIJ3CoXdATAej6uI6ojjz6Xlm58nZGDa/FKTVJOuFMjN6bBANX
bu58dkgGOcA98tiGx5jK7TiZHP6IiFu8rjw9oTfCdKJxo5j6xuIH37hxvW5PuRn5DAsfg19r/Lmg
c62tVdSoKBuiXftY5z9iu4y9OUmW3LjsLf8IBlXLSPKr97D1hGgj43WCgUfs07BTtZcI3XKp9okE
anYjnQT65/wbavtL48bUrfl3RjDF+tL8XwkZKvih3xVb90bUyDFag6phATazBRSCQQzXHXHnUp1N
CDab78N08+t9qFH9NZKsAjgrvMkt5arbiy8ykc71Cx652H2VxhpSz2KKUX6OdFQkCL74Adthjbc9
uFAbkHV9I193TWLlbRU97FC1Jwdmk6I5KBY3lV3HhyBlZZDnVHfyDitrkCy5meFvBg5i0wyhwfTT
l3siuldlhC9v0dbnzwo5Xc94XF+AMZgvn9QU1vf02QTUNV4iXW8VyOaKkqnh/ELH8ehgD+aluJU4
88ER1GZ1sm2vjufN2TMC1n1qy3fyg0KOaOKTDWMt+axPMKnKKe+3Rnabp5cm86m2gCfIcQB5gIjA
wGIbdzN3j8BDkuZr99Kq7N7Aiwc08S0lyLV712cLrUpKyZrXJULaWYOVXh8mYFi4Attvfa/VnpsR
RVsDLZoyvgBRkR8FlU70rCutnaxWLdTBtBh2E7Pp7vD1brcAsiZYB8CyZuYOLMcYlczMqRFq+Xqa
NSqjM/u7WV0RVEK5ixkAusfmOVQuHHgRdokJ00GgB3Nfs8fVB001vn2j80vlZbU+BOwFARLLb4d6
JT8hGMmS7PASd2bEPuu6gRZM3zqczrvy4Jx9mT2pc+3xDDD6kZhznu+cXMdd24NXDXPUrntQAwAS
38YJZw33tJbm+G3EEUiN2I4tYRaPGnf+Fhgy+B5yBwQ9qkRY/YDaLZ3Gc3cMC3mSuo1d4O1xR1mK
skqsDfUJGKc6XxSddnA+rSfC1nI0KqqTHQjwoFZ0ljkPCXwr2wyjZ6NB1Jv7nONiA9/WJ6Xlaz6d
eEYzeEkFbkDaFJCxsmzyorM3P27HCPoeUDQkAYHIxqfocye9IKnHQfcmY793MI4qdss3MVdvSziu
eKFCHBW3YdmRT+tMjV3mLSoRStagmWH3SyDSfZ0MzJ2h2SJ8eZvfIg8oEVGEbIlfyUH2g15SRdVN
lc7gw/jgdxIk9fa1++yHDB5r/lAUHm1bqmlvPTdFmbBksTk5ipcWNp6s+QclBwN3HBtROotY0cCQ
eSplyc5fnuSdcmpDWEuxhR4KRlhEyJG07aFrgD1n3SSS0332eBwuqlUK6US/BN+unvOeagFkzXhE
8Wo2T7V3n2wWZiUwkJC2uFaKGYXFvhf2Hl3N4e34YgY/SFV5XYE9p8PRNs+Xik4RT+KBkbiBvab1
5mF56cTqP3oEmebvGIJHjA2vMciB7+zHf25DLi27do4HTOeT0iDgPhwA8d5TkQr9xes3zprLH3mf
fUi1XUQ7CUjxENzOs+eg5n2XRAouNHrjWnBQWCStbGjAqG9HnmMtvB4w7RaILWrnDmqwJHvjurJ6
cusXELZfnprxZebt6/kHmJCIRq3FJUtBzfsNmRbI5C7JgQShjdUqETtxjcjmo6zU2jpEwt67bRkh
t/dGZKtryd0ZBvWYiWxMwHvpoUEjPyt6/tl8lp+OXFosCrLKMERnw5SnH7pmn0Bfj2sn8QztUIE8
ZdFqu/fqWKwaFL4KncNpG+KTK1hG0Pdh95ALYuR7Au1KwcY3S2CHRHQ17FyAoBaqVqOlHuWk3pj2
u0AXC4J9NtS3+/pSe0A2yqpNNLTruGWIlsspFfdKFrfWFHhCWPpXaDqTbCfFuW3CME0q6Cirea1V
ZXm4GBM8uOj+j7lIR8JdZuVBE2lYtoSN1BSKuxV4Hp0+JTHuvWxRRKThleGLczkqeGzlhU43lygx
UOUa1zEQmCg/ZU7lI7RDPp0nGn5GbW/wUcY5uzod9hyaY9xRwt8fi8WYossnWGnnYTW5h+HSpONI
xElydDoqxnLr181WK03OEUQzEm0/NtFe8cC+V+31UTzNSZG0YiZDROk0H7lrlbeoyFcTj5IGjobb
kXPzdUX/AlLOgwxWWyj6ffiJ1m6uDPr5S8HssKvxYE2osRbEp6uW6WlLJKteYDuj5SM6NGTfUW1q
cNFk2Q6evS4OT6ZH5Fz+tjmC9cmPs+hgPQ0XP05swpsv4dDmRFmokon7pslrCiZS/GKd7uvKE48E
LxLwGalhjZJ9jKIyFZLDBred5LWSyBHT0ORTX2dXx5HLcH+RbDhwoLS5n60mMcVVnk0k7PZqVnUz
MtVGUKKo/2MYiJBk37rskQFAFPlcCsZqHoypzRTADDz4FSUV1C+Vf+dlAaprwhFLTYbL+s8qNex2
ZipNHd2TZWaoDtkQ+aq80hnZcbJFxebr9SRDVAXY102/mcZI6Zl01XFHr6Fw1aAIFb8MxdzvzIcB
xD1QfKszpQ7W1YH3MpP4edtIxaS7Pe1uEQY6PrHGsybZ0LNgPuKkgHUIZGZB1EgDinAfG+ioneAb
wAPLc83Yz+h/fmb7tlim5Kwgi7urPPMkZDrTp/vFOZZhPpypjngCXOsab119z/I4/7uHKEI/DReU
1L6rbYWk+kvM4WUzFJXLQZ3lnC9IGlOLXyGOLKmJVHk3tNQNUI99QHtkcCzZpFzFy5L2BY1JwnOt
7Hroz8wwRSlpGLm5pfaoWX8pZYgQUR/yDnBIE0rYzbWVOVvQwh7TenZCByocC16+IkiM5gsCqZeM
FFjoJhFkPTcIcRx6phhnyEENeRYFeRrrpfrIR+T7vKRL5RM1cRfWiH6uJhzOgW/dDTmVJmeO+cQt
GWfod9RrYcg/zEAIdLecdUKG5Olrbf63A77sMdq6cZz0/zTDk8au5NnAd7Nu4SLZKMSgCequ8zCn
ZzHbbslIo9kK/+qfT7fdggKemmfoIdIzJS8CGPW9mJuxShwfy4JKz52zWEwFWIk4P4js9Z/yQcb4
dguisvD2nuqPzVMQIZN8Gg0uWPd0i7Awl8Gzyj73vOvz75Gdp/Jz0F7CcLyqQsfjFriM0GVqfuUI
eKk+s+SBqKEVjCN5PxwosfFBhw/NqLSyD8szgf95Bvw5AT0WZp5etfherbbZkDLvmr0+nOErSjyv
54OJRWuXbq+H6PEL2bMCScV0RlixG9lHZpDNymlmWxBZIwn74JDCxCGKVCiHSntmgVeHk9/iBjy3
eyU71lAzLufS8bQok4bznGfBgIUpjqfRwkq6olJbZxY8z3HLLnTbBNX6CtqA31sZ09eMlxvjn63H
gHFDe3zJX4hqHdnFXxcFnYu+K8oCNME6PiOwXDXhS4wEFv5wbKpuMduSVxVuXD6812BF1ElFg92z
rvbCNcX2Q4lreaR5t0d7oXU906GuNp1KrEhcYmlgAnMisS9jDKjdSbNhMLf3F3a88wNNWm4uCKlN
5jwKWGEBsSmyUu/MXbhkZeItlFzbULNI1n0Z4wb+uf/HHZLTYDUmhXTh2qSowvFviklRtVGAndoz
VZDZQ0SjlfN8acFfPX9fBzhb+CG4PzLLQ4foag41YZTKneh304i+ccLDW1M2lGnzQAv8j+o4pAEo
9lRKdUWnLZG2uhMTOelOtlq0FdwfKXqHSqRiYqr58c7CQhEEySbscMsYnTdV+5RIHfO8QzToZrWE
HYiwM26VGAP4kCXKlnNiliUuK7WAlp158Hct9J5veRNrWn8dF/E+M8ZyIsM98KIrrgJWg1lEey+W
9Cji/YNcPvleBmRpob5YDKTp1Spof9Hn9e9XSVf/5dNyU+0exzstyEqr3FPdhSSjfAdISB9HpK6b
+i6X3ByGYbWCmiYRoEqf5jTFydxNr0ovBODxgAR/6mVyZOFqmJLhGShZYhs9E+ddka8HGGJasnsh
EZixhtlmxea/sgOyUmf+2AU7KE3/GVsnYBakAKaYPh+XqabhqaR+YSkU7W1zCumPd4NFRKMt5NCq
pRBTyXb2IlE86NjLhkN0+bnHhs+sQgk5Uxsg0Z8w2Du3J1T8o7XpYdIINn1xIaGYZYKf1iWkBzdR
ycG+1UJf/qNXfiP5Y14VM4QnGcq0iAP3HiqOpU/GIkrUDfPFC0K046ZcMUqWdsQJIHSrv1O5b1+g
z+biUUbVs2RluXRjQR7sIzrKdsi1XggPGACMkkIoEASp54/SYjW2p5q3vsH394xAjyDuDpDwfqXH
sQ01+Kr7POr9xIqWRNjK+B+r6mNDUa4PUaY0Q4mgPPqNVVEUK6XH1cCjNTcxTTaZfKCB93OJ1Ut4
4CWVbxT309ziR9hYsuBRJiHMVSX/ZO9tpmkmb7lFmlSrTR5BsRWaKt7XDcfh3CiT43bYTUBWV7ES
LHOGfEkJmbo3byK19lhLGi7vRKxPhaS6z/EnhQDJ2itDbTxNfyeIHLAZXzaviQ/uuSSb2gGmMULL
Mdb7B5f37QqaHw/fNwCRM1YoZ0cKIjqjRwLhh6oDJ4fQZUVNAgzeFSnBrTC6wxtLyiprj3IuZi96
xZ19xNtSgNmcQzUcYIBbJ3+1BpSFn4rZmnfTmQORsUUMnBQ412O9eya6rhgHPSIqWwVe5Z/YJkeK
p0Uyo2w9hnkJvxFpFQlzSwaEG2C9SVIcfFISG/qnLPdt8Yhqki6P7hP7xPifX0qE+ydKGWU7a+Ug
mkhZcjWgYfzenP2Qy4jamtLIXYRvVVRrS5GmY9d7cDO2TO+tidS2i7KixeqwcNMsQzQny8+XJ5JT
dqlJd5glRk1vyKJSXZp7qAI28M0OLk3XRgiJQKUBUZfYEGhAohia0YDRmOqzcWaSrrofIif/hv1z
uilYKQ9h+uIH2fxsSyzadlU8K6mvU7sERe9Ed5/6YMmVR3uHy28R/N5jLKyUc38Etb8+i/WWDyHX
+Nh6g8FIqz731ZX0u+IhgGD0A5Iz4aY7yyexzamxzMW/RNVBieorFSrBi2YgZ41Vt9behSYRn3au
o2THO+ZSwTtUMRfUrmT+zgVN1hZcVT+QPy+S/6b+95k0fdp8US2yrT/ePIt+qPTByR7FTwKjNVIA
Pi0ftPa62jGoKaU46HIjbOjwYUg4/7oyUUiinTS1GjapLbOvxJk4FdMA0tBv1zDUMJxXqXbkvbSC
pvf36uE0WY133ZOluSyw99rUayibEDhz7vgClOHHfU/zPu2s2XbqbGxinwx9EilBZS4rnySrrG15
yU7lkvS0yktn2r8qcNU5H4wAN8UqP5DERvvNex2gYnPFQqmIyzfa5MBiEQQbYuX3l70qjnE9gC7F
qAhqMfqREJ2rVOFF08UjAeHZHv42r2njt3dSNhH3fjXyBK1inv/ngjOVVwwqdD2Cf1LP5avurDy3
bGwmEDKcOcA/Cav7SDma1kjdeg2fUkVJMcTMpx5yQ57xN7M7i+DX89HeksUhkUwzmxWclo7AC0ya
O0KV0ECuEkFvWiDUx4JiGPXVGyOv0QbjQfSO4C1GpvCcx1NRSLQE9iglQcOxjgloBp+wh3sNH3Jl
WP2zn2F57Yx8V53RjvpDc5XdytgsJoED1R3NIDjb4KUw/clpsDHjg1q1awth60SKFyRzGqKUcaKh
tVTRzT1n8yjzGjQUEGHuQtYO7NaLlrus0tADyhD4A6Ii5v8rVDUpy7d1A60b6qqRWhyydXsg15ok
VN2FEW9l7bvxEmMqbFpQpkn/NgrRcdC0qCgaFCwLhgK10W7dOP0M/XD52njiYhcnLBnzYkgKasID
0PR2SXLfaq8UOCTUoyA8RGIRh8x3peJKjuc3P36lJSfqTGFa31KrOxilka/E+0G8gGll1qnK1yUO
iWo128JxdfZYQu6QzIsI7AEtfS8DUre6AYLAyWue2RCb6lmLeA2J1zmWnmkfA/0Qh7o5PfplU7W4
7TAccKS7xyt4R5C+6QF85GrlYWqb0N1aYktgPqxodwgGIIw+qAZVLSDdX/AkZmWCA5qJFvjW1tnN
QYjT4C2h9Tk7/ph8JTPhMo2CDmydn7tSC3U5SkoJQHauGC7O0ebe1QWn0XK6xyOf+gty9C4tyHA0
mq0snvYGXhwPTy3UOhT4OZ7IfaV6hIHI6kdc4DdfCsnExaRXtI2G5/woyfqlGc2/BedsYMjim/Wb
5dqn5bQj2NRGaKUN2wZ3hpmMeVMCq2z8HrOxzPcoD5h+6GTapXZsBvWNiTQUexwgO9lpnNprJjf5
5aFZQwvsBAC0l3OJzzGA6Kmn4PGj9CS6ScmBVRaEKJW2B4URLYcOwOG4cvGynfbnCwpAWN/xEXAS
8vfRqIXIh27BIkTc9LJ73nk1ZSeh9JilaTOEUpbIjWapt8XsawrREhQoz+Ef6CHdOZGMp/ehfuwc
m4zUMSS8PiFrUH27R+nO1wWCYQNDU6wa698Ap601VNtOcIc33OC+70+NQ7MEqCEZeSzvqYMYHP7j
u9XyocpM3ZVw/N16XM6FvmmnhSyeR/a2EGzmutJWiWRG5DKamgdFd5HSnZZVWfLee4i1nD/njQWN
UkVR1kHM1pIRfilKpFAO/2xUlsu/zUccfPSrPguwE9CD2M7BjC0F7aASOvUkEJtAPVTrakpOxISx
HDB+ddZGGYSOqiaZoQjt6fHMeFovNtA3UQgGeA2ndpPN1N9HmOQXEgsWjTTYvjbkhqhqHi+7YvXj
dKz/udOoEIh1ItSLkKkprLhm1N//hDW6/EgPO9Xl2XDW8En80zLcVT7V/xiFlHXEa0hBt8Np1Z3L
vAB+iiqYSXfn2d6CLMTl+NepVXLwJY7YrqZXHOpN3xD38l7AZqqNe20x8nICR9OvGcVd+Sqy1y/Y
7QjsoU4nxe3CrhKdhxpxp8r0HoM8Xgddy+tgdeqT1uLNP6RZsNP9CRNTSVj2m86RmIoQVfTmyzKl
u3MdcRJ0zaHGwbUg1nDJqOcojSg2gHuJ+oJHqLQdCM7vRwpZDHmCKHSGLLYsqP3ReqRrwyCB1KVc
c2iCv50C6kfY2XxmizWN++KIjjp2hu17DhE3CsMzCY+5fTDpLdWsyPOJiROpUxtFxlnIq9kKbU6P
GO2HoyWRYyoy4AXnx2qH6lr9HDC5CP3IrLAPUGQBvhCAUJNSmHhDZW5qX28tjH9qOJDABtiJa556
gRfjO4gA2ejLRkJP5nFw5HNyTO6kYtsTzWG7qsvgcTVT9yDzsiulzt9bIQRn1UAWYFLI3xfbg4lI
xFVPJi+2yRaHVnaya0mhb9Mw8brLO9hDHBNbTpUDaLGRjiWeFL6NMfohNFPdeswZgRD8CLEUwJJJ
nUjcZFg9l4WwcLlLtHd4CVagP9xXFJHFQZWosQ18PvHnpJ72yHtOwV0W70DWRIykHwhIA38iPHFr
OcVrHwXe412yWXLzxD457mq979oOwqVvYQfEK5sEET0mESETbU4QFycgJJVHwl2UuGyS/P5nDz9o
dZvoFDBH8BDjaAQSVUVIOoc7DsKE2bqxu1orRKEdkwnSFR2zB0rXwOZumt4cXaReJZKieyMp0Im2
grdQFeQvENPV/Lelrihu1IcOGCmWzdfaFuTHQfq2WTt7FPgQuIi8zEIfSYEO6FjeUSNj/QMbgF4R
w0XClzoCCG3n0FcCAWgTHs4gvE4IDFeNix0zl0xW8J5V8PrwZjIp+NGFvYAwep2bGIxiziIXBQ+6
hRmDkSQcA6YHFOUYuJ7gXg2WbJo0dVnHFc2kSPV1j6PuA1J5chqWUDT0kCyBPCEaJ8YBmQ0TGm/u
AvQgCbNz4dZtDz9fZJ30CnjHs9vDBKE6oZcSTFxgi56ccuGrk6w6e9llZ/ypEGS9bZH0plZ+xM9j
IHEOh7pLdNMkDdTxj3xaaroC5q50fN8PrJZnWUwwWNSMgoo1hL7P1muGJ9dXUpCa46UA85YGMryK
BreccyVB75BrFiQkuYySrKUWEcaMOycCN6VX2jTBzdujMYDScTSrgXnFlyVqAllNBRatnLHudR7Z
jAlwAFX4xAKgmRwRsPSI0ayYtmN1JkvNPma5FNtSV/U7dor3Zp/UFWqI8ewguzW5weoVN3OYvq8x
1cyH2PqhKKJtiMqykWtR7sRAGmOTkmL9l6fEOQuvO6qVZqXhxokEeVRr3evcokfuMfVisq0OAk6G
soDFHwotJfoHR1bdSpfmXCfOfchwRgrGrfLtAkmOwCZEdCCLAKCBLyev54AYZdGxSYhxhSUzuEaj
xlWR4V90z381zJeUpGxCIvY0OLpAqoBcbwmwx2SdQopvkuEkuEB9GVVKzP9VMNBhEuHtN62qZl1H
yukDYTLzd8p5z0DxIg4g3S6BP+8lt1AyTGLmXuA5X1Yz3BFW8AdSBrv2VoMqkOIt//oJ6jMGSuAX
7DLSy2s8QtfVzrOWtX8hMyB2zf5bcsXqwS81amNSSwxOnKHC4gKeJu29WTHKo0FjBL/gP6ISykLk
HyvhPMYvvXuakz1dk+k8YizXr3O17y8/9BJMDIvBaNtKdBuhlVKVMKlfyHvtqdb7+EvonsqFpAN2
BmsMZ/dPdImokNxvta+dnaY3LcTSaaHsUHZPSmxgCvoLubKRNxhbEy+mjaGOP5jBxcnKv8hbf3g8
JFGYGm+duel2NLxYnBQXYFiBvBAJ/HAvjbB0OL2NRl2Itgq6ZXqdN4SFPRQQm1jH0ddmcUcA9iyi
jYBAY2heZAnHANJ6qBhSgBRk9DZ4pwkm90gD19sllw5vMakjhPL+bjnQGOijL3wXNjh8rWEj4n+A
BWwvNQeLuFKyuiTlBLGVYuhGZ62JREHRQu4ZYprA0V3LWNAeqJyIZCSx5FJETGyh6bv5/9ZWRxDE
L7CKkfZRaF8STT0uqSELsy3RvucUo0/5DJeuVhvjDt+eFmEjJPEWrRf2Lryew6SClMA6SjrmVqvu
4k5fIXbbnW6AVLAWjk66dTMUSHfnbpaG1jugrAIi9pLeoaAlZI0xTt+5oTq1wogKuKwJtAaq7Uvq
lh1sxJz2gAvArAuWwAay6L8qnspSgITX28ChAkGssqkKQHM5Pz9aurwkmh8tnYeodXFDCSRqp8ne
sRD1gxaCibwWOX3Vl2J4Np6Wfdh07KxLqZgxPW9/l5h5KOlwCf/Zd6HWE68m0Lh/r3p6ofxdXTI1
c5gLkACVdryLZC3zyTqbTl8OkP0/fQcZfeMjdWINekT54bThgAw4IZh7ec8nXh5cl9L8/83I4FL6
KL0wl2VdDjI3y/AxflvIRpuobEfsaZzWJDISSSKapNi3/muVeI+QmX330r1e33B6VPHynA6/T+lm
/PCF/bjpHYJghP3YI5BcGFF5yArgUzp/Uf80GMqOMZDoZhVDOA21xPLBTxyN+CBCBSlca0AZiZnx
JzzQN0da5aNMfl3f8cBgv0pmg6lXA6BlyvmuDZ/pwlQH9/fHtTMZKmwjpon1o5VZ/i6u77GtMIa+
8Om1uUV/cFVxI81dFZub/9itQLv8sHnLOQk7/4OOaugKPrqnhDJFZErvvE+tNeVpOoWM9cN9EugQ
hK2hJgojb0Y4Lq8atoq1XPT/ovzlwLIrp/fOvdkxoCXXh6GtMIYpK0eX48vYC6ArauM/bg5fFS4V
KJ30N9Kpm6gmvKPEtfHIwpTtV1nwnLDCb5e81TKP/b0Ol36M96xe5azpsAyb6hPKHfP68SkUrmAi
tFC+A159lgfqH4/ONYswwlfNFWygyqQul+tbwDbUunY76wDHs+TqdjvIrcsiBJPxjfswZPk3XFU2
84n9GquvT6cfMI85b6xdQKXF2fFFsbOl3misFJvBWTSp4d9IJ85qzsa64VVGPQ34IASuk9CwTw7m
LepVq0KcxH94IiZIHbO5dLpBVu7hu2mSP/RLwQWWRTvC8cFdH/qxZhs+oU2qF9dVSvUrKvANFcrX
wCSP6kYDFHFx8uehznPnKmqTQNxjtuEVpwzdXXT0jG7pbl7jjvL0PnI+Z3Hiujuv0ZfsEY0LR1g0
XylkE797JQGP/5Za6fWMrYZOb9TguYY2KwMCH3IvA3MqqJwOOOsr37VRSMNVfwRz5xdDCLtpaskZ
/DCRG8q7Hx0tyQBTZ6mJe4DjJht+A2KZxZTln9baICJeF5OWXvpa8V09htOOKRVfvOPlkprS00BX
4k0fvcgi1TMaYZtdJodPHjMasXrquiZoSNsCAmz3NkAPWzOqhYGKCCkc7TIeMDgH8ZoWdz/paBj4
ktpPtmU85Rt1UFFw61JmjWSj0let+lr24O6jmzKwiQOGoaS16eBrltEjvz8dh1gWNUKRyqwj4PUg
UYgvY2L94Fyg07VrkL3q4qISdHtIEP0Ug0nQU8aQ8O6RwgzSEfn+q0As+TtIWZRjXjBVt3agfyZH
BCa0nVC8Rbmurz1BDkCD6dCYudHsiijSw1K8cAwokI3+r2yXZ2fFW7UtLd45cEUDLPFpvV9su3hx
DD9Gi+RF/Ny7GNPv6r/MdU1J0BPNNv6aT8sHqpWF48b0uKgOG4P7YunF1BmMCUs1QtxCOguUSC69
DlifB84YOw7gd7VF85wWKYIDxmDSVMpZj2VWeaLehEuN8nsOOxKTyzWpuOU7lLYtBWnb9pbN/5Gg
DfVvQ4cF6F771t+qQifzP1KtjXw4PCOYo73rT/Lnto1K6wVVtKcJAcDa+WLrbgfjyf2uL+mczLej
OaxRIxYx3e2JlGki+1mOnSm054lXlLEASScZE/4vwrkDWQgy9yMus2QD6+54XNROy/UlaSp46a+z
vZmkSI90LKhf0gAsoa+Yay0/BITcjerplii5yY+WvBY6fLUbrxfkAIZPHlcELfgEYczdjM8Rn85D
6YIIkTt6WC86Met8hYbeqNEG/dl2UxMkUof/5mWdRF8VlyV3nFU0OnvIB/1wNx9OsddqR6pzxwiV
LA4QZO+5x5cJ8LgalgOQLmV6sXYtTUeTuTVeUsLmjZ07EkadL4aw8EPFti8daGD7iMEULnZhMluo
d137DDvO0B+V7/HDqa3bYvu2RAu+eqRWi4146nCgreuKEOM7xZL3s7x+OM+y6WM/lfbPz2Ec27NI
nj+g12fygtmbiANylHMkWqU/F7CWmp7mZ0rS/Au99qx7cl17hcQchkAEQlSotI1BIssN7sxkDgdy
RCNolAnLIYB+nZeKKCTe9k4aBTDuyGmwqPSbAWzDFyEpOrvZTulhEEqJSjlZ4miohKq1S6v2iTAs
RND75QDS/sFoEjcRXZaZXq67GR1sX/4GAc0zyBlE0F6ABSj3e0OwwtUdB0yW3dJdxq5jb2L6DEHi
C78j8RKevWYkieZDgqmXVcC2hOp9/HYGso3/NgHo15jZkM8AsozzSwbUTtGL+84i8wWR0a8k1xGN
0SJC6vFLwvbq7F7K2c1QHN3CbtZ85lFSvLzFg6nfpUHeneomf1rNr2GEu4jQbQxtMdhvpKs9T8Bt
dYFutdN1T7IG2qoxbqrYQvW7ljriSRz0eaI0hN6i+jmWFKUnR5LkLyIHW8zydFEISGaEKJnE03gl
6cuuwn1XvL4aJJ9LOYXf2k/MOMvpRauY7tzD1Ngg3eU2Tbx1EBMlG0yFlonyK6YpN5bhfqU21N2E
HfSpS0r59pTBwDzlRxNAvfxg2C0ZudsRJE83Q1LIVI9hqAk7nUSmrg0OrKMgXe3cCGGHkTc9SJT/
yWkesN0b38qbVmu5CmHsKLP2MjREY5I9Oyx2fZlHaK9NqoLYigGSQcnWkISf/rx1jszO4UMFQbeh
q9uU3BxgjYFeQLLRcYM5PsmJWsOJdN5OJVMNbzUHDky+eupT9IJLmO73+Eycv1FD7dQbDw3gjY1J
jm9NZHKBqQkYFBti3PU3CkxrZ0Amvy1QijWQCrSmaEaI45apPZLXJh0L/ll2aq6xiKGDGChzynIi
vh+CZ1YDrL/HFKxHhWeMjGJobTaSlFeRIinvaJ/VWCx0j3id1TuAQWIUQIOkUZK0wd1igkMal8Zl
Ej0CndATlWcT4TfeNZaBGXk2kChsd397ifDYx59p4/jjU9u/6TdVuCYRp2c0LvIHn0SxlF84kcif
rqCCgd+jtl6uaIQj2zWaWkWiYxXkNRGe5NavZzaiGBsfEWBmcop6D7TplGzSOiXReOISKqk5Qvb4
wvGH05DbtLZ7bhKYSYpYN0gX5nUeIazpde54VqPy/+8Pl7VO1+GxVw6kRglEE+/vp2a+qP6CXp25
Cci5h76QfwAq0f8nNQbGefbImMHTxAV9ILDXWo4sDIJbwuRwSTL2nR14gc93bDk6Bq4jlRwCgwXo
RE1lMmbULw2knaL2kkQuI1+x67ra6oApZbSxCMd9TFYHsiJVuh3U1Sy7Z/0S8rTPQAeqMlUEpdN/
8l66I7ouBG2kw0IUnoSko/VwJtzoQSINl2tiDfPXxE24MjeD6+xcoQubQ9iKEmJGlGK/Mjh4Dc7k
Sr7MeHpp6qJensEJo/SH1qsQct0kkUAyN0XplLvj+PVDM3fBRnkNRsnBezs3u9+eZ50Kmrt0QwpV
VsHZA56Mwgj35Val3QeegW/VyzvX67miR0ac9s4fJ1m5YzqI1AMloK5ulVGLQ/qYXASVDC7XvPgA
c2YjZe8KHjCFvsqazdVBdKqpGTAcEVpWObgkryrm+hd4gyrwr70Uf/oM4y8762WZFp7UBWW1o9Yx
KBTRMZ5TjpSbAmkU8DRXMzQ3mVrroMvGfLr/lNBc2EbxnH+pxyA9Olj3fLbEUt0ro04KotGJKSYs
+qeUVVPNVezu6Oy57qFHbXjm6atud5vF9x/0/TRZT6bJRVxDtKYfdYiKUrcnaZj4lEnux911JGUI
j4fSsjZFVruP23sUwy/IAQwWYlgM3ywdvDKT/ALSO2tbevkzhuj8q4s1aueBILt6cq/gp+0KAFHE
95Rg1BuE7cMOVUnYgdIFPvAzhgRXkc9d0ZsvjMOWcswyMeK8IGk1HhsOhb98v3CsqOHsbNHjxZx2
G3UGYP48Oq5rnaWJb/453mgqPcGHlDTEXVNsax7I7EX66PYDNxNObsOw4tkxK3Ae9tug56LYJDhK
56unxYLbhm+NGVlvc57PqD9qiidQrJz31E5GwBwhcrSh5nUtEQGHpQoFWgaxzXFxnL6G66tMhFqW
H25vjhfBTbS/yADpiTDiaQCDhdNYummb3jR0LzG21ef277W5Q9O7ORC9zg4XcsQwxmKIGbZUyDNG
FEqhIZ+PnKkVgo1dKFJD9aZkM//GqQ3HG9odPsvqKOa+V5x7EtwaTxrZF+L4r65NXdGMER5jeexW
D+6X/XyzUAbrCX8VBKDvXYQffMXL3CxgpahCIVRXf5fVJDuTh29GX45C8xV/Dtwyuh9J4wRar35a
vvqKkO0+ht8zbWdZNpaa0wflfNYJGNApjiviC+v40lowRAF0G/mC8S/JFsORwrfVYSt5zZl7hQyH
efbyZLKvOxwN4/G4pvXkUxb7QHfinbNYBpddJcVAtEeGP16LCewNXqizRZMJ09xVwH6N8LovssvN
/Vxmye+IyavDAYE4qPBLul6BE0kKmptzkOYP3KPy17u4/jp201E8FUOsi8nc1gMCJoBquZLbgFEh
i07KSXa5cXbIKi9rEH8BylK8Iv3aD4DqGUcGHuGMGlogV9gyrgSTMFTEBA17cfCdJ0hkxj/+5wqo
bEbdX2viN9aZoGmfxa/TofiTFzw7aSmzUiZAqzhmUJZxfH/ZbfXJEngEvOUIY0/VfYyZ6eP1JEps
S0y6YOBkiNPcXKsrTjhMH9RCPF1I8KfP85OPtAnSHKsrhbwNCdxoCcHuZdTwDi5Wj07ie4CVyZ+y
biOrYys4KK9LhF4dBOgv6rK7h6WwpxXrKIboh1avCoTMT1brnL1eQSMo0b3+1ZIh78tW9U9Utxhd
S5hTPHw3fAgGlQ/7pCfzKDGKhLtIdS/AQmc6vu7dD993DZUwypb+gfcPUwWSq5/gbxgRbjWS46Xf
X9GqBeqAFGqJYgwGnpKeaYy7Ggayyyp1Sl8gm8AlO8XmJvSNvkAu8J2giTc82kRLiXT8bwxLo0NQ
DsycTLo7mvB8tZDVeLzi95CcNDSSS9gdnVefDGeLka3bvTo+kSkL/vbBHUrrNv+HPXll38+jTrVP
Uv2Cm0OV0n+9ncErRCWz5K5QrR15tvAPdCCPT/CSv2PpZVDrHRoZRF4tjEcp3ixUHLy07KfztlQV
53sb+c96pnGMhG3BVovIlqa3dsZTKhDkiRnZpR2YOATlRqiDO6f3m4Ff7AZws3v1pbvMNgC2GnNg
8AYR6M4gHeFI1qFZfdRnpb8SCqGVoAh9rm34J4//ItY8JokUhMtY29xOkT9iVuaMgYHCAWPSAuWd
ffxH3eqJXnV5B8rxdGpKbgRi/RDch6Zu7OeGKk53L/bgDZIqxSTLfkZmwOFGvZDUbjxgkElqT5+Y
jmNFpIACnuJ43GeBIbMRMTcvc3n2SwO16O/Cbh4trJRNZkAlPfk9o1rhPLTdKUtqVn7TyLsvXvgZ
SAdEDztimF1MlZRW2gbjANZhVG74BUyRgAiv3PA6P8rUIMYMLnKc1XOrBchNsIPLsLsei+AgQ+P6
+F46/zHvNxuB7T6mWASeYsgSRBpfQCvY/7ue5maB9nzVj1ZsD9L0nKuv8dJiVxb2ZTQzKNjJr5lQ
W1B117/MZoJA2tsITUdKaF4MCgVL1PzacVdpCSDkQQ1o0GObxQ6SOg72CO6p+3S/behiJv2K75D0
E/vop3QMeX15Kfil7jZBO9zbWPI1Ww5GplgXmh0E4qCsHIrsivtH/kDGVKZtltZN7uV1aCfRB8Re
CqdJy4PRDRXTmsQxLrOHjxONgG5vYM+h75d/Ut59bYxJi6hn4LGHnttaJ+A38vOGsABIEOSn1b9f
ELXYWx1VC2DUyzed9XiIgkSRicug5gw77GEBuj/1+/OjBCWSYRVIWGxS2w8GrwQFcBJc/deIdUG4
5TLGaGJ5pRA9EtA+0UQaqujUM7I0GK6qbWW1x/HgLb4MOZbWOblYr3qpQNmqIbuabX6uglp5Wc+7
bRYB4who/8bdvqdpxhpyfKCzqhXMW0/G4E6wNqfMWYs/a86mGwJp3itkMuvhwYIfCq+iyZU5Rr7e
e2hzzBMkjJA5PdpPG6w6K+83gXH2DQle1JjtBYBONHq6kLvKrytyjIHySqiw/pHfXqNBS45Tph3K
dmfSmwfIKpEM3az5x/TL8WTW5hAC7eICLInh0F7Q99r0iPBUcfaCfGCQEMvq+7Wyf54gVHxVVd0c
cG6Yjl+bIJGjsjD+3uZX6sHbsjJjYzbzf2iO2GIRu7lWEOIV5a5A/tWWk/ENOmHqBijhkf52/JHz
FVR4VaGhvR2FplW00zmTK4Kk2Y6S14+MmJaNpdzHsYr49M00bY/DdPC9vkHf+JTAc4Cd8PbGuTkn
KE7UPJxP1b0zEBv7/CIQeLv++skopy+5GLNCaCqmEbcNJI48Nnjg415r9ae/doQgA8OzlCaYIqvr
dXqBEVn2pG1PiIikcbIiT1/WsGJOJ7jdXhDUhSBRlKCq5amzwHlnod45z7n0BxWrShfm0eR61cVR
NPPVtgHBz+fjWl8SWXgCZy7yybUG7WDITjAZAI0uXzTGzSHo4UIQhiGTJZSx07p2Lab/uf5rjKim
cpjN/VhJeFbfyMw/qnuoiBJksAWMYxQ/m3HRDphn9H/YWAFI76tjW/wHO2md9/8NZSZBXDK8KcCM
77+/3G7DjBhMR9952mSSU1UlGsYAwVW1Qsu8ZNU+W3QvTI2TfHUDGY8ks577bKMH523T9wA+CuQ9
w2/0AL29Jgr6fjctT3SVqC3ZqTtKNyNeVKoRy+L7ix5b0TW05obCc24JRKfJ4mlGDFLfA9supdo2
jxrEkxjMWGHbtPIDlOmfbHcVCQAkevRvuMSRJ3EoqzwxWpEIr44l5wpfE9l8HmZyMXNE4v7EwryY
w7Bb8iqc6md/7hkuQUSGxKetc0K/skMHJfoiY47/u1wuamvu8P5IJZ4ewHZyocAb+ZXSbMdg22gL
IyCihc5ir0iwefkCLRtdO65MeDwEpjaEsezMrZT/OASw4bBuwQaaXZyNfgiHYYK6pDPSIw9EwjI8
Wyfscoil3YIG5oGh8NdX57CtCEM8kcw0N8sw6NhKq8Rbc4FurCJHi06KYmx5XY0U69mGn4iLuG2Q
86Y4pZNEr7xgb7YggtdE30dyd839xs8czNgS9YIAEYBrUlRJjE2sARgqcDICvwnyK8wfv3KC/q6W
wMKATCA8qBXpD2x1JXITDiYKsRcyGYYKKYkDBCTfQPJWrgEdtd9fXcheDRyEW5ujQU532j3XeyO6
giBo/ZajTp/5mziXBkuW9cgrFrQoGnr6Xb8dd9kbxu17idPIElAcYZKhZ2xhJFq9jbtrG0pCnW7E
HKNHQadHfdgd5U1h84pNmtNYVLWmVQB4KSf+Ecw9jy/LZwFFVhAlqhh/vIdrHZEQ7r8KNjVWU4Gz
FcM7uOKoiITreR66N8c0knPlFmaKt9UMgFanxPGixcKPpQUz5QxnfYeXfD8HeevHCLKH6rpU0zuw
NIXBFx6iolyBGdNScglwEvmSuIfzoNGAt3xzo/5Juv+EPDbv2+sPUSdIULJJX4I1rYEYUIbWXSWM
S4n4tonJx2jIbCZan3OG53LtU+w3lJvyI7seuzLC+KyupwRu5WORa6S9STgzDoEIoqrnrFAPKcKd
eA/f1PyNpZhLtpSk2sKX05kB1jVvtdPGbjU/g49Yd3skgX4GyhPxeRM7X3EoVKn9EK5SvTEIK7M3
eCNwrledMt8M407YRxs5cZFdonhaYm9bgthRKwLgWMtVug3ipID0GHk5c4TmUHpolJuQYnIWziA0
RvV3m3u7qCzVhFwWOZKlYHhAtZ4Vl9YYwvZz31crCEsLywGh0vFyDcboMYoo7kFhwuNoHBAi+Z2U
gDKhiAEQVR/wQVUx0ZDVSOTGi1MgmQ8o2RUEFgLaMz1ATr3DFRGiynK2szL/KSf8v5G3g1/bZ0HO
T/19y+tewI5adhBiowlk2dnc2XoeIMy06Im6izlxveBte1B70F1wZhtkQ2cGy33ICEXicwvL2hKk
BtMJOMURxV25Fpo/FHC3zjf676XXEE1o1bWig0Ry9iIlLZ5XAGcK2xcunNAHNoeYfqE85SC+dJkW
ISehQbPi62XlKNK/Z2wjVZz4hMs/oV0IQ+U+JyfkVgA3fXOYqCPD9d0UgpV8RivhTlRnJfmpBLtG
WAUaaTXD13EGJvkhqIKDuxza1pwmL7qZxqiV7U/8jClXDj93qyhbLdjTh4TZwyh0vxbqUaeIh/Ig
+Ahu+jDVTAG6i4QmEhpt/AClgE2J9uQecRcXX2A5bzL7+Whiqs4Flcc3RHXzF/okKzU5Y8+iDC0e
iW8rgiohqxv4N4PjENGTOmBV+Z3gRsCK/O1YUlI1+APkMmbv3YWWoEBo7lyCZCuNTSrLO2ldbVuj
scfEwer3ANStJnaPmsZBUl4LhQ2/p0Ttjwi8p93jlAelDYLZ6SGH8DWDLDH89abbw2HvFHFNa+LE
jDzcODnDbd2XZf3rJMyxrmYMog+PM9bXXjt8Ah9G+5lcv8Ifs7MEobjwirHW6xvxNdFnBVCPY0bC
PsUhnc2cqETUg3vpKV1fjiTAiQ8iPBBomBvfUPcwG/4a0Eo1J+Lj8ghol8I2QH9bu3ZfqUuQmaOd
eGsoAsT1nbRPWS40iKcdvCfHvshOa5kGoqGxXnEw3s64YepdF6PVlzOzurWZgvBr2VXzwI2dmN0S
N5XlWhNdE2vW8ZiyZiP9VXrQMzE8Z2GUimvKabIe8ywGIKuM+a7y6mCZaHEq/CqPBHgsjNhEO/7L
/nnWE7+DOW+FPf0or4s2B4TFxLIpI6OuMfb8tIiG+7nO7zmNMfCelegc+jHiTqf3gP6CrE4ddXU0
hrwWehA+e8SJGpVAK3WjuzZyVdVqW+pQSfeJUg9I5vaGPo/BRYxIKt+Ki4pcqUUp6HCF2K5rpuGe
2O6jzG8u6JBmFkAOVOV2ZiKSyD+EKZQzdRC3tDzD2ueQ5rdAo7aXW//MBn0TZ+uPLsZu8UWhN/C/
ppUEtqv+quQwbRayuYW3+3nq5r0+Iun5D9/BuSLXVENOXXtm4GO/FwGk5UiwOCQtz6eG3pgcU30v
H+PmsZnWlUCDG662QqeHUAAnmRoD1xXHFTvRjFPtQXlzI627151z2eAhUhqmJb8Ad+ztExU3FsWr
nhCp1sraK3y7+R0QMuhdDz25joGAMDNHYWukjOPVBH0Pan53gWoCkAyM8QhQnl0s4YKUMiK3rCj8
chSL7epMEHz4coQDQzVtvIUsZQEV7SfPrGsMEeZcHHU1JKbdithc66sLfshn3W3lYqDaLFni3w9D
4e4Ozc64/bkyeaM8qTc53/oTYhILqMqsyA7p2L/augwDQfzQDflnaODaMum3w8Wi1888MWwPjkSN
2jOKEUJTr87aPBjjCDsLi8i8DIA9OfVpSq++kmUVxWoPbnW0MtU1UpEMBHLzUnZ8ZK/1VasQ4p4P
H4tqM85IypDWOEaNWaB6o6rSbpGnxguYDnSg3aDyT1vMncqDhvg2tS33ac36R55q6YR7GcDKZzKx
aPp7xA0xGUfEvfeXrP/XPkNRcurxJb+9d1tOlf4/4suJ4PIM+9wtHdYOQdBg5Pg/MdMNUMUeftdi
AhAtsp568yvJDVe7/n4gOL2Gxsuf2WmBnljyQ1fe0fuYgnYRzCk7MJGetPYHYNhG7xnyEa2+LoX6
ttMFXPYOAvp29JHvwW7zVEid+It4e28k2AoNKhZF3R2LL3ya+D3MunNQk/QwkCl27XfkL8xXR1qc
/eLospSnH4E5r1ZrvWQ9ZkVjhpaXDDdnDj4JvJVWGiYIPBzF3inZt+xw1bui0F8zoTcDqacWehSg
VIfYPp/nO3n2hbm2lpUJHFJOY+Mxc7mmdBjHDVl5xUs/xhdW7qddO0gTk8AgLh70PLPagH0Ztrp/
NJ6ADvr9iBBrCKiVRBxOJcn26qaR61QKKcScDByQPaRBkhitBNrfSE6SeH8qoihzXo4FkbOzXkXa
O7co2KkgKDIBWXJOo+zIMKQ+XF5U69dkpBKG+SnvDc5NbQXydIlDEDhFpyIYxD8ESoYc6YigI8Ng
KEIczWBKizdoa+0Gf5ytYtt8wx2uGR6oPdmPl+C/68alXq4ccoQhhpsbgSiEF/ALr8hnUJyhwN5/
M2vyU0Ut0/Ss6BiF+/MXSxjwKVwJVJ0OpinudqtF1Abu2Rl4qoNGLC/RJ13rHzE3QghNiyiSnjNs
wWtF6S9Pw/p94LoK0vOG4Xz5AD4bnIz3fBYMhLji3Ky9z/Liu4OWA0ODIG1wt+mnfl4/q/8kQvJP
aoEjD/DsWUDGaCPSTLC+WDfzp5C1DuNOnyPpvy53iE0YujRPl7fqynh2ReCHqmozJxNvecBkVUZ8
5jKgfp3YwR/ACf8FIE04laqmHEYvegi1KYp0wMeEpoixoLPj/g0yBaNNUsY9wbAe+89qmsn5kI45
NnQ2t5ToLAHFwYr/CY8Y56B/NtKYNT5mTYIqW8hLaGIAn0f+ozAHhXJipsqh1SnXAwnb/YX43LqA
q3LsQGvrGoWeCHplMRwZkX2IVQbrxMEIFKNyAr2c5oA3Zal+0EuDsw2ofD/LyQs2sRi+FAzj1L5V
tli4oanuwyc1mSf4AqGKSgpsc9LLVmxcF4evyhyWNM/USBgAOHbBy4N/vWfjNj+2JGLax6fzaQhk
SJeWRluq49VcJBLrlKgvoHY67JVXzYylg7mA7aesU7Ae5y/yI8Dpq0qbYBDdzSkN+Lq1OQFvAtr9
cBMy93+pDyQ+mHPGeba4yaRlONodG6RYeTXfBFJVUjusAXAFNcvSyv/3UGAXygiumHH8yVMs0+0M
3SAbW4eFx7Xj/Y38hjZpESRRGkopYAtwKutLzGGApzMhAwnCDkrQ1BZxbIYEpU2TSiKD6Zl8rPRg
BWAc/CStibKKqYZ6ywamwvb+oZSaBWC3OdTYTj6xDbbwgGYFrDmOQTcBWK187r1vN+YJMVsLGJSP
UPz6XuBHqWQzvxXMoalFenud2uUNJtwiUFsAMm96olSvpM23kL/Va0VETnG9RO+dxPRwxyAwbgI6
GDmEOeTyxt3HdW/lnPJlh87rW1qbJMqSOALMjir8mTwcSmCIZr3yqXT+Mwbtm1UsuIKPiWEa67jP
mAfrm9k04SOQiw9Z/infwh/hcF0YKrj1OGu9Kp+C8MvdLstKdGSQhZHqquHCXQH1TBpd3eMaEzB9
sE46VxmBYtvmGqxu6A5AhwvnHxBmetXxKCOUZahcUiltAI7NnTVVh0/29/YmGT5mKT12FdgX1u5o
mhV3VGJAn3n94vulbvGWMAhw7hpWuMkQ3I4X2vzzWuZeqPycGfXGBhBlEjiL1kiHewNalmTISTlK
yqf8tKzhkFWVX6LMmbO4wmDKuRCNcfiYclb/i/cACvoJQ1JcImtaGglrMoLi1H/5bp1emrfxYHSb
Dli7JNTBj89ZQ6WUt4qCNMGczkLGz0Oi4PeBVr0FLxb7Zns/FtdUPB3xC0D8kaoDOGvnXz16aUGE
XEzj2bc82F7zo5jMIwtzZ2oAJGgzind9A7o9apJ/GkfuBVUMBVKEvY7CS53vDN9V2ucKlwFvPAQV
FOkKuWjaXlT3/czjSHauSJ5n1kxmQZAJhwvXmUBnAS79ptOes3f/bwPrBk0UHr5zTLXgbh9PmVX1
qKjLZXqUGuDvtPmKwoKD7fOveaVQdZmWR3KICt0TWGa41wdiLKy3tng6HtTqhevuPLujBgCUgb1n
cda3bCVVxw/X1aJHvUk1UCCpTQ+UsYafBfS5gui5trRFwq2nVHZe9e7HVwxOZMFI4TyaDkwD4PE1
bng9DPTk9iCZ1HOsqi1C3iZ/S/G+VcFGMglUy+/vBuW1ip+/KR/G0aMafnsFi0a2eKxFFIepTTeK
7GRPmZfi8ycEEA3JCrfm58mSKZo899x9QCoyiwiS6wmHwwmeFPCQlyyY6LE88BxcD3WDcHHDasCm
GsqNr5szsbAMr4L8nr2wvxVLN03NrYrXA7mGbTRez3NdVYeV2KWLTPHQMhXonVV0TJvebZSLtsa4
5qiJa8ip94WguXFniC8uEPOERLmBVXJP3EhEoRTrwGcvTFYPnvMRM2qyAOYe17P5fBAGEueNwiGL
xZTH3PapqaObl5HcmEqoCgI+ZrFgBRp8tCz30NeUQ5ndeV3Zgi3XQMmZ8pSSTSmhbPdFffeZohgE
TLDRHk9cfZUKPt2+Pnhv7LsMZ4iGZ0CneruZ6zajxLHMKylVwG1ZcngU6G/yUfqaka87t+n4SCas
qXw9erkPnQlSUcLdwZ2EiBHnpL5OHsBdboz+4rQhpHuqPef8aXSNFAcnZvY7p60sTdO7k5NVnxMS
WxwoTddw5vp2jR/bpSqLfHSts66UnwYNi1nGBu4wak9/gYAZJbA2wlszLV3ePuFwXno1RK6+F3bC
3XUNN368Bm4ikBZe3MfTlQ+fc0/ZdL/Wt3HykQ/hQ5HQBFfkAFFM6FsG/ASoe7REN48VnbeR43XH
wW/nYbFg9RbanlJsGrDinR3pBd13oZJXwCtrab2BVAzCIfd7gfRtHaH03RaL4ITsTLR9Rzde1yUc
DpFQBygPTDpae6COzJnj0PvH2xxlyJqpGKh5EbshnK89PF+RTmmuYP05pGWfYTbPTGN2O8LDcJOY
u0hiuN+SBqVZ2fgUKGNEPYSf5RMO6soUCmasV5rDcgg7+4A8np+/z+dKbrTsl45gCYMhpSxy+lOn
cFvrgDYZ1UOFeXKsd9QCCtMFUXOjyaPe2dY1iaSDCp4aQNdYOmMCvZhYujm3XAOiFl5JB1Klil+X
Xuf5WjHmIVAB3FLfwHaWEQjPqH4qEwHOQYMVLc+o62o9J45xmXCkyxMVFupUsvNMt5snot3+Soks
l4G0mXXema8Q6Nks9CiwVoN0lZMTVJa7KnvG1VmR8ivkX7gjQa4zpLpH7shghMVRYTve7tNI9ED8
882QQUt8mki9+uvkDq6VXzr0wpTHj0EigIszWoLJQTCBSDvOyiZF418g5+t6ay2oCfZZq7RrsRlv
44Pmrz52VkvwE/dLetqRFvEGRFQbWHc/uMj14K9UMmSAA76WwmiGeWp2V9nmNo2JHl33zwIZhEzr
9SjZO5FPYJhpN4GKG2eZoPQn3y7ye1kcSYbhxglzjYz9qpzfqH0r1b6ohFH0Ng0GdF+Ch0+sR9mG
rzWZnC/n9+7rbAxHWT5gjTsilhGPqGPOyNuGD/XvlB7UVm/QRFvour/LThcQSJKqC/ItFAnw4wde
iTs5Hx49/nN2mayTD0ObAGaooLYq6Vq58IsvfwgZTxtAQb3r9acOxDuJtCJ+8XEfg3CmjziOabDU
gy00PrDSqa/7Bj+eDnb2sSy6IgOLbO7HUDx0k6DnfJncL2wPe8INXjGtwvc538SXfiJmIOGTO+wS
fiqhuAE3rYNdeQXbsrLeYKeaJMpt2ZZKi16hFvmu/Bv6FDWD4H/nHDBS7KcHoH+ivMdZYlOVBVNK
Yw9j1ZAT9J1eomsyw9aO/3Mgr9m1vvGX/9I7g5gz0rq+2/8WAU95c1CXADxLNT9mElJtXGB4OR87
muWBZf+73yR5L1W+hpFs966GxCHKnYTBmfgXZUmbkWcJJbEQuQ0RBtuXOYMQ1jQV98OuUeOleZ6v
rgP62i3xn4UieiW+wds6uNBTN2rwPAkAmgJouSNZAyM194se5O6BwGpT7xNAXMXYg5dysWSOuJNn
Lu/+rvcrlW7HaChxkRJZN9mefvd9fbEi2vLCv4r2horboWvnGk9YJyyghQpp16j88Bm1mMbsc/tt
ZSltHXBGsrBRJsA8EEZEUs9UpeFOt/9j0zEiqdkqJVhz/pUGjdFLk0ARWFBK7lNpZRAL59VducNk
TFJO3CPSsRMa5cDHPZcBq6CriaMmAtIXLdAyWfzIO8m6UDnjN0MMObuSQWIzITYWum20p9ykVrDE
xA99UbO9TqHSTYtKiKe6RRndv6/6Xk0Y9quWhORKvv3hhHIYH6H4xmDKVwKjiTr31bA2HSuKWpb/
opJsfD4rsyJY2Bd4I6ui9IVYJPDsBKftqlnJdbZ7WzW63l6CwfO70fYjoN7ShaZTZjbGivOu78NZ
VXIdqmF85mjbo6np59EcOr6ez1f+26NCVn4Ov35vTvuXqKDAiS7+rOxPTcA4Fj0n6afpBeTNqZm5
sDfmds7Ikj+9KCcJqzPzWZyfkvzDjTHNT0NlaQ0JToSHUb3UHN07pN7bgvCy2f/baF4gwH0w8yir
ArT1NL5sjEDyFmPVyurmPpTdy2ZnXLfotYNBWoa/7YbIMOB4CA+q78n+Y9puwovOLGCVV8FZROkn
dreFpjmFNPPosS/AZXoB1x+fGXJLwRs5vtu/MS9/sl6aKb1AyzCrY/6fYr9Fug+II1MU+w1s2qCe
T8A2PyDanoMTmnZZqtwwsWuUQBWBbaHWAJpVqBexcdvId/Kfr/SRL+tTTEBZQGmqS81dSix3Y5rG
zfOLS3EE/ivxEL+RWZcuJTa3vCQQvxSKo+5AvLTliNKobRmjKX4A4hgvoNWEhNjPGbMj3zmdhS1Z
qGvk4EBb7Fvl4mINZqGG6FOkLK4Zyf9JPRY9gGzLAiGYlCCsAOWS4dSMIQ6gTNsuMK1dQpAMLRzT
uGtTwRmVXx2dylS92iWxvbKbS3/BZV/cP+JyF/If3Zi7OnZ1oWmhHOIm00yisrdLA6q7lALa6fO1
DabVlbduh7kryccDBq6WeU+mQFcRtzm8KCQjZZ3ErhlPEZoF4KhWfKfS6zseJW9zUa2k8yqzJ+EF
HvNSjLw6JFBvkkuT4utk1ZAi37k2VGSomjfWbpTeopRNbGLjFc9nuKwNWuf72jfLX1um3TnUTDPw
0aNULiFTRO5YJ08VAWjzHmFgcPytWg0pyLrgtT/9LuVvbrQ0Q08wztEsTDwIURkq6iTMdONaL3p/
PuWZyne834hVVaXE6bOfYIaX4uqbihzYG3t1EY5bgCiH9T3ck304jVOst9t09A3A/YoHKdUtWkJk
ulFM/X+SqVEOMW1UWUDKePkUjh+X0fS58zE6fipKyjq+PKRGHPkYSDqQD/V+Yum3rUOrytQMkEv8
GwrrtXOkmibcjOb5XIQ48GBjO/oZaEj6mCopOS0//xtNmsQBGu39BX206gtQy7EgLuKe7qCNP7Ja
CzF9s0vc7bj2JVbW3aFdl5PqGrVpRC+eUkuuaBQ8zyNKO9YfCYkBLlW2SueoxpiqMg0NY4pd7V/0
I+ts8tysb4WHaNSTOWPnCgvlZ4WXq4RuvwoHoqZSM+8yyaiVFGSLmiNfsRNXUikv8iPMHw5O8O8N
YILx3M/G5owGLbORhnDfQB+6hLzLgseQvuWJHw0EPRvOnov6iK4Ljsf+aR6vJSeQLUUohnqbhgbS
6Rwl+w6Hbf8A1rHxUfuS0UgFbtu7c5dBybjJ9Y1mGXla8kKnXj6h+96b/2TLu0j2xD150W8p5rIE
/5scNKpQshlnn7xwCGByrIbVaDGqGE04V3JsRHmwDitxUYLWf4YwSYZVe/z4vfTOsNzw8MTk39as
b37mKlwIJXn/i6g0MoQ3jScqZ3HhuXg1coii/C41RcNdBSZuOVRbzC8Xjw0RR1KyDKlWLJ+PDUyI
gYmbsvg4/LeU0/QfsjzJ2cxb+W0cCpNoBwlENJVCqjVKVn9dyefGssQOSGT+a+q7Tdi5mRLBjRbR
vSfY0koylEuxntgQi8Q5kaZiLiHakcgxycmuEhuKRi9uB0isNq7Bc/xSmvEVho7WeBJWtiGCn68V
vtyi2wvCFGpbGFm6XzXjPJXe5tFKLvYDWrflDaj3tSpG5n/JyChm9s2X/5vMR5ej7X4ZObIoRkvh
yvnH8k8yHezwBNwzRJ+CHjNRzhIZQ9rbPyE9tdoFyXC6yPOYMFCV+mf1RsRV1EGLDqz9ZDHgWgG+
eYbNVUSABSZS718tFQbHC4U9fIOGxl5cmIsqYaBnRAsgYYCJ8MS7/uaE5MDzDQ/ZI2SvhnS765qX
wJalRgQwh6TxW69tI5ORIBWNl64H/Y6WXTKeWe0iLXjXPqublLqYqdcPIjF0d9pDsYw0zMcI8ic2
QqvMppmbI91nQr/fGueA0JyGJfLwt1FhmKIQFfwn+mpm9clJYT3NlZYdGY1lSNALzYyHQlnD5ScD
/4WW+Rd84S/gwbT3qI5lWEBeeeoOmidW5Vyj2q7gDrEaYueZF+eLBvKzTdE9FOsWOZG9aY7dLA5c
a+2yO9IQJgIVNPBUBzO9HCWnys8vpcJ/0mhApBQAb0hvzqQM/8PxCHiAIw+b5KcnLMTiv4D4lgZn
n+J5oKkNZTpqlt4AeAHyhLfGsphOKuE3Ri1kFXhOncKrlIHLDH23Y+vA3p+xFVWWwpfGgh+NpUkt
mjPNp1kqI5dIImi0X+eKm9aOR4Gro2IGS7wWYnm8ocNe4mnKSC/G9jSvftvca2H8UlLBEeBCR9bj
gduPE2u9V8G6HSqh8cujWXHTpwo9ldZMLMgtVXzWUjSUjrzEmC0yt2rvRwSj+eaKRJvd393NPjJU
+7577DC17VdM4DMoApWGuZ5ieY7jmhStfVFWsrpE3nBJaCbr2yHmvrGfsqAUkv4e/VZzGPdEY+4J
5lS9B2Lr4kIo2ItOwtFahqh/U/iLkyfk/D+TKCO/YCsCY19CmCmO+PMAw4DuneEqJh8U6n9IWBPO
oApMF+y4lBvbnXl3+0SPlcvHH4+jK4MiF++aGE6BOadG2wyuSJDSMekp9niQfUOIGlzq6jUbLb6k
kHKoAabYFX2NC0Dv4LvDyM25x/LxxXygPqk9yD4aUrsSk48AtrnQrn6SANDqGW8Ng0K+fQwcYpsB
VBtpd4gGA+zTvwhee38YSRM/sLYU6epoDOjt2lqFwlm93NlaECK+n9uvkbhdJrH0L7F3m5ChYTk/
lRLYzEFFtvtY/zg/I1nKHDp+gkh21tHG42Io2D98ND9L4TCyjJnxg2iWGNBO02Uj5c/kJdG3b2JE
pua7nHVLt+yn0G5ZFzTjcZMLk+Ih2gtBWxWlKEHQsyJXEvSEm7UnjJYd6S1I+WpkiC/UblXUFx79
2z36RRPGbgGE1zRkuzhL9mG/5R0YYD77TxCaPqPPEFuLFRD/XaH08vv+Ey7D1+NwwMU9ggTCUqyV
3RojpL/CAcpgIL9USlcXpXDXNhnDwh7+K0bZojpbz60bfLzJ1wR5r5Zn34ZXNI07E34onN/pHUKk
JDqDb7X+MpkD3M3sd/Ls6QVhXKOVcyX6J/4F6Njdab69/Jpv7/cO7VxSvfSJFf50vQwFS2AKvicu
jwjhne/N0PhgqMgP3kPR1kqScoFAy39tKoX9qNhyYnQd3iF9ZPQVlvYuA+vBJRxjMqKrxyMa1oqj
9IQ1smTj0y7Trl4lofYmiQ0Hg3flXqp1BJ8PERxmBd6/WRGRR8hvoGBAlvKamuclPhR5y7ti9Ljg
Oooq+tl9VoDO5BCdXhKyXC4VXS7pVltgKQ3rczU1tQ+GjyEKuvaid2GThp/0EOjxJGVqhJ0qlc2w
OCqolqLVcObbCHAuusguz7/IGSo95RnOMwd/EZIGfkYZJzk0ExvymCKP8B3UiVh+dtHQL/ptTMsd
y8/7K8ZVZeLt3HyFcQRJOHB3WCFmtoPwpaezyYL7MVMUgxR3x4k1JS8sT7Zz0n5iE7OTPbT0aGz2
BsNrYkkRVxO7oBa9hSUwPNZ7W+nCrvj4GLSckvrdO9b0k9RQjOJL5NnLrOxAwvT8j5a63w5o8t4u
RkmttZAkm+7oDyOhKrxWHabn99PR6M4j1zyC7z7QnsDEhWHS8vmXtQgKYHuoiDgiZEmA+grLeTxp
nH7aBzuE+CxA+AXOJ6IZyeV/ywONMEQ+My0/7XTDnoZX8MS8nPxD3DIP0q6A+5EGZ148h+ChGU55
+7wH4sG6jAdmQ/NpF+SWssD8kS5arP53Yuu+MOTZHNMKsyjcNANZ9mVNI6rs0C4qE7kLcu2/4rKt
lKomxvz9uGFdnDUBC5dvExCdvksO9bN6Geg7IHM15Nc1s7dQLnK67GjncEbWA/X9PMIax6NhEPqE
RRKhKzMWz5aiDwL20WPbcvWwhh+Z97SLI8JMfDoTKzq3HAPAm4yMr7vs9HnjINtRu4CktiGzzDsZ
S8F9UHTsdG2z0cJM9ePY7e9YEilm0KrqeDvAahZU3BelAVc6RolIBfuWFlGBcQZfHHPOpp77eO2c
bErnGsG1qKZX1vVr7xKXTXpuN9+yKrh1AhPTKRXEpogm4Cl/ahWcEsi8Ph04vvY+vQ4UcT6DBQDC
8zMqHmczsfNrUsAK7vUIDfAkdQBgkodhOE+dVX2ub2BxEtMFjKTxDr6FPytWbmp3zdhm9mqXhzZ9
Uxc6YW5WuT7nIhSOtb07odd0/FWawFTBVWdwnwVtUemmsPsMTBtjb7HG3eTi25u9/AyuioEy5KKE
WsV+uYfwzhII6HpEv0Ess2ZbV/yFvNneFmHz4VO47FtSjzUTh8re8mf67E3F4l3dVnCsjIWcRg9S
28T3uC9olUxNgwYyom+S2si8FhA3LdoT9yz9Cym0JISuJHoMYFMzNABqR5297pkkLjEbP9jMElpj
huQrY+KLeiQmTioNDNX0ZMSMs2d7wzgBOigzsHTB+lfnZSmrgvw7H5HC2jhqc1ZI1Hdz1Z+529eF
ccAZFXC+nqK9yWon3/q54n0nriDmF5LWZNvZSOxZ50UJdMkpBc05z1NjT9mqZAAC99gyhx3wdfEx
jelJrfYemaxZVmcI6xi6jpPS2htckknoFr6gE7USM1Ft7sgNsdmykdKk2iH/NTbFDM5rKL6TJ+AZ
lnNyd2xeOfQf4l1WB4j+D/byZ0t//mTUNCSVib/VLphkXPNc+rr2uAFyUk0u5hw8nKsqyiYWB24/
QWT50/wy9Txywv9ViQF/+VNtX7hzTkjr0Z6fMa9stPc1cJ1kBevH3gw0lbjGm8ZnhEx11qd1pMbt
TpAURyLiSsW0E6Cq5X+3BckbyhN9zcY+odh5ElhNGBuw377h/2rlOZZBIizk7Qzfj8ni+zUXEKR5
a59o8hZXODy3J63QNatvhXy4+6Rgrbnhgek5otcwZr/T4B/Bc/yPPGw9iEv2onTgzEt5QDVec6cp
crCSHP+quDE4SRkARf8bUAzgxCKpN807GlaGBj8Goy2pHER1S/ICe4M+9SwiWdwHafYl/i+eh3Q4
sB9iYd0dC6dDIyXoD/5zSO29F5ugCy4O2mi4+HexLODQ53O0x7+wvOf8gKRQYRAp1I6lwLdk5kiS
XhjtemfELrGyru1Ko+DY4XLg0TkfFRnLsQDqabSFxr0GEwAYIMwst84JeM0U1HACQjhmcYhjyGqX
aNrlo4MV4+w0BzKo3vRTCaAKya5U/Pu7jVl9JcvkqAk6zkpzbDf8BepIe4yzsKi69CPF3/lj6f4G
saeeZY+ckHy+kA58tXHG3eqM98ocLAzoGS+4weXavUGmMTcVlqfuyQgSLQTEH7r/ePXPDBDMoWbg
9FF7k4tjf/84nj5D7Zk2+IGfzoDeAR2292J1nd5uDDZH/xGV4pNqp6+JEDpW7uGQ4h/mo8Fg7Ykd
B8+2V9yWajdjgVeYyYlHjizDw7PFC6VfplMOjhYP9N29UQnHGFugPBRxDc8vMlalOPm9iQYLjE3v
LhVTI7Z9gkSuy54LK8O88PUCf1igaHdVr/lbOSNCefUkyLsTyhe6A9bDcWjitAL2puyi77Px0YMS
iOlaogP24ZbM7f3sQEZIrTcs2u3JCNJ9Bp9MA2K7xFa61/XgKEYLU/eUyUFijJaBf/uNhVT89GrO
US9StIX5aUgpwixbIzRNMC/r8DLSHGREHorx9ExwxMvZSk/BjYjFRX9oxRwep/nwYw/wdn58qoiH
pe34ZZMrluj/rvmqo5sVRJ9eog8UBJg+5tZ7hevN51hyu8y7EnF3hIrAz6MsdmV2RNRTGNEdsoRu
NAQvtESk7CXeHtOMOjA9Ofzyprur253PglTR9pA0P2jliezfnNvAXlvfRJnixYPDODj8HXR6dhpf
vfeoLjsE+cu1H0ouv6/wSIflGZrlKGw5KwnZMZwFkYQ2YU1jmDUHdTcMsOJvDwQ/ct0AxHFkn9w6
GjoIod3btKWpn6ENUvFl7/B3s5Ccw+yXJcXnZqovfjkVGsaEmag6aTxpl8nl0i07v5iaG6rs4BF/
xtJGCAd+IQ0Bsj6U0LVOeIsqYUVt2z8FlNY5yxLBuhx5gLLA/fX7j50mhXjuGFqUMRyyzgCfK1y6
WTNyDWZCRQOrNfb04X4DijiLqccdZajFivhqij+vYvRvGZ6cAlxjUfGj6slgE783HQcJ3TzFOJ9X
uZ6tc3OxJOKwn9FolqpPFup1/SFIDq2QtgILg1wbtBpmF6G7ml/UFVry43Smmz0xLBRj2pzclMFo
Nr4x0dJnpeF/zoNpaJDeN2ZjfNAfE/LkeUDnk2lw8Eg3V04gEU24pc7u9F13MDFmvNjT6/BJqOVW
bDKJKXZK7cn9F6jQbImVG4Cip8okFE9vrNaN7J0WbfjAITwJo0/mMuNUiCjiIrYXGH+ZY3PzexNQ
YemTfwNa68LNX9SxzG33L3QrLrNQCmdpzAs504IV9puMCOIpdbHSzEn8MDaq4FTuIvLT1bD2kHb7
SFuOKv/RN+pIhe72HvdgvReuTaMKpkwM0ZBCFtjqT8G9thmnemN7J6bYgpwiicFFG9h5FLswY+ZL
hLfNigNfUzUYk6Z7BygWR/uL9NmTFBT3EHYanSfazzhKRApQptKSfDCDP7M5P7eGu63cfXNyVNYQ
Zx/DHFVXzRWEmNgDL/T/uJPnhqph51AwlFgEboiMoPMVZ3RkUvWpVLMsKQ9f318/AA4xoeav5is3
MUSpAA+z6ICMScX9vL9nTCzD/vmqrRWN2NCLMq2Jh02WMYlMnThZGvrM7i+Dc4BkwoU5RqJB0Zap
6TzWvBw2TlShORo13eMsrEv/5hFAlgtTawi31v5YDwEERBm0TzXgjFZyIzZ1nzc3yFWfiVm2ZBm9
smC3RFB05dDm9/T1g0HLuA4KinvWErilyOHvOTnVLwcOiZSXvhfnOIGScPH96oXmKG+3UHcsTxUJ
YD9tbE7M5Yuaw2n/il4B6QFZn2VZIudntXgfN7Dk3oy2TKACosz0U9TVERQ9A8upovq6e+A9uTIS
/sVhHMffc7LamSKMnwWnnidR83oQhbEvIzSR88zvRvpfHPVpRAWoQnYR/THGjPw/dE7KNEIrH8+X
vesK+4Tk7C7wo9KXATO0A5kYhZWDO8KsFk7GZiD8v1b9mdmyIDJr8B3p3OhPtjbQ1/VkaOBIR/kr
R35gAGJTVznx/E+pkrBacT4Y8CcBWFBSMTzTLheQahlNZqKgSWEsI9CpqbjWigMfB9bk3BSzXb0Y
wq60Rw8VGGbnl727zCCMvCXg38zpHfe/kkDygcb8c7flbx7kr6iCOsnTbiXA9j+C3SBerY0yAniR
B3OYveqrq4LFur9hYjX2LsgJUGUm8iStaBDmJs1pjyxPR7Y5k93HBMcMxxtLP4RCAFUGeg3a9j93
9efGX9fQNbeGLqBo7NlMPBrXVX3WEv4GBfmunuFyqDiwZVWR8SmeGXumLYzdmo129nR+h4rrtMfL
tYvOCKSrJrUS6a3X80t1nzX80Z89nXcrOT1D3weWAStWwLj2ZnUiG/B+WkCeTeL8ZcC47shAiBRO
8N7jjD62Wdy4Ab1kvtswpTaaGsQlIBkifThXOWNSuc2u5eY2ettcMf1zffVLn7eIPgoLAry80OJX
ocy8aB4G5iNYUMi+yFDbPl39Gz/wefzHMEnqigIkdanzDJIjfvKbfGbIIi66n2qyzZrJa8FM3fl8
Eim+OyxX2FjRAhoTwDY1VL2rLr5eA14AejOE5IaPSRp03z2c/zp2a3YZh+/RN4aD1hWc47XqGo9s
tR77HbsBHld2HidYk4EFrpmUFBiho2DUFkOGzRBaQAC27T2zs535ahRPAVcKOaB5iFNWTNBQmtBW
hsqMHbj2Zl5LpbTGo/66UVrJmqDMe8yoyby8y6drwAtDUkPp5KmPHeKr+GeTT0mLH7/i8TnrvsP+
umuUJwmMcevJ+vESvSl/4ekZlDKo6O3gRW0n9gEutzt2HGnrQypWmantp+rsC325hKeFP3DadiMY
LeYTqrfjyFmAqsemWXx9xf0wnzUsElJ5qVr6q53ziuFsPYZqTeBN0F2KZupNSCxrgsZPnCo5yVYv
fNVwgv7Sh4ptBoVb5eXopwmsu8/TWxMzLaDM2ScXpAadqfYQBNIypYS6CIDNloiVWPhhdwlP2Mcc
b+w79X1/NvoUU0kKCAQaR6CAJaJWEj3k12OxC/f/bWYBVUHe38evt0TtD789LMhU2Oyzp8mIzc00
Ki4FekHpeVyDGW+MlSvXSKE407/6JikHqcSzUUSllQIZmcSI9Mfcp24EcSUJC/uJcyAHei87Be8v
F4sqqBJn/pmWvEYvBK0W9gOtCxGav6guMMundn6WWHdgNuvNvStpA+sFSQbz+ggMqvpYnUwBfG9+
gGL77QlPp3Zb11EdRSM5W4fd/T9IVMuw5wjaxZqcVgy19YVpfrzjno22rUgdahK0SDwzKsHT8Wo7
ovJuDWwiAVDf4Qq4K8qiFUlhAcqQm8k7YngzI+7ESgwyqP1vZEB7VCJTpdZMFJLvUnqDRnuiGjMn
Ufe5UC0ogaOsbcvKxN/rjL3iT6TNTeJdfu1X3EIc8oRIJ8HKsGUR5QlN2xQNeIjneondkgaKMQS6
AYRLqQPYx/35sLohEM3XFMw68Ai3C87ROoA0bzpEKXFFjiZqSqnChNQuJp995XF1Q6Y97yS7JQY7
ueJe1ExIhNS0st1jE5ZEbhY3XRqTGfgHzygT2bUtlRtU29ALSZQhW85H7MJAPGxpcAp2tODXgCFd
TBXfrx4edkWJ1U2Qz1pZ9jpyygEwY+drIvtejn1eY6U/aIYP0SyrX1BHZINel2V3KA60WCKUjBFl
jeIB4mQhATapTeILuYQg37ciZUlBASK521v41Wy9LfcZcTOrQuaYB3kWTYCHDD/2MRXqKVCJehTn
CrNhrg9nW8d+4P3L4UQNAmJRhtMnHxC/P3yUeWGF3quj8euT3VKtcVmVXYMNxsI3Y2YtFMsiJZhC
aB0zorU9Q5PKgEwmkOyKSGQqjt4S13NdMq+yKQ/lmn9gfK2Lw28DfaCIPEwROU24pOLrkh0NRusS
FXGYPC9VQojureg9HSHpC1Trkp8fEEHZZg1mSi/xzbxh0kAssBiRF0TpG55oX4IMMvxMOBFbN7Ya
9aVBPKhUFGsFmIuHqCKlZxL1Tf7MvbvcvAwGiGPjP82mUvFMw9sCNWla2EMfYIPfLzdgmHLfNji3
9g2vGlvjJcqyO4vnyYEz6awm+m52sWfSZ6VQZFmmC45PDem9qNGw2uI64OfYi6AzrnE0vj9dpK0f
tzvtEQpWP/2sBa3jywpEL4TVTBDEpOcVRK2IKk8AW51pPvEqZngBhTWsLtuOHD7dKFAmSp9S/QUd
CvOX6/iZ1h2NZq7XRMTjaOYfZ0CqClj09xb0uYhye7MCUuYpoQklMoR87gVrJgyEMP8UxBJf2SD1
vtqgw1sZUE0j1e+HlI+XKXgQLzQUuQqPpGZkFNwVRi4u1P8wa4j/fNQ7xHpa5f/UYq7XjYvD0Vvf
qiAYneVwAc7uvGtbnEkzbVdHYNXizpEdf3vE/4nat6UH36NARyZ671T7In79xq4F0xR9d3lEoKLL
9wR7s4fONb/QIc9sezm26zHT/Z4px6BRRMmJ3XQME2pPED/nI6AJeWky5chAJdB1q9UMXHhCsZPV
R4hrXzZ386bP3Y4LX6s+3tzUX0fe/j5UGPBz+hx4mLz8NOSN3EBob1+2sU/aoszIKFQqTrE2joEE
MkAakWIkPEJ7O+bJ4yf58RaFdvLUNEuP9UoNwdKePfj3Zn86lNbXeC1WRWbqlTBuu4F+1rD3jb9s
/3ssAzj4eC8y3CIVL05gPDyHAAhyBwIuDq3rqfv8o8eCyvCzw2oaW+gOGGV4S1Lj1Wpk7oBJOLNb
mduxTYcEhffKdpZOuXgnPpw+xisbF+xKopRa9X097QS9t+zkC72piayG/ZRzgKY7NDBWTy4G7JIo
RYj2NhVyeTevf+hxcOpJ7XGcfl1e5mAzhzonY6Noce7vo4Mk4hz11ZiM9j4sSxEBzwKgeFdHbfZ0
QqvoffvSHxJHouLCi/RRpob4CbRWsse89BSibE9wu3Eu/eNhcSxh1RRQlqvf1XyZnsuVg3aV5Ds5
1FE3IMfI2PMkgtGleDIK9ggPI56xCSqbOx5wywN6hAvFIGZCxWbdzclknzzL54g2LwQDBgeIwf6f
yBacUlVhM+jItsbfGkbAO4vL9S7udEOEB0T2hcryaskbSEE4kOV8A3B2OcMbf7i5JphFha+ckh3s
hsJ5EHx8JwBeFrOXfyo2cfHe/UZfNFxoE00VB0NzKvbVBMjjitMQAJaL8awwtvz+k482AfRKyJzF
5mpHkwkjtOAPMiSLlCymH14wxP/4xXbDJ+1ts6DR4cChcboZCzmFLEzgp+mJxy6rvlxTSas7k4TH
WEFz4APqNH62SMf84DQDVLj/nsQN0/fGuOqrPh8L6QSAes5amlsir3VDsGs1EMOZsn+KRV24dfBx
l+435dB406gSCvqhCFyPjxwsujlMrpKnK/WfWHMGYmIM+Epn//LaG/d//c5a+YLSCsLnS6HPuPyG
B+4e/mbTYX4LnH54CICe/LJnmeVf32pJR1CEvttZROyLw876nwnw/PoA32poYKbiPNuJtbvysZhD
UmbvWgLpxLTHJx30d3FA6pFOe1DOxQ7qTdZJcbQ0TrLvbSeQfhasi+nF74CFKgz9xLtkGO8wZvsv
GDJ6MOE4S5XKtlHvtL2/RkI+xxijt/+8lNSUJGquwk+ln+nKp2paVyoaExD46ul/v8iRQv8B5Chs
unJrXy2PVlI7mnIVIjnpg3pWTrr/cbIOV4wTC+vjhA+MKiyTgS2WFR/48SeObL3FW043wMD+kji7
qkJWr7Hqsw/EHjNGtdPCHPdiPYkGHvl4g8EnYuCY4m0g04dwbS9F86t5P7b4CbynH/MzsF2WXSLE
oL5lOFHKxSpd/u0P0BO1I+cDZonHISLW1OTceeiBqPmYvkWCria9jY2MJFtt3j7yjQJlG5WSqEqr
U9hRh/oKg+bKtufH4kD2G5Scaz85l7nw10h/bXFvMs/cEvt6HipnhDZLXJbTbzZWCz3syvQnFo9m
i+2Ev8ihxJ9i1rpIASiVMQ88QqwDdjp99blICeoC1sGHI/AL1ke8XZMMtR2yvNLJUnWxllz/sM39
bSVr2SjGL66MrzkKo8iOnwRK0qR5GZ0SatZmWQy/Jt4LMKEQ+lVgl9xKKODkjmQ0ZaUI9eDQP2wl
aGbZSopEdn2vQxztg4mxjkKLPdWx17cLalkIDBsjG47SdcN6fVyiQXHp+tS4Ha6LVkUhM6Z9hPNg
NNA0vrZvhhUM7ziPdIfJCyRmbwvkgvlHsoXDya+NKMdZBn0zP0YN7D7dvogih5yMCunhGe6UcAQ5
fKt9bUvm8HxAfqG3N7mCTa5zMUdqGnctgbLL18RqTd1CQ46jDg0uQBY9A8pv8vHa78WZJJeaMHdJ
gLniOIP9r4Ifu2+gCx4oMylGv3iQStJt3+JQR7DexU7txUpiwiPOGvSE5Gdgy6yj+wYURzHVNxzX
mp5S3dB79eeiNZ7XAcBreeIr0GbDidGSujJuTh9nbDwYp6YHTvFRYS1onBY22lGmqfnjG+kcImVv
wUUvLBal0zUMRkDxN/uiT3JoJpaqIEcQhCEJJw9AFu8BZ+/dXwGXBPu0Bd1mvTmxVQyu1YqbGoQC
pTh15z36Tey5xhz54usicNf8fxFTWP8z2OWESPWuXPTFnnMdT6XvJNh7QBiVn8C+MqC0rYQhdG/G
ufUHbA/2pqIlBJoVMpCowAmDmZPkkTrefrgrljWhdOLuu9dY2ZXK+/ZslcQoBCuDRfv6+kECldYg
BjylQGawRCLCfYyBoND2SjKjdkCH5R7PY+3dFg5qqP9KDWmdTLEicRvyIO1QbqJnfvwms/gQashZ
3o3rxqREpUFisTMRGrjIWVMpYLE3YF/5/mBDmU1sb5TZpOu5ROhOkINQ/C6Eu3ucDpzYP/m5mbZX
6KaRwVAF7R4GtXdGCz9Bim0/toNo/a8ckRId08MwUEYHFtvvS5fO2M68CemliEXSY6kdPSpsbe2j
1EeisFR3ruA+FN3UvKrzz4b+SB/eNzRMnnm1LhLmvQ6MO69XSXEX4von6qiLlIK2IAlckhPJWyui
tVXf1yT5eAeQQ4Cpg9MR9kLF9pZG5SddDTwWIe8Btk66YjnWnHQb7qimPckdDaeNek1+ThWOfM+j
J+Udil7Huza1fkv5VctK3vnS8B5c9ZVUM5lR92ebh9Y9ibPQO1ih9kydZ2+CgSVZ3dI86yoci+tO
13R9Vxdri7EB9nQz7EG1tMQdFBqpdsO5oaf6ZidD1HZr6dzl2eGc0asmprCP5BLo8Q/nUneHUs/q
DHCQqIw4diIJRRsRy4MLfQhqeFNacsirC74LRmbTi6nUv5rqeT2+s1IlkjO859bhAWDm2bRRaKnQ
KAXwHFbL45oDiIhDCXByfgi+t/PUpdpJUdb2DIXleC47ByQFMc+JXEHfiuDCMsXRiCqmaP+wa5Ml
pa2NH1hF8OxYUpnKrYK79m803pB0QW7thyUCxLtMTcCI5s+Qa0T1PzQ0DmZ0Jq19daigu45QSRks
fqTF2MRe5bf1bqVpVIE/qFzHS9R4gaEYzsWXkRkkYXZYqxw/R3OgXRnK0csDKXIb7IOzgRMAhB6x
7Ep+JnTUo8czqdCJ9lpU1ofd06eIAeWFGg2mtwG2pY7mj5rArccopooSdnydSK7rgdccD5AtAVRS
c4hyqyxHOgOJYvMUrQgFVq0P3EftpwCjJBCAij53EsdPOX0VVbLoXUi1NaeLpHJ+O0k2WQLsk7P8
6bOxsVyWRJKyV6IrhxenPPZ2ilpoVuxqK6iMWlcnwSkWaXg3vg48nZl4Ch9OxcB2GuegNrCtthw4
FNqjQfs4+Tr/XZbUZV6oD+okn6BwbQFomwrsjuemQ+UD4+uiWxrEhf9zWeRh0jGz076I/4+PmyXu
qr7oLogZleLo+DC3KQSsnMAV0DQpHz1huv8XuB1A9j5l/wH+7WL2fR9+EJNjjKtKgNklqusmY6W2
n0GoBZax/sSFkU/bmXd+XohwK+Oo+IZMfwS1H4c4cpo22p2Jt/uyowaRxGEeKxAjaDr8j8qzSYzD
p/0QCru1d3njSnXI/kSFtpjwIA0efYG3EELsiROBjhToB5wLNTUTcCVR4kEg+MOy6JYors6yuP1Y
nAt9Vm7j2pmjp+A07QzUcrSdodRNsOSBeU2GiLENypXy+IJbxgPPckU7duVNEVeLRPLFejGMDuA9
5T/eFGUL40p28orOaBS9oNb4f1GjN4tMt3OwsyRi/oODj2yxfmIcdCG5+/z5k6XeWJAUy20PLNfM
x/vfkFydEnvVo2A1J+msa51ZLGWFnJ/Zo7zuuO/XKxuecLS23fiOrOojfxLkpwQmRpIFvy3z0Vv+
R9q5/CiEOO6jrf3+Z0Sn5TwrvWblbC8xDKgYaZXYakdjntJkHqRNIX611lATTLoRmjtU90B9V1QC
toUBR5TENmtUm+DUL/XF+9BSSslGQr9zWKD5JaRzKi7B/eHLnDcjOtwQbmPfWQCP96BcQqPATiDX
Q78UFTohUQqASYU/gYmtrfBePF5RK1k7rZ+k0PPvLk7ZkbltsH3+dUJlZ8dBC+rLIr2Resx79gin
4K3mzqDzXOMpLZLeEK1llreiUYREouOEzgc0aN/KblGGN7jwSJVSFriUguiB4hpvbgLFEa7KA+K9
JUmgPmEqJG5ROkmcqr7XWtbflQrqlR35iemAqI4ifzLD2lSTwMfgRBNgz2e7uLVFUKgT3Nj78uNV
sxTArLQRml9NQJ0cuNWrWsqAd4t+D19B3Sne01g4bKsVsnkdn1yOvEWMdNrJb+nt94NmpIvukN/E
malPDhNIU1LYb9L6zP6Br58s4Mpce0uhWM30EgiLVvBh05ZnDb1n5I5bG4QloyKFjTFUvMLew9RB
45Y3ODdbZx/uYhAgGHaazelK4j2cBA3M+yFwANzhVdHFd376YNLVWmXhI1mFCYiIzwhg+WR6X5m1
aMf0VUWFUvgaIvUqFrU/sIXRBagYIXWOdKkXE2H6cLCoYt/BAoQ0eg1LH0pq7NF65nbLK2iVx7GV
6W+5ZKeSwJj1ainvQEE6Iv5u4GHjHh0BejUQ6d3uqIxvxeYpKosuQu5OXoiFYSbNL4Y82Z268jBm
XoKPNsHnbDhbHLFfpLmIxWn4K8AXosaMznAtysw8cObORwfxKZIuv3ntW3dmLfkiBY6ZasEJJR8M
YNIuKgtCdR/nNBOlex9iiZlfWPHr1rpxYjQfraqCFX9KDxefuZH7evBtITG2vvTz+vDuY48QHWtK
NRL/HPWZkWWH5UcdfMBd/wHzza4lTHZ7txRT4yVG/QVw3ISGH7KmRb6+/5ngIAiY3nuCphowiXKt
9o6gAUJRrLeZRD9iNhsg/3qwCq026cIHjZZVWAuw3YyCfPcJ7igWF6Ms8hIVi7JkT/pIaQy0vr/V
ox1Z8R4XFdbWLIzl1751LXpTMMIeEZzltPhJXqpReeQ6NQ1HQY4N5YyOEVfOiT/Qc7fjb+pYaJmE
MKGr6OTGHcs1gb5g20fBwhExj5q3d5dzE1uhOkswf4zot1E9z0I22oZvSdoz8KSWeN1hoqACk7RC
TapSgisiC5Bghlk39+vI8P2XzZv3NFTlH8ybOI8x/FtHfuoagnMVDdPLgoRksbPSAmq1IiNmLMUO
QVBWyb/xIvDVOciRKzOsTc5YPKpoXYmgytyJQDKvJwbeysn56iXyYLwu7zCesHefS70JOQFUIVLg
Cknr81Wjm1FE6TZL172G2aOAXgk3f1WUJRlOZuR8UkWUGEsBp9+0cexYPL8FTkgfJtMxUJIuvMMP
Cx9CRi0Nzqjn5dleElx2ahWBM+QcQeFJb3DZah/B/gDk+C2Y2twFGAxyF5si6mXB0efQOui98jTd
KNXR9ZnZKrigt5HTmGpZQmyeiV/Dq4vj2/c4QxqeAfgnF22d0kj+2th9jnDI7mIharU6kOUyGabN
OxU2AQb+5BzjLuvYRPpvy2/T3w8jRIhwYEnxNA1bgSWJslaWDp4/nAYArPlFjNvOZMDAYDsIxNIe
9e4QIAY9EbDy1BVviRTUaCHlSVvRSZj9ZspMmhAAhi4DC2Fvrpz2g411m4RCD4lCi0VXEdH7poia
OF45jke2A4mKWUhz/6FJvzvGNdJbSnlYi5ZFXT/ueO61tsjSh4/zxfM3KfzjLmX+VMPG7YbzeSgg
KeSio7wMnmi3iwO8m9klFgw6VSyqThkr0cCcNA1Jm71Jxxox0hbvemaQWTwLvXxH7CgzUp22MhqN
FnXv+pm5jk8XV8hOwAkyN9pnFeg03ymcO7xA2abZ80ZQ1dUHJueKTQ5AcaZoZBX2qMzVWOK5WhxJ
FkO7yHqttMF6ESgPm5zvwLSx++3QJbSQAmyuEbkEu2zfoM7bg5GovE5arK8yiauCVsj8/XEz1imR
/efcyXDjl6ALiMh41x80VEM4SzhcUy4UJiw0ZfrBoQ7doaP3+NivCvMTN7BdibpwOiNcWcq7nG7r
bwyMojIR4LjaERBLfc4mW0jtPmRoArLj6dQo1HHLvhPK2VGVVeQvbeH4mdxGoNcqR6lBrfoAhQt0
490j7RbkUigAolL1MWpGXaHctZG9soY5/0V2GC12PfFt3z/SOdQFOIC7k1SA21zJrrwtvY9zPH6u
1tUZz4wMLliRdtwIUCQtB7wINbSQMImkJHCQ4XD+Kx0KBihfP78jFyiWNFlmjNsDGa1CUgrY+8zl
o6SezbqVWKO/FKimso2RC+nB/OYEegfhv1gFekZoRalz+sWOK6XKxTerOktnhPOgGT6TL51E0ptF
SqKG7BXyeuc6svhUslmJ0h9UQFu2L4MxHsMKfA+pbpZaimTQeEDX/pnPheYVeyu2t5yWIS8j6WE6
28US89U3edc2m4A/B++8F9pWrObxDeo41D02IwyBXRXSb970AHeX2zWkWj/0n0fktWU1Q6qww7Jw
bHu/hNzS+I/sMSrSHLeRBdoJ1VNqSOmPPFSZ5Vbxk0uXdLhSwKOeexKAFvpZj3RFjdatLPGAw9KN
v+tjBNhJxInuDIzrQiCC8BzZakjXY7LJKhBkBJA1V0yYyIhAQ7KVm/lBHXMFH5k5VYAkR0eXMM/9
zojcHxeO4sybtlXp9aNpKMS+sP3vapTy6KroKKNZ9VPNounEe5mc/Ui1cK8wejKMKRWEPSJ9MWwW
bZKcum4eAhRHVaMWmGoM2TIZuve3G75cOe5m9Gz3wUABdxG51G/sNFoLA/teHkmOH3mWsYYAYz4B
x6bj3/YGeEI/hoT5IJ1kSJ2Zc6tTR84aUHWOmA066/rJRMjAEHGgW3USaGAQTjLk10jhIvepjssD
uw/t3RXQr2XH4ivgk/18njFZ1ea4dY/ljDszJGUAyprbqBZsowuOnnrG75+dqiJDOr2ZmGMmttYS
Hi7MBm9hOeJOicSDn50qNJijb2TKbp26b99rIY08uKry1oXnO+iklWoDULu2V99rddDvBUVCcTzO
ZqyYg/GG8h2KFcAR9lkoCnermmGYcu2+6UT/j/dgiS9AafyNkacgQwPrDzBcZ1m+wTBIjO/OMi6q
DawAvC8ZS7UABvGw6GkuCbFyTfu6jsy0H80DQXjvXw1LFUATH2JcfFvEmOsteopPbq8tnRIVk1YC
l2wr/gMJvYUOVItzLT2CRaewKQvmtnB00uUEvPtoNp1kapxYcSzp3Xt14XNAGsJskzJoz+gYF7EP
xwfy55IcIllno+O5+W9iv6YTQ1X6Dq4fMWFV+ahHthnlir3Zu7mZ8zBYTRXu4I6rAzQFTJ6KRyLt
LFslJjGGJKgxCw/+Lvk6UMb7tJL+qUrO7lyCq8yyeUlTNT0lfZQCKKUovNnP1iYb9DSNmpVv0GU0
DYwrO7MxcL7Tant5M07+LOX6ygUEEGVmRXrQAVunMwHbJuN/qgAj3BzM5TD/mxo5B2JeAQDcft6r
jIZikSRm2HQJT/XFPxhYvNAeDU1LQh0e9k1dk5EbOLyALrSaElwspFUvEZXF2+S1AQEjZ6f8G6r/
XU8tsz2aeFGPVPULRfJIndmtITl+pjaogynvL/9rOrF9UYSXEbBHO9vDpAH76shiy8J8ekOM8PKL
44LwG2FkISBxJp+4sgPLb2QMcrKSk+bszGMoxpNypU6Ia0PrGIvTJa05W+7RVnn4Gt3tqDuTCg3y
dhq+NhjUISFNoGF/xpIdTFoqIRml5fZiIeT6W+XHvTJ0fDl7CzWER3Atv3AvOwOp97xvS4kMKPh7
IWH7vw1/ZXbVosw+oVlj7T/Faf0Dwva9GwwWP5S0MGSlf3Vf/Ap9Vt0vnuFKY2D+u6UYMUB7TVnj
u9U8TIu6V9qXzfJvn4c0vbWRk2Q/RW5Q95JYsrbNen9n2J+HQXQ+Yuy94AuX3XjRaiErbio2vMkw
+S7eet0Mm7HyXv4UJjbWiIRiyd5qvq3FScv83gvxISc3q+wTEMz/NAqodzdS6oRm9jG3Ye/GbASV
qaCbapLWok0KosVPaT+C0rMQnFsETTIw3LzePVlS4hnLRgjuSiep2/yUXcnL6YD0nUIF1U031gQS
29q6IDqTtQaFN79ggdf5NAmjeopMS+XJjTBBJA3sHyGE6PmxicEx/aI+i7O9Ek5IlQo02zFQTej8
9V/N+9RQwon8TAvtunmQ6n2d7yrAPgxSPm1gxkG5WaYTYlFivD+elWTmuGuY+LEpbTDNPdREt4Zr
MbWbptn//sgikOTioKftQpdu5g2hTY3fLD/R3vNf28BmW5NHCX6ZIE9tgHOnZcvcX7er7pqbJNXb
Oersn4Kk6yYok6a7JmN6p7uwyYzYSUnGcchxcVH4hclOhsCrlKW7DwiMELYXpEhk6eZYMJG/GDLP
FjKLOBx3A4af2R7s9A+PzcLDmanN7Jk9yi/0FCr3K+YIPdlcX0/WErgRMIOjGTTXRX6tbSLe4tM3
sMh2ybflzlncKhEgLMxM/JyfjCFQFLxi0QNXC7Y6Vw+/8guq/+Fxb+R7/XdGvLhz2gn+dfsUCdez
6U6SM2VfEsWevFKrRb0dxabaEI9SCjQIjCa/2gbk9SNe2QqduprMvOsUx6H2wIQ0doXNSSnriwGL
BW2N0s3TJ0nYZM3Kf/2zzJ5iC7cmDPZSgzVKgX1yYby00JOT93ua10qfSqUOvOVd3ash784UETMv
TrTQPhMq5OpQDZdL9J/MG2yH/h79VDiHXq/wsDRmWKy+r9d8gVYjVVrvj/QkNu/C0FFmOZyohPs9
7tcavSjoQ6GtdXPx0BqGXKxqJpMkDqw/1faFjoEZxclBPzWDKGpXrJBtqu2HhJJIGc06ieaqJOOB
CFacmQlNyzfTzVJnB5771TbCjWQbQd6rIIWwxcE1qpBwlC7wze73GaxkixFZRgFssw6Ems0kbhv0
5BVky3AMxEFIQiJKNjtYx+U8UAk62nky+vtOOrczWlW3ly8eK07ST/gPys3TY17Vgw789gEyBOWt
1GVeILYKllL+8ctWBX0jTah4rHhpQ65EkJ0Erb2JgTgPbjtcTyjkq3cOE5QGeb+EONWVnEta2Cel
Cfpzn0UwqRM47fUficK9bvQemHWVpoLeW0bhPDfjYU30r75l39S8Sah08BCwJmMkzn5yxpK7caqv
dljx/q8cHOhZA3KmvM+ls3YsUNnED5cLFsfdeKO19IxIZZc8xgkRPAP/NgiWwltuyj+j3RUaNnvm
hO7N+A5Li9A8tcTZ867oL302x9GKRvL9VibzvwCbFIBnWuqvn3JUWgBjb0uSf0ncfb5JoZ+IKB9F
xIP7bbOaV0+4WFZsA1gjrQF4pp6jXE7kOAj51cS1mGjL6n5toCqmvWIA8T6dfYoTiObEneE1dCfp
qFncI7hGBELys4YQQVzB7MF9aagM5zLW/VCKze5vjHexwzxKDIKApaLUV2D2VpbiItcjBseRfGVQ
c7vfTxrskzrEgxGgEsespJJsdCfTIjDBWm7uBeQKA2OsnwYNEk02Tw6799p8KGEadXgHEG2pqqxl
5LwrYqfwZWWveUDfsOgjA7fCHUMMBg+PGsQyxXgSaNsEu92H3IRC1fU8AvwNRJn9q7qNqLvauVvE
JENhpvSXQ8TQfUesoO1iJlWoAr8TfnYP+WhkzjPpb7SbvFO5v2X97NKsbuoX+fEa0lJE1lIYzHuc
HCJFgKfuZBkJvFOv+KR527LYQqPZU/pa/hnx91gl4yqjP4luxubG/Bpiv4vDfDPtDGUo0qBHCOQA
akW4dotOcEpp4CEZpnzRDLPbNrymTA/Nxj2qWoRxBgnURFEaUw28v9iOjZNapERn8PSTadVrnP2Y
ie1xr4bn51zcuUFAsC3fUww9KrwpQbZf/lrwd7X+Zyy9S8rAMavH2BcZT43BdESpampLPeIrUsuf
gWPPOgAvRNNbiazOWA30kzwnwb78phDtU5nC52x9jfgrvvgHqPXFlNokORBc7EHl1KFq8GFsd8eT
XJQoux+wBW/lLG4msfTttxMBmFbhRJwPN9TKDf2q93P/iQuZUVMuUKDFag31ND9UnCkv5nvpq7Q+
NQEXwzHhMrLD5Lt1bcNLIy0RMKIgIbkIMThFbff0/GiBTghP0zJmB6U6cjDMIe57MG9neN6k6UGu
kuN77zX07cIT1pLI/n/Po7pL+WaAcJevDaUUxP/AAzEx5SuEhxC5HVYPwc1jKDXmAi7FAiIbCet1
hwVonUvgB/AhdRHNRjgpnP8tTsNGFVUZQX+l8kMTGR4+8vjBYpU3SLsxN3S1y28NEc05Yhx36CvR
MpioV2TwXUAKC2P5Rj2yoouQynIYcBCflfS+Vp7JtXf7+GdknndD0JA0q8ArrWxYDXKvfuCGh3I3
tHVyllR4plo7jAwDyhtmIIHGUgV3kCI157bBjP2NffDYaT3ECBIZGbPVB/3t1tSBfE3EnhDzreQh
XMU/gkXom1jPt64HjaHQyGajt/CC4d/sMktdNKExbOE9hI6yylw6p4vtJgxUBkPk1i/n9+qZEeuT
r/WGJxD9IlEKsv7eKMgsfDLJJyAaKS2kyvXHxjiF5Fb7wgWLm4+GxtJRQ4lFGdoPTDsqf6jkCl7N
7YueHEVBNfgGrNxh5tD64BEmv1v1czjDv9SJEpvpwGzMl/6r1CCbg3EyTMuCEqGlAqsKPO4uYGkv
CHPZbFGqKxahS7dGj9zBDRcSKX7TYsBWdUhqR9JrBvy/DBXQMm7eFgkjqllz1doB1oCKoz3zK3uY
aKR1LO7j5a+z5Js9Eh3K9mZ9NDF7cJw24KjtcvxsdsICKhWOmfHiG3GxIFAc2FKv9zbO1wfQx296
8unL1B3wjFHdN5i0ngJtszwBBqjKXgqrHhibcXMFNHNHE1BWYGDrHzukGeUGhGF/yPfpCB09ydaz
Dp8B69saZrry6mLuBX6ppGk4OrkQWAOzFDvfJorKec+0VRY+HZQ97gwmDhbXzBGFpVHrbJxDUB3W
u93jiCcVKwVuYKuMFRRUd6n7A+ZczCv5p53qQR8EUhbnuANGta863RbjxfSPOu1JLNOgSuRrWci1
xQZoB1L0WecIrkkhW4XUNCt3Qd0DBj+FkmXRkilKxFMwgakDhRTx0m6ldU/nhyBnUX0vrm2URc65
+SK4wSG9WrTU8OYmsCJX79WQbIjGzV3VsMO/XgKkD//Jqs9XlU47azsvtK2U/EsJZM9DNEf4z7m5
dWppLRG7dcmi9F4IogluaDa4tEYA0dkQatRhW0XGZ0ASUUUBLagIO4DpTbkRCVwuxdEF/YMBRxqx
YAj6RYUXxwBSKV6fvi5WDKEYDDTUaGfi0c9zTWVzi9NUusq5IjBn0ccklcm7Y6PqDSo40kggeLF8
TaXOcaXXrs3Z1YVLDaBmbRqkfprXJs/lrq8XaDHlxFp+oZ31JO8fYeLw+8kDNC2H0ZXoerwdPnKI
FmgKt2kv4dhlzfWMInm/M4y53pQDlLHTCCkyEb+c6fbZBhvhA2qQiouyG6ePSWdN4Qna7pOCvd0J
IcS+0Arumg8QlXpDPGSdk/vpk5j2kKCJ8oj2Qa3rUqTQKJq77C6/VMv8eDF9D4pTeTpEU3/lClsg
ZwjxkthZbbH2YV21LCLrPgMshJeciqLwQNkSql+TxDCJmvyhwyl/CWIVEAk/1gjuCSWQihNysPW5
ht5MI2MPMOt7vJLcAvpBDNEKBR/Su9YSee45aFmuONDC5q5h5Y7I2xCxKJoeEcREsjFU0ThiA0JQ
umQYtE21ydJIhNO8BvIutxmXg3ZOq2BSEa17yLwPJI+VlG+DkKTUms9CqbjHkMWr/lidCwohzRfe
XwCIeCku81g2bdk5EO6r29bPH2Z0WecJXPINUo0TFmrw4UZ+AV1T63ODTZE9YuZXjEtFZe3z2NUl
R5lOlIFbAXZvSfzngZ7uVWWDhdar4jwBIkgAAIMK86vzOG27Pd66f1J5Je9ESmkgB+AHLb44+WI2
0/waUutVdGwNQkCLHyqYNW6F9u+66XoW0MYpgpZN2QGG7zrUKMH4Istgt2Yf8CqRymeak3O98AKw
AGidjZVbQyDQtO77vJqqtSVgfYzEjnO6ssraIxW8KvxYQ0PcL5y1ydV51yHnZm5TyKWzVt/JAP53
B+euRhMfS23E6RNfbWRQviD6AROoyy2HMCzcgFA3lN7UjKUFHGq5Vct6eDZaItW/n2fmJqGVVUb2
e8f3zIKALiauc/AifFCaYa11uc+DVygxZ7v11zg0vpmaoaLDuZyXmJ8NPVYpW1FZZeXzNr+rBpGk
QzrCIJPCY6+o5zPmxG2trknrcNh1++aIf43DqZB61YPt3ebDbywXVxpkwPwlw3eVqCszNhzBylxM
P2ZNvuCLY0hpL3X0BRN57EdvoWcz/mT5Zf190PNt/iThks9uSK0OwU2aFZG8JAC8yBO3PLWogBwe
yr3uR77mITUTlp3xxcyJKeIPwJMJJSBnfB7RadfpGYk65UczFJPOja20SA0p79z6fX2uUiuwtwTu
hpBe6NpMTgSXuEKvsfjI4CXY7VSCMuo8Cgwfxf7akFAoH+DRm3nvpYq9OzV30Swu7y4FHHZKlcuR
GrDG5Z33R7/p0H8Bok6i1fvkS5lhZpyJu5hrADXCNzbhjRCA0g1iA9VwauBTd3OOiZxgBtrC0BtS
Q1E6N11ZxvE9c6KSaMjL2f/6gPO2QnvZaqr3TJ+6cVgi5u9j8Kl/mk4EPKe8Ev2RerhJk6BuT1lg
Z9IeFqHy8NR/sQTd5qKyRv62jtME93B1eD2X12oCgtnZRy51xvtRhQTwBZSptolxToIPy0Nk0j/c
BL8lSau5hUfaIdf2dZn3o9zLJ2xRZ7VcEkrhm5XIf4am80rPHSJsF9vD6k4t5awpvcoF4hyv+Riv
+2cx8yxH/TSw0UQANwz/XS3QFcNrirDKfP4u2OM/a/5xBNCe/z4bNqN1tBEaoSxjNe2o2Zq1Nwuz
cGjL28U+qx/fJvYJEzJBAnMbrKN1/woLNQM1CMRGj2OSx6G576vdD2CJavtvtPK7ee627D5T6m49
cWMpAVYuc2q6d7CeS7O/sOsrF3Sj3r2HgcXfPyAFiaKXhvgFrq7s+XQCq8z6pWqgxwIZQ+I+3apR
Jg6POHR1mFwg+VbKDVPI8wmXksXyapWZf/5ujquFSbrIKteYFZ4GTnSp3jFia2RACYSQqFkdeUfa
QZpRp3/xSwfrXrbSF5P/gX4c6EcJhw7gZsIrYiSSqYHO5j+ZOLUopVKrCsw/NYy2YpPVq8d4pzKb
ccDoL8ta35hclD1dEv94n0tkDnTDUPoovlMGEvX50cAxHdpHHmtcKf9vZ3Zei3fKfpIHkUeCekpg
wUOdc3H7nfr3Uhz/ZYT+XTLeKJCFjqXed5ONHHDpCBvAq9lBsFc8h7jJwmi0zdDTI1q4NqLwjczL
iq1qwq59HVmdngGlt8Eja5txXJzkPQeokiQ7yzMaL1+tVVMBG5QGEocQbXSG5JqdgWdldLwAZSvG
OFXu5SqRPPnhqYgDHrnw1GjTxTEmf6OxWv4eOI9kmPM3dKlKr54TytXmH7HPhOtGGcon0zYw8x/O
28UIKrSHtxzFybqu0IgdJmUPEhab31G3CX0t7yl65mg9JilAFfl0ZhjV98yevc13Y2OY1Q40CBjC
hbTdJAlv7F8bYwtSosWuTqYKhL++PTDyKhI0KUwwPXi9TVUlTIkGTpRE74S5F55YmzSdW/d2hJAk
xgVqd9MNK86q7WgXEU1/OpgSdgmJq0f9/wy4uksRS2N5jIiuY59utlS2UMawU9g5jIh6ifk7yCve
zljn8cjiLND3Lt0ZGSGKkUPB0omSgM6OCTPjflGs7Bpctegf/32ug0p3hPWc3wobNA79NvpbxALu
E+nRREAa27AZHbdWRNylmRCDOAPDEWQvcC0TWjoc2l9HL01kQVijZFfLECFwuFsHoNNS0UoYnxwO
DS4jnhCnCChsE9GgFnj25CEvicyxNiidvHaYGGVQgUocOetzYkfD96e/dI9GKIztt/Tvj3R8XiIO
xZhupkLOZUYAWcmLAnhV+gG8JGYVCLjjo+ju3fuhD7D6pSnoD6Gg9KN94ocrM3mVDFhFNdwVf1Qo
P3PHAL1UUyP8/FYfpQ5U5t1p+FT0PFNvJLz0xJFnWH2zogCVX554vnIn9ZWIR+/G93vufUSMRNsX
ErkS6GRO0gs5fJtDL8UIXVvCD2HDaeBkpYzqyJSf7xlkGod5QmBABl/jx6OOs50e3IRPnROHfq1m
iStkxWFAPpXyWni6NX/IYEjSjoq7cXYxgmll3kDuasYwvph3tHj4He6c6XoJDGdIIX1odjcI7gub
Wg498EGOryAOFd34t418yyweHsK6P9x6hUne7a1/sf/mwXvRRlUElfUwZZ11nekAI8NPjMpWc6ys
SDykhWlMQhPt5OcRH4Mc70I7aqIhOZuOo1gdXqJh2e9ZpaD2NfhmpPidCzbVSQXbDAKHLUnawGsQ
CBWp0wuqFrudFogMVyzg5VbtSALIsB3FElH8gHEOiZqiu++M+D7V3QWrsLi+qqh4Rrbjq2o5XM89
hdfrCgbd1HLEuypd0iXFnB5iyZIRQy1p7cu0YlC8OzcdAiE/FLMTnWI0JLvTqx5xir1o4j9F+1QG
uFkmVSO8KyME8A5MhTCA0Zk83SvgRgNU0C3gOsmA911KaJw7LjBujHAQWVx1Cfxo6H8anfe0rkGF
PEo7umZgZahAU5FTgWsNda2IJvc+RLmlcQMw2YS0eEnm3aMgGthbGv1Pc4VTHioiftXmKCIMFyNO
2HAek3ShUhSlwBNetXVNlozAZPVLDk4+AeyCCmtusXDBoBy0nzi9MgKO+lvZk33n/xohKqBWY7iM
ZGJtn+V8FpVzFl2+Ax9VYQiCqvvgvP9GjGajPrOq3qlIxmpv9NeMspugEQN6/IJqBkqzqgFwcRWU
An3Kudv6pJi9zdnGSOTFgTyrGh+R9SssrLtMA7DbmOzITlwJJMBK+1MGBhhPnm5Lfq62Pu8//Wzr
bqRW6D/YRXJMIN0mFru8yVYNWCJ8AhvybFqXU3q0N+KnOQDpRHr7tNz9lBAQzbu4P4MNSRI9U5KZ
nEKGcGgyJ2+e+eADWf6QyZazs0i7xuIzp1JRzdJ0xoQ3QgE9LICuLXfzUzcT4voGjRn1gBiBQI2G
Cbu+SIFIQki4hOwLSoEjZIFFlBOL6SdCCTa0WvBqxQgr9jSCFMlTouF5vzsFlqPqMOtoj1B7On43
p6M15l5IAH5jxV1kb4nO2BRyEm1lgHBbWEZeMuPmUbMaEVgJtg2ajblfmkYjfsMVHcK3I/R62lZ3
9N5dgj7567nlNd+ifo91y0KpKOWGtYDWNSThtMiTe/FZgRgiM6d0N17nvRxSzUzO2G6oyWHQJfGT
OpOvYF8gDo6jEp51GM6wZsvqzuZE9JmmBG7RrSFzb5pxZ16AYB0jq9xyVZ2c1afYja7I6QR+/sXJ
d0AplLkIy+8DkxjInICQYHgB0+OCzgm/HRmQKVKBzYuBn2dBF3/tZydPH5MMv+2WqIu/KKoUi69U
GcH1J0bQHUNqXihhAVbji+qjlwkXl3xeJF9rHU43iS5CrIa4HqMVc25Yg8SQM87dIq3M2jICfkL0
9vhwb9T+A2z+C7UYu4vOoQu6Hs6jNpD1TqLM04vtABbr6DBmu7HIhE748QJkwKkqMpxQ22rPgVFq
k5nI8ZzdnqwE3kx5I4uGQ5vAjlnbsXRhstk/IKusxvd/cRsTFg3DlBOsAjTQ0flunVSwwZ/8nfCw
uJGlgE9+xpSH4MoejGKS1ecH4ftXNBMQxhxBzm2vrxmtjSwE6z9Mr0DGPVOgUh/YtDYrAO4YdDEr
bSnS9Bi2+gQygSum5HmXHVrEpM2jXXkFcWw3a4TYUa/cZyaPE7JeyiIMAUClDGdjJ5z90en/Gg97
YrfTEqgGVin/SBl/7oWF0kn1mdbUgS2Q0w3zCnHNV0DlnYB9TKDW2LmnGFuSFpYls/SnQx//zLQj
swYwOiCIdgSXO8ApevFHeMTttGo0U8c1NuJbZtRdIuhEep7ufmnCqWa0w4XSNbpmhqdEe4gZM9W9
Xzx2ZHBE44dswjS6KX1gU6t+ntFhHQnjLnLDevvQc0YpiR0muvq0imS6EpkbdSYlGdBa5LohCezo
cZm+Ez0Okk0oi6UlYiDZVS93hrDivYiDKRtpswb0vAtXH0lrXnGKOoSXrq/fKWFjdPPaFXhaJyqT
OsZTHcmMqD7sFlPW8ganLokgT8k7KgsBa74cOz+tsqeUwDrrqFMbj5tFDfciogIHIHIFEvdPGy/+
n0tJY2sU2CM2Lta/Bf4sMZSUnkKlmrZx8SrKp+d7Z+kvBVqKxMur3C9g/u0j4r3ATb7TAG1o1egv
PJ8nYmxMpCvnhO9GFd5c3INN7CBA1sZ5lUCMdsynoDHrLpQ6bCkiFFIcALVbzn+UtaNHd1EOESl3
DQ9Og+atkQk50K0R4pCU87nXwuMlsoHGJo73/1LwK4fdU/CveuOXVTVqHu2Hm4DgYM32rF7Iq1v6
5hqn5CIdYoFVQ01/GmvQrub6yUVr8NB7r0xWZIFnYOiQ1iignleYqAAaZpVwv6m/+SAVa+xytghp
SSvr5pI9BZISs6bScpFfon8YzDKMt5WjEJGJE318hsHXagAQ5VlJnnzeKk8BnzAOtaMVt7F7duk4
DmtNK9CxgOISsi2NwkL/ML1jHmo/htpvxO+aYi7VeqDd9x+Bgryt3WD5lseSfyaOfyxLQyJ0aIdN
jfUubNeVzsz8+vjADu0bHbMTPWiLMsbrwJNYDiJZmW8g/ufJlOij57ZhHdJefFdMVh49zDBTEixs
bz5/HhKDJomxV44YUvKioAsodR6j0uHNDYQU+CmPA907Y0rux7X41ugyCcLqN2kmURIKuDrbUkIB
fqUkpSk5blFUB1JW9T5Cikx1LmC84VSIcVYq8MsnfCaEkFVnHFWGmQwhzvKCKPwpnnhRiZZdr8/M
jF0+SpvqtlgSeSbRydYEJQAhdgaLGbzVAihry+Qy5v35v1Hu5/IdKxD3JkqZjHcUVztwaRa3ej22
uGEsCGjV0XRth4u5V5LxucCZp64nuf2Oq7Ly7Faw5ZVMvp791ZFx3o7V7sU8ZgrKSzm5HU8FUztQ
06RciX4iBRZqnxQUHNMzWOlrgWAR3pdQx9XQ8auKGyu0FuadHSu8cezk/XOYhNyUpYgwEeecRcVx
Y1UAWxMB9DCTF1LJXwEBivocXK+aavWSnOBSEsDUKwQbHyiCuBIKiiCbpmU2JfrKALohtjj54mwG
itgly3xC/OVEgZRHtRO9wPQrseIEbeXTjBD4wL65VRxJWbsCf2fy5QJeJWYS1PffL0Rij304Rno8
78zU0zudoSNzh3AOtJZMgtD3zmaosHcIY7x4F3TG6wx5wN0Pwic2SgUWnV+Kv4c9SBhCFZW1KmVb
LXA1uqUPyKuxIyvLI04+Ku1BGw43d/OJ6B95YBKDNGYelOoT26ebMYIBTHKQRLHoCAILsOkKzUsv
0Ob2XgXLWo7jMux+u9+fmu5+JvJOnU+uXlJSHWw76tiPGmTGpkgeqVxyHjeNXQ7+XACYZkDx8OWF
ulyaDRNczICvCfxCwd6QETQbiDy4r2zm6JvA3L1AxfeMVTEGsls8ksS/J4m3Mhfl7UTyEe4JVhjl
KfL92khDyrjhCc3Pbknf+xpWTXQ+k6hrp6E6iIezvhH5UMJGH5zEpIYkKeD8WsIqn5Z7cyT0F5MT
op2ayew0lJjGuSd0mLd3R3CfTlJGSrebTr9LI/fqOT/K+5bSMWZL8vOxcCkVR70JEX9O9m/O6SsS
+CQU+KzHpuk0eq1vZY0R8acvI2S8i5y3gO/78xzcbaRhuA8N7zFHiLMC/znPvSRHsiOBirN00XeQ
oQ/pLU3LWbk7G+ckIZgdfUzEfvj5QqrBf3pqYI7oQkEQL4/ijYAZK7aq49BsTqFTl2U+73kD+fV9
fUUyUkiP3gerb8Hhx5bah2ZXJj2NiEgw3vlvAKgDzquhVZkVCDMwgmrZGneAoTsHLVRj1bk1BOvf
zcUlxY/e167sU1SnBsyEXh0/Bvjf22Baz69zRAuID1PuPll+9l52gQZGtIHHsMJG/QT0axa6JhGO
r7H1inUOnwKZFRhv1qvhzv5AxlRnG0ssKI7aJYvVI18K7/bHSv56CU13r/koPgwLJQlOEKDdlLfv
2txFob1EgURPV4jMokzlSTTgTOVfCKKXdVufNomnAR+It6zQlJH3ZARtARFS0vLa8+iS7YjVmayb
Ji3dIh1GA54VEEcblAo7EcZDbYkc+nUryiAH/29LrwXKdPuR7uxjjHEP7hpxg7HNkhWEV1TYtI7i
DvpdMrE+ZjLMi4WbX16LrX/m27SiLSxhOcDpCs9mr6PP7nu8Zl+v904iZFx0EOuvUyEYAJ1TnzRo
JMiuXvK2YTh3NKHFdApNRhakR4sxTEXwCx/OTzDxHk1240T6bbVEGOvscAf7bczD1SpsqWgdabqr
mtr6Cp+3PAH5hG/orYSIk3u65B0l6FhyVLG2N+dWDgbb39+7VjNIOlEh0CWzZRL/tRKdN+rff8LP
bvSnxI0d4NYZqKu3FAGQwWaVhccZTmxbMHbgZvy0fIxr4Mnt3jHqoRZIL+3CuMUlSLysWubqxmcn
JIXzZ9a1xDes07H94x0UmeHs6RlWc6pyi3gYe2+ED3SKfcJr6u5UOgbgb0L0wEQ/9Uha+opzXaA7
M2VMADVf5qeZmvYruYi7InwU0ep3hil09GxVIv/tq2468vznJyVfTxupJgBsrUX+RGd4g3kR9nVl
DFX2VCskAXBpr7k+3dn0lT+QuNnrXr3utNnMN+OJSELLZG0VAsLkHYKpcdR1u3kTVEfGOfEA7nzq
+8ec9vSoHGpsEc8GMKXfC7ghPXuddpoDcz2AZ7YWsbflQRdGA4GA4oqwp/xztrA0hjPsAA1ooXv8
XMEyTRGdPMQBAdPHF0xGX7rmBLigeH7RxJcfHnFFu6/i0TSUMGkDuNHa1hZVW8G1sBKBhLtmm2Bb
ZhijxHr5KBuSS/ah1eUV6QyFvjy3Z/NWs+1NXXO4aRpn6gT6gABgmU19r191oSvyNPVS1BQX2L2V
xPVKx4rtqKlPkCOqKv6LScZQScDzuaE3DGub+pO9/PagUAwZU9Zw1g7upl6Ak0b8+qKyGKwk4MVc
qSyMhLXrtd2DhBlMnmaRN95ksVxnd2/LbxMxS62WAl5hazbtIRx8DPZJE05FNrEtFj7fTlGJ4fAW
aM45xX0Eqps9FbBU/vuykW0k7WfTD+ttbSekpfTqK76ao4HfLAHG1m/Z+2iR+rp67eBy+h6idGBw
3k9E3hsobPfS1WPrdkdGH5URROS+a1rDHAnVBTJPCdVTPoCQ36POpo8O86iad+qb4Iv+6bl5kKjm
+ehCr+huKaHeOCnOSyP+RhVWTaE191AORIOriDOd4jaQUPzbNFVWxt2hkVaWV7A/LJaeOg2v9AO0
mzGGBDlTRL/aPmqFCDD6Dcy6d9W57iPIJBqilZe2xYWKfQQF39H48YMDfMuMDwGdZwK0CEbQNJps
BburBjNHFCV4BwssGJxq9PxI6BljkJFaOhC6/uOvNeFyAxXF10HU35hneYKQayKvDy1wu7HWZyhL
1tk700LDSXQowpTHMpmoJXm/whcu6YTqL3IAiuyZuszkQ6snR/9e2UE0oJXgrPwtfT6Rn89YXw0/
mKikD67FtFeUCgSF00PMjV2ujvGrXX2E36kk/ahQO24FAzXmOsa2iUmn/haV3NlGBvGs8U6inEfk
QwQWA0MGfy3O/QLxqROM4kI/dM3IR2Dp2cAr0hPesLto3K3cYIYRi2WpKVBFwu+5JL6teZ4Po/ZC
08nx0OiZDNDkgqP7HdKLvPez8b4P38iDkn+ySYK8ixkdqge8UJE+u7gK1igFDrgisC+z2rFk1b6f
xqR6wak9oHOromirvPGtPx+6IMbzPYulr1+M6qSajiSUcHAuYbhkxTmcTqFf0ymzX1qomvqAFZD/
qdM3Cg3folf+BmPZpRuu9W0kzAZJqGJw97Y/hyYyU5DJrJT7VvkMC//uuBmHkrxQtcSu/4cGRe9I
KzizVf0qht+2nX+WuNdhgCViy+1zCJGQy9l7N9ODCYuIvSiporqyLNaOj3vdsfQiOLww3DLWo8P3
YdxAlFVZXkITdemUJQJvJKjVrnV2YdzV6IcMCErEsAB60HaXRZCycMDNRKk9VAIxbWwRr7bQg7tn
1LX8vtvdy7MzzK+CMcZtyBC1reoOgilS5xFRT0vrPkk9tWoHq87E3D2RamCmHTqJRiPW86rTQ2xC
8736mgDA96J11xRudOleJv5DPhd/S3V7b4JsNSIBvmSuitxeMKMGqh2viokqom9OpNoZuybAA4eB
95Jtf2nOHRf6DIrGO0KHOyQPACN/RgnI7R5r53ecyLRJcsx0PU/mV1nc9k7yLggd3S0gJ+BKBvlS
C+1VfcH+QkJWjOjGyXHePrXZR19jdS4IBo64CDXvTJGJyRhahR4sQQxzD3PG0K6OYh1RSXmqMdrZ
Iz+FzKlZNkPS9/RPZ3ysyEepMawAjyHhdF8B8rtaYNh7RvE3rpGLfOji+726rPZiVjsDIVayBe8z
1F+CIjMYzieTiJnLUtpFu1NvnIXfYm50YIECUrDZ3eosb9MbOFJzxQbkuCfiw8y1hQa0lcqgcmaQ
ooubXEoyctWnguhhLJ2C2+ukx5SJQfUIf5K61VeyxLjlD+E0Ap8UfpGqtv6c9ToMYOoyLIhgDCo1
pfUnN+qWA9mLOaaGzw/37g8nThW3h3eoq9TDqB8ZFqFRLkKR9ZVh1Of7nVqh3BmR2E4fkk6bkjw0
EDXkB8VZgF7QTR3OomTW+BcXs2lLkF6LmnRHHb4Y8dRoFgeQYfQMcF7DE1lbgJYQ+mNCMFiDcJ1r
s61RnusgOhOFkCFCnzA4tBAZTjJUB5QoFZqWBppdMktOHxmqjTy4AAMrVU6a1jKWLFE3elNk/cw7
D+Pp6FkbgI68AF2WMKBa4sfgvT+eUGFJcadyhHVmyv25iiv4oGeoItjWBgo8TBdUbYVKHPe2SUgu
Ct6E7t+nAIShR/AmQoMu5fg1o/vQvrEBGHJUhZNiiuJsnr9CZLH7X26lFyzXxnXN8UPsFJ9/pf7E
Nsmcjt3f0/0QsaJWhUVPrMHfsZesTU3m/5BpClLDtP/EYUsHS6/h+W0849KcGPsSFYqiy7xEL5i/
/THgdMIGKLsJ7G/BecsiswKGfH9eHIPNY3DhfLjWcaWppLhpXqzyJSj+UH+morPbRTxCI/DZfKo0
cVwjPRmV5jjLNXsPuKq2MXYArJsvri5FMlME0DCnesLrLPDul1yHVt4hrysYpeMGIfmH3hs9FjYW
euJqM+0/KdYVd6Ae7ow0Wsj9FrkGvHJxRmUkkr8lrhtcauKwFjG3TB6pRJl7w3KDCZewUw6uMU0H
uzkYGp3e+SOBnY+uJi4sO2oxNHvHftYXgGNibWhb3bQb8fEhq0uehSGf1GEtuhaESuYvF5J6J3md
FvrSZfwhDaKxzeBHd5zw1lovfaty3mUxSNv+f6Z27tVoLlZ3Q9eSfffVam/bcnVsPGUzC5VSyTeN
6h3TjdyjMNe+++hhfnT/MFRrO2RjgJxmWKu6a3SWM+RfPQHn8MyV58J/lnizcVP7Gbz2q4/3mH0x
gHFLzNS0QS0fAAIMRMNK0AGXOUWvQCdCGw8vBJKr9wb/wMl5OcGQazznRIwc0L+xBBkIoUr4z6+a
vipKSDOfgR9iYypDix5iVX8al5U/m6ow0w7kN3gIy1K1dDl5s/LF3kkLqEGBevOLIoNiy+FJoqoi
EVJKUAc4Yf+xy0zboZy7MZXfE8dgIqniTBQ/d5PeRXvserdlNHeUyQ1eklzznUYdllkS6+BIdhoP
MfnNARHdev7cO1ng/at2fzoI3akTNmkepVrc+cm3BQG0mwoDiX1Vym3R3VQzfix712gxQzT6TSaS
fHqBeC1+ZLEiHeEOJ3eWOgxF9NS/txNgMkNCH3lDhWESqGgb/umIaNFieD4xBzQjTpNWyldcZrVu
R/FGZN3KVBCl4r5I2XEjSUu9kEqL4yLHpbg+CjIP1duFQ7ncXOCkUWlPITie85MomTzewVHMOBcD
wyppDrpNGckuFMrBskFBrM6d3HCjan1+vPe0EVmgfedB3+Gz3lD+hthiSxPCzCxzYkGnHMNogZy1
nXiLYHSd31F7Ij7Fjm/9y8SHUrwhWFsrlcCqV/oW6xJer9++/7TrA233gpThAtdSgbx4JkjT7tKO
9zvWqUQbjeNPCvFrag586OdtkzKom9dr1sMsyX2gH9SpeKbgdz5YMgcb1TLW6HgFl9o9KiYHc6ZS
8iSSCxSx+JYHEdJTwud0w+E70CyUr8CQ4+5MZmuOMl2l4z4hOQJmu63+Gt/177FQ+qd4Oil3C/mU
9Pg8hoUJ6NMPEL/HmLxL4+Z6uSWvpH8bxTx6YiTx2fl0I6GNy/7Pbz+99ItLbcqG3ebqIIVn1zkr
BS0ol0b6TpWzgBQN2XDpEsu+FN7PlyUsUOkO/qvyT8TzY8at5rajuPQV1J/7KeJGPDU21Z/+4FXi
xpjfS7qqh0hs1cLjBGdywLouoMruayeob87KOe7CDScS9mnyv7B9tMHzjF3c5et3MOTiGTRQI/oR
SNMkO8SC/P2YA80zI/BCFK4W8miOUOzQZY0lEiWujJoJKFFh1gj6IwnnAXf4CxkYfvlMHBJwmIGV
CFf1dF51flDPFNUVwAb15Ep83ChWPSIcUZZ9fgHH7IuwRdiC/uqidUaFNqsUHJmMhjrxGNPuR1J6
C/14YIdJruGbRraCgTjqqP5Mn+0bx9+KK0CzlUjG7/VoUVg7/a+sFdh3GABXaA6bsjiIvW1wWRSd
yeLznm54hOBYEPSBhxn2zUSFrZBnpMsVsMs1ctus4Q0wCRAfZhaspBQn9/Soej+hjEDEGSfOD7Im
Z7pcPDM27zpNcwYKUNop2us6qW3nv4VWHIws2rrgAsDaz9mf8u7dN2QQWDkSxamxGzXYMAdfBTQD
kVI57hn6TdeytORcVW7YJvh/3m6DibmQBM5TbkBf5lAlqJNTD+qCpImHYe8IHWBNoMYkKoQ63N+c
7WstFKOE8zaFtMnjdgeZkBb0WxGOI8+v5iGc6UcUMJacJpzMy+O4cK71pMgC0t2XjNnAcGD/6Q+p
4umS1Ih8X3VQEEDrJEzVM2PEMBHCvCbs/R1UOhL1fbGc967f75w4gZmnxy2PMhoOpT40qlcuirUo
/eoFWxQ+id+nMJs2XCSQf8BA0vWsnXr0h6TzYYn9+wv3M2WG8MIfnvGqn7agucyWFoW4YL2XnmOS
ni+YJcTDj8woFS56Me59pasZKHROnZTvAto2BanBQQiDCAIRMLLQ5WDIQQ0citzFabuHjFYtLMCo
TewiJbUVFmiGS6rcxw+Asjg7oXiVauCUloXBBSNbgO4oyPgobi17xRQSag+fAehQQvhKp7sK72dw
mD7apYhRynvkrFgmbh9xqrabBnoQAFBzYx2+ob8P10jgzmtz7xiBa9PQjdi7Hend1Pu9Tk7V6Plv
3RwM9HmhAheNFtmRMU8S/3XRI+KZ6Y3v5KN8B8mJv3b7eTqG7fzzjliJzrIqNq/vBilyxrUNq6nA
MkqDiqX6B61mjEK9ekELc8r6OP2Z0/X9qwg8F/QblS65oQPZqmQ2Xx+IWUXpTcFP4FQjQKHipCxH
xB5VPGMvRmKU2R3ELZTtguEILyQGFcFyAbriIB8d3nB5Df+OTlj7HeIiev+y5oH/68XJRDoVh06e
PBjH0Ta/vuYuW8yj6N/dYPK7KLr14VBZNDVgIQnSoHiq0VyGZwnSGoO/UxZcF8pbJHDmpJx42176
iYnpZokMwKhW04lbbVhm2aWQFitbHVFK1McpwTIWjQNRjtD7WkZMCBMRlo6qAmXyyt5X00Bj1TV6
uWUKHZ0anhn+YQ0t/+S8Yis/PZ8/bNJxm/t+xFrIYdShUUZs3hHKwHCZqnepGSAZ+fIRbhVZsbs4
5oZs3wGAYV2DrmXOvTSMye2GpfWF7Zo/3NdJRLCyiLwHQqi+7DAFvyGGi8IUP+ZKD41S9nPSqVP+
D5sLpbsp7sUzWVNEFIbjvnoHAm/dsLN6KU5awm0sVdt9P1v9GRxV1g8aM3PdFJmAA13ZWKf5GiQ7
IqQXMirUK5EY+LyqiRn/fKv3qHJDhLghVAzU+y22nBhjUjvxe7S+M927e9k8DQi1ZPrY9tbXAQOy
L1MCVO4FgVDMEkF8Rp4IBKF0fpHTeml9DTXhq0DyHOkR9/lc/g2DjUTm1rAJGcvIfl1Xlio8au+j
NlHv2bOYqn3vIE7leLZyO1weDhZeQcJ5iFyni7QzEbTe3v1XRZPekr8Z3mK4pfLEEyb8UXS5mM0l
HRbbFpiNlql+oTi6cfZS2y5x9TMZUQSXQpmeEpxsouMsRcOzH7OFe2h4fcZJ2iZhsLONHWTd5EP2
uuftoYjovaa7m1aGnkXUM8pI7t74huzsGJcNOq9mAuSoFMuSCXqpifGOeuyGjqmyZA7FyCkxYaS7
D6yUSnm603brLh467dK8Ri3ajOnjEMhL/Hf3DC1S3iqxo7m6KqIASK8tr16E2w5y16tngwVBscgr
iEefOJJfRM9mwW+cdn1nkBvRiJI+KlNmSFRRVq4q3gZMaWitYI0Z5sSiocXGQn5tM+65NoeNnOUn
bIhFjzNDN7IqlfMqHn3B9nlgfoRUUlX5b28//q8q0HWPHdgFtV4uZnkz+VIEu+nc/AtgGFBb5oJC
B1tuZOcwqOzt98dCPfndMIjIn5C4vA+bvAsjllHb6FmQ7fZnADqGylLUxmReRYa6N7eOvwup1JbE
bNDIcFjPkFjLECEVPPpQ/oHbRP8nWnjIkvKT8XT69sdtmE1jhZpugLBOD5UgdDqattE5fGDmGpWZ
EK9lls5Tv7l+j2yFLjm/g4Ra2xg70MAOmMnARZeZ3OYdRbEEuLK3b5IvLfWbKsY9vK9EZWC63jXi
Kzn+m4C8SxIOt3pmZLsosOWKKzTUzLehllmOR72CSW7MAIPf+kPpeijbylE8XMgKX2NJSF5iTmeL
FxTdHN43xckThI55eEzcbfkvLPpyP//Zak7W+8MoXQSlPZok0gstHV1oIqV0lEmD/fYDh5cTAAQm
xU/3kjr671De0/0gOlQhMLwqDiIqyUFBfh09sJmfGWMt/sLhPYmleZbVLVl9Ii2R7wKa/IEjy3tx
SP6TFUYpABACDLzEqRe7GaFeejOIoT3wbo7hltd497asRO1AhUPgHkM+vxUm0lTQT9kaCUXo5mlK
QQ+sljU4F5bWYpsm/pRHFmsNgphgxJflf0joDtp7gibwZ+Aclb4k+h8VEv9T1ptF4cuuR23We0Qk
G68TVoXfHw+LU8d6HnjgvYKffwpGar/H7lAlkXqu8a8bp7e9AazI5NnuNAF1iDXbo3X1cuYclzGt
xVSnB8BQCUBYU/IIVEX5ggI1COqxa9OyoNkFgQGNfWIxALhDgv6B/QRjtGUBMDczZltfvFRCTNSM
Ua/oK054xwssETbZkBgwAo7bNVEBnCaxADcaGLaHNeZoAx+h2rfMDaIqv2nXADBsCJ+ziI6/Li2D
XvzmPtib4MKXBLobU0GuYP1wv3lu41suXL4pBVbUU7dfIwOsrisVl8LKeyBJ4CDtvtKqCVUKe+CU
3LRFK6xLTyWAvwuvCclMbdcbo8sDtHBqPVhuyfh9OvyF8zKjzxOj06Y9BFQIfDdjr3GBOTAIenuf
3WK1Lu8XLSG0HiawrQmVzdtXrbGlU/xI2D8HHZOwf6ZPG1CyTkOtV9z4Ggx+FZA1rjeWCpSv4l9e
DMEHbMHBBqtY7jU71PpId+ZrHUHBYD/7b6b6cAMARCPccrW2/xbudmocwKu8fYybSIWlziDGj34s
j533hoVjFBGPIZkMaw6q/cJTUKMS65x4hGoPHWj5ZSde3jz4vmtHsN0lzIv8OR/g97UHupXKpQpe
kqb00ZSYSqwcthqXTWz6dygHseJta3TRWjuMh0JClqefDU0i12WdIevV1JZk/uqO3cByv/48l9IZ
SUIHYAV3SuA5OOcVPoK7gg9ssqjd6xP2TmIvfm+KCEblbcI3bV74oJ737N4FSdTjJ/ewpFs2/R5l
A8Ej4vq2C3KQezNtLxij7VfJE3mgW5Xi8BqmXIa6BLksMJr80ZgROrrC3r9XUQDZXb9ms7CMuzkV
AlpIScfvRjPz4SOk5fARcBPKkjUy6dfzj2IXsbowDPSgoV6KZakCUyzaykQyKsEH+XyqkTvW866F
SuV/oh3ZmwUr/TmagMw1oFhZALnLCZnomeiqVnJ5fncBO5kdRJ3s5oHuydFlwRbQd9pMNdvchQKP
4An4nLqmENXMhunZAtuQne/SocculB6oJbRA3oovflKBHDvnFnKdRxviDxEc2/wyleU9ke91aIGi
K3ACToPjlngm+Dum8yPL5hV0jgm0CQXd18+26HSfzK1+9luAWrzLOhwSuV0fSdQlc26fnKWc9SVl
DJCfqud1HMZCCDYRijirp8WPapJjxve4qKOJ4o5nXlyd/bl9WFDo2pBow7QPfLJKvzQi1DeiLe1j
Zud24LlMvwHOTcCasIzigbpLF3x/N9cUDM/qmOVrAMLAF7LQ1jRnIbBK4Apj9a9Ao7hdw3rAmCi+
joNTr3zf/X8ioH/lEaaqYTC+iHsQ2eT0JJaT4f6UPsCRSTfiK5g/JCgx2rdlFmVcIQJtLZ3EeiuI
lMSP0ux3negqdx3uL8alYQatVSsYh1KZ2aTZpZMFmxC4U5WKurY3aaVQsGruHdscbkOzdqAthkfI
rNVDkgw4m+i/T/VFPd4NhkRm2VeFc24x/fdscbJEbkLJwAfZvSTnra4s4rVxvU1+jzCqZHtLeoYU
dRX/SFuBolVKnuxcMhP7Xx29mnoLHRfl2+PC0KzSL7BQWqBor7FogWSGGkf5DW2lEc1kK35IgH17
XBTLJiGi9QfH2jN87HN846OBpOVVmrIOZe59GnW/nh10Z/ld1NJfNjvw2G3cGTeLRdRCGJ1qVlf0
7wlLFjauiJJAovivjvwISa++WNHBcf4oFLcH2mJYUcNc2pkrEMePFSlQoVyROH9isfz71osZFpxn
AmKpD8F8jBG1ex7xbu25v4stSjph4uSKrMv2HHGVkc1IfWe5TLxBElC+P2SFFefmgfIDRXVrlQg/
Pu7O7XNO0zGV67cyGr8YZRARJZ+njsqEucseTBKveAIz7yANkde4ay2TmYEonbHLqbNqlWYIwP3U
smwLwHfxb7ZpZk5VR5or/spVHWGOzh7BEDOWGPlklHulryK0jKXH+wSg4nqPSzwaxfCSI/hcjSGy
tGxZ7TB5FN6MP8xRPKOdzlNp/rW0FVxjgLK4HdQwIqJeIEMYJ18LfdC8stKDYKWHGT0i0IXwuWZ1
KWm3bpz5fKv9wQqZm7KY6Ob2l0l6OZyBa11oIY85FMSW2T0vUg7dErJeQnX3rQRSmKxnm5H2vmdq
+5Ny7ALbJtPtCkFNloLhxb44QU+qp3P64AXM65OvifN3vX1aZ6LQRlP72jHyNzmuyx2e+qNMBwed
zxYVkWDdq9AYBDy3bjk0Tv1IZ4wkalRZf0X2tA1SDfkM+k+J7IyFJ9irxDj14P63RMxS1e02P5ZF
zs4nQnNlE/BiMP/KFJ9H1nYa5wNVNRxsMA/NUBMXgJuzLqNmBCv/8iOAVq+14Ixk7gS5+KRy+dOS
lNaQe3VMLzzdwlMKcRam1CcTPismoE+AZY34qBVaKEWKGMZE9MoPmQQ6B/C4kMddwra0zQEbk04Y
tVIdIPetQlvk0taLcK4FgnUXWq8AfqZlX/FDbrcxcRK+yUY3fjEWjtVkt3fKNzHMl9cNtrEJCgSd
nj/yQMUePewUS0HAdOr3FoZrFiuvXVlaWQPTH0CKhTdzQ30D9XPZO122LExtPAdF2s8Z9uamXC9R
kO+vxaT7SzqkxjZX1iTA7lXOIRKvccgzvuy5kKy+m2POdSO3cuNTr/TMxdjgqC4ND6kHbIG7kGwT
JJf5/8297LJYJaXRpv5okLY2/+zDl7uSTxnQ/I/ZRo1kbFhd8rQlxGlA+7KyDAAhZXN1USaffgry
IEc07rZuEr+ut1TFMXt5PQr6PR+K5ZV4wibz4IGLrYGNUiDGdiExuwcyD2MuFPtM21nVB8rWbp2A
LIMPCrSi3wqD1CvOllxml4AeBtvmnhZKZJ0ORlD3UIbzcXL/Yt72T4iDp/YkzfHiSQeUb6zbAXr/
dl8HgkJcmOfiEIhm5Amvn27J/rJuejbdfRJZKO+rWgRy9tL1iwhNhwhZRKl54Qlwus7J6SkF7DdA
JYeIya76URFn0yXFZzhVfGTSKnYw9sUph96xRsO+SrGEg3N5USD/h2BlONbg6U/FHJP05M8QNQrQ
sLMO9mHpxnDSh883c+NsbSD4PcBgAoGzI3bMVBxqJBqezoUhivQZsyS/jvh/ZtyKBTXBj9LEH6nQ
XULm+K08cyUnKzPhpRzAyIdJJ2iSm+yGaiqzmKyURRbtGem6ucWIq6jkkhbXyxC8QAK7wbj8Mdck
CI1o4zFC2gMkdEjezFpkZeiiYX+mvzXuOP/1pio4u+yEp2RpVMBn/J19+3ekJINLcU4PORFDHqxF
+7+gorZeilDLI4fZqQt+8wmR5quyOCyNPmpv9WA6WLNuwp7ewYsv+MxkcYdXKn6c+lb+pQ31kymC
9gOKRkjkxwhtZS6rCwY14Eo+3BQ7m8QnkGzsNUMcni4Dfj9AJS/8mOAKCugKzBTHd5aFPF5q1/kI
/2mH1swpoN/S7ePbp+mYzrRkzcUpxUucJIHCWTg7Tk4L6r7oReoeUNx6qzVlgi8dW6Edqe4ik1uF
/5tQCw7/6nHToqijKnSiJJ4dvtuJ/wSeN/d+O8hdFktY1TiCzKV2GgBIT+d4T2M/6JVRBMCMD32L
pHdzn0svc0OQ4Hh1rMKpIUXfzn12eANbkI5cu3d1+yWXfZrG4eOTESvRqZo1R8z7iqisu67WU4xF
mbLud9nEnOBBZI5JFb6nRa05588sN3ukcpw4UtSdB/qINOl9mrMI8Kna9cRoMP/ehIYSGo05hoec
uuJT7Prssg3M5yGzNm8GvMkw4Jhp/5PDtYFBT5m+Ycvgk95m4Scp4YrZ4RdhRAk+Ijt59keWQUQr
B+Mm8naZgW2yBlv2LNgMT3iy9vAN7TVwHB0JO7Yz59ZBlgwmsLBE3Ltbi6aeGVFdslREp6JiNrbw
jsbfy5KhRH6xvLkdIcdaZhVikfbWkga4xuWykI3QWjYTtgZZSYSiYVjcG499BX/MogeoWzXZi2lR
5J3rxNv5tO2aega9vGfuWsOBYei12UDxq2bRm8NxKd4wjSKQe2Gpfu+eBkviK2A+dl431vAQt1wN
11gHbITyM18aXV3xSYZ8viKhMR7vOOla8ASnDMgxEVmmvPLdKMSAMCdwApKChkqgrXfajpywteuj
xSnvfrgNV03x/mHjHMXXfUXSRsqQAfFF7vf7j0UyGvMd0g/NiTk2jbIRr00SlBCtFssIn5Qv2pve
+O8qkng7xpfWRA+kpQERsenKQO22vHPL3mS5PNK3f3OkUaruiD06H8CNlxHuwqbXFBTA3PhwwayH
In/b+iv7XOQbj89cU+shdkgMWw7pr+FiO3/KpmYTtuGg7hUqcGNSVp8KFFJShaSBnhDipIyHZ7mh
yFshRU/9DNVoXuJrDg0cZGu10CV9qLNNvuahcYrB41ZYNO2ZxS0Jnswk2auMVDte+rL8X5lhmwUa
i38CfRIqXO+QCtXSflV7RrqC26xupf3vs5ePy5qfUB9wTGDOFaz6YIMCWByaCTLmtlDNvfjIvFX0
GIVcWXf4PZsvI6f4ZjuCOoW8xSBCf/+hrUjfcgy7f8oEmvgraaf8tRV2gExM6cYr9hBeu6BDxUlS
AcRwFrZPlnE75s2HvbIQkAOJD+S1fYta7w1MQkjiVtNwJ1ui0W/MJ17sqPLSWsdEW5uEHdi7ua2P
fZ0o0q9VFHxi2+l8mBuAPkq5wQNdjlDZ36hDZiJP4pvrP6ikz3xiZXA30nVHVvFVCX2nAGO6POKG
TBDFwNSt9OBLRmuvak8Tva6VjO4uK1IdoN+KdGlFLCFhpudST9Bj6Qe9FuOhJVDBOM2wqrSi1qc3
7jqcYwpw949dyPj5B4mJwKbTqIJWpZd8CEgtd2z24ojbK6NnuGlbOgtP0VJh93i6DgxJd+GIFUg3
/8JYgUFOQunC3IoimnwDdTDb7AgeTq6ApAgTm9hG4FUUSHeTpw23gJwBms0neJ5vbrj8TA1J6Tx8
gSFiZs1Rjt05YVbGFGSc2wWKX65q6S/4RmtJvHCNnCmxZI40uCM5xB1/ileq/VAUpxB33O3/N+ZG
vM1SK7hNGjwUly4uES6Rn8RU9sQqGqSEihuwvOagInpSCl5EfRsDZhzZSUJO5mLFZPVGzrK3hjCn
FvIVo6AxTf+PWK3eBlrU554HfCIaBQ/caACLNW+QwKVqHpJQ/cKcWeSZLeuvb3n8n0H1g75N0jXH
9aBY8Fy/7Agu09XApzN8Nedzk8wfz0QkTWyPAe3brkUPk8nv9DPZ8rK3RZn4R3wN/TdvdzaikVH/
zxP77cBu0VFNJR/XKrcQwVjjjmxaTKEThUQMd+2jJrKqnCl7wASqxa8J7oOvkyq/VFwyvc+XtzXO
JypOND2VNWbFGSI0CuOqlpgDFc3Rfz8T5OffGAyZbKrj8mTqa+3b5FbLXiEoyOmye8KJ96hKlNpY
1Gks5sxhY2NFeM0jwtfeoBoVfgjDpfRt70EZoOqgNO0m9stmg85ATWjTKdx5KTuRUk9H/NgO7FZR
b+sjP2r5F7JQBAiEXs+GpqFS5CiFm7krBM1IRju5dmNx2R6RZ2pWjjZ8gDRwc+ALOfTSCbiU4oVL
FUvduhaOtVeHwPdtaaOp3MxCfNS0aPfyIWmKNVeBc1mpWPSx0TEmsr0VDHoO25VzY+5KRF6s+1qj
Gl8e65RiWKXeNBXbaLYq3hxaQPtime9h2Nz7ExCfVZ+fAK/qHHd3KrrrktQHC/t4a+UP5f0oe/4w
ex2f58kwgJOMRfd7r/ikeQAGkGS9R+Gfn2ARxk/rJlTqsx3Nk9Xr9zjv/Ujkx8PG9vw+qPZaQGsW
HoVvThEJX//MP9uedZJhpfy4BG0WFw1cSJAvJBaBo4T/lmy8K92Hx5Rxf/NHOGFKhmTQwSZqCkgd
cLKfM4x6b3xN62beJm8+ZgYpB7DEyqEiYjWvLBZxOsPD1ETkEw9qp++mkDvuLbeemIvn+H+ckUvB
hnhbW2OM7WTFLpVY3dp5QNMRF7FGsLPgiOy47X6nTRziiBnI9jk6wG5erBQbR3h7AN64IdXlIrNz
jC8fVdt36xwg1HLinZrK19tJv7+7eSWhatdR040wMn0gWXVVipgV1OQR+OJHfpAXX9hvjkEh7kEz
91wKBo0c+mtj/9r18Lk+64VmTwF/Y5tDericvylJHF1//okTN+8dnS17S2F7l40gWtPJN9cNmp1Z
34+7CLTIMpZNXUy5LQbPiKAngMy2gELh6flZk5pCJ0LW6F/qmpLNx5QiVUE6PcA+V52V4810dyd3
N8EHkGmz7MAyPhyXwhM2m+BXdyG5Pkc1c81BLc6YXlmV+r0EZsNEltsxxNEqikL7cBnROHSkoipG
IawG/JRKQIGQ3V4w2yeKXLew5SZkwGiIReLQDwgrkCRbFeTobIvs9hhJCC5EGBvBRgLdbFyf/qmv
hvnSRDUee4UKXistWp25btKSkdPllYH8e41A0s+jBNRUMO24Ej55May0Mpqz3pMdem8p1utAOKu9
Szek0jRykxpaD/Zb4/Xli/0ajpzwlAEtQT0rVkMDBr68fnccfdEjdFSHsdTyOzcOyyKTcu2Tnj2L
t21sI2FRfAEw+Yff2ss0DUd6nOuFEfrkFjuA6yg//EjohV0ECACLyXoTpiXq1gkQ0g5uLhB9j3wZ
RWXeNzSvF/h+9Qw8YteDECl1nBrJQJbyS1PWTvWfCKT4gWE6re1AADGjdOl/xPxJkT+FVkY14hFU
ahgaB2NdupGK4fVn9dBLs8kt0qFkaeOUgZtZgeFE1pGncM8RhjOAWAqP2hQvFsUZ9jUFK9tc+r9S
SCrz4OFepR4KrtSqdPIIIk3UcvfOX45iiCDMancJCWxEkISavqBkjpmyTN0jddnb1Bb43zLriwQX
ZBllsDSCwH2rIXPm/6VTUuHOb605ZRM7DHXilKBLwsYQBfdT9FWnr1Njx1RMV7QnuD25duGK14j5
+lYSaAXR6a/qZPuo80NczLHOnvyijxuqGxYZtIPESlOosILRgz0LswsHFTQePd+FuWF9Q3F5sHMJ
V07YSEmXbvoHYNAyO5ZiyHepvXa73Ahq+Pmey2i8Z+zREJlleKzOrsd/0QjYCkrsAvdOMiOyKpoy
xtrXoZD4D6IudS/zo4bn1T4iloZ+xVudVK0xLqftu3ig/UcpkYWJUQFcCAHWTIjoDr6HElLkUChu
RlAVAHmElsa+7NHC9VZYoXgMDBlDommPU26axovU5HPULU5gqdKixnbh+gwrNj8CuG08E72HkATY
TVHZO7r1mlfin05xrs4CD+bTlDGd44Zu9C0najShLrOipXIkAxZOMYmuWw9gU5e2PtT9Xq7nC4MM
+5jJ4lmxNzgRn59RUAKxZRqBaoyXQeKBwegLE5dtdLWoDNK1kRA/CuPIbiZuwV7+oFTbBsjl0dpx
KsgI4Qg9X8t/Sc9F2EpeDjKkG7UhYaix+zee+OEyHE/CFH5pilTZgEVyq2T2d7qd1TlpAIcps4b6
LDdraT2rFTw86UfEzIAjzXD6Bib3ZZ39mUSNXNCVfst81FwkCvrhNQf5goWQffiFi6We6G+sv5sL
fKgY1NwjG7QzHIKb5FdO65dxKYzTJb6VJ7yWZrOO33RNC5NdOVe83o4wdB3Hhwtd9yogIWpuvyYf
FztCK/kH1X5PbslN0MUVj2BRm9VrQe1thK1/QzBifphOHmyUiuL7Eyq3S0TKX3t99zfOjwDkfnMY
CmqIkERkJPKTQVomAYmSZtVPh4CdyjUkVp0jW7zosAQXrRN0OIzPWSeRLLvKCeWNDIUqiVcQdgK0
EdsHTDL5+pk8ofV6OkSUWZTj8xdvfT3ldEBDHzno4ij28yIFw6DpK6Bw9iRHfamlPykuT+y74ezC
KYVk6Rnb5Kbmus51tEW5KCzNx3iULXgXjBYiOoZpKbeo7Nw6abR6l4rwazp3uUwXSZavqYnc1sv4
zsyNQIeg/2k4x2FkLjS1TGmy5+UpSGC7DQ5dTAfo1ZvAhPiJ7xDkO1JkZYuUFWiFDbK7bzAiTzy9
mqgg0M1IqBPNmxG9086gIh3xWCX1yH6nArwjPDYM5+GttfJpypbTOtG1NkTj0lEnbgET/l9coWg2
p6ydP8duez4kUnK9NBpp+GHM4ihY2WHsCEDKTIB4a024sDh+1lOr/afQNw4/VfKVdjbwLl6isdzW
ojEYWJDF1S+5RL75in9xetP/troMHjjf7voC8cvwXgCBJotDUNfjkddzpC9AA1MPZeVOvhlNz3Dn
zHUfDP+ZutU+NLEgU7cyIDavlrvhol6L0VsOEsq+uhQZJXwqMHfIexSHPSeLGHufG9k7TnQnzbN+
+u3X7abGuboKRXealDW22DSxSrqUB+RQ1oiPOgcT24PerOHSowCF96l8tv/vBe/zOMKvjf8ysiBt
k69mXwCmBc5TjJXwHlLPBASd5Rn14EQkrvwnWRGxar1sR7x2EY+wxpzNJoTrgbJJ/lZ0vtI+MXic
90trYF2zwsDgTbU/X/HWZ2w3lRM2QlUeimzoY46aNT91kGXao2soyzmXOwY2tYgRyuG2O/ZG+ciY
O9QEdDynYSgU1ZjLzKJhELCDATaNp/VCrbAAj2nTtdq6teXxx4BZA93tr4Ns+3wNuWrcZaeaHdJZ
2ZJRd3DCrOFZ7gLBkB3NwQLzMQkwclwiMby0ZFL8ZkXlakxzKt49eg+QaFEIo+75BcZxQ0lUU8Tp
PwkOzLp+hGFPcGrhTAAqy74FxeCwv50qJr8i5C/BMXHw9pzmJSOTNf9WwjigDaHZnz6w4U8c3vRV
3Jxo4r44ZqabkG5h1KLKF2/PZh+tn31IsWYZ9weHHFZnRnutUHNYvOTxiyKJ7Ov6hsOJ0KYyW/5J
uFKTz4IHR4W8K1YNMA+PCV0LyUE4ZE5yPTYVs4GuAs7EM+Rf6uqhZ+Z42Alh4xVbDEmzNx0STkrr
iC8EGN14qPE/3/u3mE8/ywVxek2HfEAHtm310W9XiD7Dv1JLQWAPfPeZ8At1BuWJEMzj8Y2LZTme
T/AXEVmaMR33fXiuAxbtmoe4bT9hhA/ksKg80/eA6rSgvr/jj7uTpplp0zwHrYOnNQTwLDaCXLi7
z9lpYgE7pYfr3qW3WrJe4BxWEdrKzwWOtBuU4ucwhQiaKuBFUqIt4Cdrfc/xvq5yhO7oUfKQ/KT+
nd6f7u8zpO/9FVFGeJkMsKho2RNzGna6M6YufcuXlwDYJ+RVqyb0OOo0GpZM80dDU+Yd7vuWQ21a
FuV+RQFiVNDW6MHYMXTWhka/k6jTkj82IL2SJhWYYF+N5xciQLYoQ9vK4XhjBpymUEGicFwtJb2c
2jvHh/DjnnI8En36G7Od/uFwZ6rk6gWjG25d5VA46SHnUkOSpynlCdZPg3KTgJQ4P2F/zhD+kbnc
UjYte/2wNZN/RrCfzxTDgKuyo76SBlQd744EHA0REy4t3LDL47FGT7C0hufC6187BPd1Mx3rldiR
2VZOg9UPcFYGo+YSK0vRGFcQeGBkomD2LZGh0wqlzjIA/F0/GVzyFBCEoYcguabZrI58L1bCaCLp
7DW9dKSJlgjx8vxh64jO+qbFqpasIiSEECiRxqctiJav+BK4a0A01dpkikNcQVXnM4/U63t04FI/
pooiO5Qc400Gx32oQLCgj2CkbX7qo9C5wd3ImnF5ZMqc534uZz9HgiZa8or/C9Jm6P8hGzyEpeH5
6yYKVqmaYMXpm3+jLHRLn3bV3ZdE4TDN8GsHSV9/BFy/6lEzIXJgWiUiJxGRkYrMobxHOcIPTZ+I
ZVSxyLuIVbkmchCpNvvhz1GgsZHpDZuO585DxUzmzM6oojhSHPWcmozdil983JAmTAVLilSYBUNw
07bYy/ZoMCQzuMVJCUaKyVXWJXOsUFMxwjLNVH6XTFANsFbhhePUzSufw/Yw7WHw+la0O9d6RdUS
B3PIFVkgddUd1cKBAIAEwx/TJf2V4UgjaiYnwQGWAaWuA5iMELSP6+y1ZGYadhYhTWpZmmWJe0Fq
aZ2g0uouS2Tb1woFDmnsZplffiKQGyV8ATG4zzYdbAmjD/+sk6KtD6oxChJIi+PUg1EAKUbRZInP
ZdyA68XmdmsobRX0hhvejOsYEIQkLE6MEWoNMT7b95hu/v7egSSQiZp/LqQAlCghm/kR48ET2tCD
EJZ+gHyjs7/LhOySGp1BMVG4qPy0ly34tV9Dxyf0ZZp5O3XEOIV9gTbPy8LJkREBCanfgDO7loZg
WQp9hNBQ8J0Ed8HodN/KoUjqeKGkcdRsy9aWfZHo6/iVlHbuOYGrNBeisSo1+4Ny6V+4lsiCcLeT
0m5R+xU8nf+2GWK81exvn54ccvS0EeybOUcazQx3HO/X8BDLURbfNRUyoxloK6yonllQErnoN9wJ
YX/+zQDrS+1IYhMXhSUHCk8uhms6ExXIQkI+3FtGjZP838i5WFfhKrpHPNRXTJWdYg6aqv9bxmYX
yZ2IiAMmxmwX/zuRDiSm3HjD8hBH5jIst07Fl7ch4EL2C6tWpy/jTfR2oQ+AFpOFGWiCdw3R0P3m
dvQ1RPhndFMhHy/fIU+NuNH/jyJIdwJ4/IBpXHl9sUCXnilVsku8rvnF1uW1QzVyHrWp6Nkn9jBa
qpDAFsBmjTLoIfcEMkW4VaPFvVfkLpad1z3Zzx7q9Uh9GzJM0HwMuVL0wJZuO7DI16GXVmRYRQar
xObwG1tL3FsTbae/olUgu/EqSiIP5H2yi/O1/RqqO9QhJrpizM4Rvl+44J2hPtVN6uOU5NVbc51+
YLP3HeKotfrpiA8+8qCrD2uqP0SdertT0xw0Uz5+2/A1nODKVp7mQT80ouehr7L0OqEMGkN3143O
auySXoQ6IJpUpYLcCg8JRF48SCr7uPvdlIc/vtN1g6lmdPsVbIsa+ke6b/nVvbO3ZwYzsi2glMIg
ENVc0RhwPHnj+9tW19EEyP8O5I4uHJft06nCatTqMvzOVBlGxugYfjollhkO3huuDRzIZvqmCD3I
lIwWGenplPI9YKfBX7qNRDx818WAweAjLbjyNo0GlBv/N/xh9tb6uZ7w7+du2GM1KMBvqV+5cYO3
7VO3OP+ofwiXOHFOZcoX72p0qgbuaaMhZMg3tkeWzvv1cKoZvvlfvH+rWSGjbqgN8QHOQdHNvAOB
AvrY13Wnkuc6RSgvs+ezw2ZtqbmV8gfmGmz5cGAqPSve3BKWaGXlurkEAsWO15+aGRsHB8UM83kL
7NsW4PIIHIYjQKi1HeQuhMCYf0x3sP59mAeIFjM3DWtdM/jzeRzkRpUdr6goFy3SF29pzsEINLUR
jL2fF3cNLOEbyAq7+WCmZjcy6KsA+RPS8pX/WSyy2aYJfM31XWwiaKSb9igI8KJ/Tw+PWVmhFSIz
+NufSrJZZbucfgkpcAd7+IFrEDPhrCZmAkYzJwMkdg10zFblReDRwxD8q8jjJ2bQO2Uj1l7ctlQ8
ektlDB7xnL4vWXgKUPOTB4a/q+/0eh4nuUzA6qJL8Yn8ias1h3+jeUF74UNXr2t/YOb7rRByB6na
yyCpJ1Szu0wZC7wZKfrcYyvFW60nPuOrnn/XrgQIno5QlVxbvGbu2nIdhbavVPZpBquUkzmfvJ0p
MfMgBvVussmaznSSGGmOT/BOD5CMNsSDiv0g4RfOeVM0DlQQIhKwEwpD2O1FW7wXR2yl6AhhyK+R
yFMHJJjKaIZwjhIsW/lGeCotV+ruC5y1gXhVdb12mDSGR1JUEOj6jE2QCairngFRXT5c0l6INemE
rFsY9QgBl+8amGwyvNQm2A9aobTFhdQmbfAOTGpP6zKbMr6kC0jSpB+TFIMhtPwp7IkXPNIqkEoq
/3/NHY8VtBY8n9JSXC/1ESzqNtYjwlckCTIZnr0cNfD9M8NAjmL31WBCcVaJe4lzzZHtqmWBc9iY
gbcE+LB5kQohOZV3Cj8cbm2lyaAP2F/GQUKdJmW9VBPTP8S4bV2hZ7yIipc1HykTo+Dk40b1Lba1
fcDP31v9nGOjBIHgxmDpRibn0QYVhMVU/qpmNyXAm4yVm96seErPopFi0s66XSWf3Og8+Er0H5dc
HUc1gZbYGoGUp3uunr2XsrWwv5EiYybl7Yd05O9mIb/zqItHGSLI3VUO0DEBAak347PLB0e7znd1
CJ4+iPNY52dCBj9MBGgb2T73cgsi/YyaAW3Levlk7GyjHJsITIam0HroC/mCcNWLUfa1bBmtABJl
1LFjxuMVoVbnB8Yoi1fDD7ONUBB5de61+bQiv7+BhBesRJQ6Wgi0av3MNjZKyIIJL+pRfgAUXyJN
SrhsNXlEPXSDlqWrZVxc3R5Crqszt+Rj+fsLTtC4RUrG4yGLCLTBhGi9VxNm86FJYtdwkCjN3qo6
4eq0XmQbby395csWy+Hd5FE672aG2Rt1jX0BBotVLN/vIMP/yugC4MLzWMGycP5G59Hb+QvNolkE
MvqDv1eqUWX42mMgkH3Wj+NjQZ2A8wX6kKRodDeyNXYP+C1eu3BSVJFjCiC4ouoUjMj1+/NE1LV8
1+S1wYeXze90nsf0GjkaQc0LvUHCrtLyIMeN8ELDKLWQRGmYlcX6OtomxK1bA/CCMtXgLZyzh5y3
sDmkF7p2x0KtKxLhBdnNJ7VfOHO2maYe4+4ZNJRXWbiTaEXzvcYqLGQgOkjgqJ8gQUKCQglggEds
U1PF3I6N4WCsWrL7km2fyfgYXajlMQWBMagL2Y3Gx3uDtvgF8Zr2xHNLScHs/o2bRcltyDtWVp+r
PFh//NlriXlqHPoddfbwc5Jeadif5nhd0n85LP5Keeiu68viGDExS9MSey+CJ1C3otfHGbtJXYzM
kuccwXbbrIVvN6S6RqdFfNsVUYfBxIr8VoqnpP8zoY6B38apj1qlu79aTigT0QmFMSlPnZQ5au3J
NmTzrHWMOxstKCJJbxFmTU4KE1i5KTAHgAAQlGvGKr2TXWWYlBwlkQ6eItg3x/CgPxvU2RInwFu8
4V97d29bZBNLepsHfqTYmANeaE1fbgsLNtaiIpMVerSObyHc7xYISCfdJ+su6Ze0/ckL5KcEPjI+
lU/EM19nCbYhjUOd7Z+G/TxjYjmSpYhHZW4eG6zVt9m1bE3Ywp7bSkSbJ2LfGrtAZGnUGrWXZyOt
fDGKCRhVqjxkjOyp43zCtLttfDfn3GrZmsM505ELg8l5UMVy57bvuf+eUCql+FcSGVIlYxoLeIas
asiSY/KMz4TNJ6W5v6sCOHGpeIAwHxPYh7LSeA9UD6CxoCVDOxtVuf4vOLCAOXbmUP58SywtYRRs
TdwJ4HPxcHMSgVK2T+3jGNgeUTDYzeIL0IAIT4fsS0ccCYJrEazpOsW9LxC36z6G6LH/CCKliYss
f7Wb/8zty7hBzHT8IJfx5hD+fCRj1dkmvAQVfyp/JFGeYxr1NOGVKjXk7QJYSAX8P0kp/qvt2y23
139gEPD4U1RsbKwmbzDUOkWp3lX+hJtSWEiF3MuFKyLD9WrO8iZjXApAGKb6kpzrSu6goAqBbNgo
FTKIz2NCJcjP1gUQ2xvTDLrixu50CYVpVlFLq5pYtC6ifpGac+dShJ9sVbiOyguYFITVMtXbjG43
IWb6dIlT1n/KKXM9do4fHJqO8AQExedaUkL2TILHrC2/jFLSXRQP2GZAtgOFyQ156evGw07U7MCC
rj4Kw371D5nL/4rJclwbiWGHaj+3RMIOBogDxHZsBLnLcehKTdBzdYNzgpXzKm+dATrHIc+GmkKK
zW6vNi2iOb1aixNPSeuH/LOwprzWslTJxlUY1ku4PgCwD8HWktJ5oODh61PRYmJBa9GgyBciHejH
DDS7Q60jZlXxJtBD/D9CZ2NVfBvK0veOB8JutwWjc7Id9Gzutul+is5UEhvGQXij3OsGA4o3X/gb
oOPwCTItN120dT5r2Bbc1bj0aoXErofXiMY6SW6YE5hNGlLKHrB1nrH230UOarbHLpAk7NkBfQ7v
smOoIiGpQ/5lWJTnVyFQ85IC8OLFdBVPyYNuwhAlfeAWS8Zg82cXUuI5H6hyrg6jkCkhZlL3+eWI
uylk3uPP4//yJm6p74Odms+Avv/JQ+GcwctWZNhaDWxKLGqbDYhQypqEszp1hhKnVbLysGWlVGCY
ppIS7/k9cPCxMOB+OhlYxOyldQkgKhcF8sxvhKziJINymSqvNcUabOtyvdTSFlVr2JlPDAfLJSAL
WFOmL19nzHrvJVgkyrvACNgAHH7PzKOUIBqKC6xWHHb4sMjzRG164NnSJkvGMKPIOGxLYjmJmc2O
fdqgutBBcJ38D6szNyR6HTm0l/7JtJyRh8rOO4QjNKZUjVAil4zXOycNA6GJh/R5WmJK6Zk8/xK9
+dthpX0bN43vMPNBo1RrREuo3e09aOH/hY0J1yhemgNSqhc78xRQk3JLLJX1kyL4ygnU2rQZ4/qI
CG9O9x6qgPZ3iuGqDS+4ysMW2c3SVA2JSCyvJUKKUP0RP6mIbaeLoQQrju/HUilcedjlJGkwM6JL
bqIM1XwJh0QSCdyNlKki+s9kdd0SClxwKm7AI+JlGRRH8FCTeE2MUYSDzg3d/Awcp8+fCuCU/kok
6omBmRdAetGuBPg8oBnW8o7pENOAILwOxqW0C7r1pDwk0Iqq7JbgC+uUZGP4bHd8ycdIRqjSWXkX
uyn2irh03lJQV41Bn5RuaYsadHJYRL4YfCsMEkqyFvruUQ2vm/cKtlLx35muqgfUtvovDr8KdK4D
XHHAhCPGRsyb7RBIJMllu/CYZcotcpwYzapoSzLHeFOmbMMciCZmWznePnJiM5T6PNMxCzkfXHQ5
xawQffSREdJkjSYQAA+4g7Ve8n+/yD49R9snu4jTyz4EMVCKfu6/rCyj+rXCFIq/VOItAiuzJCOW
3dxIC+dvwcPxRYGWXKjcAep1VJgOISmQEmLvLEtIvBZCH/pPfMVjeWo+ukYzsKzMLlT5wtYcYAdx
JWj9Pue9t7uGPlKyhVZVZARLAYLXAgR8XH29e1zK9nRMOHwC/0G08g3DY1wJqpshX5omCIXtBioa
qsFXaYAM5UlFR4suo1IAquqOpiI9RY82nfpOjHpES7cvBVSPA9fMUZokwEKcO7Xt5M+Sl8ErEkiG
TJ4SvPUv3zKh6gcVgFjSu6P+kha3P6fSqZ9U9XiuiN5uGkc1bQrK1c4Po4emDJGn1P5yFp0Qunfh
KpbryJ8prxVZ/xiVQP6YO+ZPzqmONLJgdQCV19b6eRWLaxNmWChjgwCp/5kXliT8cQKyOARznQRN
7LPPtyw/8w6QxtoQ40lX/dpSO2BK5Rrd7IPD8dEV16KYM9+bQUO4M9DlOIx6vOVpxTOAOfSUpMnJ
P2gAfzIcZRG2aK9JGz/avWrYPWHxPL8mPYMbIKh4BtQqrYMFK1++0HfZ2NSkoZ3DCXeDEM4d+zDm
pp2yXFf4u/j2yKF3h5YKyW9kaJ2bbCCj9Esip1S3LS69bNy2X/86ZOX7smUQA5OAMwzK41+bzpu/
oc9koaVE+3hUv76Df1x3Eg294jvU4u8ENSPPrvT2bKoQ0xjO97UiMEke00FPISMlpT7FJ9hwmaEv
cdB0xfZktgWDoUoCeYQPwtUGbXqk0Ev6/DSdKgpkVXEUPs8kDKyciRrZl0t6CyKGMGBzbpGwYnju
hchM5tK9Vrnfuy9SqsOSLBCAcr3cNosjmA9g2Y/LRy/LRzsItz9B7RFFRmonvlsuCPc+GcBTWpUe
wHlGXF3Nl+Go99q2tvwYhxeDcAES4gbUt3Awu7lwCDpYZu+DRyMFcNgzumX+l00CbBLuYjV9lc70
IkR3r1fBKguM1yBrO3Z5HzPDEqhfplhZH7tJqzP5/V9ZgX4JYMf0NgzSO+R0U+lxFjhSGXo/Xq+3
xkWHZziGBu4iBSe01v78v8IiwOeROcEmhW6BPA5jI9djfZWyTUBAOYd5A0vm60L5Bfr9lIGBfSQu
A7zE0NZcWQx5Ce3GFIQ9FKQtOrvE6JEqIAIkW4nw6Idut9StXQp68PZ8c7sMo3U336PkAqlr1G9U
2yd2NYkhpLUeM9RP4l4trmpg1pGs3vVaRe+hU8Tiute6kB7Y5gulLNY/uaROBj4kD5jjMDQb2QA2
ayLDWTXuZs3zV+qShe9O/ppzqsfWP7lwI+KQxXm7e4yjOwU0owdJFkzysWqXSay2eJ8zWar5sxc3
gKVnkeZHvOB30AEduO7sU+qRi0HqJfKI8r14LkvM5mmTN1Oty3wguHMm4VWT++EX1Z9PlZBNhXzZ
E5F/kc+tegW2N3PFHF5JQqCDhDoEwqFyIxlv2TkxKkksHAKSo99I2E6RZ6yUV80ADJ3Hcrvmp/uI
uLGdrFjMAVyZCvlzPJJXM/dx1R2WYvtxJ5+lB8W9oPptoFEMtE+RfE2h2/K0qMrcVCRMj3AOZo6U
zqa9Un2Xjm/Ou2kyIZj4jINVXQbeDvG9Ko5BfudmXQLO7M1bv424I+WQ/2ZjDs5+Ht4xZv5w2Tl2
dHY9og9XZFMQ4seLeU6YPalYeCBRCuyU2KIeUNnXOvju6WTbEZt45sE3u3EXOVn9Mn4TsZw3JYiW
e5BYIGOzOIa2EC87y3LKQcs57YYtlovSnKTyQiS6ykUo34DvE5/Te37y/WAbLsD/2tlp4O8xgAPO
20yHshTks0lrqgdbyXI8klULqfjZ4TTH0gaxGgzhZEiJgNras32UdJinIZe5s/LKVjeWVGHeQPQa
KlBh5H051BhCQXIU0S4MI9+rq1RzDxP8nLWwDtDW8PfTrno4FpNqOSO80rs+9n2ScC450WLoPtox
jogm9q4v2DGRxIyBGEWKENcdMuFm55E9+VWpeO0NdRNIyMJ/aJf1tbVGu1gSuB+SzKfn48Qq1WKo
BebuAKQM0Fgmw+0Nk40hkRe7JVLiMm0BI0uXINXfUX6OQXTZ4I33y0Hhv6ABRH2hgs9OS1DpZao+
sFQGZsS6EJS518s105Gh/K+KuLTY2yIVbPeLx3Te6jI1qd0K4+pEVVFNrv1+H3g+Iat1dYvN0QWF
dNSySuBrUuypP1pnZ7RblQyigIM7GYTPiaVGR5iN/udVqGuqyKszqJLw7GDZIOlLKYf6L2iBjeJT
Rcm9nqKJ7qlbdkiZNlcq/rn5ixzUdiu7vSKGFTKOqlKj74kgcaofc8N9ANoHpNAVuiRQB77kMcVq
XtkqxbDkBKzPH7kUxUJtn3/zP8CXEMv9Opa34ptK1MMyzybwAdjJECK5aiGL7pYlTE9HlH8/Ng3i
/SbNiZb4rr1NIZXQMxgDt22Byye24W6OWwxsS41GWEK+tl3+JrfvGYZbfmYZ53vURBgMEiYrgfy3
oeBsMXP4PhSBWlAxcfvM4m6HT1joCwiw/ETwBTYiWkWtBYfwQhmpgXx6E+NMh7bvLbTp+ZHpirEz
pu4Kl2+iKDrzRAWtjcrpLGSelGGJnNpuFNlD4JSfRio5LFyrRv9VTgfnbQs36HMObLN9vqKRqBWv
C1h/apZjufL7Kmuo3aFACNw1Fmht97EvsJOFqkgxxN2KPXpAxip/V55CC8qU3dDZOIFNS0aRnA4B
TkVp1OFuCZPoMGrFAm/8Jbk9LqpQK/0r7W//vf0OTbhCf/9bWt64u8qbAQug7HG7GDvu81PdEdXk
N4BHC6edspdoTW75N/amqu+mCu6SHSy1dJyDek+CRRX4qVqji9eKWMlN+fEI9GAedOYcf3egxnQo
x1OeDFdoTpFqsQFsQB84yLdkMHsidrbeygMU5x1vKr1JFPRnbzCnIEChKqMMesTft8Z4iCND1CTJ
iUak+F/lIUbE0aotrWvnx2VyzgSj8S6PiFF3AZcrugE8KOVE3tf0iSfGakzSw36+mJNtYT6Yc2uM
iiMhlUd3KunnTHYJ2fOVZFdXL9n1+ztGm/ncBcew0jSg1mEna7JQXGAmWokfnbelpTZPZ+dyOlup
ykQP5UT4NSAq56h6OKzyFP+2ogkQNTTiV6qJA0krPvyzCgZXBg2+fpiLXKiZkKnurpgKnUn7gMEo
ugggSpCNBgjyAStKsRCDu2OVsUariVDLTAcM7xHkLGydPw4QtDHOf1paLGZr9URy/Gr8DzTBJdQX
7+nj5hkFh2kHsfpVpxnrRaz5cWq5gn4lGCh32p2IDVIT9O3Ba8cyz4nSfSjNyyjz2nBOIy6wq4sd
WbCgZyCbJc9A+hFzxIDJ/kJ5dZe21NFTshWa74iNMHDwrMkBXiUkr6QaoHbwv9LP+n6429x3Vb/M
bwd+cFtipBgIZ/34r6DKNIO9s55/q/+29awadO4Hd73RKyKFtfbYnYZO8yhB3DPx+LnNsiI1goRW
l0902AURPfCJBfCJsW/0NBQNkHMlcbq7GwjL9d9UsXpCcd1cTKfTeZViLqyaD9Pxl1pt9y7oiNvm
P5BmOuUdSQecV3q1XLZ/Wg1+roOt423p/6oy3XfFqy1L34J3mpfUFNXeSz6d8/kEvmLbdF96OG+y
uTaAfFsZ2XUehd9UslFeTHvEtwV+msMzbJNuNcyYOrdb6Gswnx3KpXEDZ6neFY2TKH0S+9kPQjF7
QJLtFTQNS9jbNVs1ceIpZ9RnNWJ2vaiaiJtjzUp9cg5vOqeYaSuoBeYqfY6KYWspgPCtDDF3cE57
hW2tQKo34PZVD7MQUnluy5+KS+EsSi9h/St+/Raq4NTCwmtLdPFoo/wXAL6hpqOylGT6vIq2dgum
Hx6Sy8XrVhdw08lRMlKNiqM0ZyCDc0fWoWigxPkPYs9O0QcFHToG1PDTa5H1J90z8ClHQfnvNx1r
EvH4Utgxb+7QbDHQgCdY/eiF9VVPM8x2eK0YonB99UepbKUkxytW2SnLoDM1cZZ7W78Bo/Ur/u0P
9A2vFC4fIM2EJEX3+rQcIlG0PuE7JL43MT4SXNgcvQraMhLXuL/tc77J7DvUOEVxpg/yvii1pO7/
vqOeKUKVn9Img42ciZ6vq38ZYZeFuCG5zchvaFuCRBiZEZ/S9jx37J0p5HQAxtvNCNK1DE+3MhbH
rSeJW2mb+W9FWet4ZW+1HCX841UBWefglfj7zimNKPGigGeBNw1ZzvK1CFjOHQoF1EwBJyjCK1uG
gNzZDVxAdqXE8dx3IBUzjfE+vBAdFb2Zm0zFz1+pt0tY9VwHkwVU/3DmStDgC3URD7XEJM6OVCYr
rAjjJZeRwmFMGX1Di58Ccu811ShecScDQPQZKyBjn4DUvPYZlr5FFURs3+5Oo6BicsF+dh5j/8CV
esfPxQZJg7SwOt1vVrRwJfDTGX+hafuyNQTIYuLWO5gIZBnRZndeVW743sWVLhgsbUQn9w4vQPYS
esfx5QLY9KUasF+JcABN94muHiblKtV6b/VFgLJVxrvUOE472xH8etTf4n3DtDNhnI5tnVUn58ws
cZRq0mxFCG6bOTujw4dslwY8aJ+Tq4IoSso1UFT4bceAvYODwB5P7mHt2eYdxSZvWIMeWJHT2B1U
suMsiwFHw3eIOn4IvtKfrAbA+q92ePelPAcul3lXWj83UAILWWOdQu885zTBQS5JriBYu0kZ3IsP
BaQ26IvAW53V6EBGP86GvegE3H1WU7lpMZBCRP7hQVn1C74rMusG6YCC3/3NLhKKPHLUgn2DmFGr
7Ctd7X/mV3VHhtT4sSpe+YKODpEzRk5nyLlL3Fb+RUcmWsjP+mhZ3+uXOEqAMr5Abie0BM10f5hT
ZGddzXJzBZtVyL9Ofp7JVw6vUrptsuaGdf+3NVM68KqWKeLztvDKXbhEfKcq6qfqbKIxgAsOd0PC
RA1p5sODG1ODGAGRO/SI5XLB3iJaERqRJD6/DpUGMDWiX7++Nn4ywsqvT+C5xf74ZpaTdIP90S8V
YgUMeER1Fp/cQFpWm1EHTesSZWYoPh5P5LIpJaRpDecGD0XW3Z9tJ5m2x3rmF3I/tts07FnuRItj
UHu4n6O+ggI86IvRu3OGJ2jlp2y/Uay5ZfHOCpZz1EYZZFefPC9byG8F9wBfJNyRCF29yI5tgUs+
kdRuC3oB24FpIJWe4enTRTfjcFPXk4QVD1+aB+oVMOiIB/na4Uuyaq8hrJI8VJJ2urTcoWiKoXda
V1LfNehSfGxnHmXsV5l1HWpDlWc370c2Ye97wtrMtQUT4Q6N4MghzYJO3B1hhEK8fttWM5sieq9G
xuD7q+uKuhVvyAGENk8jC0pUkrSOegXn24uzHfymsTWmoYi4tgtWjhLczz1i4OTSYzAwU6eNObs2
PZtRzdcvU1ScSuFW4UhPP8i7S+GpPJOLg2ylgfLtBUJ9dTt93SuumtQSphv+fbfBqsL57FtnO4zZ
Ij7tR85q1hM0dTexJIXUNp8S6uTH7AuYvHWny2TJtoaa5zpIwtWJbaqfRPqHFYx5/pCDmRCuiaa/
hrUYEjhdgGEgaiQGINnvDp43m8ACvsM6hxNhLDv+Jdya0PKv4lh3H7ZrDcqntJArzamoPXEV7xe/
sUC22axk53kFvkrX2jNzEeFwXkznErEqIoLI3hll7YTwMpbOnpwvqNRU2i+K5UNbpVIofSay9+M0
MQx34YdFo3lD0iuj+KPfb6kpXvdqYg7YaWnjshuc+PSHEemosfY2rBx/+KLI2xugzmuJJDPj6YRW
2CJM+6cv5v0OEd9eM4VjuRFERm25cFEKAucxfqEEtTqURI+y7JOezNpMANkz+F2TjxoNz7sh5qP9
xrOFhS8xutB5bq9SzrPICqeonPpc406NHij0f/1JNDAjUI9jqRV0Nvh6sVJg8SVytzRw5jTun7uf
iLLwB8JrtGNdAfLCKkXGlGLOD+baMVD6Q9pQ4PHZWFhcTdVvPZKLp5oxremw+jRnl5Ie1/cp1S8R
d4UKo7H8Ul/nMOYWEqYEnbBVqHN+T/Lju+h1feAQ9fsYAX6e7H2KI0rz4oaTR3UhqruFrhXqmzpc
vFauL9fyJ757czyVGf0XPOuJzTteTNZy949QAMVyjTDXLdqYeUTpiD13/6Oc8tiVt+JzS1WkqXKc
epN89UXIJsZBxAm54YUu0NxRukKamG6IpO7bM0XV8z75EugQKL5O8/JMLV8cZ9GzjoOr6ilMlYAa
MNxAJhuTtcT3zVAmf00wOQRNfXjPesCdQIJ2mi+HHtsrC1wFMP6+9FNj1vgmuIjBgvJePzDr1DkS
fak9DgrAyHCFOa3cR5nHUTStnnxuuiDlmUx08Etzqy/pSvi8YkSI7GW6Dyi80PHX4Eyb41GT03YD
MKIGJHhaXgn3Lg8IPwPx2hccj4ll0Ky7Fd5NMv4vQvSN3v/Pe2yySyBbL+qAfzQmty8zbyoFhqkB
/E1BZMiC6cRoIVfB3mTFBAkqcYcUwSA4F9nJ0x1wfHsavuHlrdf/s7/tPAhsmCIMFCO3vWsHRITY
d8zKqJ4R61WEscsgGbQSqN9vy9pTLAssaaS8NwPb0Jq6CyHqkvc6b4TytZ0g3wL9fZ7sTtiYTkcD
CKeV0eHSasf9R4A8xV9JRmf0b0I5LCLL6ikz8xAHySmq8Ky5cu/3SZhXSZRXIhJ4PNdw+IEJAOUv
fzP1R9SaoUjfu5vht1q97GHTttWiqHO2oJRLPTEJUYj2dgaxu0bk76N+T5mu/A/h2j2mBb1oHIit
4948FKHbIbQ7VRw+tSmYrp0d9ci3335GKTLB79DIsFfcT8mJVhLMfXXFKGaMU0sY9zx4KrSfa+bg
NpHhUcPjpwrFkw5zFNxilFXc/DzBTIuHNVnLHwP7vDuvKix6iX7MM2nnY3VGoF6+GxRMGUSd3BfZ
OqyPkhh4V6gxNKnghqqdcOr6XYwyaW9xx34AHxYJj1W0njBdDXS3t2z52NMOHnRj5MlSUje1YZvt
hXsvpWuZ6F3IMB1taY/IVkTS6GH799dj+iT4MpKQF8keDopfA2OTCuGH5pNypoFpzdN6PQo+meZ5
duF0kTeZdADVWTZVLRmi5+CWPO1gVuj7+EL6X1PN9DFUD+1qn9q8a7L0HGAtbP9wP/avLuuRDH4G
tbdv2I09nKw7nlPTt8hZSmhC/hQS8fvGTIn6h7FjTY9Gd1hF9jHNIhGbya6HMDxGGaS9Y54Ta4LJ
MY2+uADuLSUhTBjpqEJGfr0ViVxM4armyThr2nylQaDLo5FuipKgcG1Sxsaa1NKnguEjElIedmyN
NuvnYtuwHe8iCexLX4+COIX6XJKQ/Lh52MFqPWB/PUPvdh1j6ibXrbBkZ8Z/9DXP5rOXm0P4pwHn
FHoAZRcJyruSiHC0iDPShHacGEBoTtV+JEyDwrUeQor155jK+sKRC9yHcD5/9CGUnWQA19+zYc+e
R7Vfoqw4Dp9RWg0vib7NGp37uQtw75igF69/jVRBoSHN/Kx8Fc0ie4BodQeZ69epluOYgrGkwigO
jUnvm/qzBTZUXP3RagDqj2KIiyBfErlgrPCsnIvumNzpSbMuCVxlFFnLANtF0Bj1QRyfUjXhPxrV
myRkLptwSW3GWYRXExXsQ0GLNjiV8bdcPmJiPmn1MXxSe6M/wxNrLju/pBrVX5HzeRfjBGlOYkdj
NDtOTqek08jC5Ga1Jfut6aLM7yoYHDmNXC36KwGautBygy6U0yazHryfTGq8JB1wqLquPPwenp1R
RgQ+9pBQ9TcJDWuI1g626hm+vYwMUKsq0+jzb/8CRdjuiZyoUR+71ptu3irAY8/9J7ZRsEejW7Ae
iBJEk1De7/+q7eX4E8wiPga6C8/jFZNrVj8WsJj2BhXvCzVMiW9ANDmKODfpWNcXP0KOiPmp7hEH
u2WKXxnbFAep8iPo0jrU71RjuwN+wNKWXfKaYZgkhcEO51shfNOC9x8gugw2se8D9LgDT5u9wnbQ
T+4U88zPLXKzhsbJwzfd9CBkq3P5xKjGYlhu4B+ncVJ5PUzCAzit3eIW+oqdsBZ/ZcEKUbuJb8UW
yxjH76yeoPFddwi/RLY/WFQ3mU6CWU7El2HdbhxhNzU4pvF4Rw7QBytLGDFdU07glX9XLFU05rzU
8sVRmlbusB0s1ypOn2VdKGAfQ/wCgneXSnIAIhqErrRkm/BF/P2zCMQVap3D/O9z+Q2s6eWbjKl7
QD8oyIhtluWjX74tdrvcRM9D9VvOEAHOabFR8473UzuGvp2Zw5St3rGiUiwym68YC+N1D5s7X8J7
RXDe7NauhINbN/yFrcwnWqKxFqLx8jcf54hvisf+gKsNXdukswbu3ALDXOJcCEbxninDCAyCW0B8
ZAv/PTaW0ge0mY+ninZiZLuQcQUmMz2RHdWC4o5ptPrTZDhe8LC9w40RX1dsp8nglsaeARY7hd4M
8lzPA/5H9giFZQD4OlhiIRt7iGvd213kFnJ2rtRv6YnugH1TcNrORvh9wowE4Vt+PwK1TuJnM9VU
z9zoQ/oP+YbKZ+4LNflypCQ5du4hBIOPAVWEVHVXC3JMg4ipvHGHG5RNn5v19ta9q77THZ/J0DPf
eDXs9lepqRy9nAjr4NolA2eSq5wptGrBHabLk18CSTCBn6EIysGaq+Z+y8ahB2O4CbUqHqtoJErw
y0H/fuHjRpfROl7uLL2O//Gs3f0vccK1LO4QxphVcCCeUZy4IDd4TNfaSIy+7VSnyOIMVLKE2CFp
kky6GZJsm3PBHYykbiKpJOThstgZmKwpe+4WI0MZtr9+ZhVkrUzxCHwpjgAxk0p+ceLUaWkBZZyC
f7aBEA7cOLs0TKJ53XN23jl2EqqCDEyZr03wrr02p1xxolrp3Gl9gc7T4NBVJUNFMKbDpJC8PZX3
OinGRs4ggJ3lq48v6V27HCnquQIEqAEVdIEc5RxuygxxVZEEEDFwuR5MJaXX0UGwU4exaGneGjsQ
3b48oAgVguDT10zDfcXQi73RGst6qWkA/LTQuDWww6DfPMHGxSXrGNtfsFdr8e6Hq/iwviky8Dhb
gjD5tY8iSTEq0BJBSWI65RZdlC0vZpeq3DXkiqSWRzRQPGGvHnCxQ80cQPyYfxBypnH7FbIxyfX4
bedbCRYpW8qVMI0/SeOzjaWk8k2iHAoDO/F3fu+wIQ1BemizuEMhyHnmGC91pgnCfuyiUf1rAI0H
MhdlWEiL+jWhyp9dgaRfkHWjd40DTZkelrDutdCrd4b7xqt/k0jv+cFHImuQ1LwhlxvQgm1mEluf
C93cFT+jqzdYulIdyGlj5x23a9xJOe0sAXxjGpYj21pWKi66er2wFTfaLoD4ret3I9AnMKbeK41C
VE6DoK/EojHqd1sHlRwSBt4jDPyUBL0QFldWAVc5zXwd3bD++Ix/CWLFF22ZG/5bgR2pIPr9vajr
70TQuSadA4ilFrVm5G+T+WG+5ElA9SbKxKP3RxiQ3LOGgwEXh+lx4+tgbKG1sSzVCT1kQ+4CB4dK
fMzyHmyFIzGp6EIl+kK6Vrhbo5txujAR3gMxszBs32WsHDBTYYJGoMc+Mo2bTc1535HAPzC//OQd
GRhc1wZ0s5xm46tu1wD8r0zSIE4RHZhdR4t4DBtLwU4jSAML34M0Gnnc2JkB3HQrYDGH+LzzCQmO
dWI0zrLjM5Abr/z9ILkodKJxSYyC/nOjPthhFYcdcu37reQx7+XEZdX6BKuoOr7n8QSP25bah4jw
qIRyi9QnHkQHQCi7GnotQaObltKk7dStGz7LhKi/66+3esivfpcJk6vs9OMLwTUFDwjVaau96Qu6
WCV0o4ofeULgGeCphW4dNzIjyjrF46ok4xkmkktwVLRyLmwZRenmGdoSBsODLpltOruoFYSvXTSw
OTOahH5Xt1P5z87Nrh3caInnihqeVYY4pYDt9KSC4bCasDFm1p3/j3XvV5TTPKFBAVXxqt9xQYQn
fZlemeCuWskBOF2Ig0Q5H0GAvny4vkCZfARjErmZV8ZUjEgH2cHfkiFpBhmsJMpLfucbVCfdx5F8
ZuCm2Uae4M82uautmLp0/oGvmRJ+MUQ78a9SP7eGxnzE6ObDJ47UKuJpQXhycaSyTEUOWL1QIYvC
zXVPwCuxoEABlK04uoeZCb8vTNnQdSIs+XS7Vaoe4k2HlrktwedXvzb6Uiz/71ah+Ldt/ZAIM2iD
R2IUgrce1r36UnLng2PqqPPxTH5Q/T/cgiu1Rqls/uQbdBXW9Byup6B2Y7SfePOO0//hsf0YDjGA
goLTwPUX5gZST1pA6fst3BxsFstp5NCd4Q34DAf6r0kH/9OdAa9z8b4yTHlpoKN8OaTh0m1K/ItZ
rkaj3wJHgCECAnWoVQEuIY0zFAr0TjNFkAbZUcugwlGpdtE0ZZTsRncKo2pbxJRmslLqyb1a2M9c
ldWs5UC8y7hHXpJH/9oxR7nMpVVafaDaPwkgJXth+hYUnwVRsBAGWd4uQBT4h+6vbBjmznKc8GqX
+x3ldkExmD4qBBw3glmI/VcuqXB3e8BB8YMi/kPRYZNbwJxNB6r5Ujh2xr4f0ERsF5KG3hVq8zKk
9zdHlr1X/kEQ/WwNh6U35Zlo9dVlM6PVQWAt07YWSIL43uwTG9VDQxZ4SBr7oLYmO1Vu5MLN1w0/
4G167QuyAR+pWL+zycKpjzO0Qa2Kw+5uotgUpwer/sa4TaIKoMrBlxTEkG6o9VokiRMHdjCGSUpD
87Sl1QC6KjpuHqofbphF3B9d9kihyxaLvLDdbILBZyTpN3LaSWCRs4T/PgodT1BT9Jkd4qzEh5cU
PnfF8zz8gFxEujW9R7DkAzATzOGIvhvJWBg8OahJhtEIUexhf4ItYFZCPpVefekGVJlZNdXj2xVO
1pxeJEluLv+Y6jcTeT2NJsX9av6QB8oqjRmt+rAs9uITiZb3CCEJG5ts7vt4ZKOuRoJiDa2yBCex
UDLFCCu3T8HTCNZQghf0bhYszfyU6zRuJGStGvBmO+9ASq4qHnOpLIWw8GVhJz1iu8sFyFtv7G69
y91PMDajgIv4RcAzXjWVUQnL+RFK1cZc4wccq+RKFcnOOhbAIfARBJv1wTtIvctUIGtHWKRhjXZK
NeQ9GrdsCbu9StORQuweW/idVRFVDmrxbgitOZ3lJi5KPEl5x3CKqEQTlOisevtNSSnf6MHayP+f
fyzzMbQFGFwC/8emrbvDNOVQIPjmcEkM8ZnI9qiFEYh91SPnpQrAhSBI3x0g1EJWm/K4Gn/PT0kN
Rs6I282IlKm5O3l+HyMhlhEz7twzNZ8Sl3aM6cIYktCpoWCIu83v15Dmn6xnYkMsD0KT8gpKW0xX
Tjmhia+nqN+iyCrm4Q3k1gmImDk+HZcQXrha9+7BOFzafi48Qks0fYqUNKUMT34bhIBKKrGud7PM
cZKyoYq+pxsk76EYMy5i3YVGhK37uHlyIxJ/xRU2JT015pxoBCdN6/kTi/HWhjJlZ2VkuxGCZK4u
zverk7u+GM4NFdP51bVBpEMtEeAsn9N+Xn773hsagAO2PLL5wxCNX6vMVjj8DbsrvrEYROpp00gI
heogbpiHD1iQLzS8FuE2Nf03haFK08azidALxEZKDAJawr2ej01d7RF4IsKxxtfbh07yLtP9IkMH
bI7j8C4vz3nDB1E0SzxetE/oKazISr+TEKEyOrwVl3e8U+gzrLZY88nEmn06qmReWzkrPPZzZCQA
hO0VaFt32bg1RTaOmHtfMkEFZ3KOtVIYeY9CGezNDNRNOc+k0ReejaK0gFb6igfOMnYZJV7LuhpK
rijMkL1qx4IpgS+cT0ZtCdolSroemMKW/8iK6qOhH1nUzT4u/E60GDeDkydL0k9YRd9bZYVV8SX3
IiYeuhAgDSssbeZD8PmvTOjHWe5w6CTt5AYMgouJuBBVH54sr7wIis4Vz48xDxyi4T9JfAN6ZQTX
Df04xki4RTqHOn6kTMrfDstJWOxG+fkekMXwDS+viG8drVUrjU7ZeMRza6yU6eNqWVap7L9jA2Q7
r2h7CQ8OfdwkzE0UDnq9lax5IgjWY94mY/XZ6gS29LeHslezwPG7rvFfBBtzeQJEE5BARPgaIE4w
glYK7u8sBsZz36fMrc0rx/mYTbzlAgws8siCdtdsdHkf1HXBBApWErssK2o8kxMlL2FaxkCTzAcj
DCjgwQeoBRiIEdVUf9OVnBk1BLD0yLKC8L/88iF5fJAPLMIwqfEIAO7d+smjs6RL0JrkvPxjlLmr
YaNTSB+yq5gZJ8ta0yuR2yWO11yvW8nlIJ0xls9/gsE9MhDtmrrOACcgYIFxi4anfn5SpduN6dpX
RfJhvpad01la+XAqoJL3s9HGdbkMCUpLay73WjGdz3LI8aAjQQmi38aKD3eoJi0+XVC1gcThLH+q
ITh6/8mwchBnJnn6aMo9T86/qQ2eOFD5gD7fptVhCFKoRdsHaL9StcdBrlBQGtf8bK3xogdxt5e2
c0PVjw8f/HcJOjGr9EPOyjqEKmXCF2pLhZpRW0unAKicdCd8TqhKvR0vxaqbw5po0fDNWTf1NZ/I
W1C5HIlhFjQV1Wf/BltG74Kfm0d24sxqMKITKcfMMqvNB8d18JNal/dmf7XXBleSTT6UYUGbhuf2
NRCCVL2SgNV1vLpWHOnOmr03Dr7nAy/hz/NfFB/g2iACagNc4UmtENk5ZMJ0qS7zB+YvSr63UluU
zxrCCL0SCQR79zfbYyeZDi+++YytgnVl4ZNXCign3nA0ptiT23c2XV5OPi8o3nrQU52ulSzYAjFY
srGRdW9uzxdQIpyeY0Nas/WwGdYNaZ3WsUDo2akQCKj3A2lL3oyHizLzwh9n82QojNAq+FhfN32X
bcvOHG+0GWJ/kZIbvLhNtlN/apY+8DxYKAmXqdmQvNJyUtjtk7iwspIUBa3nUHir9dvsQcGQAvpW
CTIJrzX2W9fjNKP5mqLOd8cfL5haWYGpcyBRwlqPdGRO3Me+x4l9bxRtKegUSkY8DqDITVoKKxgD
pznM/tjQvAVXJdTmLBadnHt5UtD7TaHzokO0H68oGzGntNh+goxjTYxXgA9GxKFpAY8DggG/FHLz
v4Y5fLuPbErrIYiM9LbuB6dfPG/aHhDPkON8LdF3kP4/5Ytsc4iynUXEXOvuMh39yBofk7M0COFA
JPAe+JVe2qkEdKNtWkHkOGta5a5tUpgGabeVucT1CRMbM2xLcatwf5wCEdNd2ONI8KHXYVNQK0O7
qYWY9HHCM5PIOlbMlJMgR9/03YQkUE2HU2Sa8ra6vJs4Re8DqII8GOK9O9KXv9ibDJ/azJD2NOYx
jSp+qa9mx2kmEavqqRSp8RH3lN4t4JyCzlsNK5rhBYiLJIDODaUVfdOnBvxqE7JCV6YpEeSfL5EE
NfTPatXxx8TMQneMnCNdp5iSSZVYueAPLZROD10I85+19TyOUEgtaZK1X8EsjTqcamg5uSSX28wd
sgQs4qBr0TpYUvdwbUlVgR3/idFE/iW8pIwwPnVwSos7FhBwmrpqG+pktuIUq3zLWUudeNabyTUU
zTvP/R/LhqvuNOk5gQu30jN/SrsDi26e5kLpXcCPCIwzLCUzzs6H05GTZyvoWHpxw1eU0GBdaiCh
dhsIhhI4o0/mfjxjZlbhkwnQ5Pw7BIJWPlAltfYsKSsFZHn/VlkDAMabb9JS1kH/xIh0RX9+RRCn
1vowEY/YRtib9BIO7nxoj05V4+SSq4pvrx3za6gLqoOArrZW5DELiP8bIHEyuBxT1M8XBZv2TZre
Ax6MYSyi5S6aHcl4PLzYQLnj31jR46gHON15oIuks5tZRhzWuBlVkWFCvIKzYdj50EMJBlYTlvAo
twml3PNzYitpnNbYTQUou87TKZ/2DRwhsC8pMS1SdEElIrH9+wq0oPKGiIjnLEfSExoTQdfN3hoA
f3YdVjOznmdiJv5aLf72rb3AXog1od2kPJBmSmkUrGFZhMtp0EzR4ncKwFl5yL8mKXfyAuKPaa0e
VzBAPqM1bawRucettKlvuSKftvvg2xbBG+58Nh09b/K95bmLAo5LX5r+NoAb2inx/cI7NfrzUBUe
VdEQqGJBuohpI9jgNdSUCb0vNFbJzHjdoqBxiDzY3Q2MT87seBhf41GYlO/BgWIsd+KHMmh7QF7i
BQSAixGXsbzyuf2NFT7UWMdPwLOxcDvNNcXMS5lWUChcXKX5LmfwtSRNc3EqA+uQNRwN+NxSApTk
EmLIlPpKC+/j4wayfyrm8hAO4wlffZnpa0aK1fugeGMRk0YEy/sG67RcKsWBE9KdiPw/+RDe6DSn
QWpnIhadW+8k30ischi+a3UumFUP7Sidm4Us8SOgUER0wuDG3XzgxsNIvIoTCAxeHruz4v8502V3
5mMp35DJduCj70gySFjrgKFVrNt/jK1gZ2CbkFadJbdcYBr8+o/WiSFQtxlS7s0KYXiM+ZMtcR7u
0baGdwkD6xEUyH3U7U2fcXDxUcrQ62Od0nd/PzB0W7/Bbn93/pFAcJlwQPDJ9VP9eTXbaLzM1Z27
sTsaeLm7+JnRUA7kRFgi60dR2Fmae8jJJOVkYQ6QvOQ6W+t3aZOxmWRLx+WiBSQ6KWzl8bNThRm8
EyYhI1I8iR7riss4I7R+p6a6wtR4qhTzAwGCXaVkZNJgHeRnZ/PPKVEqa4/xuOuTChRFZ9/7BiUF
EvawQYE+CCk2+UHen6olsa5cATGWwf31X6A4ewv9dHhRysi1Jtk+IUuWqj3/og5fsyUIyo57kPLt
MyXH2TVzcO2uJ/P+gjN7FKzafiieme9TDxUU86UrK7k4faHtM5H5lRqqMGx3WWgA4CfUrk8kNeZ5
vcZLBvPCznP0hQJCTsaB+6lheZiCms5UDfBrjeF1CB8pnXCHVkenVC8zl+PpuwgMLfLaZ+wAOk3C
a8xRxCFHBDaaPhgEdpWtTiv2HkP7mDi8qbh847ReQcRf6/eDYDPowMiIV4FvUWAzaSFf7kvRLur6
XhzOs3M9txWP+XkWMoZbLCFYAIxiGuLrJHAs9xokVtEzRlKZe8KSWzulopoWI3+iHnDVkXKoL2kH
STbgI0pmGdpyd3j55KHou/xhKgMGVQ6ZUzZ+PdA2CJgXFjalZDNobqYsIsPmv2adUyxBdhl6+j+X
jdCYRCX/FeA0j2G7Lbds7vKGIPtReITZnEIbiSAGVaD/mdQloBt5KVfH9JWpLEG5LJyDJgewjGIg
YHJl1lDlnqDsL5HoznjDczzWZOMTTFwslolSQs7NClHnXdFACjBTOcESiTsdTi/EZ7AI8LkuPHQp
/8WDKBtxjSu+XTyFayfGd0noNrtH8Wi1m8Wer0sidgKj3u4SdsUPtkTPXeYFTB4Ck6dbnfbRekYV
Z3wDx5hjYJT3i7PAytEhzCSAcoDEAvqvEKEGkICHAo/gs4d7j8akfTKRcnwUTrlyv3Vzoa/tkqST
4Vj7oC3e4hKro7aKdezzs0Gs2QWj7WURr1erLgZLI8WOPt+kByEGm/ofBYraL3hGxmTrf0cljoEX
8swMwgq4GpYKLzynffPENqzyxhnlnahM9P/BXCEn8CVG8amAPsFIF/HHATIJ+GTZ60zV2FWCbDgH
XWMv9isSCc1SqcLXwOUpdcgq4Ff8TdIjgtQbTxX50xndUAMtepj+ZTFsLOdFUHDJ2+/mYjr71E9W
KwkosyTX2ZoGl5WXhYmr/jUmljuVYMM8wa3hPfSv8h6CRXjglMJargFmCjEJZhZUD9ifn6AauWw4
cpnONJnbLPOkieellLJ7MBxcSaIoc38FtU39Vr0Xy83D8qi7PyN7vU+HxxIStqvUXd6/5CUgLA8y
IKs2A66X3oNlo95uJY0RtV9cQqR0VwGJOGZ0FCEOgUU0HlnuSmlxZkyrKXYCrwYxQD8e1Nfh5LYO
ow12uTeXb1EkPFwEa//peBzn7kA/lnffpiCPlzuMg7vDOUQfKjDSnp+cefeEI9DdJ/e1yNh0wGfR
M3YOXIDtZNtlkPr3c8aIU1wbSenXthHzK7DjzRpffUqY9KxM3fDvDvcOg/7H93Uyoog602SkOw9n
KllUJE177wVykZrFiv1l0Fw0NIaOcDLAr+UPhvcNcx0XMwz0CYrKWLG5LlhBiWmOYeKCiZ9Nmw2g
jR80vfr9ax09CWyrLRGh7h1zD9U2ehvoBuGqvNa6pUEF46gXAe0kxR6HsA8oy706sGeDKFOK/qBy
Vl7Vj6aMiRIOBDx5zm2cwRoGMQfN/c1Q7YncRxAW8dgRV299kwonkJ5WnN8ytIfdT0DzbDSSjp6N
OVyGUtYY0B7UrsSEE6UbNhNgaGwiSm4QtZQ471t7dT5tC1bVRm7zIyQX8F/L34LdPOU8z/3X4IKi
Y8NFxnUpbUEbp5SJY+0CqLeoV7DU3m+WQYcRZNYUDY2VHlcSTiqswq+64m3WanYq0YEXQHaunTeP
sDku+eEsnyxPj8vidEBTzsz1oapeQApO/HMUT+D7NT1dPeBtREUE3bjsnnZ3L5jSYW3pdx9vMVGo
K1CFHz7mlQtR2PPpsNN/SQCZ5MiRZ348JLF3ce2BqZ56HvqJX7PGEysq9uNheYxo61tx/GbS5/4P
0S18VGVqB9zAez/XuJRprGv5vvOO0jiWotKHB59anqCIUWvCUBAGyw32ijDVaibE4bcmAeLoF2At
XDprPoZAfyCzig4lKDDO/chaaVYysep3ZU0jLKAB9yFVwMRMt1m5u9/H4F1PHm3DjA8niZiF3ErT
0jmok93qksGOmkEPbNq1D1s2WfdpzaL+vtFH2E0NW40w82bz4M5cIWAn6cwxwEWqky2/rO4E7PXo
lbpkquTRALJDWaIJAHRspQ2MYkYTUhmFHxB1ajmZn5tRgxEdg3Pp+U+0+esK0A6ctH3jd6d65eyl
dlQBJdWeiITIEmtqu8WcWGUiKplREQe5ArclSOc87jN4kWxFMUyZ91KOE6u0+zwyelUT5o7qBahN
cfGP5ZhqiaS0i2fYIm6D6b1P96FT25T4T82U7V/B1idTAuTNl2bHtSbeMVXlc/2wQMzwSlaCFc6r
7KcS+DTmx1tdoV7HlQAfJWTdrNbI6dcpxtOFzcH9BR838i/W/zm02F4hICOmX+/s9qdEhSEZ56pV
e5EbX0LI1l8ygpGly/+BOfaN7iYMxrhjI/9SmqkLIIOQl1rBu7JzUn9wnhR0hkr00eR7ASuB6+3x
B/xb3OINL2myto4CyiUKpDDM9pQLIuj12APTp57kI29Y6UzYjp7KsH2TRDi3YfuhFCxXrNy5A6EM
nKvAnVMBhKHcdFJls941edhlRi7ME2mo4vz9I2a6poZGPOeyq/g1WFDoxFzkidWD83NNSI4c8yKV
/FKPSdjEfSh/9CiVdcw0ifOSWvC4yHncoRSgit/xrwv518P4FhypyVWZergm/0nEXxUYUoTNXITG
GLWbSLPcUHszDvCRzhlmMVTzNTthG54gguwTa5fXBjJMN6FZnenKdX2Tf4cb/n9rV98IbCqD4N97
yviWsnt6ujxUQTSjg+a9ZHWYkvZ/T/eAUIW6i/iq3JiMikor3eKN8L0qJdrQVIySsDd5Atd1SKv/
dFWCyLF1BbL9fwrHeWg7tP76DXiF2TaDOCSNNTKgx4V0stLfwpyhYMlHbHFLliQjUV7UkAGViVz2
reFm5Euj0jw5RqnDX02lQbtVwJm4s8vrLdreTXcbq4J/FPE52QppsdrKthnS7X7S3zlOt09nwXcn
oN4cAIR0Z72jGyt0IBiFwrI2zsfgmXEYDBFMgdY1zosKZnDmx+MYP9LR4krsz+21AA2Tcf0qnJ3I
912eHK3x8t9r+z0LQwKkgtY25YyfobB9raP5ykeGUf27mMXo6Jve385UedzjeXMs5P5CxLTKyj4m
APRpLkGt8kEOBckWX/fXoBUSc7jWEP+8qLb/40VuoE4SkN1rlI7wgUYNeM+Gups7KL26Wo9NBjdb
KF0MZ9dzgHOT7DKtZ+Mue+b2l2AwEaOCbq+jtgcqiaUkjVMqJi/V2b8/d95OjQZV2a+ztt/WBpZT
kDkaxJHI9aM5aGe7M/eiHL5LOknkcgbfuwij1E9H3oizEjkE13WTU0B9q5UMhqJgPdgJEb8MNa3V
8jpR949ljVAnFFsTTUP8anAEfDXEwKkjpojYCn9cH9/ORE8+oNySFFOsP7tN+xbFSJBXHTlB4+/J
84+R/6Ve56D2Mp/NEdJ3X7uRk71sbBKYMiBo+X8UqDUSFggLPDGmPAO12xeG6C9H7SiBuiqDAE6H
fdljTm6tt/3xDUgSBW+8c2TfOcSMhX5o6hr8EB4aLwVrPDoqTgepW8aB3qUmppcNy73EkZXMYCiX
JNvwuId0xrbLJMMFF/KkM36Q/CAYHeOlgaIoQgPJxajd80WPeXVejMuoI6Py7ycYsepCjeWY+GzU
chtaVmqxqY7tIYb02yjpG26vk1Wtzc7+HgpqKCC640lYHKo0gYiDlF/4rqWKhZo8n9ybZPTlIq2V
nNPxmxnERAKkO+lBAti8G5ZvhvCk/yZozCSolY+ZQyckW9nAut1zCMtHenn7uTEckkFyQZZpDlMh
GbVHhKDywYa34pIZ/V2sbWu2taiM8zrAZiyRu3JEjx74elyFMsXXQe7ggpZQQWgOSngrQ3yCEC+q
IIDLUu3PR3NH4upgzPTPk6IFOP+phru7oz0TpNF1vPc80hQBIyrmzvLznhM9pmlNcGXshSOWY6RR
gjsjEz28BjXfZGDjOdvkWF3238IXDbdMnkWvTg63GkrSex/IhRvXZ/aG0m1YGm8PC8hyKqAkpcIi
7a7o3GNAqJRy044Nr2VVSDPaHKPuvsuh7lfG8VXaKP4ii7OKaIUXi11pENorWVHlkCjwihn0c/zb
VvRweoNgLAUqjDStbF1bnVtRI8cxRT9c9Cao5TYAcVY0qF0WfZhyh+mbAdrbsXYzL6hIynQb7bXH
ss48sY+uqLXVvvI1hgpuAABJQW58TWSX+g5N0gCWmyaXtFHyLpCtOmYyj6QoHSw0j2jIq5Pt1Z8K
1VhS7E2ipXOCuhPEwbrZIt8UQS/fKKChE96xL+crebXMloPzHjpEhNNLCAUguYs076hKi3FOTH3G
84oGiuJs2dl0Xh9d1L9rGgE7CEXUlO9pWXf4TnLvbmnYQhE2DxSOlcJxwXpoT9vpogeDdZB/dwwy
WaiFxd4ZCc10SvGr8A/F/gYVXtnezEzcKu7pzBSOBIGp446UAfimk4QMbC3fu3dhHbfE8n0gWi3e
1GuSn3qpuMXXytSerVpxubyKlu+ZmAe8esisCoyYuO8JxR+Og7r1yMjfEWlGSi8ajutJa4t6vXI7
aWcU8CGIoINleQieuMtkL7akuz2PlOEX1BFI+09ekRxqY7kKXllZHql7jxUEllcgn+y913JB3UtM
118L2uWh+WLJHMtFafep3BU38FGy0uhDhTkMrjZtVgZNzfrmhtx7qze7XyPX/lodIC20XwQz+kd+
vF0W3XthOm9K2q5dQPNGBuL0DIhaiH5hYq7pTC6FbGbFk6jVYUjf1djQvwqOzHg1T17+lkNXpT0Q
OLWc1HTUiWwqc/0wrx8MP7m4261qjyvLo0XLbaf7imSBdOUAr6SwKqpFrcqd3eEggfuiFwykPLG0
HQaDtjwV+nBpMMK28smdC4P6RhjRmZBdmT5oAqHQk//MeqmWmHBJYKKxJiwMXybNU1cXsjE9ob4J
rTqj8pXeYGEG+GzyDAVfge6CzwIUTwRWZ5mqpJgO1xXlGtvwriYTU8vBCmTmHS0tIwSsrxbsYk2B
CT10eDMnsYIxNn9UTILD42aRoXD0G6hJsvrjgPysLau+ljLuzMPbkD2vPssJq4xtpLjhgDH2Byer
W9Qj9Q8CO19aNnphVScmh+1MYCR02ErgOGEBk45VdstOOVKipRZT15F6qC8nMT2YXDHOLalM1vJ3
sodEaI51PNATD41htmqDuvWrZtzBBfkzXHBzjDpLPK7iIeoR1Gs1PFRJKKdK4aL+PPRAgDsDGCEl
jRmToGhmOqXLqAuAWS2ShJEvBvJlazgGLQUYgfiJoj5qF4uutSVkaQY3YodL76XnMw1OAhi8c008
G5sI7xqs7Al8nFcZRYElXdA7IN3fuE6/mGiwII4Whw0CeAXbpg20I9FjQR07xwDrSjIbx3s8fC2b
waITauuZkHKXUbjzUo4+rWClaharMldFWMQ7qfpjwVEORi5DI+macbD4lVXinBIvZ9ujsHVEgGMZ
tJZnPUthDetLTdXvhynicaF5k4y8YQ8b9e8O8qvRtcqHzc1b967ejQUxr4kg5Pl7UxeP2OymOxjb
+noBwvTY2EI5mjGJGBvURzo3douV1aXENsaNPgz1nG7ts4WvtmhWPPoottedJEZOQwKx4URcXFv1
lmLcTlHsIk+w5pddkDlpXniCHOuMSsqpMsqPbYEjGI+lPJDmAzcO9avgdVeotWW5WWg2j8ZiAre+
b7fgD6gN+mvvDnrekGBZazmA22RmjtiYfQVDHtpiuIkCRNegtf/t126j9SbrlV06Qxw7ErGy81Bx
oeuZoPQglljF7OCB4bLijtRHy3k8pE7C5VApy8RK+LU+WRpWBJYnnAaVadM2pXK1s/ZLysryIJl3
NEQ/TUFT/jJqPJ1KnILRBEDqSQYRhhPPC/LM7A1h45zH1NLSvyFc8Q9bihuFcYmwRWkoMfdRY5oe
cfMsRHlacICpbQqD7FYb3ns0mWBWzn6Qw5CFsRq2cH8wGG2DdOrOWHCp5d2U/8pwmzzg8ywkdKn/
dSr2z8ELRZmzp9Yy+XsMQavuin9ndDVCjem5Ifdke2GDrMxxzuUZJRFyre7/JA6++IIFcRit5Rgf
VfS5nLwC6/vRyGgUU+il3paHtTP8mmRS34XaPOE508GrlH3wW4JdHpXs/EBsB3SYHqPHx6tB0zzw
xHWzVdelXI2irLvB+VOJh17POvLnvzHXFJ3VOW2TJ0Ot+S1eSUWrzW5APsDe9kk+Nnp4ndrfaQe+
v+Ze8+KKXQimT/9jnfAL/OCChzSpe8HTk/s9T8mdroAfaRiekCfpeSWC3+VUwMoGlvRvNYH6fh5H
MCQWs3wScsa5y5FrLLz8hzwBip6pxdR3uHXxmJllCuO1eNL6LiwW6T7iiLJ0t3BxRF1FxQ+CM8LW
0A97vmjaRU0lMcNrwRjZGQMIQzP3sQaCzFBD6Ejh6hYpo5KBmbk/TpaYkdR6E5GN+NVyxtTo5uW6
bDdbEsJzw3W+KbSNIu+NXtwszUXJsfqVAXme1pc0rIVw2soq0JgX0zw+W+TbntXAUmaMre/whn8E
qU8izytG9+x2ID36xFxsZrUzKEl4LaFOE7GRoqRDNcgCIarMYyobhO+wd85wDF2fat5rFQwEK9Im
DrVxGDvw3BRq7QgNBI35WUFPFrl0FCgmcdrrLtCPTI0nqdYn7VH4kdEEc0WWytp6H/OtxSgqie0l
7e1ZoSZsBwh6GEN9LDR3GZ5qMLf569w7SejrAMFd9OWBKF4mGhHvfq0XEx8zyCj1N+zxbDOgxUZm
2bE1O3okd/56P8awHY8z75kJX951rAweqlUSvowEdAsHFB/hDNQ2pu0ANHU9vPmIDzkukXfw5mSN
Xk2hYCWci3ssW9Jf0hP6ZYm9zf3KkEa8Thj6ANqqY/1R7D1OwHoIqpyHFCBolPyL6sNEytdelH7N
8tS3OQ7Gu5UhfvefG6Xvfk9My/HUTw90bdGI/2mYH79uPZOKnaWprOJK0nPMDs4RmG0J3caY6NE9
Xk13p4+okRljlMqP58Xw+mEelSghRWi93nGyrT0ltLMst++/zVDYC/kys4QNR6Qm4JpUft5gIiQE
5vikRST3rYt1M/oGKD5Roa9nWJWphBrHLF57rakYTClTrH9q+7hDa/E8bDwQwz+SAEBEloJNjMri
SNcVaP1JYCyT1NTkVut+qSSTvQl2gmkzFZnIiMz9Cqq6fOlgFkRgDhS+tY/KuR37iF2oZcwmQiXE
AWuRoQWK4WCSkMNR8O4gGtcYGcS1+xd8IwmRRSNL6nWokVvwEbIk56bzWpa4DeAOmr3KUtaDkFut
UHk/u77X1vBcwKdZnISBPUeU34pR3AAJoJFsrU7k3iEUXULWNfcRpCL1vfMKJQmgjER8BBrJwlnS
eNjp3xXK0JHDII0NgrgfxIgXHLHfcxkN8abRFm4ZmTfHQ+yAWoQj1Yk0OAqWxit62WUkE+q5n2es
JN/MyGN39Egmp7OooyJxEp8uF3676L8zRUb/D0zxaHiKQNaVadntP61gcC8zxVtgaNSySbgSmBd4
FRSr765P82C+Gra5l8SWpnaU46l8ffrNLpiL4J0VYlnw+XgpVanKd94qOswgrKS/0F1w1dSmCEBu
WnQms9BpHxqooq7OweqxrPvJNsPHIir6s0zp3AM/x9O+wW8q54ZbXUM6SFuJMfdJfUYapp/VUwlD
TtRkjeaebc+g1qS0ZL4jhARNhaTmFF95XxvoEcn7LXVtJ7Q4VlA8QU7TzaCa2zOxWzmb5dmEmuwU
+ua5uSBp21dhX6+E83FnFwDcm23za7PG9ILGiKgVMijWX5HBniavRT5DXqAVjtcjK1ecPWD4cSbu
AgvL5s56i1HiPo7OO3NBdoSG8jUrBIOmXaCNzLUyu+ooO5rxLQLLYhHrdQRgyFLfm1A1aS1xp012
Jc8fsyO8gPEpDqz3FiGfWcRHgPhMzzjNozcUqObOswho/HEWlq8ljlS0jYtvx4KkNy3I3GFVF99b
rxjg89UMrildSGXIYs9qGvNMbcLHRqYJYGfUAgn104JCCgXT8wPpz7ziHEc46mDl2Ssq/gLtqVUF
r5oVOUwrNHrHQbLTt/GnSfaIvCid7Xf3zpjuAt0TNZlcxgi8z7F0UyKmYz9Cpi/0sCjaJyAXoPRJ
IxMlZBUBjHMoOjJdAkbevYu2JcEap23ZH5xr9gpJGE7DHL1Qzi+qxUpltVSg1vuW+qbdG8RIy0GY
RbBI1m+I3esAgM81T+cK294dhYLUGPRmQzYhQtLYBaX28rVFc/AHp+bShlc3yYodlzdg7iWC+1LK
T12AhHBf8h2yNhdGLpqAuBrq+ur0CKoRey3MhB+LMDRXBPHj02/uAoMUryqYiwJPdbcQ1FHVy9qC
SlfbMcSUWcomiCsCgQFFHxAArubWAGi06XuvwzXw+MhdlUHxDdXKNChEO6aWQdGhiNoOTSGaV34f
j6K+J13ugX1zCqLzcVLzIdGTPNTjboiTwnNcIeEvba1/0h2+s1op0qW1FUvWle4kWgWaMBgy5znC
rolhgcoqmDCaQ0mi5NDjZQDYUUg7ZOnhqD1bJ+3GdclIK+zh5LdN0BwshGbqgt399QKo8Xl6ET1K
f8ULhnJ96nMKpmS7mhY16IJtweUQ9tm2bdyqlEV1apFrboLcb0ZzzlbYG5ErAPKq+6ha1w6GkTxg
mfPg5fQeFxKhOn12/c+ppnHYVRkR7xg1PAi9cDJOUiy8JKJOKeVdk4uPKko1uWknZ9o87wss8HbA
7hD46NA1M18xgdzIbgDJFaYlytdYeLTCXJvC5khNPWqcDzEUNBNfdIkDH/Kh0G8iaZPCSgZg/E4M
fdr4rPBf8I8bWRvbrEgRHQ4L45FMKTU/y2dm3VjfYjs2/GgiIFlxdAZmU+ISmPmwxRIbmIkgjw8w
yN2HViGCYtakTOlopOlKfUVX523E8k7Be++SHXamzrHsEvoX6IOLR54DOBjPSxrTV+w+/wj0uqz4
9Ke4IJoFWn3STq3FMqgPk+uDR8tbzMmi+clzV4wZ89ErYQDreiwwu8xGQLwxINm7ByIR+g4XhbIP
HAkTzaYDprJ89I+ZJednCiakShwvz+7T+/+g9jXB6YoSnl/MzGP4ongj81LZPBBfKOIIlhX5GbXY
kGWW/YhW+1xeqdIkFmW5+oiDthhPP/GadC2k113aaVEDNSGhsNM/y5mCub7/zJVjS9UUPEryLgfS
gwHmQa9qQ8PZC6eiIl7mmektmzDQ+uiaz7l4ZbLy41C81Y4ePmIGOkL69FZQoFWaGYjg8TLPfV+v
Wdbbx2L/q+vz8vS+wraVlytEu1rxBY1cOtqmQF8Gzx02fnDS+Eb40mqEedrGl79Wgemz3TDTFgNo
BPjpXXcYIR6B+Yj4DvMmopAOyfNqXs3nHqp06mkn9UAx0R3jxJAUfAWttLQFEai9k4iiL2Ov77i3
HKZ9S4s59p4QFkjCgSYkN8MQLK/wGz9kKvezbVn1lsQm8p20b2XdBzSECOXS/YzIERmRQeAOHCFO
QQYF4QxDkbs5pA9DtQTo/uNkxCHOscBfYubeNerJKtI8i4wkQWQN84nq6wuazVn/3YXWagTfWF2W
v3uF4MyabRAKYzvun3PtbjREtY1oPTj/FH4UrvBDM/Ma+6Jr/WsNtCAaXX5DwsU6lTEFdJM5TTM8
S6kLEN1u+2QEqApJW1QB6e86WvvLvywNbX2PSBRb/iMgNNOKUslUrMNzqMMl9qQlUC/mwksUh/XM
AMfIEvvNWrZNQmukVXEMrH6Q/DJboX+tUEu9C4KUtdgr69DyCm9tci58ji+kpJOQs/+YMLoLv5sg
BYlm3d7cONPKV/SCyw4y3RAWwYCSAdh7aaoMgYNTSCqNHyiYzjIwLqE10ewANG1TiSYVdpPvMlPK
u9FtdDrJb2W66ok/aIbr1kE2xhKwtkhVz49q9YYeLst8Hq7Y4zo227d0+Hlj7cSjn1r3iAQsBPkq
0qcYLDNdKWcump3xZQKw0eelhDti+X4f6nnjrkm9mlNW9TsNNkdroSFkt5nKVpiUs5H41Jxb8nT4
oDlNa+JrUVEfc+fpHBH6Zx1TBD5rfa7DaWRws8aQsoHu219nmYnBKr1Uzdv7N/XBsshXRVJLm9kV
BF59jaaz/MTWlvIbzeOcU11nM3j7vb6pus83mgIEI8dup0tE4kAg+1QuzOjtvNjXpuLz+5R0WiPc
vx8F6P3oDpUEp8djVxTzQIHDX5U+0FG7E3p7e7J5jQ/qIqLyGjJ8IY0pYTXLxd7PaRDFWP6FGTgn
SKLh62WrA1GLKhRQd54nBECGC6lZW/9590ikyNA0HqCRph8EqNsJcanocjOMWKrliVjqsV2m1LHd
vD/At4sdYofa+YiCiII1tuyOYb9Affy3EQ6t64eie7eWiGH06Symo/K6UOBiE6jCLEp05T+FSFCu
68SevASMJMD1M+SEsN64X0L8o2lz0RQ6KS9FltawM0FfY9jcaJZ1NRDK09nGnygaF5YhB/k95k5H
ityUGimmW5FBs5CBxJ1CrIBtAuBBpGITv98Y5lLsw6oaEPjY/hy57gxNt3f7sLaZq3/+15aZUY5N
UUMXTO/n2jLnreq4ehzBjJnC3YBDwuHCrcJ0Pte7p1WISDV+66rRSsFkJofiu3PHjDGJ85XVJeZs
esqGJ/T0vx99p7+OBGtGnrQY70/iOqctqRoKTyeAmaQRQtZTEx301YhKPpZA2E6jlez5pSvrk8HG
fUQhRHmIfOcxN2rmJEO9s81LdHBiNLdzYIK4Js7ujJ0NXXFcWHXhkgx0x9sxU75bX7K6MTKbt50y
6qiu5kWKpCkEovCUrwZM+l/E0us6FYsxqDqu0/kta7Y/Yd29JMw8zw007pwY8r72M2tzkPtcdRsT
F2laWuJzmgfYlht/DonBmdBTjz5ynsoqyZqXP2C6NWbZXYbfaSkvFlE/ZBwPIb7UZbFz+fnWUQIG
dW2PPfGyfGIgGWRe0Oic/69kCpPyqV6gGbcWlN6LD6DV/eiWC2U9hNfNIOVYELk5iQ8x91YusSyX
ADgtgHnv3N6tkgSwoCmjOW4/oOnFWC28sh4kLh4FcyJMzjOVS+r67TELruxqOKTP+F1+nuZH/6YD
2R4LGF3+7EfAblEvNlfbf1WMzoIcgYUCMxe6QKxvbux3UzSY4bAv+0n2oIukk+sTP84y7lUzC571
HSQrlM7g9XWovvPLDSxCKot67evLI6Awwj0rgY9PhfSu4sQmEOrH01v589IT79ITk8qjzU7kTOWu
ffUdShiX+dPktdVe7EJzxchUr6//HSPGcEi/wWxzpXulx3gX0aXR7uA5MZXnZF2bgsT/98Dzukkl
0y4rWzndazoCRlHv2kHsHBL7WJAq83OdANq0lXAO7l3LaY2pE3PXuVClkcYz6ErAZErl63zwGNky
NLU9g9HVBxtpqFC6fwoyjIbKU9ZoDGtInT3sdUF0PJOW9N0/cAbAf2N+5jjP4TMPl+MRO8rklHfi
PcHAMVGBR8ziyE5B5412Wo494zL8VdBt5ELE1+9F9v2j3s4bR0TqaTJjWbevhQkdgaQ8zEUNp8+R
VSLL61nP6vKpDjzDzp1y3d6V/iCWJ8lxg6bJhjE5i9Xi3OhLs6g1QI8bVZdqA4aEmZXEbdgk9nqR
YO9QLzIuEd8WFMzbxcj0Jtt+JqrJHApx9vfkdgJb4MpwD+4XPFkY7Na4yWVH6Zigz/JIUNWSv5Q5
3X2KXOOyEh8eOKmbchQoWr1rmIE9wSW39dhxxbHWZpBXPXvHiLi/xSu8lOUfS02/4pByWZ5ISxR5
g/Ois7+bspm9n0TvUo8MpzWEhcu+qOUPnUGbDpt7GcGo1vCt5Kq/uOO/sc4JexRWCiMd4DBzdH7Z
nsW+KgH6VmphHV32VlMxZiumMc/LW0NEaTifJ19BmIK/uSeAiA2qQ9Fh4xQU3l6AQdumVcrzVTOQ
+BnAPdUYDvlqHPYWX1HzXrv3fkyoGLw6rUgp7/vyA+mWCAuJF74YPfpNKXjzj4yEgTDuuoPttkL6
ttHOwFeEE9AuJi7vgACK75bg8rFkQeL2QSSHvOkIowpTZRmjEqhi+7yU5/EcjTvELW2IFTuSxUZu
pAO39T3YLiXt9nZg7qbqLiwmbL8VMwPrc11XmLyqZXDfvdrFDfH2EV8QiP0huMKeVohMa3/5M8YR
UXVbtim41dl3xlNkZiIdKEYUWlL7Eo0bcoR7mF2ClX0B/nLkaW1c1PNGaVt/P5M2S1LRTO67hKgU
DKsWAhbi2noa8/Y4ctQ9XCJGo8lEBCSPL1/9hgeOW/Ve6Z17dd9vw2penoLZROoAsSqonqmU2D4+
nptYbrHTE8UPDwm9FutUm1wstkrrXdNdK0plQsOXEQaERlSZ6VSaxP5HYD3YFvPmYYg2GD9DiQ/i
2pxJl4RUnBOhYR0AXmx81O4ki1ToyQbaXw2yMOCcc4RSo6JjvMSZDufzfh/T8yzC6roMuY4S0Udx
wb2Ua3amtwf0srN7nOfMdI5OOpzyaNhHd3ew0s4KKFCJwpEIKzCpdgY1r4L5mk0ByQUT8pvYI/HO
c7yhYeBSRLjvaTpIR3xpoMTH1HIsrpIPX/aBlK4C/ywwSzN9BSaBbZlYDLgR5M7iFUAa7IlxsYvi
rVLwLHV5rMn2Q9l44/iU7P4pKOS2E5hz90Lm7DHQlBP9ivFtXP6ky8smNxM1u7gRQQ6KH4lloorf
TZfWrS6MEf4pdmf3tz/bNPRASKM6XGvKpVkgU/LynMvYmw4wn2khihE+8pnHJnfVMAscUjbt7Q16
onIGU1yqQMAkwLMxM5BQc+5QUGsjTlzCS7apbr9XilMcQU3i5fU+I7aPdS86fapnGHSXl/UsKfZR
bPbz59EHhsKhJhETQCnSYM0+WIMmOm/hJhvnY2H7SEa0Fg46htxb9itdCbfvlE4PqGzPcpOJlT9P
Tte0dNCIYvI+I+pUP3fPPQLamuEHJklUEqgAhi51OsZH9JoeHpI2756BbgpY3UzE7eJkit3i0GCS
qC2V1OkAEw83+fhOoNs3+FMEw4I+E3ProAEN1nQSrcPAxvhjxdkC1reXTbYJHMaJVlQ7dqUpN/PY
agN9yFqix/0Pf2JjxQRH+G9oX1Ts3qfN9R7dvsjrkheXOm0enxq7+juNWSvF99HAyXpWycylrUdq
HVlGBGj3DFNcwMoicIxkmfiG2eOYsqJKtqCffuKdMdCNnbGYuJc+RFuj13T6xM5FHsqZnt844dtE
JQ0T4c5Jb1P7K6PquGP6xdpuJKDtdycyfAmWtD7eWs2i7SxRB34HdZAnNSI7IMAFG7LjNWhy7JTv
20GvtdcwJ4lh5Bj7WDyXCgEL6yGD8NCU0gaOEbwKatIjdyM0zCwQCOb9OI6ME2zjlT4m+MHFh/uo
LyOSsfp+9GxLWymJMhHhop1cm9dPteQ915I28bphI5usCASxlX7A3V9n/DeZ8SqtRUemm2qOSnbI
FZOSsDTJLP5f6QlnxnJXktNhZRRf8+W/PR4p9KhUXH6gO4+6M4McHY6ZzPEaRil5Y31pFTxkkYTu
LsodRXa8Vo0lZtn6IHNFDH6VTfUkQLZMijxq5IeiKx4KEn/6g8xmuRl76HBnglWFokl/dlVvoCgx
xQsh/jsu58mIbssLeDg2eAGA1op26Ay0EEjF5f9UYxybZinnqZ3COgnY1+Mp2VkEu6KS/PEYN/Sj
CotnaX2T4Oos4N0X8e9jtt7hg+lu4O57cRHJAN0F0/HNPzm71d6o9yhAKOpwChtYdkLB6it49okg
6Ckh3roz8ZWUdIc0GPQugxM0eLeYyNWg8mtaBsC7WOjCYrZpgpJ6yVbkvf0+mTnCy0V9VQcgKhU0
Cv/0eAAALAVQHy6x5vNvz6JPd9KoszyR3qqVpjHOiifDYbsnqiYFiTBpAFuR1j+fXnBWp+1fEump
DqJB/2YxxtjDd4lnuJ83aHVSIXY0h9is44jY7kjkKYmCdQUSKk7mESO3aSUQTezXzyPrm6oF8O6B
L6L7FnYLogiLyaQ+if9UqCmVsEO2Pr1/eCQtYtgclIEpZ3a9hXkBpZO5os0qBKgZ54uWyclyqOUo
/sMcyTF8YEUotejJ8xFGu17DwatMC7tgky9zLUMmgRmN5orCbxfE+RewLCr0bgTRvWQ7KtngfXOp
LGdxX01om2L1a0Jjg1Nc0lU/0TyBGaqAVWzeQmpCsMUp4nEXqr6qUvArkL8VCRiovBDXyHhvC9Vq
dRGmGbEAsjdHcbK2flAcnXBgIYRp8BxQH97A3ptEusfmGXNlEQDsA6q2BdX49mYWAXG1FllK27Ah
Ry9dir0nRg6WcG7lZzY4+9RsHs1z5YGsRG+KTA+d+AiIq2kqfk+aALqFTKK5TVADXygHFH+xx6bM
I9LgjaVfAgl6CYSSWFZ/Ip79Lz/Ygs9rDgfGOCMW3wy2oaupFRaJqArbF5S+VHBUgPxUygXpBLdy
7gfLkRMrit/3quvk+ux2Bhd+rTCHM3xfpVbcGDMajW24NTr33MTTGtIQtfHasu4NqVlSFDk+MZV/
fEK/4VwH2WJ4voMye2zAKN5sB/H7WYJQMuoNXB/IzA9+f4EUEM9M3+RusdEJjwSKggTAvs9Lrmmv
I9b2NBb0nWhFYrnxxxXmK2B4Kn3Qsa4BooXOlN69GsS2cmV2VAASizo4i1Alvf6cdWjOaFfj6cb5
q1qg/mYzcbyDLaE2OJ9BgIcEUB5RPknBdDle7MOXiAt1cj+aOtM3iKBBSALrq540DiFjAR1fv0bc
K89fwQd3ue7NJpkc2ZUhGk4QyS3KFyeTBYuSidBFq4z5puuuFRUntd5LLQSGK5qEP4XS5GTR2LYN
Q+VzqjUfdnOYOr8DvL9OA68Qu+Ft232ZKt5330TlcEhAffvZzl9yykNm7/HFyeyYcTGR2aZj8I18
eltIkIQZsyPDqbAUh9EFKOz9DTEU16m+CJPChUlb81PG/LSuAVGY570lKIqtAcDdxsmOlQTG2cTm
bUdhcBO+8Sfxr/WD6gLyfFWP7KuqtMqbtkcFdwigk8AN9z6QUYQDY4x6+RY5woscFBUWUci+zYEH
6lQJVlHpyeFTV9qHDUi9vZRBMCVsr6W0YHlulkoXNSK+rGX7T/71JlvEe46be8k82xrriQOP+e5g
4/7UJWYMBHqRr64NpGgmy5nj/dED9Yk5Zs9ZwsojPjW3wN1AOanEnGEIXMHJrLzRaDhSZGXLobxe
KTkBLFqXOhrD4+I6G9q8nDFzNVYGKeCqzQrvBXhQS4sq19Ex0KT686xZRRji1jhNsJI08vYPuyWg
jSMxlr5JbToMAkrsRYLmTkouCTJf/yDqQOCGQ+26QMLqjw1wqZ6mTd7pggKfKYKXfLgAXkMjoxAI
GVbV6suUA+2g2sEOV+n+9uZQv3nbsSgwDAPG29+qdLZwM1xEsk+frrHIV5reGjWXWi5j1/NB6Kcu
BxvRY656EsH8ngvOEIiZZ47e9y+VGQCGPZvw6sAHnk84a0qQJJ2kY7wd5QkVY2PzFRxSE0LPqW9G
ql2lY4yRCwgZ2qnTA6Ba7jurChY4lrqgJz3P7oGGFXEKbXCOiSHGpOwWe+iOGUO8QhFLFVzajX80
rIgYYACtJN4TJMdnmVNGsO3FQnhqhqgz/+gLkICsp6fN8fIWmrdAwFyqpch7gfzj41ckjt0fLxst
3G6FC28ydzbbioo6cXttYCX0rqxMsppBoKbGnMe/jbKlmUwe7ZYSuxrixv1sIGlrRl4TMamDrYyW
kxAzP41b/BbfmjAI0BttkDB+USAbfoISLmIfHikvAd7JlV24CJ4WsfJl0V46JZH3lULxzdG8AAVj
aAF/TIb18QhFpJteJsiGI0DpwlAg2ttrIQXXRO9gJ4Lyxvo+tDsxO5AsrOz4ZUXJ8KvnmPOY1s1N
ClJ71d6IevBaDyZ4/6UBCkjLJqE45TlTsEkoOudD5nVgxq/wd+/CdeE1zan0yN617DutuohU2cbB
XoScAPj/OVtVd7wo6/Qg44SeG6TruScCbUBjKxut5xf0e7vgLL+B1F4rIzFOH3Ub89tS18pSvfMX
UJtPDLUgPEOaGCiCA3eZqvvFrCbfaPB1XleMbU5Sj7qSIzD8NOyIw/lqBRvGf3b1YyvO5CWJ0ZtK
6hFu2ocWhVjKHQX793JPcyeqgILk3JjpT6wvcFe8XUPmLC8zvYSqcEbdsCWpi5zfCesPQkSO48Pz
UjjS/b5N9jyWXinl0t3x+u6kDVWXymmt+AaOD56ENxukbOodLV1ktCzzyI/VGGeRMHFBw9HpP2go
ssLE13ZcssmyaQjPVkSbEeO/5QtYL7fyS9TY1KRQm+qTWxER8MY/2NB+DvuTuyo/NsuGxwl2RjH7
Vr3ihmU1qC/JFlGUbKUXB8tsVNLS0Nm2738nj0r6dEAOm/T7A9oICrsOb0bAkuVaNAXNKf1TDRp5
XzD4/u8ocQFej2ij3O/BIIg8H5KZaGGRTZpvF1f1/cuoKX1Jyo0e8VBa0mfAPkcQutWaOVeMf+az
ofzDXMJYAQCCjYKo/q9tsrrL4StYJVr2dGuHOwAkK23U7BS3L5yQZuqwTuflXUbPRrxF0F3m4glk
COJrwqZf3lqg2RkGTHS9J9O27zvCVzUJ7lnbeYkW7p7D5/uWOUsmdpZKwqkwEL2H/j9DRZ+luCCr
v11wieniajsSMG0LMqfagnHLQ3RC/cjuQY+8Ivy8PPstkbh+EvfOigWMczFhBznh3X2T4F/kxqxe
O2pGOxLWdRM1GJ/VnAOOE9Mzm38S7Z7nH+X1vjFSRstExehsdYEF4mFVMUyBWwZzaPocbnFN2FQ5
PqiPdMj/+ItdjAnw+q/mK79oLCqVLTq/oHJFXdubKl4G7t/fFe1Yn0NUs5ahGXXamS5AOE8dtu47
r6ImdZ6KpLQAm4UJRZ2FujxGCOpvI2oJ1VZvcml6zDcUcoaKqLpk43jsZMhLokhvV0N2BbYCsHuQ
vOQ3CQeDgRqdmVy7OTvUq/k/WcuoeUnoFMrN1gMVW0lt9Tjgd2vLzrwPjZfCbq7VczdHGvwZoENO
UsdR2kF3F4yZtm2q+zdZ1J9mrVN3YMsHy5STPpT5/2w4jjHeVgMkogySLs+O37YDcDpp8m+zwHSD
zotusKv1YzJGoYKjplY3pLVnChrKZQ+I01MP/eK4Mij6r6RA2tY6rOOxEGiZfyZ3DX5AJ8cL0qya
slVH72G/gdVcawPuUDQMMydMP3fs1+L3c6GGEmFdaERsEZGgAzjq52Ss478rAMwblOCanPYX9zxk
Yn1Wpl+clcTaP+jEJHWxpO6rQhRMbyrSlN+K6HnZB8uIgEKJnetJiPqc38f7icxMSjyXOCVNdgyZ
E1ayppPJS6nJswgPWrdqRQrnpJ1zbI905KS7vxoyQNtEhF6TfvIilKQSBO0YaC78hwuANktWV6cN
hxtcHcde8TEg3nWhwCWx5LEJtGYhNfipTCjZTgP5vED6Z5zHFUdzV6SVM+z3zwujdfWEC4zItST2
2IgL0NJqXWcw6kLCDSWYkfJREWXzoGfc2I3Hl279hCvsQ/pgIHBUT8OPb6aEmjN+gQpI4Hm6uDsx
U/vZosJkyfkBWfQSQx0eM+qztp88/Weuo95kdfaurWRiDdyRHxOq4fbA+W09siFklIv0ebAHEw2g
WGx+HodUwRklFEwJduIseVG17UECfTOGCMAfPZhJVarNovD3FcE0wDe2Qw0dBBvvSAW7pGCtwxIX
it4OkKEW5oJPufdhZpVDgvmaD5AdhHAVbKeBeBa+dU7E5niV5tyYgoX3c7UBYEh9FVmkyCB/+IDn
e2Zmnrx5543N19Hacz+fx9yB6xNNSDnyTReWxyVQk3rGtJGs+xf8VDoswcUpR2fXsf6fOqXXoGu4
i4GZUSpdgTYlkYEYKzkF+e1ixXkGI6xhDJHyRUlEQ63sJYw/43Flcc2uYKMsYSSrICZCSBHIeWqA
iswpMx/K22LyOorF1HFInAXkOHUlXmaa3O0QCMI+X+HomymaYY6SYCVPm77L2N6gCPqz8kTmoply
O7BV1lIRcjte6Hs+ahV/BlYZnx4vu05Fi9KPA/2HD/W65ELTCTcZnPAuBbPr1/+7hoaxJjAQhHl/
glXgUZLjSfAIruVM5t8h37H4XOQiex1egwPAcfGAM4g1k6/WgP2++4XYEd3CcqVqnhQeXx8ejqk6
pBC/zhKlEAgjzvhDH24IIDsFU1uxUYm//iTJ6M2h3WZJcN4M2V3JumZqCG+XKBx5rulEFMGKm2tx
vwTFk7NwpEhZ0SqtiQKXQbL1GATWQTPMwPUNdwyXkNMw6saupPsxZ6yTGtP/VS/sVFqnWRFf44X8
0oO48EiFamn2qksVGwRbchcoSwh49xIMYs5sDh/Xckzy36TmXsY9nVnrjIpuJNPQWTbVuNAAV1nY
UkcwReYdyJjI+50c046isf0PkQP8A6Lr3Mfx1ISKKbEF++m7p/sRQ+JVXuf851hLuOiVMVMjPnoA
0wdwvY6OZDFQNPBd4Lz8nVya6RAJfhBVlCD/aSGFXd06ZNFYhHDHRTO17DQT0NUeVrL0VN+iaQ7E
NoUYOg/xOv05GrP8IEsHaFt1iK03a1lBBwHzbNw9RQHqCD8oqC122iip0P3aMCjpvz7g7sT7VmEJ
3nhvbRNNs/XMsyznyEdzUfJtJeavROaKsEb61IGbT0mtjAwXHpYwjhlyC2Zt0VyRtGa1Q8idX17W
+NwtpH5jqzfsbs2uoiJzF9wEv3R5pOfkkvs2vFBOX/mP+X5RXbiZOXhDbafipfnFZ2l2BejfpYRj
gu9kfZwuNEG+CAR+nnLCrwr4CLvwbJZbeAWCI0D/oIEhXc9/L2GXTItJ099sPruy3m6i6zlGy7ZE
2Q57f9ChgelhCceI3p0ZzJtN8W4Sitsymv7lLvZ6p6tJjAHcPv/vqzOqWFNCVYJhefLgMC/Dpx0T
+yVtJADrRXqoF+b6uvFoXDyQCEheTMPJ4yxCeEcAqO/la2xQDZW6yjfB6d6aSwFKeNrAfH+DlMD+
w8ChKzn38eorIbv7GBPkfNoMPFbJ1agRfaO3dufTdQKAkBeSZNuOe/JDizVh2bJXKoq7m1pn0/PN
BTT7CDl/m5sOt0VgMkJJbv6Wxmx4OHK8rAl+u+ZxzaKvGJJZ6XoTFr9VV5HI/Y1i9bUIuA2wf/DP
eRmknPVwxntNnOj3TlqJ7foOILzUBrKnapOFM7X5XNVfVeo+Uo27nOmSC/aXG5bUjagNec7/ta8L
4wVqwprVm+xX275recdDjwKNG1YE3a59s9miR6ztxMgDCH60IRa7Nb/HDHd/80AVUXDP4VQxtk21
yp8dafQ3fj8wsbobRv/S6FAxgPM3OgYk2nFNMQxfUKE4d63nA2x6LT/JqNHDtV3PuI9MEDJroKBq
8FBOpfG0QfmX+pWdPVMiPJ9XsSz965D97W1bEkgWznFgZFA0gYxYvxj7RdCxqXpz8oMAlPVOESTp
0De/3zwq9Im9mUJuKeHLj6oitCIrTRgeKaVixZYeuTcQB6I2xt14A3EPcLRkKdpXSrd3hpKV8qjW
titkzOsvP0Yp24QQc2Rcv2vPubkc4WlSyphAEVnPSXt2112U7mUsL/8Mcd6KeYkX571t9WzNNB+b
7uEdLfKXMFk3lyYwWCYBa6WUqbmRrBg9YQsoCFjxwJFYUIJvEtsG2YCcUx0aUh9mM1JK4sN7x0/N
lUF0RUXNLPQxr2ZGU3HQYnicbsryMuMfYG3acYoW8u2PDejNyENtT2gBrPfYgHiBX1w6kWbaZYjo
zaMy3q5vWaD41QbIaZO3BoyZh44hVkx460JMH8dbG6bG5tEdadAjCTT3fV3pNRnsRzeJlExa+0Kb
F/zIvFBnFAKhhRnZMGeDvsD/SWgbDBq35cUOMqcgMkH4GKoNgiu6eA8kSt6xiGAfo6qW2VDizsEQ
tKqtrCG7pjSnnGbhOQIuZDKtoIChG3xReXRAHt7Mr9LkJtMqxwr2A94knhK20nv6pr20PmwhbxqL
cUqU+WRKI8s54PRajiE9gMBDgL3e+R9dqYcx2MummwHQAppH6jYX3D52SFU/8OQNRRE/hZRwpIHx
hS2oKRFR4CUIxTv4VPCkW0rSE6L9hsV0e3imI3whbY5Iv97Zb2ZbmbCslTO7NMh7RYwODJN3jVOQ
kbwOnb1yzUNY0GAS4EWzTKfNM/rjjiv9BEtOCYV0FfmA0eE8ESalToJk/XVWVhWGChWb6mFEP3KY
fJL5p6CpIC/gI1ZbiFmvC2jI/QhBTjZf3py4bD3QDG0jxa9EktOjjRoxVtmjbw+cOHeXyouNF6RH
lAPtemslSIgmJy1eXdfwyG5Z+VpgthpO6/zolM3LvTlL7/t17O9Js1Zrm5lqVRNTcdk74nU1VSdQ
09Mq/+QQdZi/w2LExBItH3Q4ASjxdat8OwwVRG9yxszTq8jy2L95DcVB1YpFwICv7h/+sJSHBxzu
hc/i/EItXXUclY5P6iQen2Znk1XIsSbRP1E86wcAadB9hRnRSlg8gDVTU9qUTP61gKzgWmSdMWHn
FY3t75YgqlEQROMS1cF8TMjwfFZDgOFYbltsMjxvsJCG8x0sI/VfXM87Tdk4hHE01J3hYVp1+pk6
gm/mAO79TR2RicN2D3Ufj+Tltf/KCqq/8IKrYjkIBdc1Gl0D93Lvm/qLWJerxztptT79xLUsNUin
T3b0fZyWAG2j161Cus+bQvD8tTMjUY09tLIHRfKlQ3BPYOw1V1TL+geG5byD6/5xlP3AxbJl+FGG
hddkH/XHAHKskBz/MGpNE8C75ugnkGKBPLO/jqLZVJmIwR6TQTxAlcyTSMXHX7eNVKM3MCdwgO6v
DKjGut2VKkXSW1/LBQZpVUKNWGwz9PS/EF6TqLAR0odHKGAbC3RGJnSpCZnwzK2Q9j8gEnte1FzV
1jpT676u30NyMYyQrMmysp7hnLMiCQpe3vGYrMgfnchGZ3UImu9htQSxV3QLIsJREYJdMHpsYqjN
hWs1Lr7+SOFXUvgsBYI22NwtRhi8wyY51S8sxnAjYfdpD1VjtUstqCZZxgMYDNOUiEWzeujMZ/fW
CAJIiSdHQYdxVTLNo2JJtFaP/BD8FsZ1zo4N4j8XQaGwUnmG9G1sGlZ8TrkrYlEXstC0DbYyynte
E00J0vBbkhlqIWmbjKVbbLN9VQJWbSzabP9ENnacDITIbH0GYMfqeIbE85sDKQwdYw/ydmry0oph
0FU4QTxwAo90myqEa2g3hAOEgfQL01CH0ivdIIVvHGrnOLmri6MbyeunoFrip4w4roYCkuimwg59
LAxsN9UFqoYCy+Sv0uDSKs/9KSvFrsGxHEGWdvrcCY14/TOTLWM0veU2uo+RjevwA7+aRTWy+x3o
NEkNz36+l/4fS/l1vbgw7Pu7kdkwH07+4prQob/8RMDk0chXQc/9a/IbVlN9kL1bC9ec3Fl8INcW
xPNyHSboS2U3TWfn81c/BidcEMt2y7x+wCKYuZsedpUYpDN6OrZybkya1UsYFDVUJ7CU4cBcReFe
MeKHLNW8tNy3VgNEq/tInn0LG7PoVBqOTaNb31A2WToD+VVdp6t4+vAyIeAdLuPrs+xvzii6gg2q
65s3z1DXUkOQgOLnLzN26W7P1aMO+9WhL0EHm8A1FP7fXBxMJ6YtW97FESuxO25Yd68BlIDgBF6f
tJHSUSagQaI8UKbLh+aj/eCfoNAqy35HYWyXDUrgmnKCinOhCSNzPlWpw0V7J3uL/NVVegO6piLq
mrIe0VLjcXehe3xYWD0nwWYoI9Jvn/vcKpnu6QuckjFH5DPwaHLSVm/BBnNzrtinVtmglPzrkik4
XE6zmc5rfGRd54eujwSiWYmjJiTd+LVwoZIoN/Q2/Wlel1HoHbS41gIe7uhzrEpECvB2k/RXJ1lP
zGEKV0FALDbammvfKp5N2Ku7NspJpS/CePBfhaTUz3k7ZgZ+Zl2CO7Xbw1gaJR0Aot963DWNqcG9
z1XxQF1UKrf5Bb0n+IZQUIXQURQv2LYjPAdfkr+9XElOBzGwiTNB4ZPX7tEMj0VkPpGrW4KEMSGa
QWbf4HWPW6OOM33E+/HeTyLwmky0Uk+/bWoxKRVv2P7bj5d2TSDX+PqmjRfRlTK3d8IVE9j5OtVr
IulKFB3GbxtjvxRyDyLP048AnGzLYXRN+sfTxcii4XSoBS3FvGvC/TVwf33MPKaEXYI44LJgfXNl
qeF9z2IyGLO/BkaabpyEKZgMLYl6QzwnDjOn9X33LZR2ZuSwJPNUkCJm7F28eMSJChNATircWaZL
uVh9ezdlXqpE0gwckLcRik4PXzld/rEEbjrGTMzkrMOpmIwwdn/BdYGkB6N9QOmtiHqTeT0tlrV6
TWRyjfa3Lqm3cenhxEvGHMbetoJxPh8bf9bV9tZYCiCCR/Ux6Ktjh2e9qS7QgTika5/hSOg3JJk0
lg1WJO8yzxyorPKxmwx72+aN0Xl9R3Eagb1UvWl49N0fCVTDTcn/OkaHxC+x2Fnuxy+LIOJqZEYv
SsYI4BXR3ZngS04N6z72nkuh6llEKadtgmMoriz9Xq8a5WD7w/TLwpFagT2oJlJ4+yfPMcw02plN
c9Uhgq2+sDc1n9FNBLCPlsC0Wv+NMUT0b5UTHdFs7G1n6XAxdfVkui14mLSI4LmGGnQJmY84/j3U
vrB40UBs9WCJqL/3VksDuNm+IcqgeGiiJVRknj5aQzEdUv79UvDrIX317cDVZOBMsHWH7yhmE/1G
SzPgNujblmGEmmhnNyDj8/hRGynYOQVnyyM1CPqB5IM/M9n6wOPegmqZMitXL90u90qFs+6+uBre
jWxmydPiCfIbIz5ECZtatExtdBmzeOmIdXYpnzHuo4OhjL/Cn7c2Oc5tj8h2r01Wmy7tGdq88oIP
Adf3Qvn5kRZ6lrp4WU+bD5QhJvvqzM3bnX6tK2RxKNPCi4wfKmyJ2ekq7KGBaq90Fl6v+LiyoGEq
GRDzJ3TYdjZeZIyGoIG/B9blXIWSh+9WWYlhEzGORcpoi4ODUmOBLry5+NGQpQ7KHQNTJ9ltmHrF
qBbW5JczLKlKOcwM3PjjZsjxYigqCgppg5HxVNQYqsNLPusaRrPxO8jNSGgUuE2Y0J2BEelDSN1e
9LL3dreBeso/nv9BbLNUmW0EYRrnd5zQr8xk/e0V3nQNbNRSXWd5v+7y+kOblccM7O27wajpHJQ+
VLDp8sX2AWqxvSNdCWxNg9oZ/6d0eVAqCOA212ocF22pY3ZmT4zcqiHjxs7vPPmkFEl5Er4wyE8K
LCI2sQBE9tKDEZ/FYIZxPJUlLQyKAa8mowyVedgxDqgWgcTTQnpUsYpgN6u/KgPPNkVHX9jRxRKO
s0x2ca1tG55NHKfbyQjPecNYkpt4l7imIrMTC5dZPbDXhoofbebkWfnw+a81BMc7JtFbV1mdmsvT
dWFNhA1LA2ZX60eL/6FeBF6R7dUlxZd9+640g2DORQnmaBCua1liZMaG7E573/A24I5HsgwqDr7k
6tY49mLSGlXtourC3d437E+tA6aIYHN2oGpOJS+7bncfR3SJpGTSgEQLShWNloszu/CXziYSwHwH
Et9U8kMXLkuSduPgb/T1Wk1NK2/tjOxIyNl38Kee0MXwaVEwMRA2Z1a0TY/NhvyyGk5i4z6smEFg
Wau5KvC0VkCCZxj7qRaW+U1ju6kiEZReUIuGy1VcoLxzIL/C316Dybp3QAHmRiX27TRyHmABusvZ
e7NelbIuKM/P/Lltn5FAiQyJaPLMcYb+w4WqHQy09sYWZ4tOV6/zBY8UDsUIcOSEQFq1/UGcpPOf
g+HNYDw8k8/LoAkln/OwWYOex5F0MSkWNt8ZyPcMCN4cjFw/lpjL/qf1FUuH30Zw+TOU5IECz9pN
Ei1lqtObGzptwjCVCz+6NQjs41GBrHtYbXnCWHnq5mLpSYqD6/L3uC6g/7bTt4f3Xl6+5tI0jX2n
CkESmJvJAveB3ai+AL89QyosXGhv3uRkGGUk9rgRKzuChIXabSvv3o52fePicoOV95h96COPnPoI
auIJ762/QUNdXJmoDsVNg5WTr9omyiqTjMHVU+qOqNp5GyG3LMh3gdIyig9qezEn/odIJNJgKpto
2weYfsK5knvpZtLvCKIJp9vJegGMQF+woj5RLAsZupafCD9qd9b0S0s4LSFUEuL87eOjuAEf8hA3
jc8TCFXL8VndU+pjaS0T4VY/a68bmQbH7NnJA04yZoiGAxpvXCPQFaNePvEtOSWH+25xTjMGVYcO
Q2+28gO5Do3lkwRVZEl5NbAG/qbgXx8qtzZahPvxGlWRUuAOkcYoPQVAtaHvX0cdkum+eT/YlUjw
Au8IGHI0acDtsfKeaZM4wdpk9ktT3gNuIIkxskXi+zz2wD5ZihZNePPrC942/Gh1j+5dlIeLKSjM
/11b7XlDqUbieyMJXXEQ/Mdy7NoyyI9K/IdoxJ+Dj+JYc2GPvw2OJqutvLG8Mk3Zg8JyYywVPRlu
8ScdZeFPDNOnh+pahQnsFw7YYDimANpHL+oi6b0aMyGGywuc6NJD1corilwvKbZdVJawDKLq6tIc
mrV9Ar2sbfXQdgCrBix2K9TtRczOV0cGNdXVafwINaHgkEAno89FhmCFw+InGbgabiTpyTewAls8
GH+alXCyXh+2doc9fzI3XGeD4LmkXyedO5oMB1rvLpYkwRtLGOdt0MbqOB76kDc1r/0Tbw2uYqRH
t1wKu3lgcbQM8yutj5NadSgCexJSxYCn4SRTerDtrlOH6oJyzsEf3sg8AGHXaultCGfLKvYHVQeA
yly+KqMbbX0iebIRjr1nuv+eP6jEqcnLl7JGIlR7NUHSdHVKanTRXH0W8mDsTHNZusLGYQM1RLtn
nOBFDfHOeYHCpEfywCBTwDKNz6Gtnn8ovMLK+uJzX7b0whr8vMKKnnFVOK62UWsFJi9uCtFQS1KR
ifGgwN3xymGmtTw5z662XnYJTmWMhtyknHni4GzBD5L43RuvXwfdwThofllP8s+hgl3aMYpd8Zfo
NYmAqRVxFgk72ZOzGsYV35kGGImbN86zIKZKccWxydJAcevbCGxWPD9i4zIGeABrr3U57A21MUza
PQbyDX61eETBffnELFO2wp1VMw+noTZ6e9/qdZPc27qe/YVQ1B3bon5Y5vLzzExams+vrZHOZp7o
OHwYUjEBDeLbNs9Ccv/sDQy5nODWBaZW7+AjCR2q9/ERXgDBAoVPbtLWndWcwJHfC718dEEFN+bX
wTeICOKhd23v4RVH6hZBGfDPYZMXs4B28K3uZKioFjv8BhGe2c83ry3qswvTmbcHEr/xxCBMFMXl
zhhFISE6pBvu1LnzUYz2fPLC8O9XyfB6vcbFLr9I2i+o3lA/b7tqgSrPfrrhsRhMD0VManbD1sAA
ynrn0+yxEfTE8gfdKHki732C9lzISGHOLSbeTt8aYl2f9Mt851jbrvJPZjqGjNtCXSMx27yDKdG8
k+d9Yrani/oyMHRFL+YFR4a8Pd2mDOH2zxcKivNHCZeAhcFFj9BeQ/WXyS7vIP2KS/no6LVLLDyx
zz9GYVIsnfueL4bGR+HxfmgPgB68HfU97Fk54Zmddc9O0k4OQcs4tP7u5fzAno3i6FBOIvnMUByf
THYrRxvwxqA+tYooKOeXhv6yo7aIEYjwlaAwKUMKej/jm7u+YOkuMQTeRgmq+ysDljelFCeYEGKZ
yJeEgAlOYjf2QYUTGgiD2KU0g/52AqWmWDbvKNUpahjzjXHF/c7wzX7Bu3vOMz3rSbnYIW9/laab
+xRAymVWOF6P3jSTK25Pi7ni1Ef4EXnfTM1pRoKa/Hssb+9OiUZvZi69ckG/qzZWomAn4nMEOV/M
qPn71MAUPM+SUaVcvlH0v6QZrZbM64jBy9/dEJMEORpfF0Ssm250PmnyyDgut4kCVKkIRyR9j8DL
epoOJ+dWuiZ2dr6+A+Yk2iX1F14R5lyUrbnDnjGDCJyRMpPouTlUQQfXLrYZFH/IegRwOVKQaJPP
GSAm2/l/PjVIZoRd9zvzW0stGM8AscdHQdU38E49Vq4NwSkcFLXclHLnuvlg02lFFlCOYFV/KtOX
cRtjiHpSNnF/XPUV+U0DYXZ5kMpAHSgKKYesmI8xEwM0zCmjSg1/fQIUmFHCCJf6X8JUV4OdIHEY
iHRo4G24Sr6P1TUyAGeWw1YXebWo+AqbiTL+lzjg+lnD/S/qMXlOi0swf3GkEaTf7drG9IdNdEKI
JYxXCamvzF+esu0IxTJmDlN+RJKtwLN9DqRkoji0KBu/UJSMOD0mlzF6loe6pO8LJWEFR0e81gi/
1nozV4B1dod+vmwwnT/eeTnvfbEQjkeklH3JitXcv7cH2BweyaaWTv2DeD9927AOAqEZxq5RGgw2
8g1c2mhDOi5cVQZ+oX75oAmOoInS0SkOBZq/TfAKv9VWA/KO86zI5l7Abt/2KCl5FPgcmJh/m1so
Q5/hii5MlgYAdaOVmOV7UcQnA1cgFFRByjcsNoaiF1PFDk3N/mWGQGDKgDVHqQ/Yrvhhriln7cvD
LrEKY4LkLopyV5W8uJtmC4v0on/W663oifzjTAdPnVtcLpyBuzW68Mf2oGw8OQoqhtQdp01ehNyc
0zZWzNqoWhhl2xllUPUe3kh+MXXNSxpNlCMn2klYKOVt4tPgCTNtsVfhekeQZ7bg1RxibGYXs+hg
jix1oIL4HjPfbLfGB6IBP/ohLR+8A2tcqMcgiPuQpN8MPK3iCwAyD7LOuG9ZP7ha1xROMNaHQxMB
+vcbkkHaJdo4nVIjcpSkeow37IPVgd7l8nK2qPKkcwVnM2I7v4L7ndM52GhB+gbbhdRTJGHdAL9c
yti90mOKBT55eM/XgxuWb2bYdxKwrHznpFG7mupuvMlKqLcSwJr93clWtpv8Q1BMItaMKkuwuN1q
cZG9b+kYcRYG6cz7IjiA5ZqLijaH9EmWYPhBWRZlnBMoLFXaNXTNSxMg3MMRUV+xxELR3BwAIazg
vA2vhLS8dp8J6yJqJvG7v9/SoRYvqh9wGeksVEaa284/dze0AqQlmAHccpWkfIRZTXQL4cRyqlyC
GIjpFdrsWwkHdJr2pWzSFPxzeQmJ/Ey5LI6UaahsGPjCLFMH7xiVyRbubdrGq3OFRhhle1hibJ0t
d8b1ykaV1O/UT9/ReoS0ylW4lvYCP3DQgrtxQX8nYY0rJtGDM+jaXWbnm5SfsIG9C8kdhEkKpYHa
K8pfYXAyNZDzvhOm6uI0cLciyPmWorL9czBo4qCokbEIGRUlBMFREeAGzV41FMotoRfjYzd3FWt6
iYapOkgWfACdWij+3cNmp14st/v0YpFSw6NQlCQDC70Vkb9JH735ulKT1Ibl5VzLaQu6L396tsaH
DIS/R6KQwKcJj69wQv72Jb6oTi+gXnJCVwVqAR4sLfwgDfZTC9n+1cCQAnQVXgWwYvaBp3AQG66c
3HLp+2js2EMKLI8bVBQ0Tw2gkwvvVlDRPZyS4/LCvF82MHq1uFEV4v41QF0b//8lmljH2Fve5Z2E
voTZZ3IKXcLH7Zqle3CXLKKrHlWOpAGJKg39/SZDWz6Gf0uu6vMY2aQYA3FKB1SENgkTvJcTVcV2
IxNj7vVQ7yF+go2cyFQ2RTBoMHPQlS50n/CWgtPwDLoDx8pUW6D0AP5/2PO8P86+4KxjBx/Q37N4
l+TfeSQvVU7LLAwz6odCHufM+bmcJUWXKcCt0xjBAkn1cgzdgoJ0e0TeQzO0qRYbcOYiAd5lgKrp
kb76Ygnck870ckfrVSz33X3oawlOnyVvO/WYXXSNicN6mImq7cjg4KlHgC8QTFE4nfOrKubXF/sQ
/RowlsGjhR71ZoaMxp/Yu1WtPi/Pf/FAExOrvVkpa5EjP1lUXLOWi4p5s8rsusL10s9yNXz/8WWT
GfkbJrvbf2CJlzvKPd7rtF2SMb3ryQMm807ukpGQM0IqitgWIYtJyoeaXRijWsF0blcACrpL/FnZ
YKO3+ppIfS7OVTNK15cwXOGAx6LOqM3Q/J9E3VmdhjSUQ+ABUavPYjzmcG23Dj2QX82P9oaQ3KYB
dGgSz/pwad6CwYgi7fTC/zYH6OvGIYCwaqBA9vhgQbzUdyNQq4XCuZeJ19/aXjWNaVIRoCcOJwhW
e8Ex4nRsMmL5y2OjFYmvQ7emz3lDYdr8pMzS4RSlsVFcYHP8zNpvyxAJzo1HV43ob0Ocyh66MtGy
frubtfqyckdNk+EGQPEyX9t8l9oWVg/Y4CCEohjBQ0IRdEy/ccck+JI+bB9WrhprqN6lKCrJTY6v
ADr7Ra9eBFkPw0j+Ps4n/TIEPY6txGnA4kPl4PqJTtMPBa5JFU25ToRbphXBDyWdDawsh/W1jf1B
+v4B46w0VpelM/xEmmBg5HN4t7F8zpDjjK+tV3OvMDmD5PF2tDR9EJ8Ufn8sWV/ST3lxNwG3rXgo
ksCuvWXNJNyWMoSEoe0vFfHJe40zcuKUx/7kpMVP3Eh9cKQ4/25gkIz4pCdhaijn8jHc1jtDPuBE
gYLP3KPcKRolAR9Yoecf4JojxLISMtd2QlwdRmtG+7jkJvGZI/nZ92Dk9I50xOO/jDUJbmQP+ru1
efvjcyaykK6sTKk/sHPn2HEGjeDDRgvNxFxAWJ0jB9T1YUQk9yj7j4qGrmsOUC5g72xDFSDnX4ke
nHgIfcOjnBXMem9iZIkNY8G7K6pa7xC4BTaXDgeCbYstFR5b/3YEVVeymYq3VfHHnhsAns73kXvH
LpqroChw/eOiXB33qEgvLrPVpmX/CBjeggtATcLxSwyknqOu2Q32h5lDfgNzYOsZv+dyiDJEUoae
xcliLXifij4jG87jdFLkwIpyduG3MGE68bsg7O9nXOaOxQhFT/SE2DRjqtpSmtZ8aFcb6X5AiTlY
xW6ijsh5NDC5dlAKyC+SyWeLeAaedgSTlHNbdguvvwOek+WLA4eqU37KNuWCObvjq2/jsaofbQRf
GdhBBQx53XFhiSRRAAuBYlHmnFbsFOTn17cJyhrMlFtwiG/hQl29q5kSpGnyS9Lq6clmmGDeIsYk
Vnn3ITE4VCqEW0C15ECdBUkNpVOQFm6/KXS0c5kWwrYn26tsLA039nVlfsYNG+RSXyCLspnVSScB
aw8jh0s9ro/bXe5jF6v5u816/JFU9gqS3ar2uKeNJdq2hZd6qAawvo3sAXcDmfCHm91gC3RQS+yQ
RJKyePbu63JPYyMOV+wntsVW0NQn/UkImKLN0rZpMpHhi/xaWb3FQL5InsD/UP5AM0YSKIl8dyxk
AX58Mbg4glaoz94VB26Id365392skdi/0VQTcnleULaQ+oCgevdEbfQJgOX3w9rXasRgAtY01ITA
a+Q8abJQQTP7rP7ihL24DJFKJczvnrRvBcwGqa85CUrAXkTRJeDHKqDvDLFykP+CuMEBURIa+sd7
BYu2t99eMikrwWsIfJx0vHa3tk8X/xKfxvjx2tVMhSl0szgkYLmWomjPjsCRr0UxWs08LbI0sbR4
RZxzilOoN30PigwxixF+izsmdmdc2k3qaZ5CgcDWhl3FU5DWo9cf0UKmizJEFWr3z6DIXLx3iWVv
mH9QblhxQRdEQjQpOmzkr6ywcY3IW2dA35Pluq874GyHnIyhZKilQIkbw2vuaY0lA26NF15HhgNz
ZdjvTamWmSLIBaBuuIAWImm1uxqco9ffCtxRbEAEkBfbaFk6RcWX4wc3vpnxsX8Tgil0LJQ8YAKP
P3YO04uCGqPWOsL1HACxFNyDMVx4c+776QgPSonnXGkyuQLMqJTeYTf/KzEDGh/zbvYrMUtQDGY3
VYcEL0Kem5/4MoO/PhfpVmtDOKAK4XmIWN/Us6lWPWXmqrv7EioS9hRAmXE0XLVYrIGg19OjjRjV
icSFSbbno0WNl5dBJZIAq0aKkpve8/UraXqzkPHI2tb/QkDrb46PsuusV71yzcsZSouVSFLJEycy
bK2zMiHvxD99UHcsd3kgmr/tpn/4ed9yWU97wU+DdadViVUM0bZMHTftUDtPZhVno2ERI4zca3LR
advGK8zX4pyOJnNcUkh5XgRywTkeCvba9zTybzaT3rt25chrDmROEDk3l2N5I1pDgKbvgQ+oUSNH
k1VEj/4oiUFynnf7xRxVY5Eptcx6qq4Tm4S1N4gevtOfTarfp+0ealBkdZXi2w8i/pn3pvx0zYob
OxsAvcCtaIzijhwHIPaadALttblCZfOqJb+twREcZSpbuc0saswCDt6JsGBn7LpCWYBz0hIdSaw1
q93KCg4WJyC7s0QAihKtevUKX/lUszP5fDaUhBF+SbcfDs+I7JBUixltnoWBMTsubixsEdtDlFLH
nTqYkwTFPssEo+8iNoAIIucvKDf0qR5Mekgr/bkN4bi4YBKpe87+xgmQH8wChEi+IzGHpXuswY6z
gqH3doYp3eKsVtJBvgkl17SsI5voa+Co8ex8VYW9/srVgwJKbmNZfzx3wOIR7KfEQFeKDmQJWREt
2Imyx1KV2e7znPDPADI7J7IbsJeDr1srxS+uISuoC/8fbSGCV1xgk+YFEQmj0HQT7ZwFLqaAjCeA
xmz9QygqfUXUYRuDe3zLvotW37EQPWCrfKRNpC9cmrcteIl8Y2mOaUvWwp0B0R7Ynz7SQE7S/C5F
soi1kbJFFQHI/7gGpJ8HiSocPp4Ry3Luo9URZNImXLRVCiQym0opYxTH5B4/OstKoFGvlTSg7RKA
FV+p2Mb1IQNv9Tt04CtruPNXg5WYJXalJ6LOHP+UWl0LFkh8yRjtLB8ih3EcdJ/IF4/iSbNxmMEw
wcGdU60iSojpzYuT2WeDdV/cx6PPBIGZ9Vfpd5/Kuh3nYy6Lzyev5NbhmoRK03NuaGJ2YfsJ9I+F
NAyPSB7f1sLBnUszbZ8JBN4zzoEwd0npHkzo1sNm9hdeF66arKz0uNr95VGpX8LZ1R2RWSwcPdXV
2+UgVEj/MAnoyZpeNhwYrz5OiRNpyYgXkc1yAmaA4J01WOnefg2rtycAzDEomJrYBYT9QF1ZVtEg
PSxcz3qFFZgIdI9tXU8YDGrcgQMp3aKEzS0w3n57f0ObzUHctJwFPHNH+c7B6oANHltQZK0gQIeD
kOXmApPHMNOT8UcVIAT5gbobP9UuF+MiWIsoCtfLwZ2l77wueTtxROGTboTh/6Qmka+DGlU7YeMc
WDVaasIj+BSqGMgMEZDcG0jr60msAY5TLpJAq35/i/C02XLJXg5NILgrP+0nQ1nonJfG7pXN9j/1
NUWWjnxXY5QDQjLYJ0DbvBo8PG7DGXkuuSxGgJz6F7GGrE4mfUEa4ob0WtbkaHqX3GGAfuWkC/1R
pTWYf2tWx++B9qssQagF737q2UsEjMfC/yPRCO1lyt5z31v2Qc8Bf28tROnV/WqqbhP5AQu+DGTk
tddBKNwuUA6zk4DxQne6Mtkfb/KA3RsPLvmqn9Pm1fxxjvwdAiTqFQzj4MVHoN16an87x52X6MpJ
kolmcNGYgkKVsr4wn8k75AqGqf9SwgeVVYKeaHTEQPBaEtsdzKBGB53WIFocZsyXfo871JTqPVW0
pp0uBJW16KP7aFQRlNLBSZaSLDGpMiG/tLEM5A2kW/6MEYQLxMrQ1ihuD3NYokjtUPNPaBX1zpxA
rTMWyVMJP5AFNrhO/aK3YFQl8Mqd42pavvgWGpYdXAhwfja6CKL0Xy+y1/xoOvdYPfhom08bh0DB
fcw/K7uNcpEmmFUwrnD6GRZwKxSZqQ9avSD00I+12wI2OKIQrvLfHkXzoWIDudVEz/h/Zjxkm4+W
p2/fUfueOgPjpdHkely5m5GiyiOpmtz4npxu8OIYH91nHJ/olcGjkz/gt7TcTeOhfZ5BLI3iBHNV
DP+RRH8ZWLHJcF/tSySsYWSmYUm3HwjAHBKyQnOkQPT+mID2Nj5oDjLXtJFOilujTmrhZ6IgFfCQ
twK957k0GOpx0tK/ML9qHcu5+UoydLBxXfqAs7V3dccVDYIqftRtMQKUY/i87lI8VObEnZcpcFp+
NPEQMLfST1MEFlDU7CLn934UiMlFdgrOgXrnAzLNaOEe9KWjcgtE4ckngt8/HpYhwSQPg07Bi2uK
+fZFRHnY2o71gvaKz2/3nwxZDqLXbUstGwwGtfOrR5KtSkOQXY759ALOe53GiV569rJEZsyv4aer
PmvgUQSgugZ1F/QoTcUECQkBAv6GQaDFglP0aM1BFfpjQgH8pU1P5Dzi+moy9rCHSITX+4O1taPQ
zxPaU1jGeM4b2kCDfEbhDW5i84EcYpRLQmshT1JLjXt5MlAIulJ/M9kcwbTzE26zaADxjkchaJdH
h+z+U66lA9DqWkFB2ul2U5Mv566w7Bxw51dhV/3zndp4u+axP3OeyxVSuYhb31ODZ4mhrnRfqHMV
I6FpgEcDnP5MbgrjdzcTHCIm3KnTMIcaCMR1EsI8YBLq39j2sPF7T6I65CA4kha0Akon652xzWME
v4nLfL6fwHWwA/CKDzn6O9Kp5oyc4Nu+eoPfdXhLQchgc28H1V93Zymi8KHfAu/30PPWVVUki61h
VtmoYg+GMu54XfmWhKgn+PG02HY/+31fgpbIK+ZyiK2S9oZO/OxuAjAKuzsypY6gDkSqw4d7kTvE
MKq89rZJfIv2/u8Xta/r/CYsKzRtIb04b1uM7+FbBGMN8w8zOW0m/YcNXValJjyF6KK+ClTm+Vla
pOzT82w77RM5hRgjf4tsmgtPRhTGE3Uw3SBQBurTmbElXUrw/Af39OgLhvLl72ZL5NxaD+bGdFX4
MVRNgzJtV4rktsPQ1KTlvqvJzagzAyfh236+mSWMlJR+hBWWNDVR6pnHmG9MGH9mI64+hqswVt//
stfP04aVMJvb1maXTE4Ol42xrG+LXIlCN3cEue0Z6+Qkq4KZNpHnGoFizYCOsklSvQAGVjlDkNVe
sPoS/7unVlxYOJSw+CQ3NSiDlmwJyNGcm6Vq4okRO9px6TbSGHD3XRLVIWq8m1PLatQPXAasGNRu
dF6hdPmL7UIv6B9MscFh9Ksbrh42tQfIihEDcDJWFxVpi4LAdg2V5jpHkJxvMw4Rh9tU1w99qZoa
eReJKglE7XFJWybLJ98EhA1N29RUeFqqagOMr+kEuoCxjsNvXuZ0D76EYHoqJeP82zCT62oxnPbU
lGUrHlHPZv4tllLVesohpHXrBfkSq3VR2B6Xju2MondLi6edSvfw44eI1HmGV31uEiNgLQewq0jg
ywD9yrf9G7lwkxzqYFSURCu1fBY+yl+1ewsvjBFcrRWCryesvnX/EEn+c07QW7OCjRUelAERl5Vd
sQ+av5qvIVN7mXfI65OxIp6zLW8FNp+DkXRM1k78MjI1DQp7g49NBl5c1v4QXQ9Cya+m0NsZbYZ0
cSy3jXV5LmntGFH9Ktt8A3EPtU6tdCnTw+4nL1XZxMclcaeqgBheWBXsMIFQCHSXr6g4UBhqHMe/
x59NO8n1x2UVcvE3t7+Dfxjr/h4Ty5/ga2LXyf1oU1DELcxxq3VMF3p0EpE8Q2IqEw/bRWyFBaku
Rbsh8LIWy7Zr70nVzneVJSqIGkI7F9vpimxXPghWi0JhTL3XlmNdRxCwxT9S6COzT3pY9zL4Adit
5fjx6AIu4dCOHxMhiCjPEvjyQGEpbMz/Im8pxgZNqWWzj6+JvBpowGj1gG8+/eOt81ER4oWTOdIe
XUgeL5IR2GNFi3Z0AKRQv7bCvN4G7y/PR32M+V9QCV6WyTgXHFRFTHVi/p2ekTN1RRBgLVKj040+
dDTRRVXoPZyKlh73cewSe/kECccGVLJhpIMGWaO8ywG42hGFp2R9lmu5RogUBPLtPOtd61zcHQME
VRltEfISu3hzCfNX5pMo+RONFzSkIOuhcLg35RnfTAXtEs0LnloV7r5VfV7itZV4tDcr7JIx6/HF
aHQA8PhbbyusjVpBFtHfNKwr5kIzh7MNLWgvu8j12m0+7lFQRz90X2M36s8C50C9EKy7i2CgwIWB
9aTqRPNeRxDyIsHc7xAPv31cqA8in5KAApekMysuz9Ft79onAy4GHgV0u7ZaoAdSs2QJd7aj5akw
a/oyNFVcJS2KFVNWuy1bts8A8owiGZTqo/maba1mjcgP8EL0HeeEg5ydwhutyeKfwsopQqAcI4Ma
7LTjHrr2P2+FkFboGP/p4VfeBM9yUKgIVtI98thcFAIS6lOXQzfLh6w8NXF+42oa/CIH1U28oFFo
lMlMRc1EH2r+u/bY7klLPy3obQsilNRR1GU8LD8/G2fE/fjODn7R7d2nCTQB70Bn/ImsewLzw6Lr
3bVW02H4NV8bdwKo5Ge32UPUtotGIuYT6OmN3c4cCVken05llJL5mgftIEyuqc8ErPmNIQl25prc
ihD+i4x+CDHQshQsfD+NhIr7Lq8R563sEFHr9lGk+vtcrGwM1lu9IIUYTP5Mmf9us9/PJVUbIaKX
LbF5rsM4keyr8i/s1/VAo2eJsid8E/iY47BRDx6BbemuAOx/BWv7TEPcr9zdrJpOaUcJDlVfCcLR
2CqSoV9liI2X/IlTGbsAP0H87OMicu6Qa0BZtIGbavMb4751+i9Jo9TEPVpqA+l4vTniOvaHb1TZ
g1NZ/zQW+3UsFqDESwMmK6QBBjM0bX0XcmhOw/nyGVUUlwf/CqbQm/K7FZ1K0ToRZIo+Me9D4v20
t48RlTGiYsAMYUY7SiLtksRli+olof/lY81CU3BB3Uu4JPB1nqsbIRKxWjFcGvt22rjqNQUOjxnp
UAMX9ale4lZ1FJj9p/E5gGWaFglUDcLEdU6AtuuNC99aSK7qotLXaAvBqvt7P6Bd5fUG1qeMyoDb
P1fQ6ki+lmGO0T+DzEvt4Gfi5keO2HF9I0VEk3eie/T2Cd4z13j1Zw2rKdUu5sSTIYoIZrtf9Rzd
NOLJy+VFy/r+OwX8Z0+W8GWYu2e5VDwhQHdI4w38b4Lrt89BhvMat/GKu0JW5HTGq3WF/rqFL4KV
j2kKLH/OT51+LnYam5LIfGge5F8nFhTIzxxTuAKGb91K7qXsDx/esComO/Tiy2lLwIjDcsXlRXKo
Syx8S6NdVTzHwGwMfKFC5V0bNNOGvpIa+uDp+4TIj2YBjq2NP/iRDGJLxXf/K+1lOHri/woa0LPW
+SQ6y4BpEEHA6nIW5y8PU1ogHi0RpFDSPv3ql3ldf4RR9Q30EVmdwdopwOsIbSa1XIXp/GQU11qx
IN/FA9PP8XbIh5MHcRWav5fqdcVn4qi4O9q/ZwMjksn+vrt29LtGuDOuhBlm702A4eWSS8bC91Ho
S9jrTIqTqJIMIwV0E5ZZfUV2XBRQPNQpYITZBAZF2/VHmgw/CWPy+rvAQBPEKkr4UD1+oymgFUMz
i/7fEwRaXVJB72Nrtu1aI3Gwt+gQ5RvDrs6RY76s4r/0xYaJQsj7pwnpZbvGgQz5AG4rLiAQ9ASC
FBHJXhfc+DJrnCXRuD6HKPZncNtKZLdXwA0oKB+2tEObgXdRsXQnF2mtE1VuthNW7mA2LwXNBclM
FIlM4F45ldtnAXVopsc/WqJYgalqhYG12IpGqkBSRgCOBjf/Jy/xJT92g2xL+R3atCj6zfoft3OG
urfBjzDt/VlOzT6bh0SJWVvJlbcKqJ9pnM8uURmXAqSpEdMczM/lBeVBLzPMC9YEEN/5aYmWXYgh
STuJioqULIMFIcPxGb0yCXerWPaoKVyVCtfefhIk5SUh7bUODQ8ZrRugrUodcKsvrHbCREp+KcGs
k1QJTzyO4faItidSAdFDZUTX31Up3q6M62hjqKpuR4lrsznJiNoZE/ixi9NINRxmXn+j7KSMvRun
TDbgZKCQWSOsprhh+yBQQ9/NCOJZgBi46W3loCkvazuT0Ps4XAPAJxwIEuFkCQivmsnfa+zVh7eI
iHYn3pans7R70C0JXJ6U1FA+JPv7tdq3ApRc5tskZN1twd+zyF2uqqE/ARuu43immLz7rLhMRHly
qgW7P/UWmgbhVAR5VgDOsQtNBtpzdVPEBICd+hB9AsaY/ELGsQMXupLOC4P7rq4P4DZ5AF29rkQW
HfZIpVdSsIW9aw5V85WC2Frn2WaZ0C6R3+qPyMGm43gENQR0QsGTNDm5yaKHYqTa59P8fy+0UI0u
kL0xiUqeWtcB0lpmlu99bgxJ6AiTu7l+wk0ihrkQph3JwcavDzMezzc10fXKONSXxjBcvQlt68U4
zqdTjQxFuFicrOK4OOX7JyWz27Zx8PuJ+RnDRvogEjMqaeZDLHV2i0W3E12u9IyElZAxshiLvYIF
J6H3Bp1UNqzUze1KLDfk0wW3/MRN7r1yBeYOYjXeLFwV6cnCtqEQ+jE46BpgNaKcSvd5N+R0amsG
6fmPGmwy9zejiIF38YV0vrEjbJwy3aV2KVGxOgl+VxJ6xJJB57XtvOh6zmsR+Ybr3Zhxro2zjLYX
uHwYv+9AKliehm4u1pgFeg7iqVaUyVQZTiEJBGdfgxfRODXoRK+kwOf4+vhyW3t7cUuYcGbnLP1G
wcMEJtlIz8mdfo3QBWznXlRCIsDPhw2x6vWHQZu4cSWQY+ipSixmqh9EqDTJb0UB4iX/Sxf8EvpB
B7fKZGkDGcWrt2KHj9Lbhsqtu+B8NfL5Fw/8PEiSxRXwolp5u3NOcdJbubhV9LUHevnYKpATyrjj
FlFKCoR1ZzgLclHf5/rSHAaxMXet2McX6WGWxP/lrIe9xfOdC/rLtL3OnoomC82820NCnBUQ4386
3g/IEgWh/vPAupiXsWx61fow/eXn6JL7a+xWDSpWSXEAAo7GPd1fnC2l9EeuRU3bawD4sK0+WsyU
b8j6MdXbVzSseBd12ai4+Ef0MO6ih7vMZINR3J7GxBCrjovb8BX1FLOtoALaMqTJa/jukNARE5Vm
7Vxp5M211R5ozFFydbPC2CLZL9UgxgovhFZyJyf7XESIo6jP25MiyVRvSxCH47zD022KZ3e7mUDl
mNj6D7uSvUfm+bCxDSrLgswnVmpe2es50MyfGRBawM+c+LttJidqYLi2dI50aBV+nK6coweXzj1r
3kVFSBMhI+7ddw0zeSgMGYTR1l47qqSFMlqUY9e47e8PgEghROg4Q5eHznix69uGbxCtLS+0DJyr
ZGij5Zlyg8INV5Xtr9lXWfYClzUxjMylsTnCmmjQmUUowm6IRJY+6aP7wmH/zojA+2MCfqdujIMn
iVWiFfIpBgC4QCc8hyO79D4p5YskV0Uk+bUVc//zUOg1qIyEE3pAREGGBk5QMFRKrYY/bczpz7Nl
b25xbKMjQKpui6VSUiaYuPIw/Y78nTuIcqtj0ROsaCdegU6blOeR8EtdJh64ZPblTEDvuen04QB0
N6jCZM2Napxg1nspKS6rrZPPKH29rdaE5SCCFsFTkwmn+T8PweEzA+JqIDtZKnNlGrSl6CaEiED0
F0Pc1nC5cEUuonVBrlNUeZ+NjhrKJypMpApMgbKr2CZQBI2x2OKRALOgL4joTEouQqdr7q+8GTUW
ReMDFj76Y9tmy1Bx36g3ZQ0GWM+9ycZHtWwqQFMR4wjGMzMsXGRygwEJqNIv+HjzFpyPFhJ0SUgT
PVCh2iWwPlTBCjBNLxbibnZEPH0MN/gHtusqDkjtrI6LgUZ9N+OLClAzNBhEQhEYZwDeTYJplh1I
mb8e3xuFhFsibaPCH0Tbv1SR7zPGtOsophii3nzWziE9hPJ3jmwhoOQw6l6pnA/v8iY748hCpPiO
FohX4ECD+Z/3CzizJLwBQ+/DPMuGoq0RNb0xsKAV7mSZDgkuyWr2Nd/EXXSwTyNUn+clN6unxKlh
o01Zqv9Rm0Utac9fTadoMQL+ze9XVGpx3cMgWwauPxVH7fbNDCQhkb1YNLJnYwzrH8SEftksKj6j
LWmOMYa/Kv2FZ/8Mi/2g0mQVBrfzXxc4u2XadS2MLBeK9a8HFsnlVfyQ4znTU7DJz1rCyzN9Ra8V
Jhq67KfFxuNJDcNpN7v9uqZjMbZ/X1woEaZ9uPYEJCvtJbmTShHZXOmLUTq0J6dccow7VfGUSPyC
T8CGrdwVVlIYxlXdKvyAu9LhgKZqTOW7qnENL+BMIczCg2mwgwmSUyM8FO8C9+bGNGeprANBTOWN
57VTs7KV0PMglzkpPNWXCUITb3jsS9vnCuNx27o3lCM+FeVHl/5yBsL9qanKkPB+kkEzAiiKYwvx
y2Yk/Eo3BbjrPjdb98VqYqdX0gggIZuEFQvHFVh7/MYNF3kEyzdV45I8PRJ5g6ISGD6oGWazUUAR
ItPy7FPkys6RPS5T3fD4zOlXnHDF2Ka2ne2Bxx73lhF9DG9YcQm9vTmwsn//VinESBWRFc1ls9Td
LlLMyuwsBelJN9bdmCL1Y2svXU75ru3kN95iWAs/jOx0s4o1E/s/0ylKbHE4uh8P4mJTS/tgd8+b
IXi8kqdKD6jUMF3LREzSv+zdh/sEZ1KiRU0g4Rd58pUVWp8uRcEHYTfMzxCtQuIKZKz4Z/IMg7jI
ziIhQKn3aMMYp2Mjy/h921/KymYm+OUwcHObx3PauS17nWvocDO2OVvXGRMw/YDX4Ik+iT5RDBL1
dNlGCMsADh0gN77LNpLjQ99WkwACy7JDfGxYB+EdHi2CtMbyVklTutKEHAZSqcclZePfhQLubmJB
vtZMxVYYwUmrIYIQjwa8SY8W0Oevu90GpAU54x5Pud9p9FyZhX3W9ZBj/w4K0s4dG2qawMKOzSj/
kMJTLalO6Qevy75gq4j+O4Ngs3yA+MnbntxkV2iGeK7dMfCa8dOpgShhveHRq5LO+Bm2G8itDen9
Ni95PVLhfgSgL5rUH/f1tIjyK/SR1uQMppp4FLcAMApXC9BOLnzyC3ieFlUOv7bHgbORKwcKQHIR
wGCog2TkF1h09LZxW3nSLVslGbV8s8BU3tW0R5MUI53sLr500uwS8EdLuXyh5IJ5SMSitpYx0sKM
1UOp8ZApPH84HSjppVaRx0Or2NeJ4xRDx2ugzxKddVTm5h+Uyz2zlX4ud1mlXzDB6KQYEcFGQWfc
H8X//zLa/Bz7qDhgnOZ5dLpT0Uu9N3VcNDt/QdDIf5qkORfnXe3vNaNafHvKCsogIsB91PSnIpIL
qo7r+yccim3pGRtkwe6uqvLQJMZ6csxmPTHL1vmq+MkZUJh9pFnuTEWryUz+/+kX0ZRVim1f6oa3
gTUQ6YhT1eqe4BgGHywcAKlBoquHmZNnVYWVvsoRjuZDPqebZ9yWg1xKSGqx1l+uF+P6wk8b1B+b
PAurLtaGJeC9jwwFVolQgiCL9FKs3q/lsUmo9CS/m9dzcmXxuxf9TwpogkfN8VDQIezM+GN/IquI
ymU0a5JXDQEfHwPi3EQEPkZ5TjvwhbOs4MIKdKAzx0C2J6RzDO+MFBOjX1/TBtsSxv97fiM7p3Fe
jjgax+9FisvzpdOj0zxN75J1y02R7s8D03Y4q0KywHF1ztsyB4Hn5KEgVAllUFsMcLo+qFJhh6O1
S6Fh/S1Gr6t1SsCwmazrW5A8KGXwm0iSXlv/B6HWahOBZwgaEVPlw2jEG+TZzAHABVe+O3eUIjgo
S2fApHeGdS8r/V67irIHLq62gh9rBXDw6W4OjiwGCOE5MPv1M89gYfurNljd7HqZB+JAqx9uIJtU
EAHBJZuGDR873YdZEdrnaTHWZmHOuU3hF8a/wwn6KlYY+dnAoymul1DQtlRht6y+jf+yUgBULmqi
ebErOQZlxkwfLoOuvXUtT6xwN/iKmsshNtTx6ZnM6zvjgY+1U/0t7J71Mwi/b/nBhQbhBl0HyKm1
vzqWh4HUAs+LBArANP2CKJcovlScPXTng2OYV3z8TMWIgP8iu9Ut/KkUvUQmBRulFn/ZErQoo7AJ
9b+97kH//+yK/b4CP23Q2Ro1vTGr9cBZvvPza/bcJbDNk9kfW1wJG5+BtQS0GXaTt0zV9npKc6Jg
slGN8r+2+AdEiVlqm9JQ4T90B+h09gtYNm2nQ/bn/ek3/7MjIReH1iQn5XxUwNj1U98JNeHnz0py
S1PcmxgccTAVl0+huCFn3UGMVogSDZHYE4FDy3FOiMIBT/gxf2NcdXNqXBdi5Gxnq8q7iNxIJbP0
ULYozhRVz7ZipWI4y4OmWb4uUaGNgieWkz1yghqNwoD8MI+uTYk5sNKdlD4Y+1lKSxBepJKMw4qJ
ZW6Wz5bfNhHZky6EyDvcS6NYPTlTAHjkB07nU/9J1Ehs/ioRUrpusT/TAB1DzHdOD6L6ITpaNdwe
RjA0iHq3CYKp08hIiDsKs+WfzCDtUsEKQfzIE+/n5dmRuCApIRPDrcwkFcL+9L10gAF0kFFLWg57
tyNCVB6T/x01ji0dCueoS1KqJp1PTjrw3bwBNIzAyalaw2f2HS5ssmVUnxNuHguQsTMPC22eaZtT
7+fIDTRFQT2XOMOQvj6tQKsv12tzINTbcgC+O0bnwT6TxkPzr4OL8mlN4ibPZNUthqIX+85AJFvW
/o+UAtbNNHajbJwrKC/AeZ6PoMdOCLHc0oOHt6/vMiyvq1ojrK3oygi4Te9F2qF1z4PWPr3BtLrY
0cd8unpYrmtJp7guEDiLMaWRrm4Ra5caRXCBndaY0Wt9dtjf5dLezQaFtLc2QhDcLwf/p8TI4xoF
OZr5AwFsothsf0apk3KsrBtBl0F+ZDL/6XH6RQ2IOeh6kWCAZjOvnCn0Q6bQkUqZPpQti4P8pKgG
0t3n6zHYMZx22XiBcaab2r6rXiJrJs1z0VauacU7jljTuvlJAWv6R/h78ejhsPmeRZ7J0TU7ILrC
Y9r7CYK955cOHPn8xpjtWLcsa5Ol8DyYYm/EX85XKEsSTtjkVMD/iIZCO6ay+QS9XIKKiHJWqfMS
4+F0EHWJGgxkH6/ikCC/vMbNXGvMYp3+8gjo9ZZ4sta/f0T+gGUz8v687UP/xLOgx4iNVwH9RRt4
3TfSYCbohx+dLGMQW4Us0Qdp+YPX7zss+4QOem9UUimNQPJaPkQL3paz3pT+T9GIjFoNVOwY+9fC
QdP3mR97hNU+jICy/u0pNXgdy0dg9DArpOBQtQx2EB5rvRnGx0X4Tpm5g6QpOlQzGjaW/xxzse83
xyiGj9/gzaXJtx/1Wqalmn25sqqWsouAsGJlD2RJ9FqLpiMW27BJHZHNKIHsEJtE8V33FZAVmriy
NDRepf6L2X4DkEsCjXpc7O89Wj4SZIEkw6wxn6h4sPMyNcpaXIXXlWAsLMuvrhkVZ8Z8bDvR7ISk
QdBbW7x3pCIL69yAtUhV3zQF9zw2v6PZ5682un+Y9mmctMtV2BX8T0qcJ2RipOrHZhCffOqonszG
eGalqvjuyDe9c9HWpD7NmpPOE9g3WvMw0+fWW8tFVoM7VJJhmhGcQeLvKT4XoWfCvqwzTp9G0C1m
szoYI9Y54h5RaWgx6Xg3VKur1oXVb7J2jKr+BGEyb6G4nXad9dR4Px3srv+751IsJHv8osuouX49
K8OEv8d38f3vd8NRL1rooRKfzbibcRGD9KosbU5BMc4JF+4n2DtSsOoo9UZv7Z7cIaxfQ4GC4LCF
VrGmKGb3zb1EXacOJwx24XWhl8MGsmzp4OljQt1jstF6SDlp7n8d2PbbbaefIWrJno8n1wHxNB4l
K0EPKN4at01GTIXJRX+s+1YnE75t7G60ajYnSP4ODRsQ7A7TtQqtM2xq/R8rmC/Ehva+GH6a8gWU
n9H6FP1aOxS6kesClXtvuxkMyG0oIQtxAWYvHNLDc5rCP6Aqu9BR2YoEZI5Abmsyjltxdej/+Cz7
ioM1yIJ4Lm5CyiJYnVpVuO/FkskDoaTrhAMu8PKImEgizDqE+INJdF3Hj4ipYjMKrJQOrKcwi8Gx
BLS53r8uV0abSl1Har8iKJtOGK0jx7IdK0dSvAMPp9pV/OOuHdEklOVRCvo/bxZasJXx39DvLu/r
JOA1x0cZXLkihsMswtEQcNoV3ziOYZo2YsuPVu/ueBnyfkw0MjL1MbNJt7BRDSFBjjw5XUNR2j3Q
T8Vpqr2PIk7lPQg1qD/AJEsPImZCLhvyI3CbmL34rdjs1ZjHHBYb0K4Kl8r+e6T/TtZH3PbttheA
MEFcwv6GQr9hGMtUnmEjG2LBPdK2Ps+3OZxSzS2dlEawKYp6nsRpbJiXneCHvkj++PfrakvwJQtH
tRb+u7MFGVebvC8RHQkrd8efRnXGpuunDy35Ywg5dYOSO8G0PTQgIbO+Ma7iS2aiYOATdVVoAQ8y
vTjMsrfzNM+PwQSm3u0ejOcrt2A5SBA0CzwpOlDfg1sS8OgGVFv8XtMbGWlHGJS80PsQ+zY9+2Gx
2gVOoCJ7mKYeKjKNcsZPiTiMkoxHBUcBuTF824lobO5+JOy4d3dV+BXLzlUG9T+HG7ETHzZcuXbq
C5OyPfDMQcBWVqAuv5ziQ8svrDXZrZoURZB0lPtRRvOyWAFAY6IqibKSc96B0h45rsSJgP2MkHeq
xYiFlKXjXhQRqy4OAvcy4FDI70a4Qtrrg5y/cD9cjNKLIA3zj3DUn4OXAuO1XVFML2U+dEDjbgzN
QLKpcrmf0GUOb615mRpCj+NtRLd5Wf+PRQIw8tEQbBFVDTH90F+7Lq1FkWGuxQ+/VaxibGTa+eMR
aDaeRsYKIe4J8mhujH4Am4XryyF6GQeedd3ojhW/ZaO3iFgJpPLjamv/LJPgV60kgYqYQc0YSrhb
vFUi9T1A5XtbuYSRqP6fOQKXachXEv/lQ5bwvh1b2W5UruTJMc6w9E5+Pz8yEUcQy+Fx9ctZ/o0g
I3jXMciyal4mez2CGtoQZqjk3/J/NnraG6FXXsP5mJnM9RSBQJqm+0qxpgKgExkFm5PxlthUuGSl
Me/K4IWyg4Gqv4Su5ZdeMeYr0iZWCS6wVv8HmV1VNPJcx368Hue1vDxXzuXJLcSIfYtGXBKfR8oQ
rXNgYrZb+k60OQSJjnX6lQQ9BKYB7J4nZdAz5TurlwJ0u2L76/q0GXecjgwsJpjBd7GWF+SWmiSO
fUARVhJXF9s4ZjRxiXY8kgenHlATnJoFtRaQa6H2YvGMH+xR+GTdU5mI0u2v2Zjd4CEIAgswG1Tl
4oDNaIE8UxnksBVk5obtO2BPC+3yQSYDxDq2FtjI1THDCqN3neMiy0GZVSbTglCi2xap4y4Y7AWm
u6SuVLjU3l2+A94t4bGR6dcETIwJGpWc2y6XWetyh9NgWLHuXeQYnVRvnQueH4NBeB35YzE9nlRU
vlSCfTQw8lIsXEQLPmszwy/JPln+eDYsFghdeA3zqowN0hq8ZdTJaZx2/c5SVjxSWDIV8fhDlYQH
Bs5HJ9wkCnmM6L/nyoVCcaRKmyIhPvKDUFGIkhnXS5M2pPOt7J6op3uRxKHUp+TD3M4LTx6IFFik
Cc6XF42SmSvuMH9dld8DiAwrvZBGxrEjYNq4cp+rU/uv2JkgHA03qv60CsyEw3Y3tJeAlzolafD0
/l6BQZOXBDxa9cmeWCh5z0So/r00oaRc3/2NoOyZog42kgzADzF5UkzF1WvT0H4ZKJxY21YUu7+F
j4hXOgV7eq8EGO/XnnwYFPxpqbDvZY8+YtQpYrtcv5xMiN16O6NWm13P43JVSKYfmRHRNxj9LyL+
BRfeO5TSId7EunzSTVDyfd3Y7pl3FAmaQRgjGYsRK3oacarRo47rp1Xs21v/ZI3iBqndG5AykiqW
AiqGRzsjSOSxUbekzKG1n/GhszCf3VvhzFxuFqdikbbSo/mvN1rmDvJx5vAO12p+7tUwiyxqHU3S
iKgNnZwFntjwWwfNDTYc+NUXW0Mpg7KFnkd500xNYfAa2M0dpqDembFX/Lw93CHKDomrfEQaRKwG
LoJZkoDfElOuzyVYHqDJ+8+6d9Sb83t8ZgLKVUboNjjdtXznYNA6d7Gml33Y137Yxjj9n8Cq/lSY
3tw/sOmcUlBOT1StcbMBWBeWTZ9U7n+lILwxfOFnRAmuoI2LRQi/C5zTiJO2vLYyAwMWoHpe9ztc
95y43FdTJGDyagmRwTRFjUVxLjI3X2XXNs+un0Lr7wRsUhirB/Tz8NFIsNFC74a1hmBY1zQ4EiVq
4ch2UMWYaKNSfzK+c9m/GbfycdFClQOVLIwGbuDw+UXmm4hzvpnu82XuPRJDNfRam1rYFoy7qwK/
fX8dkba9pDTL1I+gTzSG11FDWX7JQz67OFrzkLh9XeUKsTzQ7jeIEBObjUuJlPPIPZbL2CNUUIFX
3K6zV4Qp8tdeD0tGTM24UGdBaApMEJurV5ghKeWM3G+WWOtUYbxlq3zO8DnDWUvhRku0OVk1P8Jt
nt8BaIRdgc4Nem2LggOP6dmkC3GmAprd9GPZSjfMFpFFk3xu1h9JT9bJMNaSQQDPhN33sFL7uVxH
4qyhQcTpp2JHZV8bGJMYI1QG/QHWGyqABcvffLc0C0XDRUznBx7TTiUkUwIiTY/3+KfHQVbmZjo5
1HlOTLJo2cii6Bmf0AfsZAUAltiaOImmTlzHRyEFlfstUGYBhCsAKlG067v1OmNg/7n9/rGLvyeJ
oS9HiIe8Aee/azbM6PrrgWhOXPnvqJ7M3/4dGZXLDkV8UFVAZxUwMxOclwRga8PoL5tc8krznPg8
Tlnfz+OGT9GnIoIo38Hk2mAR/wdaSGtAxWdh6ihux37uy2g4ERIJa5VWI30H0JwHxML4leUmQm/2
DgEf9FzIpwYFUnh0o83S6j/hXOzomOLRpSdP5Sodcn6GQECu0JPlA+mq2j6VWPEZpJ5onpvZmkME
GNqYIs96WDHwtt3VZfCbJgdUUoZFjTSZAAZyOhkoSOSlEA9vazhbqVHc3xEew9WaABokecAE276J
HvhAwlCS8++Q3L1KiTlV2baM8+pg+XAyYEtN+9wDGbWdsKELogVwevErZHOqPykBMR/KGV+HWLaB
iDpcfB4r3owQoUr5XtYKRxHquuIhlKvRlDNq+Xnt6mAzW4wx7iu+nrVGWRyhxEz+OmQNoaD5toJB
EmLcEo1Rvhn0wnkrecryYMYSQEtWBANfvfafvJ809iEf2bPy2YgOugjX7fsCXMejayLHqSCNxryl
5m4naL9GIWcn6y1IdHpBWBqPdMqA5swVGKdW9GLSX7Ws6TzKC9QlilUSpMMxVqEYXbFjEGaNOWf3
e+Wk8OxwR+acPbU872Gw3QwglXHps7k5sX+8uqDYIAYePqbkj/wRe7EckWiyCKyFjK44ACFO8BVb
U7AVfUHJWpAet22e+5koTBImgzsEl3KxrQLIQIZHfXJR8B9oOX4hKrP94RwunjASaAAWV4FpwG96
4i5hgHfiByuxLSR6g1J4CgPorSEO1+zbNtbjxmNc+VaTR9Depkc8omn/ifoo4tQZVLS9dd6/ec1U
6BGgDpEcNZbhfnQUJpHADA+illnwvg8U+pAJlmBOJSgwVxHAV1aGNfBANwS4+3Hr2+If85JHIp24
fkOpfUPxjKiVb4+XR3u+pzzafXmg4/r8l+AtXw8kiTekfp6vFK33BHQFOye0UnB+2BvHTaHJMlWW
7uV8J9e1/nOgpZkJaNVV0TMSxPECv8eF/XLSgUsDddfhz7HG9v0d5YiNMoedr/ILFYlUtIuz8tYA
fyQ/HrfYHj68QVK7JsxvmceWKA8y25e807ADz2yjmSBxoI+KKbu/S91wMoo2GhHEZ/snsYgI2QuT
blaBWPKRMsqgodpqB/xWxK7s1igbVAEUIL38TUvnm8qgqdM8HGc6KC7kmx2bJ5bnuHlapuVYv6Sq
ye6tw82QJAZ9Ge/yMk+LC/00WEr92hLOZUX4SmcT6Epwj9zfLCoSMVU4OhI3KU77Tr9m/3O0+6Gj
wz+QwJqfuYaSJ4qco+MZhvQNoxclf/mWXfPTZGwqcbQUmPtKrg33Y1AErT2K1ftZcEYN9//xG5vq
we5vlkhKa3H7KZjdD7LQ/S1s6X6kBzG0i+9jZZLIC1KK5E5GhbhI1t8PItfSC1e1atPS7e2X7mbc
vvb/5rFuIl9vwbwXlcD+VT9JDhlKA7IVXjaRxaC1sdvQseyza9UQDolpIvCNyQLoVHXKNDaf2FCT
supwklrKawangVhCO5qZbLiNtCfCVtY4B1dorzNkz4/83cfdujG5eOp1vjRJ/B/+ijHP2T+4xqRX
62A5sl4pldEzWWn5ZknecLk8bKsnjEuOEOHGDb3LanJLzRxU4rQKnLOwZYqvEjaiuoylDC+qOcEu
a3/JckVGLB5YKbuwJMSL5FsEg68jNp70URJU3DgR2ydW/U2GLhY3gyPuqWGl2qiBB8cgJfGHdCUM
5C8S9/JDj2+DeAkTzC0szdz2q5fBEcXP+Vn1Nfz2M9Lg6nHsN5EogbFuTfppILaYg0FT6i0RYKPD
+8XgSnQced/PzES2guX84zfaOP5WIKTWTS3DuNFXY1qG5AVkrwVDto5q6CA13/u3n6mWdxV5vj5+
3vTn4QaqqggX8GFLopFIuz8bYAlOinyNv36eCPvqNPVIWH1iDj+Imvo+oicSh9qHDrKPGSDqrD0t
+KDT4g/dMdFjIVQiVYWg1XJr9ftCH3rFhH/Iuuf/ZxT/faifNJv5FqLgOhC1yQbFZ4n6NIxeQOyH
CBlUvMfweggmsmtpkwVYpBfb5bNAtqeOQrKqdWIKgYelCRAIGEbAxc53fF+zMxiUC0Gc4lJ8rVsw
LDKEBebetho+xhmJB+o0LmXb++oa1j4AAoZe7coE93wK8IuRmRkpojk/9tYxjrT4mXBubciTzWsL
yz3E9pLuLHhrBwFI4EB6OgYwVcGVWkLAzzkR67zvg5OQJzGmgRudxlMuHVw3r73kaA0ouwlDZrjH
m9eCTpsCoRAFyS1V8trQJ/+A6qlhDlfWh+krz763VBJ/BEotOps2MmvrFrdO1GLbBg+PgqB2aYI9
a3e8Ebe2fR3MFUFDbWvvuHDPtlx9OoXJ2NIiz9XnYiIa0Mmvfbysp5XvtPsgyjiWHF/hlDG25PwX
5qyHiaJPjo+WvhVDZ5TznbY31rUeg8/zJd0JPGwojF/RRQJt83Eh4iGbRXsA87JfvEt7aq21s3bq
iaALv9LlldzkVahteOchLxavwhdQVBXTRlYgnTUciCJuyM0UBvkTKcSN7HQJl//8d11R+EzEvDrf
1aTmoDBz8Av3U5gBVQvdwDnT+tBgfqCiv1TFPdLr3hVFSCqV28cViZ6qDhT6P1Vxg3RmEo0yGjgC
3NNJvfS4wVMuwKPa2Y8YT6YxjAR8+5rxqdIQjmCeJ/Ks8tKhasoxFNK+JsuYVfF1rg6qRrKn4UIc
I6iZlV1D7ak5jyfmtwG9oRk5Wkrgk3elABtYesBtPEhnTFdQHDj9Jx4PTTNuwSB3lumx+NFNNTL4
0W/D5sm+91m+sgLNlBONg3Dp8U/HTQEtii3L9X7uxhsUc9WI1pJwb+WwLAJ2kQth/VOfPnlsM0LV
KJV9yo//8EwTWx5kX6/xaK+ck9uFpRosU9Zmbiusgf+Fz3JkmQPuHGEAlJsM/QMmrDCI+W4zCpPy
J2qpDVPE3tnbyGd7+4OdmYENmAkI++C2TACWpYL0RwRNpChMkvFEYlZ5MqrTMjbltYfIkwAHXNsS
trKzMZzNvCH3fNhbqMgGMqmGFsYF0ry9acYkIh9CCjcGyz7gKvtx2Hisnrr3QoRV+ImjlY1BIdol
lSZL7SfKySU3unsjOO7DmQqELg5MsfBTRshBJRrmjswA//4HUQAGLhveMBOpXacEFV4kIAwqAoBz
XV4CwmoJJ3EsjtxsgL09cE/WCroh/hx3G9wnPGhf+ZuHdBQzVRXSWEk3fill14YlQy+HrRlqgWqJ
V2VL6sZk4ixF6GQLTR1lWeQm3bEouW8R5X7qlUaWhjLxjkQqHXUZADF1viNMdHJPXUCp6OwCy9g7
uhasBAnfzE6g7QMYlUYy5FYTy2/aSVguVKU1ICkgs37Cnqb/3qu72bLnioFaxNo+IqiVwn57FaAW
qrwiGCWzoXRLsqrlYdG+ixLrtk8cx57fKOoti8hxTTF7JwacA/TpfokMYlpUjZhE38kYlunP51Sh
4aZ3MdzRWGsto3usCvm+zkKSUmfHe5agzRaBezbKkH2ns7wXVt01wKZHNSXiadAbfwpBZaUxXSWY
CwX64bBT/+MIvaF3gwATKn2rAMt4Y46/LEL4eTX6jnJasqDsZ54JDKjnjb8CtfRVQ63vkXhl2Vs7
NyI8XW5DKNNF6GX44dLunu+xc5+ROcQJinHeS/uPAOi3IqX+fHfj+aydtYmYSGYxmMDdIv0tilNk
7GLxXV0rucf72hOPE/a+Kpsn7HbwxG8iNThMYMrJw1P1tYKCtLXfP6p9tWpbG6RVx1IQ0zsgKm+5
g7xQqw6R7qiZlrRBdtQfy2GIRW5mKgR3c5I7Oss211zYMcmYaNqUCoSrB0eEOgL2ff32yXwRNAbm
O0SB1VBOnc6oRtg6J/ThV3WVLHRm8Q+RejGAEdsm+UpPWD78J1N2Poy532HlX8bxqdh5koCWi7ym
y03EuWhvVhvq1ijuQtQbir8rDAlHJlycX0w0iPDSxrCDu6iMx8+rZzNXTQh7EspPvFmhXPSCmhLI
KLEWOF6AmvNLkr6VcKzxlHLzkZEqC3H6C4YNU4yQ3LedHMbLoEu0LdhEEgWHcI7R0D1yzDGHQ42A
g7xIorEjUtW9ln9TfiQyF7STJRk47jQTy8YpJ/tHUE2oLeoF6LeudhT+alIOqHhblgIyAZhBKkjZ
p86qu1cA0tdpSP+kiJNMgE2ppCfDPCG2mEN9HqATHv3Mr1iedoJiAr1HIU2S07/XBh8OWphYNUVh
OLi7NlPWbLEUKx1tBplrsOug+KkWL63DdlJ9bgUfMBnycbS8aDDncXvGSWHpSGgKm0lj+6C57Fyp
RZcUMZ9n4E8yi7vm6yNaWNVUbiX5MELuUeNfDN4eOXMmiGark9ainURDxJyT0HEd2BiloYGsvLL6
BpVmjzskKYDaAPJioIr3numdvCLmdrCgB5v9N6a9QeX3I8uigJKYwOqTFrD0FElVqidqjwmULjna
tJ7+swn5lzqUGRoFcSgz+/Dr8Io00w3ifcdHB6M1/Rp3DqTXT7S34xkJdI2QRluDD2Sj6s9LiL+3
jpVRqGZ7AQIogQwyxhGdzTQIzF9GscMrdoK+ztosjSsb+J5QveUk/4NqMaiO1XSzqRXzO+1KSzmA
T3ibkhU/stDh4aSv3CaCa5NopFG4Ythmjx2qrMBZz8q1YN6oYy538IFaUlHA8uFPoGcmlCzgR5pn
4a2uqxq4//iSigRHvOc3bKjAmzs3Lcy2q1b0EbyokmpEkLz/i+qtzB4iT9ocAooLGS2CaJF8X9jj
rbVJRWA2puZCOy0EAdvUjVWGaQGlg+/DMgOGrkVFTP7/nmN0Sq+5QcAjxTpA3N8+Cd+CQzogX2/Y
/U0wtHCRNrF/og2NcNb/tFdJnRa2PaiBj+PsM4g88a3bPkTSU6AIF6TtFWjKJw2fq1W7ARmIRd4O
HwnqQB3+qV/UsZHmYBAMZy7SXP7ualYuXyAVzIBLhhwucUtl7r/nJulkhfLCmunXaIkV26dfKX9f
e+NZo6yOSkw5UBf6s7AhiB63kop4+BS/BvDO6Vx6szDUH3ya0Uwsz+Xt+e8sFrAVMl7cNlm+p73H
Ixp4VmUsHxSSQnnaPiT+cthmZpPis4i4M9hsMyYj4OP+DMuFBJfn9qaYHVb6hLs+fnm4t+TNTDbp
tzDktn1I+4LFJsE8YrfOLDBkyulfmOfGP9f8cxpqTjWA/VlKZbIeXprPkyfO9ZRpLib9OEtDdp0n
Bqd74hXCpzDRE3sNJjvcDTuSk1t0iAnXiA+H9RBTQqOLX/HTA2OGqZLdmBGpopRqLloHSnwm5eG+
pZnctko/O/O0zv/dJVWToGGHLeVIE/hhLrwNw4NDbfWykKxZavrfC6B5HKDt4IhmFBSYAY4kGWla
Sk7h2fzSHEhaBINXm0bKlLy7UYtv1fCpY88NnyWXwMVFyrt7xDvkdRIGIH8Ln4V9VIr1mH4/q9pc
F4/dQ7fY9JMhmTkcFx8l8Fqb3gS+H4Bmb2v/tWaYimvZnDEKFEYsW9uecc3kVJhK2GMzqrb1kbFI
C5/kc9P7/2KxHNT046Lc88cr1c4iiuaBjKPFLkPKucCTXJtKueLx4/KSURyrpWdog3gkhLFZseDo
V+W7y+92Oc//8U8/EQ/Dsy8stz1XByelwic7FOCLV+tnzpE4QZTCkv0sE4IqiccnxPKcW/50nV9X
FmVrxAc3rTt9YE72biUAvaDVklQdVu4nu4j28QHzKGtRabT/R4MBqyXhsQ7UyJI9DFieVoZKgA44
4R9TgLPb9RI3fMycBWZvYEFPM3uVI7+6stypDU+qGYZuPuiD7wMQnwSaRI6FGV6UEqWre6EiNcXQ
YKYyOtpPY+1YVR/VR+2VkCnnFYz+h+xr4bq2OXNfd+rpTUAfQ7uy/OZeSBzFdToTroaZh8Axs8+4
uWXD+O9GXBfoAjVfxa4CBHEr7zLTOGXIxnJqCJ6RoLXfrV0UmVIq7xqs33iVyA4Gd6AyHvGZt3uL
lLd8A+hAuV1i/Mx/GtCUryj7u2WHAg0TTsRdLHHGQ+kUWUC/moguNG4bfb3Q3VpVJbUkaWU+UYD0
qlgJ6q7u7mW14znqFrJad2zYjhg8iB5MqZtgzSJHOMNfpGcfvReBZwU/9c6w4VjeKKnudWcuRh9A
U/kqX1lDs0eXFL+uaX7oLvsB/obgBKOH4e+rCM6vrcxgMCeyWXg1vKC8qnR5nzKMTz43Sda0Zk1Y
Gcdb7oB4QQmcKWHFEGBAguRhaz4lWmblOZF7el0sCcUNr1zl8bzMnWL4L4udfUvJ56diFXFZm27E
2ayEMUA1fC3kIo1XIzLUXx/OgmSkblWVkSaAw4s2eID02GBmgOSNd4al+5Qjhk9mlcEiHy47ZzS9
QgMyNTDK6JOryq2idFzcVYcUa4JuNR09sfGK14uxQoaiYFd8RT2o0tP+JgQlEm0ZKXhXQZG7Cv6m
LEpQNCkIM+plKR5oLZv09GWbrJPHc5Oc1zek56dgephsddCHx4V/bEFu81pOfLxivV3lhcxx5zzb
TfQbw7ut89kcpeBVXoNFleNOia0MtCo48jWcQBsxmIl5p3w70Ixi0rZyStmjG8L3/K9q57wlzoR1
er34V2RjaIvQtrzk2LNI36bPEy8Wz8pGwTlBS3DFSnv4UzsSJDcURkQc8Dr2d6pLuyimoLrFCS8d
HOOc7agmPv8nlcqEktXq89vaHwW/+NqZ2NWv2eOfzV1SrdO1vbxtl3EiGhoAkG1BDk+CZPhs/BV8
H14FYzahcWJkFHQMLQtWuyOobfwlgu+JJJd+OzKH+7dl+8hfzWCIqzXmNnIvf3lF346RKY8NfFGd
If/IUCZXZ8feinYy6EL43BK2tgcmm5u1x+APjeC7JexmMVKpkpVF/ioZ0aOaTU30hZFvG0Gspas2
MIBoy/PKInYNO87vefmFdzjg33JqDxisopUKcYqwenVqmxkw/7agxKOSwXIS6kM+yIlhei5VsLf0
VVrgqBLhAURTdWdGzG6TLQbKRN14qSHTrNb7vpzpLY2am6ItRltRhVN1vpnqGtNrivF8BCsumEls
k472u734aLMBt8pCyIudZotWWhWX2SxyqeaSIhs3tzkLPP+V3HQSmQhb0DQaS1gtrMcW87z7nxLV
VhKctiqoVW+LtZVMMBXDV0BSe2MAsyLwrz6x12W4VCDpwhu+/Etr/HTZu5ssV91HibzgLXpZE3Tv
qEUEGpTUGnCVwI9LYh+qmoYdi5DSwayw1xiZRRmG06MoWPqyrygSHkFrOB0h8H1IXqpYuCvgjrus
/wDZiCKLVm/dd4K5PmyfE6hs4iYiEt0aXBNLzhapQaDu/TUgONuyMVwC7337VktdclMgIv5gpxub
UZYrMnq8QGqpXfKQKZbh079Mc7vsLpB/brd4IhcX5QlGeKE35fcABNhxJeownyVmv16WuqSEJvKs
rZ++MalhCrkGWeRp29UY0BKTzP/+sOjNcwfaFZku4mwwe/sX+snO6b43Wz9UKTv7jyqS6Qkn44T2
Vbyhoh7u8L1jeBEIgu2wAv89bNrKw20rvE0P1lL6wQLv8kOVFRNTigMFJxbSAgOa3JZQWOawVx2X
ZQFnlfLnnh2bgHdQcs+rdURFzAGHGTAgPAl3gsNwymOj7IsTi3Le7xwZsuGcVQkrXqgOYj3hgyNw
r1c7sDcfLf9OEEGWgKUlvHGCpLlBy4BHD8ratFD6NfU1UjHFmQfVbRe2s44QGcrcqcJblrmdHKGt
HhNyn8gjXS44ttAfcvP9187K58DZoqld+0DvVmXtdNH8ucTdKTy2CaMTZXUBGMvkoJeVw49LSiwc
ycbFSspeVdmsXFpTT/D3FNLTAKAZTFQ/lLSLPOfxUlXN2dBuK8ixjKOlcMlRF8Mxjfq0qO5YyoES
muu3wAXx0fjM/KNzXpcHK+0W+kzEy8wK8mYnIT8bD9kgzJPeF9JEsyE1aB7YtZNKDQtLvvcR2jYY
J6xzjQC4hAJmwL7gtLEDThYP4U6i6UH87OxXNyVB1hKBiKegF+0C9BbNNDtsugQPsG0y0uikfx8F
wrNFbMKi2o4dwqmcw24iRLQNLfPuW87VvIFUfbxNFSugldFQyxMrji0AZUHwPuX7sJRSvLMgnhip
CRZvu02kJKRYwU9vI25xyZwbuGhfKiYemsla+VLKCUNFMyVezs+PCrlvTrkQ4XY+/HM4TBI8nX7B
2PNcm7YL5nkwDot9kl9p2LfPRokwHmvuvxT6V+AqgJw895e2qSS8DZJb8qjbboy2COucZMw0mub6
UDWyyA5Hy41zqJJ8vIHgd3BHlHkUg8O0wFRBnD6jxs2ru/r7XSHJuCSjNHsX2XiXow5qQSkUc5eB
RukAP5i5cF6/bzTzqoQMNA7KZfrefQB2AFzxLukP1PM32VQY720GAQxqeeUPglrpAgxex9uqzXVd
YaC81+OliVXraTMJ32fkq31sShd+jHTCLmYMQB5dLNa7SZcS65L2FozAibfmG6isWFULPG33cBan
Om6NiuNkOp7udcdNFn771rMQUg3INzuVAJXqkujBx1CmkaG3c7CguTVZwxyNf1hGfPga6Ki5PYVb
4oUfIiV0WhuOCy5ujPE8LmTPft9ggeFD+n+dCcsjjjR1qtQmsiWhC8vWtTUgo4ooQNjIdX4mroPd
PschlzAmAJSnmHm+ED90VEwwsL+nZSPOjRoWz4dzTIkyZ6CJfZoBcv7cSnC/Wx04v/tPY1VevoV6
aLaYz9ygwt7FhcwKz9LOSVMjyotFRp2mbUxW1wEDBHNKU/PfHQmvrwA1MGbz9mt9T5hQCqP3fYlA
zCayvTvqssLJG9ZzcXHnI4fHbckVetPq6j81VmErCIGzB/ZaJ1fKrvViYwzE4TRRb/ILlZ2g/OtM
l+/gWw27JdGo+DW7INuzHZY41mEoyEeMLfaIs84jhohzH6n4azA6kW/ySCZF3PUrILyZ0xdkolH7
QTX5ILJqpXSKRqRASkFqjqYFwM98iav4pZF5045XvqNb+HApFn3nD43hSAMIPrmnzNq05oCFmK6y
uWOR64dMkcXsYvTucQ+a2aTapRVsrbSUr3A7EiLfu8t1uQUvq/d4abXYk/y/OwyGqxZwxVvWsSoK
ZizBExd/5u2a+EqEgeLdBr2w9x5FtF2Ec93+mKnAdEG/sd1KBn6aP8xQw/HGl0a9zjrRe4Z5DV82
5PKoDvt+iObDaMJUcs//CvzeJ9a82dThsluqyjh19e0KQVXjeX5pSdbvM7TREyYAFs2um1urPv50
D3VyU0nHOinIxkPJ5FrAS006hnrTqJrCSZh8Pix/h7qEHYNYb7xBGauVLVOcMZwqa4VqqAWLp7qQ
iEdL3Va4E78k9Q8Jvc7t0Y4loBFV0nepbXTcFrmozvCr5o+15o+ZGtJ2uiV6ieiHJsGUjvRa6Q8R
jgf68fNEcP5U8F42G2SKeywYcTIaGl6bukEYD0jPUyuscfAO1HaS2UxXESNsmI+Vtb603wcJIcY6
xmQF+X6Xq8hOeVNuCmRQJMZmB2UIZWd4me1Bl/S7idMK6YEDfUPSn04rMnQoGG0wQ8Murh7GevDF
QEsZA2S8j46+UJVzsSOLV8XxJo912bE8X6SYMzPtkaly3HnarE+tAh7gRjYfY+eF4C06+3oSDMEV
mR5N0W/JpqbHp0VMeieky27yaer2kAbAYhsq7YnmIrOvs3H6CY4QGEvle6l5O278Vxx/BrqE2Byz
Lv/Wbv9J+lE+oNSAiakyp7BGYwBW5cvxlxUKSJzudOGgTmMZmqfAHqdtXlvvd+tOA+PY8QlG7bTq
ExJ28E1OZWqpq/TiHacKXskHvuxuTYBpdAvSRH0ePwdFMIC9yhPwJWV9AcECe95DZvEIR1EnJReT
3YX5j61vqv/nHm2+/XhUwcDh5PbxFARPioi6IhDgE/WeEZSYRaUTbcjQV3IWEyOimkZ3w3/6fXK+
AAMcOeLyKrXgyIcLDaDZP9bY+wxznREKPThz/XIHNgl6pDDjXd3dzdPeOWR1fsIVMsy3q6rbL6y9
3N2eVs4ylbRPQ+Dgdjp6UZbpQX2zQS6hl6Sdej1O2JT+WzD5vWIp/DwLO/pR2ogs7a6iPBHeIcBg
dUcFJ1El+V0VRCw1o/G5VlvMBO5HQiAkO/txyYHKajqa5zMNR3DDgkDini/Hp4ANHRKCpW5YPRE4
f1GTuluzpmE+l2NcS8X0rnJnSRiQC9TRr3fRpCxRFhdaV2Ft2XGzlD086HUQM+atj0ZEnrQ0zR9i
hg3ZLYe/rgFj9nCM6wn6Q/viD2dlvEcW89b8aoesKBtff515ajLXw95+12TQ0F/4MIjvtf3Ydz4G
2iqxjEy95yS4f1lQW5K1FwfWuhxJxA1de55oBHZt3pDrGX7sjPA9pTUhHb7bwR32NK/S4EbtPdPB
XRd25GD+V2UzOWisK/wlo7kPrUuegBGHwtAANRLr7ThvIqYb79iLK3wGXlZoTHlJFFm67PMawaL/
VSy/xNxo/gq5BnXoquzj7lfPdXgT08twEXAfCJC8hLZFV5HvCfPljiy8X4RQrYRKaA1Sr0JaaJVR
TcoidMGX9fXPTE++MljhkWknbM0p+mfQle9MH+CYHDoC2L9ZmaYnGHn3+PRDbaLxzBlG9mCbqAqF
79QpXJYA52Zwa1JIBR4nRImlkTYtkg6+U1Jh6PFU84EXps9CUZaDEPx6RtPB46Ii6YC9QIVKRXLY
SZcarRAel+hnkxYaJFDcmxO5uKzB1qtQP18T5VP9tdUXmsIcDCapzc9cu89hHGKLYjNgkIPEn45f
ZcPo6DhRlTSINkBqe5EV1+vwP/n8uf2fu+pZ35khMdEnma7VEObzMHUCc8H5Ednk6JO1dgrGHsYu
fKJVoUz9aytjm+J37UIKvzFMYI0LzKwboIYkMJG0kklNKHwqMtvt1HMqirf5tRbY2iMmpE8rVjHF
TTYjQMu0asQTbpJTFpsrCmAnRu0zyrgFQTxMJsEr42k96cxAUC1dvvIukEPtovjqGCc+MQ9xXg/H
XXowkMdFo1rvf/P68Yn6ANc0wtpqThDPdDkwK6o7m2LzwF9g9Uu5Ijrg9fLyiTL5+bDHd6Li9CAv
Mg36j/4M2bhoCl06C/jX2x3CfNpLjp1E9qnbnUtG6Gk3zy7K6XOjfuQXleRHwuiNtfy7IlHjAUVI
ggMaAhIfbzmUk0COAxR/ln+CAlIly/yC3unDhqTI1OHJhqCiYM2r4wrXLXEsyqABGom9o9rDuPPS
RvbhdEnBjJq3wU0Q1zzVjhfGLO64sq4BhSf8PCJes/xxyAZU/ixALvyB/cAh2Mj+2qNWoiSiA7Q/
J9ETar3P3ki6XIr28i4soVaJUgTpq2bC0QC/rXXhSFTldldYNooB5a4npkX00qHAauw1I3HZMd+l
kZ2VSOOUdMvgfRWT47QB6HaYd1UxhG6lE42/Gje4OZw/p5GtxHDJb0Lt8yWP4KUjC885DgzRI2BZ
O0iWtyuBEUjgr1sOZTjVlwFMjwuytEWPRkOtO8O/qJmDHpurvi7jJC1WLAQGJGaBdMHexRelWuHj
8AhoBnpeUZJ5U5NxQasd6YPFmKuCq6CSi/MSWnB+6Z6AgVLEOAPgtF/yeTKXnVpxQbtFqAlAsuKS
KnnP5zMSVNwdnIKoOkehzQ5u2pmhA+a46tHC9dsKf4aNawcKdMSnxsN7Q79futNSDRSmdPK3ePfK
eojdtGm3CnQCCqLycMoLDtnGTVw2EZdGPPNlp+Svd3ervTUk2m+lgMeJCtXxylK//0p5KISZotPb
Hkj8HOZ+tsjRCgSM1xt5N9bz1ufm4g2kXUgzZVrVbTwnWK4b7Nnul7bg8TC/T3+5l02StXZI6R2c
MzBVcdnCdLronvFl7MPiJWRpkm8b27PyLEByr7XFbzNVKnF9Mn/oRtXIqghxhPGNLgBpLQeL3LG2
jF/HaxK7vN7R7HyYKPYWWCTvNDdudnwEQmkDZdlTQeFP0Vi2sMLutwPOLRKYY6HT1RNtuvgkVTI4
mba3WsP44oGSVkY9UJV24Sc8tkliUx8V4cwtIAXS59NAiPMgsyuBMVfnZl4wWpNzXmIW5p1E/NER
ezc00QJaPNN5MDMA6Ghpg3zJh1pWORZd/pqDmnkZjX4HaoDdC0eTgboHueIziddNcGDH1tjF0xfS
FDxOGa0G0a7c3KuQTly4uzNcC8ZwmnPlcDrv+f3XjCmHvBYkT4g6j5Lxdl/nwLSrKGquXpoBrzeX
x+fVi5ttQI2qJqdcUMzYRPG4PEj9HSTWLjq66qdUA/EAO/ZFWK+R3yLhE0oFq0f9oyPbh5V2eL18
/Wq8pS5oIhreMTLXgG9sTnBQCd3fZJiHq+GQQT0FyCbdJAL9fWhC5XOfM/UX+Dz+e7KOLsjgd1Bs
7dZVAhJSD5HH8BkVGFTjSuCq4gWufNTS+fC0Tjf5Tc1btq50n85tCYjbe/qF0NPitCnkThx/mUHK
TFBfQxxOVb6i8QEKuJvwif+I+u6rUX4VaGLbPQ+JNR1CKOJBFboCOdtdJLDr7jQkSaprK+dc9ZUA
fDU9Z8+v2P3hcXuYLR7c/Z7LMawYoTKS3EKzeRax3yQxln9pKwn9OTDRepDkM2ujN1wfuoJVP52j
KPhkBctHiMR0I0f9Vtgu1puU7k67coAEzu8eBnGidOO+5YLGlCGnsoBgbnQzMSh2XPlvioyWu8iW
sZ4/lyy1OxezfSxnuYZnwyF1Uh74J7W+QMZDXCQqzs+4xEUI33owx+kdHR4dlbdr/SlPNQ+8Brru
BGi9P8fP3Wvt2kX4Oln8htrYkCpaCj8yRBLWQRiEKhTWw53/cZ879nf2kCJh8raxLh0Q4UnuccdQ
SMvyw3w8aOdcAvOxVmVjKi3K6RUeMYuA4lZwptRvWDAKwg9QjMKv1gOJUqrtlfGX/VUfvJLX1tIk
iMStP/EcrnD40TwBMxKjS27kKmhuITvvUb84lJC6c9MeRhEpY24VDZxs5BMe6SySPVd66W7SeUe7
I3kSkuLRMVTwDTv+e4N8FymK7JgxATkPEmFvl85NWAm8HGlH9B0RcPB2vbUjrJIU/qvqPNYicA9M
Az9wNL8vPmbDlkQAn/l7tXdRQLSYdy95K0+ZwtV7SKRDn9iMHbDrRG6nj7oqPeHoro59VRHbPfnM
JwG7TIvaXzP5Q0s9Zu6lyGda1Ize68EH0u++RD/O96dP6U4bTxPJMYU3aspJEPMwXlD4tKVXYYVA
G1lqP4DKFZo9tVQmt37HS2UOEgmNJmMyHCBVVqVejZa6dGIYGFQcui85iEtzF47SoMfAlfkH5RB2
M8NtPQ/8Blpyc9vQkeOouG+Nali8rtQKZgc4F4k2oCUh1/T8KS4FDKGQ7/kXnxgMSZF1bI4RkQbU
BaM6e7Se5g4UZk4dKykbtREVzmk/Z7kSxVnPkOjKIBwmmXfk+0X6S9ais1LtVaeVuLccJCNuk++8
6YhEGHCCiMllZraaLITbNO23EhIFDcBywQAMy2KZsLmJWlAhW5lKI2heiJRbF+tXXsF4sPpi7R8H
MyTFRHBs+/felci3gzuyr5X3Khc2s5Aqatpjzh48/2iIfM5K941G2qLdBDwE6li6JrXCefuWarvP
c828TCEc8uA8kqvOnW8mubvbMfo1eOXvsrMROgHBFaupim3fX9i2pTB8AwAAkdxCzLjF24UyM1jf
KX9dr+oy8TsvMlm1jzdcIE/g0/duNm7DAuSvHIjZaakyE1JmKxzhhRXqzGUo7NNNtlfsWC7PET1l
CflSucsZKJ4W4MmhFHEC375Tm9mD7da6MKx11+x64TJRkUlbgUR5pfPxrhVhG6Q1bnr9oCGiEJX/
d+O9y0Wyhxrug8K/pJNTi+ZyqEqM5Xeal75IXSXra/7nRYNTFtPxCoXQfgUTt9sx7nt/VP+cLBbD
JBCJR2ZftT87fsth3T7lUK/CF+eW7beLxrJ11+feBl289XF/3zsCF17Cd6Z9S7jx9PQmf79smf3V
0zAMsm/QoqAgcboTMWE/Ed48w4TZv25M6t7XoZbqb9kqBAa+jrvfkW8vueVQM+9HBbuqsCG7ZAyL
ytqMJgskxgynJy7FK7n8Xz6d+gezRj8it4bn7Hvyw7qif48TRGswz6p4ArvadKFn+Bqw3jMZuOBk
yHiOh1Ciz9ONMz4zxUoVIr8g32LoZHyZm22wh48YFuA6RslspDsCtNdYqh04WnRk0i+kBpfWRhUD
iY0PluikIF9VIrymfkmFr9g2Eq6dCJ0Pi+OixgPqxidE3AD3uBMxxoGMNL3E4EOeh80GfAbMdQwD
ZCgzTPRVpVqUugKwTq4sWjwvGGneSYoJaLDzDOPU6Q09AxgCYuPKrh9iuOKt3+VhlR/UePLEKGed
i1Bx0cSKbq+gzRERcPxqPrXqfb/pnlYXrUH1OGpn+ODn934QygILQkQgs6f7NPePi6+tUBj3droA
5no/ULnae1pvPHuaI0+9Bi44nz+8xzY0HjrS4U8jOZ5xlOUJYJqzPyKPqmA2h0KqIzF7Ubk1W4rx
STibW6ObbOalsncDCcj122B57I2I/7+k2IsXVpAoHB7sZyRAbyFMlyGiopPYz5tcmJQ3uPsQY1Fv
b0f/EKmjwtawoRr3HgOfTtE15+Tv1Rr2gxYPq2qyfdSoqdnDNiBB9HU/lM8ThAVDCgqhw0ft4gvZ
XFwAzIPhxKQTvacTlJjpImhjhvTTlzGdRMr3I69LxvEoZbXjQcI7XPicmgY6eElTiwge/XZrDn22
rtqPWYuPOQq6xdDzcX1/q8vBmMVz4an7hkSWInINZaWdGJNKpcXTzuomIPyI7UymBc0dSwtHDGc7
pgVXo5ri8B614ECXHrZr4XrZj61BKJN062MFdXE48SR6X2N38cnWLlpLIh7Dxz30+0mfwGm22+ou
cAQ3wV0Ug6/yJYl8Filobg9VZ1mZYFCGablAzmMeqSeeeK1LSymk8fQpD2NCFUswDK46TasQqRqT
4rYM5opx2dabGoPbz0BZurpQdrTwFCTuzPPCPuKH8556C9PF9Z8NnpO+U4e1lqtduIvGT46Qm4l6
97UCDIlamMpTO1LVlBhvSXRyFMCPRDQPFiHZ0Qc64WfFawH4jEokFOXS8TUqEr91Ud7QpxQRzyre
BB3fCMq6FArvMXZ+L3Xq5Oat3MWbFP/eybm5gbrNBAURWXt9tfW54lrNuJGxKdRjMsrKQ6tJaFXf
pj4w+61AqAm2WO+UJNa9ExkjyA/yB0JUzsMMNfRcEjvy8K0E169fqaYm6EDA7BPwkyNAPqFUl2zN
G4BVskQVpMKshWiyGjgyg9pVsYCffdAze0ZsejN9r3Oz16THnR29mJRYRPj8DmL0eIWIe3M5bmKA
dHKEm1fMGrbtZMxO58ur2HF9uXcnIFhkFKkEKSnbNuqdRaDe1sqLCtQuXVudpSpaqoN4RIki/ISm
He+oxvyudiMVf/y1xg+Mq4YkbGoaHHQE1TXHY2yv39Zwg8Zc0Hoeg3m9nSBsEctM/moSY3sSpsjM
2hq7B0HxA38G4l6HA49SF3F1YiYyIzLl16brl6OQ35LHfHkZqhNcth8VXfWTfcEfAuC/9eHI3ghi
nrhSKl873cyC6EsoWCTnGxR2ibRh4AUxyJLObD8yhlxNDQg8RXDBTjdVDKi6hfHtd0oa+z+W0DXO
0llg3b4cLh08IVV1syTU/Xk9I5NK8FHxCHum88BfXNXvz7UA6k8+9aZ/+8FL0GLfnpJ5El2YSRQp
mDIJzBsCZ7dCVPQ0x8xaE9poXTR2WuFZ0MHF8/JKB3Gxi9Wn9oPDPu8zfzhaidkupM6xBOLBNME+
2Cg0kXr9EuJSRggr+3+XCbSi16ZeRGsTfWeEjJk8HLaZ2ugH7gFZZ4ngJa5wF3eCnUXqICw0212p
nmhAsh7P1qC6M5Q69v8XfpuvHJ0dzlgsAvoHGTwGUOnNXzW19PUjAxa3e/qQZPgaZFg/uBNs/dOE
O8qrP0i8eyACl2GqA1vJ57KlMFuYzIOTjxT6f0PvAbwpXw9533KgkijVdXykDd6NSdHvUD5P9h3c
uYKTvuS9TVWP1CZ1PNVvcU1TjrxiEqSjIsWJ3JjdAjKjn8gvFQF+BfF8FQaCtOUQI8eXQhK/DjPC
f1xY/jKqtag5uegxkQrF2HqfkDWCMJQ278rvt4BfQ09hls4dm69NR7JROQVREciDmQ1O57G5S3kI
g0m7XsPYNFhroLiYa9l1W9hy5UdiGpzGZ3zWJs22HKbRAW40iaMgWYZ87LgUWrDcIsvHON9bUYAS
CJCMq2oUU8Cz1qyWLxvxY0wQWwBSV0QQOph1Hspvd35tsc2/fq1deJjdUVe8ffmGgMeJrr+F2qsx
rI9MYOg0pmV8btaQO+qrPjMD46w7cq1bcRmqGWa29lkYMOoe492llVHYPJN26YtLPdcP42I0HEC8
iMLkkhHviCAmc2EIkUWmhO5uBj22HgVvlVr2AjOEp2ep0Oh/ygKU3hMJnTy31Ep/kisdPFkIEjBA
us6pVdWfbmUQh1e1OuFXkLsUnHOuhduGrWtBv+sDzR0uZWCLndQXTaKw5vhfq+7bawGstcE0ffr3
jpPMM1fBZuKAtk6LXC0sOPDRnohl+PHaHjr7L+WTuqXLeS8Eyyp94zr4M6JZvF+7c4x/c6PnCgHf
5SUus3oQ8/3X4hqd09uUz22pGlPYg6VxVjjTDi2znVCDUBwjKO8e0bDLyZQbIdZ7PIMTpCFR69y6
fsOggoZQnWXCEwdVhmHCoabjKR0yGBTCztCg1V8yQsZrBgLOyUXGgrtju+hi1Akv/jmVRCiceuQ3
e73FIsNlTIqDlJu2G123k1S4hU/IwF1tm5Up8ct1BioK5/mivA7FfUqnYVHemS76rFxAkAA2Y0To
M2orrJmQModUGvB7kGjAKD8iaMCypOZPNoxnV4m4GKHOy01PntoN1dSt6HyyiSFHU7W8j+1DbxaD
jg33Uge9A3r0XmLYGwQn5AvZnCjZ1Ey2Jv2d7KT9omjNQ50znko7DOOlfqOr0pQxTZgRuh8vobAA
ajjL/AvWXQEjOQ1HvtmHh9Ksh7ezfL6sE++J1wNCCrdDmiVcEyX5eFkrEKev8IN3cRYVPVi0pRwb
BWxpKFw1LugOgZgUFmWDJoRnDKSvL03P96fq6Rq7KNkL+s3aS5HHOZLQIYD4slCdNFnWFIEuakX+
XbpUJicEBXRK5mZNOaRqIjMEZX5y/prdPIC6C3IlxO4z/dtYdhNsdkhpyg9XFNHwF2QwSB9+8DIt
MteSc9AvO/VaSGTX98ggtBGqhePQkAPU9/Dl0WYpal93FOPTZbeGT6ozxsSTNiEPU5yeNS9JUQ0/
8DzvsVZIGb0w0xMOxesmhwy9uaxxKASsW8rJsGujtCFWu+ogwkRN03Od0aXUyZeSW3BNEk9L/pvb
WMg6pVaDx1CuDSERFfq5cJD90KzcaUJPwdJAefY1p4/2vUvY5nbTrJXrVNllJXSDaajXlKijsMPa
lCCgLcGK0U7fCKYHq8W14/r+x8f4LxDZTD7L6jBNYushYJe0MFqg3G20iPUy8OPBaU9A+n83xFO0
v5KdWf29+fkyjl9R77S0ycG2dwGx27abkOLwnb5iR8ijmtpAabrGi6mw3ffyvMXCc88lFdFp0EuC
jQupUy2fte6Gsanp965Wcwkp1Wx57U1GpCAuJx+LkSZUONmT5dHIx4HPCa3wwh43BDnNtecO1ENQ
1ldEmx5eVXbwmJBwlG//5w7y8vlCqtLfLsIY7lrJUelnyNgV7DYxvI657UKAQiARt+RlNLQuzuDe
d7AexYKkI3w8YeaGfk9p/F5g6gWHQMRUlJfiXZFB138kn/4qvi+pTlvt+tXRZT203meWZG1fE2/n
f3dNaaoC/gMD7b+ZLx+WJI3gmoazJ46+lRt/OZ5DD9FbKI09tMvz5Q4ucs14L2ZHOpbXB4Gsvi/Q
nl7q8si2BgozT571o6nX3zxl0giq8a8MqrDWneYiBSadF8bB8QF968XVF7apMt9AW1hDiHN+lc++
/aM2sw397boMk6Y3YAh2u4l8yNMZKCpV/bZIbRFQV1eOxVkCwrTZWgzD9uMEJLq4/+DJA/MJ0vXK
8R0yfF/ocUhQIrMLTt/1B52Ig7WFXjJvbTeBwOsPxAe5TUKLr0+YZDRVcuwd1R7sG0y5lFK6rXfU
MN1gcvapje9ZvWjXvz2aB+fYDhPde6QYzetT7NwU4dmGcYzlWg9uQ4Vzu4t1IK77qDrj+C29oCPp
UyRVbbHPZpwzT8EG2PWUnd+JvuEq1lX9ZbOtei50pfVqMNygxTv7wm7xwz33XojRAu9LScRTCA4H
2qTYIUyu1+CA1hJWkf9eZq/9JI2Nvtk+A4W4h0hv5mLlfIA0tanb3YI26mqmQRTH3OlWuKNZfxL0
/VszgGdT4/G5Ng0S90b/hgjGUDmWIQaB2BNNakcwaNQMUqXq51RdVAjsQdNrTDXJ2eFC3VlWyAW1
FHbfTWIvpFJYqweFigAgIIHDviIlax5Chup0F9et/BKoyK2CIaFHaqZqcs3UbgSpVG5FlFq9LZAA
vXouDq8a8icw2ZGPH0+9dhZMhQ4nuF6LjuMeTaCFY1L62xd4ubLaHN2q3t+b4yeg3plPv2UwMO9X
KO7JAOGwc0eYW7GSSBMUGZda/63rTeGZ1+4XHYMXJhdu9CcmiwxzSkIk44yY87Qg4hLDqekRQV0P
0AdpQ4fhMc+x+BNRImins1FvdATAMmE+KON82dOGl+mTlwEJShwzTdl4J+7iU+qp2jA800CBmjDK
l6XB841M6tngWey/WdbPP5MzjEr2BOdAVY6XL70ASffRxqlJDAYtBdZrPDHYoQppDVssFryusnAW
Wt3fkQ1kiFwtDhMQEunlZ024utyur+ic6+ZCX72jhuXBtReDqGawhH8zoWoFYdnVtKtAMwDUdvU8
8oFldw+FNE1QsgkHV8KH7U+FWZmbVVtDDhbCm0SNIXK41lXzX6+T1OQi/hhNRZbatSKqBrvaA9LC
rMVBXYZqhQeFaPWb0TTln4C1okEmpatAmqiW9FCEE2RmQvp91+FM8i6j64BrS0nFxIMKhdN1B6cs
0zJ48/HYrlAyDcbkZN7xBBf/XV7xi0gJPmw+XFGlBlu9L4br3n8t9HgH9tL3nBaAx7BzddZExgHw
LmbvtZFcMr77SwhnuzUN0qWP5vbbSdsx3UqMXPwhRGevOiN4UfkzmiYoML//WHN9Sr+8TEaI+boq
jmaApW2x0/ZzN/IL3y5I2+rxuhMzYBwvwJqPayOevThsZfq3lYU//tmjDg0cMaFXHrWyWJtNYY1I
rtYbB/Is18BW9dYznrVCLZ3XJyWVKQqmT80AD0Uh1tbjjVvBk24lWeaBmW2HCFeNOoMAEMxOpRZS
R3PnPSZNJZh4iaS2txnUr+QX4Se9pUiKySo3qaENXsFGd9fDo/fwNHE75BX5D/Niby0uuDGVCkL7
ZmbxR2oXQJmG92SxZdT2vKZ/BhSt0S8JeflKCt/b2qrWsoPpFxd/wgFxXWGXXmU9QZtBkcls/Vn6
+yxomBnWdgrXjiWBryOad8Ol7k1r7CpKASD4btrZNwSuJfrXDmwWe2fR+ojKx316c/B/dbQFpXZ8
Oze1+/L8IimbLJ1BmzlIBYW+QZwLWByhUoJWzIWovUWZgq2OcCgxt5iKmgYhGoi65dSzNGlq/AUV
GXouOocl3DWqjrQUeZaOQzH9TDhX5ArLT6/NLrXng4WyZCJ237n6tieXXRMqg6LsYFCMXd1RquHf
9e+gGD03SG/8m2Tg7hZfqGGJ9TZjjisGGkYLILql6bbWOntkbtbu6vnsXibR/fy5+cemOv3O3F8D
JrlESGFT+SBCJFsKnipliWQXRDRziIm2f+YNhfDQTUKtVTDYshtiTd7WJMwCw6ZgZZ9LSWP26+oT
o/DGz/YvELwE6KSNm0KqdawstFF55JUPKTZpo5WWwe4pDYMreA/KNsrvHhPQZR1YKAxF2vdb8m1I
tqMfiYmpaaoRMGRu3NSEn3jm0+N05/oSzaKC5ycypSKwpemb17ql2yeE/9k7eyN5hHXDThSuuARS
G1d5hcuSHp40J3hUTtqGr6u4L63NHC0p1wBJ/SMuZRwSiByBikSh+IdgdiVLAMhbrM1vNYkfVyR9
JAyyBk5wV75PodNONt0s9F2Ydg2iKw7gra7a/5q9zlxHJyhYIwSnGf506zkEIA9XdlzFtMC8iGUN
uYoLFW7Qmwsfo8PN8a9x0GyIygxwjw35p2oQiYmkthbRTGtlMcICAWF32JPKkmcikZxXFmFQSqmQ
o3Lm4uC3Lmx0tK1qTKq+qt42y0FcEFWUbf6crEUoMvOJjk3FwUowYil/8Iyj2KGoETEUGVv6idb0
RF75kxcuUPJKcX6+LkKEme3uXHGJ2neA4w0ohA2wi30CR1Qb99Q5DkvauA+P/+XRDQw3+Srde/z6
1Rf5Gvut9mZblWmlpPbwp3Fz9RAl2vBIy9ASFL1JEuvge66xqzQvJW0MuEdyFUyQJcjB7vIdsxnr
4x9QkTeqCP88BMWG0BtzqdMbmhzfdE0YzVHorN2VD8QF29PriJf6uINClrrqeVNkxBV8rQdByAD3
+qLHQIo0zm2TgaSDTgMopTQK0AVk0o0V/HndKRSIdo/FIypuehuu3EG1xc/ZfPmMiUSn9+/yrBVE
s9nwLQ58xVJ/g21oNc+wjW6EJq0CiUlZyxfMUi6dZ0aOHSnE/nvgRP0KkCswC5Fcv4pLTWlaXbuF
Pa6duziQsuIN4boD0Y6NbDBk78+TxLPJYVGKzFQOFeWpP/OaOxC4OBuPM7RigpLRdpxEH/LxcSyl
NEr+cZcyBaUBzwOZosiIIaPMjIYqLaN3hJ4mLLcEqdz1oF2n2RcSlUVEaPjqfhBN5frtIFlbV0DD
P44iCAiQhErd9yEFCOVNry0IWTSteJFQm9ebg81/nY0+1+qW0gtP10/XIGoX8BvyNwnQE7KJPjCb
NhbgBLM2vTvb7Dz1vEDEYXTqqq/6HlXadReyPyBFpSZ2qbLLeaTGsW1iKxqdb99/B1iJM37L8qek
xqHMsj2TsO/e3l4gFMye6/zAJhgpo/UXv6KE/GIQEo7vLzhCXnIDZXvDYSOLaBaJVtuNpDP9HfIo
Km0lyu5by19zPjQ4E1K/pqCJkPikjVNLb8P6LT+JzUapThK4w3Bk+mF05NgF9jdhRygBi+bL2lGq
WyQVHjtY10kQTpa/uD+mVGZISzA7gd+NeUJfJsyKX+kNvPhYMAx5V+Iv0u7UuY7q/G7BJ1EV99nW
tvRT4D8+AI3AVRyy5A/ajj52rupIetlYXCW9cZj5n/fhxH/DmtuUPte0SnurL3ouR2jLzyOtXdsi
jEg+KF6bEsarlPvKwzT2F3VUp1nbnhT4H+Ne7uD7GZ1qGJkAPMFaBsFJjKA+FOkLfhP/jcm2DE2g
9UufVMx6My9VYszmDNg6OhS/xzTI+sZrrRoO2wj7C30rSMAG9q6rjqtjcCn0R78KuEjcFnYlEXzg
S3QVFJV2iAVqgva3Bp/P0ThdHURiJN4iPEu9/PR5gS1uBZun64/XbzLG6dJIGc5/7Rjl1hXKfkWZ
OlDl+kNLarU3WWzrt2smGi6VkRd/PAXyp18sTDoAP4K8BI2pLI5zprzE+bhaHjimKP9w1Q5UE9KC
kzTgHnmSCJHQZgDaoXTL/H7l8FGjVHgs9oU1+RLPzTrFkQZr8nJSm9+Q9Kosuhoj+zk/8XGfrOqa
eFtsr7pbN3HkZ/AqhejxtR7EyoFGjbcp/SOkOZhecii71HXtqHGiu0h2hs2e08R9WMpLBip0cnI0
7vInOyzs2beUemRoUYovlchpsECkiusYc9AINMLAFZOpPsDtFFboBwakdcGnf5lQFBt8fsVNNKLb
9hiew8i/TMIf1+4lm9Tv/jaqXcisyfZhV7zaxg0l3aofDr6FWJV6852ypQcZ81rv8W0I+505+rFO
kYtcPjHLesGsrVapQHLGEKQvSnjZZ2XQci133PxySfmNsSvJw7Huzg6ffmyMd8X6NHhNCYXBYzhC
YpYQQRAwpiQ6oHBZ4hm4IpQg3QkJnb1IG1HmasdF+H4bjdbHGqo9+T04IO5hLPZDApnbP3+e+Uto
2eO9UbQg6gcOISwVy6eRKuy7XZgJFB37bYq/Uu6JaenQsE07C5G/dpy+oymWTqzvZgIOrQjmlWx7
h3Eb33ZuBcwSvDoRbfUtvNd/VXgasETRh7AlRDssJ1b4yx2WwyTSUh0HtA9QsOaujj1RmVE3nVs+
GotevWsOctS/B2bPlNJA3N1zyStIr9Rm/VEiAChDW0BmMPLhzbYJbgMgMG633fmV7P0bDoqJq2oa
US0MNQPHixBG8aR2TfT+eb00bcTv+BuVXh4vWMApJRvKwVa2AWm0MBqHCTGKzL4DljRSmt3OIUbl
+wrTtpt8YBVqiFra9RjKNTMTmUyvkqH9lwE7xr5Q1u4TR/SLn8ybc4eGuMFbP6utJRUYiYvstLYc
dK0mWX0M+elCAAPAnplfNQMAhmFLS5JU7qNXIokyPZ06rIiM0lv9SpOamZs3P8NcObCZQx4wsW5f
rF8T95AiWzopL4Sb5aRykATzWg5wEqHmAYZcvnjAVuXcJxf/ldPzW7G9Q0mPDBXChF1SgyCa0OJk
Y3V4DON0ZJEARl3yhyz81kdIgPGYpGdy0OqZuAPm1W3i2XcxrBOYxSai2Avw1YbMBjvw5JzPWTkI
HxOBIOaXgfdVd67ru799JHDVhMrXuYu52wdwu1MwMwknYMSTIEsCgqgpaoUadWjsTLv/7VXZFr6I
MQ6WxbC6o3xecYnUqMjuZa2iv6UIZ7ztzJxPiiCf7Yam2PvwHE5BjAT1sLg0MLIi+3+pQ8nxgsxB
ROsL0tx6cg49Ktoi3gFFDvn6ZLi+nxGGnzD0NXWyeYO7pyRno/H5kSJZYFON3XBLWRJ+rtnmCheI
V+4PJ9lgEinuIeJI6m4OSomVF/IcpX9L15igQnrHq3Digp0BoN0L1rys8jmEUXVqc+S4rZrPJ8e9
H6Lr2P9zrji2zR2XDHTnlAzq/nARiaEosHPKUZmiA27S2ETki6TRtTmStvxwFnAkYF/kw4UNKrAt
axr2MEDrsZDcbvQqOcY+JYPP55gPE8L9DJoohcdoJp+5fvf0eG9Ph+yK2fSWV7hDcJIrdrQ+ZeFz
hWjAbN1Mc0wegOxMhsOcK7Tn1OjHTvGnjrrYEdBL13s6/1+GPUrWF/NgHdK/Fh63HgbkStrDFtJQ
PsRSe7c28973FZr6hmYqU2X9kEEVNGoTc2WdjZMMRX64wiwIS76HhmdewXW+mNCpVg7A0uF+lhLs
hpjqQ4G/shDKotcxCrV6MxNFSnYE0m0kUdUMDCdv3vcCCe5y91lsB8n2CaVj3rTPQJR5cx8j7mVI
9+kV71L/NKx1Dg04aWqTk6QfxJ44wgL7NY8p1vbLwU80dkEZto9cuWZsdcf4f38+ZSAzF6yo4Ugq
gGstlo94ftyYSOgs0qq/y6RH0Ri/q3xjyxLPSfjNDFHC9IzJdDMKDMULryJuePQVuHCPi2eXgOxq
HT4zwrJYyo0u3YomLPBUv8TBsmzljzg0nnT6Wa3bjRGwfV6EeGgH0MTxETB9DAFHS0P+gYerEidn
DQpF9aiNJ5/UdCktBJ96rikpr7I94qAmSH2vpv3CDP7WikB+oqAyZaPNmEnWdnY4kP6M8QtdqxFD
ZyJrOHkOeg0EOqFAK84um22lEw6LC5Huscvcvm+EtJGgbxbnWU35nv0yGTsen4+YVV9MpRshDfeb
C+ZUV9/n5r5z7aqY6T/5Tc4FJx9seK2v+PvxuS3nDnyhhq9hMus1sw1RpBVQll5aCwJbHZo2iaqI
6jOutliVCwR+wVSw/NMHKNxWuOG7NYRe80ZeSbp+tEznrp45vcXsU4kajB618FABYTUf+19+V9Yr
wSwVEhMIyXKjWJEoktdBaYU0VW+vjqtaXnzoldbNTM/exCpVpry6LDBW0rg0WP4zoVUL/sJIAfVW
PJmhIR2IsvN65EVic3rt/tUmqpw/DCXeXnAXiZIZbL8ql9T4jMwh/M3cRkDfb/JxDBbQ39vItGJp
Niqc7o6m3kxG86U0eV5kiqfA46gFV6y2nyeE8DHZW0eVxI8H3ZTM0WopZXod7OZxco1xdVL6/mVm
TI8e3Tsb5dXyaHKjuLdamEn0IYLBrK2W2u/UcERxm4wL850YmS7LCgJzHRDzifnzGVW8PHI14L7+
PYOgtLai3IfJWrS9U5m8BLePN/OjgnDI+xTj482B5zqU8RxXRst8ZZLArFIbljOCv5YRvZHpfvta
/IMevhVaXtGqIs4pdY///lzlsM8+iUYOig3B1XSkB1f8Lv+zClX8uVbX4wYju1MTsbfB8+AYDsob
JSOFH9MNXsKMqObmm2az39+jehf6TRTFMB4r0N68fgEWt9+l4WBa9iNPQtrv+ztyx5+PLJeaFrqH
7wxU/qHSpJrVaNvn2RAXiXL8qMVR7hy/+sGKASs+EIwqVgFd77moKAWPRSMGHMUef9nEiO3jlNOj
x7k5rqdDvuuTsRmV2Uzrz2zE/x8oJODE4kL34qNf+pc7zDYhpcxc7i+QUg8eRr2X3ZGzKg0GCkQR
51TxBKPI6+4eAsEQDszOsMEcz106qezZxkMMO8q2mDy2pSSQ4vVr5C5H3WlgFj0Zf388HyR1fpYC
ZhzZfCTrP25nR613RfD0ODQyOC25mA46L4QNHbfJfvcNVyTXqzN8p/zrE3hTf6MO8TaQsI3oxrPQ
UU4sV3N8bmf4qCIxMNunliWEBDAb+TNoG+Tqj+C6/4zT6HFI+px6b+wE1PWQjKPU6N4WSZe53j/G
VCH5FzF7bskuU9ysSkZODzmL+2SOvGPSF/IMCQLei1FHrnmvnl6TMqVeaImaRxjhnv9Gzgt6V1BG
bJBfT/kym/CZ6MbuNtRPBuWrePNZ2CohwNzF/Rn5nAAU5E9Jm2hOF3GQqYD8ifHzg2NE+PhL6ztM
ZENBe4LUvlqiygyYkLB/AsAMkau/ukSUGQhb7Gxo63yOGq9A1koQ1UUZIcrrcQUU5D2KZ1xKbpu8
1LfyAy0I8pyTdwexh6GYP7MdQf1HtVOc7rOn9GVFPr2gGRivDAwWsTpv9y44CMEIrbwBFsRg1sd0
XQZe00L7uJu+yY/r7jlSTicL/Hm7AcFutytzZctVB/PFVakQy6WmFE8eHx95L1KF9igYFKZbX5IF
2HMmOiX5c/GDGxqwRpvi7BSwYjvOFf0MDsWJutuEgJDZ/gCPclQmFoHrsi7JjEm5k/IraIojKJUT
t9sT+zCUC1/tGKRKYArPMtTm9BkH6WgnVBdNgpE/TVpEXOzUtqYsr8B91H52FSI9zTnUp1lEPE4t
NIEC2TjK6Er3ucIwflMFSFp2pznaCLCYrC6319FGLuRtK41UjtpsI6KQEn9zEwrbwIQ4K6qmbJyG
rxDVvRIikTCeFBLqaVvobvlgBr9eMOUSHrUCk9yIW+YwEt33W25+3FAyWHVgrSXKkinTW/8fp96r
sG7DIxm0+YHerpOAj5TiZx6c5kRrMpGTqXtyCdT8fs2DNBLBu8h+T80pf7cIz4yuwa2Y1I4NhILf
QPfqGYXmqPy+3hbNd80tytbJimKPpNmkV6ffGlwCTGRAZHplonSY8pyGC3gysYKwoiY3IKUestxV
EFpVhrmhLR7jpF6x9OHdOgUJBbBnqEBGfr03puLD9ug3S81+OX2E3k58R6H1vwQlmbTiOv2Kxd/r
AIIeXxg9GPEkyB56RaWsBxNjEmnDSFNcvjw8qZWxoZ4iyYnhpXW8gmNnwqZj9j0ddiDXLa4yx1Im
2KB5QWL4Ro+VcPhH2YCS/CL+60kj6hPgXjkUWlFDBgLdxxs8P89ztOf/LQlwbQQWpM7/p9cMMFhP
mOqzcaCyb/qBhOd3eU/zpxKpQNCJM8yudvw74eAxys4kwHeVjR+sMBhP3Ttin8GHBILx6+8x7A1i
X59tqSRxzAm68Wb0AblEehNBZuncP1YXU/RhRU8u8fHtsiGQp2LN8DoJ8d9HvLnD4aF9nAriFXZS
pCW43G59zu3VGGPKZQDVgC9mnPWsnVwIFpbyMCi35+jL4b3RYxMcNqiWDWudFo9mAaBfNSceMgAD
O2EGM7Y3u02Aq/b6AULWl/zK1cJKyJfb0avk3Ef2KC99o6wmeDABISsBu2EKyr4/alG5VYlNiY1u
fIHasWBVE7I53ouQq2eJ9sFoOEP32eALOtKgmNxYyjqe/kCPbZPVf4S46QyCcMc8shoM7F++udF+
UXB7qzWsKGZK23Tm6B6EfiF/2ftCGtN5TLHPsxad2MqbNF0v4ohMBmFBoGcrgG7OZT8yN41Hat3J
sErHE3BTv7/wx5bhRh6PQbk/orEabYk9sLwQXshQDVXX4tP3mIihjbMPELrRuUB+Fa0bX1cioPpy
v+/oyP0flaDEytZ/sPlhqLSnNvXv4GN4hEE7uW0LHOZIFXCaZpS17AknURgUm86E8iRu5JwzlKM9
WF8EzPO1OQgUHje3BmLCVKW1lA3ySmdiOOGDSqkFr88dy29zfBRFk70qC/lfhQTfRHz8Fs4KoQ7y
Ax/6epoYDIgT9dmdq4MyFd5TjoqnqWSmI6zp4cGGqB2oCYXuQAmuYC3eeza5nOKa9qcPEOGOXUUj
yR0rD1/T3ol/UeHsXme6LrQVYXR7b1XsxgXygHJC73qYrwDgUoPBdAsfzrtEOomQJVRiB2+1dEm7
/TiN+SV5YdDhfQBoXKGFEefZQiXEQidIOju+JhpNMDJmZpCQLuWJ3Ks8zS1OvoWaMMYzdVwnscRS
1gyDYKuVKsfJBrkw3ESkOz1+NlIQ2tA4aKLlF/YS0ztZX4Yi+WXf0eipdd6ezAlOAhAZyLStJy2G
nfy7RQaAUK+gIkenw3pqdAHKeCXHd6zAzuytudgRq5/t9riypNw/HqWvYVhQrVGA2OLgTdyHcPOP
47wUZCm0sttmTAdSsYxzFmBWLlKdG4bMg7fmUb3/9d5F/QFBHIu3URdWevDjgeQqrHYzQmesxB5i
X3njsfKvN6D/bsorU5I8BX6QLTVdVIKuqaakkAMdgtg+4TIX4KcMKFNVOATyB/QFgCgqFOhQln90
DXqMSlr6quu4Dz/lfGznovrwBGWnGEoNzB0wH3q30m7KVytDTshIpadQqA8oXSVxTxjv2ODaSW3W
mFv/mszcXzRvBsxjRDwrasnyRqykyfzy+smHNBAoN0nL8txOtfk+HpshgzRFPx2NQRlCwctkxHaW
MFJRKqKp2GqgOSGVkGKhiVhcBS6nsmbHjXzBv+TLe2cWjpob6vFUkH4PROc5Zanx4TzCdrSnKQgK
2tJRGexqLYklCCMrulS6jN45sV5nVaC1geNAKgL9B333tQkHAMAGTea2yIvhiX3NO9ybx3vomySo
9b9mWStXHthkoa/OCiCOQdv76iQn/+z5hFKo9fGjirH1NAohH2C4Iy8pm/GANCHKZ8eLFS2hVkcN
vcdcP3UxF7Fhu6JYj4vzUH6qGW7TQ2Y3Ok+OmPOyOxcoO7h76MA3+Fih89kx8LSSczxs95gO3buB
BvUA0OQ3NB+k+Urf/jOyLB3XYfZN32UZbq5Rv7hSb/3YPElqFGVELzRUN6nMf8PLDUffCO+PSK9a
rVdHsBUDPKsgDvvhP9Q6T2u+bYdpDDrtJQ0uPZ7D2tTJhj9Vn9uzXO3aPcH8hINTGAgjJ4A1EEoW
cnFwTBUwYVEQUnvybrq9fIYIlK7065mlXb/kkdEdH7Or+Rxk1yBhrbFLhz61aVw1UtOns24kvGBd
gMf+Uub+l69LdC/CtYDXevuIItWuubMSKwI9OWbLt1FFyOv5A405K3Dh/0+ZbnSSZ/jKobsJXh6B
TQMHs3s7tzHJnSHm69oiRGvChcwMUpWJhyqfuXORcFcIXCrImmetOZqEd3BfHsNADl5lO2JZAJKC
VYgSAAG2kFrYWYhL7DREyNX43yxblZ3h8CpWEXjjTJh5O+LIwysADKgVft46jX/WRiOAC6bD8DvA
IV37qnE+4QfftWEuJXl3tnabwokeTGcGKwUtG7IS1hwjNufLgImYQFW2QKkHIGrvcWNRe+khQPQl
ODfyu7QWVCkfPVV5UNeoX+RSUrOuB2gLeKKQZMRUBfYlmzs97GAN9B3z+QxWzGMx4VvftB491WwL
BxBacoC90zeeH94FoQlfcwj3BJ9kEPE7iMHJpYS+7f7dUNa3NDSfaNc6pAiof19VotOpxPdGwoLQ
ykwzdNPfgS2xEa+EmtnEr9ngUuYszR7o35xlOGbvNvuIW4YbCpNM3KlJ1wZ80mIS09f3t0OEC7hE
0RHAQI2kQk+6V5fD6uVSuc1N/W9XtPmQb/jN5UppP06+xbwv5i/1x2DOAI1xJBne1xpeucf6fXYv
wV/h0SBOsArPo4areIeuwioJ+At4sAfJEwNgTYaGxku6tkREmJIT+zFd2lTnkg1Bj8rWVKEnjhah
idKMnphG4p5iTTVnzXN/7PE/SII+88l9rPLnnkMamSl1VsAOrUEjFIFXIfHDOXkJ6mnEpcE6w6Y6
jNg1ZBnSugMdAQPaEcoiSd0c65Ops5qg0dJ5FM7LwQxXUU4tCgOaG7pF7bD6HqsOkvuScWuvSWpm
r+ZToZvu1eyJvTnov448Nc1jzfK45KiEMGlgI+fuwHIvS0+1IvpanXhceLOrjk9Adcz9ZFOAX2zs
6nK4I4RKcG9MkUhDMo5THQCTc1EqrATsBTF0g84Ews+ICES4vV8u45RY/n7Nx6l2EHnkj7CVJBj/
mAp6p1U4KsETP7kNpYhMgBxowvZ1Ke5j32nISFmIX8e0oJtBr1owznXHJXg8nvlT0ue59r7/ztC4
LbaBDF1TWg0OoTnC21X26s/w2hKeWmuPgiSa1x1a2zFSwK6pJWIyZp3pbOnilIQt9dPAhmvHcYm6
5OnYrlTQACL+raSpaI0v6Rsh1fIsHzCuLmHMAKfIWhf1I9iuWjtOzGarq4LGzzj/Iu845HxQrFBJ
IFa3BesoZtGr+OEjp9n3MPg0mAsvSyogFpwXmeK3+eYwlt1fzUYE/iEFl65oROCy81yJGdRu5kRv
lbdIIkR3jPgeibL/BLrHpmUbtFRoEbQyFsm5qKk8XnYrOkQYOAytag6gNFknz+65rA6lmsHnnqeh
6Z+o5+nbSIjvoqxEAoEiDknV35npsQ99pdC/it/J5nCNK3L8N48HwfYEst8euy4pZsRIAtqHRBJb
pZGnNDvcfH0R9KRHdygkO7IE4Jl6IZ+iNCwyqIrlXY2wRd3k4TzhPRUgXZpOxE1YLNj3DZ4FpGF3
q+YwzVR/G6cyFrq/5/iKwC2f3HNv9jOmTuCXo7U9ro2965MwmUlG18cB/RDi8FSFex1fjYPqvV9E
iILJjUzIc1adI1yhZULP9c1hBrKp+KOI1uGguKSbT4+Ooxj/dTB8Ymz9CwlJtuqMg/ACCbysvVKu
HWcLvsYpf1EI5O3QgS80zdJ7ajaKqhrPeyoCLWRwYcTHtNfnXkdGoP8IleorBfi6p4Vn/lQRkHm3
LEakn0Rgeba5PDVkKzUd8MQ5Bvs2b4ak0o3adsC4oEhj+CWWx7+ttIV1Pn+GL6rdX/ueHTM2en6h
oMvXyGkqvYQw9wgUtiOpCt5o3R/mem0csSAODURyB7ykHykFnW4x4thcKjXPCRPxLM7c2jit9aI/
PZ+XSlB2rCUEZeTUT0MwOj2TtVydehnkx93Rsui+6y6V+rFzGOu7ebkzlVHe8Sf1AdHDoR3r73Jo
M7KuccR9fLiot8V/qOAeBeUSD1aXZvVpvpyul0260ZkcGT9fN6L+N7+Lm38bvPrpBUh8OnaJjvOx
pkrPjNCti9TdgUuLGMFlCpRRYDxcabyhHFCtAhsGup7FjaYtXllKU2AMncYjphbjCObMhA9Ci0lh
NF/wX++u+ten/qoNb+/sPmeKkT1Y80zeOA5hdtQNdc6MVtUWzkALXTCO//QvaN9UjmGZLwNb/C5E
MGX3VG4xmg8fee39qYfMNBCATACwKUy/ACJWX91Gy/HSyT99xE+EOURAAaW6XMCAVVNRIef4l1/C
Yhd2YkgYGC18ia0bdFkyV4rfXrU93GFeslE6DfPJmqFE5n8KQRYqNAzizlitaFzk2+3YSuv/1Gef
KoXheiRYztiK+0iAGJNvC8b/Ys7vmczYa89uLlVNEjFrHnQOFijBqr9Z+TvyWdgqWf3whVL+vSoO
1aZOyT0erC1k7VOQ4/yLOhc9LLM+6OstH7eGnnjtHqJ2iRnArf7Lyp3InbaF22yBKeZ/2haWTEfa
fbJQ1gtbDiHnKPxKqS1z4TGjmnXmVhjcX8WnKmSZKxA3vI8Fvo7GuUBlWUEzm8jtViQ1oNdyfctf
hNeDj3zA5TCJrgV2uvpjJRHEkfr/aNsO8uSBJLseIHXn374p3pwb5b1f6156hmXmFnmmqKZ0qfQ0
Bzxx+MNuVCBG8KiGKh1RyZp8mPFUtnj8peI7ebL1rw1AcXtF3slYLcFF1EE7ORoaeBeGrhxisgtp
TVSo1xPQ3bG9feGYDuPM4Kn/pMieICcG56RuQwUX3srFPg2m+fucPcJ4uljLqeIFaJ6l55EebHau
Xn1pVb90x6koyNBL8ajXlEHZWk6I7Dk8Cqrq2rXNtW5s98MnnPBtjY8Nl5BBjEHHjDLS/ry5DtL5
pqMsEqo6PGwpwIxBkq9vy/Xt5LY7s5VEckt1VrKwZ06KTXrSX9XvKAJu63mYHiQ1rKTgzsKfix+Z
rQGvGHoZqjheMLbfzNus5eeN6ag3qTmgp0g4SsQ+mXqirYfXNhBzs5Kb7mYw3aNEqlL1j4EJEHHE
cxq6RP3WULyDL7hWiRmkFaO2wq9G2v4y6N0IbHlPKyolcSCOr6NC8Vpqu722aQxDtg12HsQKN8Bp
vy8aMT3QOIdFxJnCQDBiYSjmRXvPdtojjH9aHinTjnx00wHwH78+3bJNHyJLbnZgt3zmFnescNuv
5G0ZKx/ddsPk6f30xmhSc5wnYsSh/WWuUr3fNXIR8c86yNSvV3HJnc4k/gDmQjjzD8livAJBCL4y
4zFd7cp2vPRk6mUb4tmpGxkhPHFC8cT/vdjExi20WkJYvQ+KXIvKkh7lpmuqdo9gzSBEbhI1N6Hk
ZLlIey0q+8PienXMKNByPrVV3st/cUchDMLBeKQaeWjJi5L3e7l7WsyQk1MmrjK3rlxNY9KoevwH
j9xbFXpyMFMha1gY2Oc37IISb5P6rCOBzgz/+GsACFVEwubGCoP/GIgJUZjw0IpHHLJ1Pt92HtAK
ElO2QNOBP6UKThUNB2Wkb08aFOFv+F+wHfTmE9ramMvgIP3euFEwn/KSiKS9Hu45llnyOtDqtYOy
irW5c0gyLq+HUx6PTEDiDwAcWc8628WLICEkLdim4ssj91kpeOS0tO1t+L9iMvp/xTXblPCmopH6
ze9bm09hna0IWvQq7ltFXL9QAReE6CkAbjIh4MItC9DSspZRdHsZYzw13deccSPc/KNtdcFK2dFf
rEaDzH3XfVKJhDVjJfglQ2UR6OFsBXzgBjS3GA7DeGOPa4Nf+Ux7DJTybAebcBx7lQjxzbn2pkSB
/iOAtHP4WDjx1UdRyuDjDVNyBlAwAnNWk8lQk3OM8eBa9UhtXIECMAt3QjyqLUC15366vBwI3Rdy
5cztPPfft6dDqGiVyxxB7Hf2XBA2l2YlPvEEZndDnCT99Z1wIFgwihxfa6qmqnTW5lANO3ozz7nr
BHaoXZ/XZFyh9y2w4iWFkccDnqL2ehDz6w3YwN+IIkXmkEC5lVY/TVM3nQ7SVzQ68rP99Uh6gQyd
KSJ3e0WljzBQb7+suck33kRtqwso9DkuwZ93zejGjoAgLEjra0KEvypBJRmWUCR28UBgMdzT4qRL
imUEwYyJw0SmyqV0AgLC+jc3RUImISE5i+sPj6/qPwmO8jqCXfKRL4eUJJnYQ8r0hMb3HuypnfsG
DMizCiLQPBvLXDGv7zdcnQTr6NRfhrUTg4k5sYxWlt2sjOpF4Hh5rcr9O2ylGptelcOs6xf//WCU
BTGRJk6tcGM8h+3Zfu3a+zWwnJyT6+FrX9DdmnK8UeW89C8Bg6qhr//rvJxsJkB1uIBHPHSgzN6S
YIupDTmFj41+RH5BHVY8ZmCuxboS+JO5kwu5IndR+DJZyIs5OoJXxpFuZeCIB8ToM28i6W8F3siG
9yt+o0XBaPZtYUyerKZj4oaKEn7+BhM7YCAHYSKdwRvazZMRt5OWsH5waKTM0TkMuJfVxry2pVB2
qkl5IBC2ZqxDWTX5qWRNxcb9BcPTEahiUSPqtZQPg7/D1jbXKUHQOhX/txeOlbxQKoAAXwpFb2f5
Ni9Jg7QvaT3fUsLUzrowf871pVGqEdtacL9SKPvILng0OmGh4KPJt+Q1GR0gK6flUc23LTNmBLxq
/lc8XCm2TDQPBsVifQ5RxeR5D+kOgU4auPnqODAGWuLNWnOJZvajG7cdYZyJq3huz6CAHg50gZzI
2uWTS3LUVZRyi6U3c46ksYOhJndHDTm+R3RwRaX+ztR+Pcq2EmAq5d9qzKs6xEsP2HLfTjc90BwK
akLCJb6oqhOrFUvbBTFBirdwYOUJi0tVmVuSmS4CKy7RulunJTw98A6YaEmD61TrtOXN9Gtko/XU
fZ5+m2v5zRQYRNEgEhaFs1J31tzUtHyiNJOJQR7zxSlI4un9LiJGqLiim0YM6ZozzjUjDywUXhr0
D/HriropW1OYwQlx0Gqwq2TlpOv+He5ZnIMjnjw9XVNzo/BQ+yAjUxgZvuDkkqsYf8Z8K+B3xhSq
z5NWSmvAv4es5ey2j+k6i8NI1XYbL5iBhmr5FPbOl/zDUdfguiqQhr+c2OBH74/L2z2MXci7tuUD
WBzM4eMUGDD58Bn25TFzNn08ydnZPeoy/q/lrWD5o729yYiI5lRSFfCtxNj+aTYWqC1uw1w4I2fi
MFhJdLBuNeeVYfNR6CTbIKvg1AA+sN23DxDDAJ6yEDlgokKS+03huQfvymJVogQ9ORUy5u+cRZeq
HcAWR5uAfa8fPKsF/zz52HhxnNeMt/BGsS+Wno74ucv1HEUZwgsx/HGyaETxqlgujS1oUMil6vnj
C6F9V8HGBtZMuxoHGw4OEGTTucPjXpQSC58vhCEExt0fptln+d8sKbLiKulfqDSLn/I+P6l9LRqT
HDqd2mQwgllJY9iarWsShdWrIePG/Iw/GxfYKxTuSl0kTarvgXgjdwu0MHJnhU3oua2F60iwjPZ3
xnTM+hsU8c6lxh6GlJReTVte5Zlbqk9IBMo3ifUJiwfF2dqAksBmCVKQjocoPu31or1phL7S9EhI
Az2fLnAmx2hqI1qa9JEcr61ZSXCmO0xa60Bnek+cjlmz6NXy7Peab83E6DeocA38tUIllpt9D9IP
Db8/uU6gGQrGnpQepZd9s0I8+H9dhLWn8BqsiX/A76AXV4/9KrVVEt8LCyz4LxilvFSL3dwYJcVj
lHiQV/fjXvJewzfn8IJp5HZcKmqmzIBiA4wAJTn7KNVh/G0Mdy+lRe//JIATw6/olIOPKHKIBYdh
ulpkD6KUSmWgqLPWpgB4JsMBKmHKu83rYnAuEKSgwj2vAW0mP/N1ojWu12mZ9M364tLcLUCYAOsW
9Ji9hhpXktGejQUP6fYrpjJtDR7+vnsGSZC8Jl5L+6vRC25HXgNjO66U9ClDPwbNSYyrg0yA/Gpj
1lrxBO4bhHD9c1Ihowy7rv5EFVywmjCXrYIkXpbqoBgfjJFJuhNXP/BkS0j70Xxo4VDj0DS28PaP
Pr72HQEKammNHRyxmASfi2MDmojoN5TRUGWl41h6nwJbWP7dwzrclIP1/5JeNQOUHrni/+pHEniF
gcFnkDbXIniW6KrXxY2asqD1Z5XVVHkZZDCsDZAbF0Gv/wJE0KCj+qHNZL+MkYFPxdj37DkZk6rK
R3zi2Th8IwOHrLqwGL6+VGhwIeC2D+m2suEyb9blcFBRzg55uJvRpeaK/xqOPBz3Swf4D6MhJnhf
8odlAe/CIRuxqBab/kHqn9P4fki/eDMEkJXpObkUAI/qQBViPDUUIuMGAAninADcW/6C7fn/DTH/
vLDP0+h1bDNB6w5Ct+toONdXOxxurdLdnIuf4QAMaHNXKKfd+I9YkRf0xduDA0/EG7Du2n0FB0JR
IGe5KaC0oFquywP6tui71O2UL/5csUaES1WcCrauRS/F2gid/Ld3ouWSh8y9R8ckN8qTVmIXsT2s
A5l4X1JDjAj+GE4gkEediBzggV4oJp6g2pc0BX7RQyk3h3h6aGIUaj8e5GrfMRjFOtSip6o13/C0
D6OAj36Cli9Ub4AG3bGj74hPL2C52apVEcmNk7XaZ4VoRkRoco1Z/VtIsT/X+Z9HVDHayZYyexVQ
OJFm19Nlk8xuakR3W/fPCZe9GyiyJYA3W6mkKYtVuCkiwuSuoeJafOKVZvRe2EXk0oc9lstpshfY
MtyoVAKFGv1JUbBam+70HOe59G9JBUB0el3/MvCTaovZmkcZhazzbmdOrXw4YI1DPpkj783aqXo2
FDJ7Fo3aQqcUiiRDqHQlWmIhgvKyd7kC8+uckeQN/qQcopZ6bMfQ7pa3E04XtyhFU7GZR6u2i8uu
xvbbyCYtc86Iz2m6L1TDCM3oXjbUx1LL6kBpsHd1XUx/cpnebq4mCHuEKzZqf9uLKKtNjaSOsAml
auZnJZJtGbQ3cnBFeHdHp91adtNyK5JMn0DICoL1fDPf4z+WLnbTdI2fMr4G6NcSC2zNLEZtO8X+
ososG/vhUkASxCyhNii2MfEhyYtXiIdiDXhINlrF9oEY1/zQ7v8EQKyYBiI4UfqK2zNO4Xlw2Bbb
tv8cB9U+PHBs+LVMmjD91ro0sOjMkmB6Ml1RGBZn6sGLODNs8rOX9dPxtMb/VLBDLgJjTf9ukTNW
Ksx52opB2S/GQuJ6sy0zWD6X0LQ/jWAsx7ocH8LIaawz017TnLHDocXwb6XHrxBWDQMcVwWO8LWJ
Z4ZmS0f00NIL1e9gx1Ftk3u2pRVV7i9POJ9fG57N5WaTAH7GvddivUVq8Q/wpQkh4paR2LZln+oY
cGFHwjAsdEckdvAIxpEdo8+r1e0830/90lA+bnD33oQbevn1FZ+Cg+rPL/BX/QfK3I9ij0HHKvk7
HfWSfbHvft0FOQBHJe6XpDBcO5T3d1G/76jo2kojIlavz6et/LlUZ+74DBHgDBScLHH0tRx7q/22
URLVa9PPPTIqUPj/7B/Uz/hC6dOh/TZ0pHjqIrZ2N8o/rm1cfoUWpUFqU9t+4yQX7RYJTdE4nTiO
9wZ/sjJgqSDXznmZ4y8eIGoP7Ar/e9sxhCLTQ0PbC2UvWkuyqR+gtFBUL7WvwmXRqlwmgwmcxPd7
ZFvU4gLHhd016ga7tOobA8TWoECT1YrBxbk4IeKAsvuzBB50pxjd8HdxMI9ATrD6S/WKw6FcVCK3
jgx+EvkF3+ggCavsEsLy5nHNvw0ScoNQmfMDFpUtpbeWOqisC/FeOC3xNtplFK/Yq9Go9H7O6xJe
+IolLmy1O41BVXCzzdx94+e6JHs3SKGyzeuRF04hI1L4wt7XHqnWmx+EuiNY35JN9q0I1aTx+Exu
sMU/dZ6zRF+lBkd0PCPhrfW+cFdMj3oPxHOuQ+rxotMbLqywE8HILtGrYWb2fY4NuGhX4cpvBtip
rpi2BniG5gprwT9RX587PeukbBxsXYo6RiMhlLIB4QaJPzyf6bXz9qMyh6vSVcMZ/6GpxcQ7XUmV
2cVGTtgFTPJBSF4GZxB3+gLuPlJZSmrVZiOyIpkd8GWkKs/HFufga1Wfm4IU4IuvDymD7uQhmCFJ
iMgNGZctEOw5gUd5DH8M/qE8WlGt7fQzFCfL8gcCYT2GZ/OEFoYrwB2QOqsbXY9cOPXcN+u4i4Xa
u211jo64Ow9UH/5PUGSMHLeoiaHgTXMIyJ3v9XzEEeY/peYd9f+Mvf34OQhBF78EpXlcLtKjJsqa
lMgObhHPu7++ZGmB8TpoEA4WieYRy9eF+jw5gZcHqjrLn7iLMznDJcWeAM+XGQm26OiMBvNHHrDl
c7r+YIsmvszo1Su1EI8qGkJQdNC1JtDUPgolfSIUsFZ+0WrsXslw0LUTOsQEyhdTKztjv8sVRkiC
+0FJPIpjC4FIR2avBYn1R4lK+ovkvqRdleiUI3GdVnQ8nXgPhYtJlSNyX7iY2BN7iEKnrj8ineP1
97YK/7SdrDHDfhPdMEHBLGbLu8Ojc8OjLSXD8t3q4FRy2iY8ktPW/pcvwtnIoCf6Fxdgb1Jksbab
ohaf32U5IyXVtUN5eu2YSiqNN707jN3A0UXOL/vqvqN1TUhtF3tMH9h1S0heRk4buBvcmeBtKWTM
kBWnmkNBCM70ZdV5ikLAe4NF8iKKii/Bk35B9qMa/c09EffwJ2oDWfCqVyI8ooZRusWFOtUpnl7l
40G8HFcEV6C26ucePO+Eaf9HrKaSfy1KTY9XdX3ZY62WGRIrRmooaIFJB2ga27HBJrHTiMhbl+1R
VmhXNFqNEhSJY2YgYx+3/3ezOOZ7pFTa2Qm96LGbtKjwr160E9LQi89Y9rQZgmSS/27cY/w1KhaC
84hVFuUpPHls9ywhvfBNgJ/+uowl/F736+RTAbNnwx2qy5eTYp5zyxOJ5dpGYG7QH1Qd+kLFFcBT
RjKUx5qsIvLmuYp1HBLHh1ICuERKb5iNeKImAqj3mGPfP5UedOnqrOszuEoUzEQsF6XiElzkwWdF
IfqJqkfijruJJmf8Vu/5ue2a5ha1hV9eUhFAdWXduYAcKvMCnrq/9vzdFbMoK4dS38dmc9JJjT2C
0Dim0q7Q2TpcAvXCks1bc+6Dk9VkMMjzrOkp+A1PQnKD1sK7dUXr9qsn2WppH8J8Bt3Joylso0q9
abti/8upFBLEhYqpEwlOWC/kL3ikusu4JR3M6lvt7JHuPdtxo2SBHDoNDez2xFnVoQfropHg0sqB
xnrSptTT2m1XKfrfn3uA1xD5qYPsZNgdolj0VV5RuuuW32zIJ+M4DmQiwNb7Z1cVQUI6lV2WjYUp
qJnJEnsamL9EVvub9PbIEa9LyW71bMvSvTd13KSsn5ytMwuyy2J2Zf2XFPziMyH4G1L7uunlfQQ9
JSu0B34gl8dOVa3NQerHmpW/JNiHAksVUdOktjg4AVqfISkZsVTZ9rBnJ2L58MkpVdWvMemPuO4k
BsDU25cRt0EdtkrEx/ykQEkjAwPUZXMXRrnui8wkOPfxrHiCkHlPvK1Q7jY/KBEoAVp38/15JGjp
ah9VcOlboqvT6loyydmszrbUY7lgiKpd2snkkc+Ip//lu6LzYV6N7z1IPfepGBWzPgVvVmBcYoeP
tNl7VSNA7hwD8qtmDIfBMnGiCU7WO+XD0KKrCR1+TSfNmOXo1reB2Xo7aKPUyifoNTfKNGdV5L/R
7yyiqYuMMWHni5YO4xn+kyh5088T0bIFOCYT0GuqJjgARR5MaMvCs9uEb5rSIsppI3CHkjYGAXV8
ttFFbGWDbOTbi3STnTbggDdx9yRRluPKrIeXDGJamlwDVOwvPZuGfx2QRfjgR6Eq81wFKNWTvBBf
fsDCVrJp385kbjHjFXyxiuEcyDCdclGDz5vK7/TiQKjcUfaMyK/b3qstsdyj09rrX8v4PIIh1EjA
Xn3f0pRMn8hjnUTH/enSrtXa58koA2ji1XOY2QGbmGOVE4nU+/PHLqOAD4+e/racO5DdYtegapTl
DUDXzcReN0alX+FVrMPUy4qoDXYuoQ22nOnbH+/gZaYPWaqMXGNghQ5q5fD4UAgtV6y4dQcB2Wbz
swquAYrON7h3w5PjyzNov11lxER/DgIY/s/QgF2Xj4WIq5TX6XLz/+Co87tqSSBddnAN5O9UjJAT
1AsE5nKBUXPeMYaBvn3xjEkg2KFM3sWI7ax9yMytqTK7Fh5U6QCglY2E+0j7FLIBcPIwe0h3DJJV
PSirkwxjoM90dlwTKD2X0Piba2mwcvX+Bj5HnDZ8A3jhbeTMCeHl3u0x0odwGYBbUBbKpSOtggT4
84mQt1ns2uCi08jzFcBEcfhIyz+L2w/MvTkgGqVcjnFZ81MRbqvdAHJiXSjCF0+XU/NSErSfrJhx
BpLyPmbgnD9/PY7IR+9plE57u60HtfLAvqk0HXlEkpW5XTJKlvoaETBz9UI+WBxvfJJCKrqYxhpm
Vv8+wjYNo/zseb+KYmxgPxu3/MAimEetxnRjwX9VHTJ3I0O3dZNFcImr/LEN9bfEt31aBkgyRd3C
9cH6ZCGU+x5H+bzc+pwlZ5/ccfbVCR4hlDGkkVbV7TwPLORC9v7+OsDK8HZ5d6Jletn+I0SYvULX
70GXfCpLZLo4bOQAD+HRUV0Njv2xqWXzwPoWJzepWvY49oN14otf/zmaJJ4Q0XOlhJwFgvth5W4h
HPwsBfvBb2EkKb3P5Ghrl9kZFzC7u+HH71ni6ifUJdVLBpgUmHS9f62OcDxzMLTxPTJnapavBka8
W/uR196O2NT39DV71jlw4SIrFlnoelUtIVeYCrTLaWcOYtLerFgHF6idlleFM9jiFeiVFcyykWQm
/n/Pr6WOn8m/FeoLuIFQO3ehWiVrdIEPswHHW6+GTpIoj9ZLhPuQQT+pmIhgifzEKm0aO8s8q+xz
TWp/whF98b5AGk3IVk3/puiQ5/ROxfOX4seCTLnIQGuFEzJfTncEWwlv5Kvj8qM3VAvspv8ypNqb
f6BTXJ9s8gEpdd3aAKDmW7hw6bS+s2Un2/nzUVsev6kqB2NEhd86HBPQ5zuFVm0D2oyZgS1e1p3o
abuVo4svlZlc+Hd/jSCndly/6x3esS/oQ20KFC9eDwb3GASjNEVqteEuvMGjhaHAGScxOxSDAeRU
cpWt2mVPba33b0vUxAMmRRFKbpiYyg69YcCkH4W1QtuOvlJLd/G8EhrhK3vEtXHzRuUeF2giV5gv
9hls9l92yEUpjZkdk1XpkKU77GQgH/LCf31fF4AG8Ed5l/d/Tr2DNflma5vCFwmYcOOr+JGrU+R+
ggIci3ZFBWyMqc+O8p7DtU4d4A31AsKlH4LsllfxgZAgn+dAOYm3+EzSQ3KWhkuI1TgwX8lH7EWX
5OoOy+xe2J5l9NE9faMyqvg0wcSvNvXu/UsaFl9yI+BZU8v+JXJIo6rMStsgBe4phm9V4KJISN/2
PeajT4bsx8PrKsX2qRdHUIRbDMF3lGmG/oXttvwhzuzeRmMvGU7irUGci9uVeMR7wZt7ZUhWXuhp
Zz09ru8lQtt6KLrO8Aj2s4M1C0RgIv5j5Piq12K/acrEtXhqvMHU15vt3sznIOuMJvkWIeSJqYlO
DiqxAeAJBDPRVH2aZpr0swkEhc75/6QSzTcW+bgGD85+zIYaKx/QD2OG2PKAAqIp4T6RuXS7BtFf
0eH+HAf4nbAslLy91/UCbDMD1I7FUO7KTMoI2rVyPdZ6DGlqeEQJSdbnoWrFLv8YxkHzYM2BxoNa
zDgfQ6l25AG7ehUtKqeo52LMWPPJtvCOW/FIDdYkpUUQaZPcigMbbJXk8g6QBOS/D+LzCuVqygYI
08BLlKWPM3lGB+3wR8fUO7Mydk8AjauyUBfnE2FYJfb2yrWBIbeW5+fgBHGuUfDFtjKKX80S51Bp
dXkjhc/v3BnPEYzy6vE8WNq1qqM5NaOXE8C9aNRpyTSTXxL1kwS6FO2G6igjnac69OGH/wut96oW
F7NqNdFXzv1bnpW2OdT3RGB/mrt8cmIGWvhBl0m1KGtzoor6DWyCCPEsaqps61y6ftuoRLdP2DUA
Ba23ifFwh3OGlRU6HoU7/s0X+d/t0ugX1BlUuGBEQseQSlHT5CRB0R8L6ezcGZ+DsDTlJIO80BWo
sYMT8w4ftHLKBiqvBXXP9+NY+eDOexl+6KbQQsbi/aXu4idBgHSCsX135yjhcMfnrRy9qjoZZFA8
6Y2HXBuxJJZtQdS3QjHC2dzCXTcMf0f8+6l+k7FHY3YNCN3fxEYMx9K6rEh/r+4MLfgvnq4vvDgN
1+zD6WW6gwr0WFs6nalbNp/4Xbbcmp+OWfMxE6pHC3gjbDLAuWr8D73l11DpTlEKi21+1/4DC+RZ
cNodEDH8c6zLYI7wxC2C1OomRR2LMLokhaD6baOIe7IAKjx5heCr05aeMDhq0KuVZmbzSeO06CRu
zaHUDMHaL0IvQSW8qonpo0/45jXTsa80tWt/Q31L+WIAXM+ElT7yqOfzrXMYQlEaU0r5sdl76XzI
GZz+MyrvNgb6jmyneE7PFSopixkrSmzJ7oifdbsg164yaOqspdew9mfBjdu69sgPEtitI0DMprdu
tUi/xFS2jmxgTwMjb743J0cD7onI+qxy0lNoFLdCy9myDE3cfQ7cmkuPQXFkw+x3diAXHHCQc1pK
wca7FNYuw3E8oBIpequjvHrMfAyysTkXAZ0pzjUbrOvRtshVNtVK5yeT1tYBmjZjZhumNHHF/zNx
sE3gzFCBR6YPZZ+G2NUQso/1Gjo+bIbiCPQzYD8bVQLACea8TO+6Y6ahpNRcN28l2DuA8aIHJuE3
ZevgC6rue+HckoVAUTN+7Q6g34NeFL4VhpzbIfcktJdsdo+Q90FNgt4sXgxIMQzsWkbUDzQQ7KSu
+NhhLPjiL2KNp5W+eIg8TIZyJZiKc6TnCf2ZEPXq0LEoyJ198ku9iyBEiFEo8kDgu/JbwtIE0xUl
Z+4exJKN/9EQsIUquMmUkDhahXzJPAWC3hMH/GyI7w6NSHMb5IVKf6INfBandgh644OsmQ4fYa6G
Rvk+Y6AImTb2e8g4TzKik7D0OvE8y2OGx+anKsLxGMPW9C+GJWFxN/AYf2dqaqMlitrP68d8n8NW
qCRMaoGs+bY+bjru/Ut1CwOAXUPmE4qzxI6u5wc9q6u5tUFU2ok6XBFUD74+F+i+e8xSFF2dYzKq
EKue/D0WZSLhi0hZtioscQuEFb4VEUSaMQX42RAAllqwxa7Q22bR0C94lSLMzzVFK3I97cYeF3DY
Ow39tVA3YPmtCIvN+QHx8vWIY2fO0SxjB33bTHRT5b6ncXnkoY1JUuFacsGawWkS09pdeUw65GLa
kVjYj7rWC4orZ9sDqGg6vqd2eFkdhS2AyyYRUCpMW4zN4Lb5xtcm+6tyXPACcqvGdBm99I7QouPn
J2QOyo8ElMToY5Kiw7fQZIyOod/PNCGfGx1BKmiPnusDfpXe7tRiaL+H13qjsL4IDKzU7RkSDjc7
sWtjV0BzwEPUIs4EgKpdLVcc7eNbGzSaTGhPhlS/eLtFDFZetWcxtLrjORF79uOBEEDs9JYhaA7J
7KI6Tf5hmS2ZQjmxQIUvJGxoAcoZsi7uUqH1E3UtBB2P0vvwKgwfp1H+uVGNjG2HCrhgniMsZTl3
1opt4OEQI9o+Sg9ZwujXnGLGZq0Fp3hfm8L6vJKPh6LzQ8UIh6DeuXVQlnfWXuKbnwSAGdV/KYka
Ru+ZeN9aUb0nEExj82oLWcrCicIBo9Uis6gFALw28NbH/iR/34nkPMs1KRea5cWuei2kLPsAB5nq
RN2tyZUVyqEU8CWjMwDDRwgN5hdU7NoqlIK2uRGZJXVPh4wxpaEOtezMNd1WI4qQI5PFx/FZmqCN
HOndYoCYZI/AHQB5lxcjbcTpF/ShOQiTv/mFRvLAJdIg9lVZA4uyXGI64DqBHJSHZciwXXdj3ij1
9B9OU/peCL6MZD2/TgxAt2H/eT/BHXB7dDHlDxrTV3ge+ViAcCHsm/VTu7NUnxtjnfKrx0KKYee6
kLAGaBuAT/xT8+PBdGQ+0XE61XRoZ9GPc6GAbFlGpG/uIyt+dRO0zT9rfhDA0R5XR2bfQjzR7bIE
NkhvFW4OhNTyYzFS2cv0r+XR7zk+NIGMcbDCHxOnicdUFIhgVwImWAh3u7U4agMIdKprXpVeRyFJ
9Bam2DngKEpg7+s5qfXmym9nQpLQH7YNC1TDBpnKu5MBLFd4vX+ILQgpSvTZJu+5ybvq7N8BgsAU
C1+7mC1QBrYAMdZwdmTRC9BPX4U7rE3z3MHbjpQ1NZ7Nfpn690+bebygwtx+smarJRJJUIc0HZt4
TxCB0sdL+yL++60j9O3nMsmaQwVkwZXZdHfGjxHoKkETFggT+hr7BvWtO/K033VSmv1P5uhRMBIa
SzeEf3CPhbzA0VsAgPMC51Nn4tACxhHsdPpfQpesip5uSRsxo9wbk+C+Hapi5nnZjT6MCCoU506N
z56nkmIUn4TT67+P6jsdUkAOOONuaOE3vD5b/pISv+MkbPtRzFxH9cuw8CUsPg+PKWUTE0qnNASr
IdHOsxJsZvcrOlutogtMpA6PYRIH+vldGUT3/w06vPWjj0Kdt9N73fhe8t+bLhPOzoTBz3eUy2dV
jer4QxPiZSKa0Sfb+d6binQvofmnxRvec0iNF+Gk5pDWvmtV11gQHuYJd2VwDs2BuP7/2OLL6sam
rDGkkSG9CQmfny0MUz+Bpz5eYFrP20cj2ocQR8XTI+vU9tCY9LVBfmlkfMCWHKVK33uIOdN9q8XO
5ir3sHBxVujDleM579v7BwaOhEHYcEpMKo2TgGQ9H2awyTcNtmIULWENbqAlZcAKlhrE4sgARC2i
KrVM6sIgKsvcUuqnnZPQD28fJwFcs5DgZ8/qwCOcdu2fJ75IJfOh707Ur4XaBVQlKhMFvPt09qqx
0MijB4rgAQaZ7d8UVaMsfAtehbrsuan6POru1vvyPDzffRyeSfQ96x5TMvrslls9ThZ/cUFR3n3K
C+onK/2xaBiw/7fgc0NCoxOysKTYI0QR2fXloIjf24Zjt5GInbsIMw6Z6TPW8x3i7Cr9LOW+dw92
wfL5b13qYMWbtWQjkplYLACri9gy6kjLDj6xf1B+OehdVU9vqcwGrva3HmGOMbT/xIpQz2rFETnU
MiM3YAw1ESBmz2se7zQHTUzZx5Fq4g/PzHh8GDY9l6ykU2MfjCF6aHJTIMdrkgA1QnHo+lmddijf
4JO5iqSXq8UYA5W5R4Rtf/51MAbhqkbUMPIDmcwtP6Fuc0Y3OfyWM1eoAlkeQSwhStdrr2kJiCzS
ro7BJ7aV21wGpt9IMcFZnGtwAVoipgCz71Fs3B2nxV7HBGW/rNj27mAzR21bQeleE0oURrChtmBb
O4mlNVK8/s5qTxnhjb5Hy6gYvVLpAy/3hj6xnviUKMfnf+V2QUWkeNeD7DQK5DcbKeU9fcIusHni
aBREeND4rseVTpy7+K9yIkPaiyW3agiiZwsdo8Mn171pAZtcHxu8u1isP8XnOFVGS2h1osCQ9jIL
CtT4aJFL/BpoAZTwC4Bn0gaeKbHsqESvrh2XtyAQqJSdIZpnkPJFDttHZQvhculQ9GRAV1oi+wbM
eE3DVY/PU03p7lciAD2m05PuyN9Ue1wmGq0Zqac6LEEu4L7BBcmVn4ElPQswue8SOuKrAe8ewa8w
Aa/7TUdeYDfG+yPinrzjEWUoDgmlkmA7ofMZNdB3rjy9ufXvTVU4BKAJatkSf2L+xmYG+VQ3oA3G
JDIGUUF5+cGzc/wb2DWFrW9sNFUCGOYDWSqOWRam3XxWc2qHIBPnFh9D5u4YfnxU84MpMNAuw+JO
91H3TgVuG5Fn22XVEsasCbuJ8rt1G6vLSNf9PrsKDRVq6ddId5JiF0M8SIsZBNZLAmFVopm2TMx3
EBq8ujsO8Yrkfy2Pd1MDNYvjiv0vCnDa9qVTiYILvdXWxkGHoz6YJKwp7qndAFJG/r+wq9QrW3EM
TjMNNt5w9Ap5lOQQ7GY+vGCQnhKmkfhEeTP/zoHhCe53nwrQ2WfrRulN9AS5ZgEsRcsJv/EYVkg1
9ciOoJQ1ElSu6WbFVHpI3I9R/SKc3SX813rLiKSY4pGq4I81fb0uigJ1TO49IK120M+9bWKo56me
NVbreaFZTkJBziQjQ1eMV0xNsF7RaEQydEESj4NK4rtmjxiRgeAjnHy2ubxvV/wB3ozEKLtn9p4g
+neFFu08nNcQbRnEENNwotbWisBjKXO1oVDV7JIYa1eLvhpod1ffD1ocLeiQB3HMTXEknWvOQxGA
1sRoV90okQ02CHAc1A82DxtSWgY4vb1/K9Ux2UVKcLIP2wEyXiCPWLwE4kgipEZpKqO7DwVdxp/k
zSVX26Ex0BA/a0UvNtYBbkStQv6Dz3XnASRNDHk16VTO/xB00o//3Y6c2wcFMat0tf16RE+swPx9
nKphS5RbmOcDgObQtBRrzU3EGLTSy4xVrNio+LczaGuOFvhUYZmRD4wjWlIDyNncTI3I46AnaadH
daWjjIgoBck9JYQRdvrD55n8fhNljWae6mOSBeyrXuWzvv2atSnydrWabAVsIV0tq4owaLJUeuGu
og7lBcVEIu03HFnfKq6QTIcj/funSCOD5g3NTOgSve6fkCC2HaEkQnBbPNurkvjzujPj5g2sr5HI
ae7N0cm08q8HGBL7sq831e0+7BrrWAgd/GCIhZ/YwCB7v1mdCj9VckFnqfZ1thg1cpsWz6w1d0k6
Du+YHgp2nBUPAM37AZzZ3koldlgNtJoHikFfsqxIO8IcIJk8N50O7WmRaPrF8sZTrX0tKwnFZHmH
fSsLzve85msX22WV5A13Y9qdALZLEkGXIetalm776AHdESDMORQbeL26TadlMNMGNv19gnu9MM2W
lQByodOl/99PMCaHyMjXBNPa4eHhs09TzAGFDrry0wRTsDZvbeSAtctBs9an08sWRNl3+WjmuYGE
OsdhGz03Mz3UHUBCbv4HNNEnY51bKJouyj9V+IcF9q82g0zlVjDS8o1z9foE7zlL5a/IAuYCjfGU
Nhd5N614AqIax4U9egXj9ScYEfjHGAoiusFziS1ZxEW324cCgFZ7Ops1iRTRMaCSNSgtuxxTP3j1
fEAWgl1ph8BsBm2JcMMuyN3hMfTwm56beUSPlMZf9jHUP+Z8PSH5LgHQy/vJewQg40m62hz4NGBk
NRvLNW3ghe2j5N0bRkFKpzX4wYfn4WXQLJUe+wYpjGyR91oHOrEJtk0JFsStqSzWjGcFjVHWok3B
4zVeXsWB2HjQprYQ4EoDWWraEpzrds6UtwviXtdOSq2znhF1uzvyoCSvbNMHOlbeFzSX6Y25Hj6j
IECvY2u8wl4yJSyT5QfZa8X+FAZ4nxBNkS1X4uwi4klXo7PWUyf5tJguraSq/0Yv7gLYEQLsxGbC
2cWmhFAphRJUc6jqVHlDZRMowGkbWMtrkC9qR6gY2hK8s3FCjmA6BVZBDB4vwyuVyJZ6yYYtCG49
GHO2zUT+UkaYf0eBa1DffLvH4MSWB4zTOYTKtUcX6a2bewbKt4Wn1ZrETX6oL0C10197NMtQ/8kg
mNgDpbpnd8XOZV7QJh9Y5iV+TQQ6vmsxbWOmTxiPye4l0n+SDxVn5oml2zJdVuZHCZc8tgLUbF4s
/qdzHmBLnBBE5oiiA/oh/U2Yp9/2Wlwj6a1i40gMQj1GQRTA3rloHYF9fSdJ6zR1CKvbqF5r4RTB
6xhtjextvdJ7cDhQv5FvZfLT4mt0tZUTFxfiSkTmyzxK+uwfgsBOcYDuk1uBv/yJAXRldgDx72rR
rgxUa8W50zFVio0zMa0FzyFVcl//PdXL/WEku8gp+kfIme8r+YMIwVNZjig/y/yEDF9TOlz3ghtJ
dkvvbg1qJcnn6rCC7jiURWOHT6wuUGX8ICGcmxkIw+dIGCeEkZp69njNYI10h7PjlRZMP2ZXsuYu
Hyd0EuI3qNLPPWTEyP+6ekxoWE61Egl6VsbpuZg2SqGarVH8u3oxbVpkmZ4PCdxvunTpJxDo5z2l
ioYM2rSwhRZ+VrZH8kiKhk40LFOTvZjTfqf3NOYRhav85PJrVNxKW19vd6svm77GTaa9jnqjthoU
ROkXBCZnAmYzQ7iWW74OkJysYJngl8jOsYDDkz2DEYjLCmVQ+b8fLHgGw9QJtYXzfqxj+FI+nokU
dhQVO/Dp3TihMXJTdXKWX+FgIj9sAcCEYIMQJTzicCfIEQ6YzTj28UT/i4OFo2y7llXwp6AZ/3SS
TI/RqrHnqKcgHmjDkYRSLLmUpV8NwS86M4EqloLtgCA7qNj3UC57XQOQJF67yz2BaQcZz+wv5JG/
cDVyrQfrhVrECPUG/6P5dOuI16kFvYugRqj+NhHkqGB+6Ni2LQq1GKU4s7f6KfVdQ/pMR8tqBxy4
2NG4FCiRJvIXWSkTbjvuAS86s4XRLEXDJ1koC8KD5LVN/UjDV36oBVSbpFh8GJCm56UyXyzmFDeO
uDi1lKiygdl589MxTK9LLStJqyeD0V7KGlPNfG7+NK7GMhdspY8H0NkYPqwCyP8KxThilHhToRH9
8sbMSlO7grABkZ8kHYb5g/PfQ8pbUwPuqdQAwHbMt69x4P8W5WL/2FWMgQH6wK7MltmW8tR/5jid
6WaoXnynL+LFz1pqcMX5aJeDErGQgD/JxhSOeNm74EY9ZI16bQTawjPBEVyBThT74fzOqEViM+to
B8RLunlBZ9TwC46y7YhVp267guoWYBj2q0YdCu1Dw5eF8s49krimV+3221nhSmHm0E431CP7tOZy
MufNDnt7JAVvHMU7Q/9i6nsMdaNPF0P4tOrqfrCglq6wowkX/ErHtd26h0FlLaLyWJoib1zvZhX1
n/XirWB9hIyf7lyUwWdjacM32mCQMDUofl5K2yDayXcWWmjJj3kk/a5HfVT19me4PeAD/U2U25hR
jSCOZdpGp78WuG2jK6hUtJteowevWemOYY5YxsfcmKaB9fbv47a9Mul6WbsnG3xOBa1Z7gULyEN7
tgrhOMgWdYZoLudelk7VYqql5uxPlq941gSX7spYkIgMw9G0X0omzvQxVULyODhLzW2H8ES1Mci6
g/ZXdM/R7xrPducLtc13YrRz6kz5SjWdJNwvQSpIBWkwFQmaz+KTwu/n9bKthNZ79tM39H9j/yYl
10DhPkxx7uHxanoqUTLAWy+B9jwBIQPccu266YmeRt2sjIylXieuw5r9R4h2fVsqtZhwN/nDYipX
tlC/ruBJB95FJJfJNMgAa8q+Pc3EDzWgDckZJHGgcx8i95yglJc9cp0GR6pITVdd8jHyDbHC1Fob
OcTygxS909vNgBO4vn++UL1xtA568ec1pwjqpBttnL/NWBLQGQol50nto04/VIglvgCXv6DDC+ZK
Yv9tIYxZVvpcan8vYvqT0zIfBgVq7MNkwhm/OFAVM2HgzYgmk04gjxbm0IFChi8ALcosQB0e3QcI
7xycb4Sft7OnolE2i7QxKt4cfhQH/Bkly3pBKXYb78XCzur7Bw+p4onZh8gGhBZPToHPC1VJiAlW
IKZX99zKTPR7xiODFkhOo3t1JBa47L43xqCScSJhj0Lrcc4KfgVXRZiorIJQURZRzp/7pXZr+DOn
PMzxPYn6KiwtXpruCuO6RgpNPCE4YWP40kbFczueVziC8hpi3IdErD4vmgQySaYXOcifRJzB3G13
BHslBfbQ+6X7/55PINaCLak8yRRh+e2r6Z4UOlnMf6nd/s3+5tivuFn2Xcao53yS2cYj1lJLf8Pu
GIn7C+Rv5KZ7tLLOuXOpf33ojW/rglarmuEfOcPkJLxpMlYxBfGLUvR9FVPqP4uH+Y/eqM6TFmFj
JNynWJTMbVC0P9ctJIWzmDktydr59Ck0bmnq33NGRBHokjnNbMEQoXMlnBv+6K8xXNOOqT4O1xbW
dH1PHX1YCsGMEWcFlUSMqNv8irCrrzfhZODr+zX+7TtU8jVTqRXNS3MezzXzwJDJd7PJ14R3z6+l
9Z432Q2YXjLrMhrmuYZLL2se27SaNXQbkNGAt/1OXwAGqGmLilIPxO4pWPB/4ERdYRnyXDwj+Cyw
6H2zzhQuNY+xVvDsKEokzbjB9XLN0bZAX9CJqsdzf7jDdvnA8x1pEDEL397PU4euDGRTEM7c/KTc
c1PhuZzKSyL1EB2zH2rPB68rkvNPInCS8/2ueF4T+jkKQuMws5DZ+v9hRm9Gex26v/ilDdirMQCZ
N6dbC7T9t5IR8ZXmbSxBJICwn913Hku5nOTCcVDtHDfNy1Il8CbJjFDd7PAfLGN0Us79lZrOck0R
DmfPSD6n2/2FYtFHDd3aaKwGEMnKnAsWMlwX5nhNm7gyp8dj3VkiyfMo6F++PhFihi004gCMGbZ8
eXt7ICdid+rx5rROhRjM2WB0LER2zljyGH9T9bdlTvt0ZQEwkkQPpK3AEGuwCufwcggkOkgghU3o
WtidAEeBjGriWwOrjHCuKM1SwM/BvMLRemMPcALMcZfkiJnEbTBh1NpuZAXVUcY9b/Qn4O+l+bms
wv4sBPninGDWXPPxme4pzVaExpVPeIa1dzZVyYg80ZFdjktjMDoN3LT3YlPy4Dd70Njf2Pw5uFHe
n8a9T148bnHTThRshvA4k7T/GFrI2Tq8yxg8/rhMLg5PRjZiOOprE23OxXPT6kWiP7gv3xyBFOcQ
sFvCgKrSa2GX//WuP2RZma+H2fAHxeCUT5nIK6ofyr5vtnaEJMsfSPRcpIetLauXE/qZXIGrUBbv
5ViCD7vpNV/Y+Ir+KjkMOSFAVhN2ItvXcO3FUo2CTshTxUQIE+rNMaO8U4/oiyC8v4TtRcwe1zxi
z/NNxNpgAgg8ZbgfwB7cf0r+Mk55sf9ziXeKTXm+7P8QONmuozYfEGIJX8YoGCDzlBFkOULxRtSj
nO2PcnEukShoGBPnuDs+gglzjPxRmLy1gLxrmi+/umh4DvQLrp3Joj//ScsVVH4nLpOJiAoFSwtV
pkXhm9Yx0j+suS/yuypj76e7ZX233PmQNbn6oPICU5z8/VLeFtrRS+4DiMwCvAtg90s+OUY2fl/l
qxZ5N6QMNtdzv4cSvZtICCSlhHTOFSsi95NiF5nb06mBRdEZLHsSwlQfuHr8SzeFglcsJVOTifQb
DmxGLEXMNDfP5NMf8bs+CF3pNcVk5saKzt8PwlM0e2d2NTAEqzoSzm+rshpKNB/THqgs6oIYTHGL
WGbLdbBSKeHyC4UEJ7CP0spzJ8lH8QIJIgqAIv8S+1QMlYXRV1GvFL6+GowAcUtj3zx4YSFTedIZ
LdmY8kFonP+yaPLk1blu3gSx7qI7i4t7LfdPmMSdtVJpgO0mr4AP13091MqAbMwgZ+CTWcmzko8l
csf9tP2uuwBGtAApV5lfWw5oYqVpmQIu1ypnED/Re/a3NjlsI4WzG8lWz9ncVtAjLG8mkrUXZs1+
ZKJmNOQQewbtUZ0xzF2GiV/OKZviAloo7r1b8SaRYkNC3DiifpiItDY54G+nHIrz/s1ECH/ARjPF
QHRRYdHZ1EzRbD91HjxWOPg87JCTpjxs9w6nb+EVjACmPmgcBcOJQUDQO94LctrIToLqvbJqPZxb
MzezW7RLiUVNK9/RiRJmjF5CaWHWPcloJ8K5N83lPuOXMSiCCZFy8HHAEpiNj/vi0njegDrftNYS
CdHZxhHmDbQq4dH819KQrThy05lfa8KqNuo+zK9oV/v5LmOTLspx+/dKkp5IVNVUqDlwaeHZAkMi
23rK/ZxK7dMMtPMyCkrJs7Nq+4+Ptc0Nk2NRjrqS9tAZGs3yl4x+jCl51esWiOI5yN8ga768Ct2M
ATiv56AMvf3bBxEzdkGavrdgKAYNTVhC8XbzIZhiwRtuuhBjSSkTB5wu4RGZaKgj2IBjNYAZatSN
tgAjdFNkowbxC9xTLp8mzV9NE74pdU7hsRhIOOiZZyfmnXRvH7t0LkaFwHa7jYA6sdmtxb6qa4Zi
CQoq5yitpAm7hzBQ6HmPqK18jTK+Pvp8TGQ2UJC5XjxjRjFCvFSilLpr0GD3R8IigNZ4y8qUstWI
z+BZSVya2lkS/LvUwoC43NKzrPoO7mVbA24Tv5JdCkuf0FjGYqbg6/IXO6WsoAub5WAZ7MLdJTkB
6XOFJtWToMWt1GaKAcP3H+kc2rsC4W8F6GIYUTBx9NS+FmBjeV+dpZL9BRD3MiysCWOC9uwQt95V
FdvVwOQFGZIKsU6hG3X5LzHLosbEYCiBATS9+fF4PM/Zwhhw5/zvAydxmnP66VIA6gFlnJAePV+f
dpZbJV0s9K74neYirdoHMOwDXY03KhNlfQMIsCOkk7gLhPFRnlqMxxoSBVhyEjKlGJZ58kjVBy0P
HnX+xo08ZLO0+Hgfz54cetILrkKKrR3QVYSLb4pfYL5Uh4oAeJwrFI0MxzRvi8wVcD50bJwPN7Fq
3xwl2vlxxDg/WzQW1AHDNlp7W0qth8K73RYtgNarzDh/k4A6JnSvDKnzsQJrKA78icHKtP0t78i+
JfejMH1bfoWWqy7Rg9GHZY8KOcNAxTY5r74gnddJ6A7tRVyzd7e2o1G7VXtyvT9vFj1476Lzy+rp
6rY6XWpPM0U0EpxIeMq2kKuYhweYwxI/XGo9w/geyL+AUH2S6pka41UFmbOyupy2/yjRdRds626v
24HnlgR13NlESiQ/50UzvS6opoc9epdlUQQqmJPeWhBmjTOGEWMvg0q+j1tHwoDWrfUQmREnVhkU
yj5ZV6xOXUWFF+Lf9o9Y4lmTly3TfDJ7CqH6hthp2xzkrquXwcecbk4+5s6Gd903gqENJsNd9she
1s9jXPVwNVjsajatHTAA1rsyTae902J3t1cE1efHCtVnnxm5UJYGb0VQRK7uPKAhgW7+8WhBfy75
LizT1goSkVSxoRXUwL4EvoD5IXEC/6rH687C6E5+x/tgpNcAvYj95HI/4aFOH6Zd+27NKXrejVhv
DsXQLEnwQeDdgI4E2G6IjpbGkvu8y1Wmg9vCfjaHUC7g7V2am8SRERY83UnfBhw2xKJ4MVUZSzge
lbKqcBADAdyZvQY5VdrZ+FmV80gttS2BT6dD3rNNvaxz2juEHJgqiYX5z2jQywiYjKvHdP+5KlvA
+3No7bK/srzK+H3XZiSICGcJqEDuhe+zMzU65NC6/TPHz+W+7RB+HaXJY49oihFRX7SXqdZqn0f6
urAFLHwVpw+bwS+/xKPWj3nm2G0WUIjBHjGhhi2BoLvyj+GwuP87LQaZUWzT6MUYyF6P5c2Xr+V3
/0J7hz3NMysm+ao4R1nWqh7YHb+afj+cC9XSZseSIAxJYsYz0TBlx4TZjHJ0qouo+2zebV7wAxFB
X2F2JSvw4JTCHD01BDzv+hS3mU/Fn2NghLGDW2XrtR33MravM4+Qb/7EY8LRKBqtk4UAksaPvJFe
HCPj5mZtcSw2Ivq9vNPgLKTlqTFS3prd8VR3vJNJ1Z9kRqpA13pI0Na6GjaN229B1CKjYXtj4yo3
3zClF7WP7HNi2mT6kVc3oBtjAJ7fQdIQREALfo9av+Ive7io9A4Ni8tesxbzCo07R2ij+Fb2e0o6
aEHWSqw0B9v5G9s5gLtpG4eRq3B7xyPdluQpoeOcATcw/lFPGjuPcZf5Qx0Ku9ZcbfyjPcSP8BLQ
UcsGji9CpVfj70QaTvM/peKx78otCAq4UBXZXs8xTc13vid8v8GPT8KH9qTBiqONLOOwLWYOu4L+
GSAckOUeNZWRZ3hb8Ar6KMZk4HW8RqFkHG6qPJ1wOmY4C8u7UJ2dV1Q6t9hhneDMda0uOvTlYTrT
6XVE6eq+GJqHO26xJJCJqOOhOzS9oERBrWtCZ2FptdU5H0jcimK8X8Z1Ka9gwidd+pxC2HxblHSz
cBTdtyjCXsWlLUq2ilha6YLhGNXUtMwTFKMtJIvJ05J//P77MbPz/4oFPHdIluLMVyv9w8AcR0ow
GuXWc3e64aRtcZR5PROq26sjLUOrV6b1sJOuUOM9Bdw6zY4qIQtI49Cu4NgeO1K+W4XTVJ45XYrw
a20jRZTQ32BLiHUo8Gr+G6+fmjJAIhUNVLYH8AI2UhQIAFhibnqMp7gKfoggPRkWQ8LfrljXcGyv
PQoLc54TQ3aoxq2FYYAJfDkMqHNYOUdfdPPxL0YScNqKsVFOPEhw1owaWFrMjNa3GDR+2YxvsEt7
FSxBwqL7zQp8KhEfVJbuVSjJnb/Vsb0HqqVCP0TgIEx7S+BCNPjnnTuu8mwL1WgMh5vMWndNJYyk
sXS16/FJycaVMHOwRV1xxGJY02CKykoSGZL7DwbbxMZgHpfL/2fXUhYPfryvamRfv/h7p0sQNXUI
UXbDw+prQnbzDx7ot8LH9AGJOVJ6AovOdy5/3tVOnsbwcrj6fU+brXWIMqjsjaJ933Plhvhjeyku
3eIj+3rU1xYgZnVBTTHY2IDEoDTYfISOoDm58/wmjCO1yj8zbCbo0IMGgAUdAWlbrA3mItpAYWSF
7ADnAPYD24OcnyqTtAdpIvHZo5ZrBe0wT9Tm8es11HaC+ulStCn2ndjNMTPfbzK61ttpy65Ll0Nq
f2j4Q9AxL76frxum2iO0Aq6TS/glR783UJIQFTYpZd0hDEccmfHCjWINAdmSq7ByQjz+vjwzWFf2
4r3NEn4ERdzBWWaY8eEwgmwAjdjGDqjHwLQtnU4dDbr7KoukBpGCbB+ez+t17F2875IMHsTvR9R9
VZNQLn9rm/SUZNENQdFu+fFnIwia1EeyeihpHHGPPMD8q8PVINrY/LdRLxhytBzIvNxmWZlsM9DH
MhpjTa/zM5gZ+9RhIdacBQJR+fIQnYuwPjiy605DNemywmoe+lTTvMoA2NnwqobNJAe/cO9KvF/S
iToLB/d2uwg5uD9HXOn1v19B42qrFHxYouQR0pNQlTtatpyCA04M8abgKpktIY4i0QZF2btoKfgH
nsd8B8B+zkGAV7BZDz51LfnsvGeK2uZ++P9nxdjT3sT2hYEjXf1HY8uSJQjK2a8UxGT/Kt7EpSqP
ErkgI4Hgw1+mjGIX/dKlSi8btsrKRr2LFwjnC2Kg+Ybqqljmuggfcv7oIMewz8sb1aBseJGjOkvh
HsNCmr1cx95v3ZLCn+F2DZMdNlxjn3u6J/tqaJcZTEOofnk4fFMTWJ6ymSF0C/v5OG+1+CfN9AQF
W2M/KeShU6aKLPH5IkTd0NHkkYwbOaRvq6uZp2nQy+3ZI47ppSR/a9TZ+rzP2ildzvlOQPlkxdQ+
BOBrouypr9jv5w2yFNBvYgWEHFORdPhfDDwg+WY/WHKIPRqzNeCrgISTphPmMGvD1bWqmK/zMtMj
4+GaYDxJ3bX5fiS+lEfnM/v38whoIEGp8/OkFKLAlQn9/HP3zqOfMVT7VD3n1Gtt6+UL3jfYf6eA
8wBbn98L70eJXxJMalXHPq4+VhT7cM4ApjQeoxdu/8lTg6TjQVlDxIt5Z81YkYftPaR1HMgLR+UU
3OydansiwYFU+8APEtpUxRbjmXmmTqEO1JDilGio1a1PWdX5zVjNFD6klMmOSNiPacV1O6+hHMo9
19x7FB3xAycqztvjtaDxFzHJJhq6AapD/131UGHVGmYEIVBv/0Ec2abLw9w2kE6OdB7eENS97R7V
FRjH326fmCTc5/kwsHalmOG18ZlW43zRhuWVEi73feZU9366dLeX6xc8Why+dYYyAlYoK/K1DI8I
0UvomRSmDKdSLBJDMfDdkgwimjbvg2py61s5y0cRrTZ3sk7qho8co8ARVd/hM+Qpomaf+gia/vjt
tB7GOn/6qxHI5vHPC60+3WD/Cgvg9ODa0FAOb5Il74gt2+rMMLBQhUZLFkJ8p6TLFQYvMVtbjLK2
sbLoGFxy0kvjT6JyTzzGyk7P/x+zgXQpJ4CLps+MrQQsYa5CERJnzbYsQhHoii/8UJx/TolX9HEM
h077qCeYD0JZlk8uFdXTTJROt96agC/kOES/Sqor6FFUZYLALYzUcYZNSJlIh9/RAHvhSWwopfbO
XV+xhvriAViYA3FyaaqqMzYUsXBEvTNoUxUCD8NjkjdjKScXrI5rAwznNfMcWNwxB/7J49T0xXZP
G6nMQkAHsmfEQNz9jXlgScaWf4WPwgMhZyXyiZ9Ypqrdbmtb7DElglHMx/GJfuwM8AtNs++I/rB6
9Pc3+EzvqGWorArlG+EXQAoiecHpV5JKZwTtyYZq+4MFA/D9Gc9466R82rILNKc0r9mO/GRTQv6n
5LB1GmyZX+UdgRDxu1qJrMKGosWft4mfQw7RnUGyV5gPNoXhq2iuDTqWgwkEwxWcfqf6uvOizFCI
Vy2dAMpsCY7F9C6XAwvHI/43t1INB1gsfVVg9L+Ih3RMgflFFeepl1t4Yi7VqmlLRtj4z8ndTC5W
BtNHYAjcqWNXPiLBaGQ6lMe4FY78qy9FP1NLTnwuiAr4c7F5Bpy5wrQYkhJQLXiHluUmWDYzbvLF
KqlNJid3OTVo+4n3sGVeY4+S2mImdRlko7+0IEqMSsN+tUwwrT7rBLMeqw8wEGSnZhvaxwdBOnGk
4cxoipbhNpjHebBrZov83ZkwpIiga/cFSu2JGEpXT6/8kjdFXJW+varo2xqGxgicvpqOujgmJF79
UAnFleB4ZVwvT71nzjtpxEhc8rmv8u0zErkhI59yQ40lQ1JkU3j8ohapK5k9pZm4atHmiuVEQbrk
zLwAbydeldr+guhXSl2GL8N6AjkRRQFLWA1jTN2kU5Folt6+W7XKZKuGM71QfG95vS4EaNsjpAXI
J0CmB2w1Z3YSdBCozHjsJbpI2svd8GWaloeBs7/RvanWjYgzF2nliD16bZZMb6imo+G2dJx4el5y
NQko5bEMZlKzKjYrp25kETZNdfbW114eYwpBsLRIcdQ57R3N450gvHcfJufjYmBRBK4Wkrrw8+LX
W5sit3WcoVdvv82VnakmPN5+EYM4kZ0QrqfM3u2MeZhzYW6momHTWD12gJSYE6qUOSsBZJYmNytb
6nHoqvbaTFUHW6KJVo2J4HbU11aL1ujruS/o4Cf9DmbTz543DpVkotiKNlG4J/YQ2g7fOtAlKYqn
VzO/TREAURSzjuZAwjsoLaM/sX+H2ZlzJZTnTVoFolXZhFczClPzTRpnbbix4LxafmnrycRlriC8
SieNoZ1BNdyZObXBd0lQDCnz2ycOdtGtpSfrimuMK0CJzxfA8nCbG1o9JTmOzcHDGyDEaCf/GPvk
ILjz35tOhKO+f3Y53kZeWZ7HkGNGljfgRUlSmETAB+uykEzkrGrPIpnOsUaZo82BwRc1Arue1l4O
asc+gpneUY6rCk8Ku/DGh9CqkBk0DxPVldH0LgSpu5tTONcaB1O5k/QGI49/ydDXsFaanrr8dQ25
vb5hcL8DpRzIN4yut+R54bK8BxKmOK6d557Rf5FvQMnNP57qw6hymaTPf6i2MmegK1vDqc9nu3h0
n2peo0GrxPSo14g6xoeTu+nlzqws/QCcauTHyve5usl4HrFsz6N9IwKnCA8JPsBXtBhmyPqNrzVN
WEtqvhDvNidoJ0DWv71ncgTfk/hsIB5eN+IEcdfRjvnH+pPAKrCf5ePHH/p/XXkKfO5md59wjGPr
fbZ4k8SqKLhcmTht2z4ItwjtxKSZwLd1RYAIu+7+/ljS7EdfSOf5ok1CIOwZa6FDl1paFoBChIUU
la47QYvyonWS9Lg/Opvpi0rHRnxxrKjgQ0Bwsk2/fYCv++5AjpvhLz0WP+WIW9f9sDUEFTs8Ldco
YaI3oFFuUCZOLd3LRjUuWp1yveHxbOVFiXaBzOHhiyayGwSOKHjD4/u/cYbLz1jcyFS2QgqDXXJi
X6rOznEnnyyvskTwpHkrKUC4Ewb5KDbwkoMnvZrXCjUrAef0TKcuQ0BC5XnD9Ohl55dkR5Rr0iw7
skseaFYlzENQr5YeF2uETt8NCNdmdfA4kY4Bpg9GmsfvHRLyKe4yykXHIoFqe1o5FU03MFUvSDHp
AhYuBfZbHuMw7fHmEQGBINrwfs4ZdANMYs4e3N8TCCcsvY1V0j6cNIXJPt1xnr9joEfTSzYmRzEi
23i6BvFV2zu5PwLYkW60MyMLp1i5PcxZu+kwLuw5HoxGyN40/pTGnKeiR2vd5PZKDTJ1J/OnXxBk
tgVnNGf/y0nb9Nm8DuAOyRFYMb1/YIoXU4gAXumHqlNLzEmRzj8Kb96P7wCJvHvL7J6m29xHbyCp
hvE5/jeur8SP2VnxDSvgdCjdjL9JBnt0dQgLE1GgzTwo/nSiFRYx+lZiknmIDQHAJ9m6YFnOucV3
N2I1yZf8HTCLpeq9n7HxtWP4jLEFgIZ8Z5lzLDjVdr8Krq5v958T+7Yyu/6pBpqcvGN5jN4eRZKb
xa9en7oVbzhb0YNBWA2ExkPY/czVrqzfeG1uKNhEU/4oDgeraHZQGveifnmWVGZ33cz06yaBWItt
bvJL0Y3e7JvOVX2h/cs77B5hug8gc3Gg7fu/ABo16NPVm45hn7uyGZFCGzzmJrVUE3L2oycRr6Bj
SaQxYUP0SPJxFBxODuN0V63AxdXGC8INyxbWekkRA0Wg7o+y1M+JpyrC4LszUWxdfyILkjdKRR46
vgeL3pdyv9RXRtLv2RRpY4yVmBgCHoC6pA5MG2a7oLIHusrKwFaEqt9vb1HPbdn4YVY1OPyol5pJ
LS/z3u8WBiE/Uqf8U7ZE0hOuMEeYS6pxi7RyIY7WJ0b7z1GYrH6inazKmOBYBynq+IUBouVP5Wfw
UMbTmjfx9H72jiq9RxXIxh3q7fAqnjUiHeuXJUI9xf5d+PrioCJaBCe1xTc7jD4i+t1r+m6GsXVP
xOMO1C5/RT17XCIqWs38WE63sxKvi5AiCCGvrZe9fqH7MLAnHmjQL3jGSovy3L18zAFla3IjzVJM
QCMZv6jRbVbb9KpjqDQfKiu0g2j/McQbU3tgNwEFb7sI0FzMYO1UhPFAJJc5+y3NQFxHXfCkSoeu
P6dXYxbiZtYmPgfUpxZSrwqPGovy+ixuBxX67z7sLedwPa0h5aUL5wK7lOXuXwWxEXzYpDhRDS7u
BMDkHuEb9WRSvJVNKMNbztSafjqBjcXgJFouqCel4KD2bSEjOzWXZOuQyOw65cNn85FsrnPEgbFC
FGybdEl7wZzDacNpUtDMN11OB6xTz6GuerGtOjbRszS4w+igZTIFRoz10vluL++q2iWEUDy4MC78
SnGDzSYyW+eAM2GdS+L07izHs8VPz3yDdlbzv2OZxQ5dZPgCyy6uyelruHGT8nKSNUPqKkxlaOVS
3epiNyNeOD5SKuBSqF2ha2cwW8C4np99M1GvCKtKehKvx1W5hblSm5QgmIMgc8j4+8jVq1fMdIP6
DIrsJ7vQ/w0iWFNqfUPPlDfaRIVGyZF35bHcww4f1XvNvw6BCg4IUo7RyMfWJ8jzReGOWF5O3vcQ
wVaUGiQBmsTtZHWypmRTNqaAkW9OO5rw0oGJeCZ6Og1mAnIWV6SYGINHtAEypiHMB720qmhJ/mOc
wziyDZOEu7VTgGtfecpIz7JCpXskGl9H4gqt7EngZZ3fsRMcIU0uABsZRcf60M33gHgHatRZu51B
ZHEKRZrxjbc9DbNQcnHgY8slMzofi/WutDe+/pGeL9OCgh6qw+CnR9MRAqXSQCrwfTrFhTbg44Ov
qPpNSO1DkXU6WObMLKNkovrCa+W94hBUqIKnAz17/Uam15eZWjYT2XHvsuBNLEG5fKIVHxm5Rf/V
yGEmhcrzLsftWX4qfkIRviHEw9iH9FPkjvYFxaQqqjIKlTyFhFLz4tge8UZ1wWsRyPaNzd4YrQn8
xxKFrJZvDaMndjOxMkkybX58odmDTN0hMLwYncvWHKHavSyFsw2tkxh7Rw7x0CKIjsb4q7/7siO3
8BdxXWmcAfgz02ECs1g9pO1whoD6pYyn6goDm93sFBFlJJyZf91OGp0JKtHKD5sJ0s3iPJVmhHQd
/50Fzsm66kZCl/fEjRp39pKqStzQCY2OTfoxhAkst+EGzR4vKt6aBso8ZjzndC632AAn4uMEFny7
FkJVQ53QeHXzI9pE4zEzpsyOGVZ+flbfmgftu/yjSlKaSJ4y4kZr/1r/pVTp1oG2X3bPRy7cuFZf
lNcb263qXBT35tZwPbFGWBOiL8xpR10eGvtvzGFDInApv2L9mEPwHl8L0UsjXgiFTieS0skfsaxE
0sF7OngZkgFpZ8vVWWWfofF5BKYLSN+hshvuXI2MbLVFgTqWaeFDfybn4Wz7xmJxFtfn4iUGuEOA
12Bj+ovhkb8brdA1uPKntY7lRh+J00O+T/6XDpvxOFj75pChhwacFpTz+s2THejn4wKR5VRAMuML
j7hMMMa8fIymLzVOBagWo5f/6wDbv7ykipaICY+51DzSXaR0fHfG0u17Kr6KirjsdDeBhxBsFW37
AL53BTGqdbPWO+WvETYxLVpN1a0SiGRg5eolwfwL8OxPE03alHE3W1Nhi2BLIKxkAOFd8Kcp/yf7
0glSwHeBmJejB+DBr0FzhwJOb4ezVRxjnvUTx1xzzgGSucfbLu9wwD1BNe3q3cyDj450J3Th0xSF
kfdFpKzo8WVNusFtA1vfx7v9KbSl/WcmJ2eYwyKi6X4b3bnNohw9BR1NL0v/puHWwLcEWayujlru
iR6pF9mMqyk4IFL6wP8pjDHubE8ZU9bjU3es4WgdQGRZZwvnJXZfOmKWDeyau0PwxJq2f4OQaZgm
O9CfrN2g2kcLe+5vJ7ByMMtL9VuBrSSLkF1ZttuUH7SKBxohQnOZe/rpsDSjgv5WtEX3IVfOsDTq
SPR8a9jeFUiN7AArc93yPoqwE+uMdIDMI9bups/YF5G2WqqQSG4AryYCo4TJD4xzscBYmYf70L0a
MS/oUYslCMPpnhDRGdvOyv75F6wmdwg80imjbwjbH852XiCYgdi2aZnOG1PcsKKTOlMtsv4ylgp+
N59w9K4HfcKHfN2Tx8eiSONrck4x/2QjRt+B+4KFC/eC8s2KQEK/t/jiYnaUCaKlYvvBL5Mu1Pa7
jUtdOrM8ezJPtb78bFqfqKd4Kks7Ct/0L1iiNa85Uqn0aff/HizZhWJlgIC+OZY403vjik43V45S
6NFBdQNhyjqU+2iAu1inR1Lu9ezn71nK02qBz60SmKxP7jTAkPGdXVccgvYlCnueX6zkq14dOe0d
xFiNtJnJEpZM2stgCRqgCbtaBcfejq+4MKj0uUWVzzdxMXMkudjoBOLdWaxz77OkW+mkIKY0BmK5
c53x5JCJ+IIEeb4SvclULZ0sHQj4ccPSDN57DuDwWYKknXWby2iPMH0aEgMaUcnT9MX7J5Tq9zIx
QaTncaXwSKvl6A48qL6pvsDWhmWQDgd58jDyRY9fQ5c7ijFnVJlIRhpvzk+QoesmTxsjiGfE2i+y
y0YrXOLTUZipLi5myR0ILzaBx6yrhzmTcgCIEaX8m/KLHXAbVfXMn3qbH3CN1ajb03Z5ZJhCkYZr
G8QjwElpFEb3hMyumaN7JzmB8UmcExXIZzWpBQJY3XzIcAfceD6pawyGMY5BB2vq1Vm1FlPn7NKy
qmra00f5FOWxJIGrJHbYDc8oBPULaz++8lShNpZSdNNtHGtRiUTTH4NONO69LEeNQVvaepScszMu
FOaZWu+FWdNwCXaz8bWSBBW/H2Wgy2Fbnt26Cbd3ZnEARjR94wox0pIvo5rZ0RRbJVLMZC4FDv2c
yYdA922rhQChIVSkVs+FbZNucoNe5fS3uEYza8ZrbIK1y2VYgV/OrOm+9VjRL050PNlNfXSlm1VU
qk2QzobEl8+SnZsYHmEm9uLyY/lUqUl5BTzICFxujv2iDHNxbcyJ4pDNOrEu3GJ76Iw1y9iaOuLq
q62mBw0GpnGdL3WTvD0t397SR5lzTszYBI2bTZEDYK6F8RJfB+OKMqNk8A9i+ycxPPMKxCnSqA00
IWkuTyhf4UptO80zk9x25SHUSLb7FYmKO7t3zMi6I8q3sjokH+gBJo450n8DKw4XTxUBNZC0StEM
UtvmP4aY57D5tZmrwHKnURjI1SlRSh4xHEnJ9kuycBtBnnxwlcZTw0p7QM+XzQG79VFFYe6PNQ//
M4c/sotC/gdVm79Jd62Ex34Ye3rSWPuOWHQ4oxOUQ6t6sXUL9StTr4hAhLiT9aRGeR/fQV0UWSgD
69fo9C3txYDrWYDBwaBvyi1E8u5AnWd/eWKL1uigBLlIXilRD2C/dVlUbBNmVufk0qKTW3xJj1wz
OWEItl2ErJKR6pI2zA73nWXRSezW8Rz0w72NzxU+mlTVzqqKhRq88cajoy9bG4K8CUsSbjee3QLM
iI1FY4SYraTafr4QvGr6+M9wpqtYIlQcXHfXcFTcB77b37ZCnju6oQGagSp8oHhra8vudA2XLrbj
yaRNCQkiiZMUiSaokbGj2zMULMk+s9R5LlzeXJ74DuYsSADkqak6rodfYUPejr+iD7luZJe4KNRA
2pmgBz5+D7tpvs1nFLgabHQ3lCWZYqFFFtl2diow53XYzFN69yPjb11ljhTi7emc2P3jdVDatQ4Z
hRJsR9NHj1QslFAcBdonW/DeZp9rhzGNKt7i7yvo71ydMiT7IKH6fexTG5x7OcpwCGTc7QP5nv8E
NKwhsCt1HX6ROl1kGV3qUBbpPop7GY4OQKvSUt9NU5k75vU1Lw6xHnydLOLNdkYMS8wnrWIiuXGz
XesUujybz6rv8BN5yElhu/VLXJY5fcGTsPd3djoV03Bn9M+ZtULBwcvZUZLrkEPg5CkOpd1xudOn
NVULWt6QycyRyWVf7UEwim8PPvuadFKl5KZwRw3zo+YA0lF67iw8K35oIulYkbYQNr1MEW26CpyY
QN7MFhY247gOP/x0s/AKWXyA9ViZY4HmpqsG+OsaPWreeJHuYHMaE4Y/7XZVhNkGbvhdBTVR/67S
+EvRo2ugFkEl2jXCsUg4Ksvaw1Yst5KnZeer97LvnPA6if/VlIBJXNUTq1BdDAF8WnE1NwaVBD67
/3WLY2mPZFpuUfd6DCyyeu6mT1SvznoCX4/9FRS1HoEsq4ALY0E2xWeYddN4tamjjBJAoep71Dhd
OyeQT2whOx7jBpdPoWR38bNvZmN6NBY9uEQQcQ43jhNsm1ra9YQXZiUgwy0RdHA2WqMp0KAkIPBF
xX0YIhwrdok0VHm5HWZ+KtjeIvaSaF9g5Y89lTlu2ktY4iaY8qnCDTFWifZ97wU+yXp+V/hjRyIF
rHV0EnGmCzpxqYCljgzjjA51WVsXOUxMuMMkSmO5iFY3/qB00JkrT4oOeflkPxI5Fza8icr60IwE
QUmFPFXr7we3nUWp9WCKxD+GcWmSHMLTiucXJBJlkKu2kOlxh3ZiaGb0J5kBvQI8KJkYZQXmi+pY
JTqTZABDQWMREP9n6vcD4qw4fWGAwEYb/delbU3Xyf6O4vu4EvMYWaFsYYER0j4/lj86+49nVmXY
t+Lkihua5QeY990UicKcS0cPA8XzTHir3B9YhoVc4+/AxtB8PGzr32r5b5kuimiuSZ3SjR4+Qm00
l99yhtpP6ga2aKcEqG9HxcL0t55hkDcJ7zOkBtgjdYX0gPV0hQBkzPR5bOjpZBhMS6xh9eYBabm5
dBTNatMGNcF7utrXdicPMAB/Fn4cY4qG1iaNoBbCFcG1LQj7vdz6EWUfw1IJttlI8tBT+iIz0URj
lqGLkU9QATTEWMwYBX4oV+Ryhq7GP6SsjyeER206mBKJNJNm5h94cSqThGSPHr/6RfiATmD46KGS
NkALr5JQy01dxebBqWpvlZn7Da2a/mnA5/0dIa4N96hrdjbLou19sg621VEKWQLOOic5QhsK9TY+
dYM+3W73sJCWkutcSoauPke7c9YUcAI9vTHjeNfEupikCHmmpqMCj6ZYXxVDaTYtc49e5/7fJUDu
kJE5W40pgVMIqWwcQI1kbPNhpb7TJ91HFFFaQgEMDSKnTcJod+Zd4+8pUmQrPRolLrzNiSCqsBzd
xMVPdJ846NA05bObzEnxUE5juDedQXGEsv6B4xsPdqX6W+wnrJ7LnjxLG9N7SZYNpWy9Kz+hEyhW
vXnTfnLRL8+S6LRvwU20gRZJcWkGuNCP2s4l2Wny5zon2QzMffMTfkR2A1gpAs+6CdtFrfugs8Fo
gA3kZFo2WpsFeYBTLnyQO9P0dsVFtSaOBHdY4r9cNbGfcVpL0kkvDSq7BJS1qeb96MfDDlzCWVou
BcS4uhnDlw4JRw/3Elc0oCxCoQ7Tn0JSYZZKBCHfaw/cV9FlydRu4++audaPSb/L8va2mNnlfmHY
RYu8yso6+tJFwl+5nFJMcy9DdZAcV7oMQmHpHCYzHzJrGsSb4dYF/rzX9emDLNQq7tG/dynz+Ha3
p4VqOFJxVxMFSciaTQFlHf+HzoCRQc8Jl1W+n4mX37AWU0MMlfUTw4VYB1E0PWlTBkLGoAoHpYaO
rcxd/6qUg+4jmji1dn7DrnLzKmKFEfwDIKr1NzQ9dLUwTu719hZFHXsUfaWsx1GBGxRhjzQ758wh
IoGGB4qzF/YuNNXmBQPDyjj4lgOwqpX5NDWf04p71BGupLU+ohjZ00Gd6oQSBKvqoiPJquRaaJ1g
beobqeFz/9QjvIe1IDt5XuDOTlCEWdyl8VFIYriMiRK97aKms3/WooJdZLOrCDNFXXtibbAxTlFj
A+aJtvJHoos34/DmLXT6uNvcgggSzbMN7SnhU3hld2eRC4YRIe52ahI/LfYv8UT94h2/IlXqWKXm
E1BGvA6UN7/QYMflr2IlaWh/gPx8BFz7fXnIgyj91ZeZEvORy7ZCkglfqTOFfvB02N0J5IOjszoP
NzWd+LsTrTPEFm2PGGxlg4M7MRoTjeI8Qi0s0AvCkUAV+/HGl00kf3d02VtHKyQGwzHDFmKp51VZ
D0/QgbZFU2af+Hl+9asMUQyLXiMgH9NVlKAKnufnEmuYOQOwNbmMldk04MlLEB0AwT1lwR7zKGvx
n1B3l1s7akfa9594uYI5hl2DXJUDEaRlxqb5M3t+QOwHj+/VSRaN7o2z2Z9rxPvrtQvpea6hLGty
I8HjcMUJYy7ztln5kiifQqOwBo3TZFLR+z66zIJPqdLpL3eT2rHT82zBU0hxOoW754Gb+G9jiLrf
dBh5f0liQzm9yYVxHseXlmnsICFNhlR4HhLLPPN7vL7JdgZsguhWMKrVZznr/lTnVKpNf5kkZbvV
24F0W9US4b5rXnNzKksZwrhhXLrPeZGb8/V1Zf6xJPzYtwrcoTxdqn2OJyGs3hRI/SKe8CUiHeVF
VcC+IrBuSITs9+/hKhmT1vmeqL2cU8X9os01D7c4DOkiMa1a0AvSA5UhbU1rEkdg8A/BDXImAx89
RalhXEZT+i2U9+AunnJpW00BeMImUOS0XnBjwqQDglwD3unM1s1Q9kqH8Ipxq28LCyPmnr2J3p4X
joF5FNSzdI+myOcNpSU3v4H+NpBsP5Yg3Tp7VkdzNq0V/e8GyJTvmcNrKqI1DbKTJK8a/82ISQw/
Rr12cPcA84WKzurpByX4/QmSHIYI7Cg+2B8lZnHLjjuIjjq2GBU3iMaPrk3rVOhnaFinrah7ksvq
8CMP+NrAZvEpvat63ts1BllcmvpxzrgBQV4wvhz02Oj2BL/16CYLkEdfVbTsj/amvrUxtMeuxAo7
Pxp66qTFxfgyL6td4tW1f5uqVj2+acHA4MSX2vTGcwFLJy5Ncxw4Osni4DDq2qdhp77QU2v/JV0p
+fEeNrRtmeajrsyIWAiQrynPGiJbddgqA+PwNfokS46HOx49KNWDK0GmT0EQJpFQ5RVS58nuPyYx
tbWKRg9IfXq30bYpd7HEkOY0xq5PEPD6Ypn8B857RhHuOr30k8TzFgMMOqUiGhi9RBotoK4fQFGX
K5btGX6tx+baJwSeR8yPpP3RMm6b80U8rLM6yxFGSpoYcOW6IL/yn9XMKEaIj6G/TxDUVIj3MPSn
wfYIHFgr52ba7cJvFYkBta+m+MAiNghfBwEuhu4NImB9yMxyrdsK6RnNWP/cvx7VItM5Dy4zQZuV
9AIl88Uv+HSickRQ9WGry7+cOlXl0gnqKe3l1enl4v1Kh7pgFc30ZFOgkXgCisxOQ2/BmI0u7YQR
KybSCH7/o9VMJeOB6+1vT1wjdGbQB+6U9pY9lt1waqwXwCDPayabreNAYpO1XgACWmPWY9loVjBI
EtTSO5BIlNAWu9ZdhkJq82mfWFBgBYeBXv8diVMkbrjdd5b5r/RH9e8KqqUtlLR6n7QDhSTEaa+h
bF+JMcvUBlQf2z7AItToxD5bVRNimhTl+RjgIZi3obj5zUhnITXEyt/yWA5yy9Z8NNNJv91jjdzb
wx1Byp4NqUF/E00w871Gqmkj/dRCgrwuvd+gvCfaLCzYEXb+QvhXE1oINu93E0TFZBVG+i1HF4fd
8BZCx6ST2e2B/Nq9lUBAKMqXSKfetj0hMQ4k9vvBn98zOcVoWivQC9q6nWp4Mt1eAYHfzRe0G16x
AGnwOgQER7tzOfclmktpfIWg9IORjneFUPKUqZ8hJ8z28QC2TOz9jV2Aj4zcCjN1otpJUlZlvSyq
tORBdgh8o3OS0yynINkZ2jix00VOtt3K0L1MNy7MVIIOAE4/ySlT64QTiMcc3cb/SpZgX39XZKHw
hUJWu7gCBWQsE3NHPhchRfsYFSPjyHR0Dx3SGYBdEJz+XZsev2tm+KumX2IISUj9+6/RFpcW0m18
kmFfR16eNfbWRYjCfQbiSQ43zVxyBZU0ZTOREs3e1/q5A14FE4uU9+41vN23i5grondgUTN/5Dza
XmAYGgD6bJZASzHWz0O99Ucn9X/2ABl+vQmRXmSRzWpmP8X3NsrOLt3QVDPZ6Iq1do4JDs2zg3ML
TESTDghm4YP+dvsufszqoiHlhA+VqMP0E+YY2m0/haM/MVJ3Cu7eBapm0qDmsH2yU58fsO/C0gln
zL/Zj1ClZMR37ctis+oNVMltXnDlMiLl1cprEl1lrhe8Y0nrI10dLCNMKnDrdY5pFygsO4ychXtu
81E5IHUX1me4WD11nmCJDMi0wyC3EK/TKgMIPjPgEKxS3BUWondLtZXgWQOQrPTC78909o4kjrcM
QCujBk/kYQNvsScztKMlfXVYzybcn1qwQfliCOI1mqLGTP9SV/rItGLZrAW8V9bDxFZMgP3V4ITc
tVvj1Fm8JZv0rpEAXuj50EZ9IoFlT+QeMz3GUAI3whj3V6xl/QXLlaK4f5mo28RhaOmkBD5NUIwL
/unj+DrWhaZJUHI+sv1Af6OZaYQC3pgREauQlSjriFMLmDIBuA2E7CZ2cx5G/g0x7xnC6kOB2Ord
gR0XyfvkBUA6VheF9o+0Kw/DZS4iJMmObBICAIR72UB5riL3qLYvFfWwBP99jWJLsXlDX6oYBwlg
GsGzALCfJoz/iXFjGkTHIaVidAjyho5ryGckkU8jmGCknHOtHUjZKYjkEa4TMOUaIwbRLohVK/j3
pcNl8KS0Ff4ofVZFh3SbZnmzYxI8yaZYi1vdgZbqZ6vZUmRDSlR9cJNGR0OOSlfrVsGouFij7fRj
G4EFfZFCCSMORWvm8bKrA1eB4ZnNuTKTKrHCowu5YAIhwhdl9joZW0LAjEigZr6khMY7/07xNyqY
OvrrB+YIIMsxsVHYNll41yyoJcLToEYc5OJlro4mpCcqw30kp1sL645m9QY7UGR7P+W1LfMIkovs
X8dqdXo6HIWJd/ph6SfzpoecuT3/inOCyAK3JRrvh8OSPfpQ8jqwxmXJ4eF2z29JsfRaebCAoSDC
bMQzMIzfIcZuY2npqad199Av9uQVL9nd8f8tKp+vMRtlLf6j4qTCVfLeXPo1NRYEpFbxlEgbD4yO
DtBh+toAJHVsbzHFQUZ3ZW1NVAF7Y6LeEIw/24+op1ZG0sN4BT+gOERXwU4XYaheWs1DxW9znilc
ZDA21tBoyUeosztBNxRs1cfIkrvlEsBmWYKMuUS4DzMfa5g5/CXOHXCs0M2BdgMS/JzBpGe42FDz
9tTVSKZcsujrQh3UH2QYdVGSiWpqkADdYVSMPLEX3VpfjDQLzqW2bgHaflXjMtidu91WYCE3SFVl
2siegYThfK/HJ45jfEOMAdS2bAGyuBbUzIhB4vfCmo0NdscgLSbi06+EFGd+x1YgkshviMwCM7eE
y6coRmjPpFEJC6+GiaRDY24LJpnCkcw5sDAkIn7IAK4wDTJDdSHq5n/j4ii4P4/9/nuSFDuQqpY3
osSPHHPR7UIdvbo9d33XrVnNgA/T0xwrNnYv4mGCuodGGfiwd12TvsSeWKdQovrx3IJVPngkpfAI
PjbeDxkv8Bt8207ltCnFm2an/nOPadbym3fypl9swoXNQk2zLkFYjLKnH/B1VC3SSqxdMIIUZUlJ
lRp1TQMAr/jESz0IPN35c0ddGxt2z2VEgCxYAWAT8T9bwrokBUq9qTlHNxFp9BDVvuM9j74+OS73
aYPbV1gjRFAVJW5HXdi9hslqdDL6X1OtMBMqTWvFbxcLG3Pi1mGSzFQHxpuXyZmyR2Qq8P/OwnM+
j92QAgP3x9D4/Wkjo96LMplLIZTVLixa24Q4q1jJIV1KC9R+82fAVq3GelH50pjzkrnqPGvbbzkG
xkwm7p2TIkCyjvfa6T0ped2kl6rqtICiZyVPRoS8q8+9TV+20IIgbqs9cyVdgEkPKwVL0nLjsOdQ
4iSstPNxcS+KxK7lWWBLJuEziBQDQ/K6hvwLsgAhBhS96vnBk9EDyCBJ5ubh2W0gISG+KUOv00Nh
tE7IgxnHeLr7s3lNQ8tnO5v1kb0FWa2pkAIIdh78tSsY64Q0en7Ya8KqmJIrf8Dfk8r7dI84uRF5
NUGLAZxcV1rIFZIun+vxeiCpkMkX2ZFWzFAJmUSVjiXvCI/Echz/2du9IiVnaMJH68IH8bcq0EtE
31eWcl95Eqg5mK9pRUl1tm8/n0NFWFPv0TsWfA7wOc0K1fO1fSg3QvEfajAfQu64Q2ynmGagYXoR
qxgPfFUVeWms1MMMToEvtHtFuCdTYTeQzwKb50y3I4uIcvNMZMkcE5IBkitji0rbqJ0C4frg6+Hv
JslJszpGEZVYDMHJJzLpw9JUWErTy4WIWDYAaX0LbE/rQFZlZ9yDFr4r6FVoKnW4vR2Z0NMsYZZl
w2YqaFLyZC7kBSGtKYaL35bAeMyhpuZrqu10Iifim8UUvfJGepYUrO8u35FGueJ/ehirABBsjNrw
tveEw/nKgvaA+BZ/XgmU8Ql89U7Nbm+3WDEFDQns/vi+i61F/HZfHk5eS5e6Woe1DBkRHVKLLl4F
+9LNiEVlsi0ZX7TmEOTrncxDsru1jFUUdxdHsaXTTmSYyRGqKRFFFPjrxqynvZJbmRYRdn4cU/vv
aWbjEMOSZRd8nIQJMdTUM9hRcGH5xpOSVuyzJNOeH2vNGMG9ZWrguwfM7iOu9vzYd6AGZbePfBJU
BhfacJtZYcFldM2SVh35p2V+q4Sg9REPRq0fGwTs4ICKOBGHNkmc4wCosi2FM/03L7NCnxcMhI+Y
mNYkOwxoQZZ4pcE5U888FnCdbcTzzKCBsHHPT+r9XuIkUJ1heJcNzD12MJ70UDeH02A2rVqJcX4S
Q9XoUFqL+WMp657STF5mdC65xUCaGGHgOuzxGIN9l+qM/31IWZBoVgcoSlpSYejCPoeynABk8R44
RiwOIG6dg/g/ZzrvSfa4QrUbkQGjdYzc5BT8PQmqtccDosSad+tlmYc6h+mPDNQmKbmZN2P9Boqe
EsJtFZCMy+q/gePlnmVwGZp7qpniGV3FN+hpEGvnVaJ5G+z73aFeVU9HX83lKVXmVwBfIu0WIKoR
miQvu+8GhpnZMI4TyXEIE6XdlzABqeJcxnr0Kxs0jY8OtPsX14rUujEOTIvwiUeKInCBHUTQ1EBv
vzqXETosuQWiWZs+vFiIESihxJmKm1mXShpVUqLQoio3fj+Jhd8QPwILAwCcd6fkRSM23E95ezcN
uNRUdiZua8lxne5lMqW0d87L7fi4RO051ivf2FyhZhhs5njcWSB/Nzap0y1eYFmMNFB1Il/TMpgd
cnhrMkpmVsFH0w5NNN//WdjUiTI/vOI5oe0uulTSV3oSvhL3pmBBqbfgKI5IJRFF2Bd9fcimSZGj
+90faIe/WmL42JVPKAXHQZ0hZNYhg4Zt/es9xHQpkPmHm9lSMYqQ6l+Jnb6mEXtDMw2lgmXWK2ZB
ij9+0xm/Pg4XV1bxcgThDPWj2TkEGfK7GoBTIaUQ+Rzn0l/8AIjzYCWFlROO0rugFcrFv/+QnvIN
q1kSDgAAWhQ/EynqYMDEvVRlO2EcOr85CaXmlwmLcXY/3YUdIEKMLl/b7/ApGeZITJqMLh9dk+yI
BfUjkIrpu9gGYiXRk5k8leBGTdPiPs+HTFUgsw6B2NFXbbIf5VR+NlT6dOyAk5+xMctbJNFubx8s
ylNC4mSxhmH3fTafp5v9sxE+D1jU9xc+Eoouvfh4/M4QbHYwAV6Na30wggUMtKWv5bsKDEvtnhgf
tQ8FJqRi/Aw418V4rJ1jO9ulL1KStk6JzhGKkhse+aAqqEKHHZJgcNMJpl9xtsjxK0qr9kibVX/d
yjq6mp6ihEQVpHVMWSmDXzPVgLYmlq5AkMdxBkDtGPJLcugxYB1zoKphXEPipeCc29u/Qg4bYz6z
DhSlnNkI24is/uuzaXF7WAwvNup1nosPPn/CeJ1/t/8c4Pj911hfbrtmHdB2UCCG/xiHW+QRfleE
3tUGhMzViy1luuxGyrPj2KSY4iRWujSc3aQK0DxwrX+lzzcEf3tWLLcrMS/Y0B0aP/wex5QI8bD9
ZO+YFKUPd0gVB6Z4tneawmljjMM4MWYMbGRiuHWoelGkrNbmNXfhSJT8BVxgiCXGtjxzGLcYNKgw
IOS5kJG2j9baOqjsKJ4P/LP4fEn+q0dmLQR7bzrTvKCH78ducK25dUrxud6gH8q02M5U+lJQ+Uh/
gVv4NehohEKRi1v+85SNFMVxXK82ShelE3J3lKEBAj6aox4il9/uTbaKfcZ0k7Aaothk5ZeuiSvA
JPueaEwuiH1vEdF/cvZcT1yy5ZYxm2G21qumw4BUp3apB8xXGgOU3nppONGxdAgF3vltw9SpQmLx
lr2cuFGdTqPn+eA7KfV77i4DagX6RIQt8Zlz96yKaUbFLAluAbuHX71cZv6yeL5Q5waIA/pZwKEG
dhUoOzVkrGqkAVHqXMKSVMzHYpntlDxNpQaDc2cgRkBnU6l7XmsCnJHqsmJ73abfm/3Lk9j5ZLl+
N27gn20Xdy7iaZBI7WbpaC1woJqzqJaCLBcvqhyJBLSNX2kvuvi7Z1VOlpHf4e5jhN7/95pS8PhY
rsrwvjL2u19QHz+4Zmsxc9SJWoIFc7AqW2yxGQr04+G5SaqpvQx8+l6HJSa5lUBGmlkyecNddCiU
mole6e6AZrw+smrtxeXixE2+PBsmyZeq4Y4/GLKIwRBtGhSVPj4/PtEYGHDMOlm6xOusOgPuY2Eq
PsHXAeJs3O03yr81dIf9mcoLw1raiBnbAy/WK8YbDT0b8JYyHBy27X6EmXjeanDocS5u97FmdTIz
rP6BNpPypUbnflwco6suXByO4tP9oscpk+YTFw9kuKSF/p54315JaavfIfyhCSvmMDvLF1ES6+Vh
FSjfrDLIb4Jdd5JXg2Q8WU6WjcwNycl9f4SFCJhCnfIae/1aH30+wlf7WU1ay5hMk5rbsYu5Q+sl
l/WdZiG5p88kDfsp1lbGa1cItPQdsyUmihmKGvIxmkkCEgKVCav7FlWPHXoFYzzOSNlFDNzv7ghI
L+OE0CuYDllNMs3tDA+QXwFf0sI4mVtyNMBWskK6UHSnnPHgqTwerQ4q3zDxW907DE1SE5OktNWa
VM0t/n5VysZmOkx8NktPPlhq1XA230xb+jfg9mgHQRQ86RyeyJFh/6W/vJcxWNeXwKPML9kYXQhL
oAmJdbGd3lLVXYEGm+gXBeDhrjLVhEbi6P8D7dScs7NYQUi7SrBj2yb7Ea8sziOL//5nmfBdMcvv
B0koLYh+lWciyZb7Hs2bg5C4ciI1w19nGYLU8MeLS+kEDmuk2D18RNiSxdC7zHcLE7FhsDEcyfqX
K4o7QzSPrMgg2habUcnV3QVk4kN84VR/+p23NjBjOIaovI8eo31SG6UXPfDZBwmPoGfsgmuPAFV1
EFVU1Vr0oHmxXJzHtnZs4ZZMfxSb/w+nb+kgIGDWYlsQRrI7qpH3EpNZpDwcZpyI0LD/5RwqsCBd
rWk9k789OIWUit1hz4UJFp/h8FuzAEZoP0f5BkNywr8TxfRPY2+ToHKa2FzmsvURROl6ZE8/9P45
i+QT0t5OL620HeEz5ufM7cWRKBDiKYxfvB93zX+8ZMPsYSb/bDRqKHLRX7azN86LLEwS+Hcb/EoM
fG7PjjpqZijyIVE/1r8VT9z0nw9xjI4JtKKoGkqLyRxgEqhYUFFC3tGKBUNQGTYUuTwR6BrZXWlL
aMoAjETLKATSAatfKYaJ/5FhMImUQkfYbyoAcBJ8pzsA1/RKH56hh0cnhPYBX8B/m+LuO/nP40Kl
qx8cXaH0iLJoGwZZoBaUuGFwQ77m/cFjKo9FBJvcE/eQcMFI4botcRhh1QLwiIllil24gwdpRnX2
zFYE1z5jTBzbm8p7HpR9Fv5D9+aR3HVEfMYln1G3o3Qh64P8Q59ozV74gPtyY0II0LvAsoDDnZ8D
/Esp1m2gHy6vxYDVejDD2TNLrN9bNTUi8KXSDh9mvXSLJp9YFfUoHNFiTREnqun9FKSV96simz8K
yyoST9mvyhV9G38kkVrE3W/xEcXZ1WV8pZv3r1m5ARkXF5DJ1FM2S8DrEhRZ8EmW71nMT+7gA6Jw
3YRiwbKPrp3TFbV2sz3oUxbvUlr32Jhx9bKgZhkaqpUAsNqJT7uUGK6vdNGiBLrly99VMGTJJwmT
whvocvjnUyAe9rGibWgrbID8B6qS5v5+S7XNJhoHiOQ3w/Y5SgQMCrTjcgs7yF7HxdAG/EJo4nRd
rXmVXSmXSfeYEFKUZtVJjLdH/zqZq1wvYR6KVkDGtJ7jFkVPRQUAh1LAMeBQ+/nYab/yOF52Q8U5
1pNcASgKkHNULNm73tNgXu2k5OrmQXxWEVWFh9/10gAv6zRdBv73C9lUtY8NsKNUjWQT3wj5agMy
/UzvBB8wJbJwoSm0mYdm0Qb7ymgQYa/VLeFVL0gaTCQDaaTMvHL/6e39H7kIgw7rqGhMuzR0dLB/
8QqDhKGLdQvQlS9NmJKlTUQHQdDK4MZgwEZBJP2wfqLwlDV29jQon/pQbspSeM17r8/IDz/jCNvI
LW47e7Q4+rS/c9Ik7LVd4B8aUxfg0sCqxvHED9GtuWjsJrKym2p/J1VoLjce8B5OKld5ljQa01zd
OWTfWrevhn3awUtXyyQD3nkXjNeiqNxjAwKI9qvv15gtHI0VSavL3AHJ7lKVwAyuKXj1JqZ47Nip
AfXY2BKlaB3XyTytGjulHFy4J1IEtkE5uql/phTCnPIDox4IBK77RAgORfeE4tfcMNi25FTAeKyB
pyBp0wbNJQ4O8F3bskCf/XfNY35+R2sqSLb/A84Aq732VXUQBdqOtIEI4jMeVA28u+sqN6Q7AC9P
5pchCvWIbKfaQLi9yoOlJRXtwa1Ec2lwbQVTxRg7VzdEij9In1OHnyXMhNxbX7M4gbebM3XBpt8U
U4opA4D53Sla14SRRdosaValg0AmUgxzfDdmO3Z63GCK53o0ri3KK9eZ/rq6jm6fJ+c5ckurbzxO
BZTz6KwD4WwX0+SraehqQciPRh750xD9xfubTjDbueDIro7lQBZ837uADvaBLOZnaSeEMoFpr/ak
a7gP0kQwM/CoiDtW5QaVnDr3frgmSQvi+RW2Ma/YSkJ5akQryHva+FQkhGN4pOpK/gRk241h26/R
3Y6vsy0LVv2ptFYbtdWVRGO0Qu8iY7sPy2HYrybVTyugiUnL8Rz9qF74q/Sqrpx+6xLoNw0Pa9qL
EUXyDjRZB5Bf0Le4DfvppGhKpUmtCBuruidNyen5XB06JUwGRnPRd65zQ08r/QkZK0RJ6dSGrl8c
C6LlWEFXGbhRMwvdZot7GSAxwMXkC8ZLjk5Cl9BHua4p8iPBRK8FqP2/7bpnIqzuajxy/Epsxth7
K2LsZ8EnXM4ouWDhY7KZss0RMehDO5QWvkJKbHNtjdCWJ6mSMzOKCWrRTgYxh6YM98G8qi34UQ+m
P2gXeKJn6qMGWF2ZmMYR4DWuCq1S52jQKdtWSMEyTDmoQ8u5acIU+ng7hdRH8QtMz4r2jzEUgVH7
Nt13XshwxESLtMQdQgN1VXh/hdXTPUu2gc6L9QI2uH/QM2/oRmVjrAKhwuwCeTQI4fzGGnldWYW4
7rPrrv7YcdEZAWJWaE7DvrDnwUCWd6hYO5KpcFk7EidfTA1gyZob0PpmJ5pSxhiBh/l5BqrRfy7K
pqz1dcf46tKOW8VXPTE4gVDukt5RFdzJ/NpX0RqdfLQltoj5Zya5O2dav3dh4YE1gYU3wO2HgAde
Ex4jd9c58SqBJoTShIXAxjmzj2PbU1YN/CPXz5p/QlDtgv/goTT2yblcBYOliz8E0QxVPrB4vaUx
Z4cbuZS2x9EOHRduGQOP1qINK9hMhEs5J3lHnDuuIDtxh2bBhO0h8WKQJ4pAONzKexH0ukH4ezE2
6JInG5W+SorvLF1VVms5LZm/+Yka1+g01j0RFV9IAs2oo/mRt2FgqLnarY3Msprz1zFPGEOd1J2Q
LRKH8OvfxCSaYH4CJm+nBBBtlf77YWk/PGDKW0oWohBwSD+tYIVjQKTD8lX8oL46yt3NxiaOkZe8
GeLDekj7jxZYAkVEsp7FunXkAHcM31n7tDyl0ccbtyByyg/aPABmVTLTOj3Iwz51ED4+4/7rxulV
YIsCc4q5PR3RoFpcJ0xnl2Yac9In991sePX+8KrgB4DmBPRNQzGRBFwjLPMQEhH2Srb3oL4+mw2B
q5qEqmomBi/tzB8IujdQUXkbA/PPd2bW/o6/4BvS2ix+kwLzI4+eKM+Iy9eDKXdj09bDxv+s9pu5
VUgirC6q7e/CJLeleAEb29W30KTD2xfTQQfblopRbI8EG4Yu6bthCtLOtKleGPaOJX71+s0wXY1+
d6KNQSpC72T1hnEJNjYYXk6p8HfibfsP/whQH4CWRaso1PwCtk492n9zSeD2biWN0ZSlFGJDWWcy
O9TCm609n8GjdsM2Ablu40nUrgplkVfs/qWfmS58IsMNl3/8XNtRMV9KYL5Sp+7/PdUNnJA3DtH0
hbgtT6U5q+vM6DQOw1QfI/M8btQZ5CD7WvhFf06Cq+MgXJWiTAPWYgsREKjpV2FsRXvTlsPZtmYJ
3b0dzPtpHZRsg4ul3q8tYyQV2z/R/Amxg65mcKh3Ph9SuaNeo6XlsttjUKTzEXGTcqtEbE2BSaWt
NPf2KcuUATQeajmNS4BWR8tvq95jx/DmUXiEKxMw8Ik2bQ/p+aBrMhOKYFxftW5O0Wcn++PHghmr
Uci4cnvjXimx6ZznJakVtFAvCNjRGNw6VAcXeo3ouJ7NVDbZFeo4D0lXogWPlOMHwaMUaKnfzPW0
ElVKAKKQWG+MP5ZENvjJKt1rnqpLAtVg0yX/7b1wUwKvlrLLZZ50s3clvGVgm/3dwPYIYMteKfp6
0JGrKVixpH6jFmeiTVvNo1PsoSh3/U1KZyxDj0IlDSZ64CR2dZcb44bNuO8o6jT9/Hh/rotpCEKs
tLmEqUGN3yPOspsukchwr9jMvFyekpZ4wqXueDqkfZ9c6znR1+QYtce+SzDEx0JWive9oFSUEOSt
jdWiS61tOKMPHlvNMzh8Nuodb7nCQ4wb0eZ11e6r5P9d/R7wqweW+p54qKACPhIkP08j9OC2HXwu
UgNzoAVncih3OqNqzLYOObxQls2jIHI6Z1WV+lWFr79YgNvG/Gk/4QbvABk5X+cgj6VpZadJP1q9
pWAQbrctQ1ZHBTFa3OA/vcSPbiFjL5yYOnOcICI/jwQCnch0N/IcqTWGw65DAgXSI2yVjns7a21U
9UEC9KTw+X1y3msatnnPKIYrC3I5sYyzqV3ZuIQzP+0QbO4xPXUT0KWd/x8hDh4fp7H2Y0HP1ce+
pGW93/DAXb/lUXHNLtmY5t/mGAvCx+y0CJN7r2bCymbItJDTv910weCKRoLxb4txHDagyI8cwgOz
n/XPKvugWwBPebz6kAWCm2hxFRkf9MCfoAzq/HUlXGpr6+npqfszB5WaUq2y4oTJwvhBGgTrWjnU
YkvZLeIsKvvwiD5f9z99sxmtljugkG1WiaaID/4ZXvMUhcTpRT9lrPz0m91mw9He5ubK0v6MFQMs
vsDHJvZaN6I06qryGWJx5/5XHuZzJPpLB+PkTbSjphJRyvwLd8tLmDFbbSth7tussbtJtIcwf927
YmWj8/jTihrdi3x8AgLhWAXCoMLwLqxXIW5lK8lKulULjZ3znd/Pa/6Cl3TxXUZm0wqM2Y8L98Yi
sOFXQxfmSbYku8V67CNQIumClEXOJ5kSRqv4S6fBr3r0n2e48+LSkf4OTUzB3VCtvImIa0S54jsP
z8/d1BBOq9jiJW2scv6qz44Er0vlbozj2yAAHqpZiOxux+HoyRgihaUdkexeahZ8UveOD9C31U4D
QxK8jQgjD2jofDtfHSojKFyBQ4PQlwcq1COuLZ2UMLxTasMX1e2RioLUECRW++uty6H1w9s+R941
dmQ//FwRP7myMJWrCynC1z38Ruwt/3p3/YAljnS+tk2/0BqNKGcOcRzerHBmQpWS7mkaoZrtQG9v
uJcNRkwN3hOuNzY8Ix6dMI2zCvAV8Bn1VYVnyIhJomK9g6HtqMgrvRqdLa8SqQbL3ce3vh9sGAsk
gS2yO7Bkk1prdgvfOIed4Pfv0NEezrAdZGSBQvbAqAnBQmxIOsyZK3OqQ8h8FDL3qn+qzc65rl+d
V9FBaXJvbjGZ2M0rcwH4SRtGpsdX3XRuCTBem8PU019JLOl12DuJ6D3w9R27aTcXcR5Sk2m/aIBj
gqufoILwJuWli0oSXvp99NDJFD8zgtImfsTCpbWCFas1KvvrbYQAWfJzLlskmZmkPjnwbNrPKSKr
n0GvDW/HGlrnO/vHBuh79nQlL62LfjnfwGYNicKct5S+Wca2oRRnoaDEw0d7paduIJ4jOxP2HgTC
OfnDhUIV2Mitn1dBSW/ubYswYtSrYNvREl1u3I1lr8/vbG/mLG0+vHTAQSwOkuFi3ASdiqQZAjMU
ECfP1ZwNE6LOC3S3h2WOGgznZvPQ6rJvmpdpPrrsF+iglafiqfI7wlgB93ZC9izEX47tCoET8YTa
f749et38UVOF54Ug/jtDbMc0NIeo1Z8CGKIIot5+4nmDmNb5M+yNcJtWWEMdjdBSDF7EysYxwpQA
lLyzMZZwVZgkDSH+D0c+WnMDI7ysWS9S2Bgrur8u8/4v0MwTvtXPP/riGFN3OlfT0WVB/Q/HzUmP
p7p3FATq7nXTxnFbiyZztR9EGHM00fGECsVTxB1bDiSTUhOsFprqMa7jLLWRQNPHzJbCo2Wst/TB
X3ty46fOwHzsHVUMxLVhWvLO1NhI21QiUF848Ek13Q1yrZd+zG+sLiB0uGIdzmQESz4qlFQLMRrw
nmQbJx4SDyMNzrSkTvzIS7sVx/De5e1SvMM1MZgexNjfqBqT+syei5woQ9Su0RveDryan8OuntUn
+1u1fHbxyWBnyB0oCdUfzXa0Qpm2qNB1Vu8BbhBJAydWMFlkO5EeJli1K2ljPkxjMI34XEWeLgNJ
iPMVs7JV8v3HlZw61PLPkS1cqwk9A0md38TJu6AWEo6ROa7/Bqe5QKYICRl3xLiFwMX48R83aKcK
3CbP3MU1N9zXb4RS07Oof4GaaqA7fUFpFR7P0/ObU3JBV1q8KhyhysEaZ3wCAbU8oGbmRHBo/Apo
4rPPpZdQa3NsSJSRCBncN66Eamq9Y9ezq85yQNW26z+qTOmEN0JDe6LZ5pgsu0x3t4OIxWmZmdgO
Cg/r9/PQbrv6CYQPrZQTxiwyjmnIm1wxYRLCOZscB97xGeEDWJdtgaMnWRstoUtrsRcue5EP79Iw
YYrj02nx/KUQlzlLgRLKrZdy4vXj7A4Fn+5m0b08IHn7x3FxIGqMaAorSv170N6I0+KCKSM9SMUO
M+PRjAKWCGnj4ytaxVFNsCc8aQuGaoyIz/oDfWf6ryNecrvqd949uQRtd9YYyqgemSLOxhJ/Kzt/
4ogtlAxdTfIoq/YnfKuuQdQe0ILOKLamsfwF1a/yHhiA21ivHeO9ZsIquIn+YbYdLLkUvOaw0OI1
yg2P2w35fhm83Rr/LECtvJsCl5I8LCJ7bj9jlnxJzPwx2G1vCxdeMkjIHQj1wpy8Wc7TzlM4UR9K
pR4LuPRI72O7trKkLXyq8CbxD3tOoKnx20F3wtPpFwIFuQEe3Ymo5S9Qwocx3aLlxJwa0NWbuo7f
eSufgpRAVm7c2Ivi+I/EHE3/e5f4TFCHCcKkfqeqnuvf6lhTGB5UjEQf8T949MyiYj2OLQiVua3f
nfRCIWnKO/d15wlW6+ZhQSALQHWiZlUTg38TTac+i4WHQ/s+7hFIQSmPMntJlf9tYW1mlsLAUYhD
cBZxVNHoz7iC6z7blfgYR9N2Wf/hfIMQg0PtrSvYQikou3v3Lru8A0ljdi5w5zWXNChOubKF8G39
SoMIMfUYR8pG+UJlzBQ1DDmsFvZRh+rxxpT3xnbnkDERnoZkIuSS8fUnLpRKJxjuq40GFJECSXqE
bfisZ7GCpMSvv5RsEDN2VbZlPyUWwimgYRVHGnYlNgpSA3DIFIDaxdCR3l88LSTd8QaTyF31DsgZ
ZT6KUk/HRp/hAWHbzteoPWDPPI4Vu+ru35n3Jr9t4BAYudw2lQ8ocwRLJanKVqTfAJzOkIqQy88+
aDiXSTwmTV1PvzWagzm96hBCzOfcbNHjM6tYB89PEgsupbrLLnzBav+gSujxeUP7LcISn57uCi8b
N1WM50ex2Y7xep+xY7fAoPsB5dhSUJfddrtQ2pBnlNF/9RUq58U7NKWVR7lKIoQjUZ2Rhijc2tOp
8uzzOfEStQguL+T8Czt7C9crgDjHsmB9cnskZQ60sq0A4luZMyRQ0WWYBW3awAk/4ad42+GkGD/B
ecrlCrUaSGdhH9b00imINfWyOe+SlgSacaCnANQhQhqP8gLOfFY70DtSoWEx9MQGQSjT81dNhHgu
Q/acaczL59D7hvDUopjl5sRnBrWPXJcGbD6BMlOm1LWWzHiaHmVJnqkszsXDv+Eex66rMsHaV0kh
m2zOjqx+NlLfJqJj8FBXck8Y49XFFRTGnyECCCZL8dwdQzaanTI5loNYS4PxzRuYd62BKvduCleo
rvlefb/HWMiwtMst9li/fGwyhrBIwsIE1+VriMQiwxFkP1QQHJvIilVrmc2V3b8ryeY/0CqttwA6
YZCtb5YyUfXEORIcdruQHaapXLaGA2YJkm2IyUHgmOiGT8BTbzPzoj5HFbR8F735jm6PjC9SRbuM
/Ho9oApbdEGOPdRqXCYRL57TTYZh3r682lLsPBFpEZGefbib7ip/AZ13c5NTux+QUdsVv8/u9ND3
1SbWZcMnX/oAQ1PwaJ6/M4QrVuUcXs2Vvhqn04UDHFOXwHpxFzyPowcG0LgB6JyaKS067bQd7W+/
dLjuUJgvtJpgx7HDaGSnpdj/HBmWZKic+ZsiKuIsQLg9AuX6wdW5Td1Z43Zq9u+bdCfGZlsdCjXp
z47DSduGv9q5J2FrkNdyYcHRrTKpBxIJWw+jqiXkFEvqp952jONU4KWM7FYzmQsBHsFOZ94jk5qu
SqM0b0MnfLcUrgzaM/VQhVxlQqqkjyYnH+cyuoJU/UtqCxD9KXFXaZLFPxokYNUyezdxwa3VQA+S
DDHXFpsGwkKcQ57IQT+uKi0Z+uYc7POWT4pfI5QM19lP9KrlzxcGdkml/ZF/eC0qADVNNBLbSTAH
OhdRiAr8noXL7s16Gz9JGZLYXuKgYyCY0kWyzTBXTRNbCi62Hn9V2YfQTTQVvwJWcqzmVynHSDZk
YGjRQNnaz39O+FaIrFdt0pUNCexBwzLDeyyeB0n1yO7wMJcDr96USOG+d+9JU5ZzLkqXeWrmoz78
0pLEDKFALpMrmyv46ZEbJiu+wUxYbtF4VhO575cpsLeMBPLCqnO9+YcH11ddcC2i2IbeTlQPDxLP
x0E8xnqdKVl3zcma/mMsSYJUcj/Ilu7+hZG2Lld2FrHaY2k80CrOVY9y5jYSpOl21fH7t7RIx1+A
Njd64TJ3DRh6Ryb8zOgX9rRxy2rjMMClw1spgNualRxouuHGDE4CCjAIq8yKyA6I09Rwg1QWN79o
+/5mvlQ4NXcRhFN/TVHFK47vXU4zmRfo1DQyflOMvB5XGTtLJWQJo1H/xpka8hXWortSGyW/xe+z
bY2EMmsSlN2SQkgFOt+cl90ttyDY/TiJ86JXzN11nedtdxp4MpcnaDAvxEHmR/OumqjgydVcHl92
ngmZ+c7C1Bjk/Y13V0MC5974xQij3nLEYndV7TaLemB5z9GcLOY2w58N9kebWfoe9+8aQKEg16/S
iHepcrLJiSzL4a8Kfb85doc8uAZOvTY5W5bgxtNjFV2XMLaZ3Ge+qfIFs/zu3FyFnCK7mEcGEB1V
x7MHhhmxPVx0AiWIVIMwgh7c+szrWCwBckCBHDINPCWUee3zUDEGTQDoJm6K4+MvRZnN7q2ViTPf
lLtYo+iMLQa2TrDWTRgIzfP9MP+j6GiNwVeJu0CesEu5J9relaKVqYMrpJtzvEd8sze9v0RWSBfh
EZjwaMxXZra41JY6EO48r9AOfuRyfF9WwXUTrprjuWv6S2KJ+JW7JyFuN9EA34p96mcCCAq2ug1B
iWhj6t091lhXCJlCZbKTxZrGhAsGTSxwKZvbRtKK0/AzGo7pT4B+/c4is1OyJ795VhUtOHQt2N7I
/885MQRNvXTXzC++wZq0RJXk2AvNU6zMoFudOZXcLtACRJniH0BbEiStob8s41gPfT2e3gZ8PnTJ
8XXdh/dqhV11+2i3kcWY0UaFxMCHswi5Wh8iwj8u0YNFgYZWRQWcyJK03A75T2NKlqcTqkJhTSXi
uMNQZjz1tYCuny9+M8p4kX6OVQ0NGBgjS6zqa0yChqGbM8ndJ6rCCYmNMrMv8Lrh0d/zXtx7dTlW
hnBVSR74eaKtoVilK9ej10Wj3B9hmmjGs2BJ0MnsSOuFPgqufqLthveLMK7i0Hw9CdFVvIe9d68U
y837Aw+KpmHxwkOgr5ekZox1iTx7fkd9gwN1Ix/+4sx86PA0C4k3EKe/XO8uLwZWLRkqVqTMjig7
6Gl9oQ16y+txcfWNTZJNCliYh2nWl4bqAdv/NERw4dS0ywRS6JYtYQ2ZZdwQeERDSy/HTNt2RFWq
B+y0gCX1eua/cuXjpdtw6uf/AkVxFnOlZjZTNCmgHeTeAZkqGiVqfgkxNYmnNabcAUjjd8BrSekG
qUYsnEr6eym0eS3vp3v7+vlb/VqzQpb5LalGZkZ1A8tMDz8BRO9apjn/gg9222kWLo+3KK6Yqqlf
H+wEgSsWEBoo0KgjEC5pg5fuI5c9SfR7F+fZp2AgHsUr5IKQ0NmwOEy2MUJ+1VRUttuUGrPqchYR
rIqNtFBM5uKhrQTWsUB33yAmncU5Aiff3GSYnL3cKCsyRZ49IwWv4ZKAZWBsvJ+5DYOrJIXecVeC
M7YCR15FziAH6wCZlWRGSz2kPUUwAP1hV92+drxR6zHzigtMElWMACJIt03/dCle6rSa3Jc7r305
NxLvtuiGFC4c5Cw90fChk6vJBaUtxOcBrFJ+ZsL5drRkxT3c+WILocpP14xdXlevxIKLCp557ec+
PyYQdltFRmTq3wWE9Xc+J7r3yMajRmjP3uQl31Hmf3u5zgmQaMwwiuoo0FzQpuSj+a0K2MPYH5im
MeNTFgeoQflbbqqftG203ebIvVWfP9ojlB2PNptbWKDnEPN/AV5x4t5ztJCgW1OzzPnYvkjA3FiF
LCyWLl7FuhgodnAsDWM1/DLs/DZZPi8JQHd1+L2UNNntqyXOQJ87koRAF7U6lEKKYD6biR5LhKbg
DFunXliT206Be4QVxegPnhIVTYBsncpvhG/EWMbVqg12h/vqTam85/L1/CHv859fgsTMkVo//QfK
Gg/MDRxTEBDFmUez9j48AlnQUNdD6j7zwr1NuZwGpCpF9PSRLjBIc7c2AaNrVAt34AsRLdluVs61
vwPH6nZ1GAGR1ljk0UmDoS13mTUqr4p7pTxGB0YLBgz1XfEzsen4VgGUPuZyhzHS4JSwR7pE8tLm
4U1P5RnjsMpwPgUNDbcTPayiYPHH2UjOjaCj45YNL0jO77Ux0cXSKxqAQ5n5wgxf5CWJRU892lVy
hkEffqSd66MZh4j8Wfu0htV0Z/wdOW1SrlB8WCdwYSGVU9y/PlvU/HyIfHSM/SCpSs7fxrMwSxrc
fJC8ZEcvVcgCTaQV3XUpYzdeovJvjx9xmU523Z73BslQY7yevEl8UTDix8Iask1nN+SJbTsIjLRW
T5OUn7UZ0+sq2G8UkfT/kfokk/YHhFTRdSwZyZJjMWVVci8bcC/cnj6a+crpLlUaIBpbDWNlDDlV
IAbicp2BCrGAJvNEjlRxtkbpj7WFAeQ+RWnO1vXf8PR/hdZPxejlSpNC0Nj23F3OThjqrvR10e6B
i3P/3asycK3FpCvOSzPx8ldK7Q3Pld0j+EQMhnnFHZ/Pl+5SeAWDDXWHMdaYlaU2U3OwCa/drxNu
KoK5mzypvro4pRMrFTvpOSa5a24cjJcBCctc8L8LfGZL/Lqno8r6wsvtk3OqWrC31t3aQBB1JVOS
EIdZ/cWiKVcguC9i3XWY0mkHiLOzNFbO5QVUuKpU36jFYQmvsXq89/MHx2BHZO1Y6N7gQTd7Y1Jx
QXLiyMq6iQNEqAoB4U1FY+1XPSU46T2ude0htNDO+Deq5Xtv/ZqCqztW6uF5e3VWEPl5vnOVF5UN
TDWJYG+kNS67opLCLGUOXueqx780RK2XA2TKppoODmDa6Fc+sQmGFM/Yt7kBvSAPoE2URBvp6lpK
Z8oWodgofyLIA9G9AKZ8bieoHNv6plTZYsCIwbbw2IZmhWcxkuxFnJIo+ZsXbTWR9Z6llMgrujDz
i98g+mBhMuygU0PUQWpzJItBo1rRTnSrtwj8PTMHY0dPp763MlDS4HCln2VfffIV9Y8Npvovxfqo
3bnlsJyssTF9kNsYq5wKyF2K5GTwg5N/MMX9eXS6TzF+q0JW/FcznKA9afT431yiKpI01HfZqTlz
WNF5g92iYPCWdM+WnhvkPG/yafsZX9btlPf82ZQEduJdMX5QFGlg3WIVGGt54ho7E5qROVGJ4Psh
M/6mdWHxUpDGcvPsXszVDewY9UKOrj5JV1T5X3j629Ms9y1W8dXppo+rUD3MzeaM6+OExtdp9dGU
8Alh+Fr6l1RDV7OGltB5jkponnftbLDAZ7kmEJCw1PBH51U0Rol79VH92w6PV4CfflXMBVNAd1P8
IKWkF9u+ipAfVzqnHSsZlb2LIs1Z4zHf00rjG2A+tmhe/RQnrpdS0eiwbHPoIE+aHV9W0pIR7gZN
ql4rtdqDG90ThuPKIHtW8izhaEBUvy5MvxNnTZyeEC/bc6uUCr/CXsZTRJAIhXgfqYTY24+Hfv+M
pzwXGipAXDR60YtvqauS7TK+5ctWi6xDJSsd+NdF3bZqVeYgERW/rx/EH3kYhaM6ghpNv2x864pr
JVtqAXzeuwX2RLx3wCe412E83qN/OpUniBizXER9aNAC76UTcooNvx9qyI+vxOQcCXEfFNeKnhhO
Ory+15jai2T7orUD93LuqsoxUB+8Mx+zBm54d8cyQTvQuYIr1H4JHtZ6KxzOosvqpyf1RqF18GNQ
8re0DruE5d8kTM+RJJW4wh9ChNOOrBFjiR7UIT+IS2svf93RtkZhuctvxs9qsD65JRXijt2vTg88
vu8bVf9RtlTBVYme2pOSJuS821+CMxgFloR2ZroyCDD8nBEsEkrvsozWJFQKbYiMhh6fqP7KnHYx
D4RGebnwGxcSg69pRT4Uf6gIK0ipUGI7pnE6xW6/4aPbIL/zkvEeWJ97mnTHNuENyZ/TvzX5URQu
CwoClTx8Ja+q8llaR3yI8fPbUo0HpmMhOGe0fC9IjWuT61bCcdyY9YY/jKECf3O6zt+2LPi1Jkum
NAAYwigcB9hz06tFzIxhZHsTk1r4X6IHB207X4JEhFsNLQetNMEJteZ63WSZ7ryH45dKtQJk4jvj
A7mf+tb7myu5m4ulTFmnqSCOv7ZO/y8k3DXVwqhVWS2zT/79gYSlGcUGo3wTaPtbR03VO9iQTZwr
Sk5H+R7OxNLYvSc56iAZrrFOjiX2EDsBxlheQ5I9N4sbYkU2ALNFtcP3kIKpxJsrivLwCaskolEi
nQd2LCSP3+s4AP3zuPWIq6Be+ufe36oL5jwwmcyVdqPCAw74kKmgb5AvvPGHb/3MGEavU2H8ZSrs
23jZVmqsJSzK2gHFbNPgtxFY4OzNAHZnNtQoZjKZgJdivTH4RvcYlTMXUJWY2RcSCP0I/GDxeSOM
H6wCjNLoBY+pZaDRsrZoceSypearz2xTGyo2nBSnmnyGEEA1iUaegU0ni44HICTkfCrlMiy695Ww
9Y+R7+wBcHtgOKhvuuwvHqHvCMj5ata68cUwIOxAbLEizF4kTk0Dy/tlUhZpufL0P74GBOnT47qZ
TNYmejS/W0/u7VhbnCwU95pJHU9fQZJV5iJT1l5STi1gMVEtn02zduEc6QoGzU9b1cX5OljBD1DN
wAtpe8575PxE6a8HbXP8UhCPpAdQ0PS6owvvoSok/waO0Xeoc/FiYxfUD0fU3HI02GzEdJ/yjXmK
PH12s08eqE9Ibz178TQf0QPyUeYXRlVfWOKuOo8aISFoFyMft+wCn6eU1+wo08uRXQKKk2KXUzpp
6WSKeXHZ5uLi9M/nGZsIPvCp8PraX/aVj1l6GBYgcA3dB0GllKlmnXz3Vq3aMQoaMhBqIljw+jrH
o5/a0u3Jh/B0iBBgvOB4CfWdZOmzCPAkI233+Q6mh3MGi8/H1dOysvaJ4+G4hvUF3wSSWuyWO/Wv
3f14/D/N7svhdv95C+DZ2zf7fbBGB9nhUz7/hjbFcIeyFf0X5veFBim7Z9JAWVp+8loYXdsR6mRO
yzi7CUkt7FXvZBjaHIzPKIe4lj9HXaIyzZElCe61RXXQm/3fPaslrjtlBNG6g5BSE7HVczacLoOt
367fIz04Mogk5LUJLlSblmhj38q+ID2aPv51FwZ2EealQdC2ylI+tn6rSNi2clHP4CX0nLOEBT9c
SVNzv1YMWnmeKUPheSBE2++WudJbXvwd1dSr09lQRgwbSb1Xm8VmO1bngLdk9Q8dB3efdSn1GvMN
AFFaM/qlYTRH/tIHHrGquELl/+uqMNia3ZbJRD3finTbcbM5ukxg/h6q90psWaB19QINuPw04aHt
oW1Fae55HtKQmu88HNAb3Edpn0V0efwBOoujzhk5S0ADlwwdVDzHoDg0Joyswk5yeXNp1xxzRImm
EUMioizlJyPuE2LdLjj/zb6/HMH8BAuaxc5Ou56BAOH/QeDbILHcKaviqLL5aD5TSz/5fdtmcD0Q
9tjUGRkYaPFyoMdu1/s+9sO1/u6HAyeirS1QempW3H86wr1nHU2QaYhq7iHidoGv9mqHjoe1A3Ut
57mb3ypatxTTRLskgsa1undjih4El55ngJLUIkrRigz1pMvyGUUoNo/wdwzlrMmJVarWnVrDYyWw
uU12LQDaF7aZURMqz6pwkY0QcEvzshsMkxjGumuK/7THo/5bUDRwKR+p7W9pug5CakcZGzSW31VU
k93lXCZbBJ71DxUlc1AJwjT5CHfIe3jnKuYciQA3rmA7g3dNL740RSFNwXFTHSS/5sxrKq0YqR8e
7f81yRvJ76MlYq0ZfqH6bs3+1M7UcZ7daxDBCnp9mBZ1yCJOpiU6fqyFBMWttFAp9yHtwb3LVoZr
zjHGQMnUfh7FDQwfojUj9k2DhdFyWA9ml7Y6reew8RSHKrN4Wdk2LKM8VnnKlVEH62B8+znARnLa
sRwhaYVZr0PPlY5+mH0S8v9WHYDiefOwGfnXpqtjAncGxhomygfDW87Z+LC9uKittXhBaOb1H81t
EhmJuCaESsA6zDA6Ej5hi5eyUj/dyz98hOLnKX7NJJi30b2GdRBVgCFVaa3dkVIE1Fh0+V2ZFyiX
4Q0GkKijnpDzHoaajaco59oJ4WHt0eqJlKIL+w9btDkk4RppOk1k5LgfuFVx6sevDwd/pcT/crYB
1pRnh9XHu5SgMDNL/hj0twPwcJY7e3uPO0qE6IcsxFSvpsWZ3k87ym8o9Kl13mJfvltB0zYfORsM
C+hPhTB7a1FckhygJk69ObAH7zYAxWWI039qXIz4EjfqYMMAOX88mqdxi4vzZy5xojsEKaG4Q/06
uNNMolq67jNh0Q222I2Ka/MtCBw5VOpy30L9eimS+lWtUbBigUXApKF79yO5uIbGYpUBQUTe2vAy
V8t7CKF51qemt9UIcjrN7/0BcRHb14wcNtH30gLZsOmq/AEEcMqOIzQuTqFSeXFL3CYuQyRibHd1
1P3nzPcaAmOw7Fd+dlSnTI8NY8aaYwqxV3yQTgPqCmjGt5svTV+G6SibNPOTBScGwYqI7g55petE
QCmLgZY7qowAxcAJHMemkDV8v7mUFCw0RQQIMEnQaY0mIk/6rch2PBLCm5e3ZmKx18MSEBfmsy0o
tDGSFo+xZTnxIA5EfjGUa1Hh8PHLF3BfqkgvX7+TJdjOT2Vv4D+SO72dCLIRm4asHQ4nqZvaoCiy
c4XWqfmMpa4elL0vGIzz5ByMe6x2ETY+MkfGBVAdwOXhzLoJMe2TE5lcXjAEANUvb2woUkqfKcVl
JwPLdTPC6GqDt/d87h9zVgT9TrQQ8xJpu30H84pgzSQJXT0YnWcz0HcFXIXobEjVrHPs2XqHdP3R
ONlhIPEmmgtkHSHJqotBpRBrSqVjY8PKvqxdiWkWAEokUQRL0hJMtQLVw7ZXXnpj7pgtrwHl1xlt
klMUnR/i6TVRVxkv/IfEURHCfmKLSVgdeZ+Ej4N9h7CYFBAKiT7R8wIOkVvv5vomFgNbL0DH92Cu
7TmMCZRELilCr9aT4HFkVkrEgTGVXN4PXm0kkmKcDdEBVxdQUoCsE46hFJ3n74UI8SLU/fayzTCF
UR6jkpKDUcqGVZxGu4geiF3lfuVgJsCdlq/V86I1eIi6PT1HOJzV94y1OcupKKoxnsBLPoTngtcR
jntxXfvYYbk/QapSlbQVmR7zGFkNPXEY3fBR+J3We9hFT4oI31IAQQFeaP5gFxS/2MRZcKMVBotb
NlKpGI37V+6LLo4XcPTCN3tKB9kdDaon9QHtu9e31VdV34fwD8uwNnmC5PP4Ih5ROEM2gWXrdd1h
BV7P9lk4TEZWx8Ibpl8pTAo2TWKs6MPYSzYpsPYtb4WOu7HJEbC0WDmY5D6rffHJ9egMYyspsxun
c1axaoBNpRkFEK0wvuWnUA5sizpj6Ktby9fun5Q3s8O6k8Xz4MdykT16+0MGbn8W9HTL4LT3Mb6V
DYlD+JlDmboRbIi5a2U3J4Q+N3dRz9C00IITdtFuY0oYorVlWAD6bBGtIFhrOq0f7ULE0f7dfLPZ
0juuHz6w0ewnAJ2cr8SZIw/CDlRQfMTaUOCPHQmsME13iWDqir4oqc34Dk/M63z1pFtJHUhxy/BH
tXHdWWc8vic6rs2ILkQ82F6VVsiwQKGAzbJ3xXIZLhLezSbcN+PwyClJeQu1EZ45RmRMLCIXN+2S
GZAXFZ1KvURTSbwvGVhhqOQ1g7NFn07lMXOd15TvXEo2a55l11JdzAVp/gZTWMHeKWc70wAcv6CG
1a9iGfiRIRdiEqrACgfVv6oeFfnYah8urrSoM1agdpzdCFMjXb9hKyyn6yVVdg1fwwUATBO7lpmP
EcVrumLmFEyQWu6+LWwJJ1Kuj0TIihbiCAZBVD7NrAgiZpLaPboN5dw173qYqyW5xVlaIFXE79T7
is1ROKgFXLK/x24C0OE95763Vmv25ZM7V5G/sC0DYQvXCqbrvQKJhmOehNfTYe0mhnpLnzzaGtMB
lURprwniWagBUmEwwbdtsIatxTkHqHkCnSEWDUK6Os1RoR6UMisB7KnAV9bNILylTlQM9B9aG1On
BR+M9W6JMI2o7eXPYgwKgBbKLnlSFucoGxITFSkzUalQjf1bam7ZEhPDIXegcWl/CMBO9FvF976L
HkxYu4MwcETRU772rajcY9fKIc5+KsCn9McLbanu4IyY11dNXZd9p4M9zqZi7oic9qNztFE6E7A+
k255gxkW/6Vx1iKAMtXFkh9AQ2+wTl6LTS+vfENl7BLH6uKahTp8CMKJ6T9ew0afa7hzB3+UGHI9
Ozwc6KVCWhzalSnNpYUgqDJhHffZqjAKeA3It44OpIMHaIdteyYzonKWmyPOARxqzmUF2yOw9eId
VJkbdyjbjq2Cx2PZwAxQIXG3JHx1G/EJI1qA65D2S1oI3KKQcI/r4Zt2pHd9WSXqSEb1qlCyRULY
tVC5h+ZQXxSxThLACWISAkzN7U9A8WmPLC+jhvCr6JeruZKoqnzpRMvqpt7lhvH8cwfQb4Tgw+9D
cvjK/FtE2sAo0B4rsOIhv8gE339Pat2dw5J3jgOXRau1uYuV1/yWrpKaJy2d8JQjq9rHdtm6EuQE
+vMohcuaOT9H34l6cqCPjaXSvT68WhLVUn8BcqmYKA05y1UjmL4r+U/BmxIIQYrAzExm+7Y+xCME
jWJtLaMQz82jFOCI1Zh5PakiX5bVqx+GO8zWDY5TJy+qnR2uzK/LuFUO6N+EvXBMwBeoj012ig90
axWkOlq2kTapwcmCpJKumDG5X2mQo+TdIW8D6u3wa7D0ICggV43hI/u38jRLQXNi8ojfbGbkwRh9
sfWD2DutneJ0lxV5WKguVK4W6IOJHH/C1fa95Py+k8r1hEp5uRdoYF8rciAQd68k8qsuN/PUC6Tk
gEQkVoV2YuT9tB5hB9sq5E63DsXblKzo8ZOJUkhVirt6p7dihBVnt+u74ogOI/e2XYJOioSLZaa0
uqW5ndze0WroOZzIZZRXNz0bRQG7CNtDLzPjN9yjkWWtcomh/hbEgJDIXGXPJmX9XPTfAjx1VOAf
fjaewEox8/fvqFySEPHdts+5gyauuhUrp0Y3vekzKSLqJvq/9AVSGVhNXMaAQ138gUZiMtz1a+1z
jts23k03zuYvwftSfNeDAtp8iTnWKXcNesYjRCePgErf5H6zkJrA3LJKEtF6wU08Olq9snzz47T0
XQ3/f1uNYvhfUhaKyxwirVu8aKyUOQ0a3dFD5pxGd20c6aQXgCVlZJwqORMfHIi/M4viyjYy5vaP
ccYrxmXT4CBRPO25dZbwTir5fN0OANB3l4ZoZpyCHhM3RoJAna9++YhAIe3lNMqsshtOrvOtB6xz
pCRopwnjYIAswULLgl20mpaEq50IqV3hToCMAu5W6UlGikjqW7P4BUCRbuDAVwew3FXkOPTbfn8I
a7GLKZ5VejSPqKKdmA6GvlakABFG0KhsVYjT+He1IHMQ+w+QCtvL+1P9tAa19JEhqenZpbcFth2m
tvdYhR8187imQ9epJ3K7zXu8b7UNs+1ibmzHhFyaRLJXOgHu4p1B8AsilWSjrCWhXyjpycZ9y8vM
xsPOuViizdN/vzJPG4aocudEFyxm9xboFzeZDtP6DFwE2YAvf/4PId6lrAT01DXh6iTqLP4wC17E
CkgUsfakQwhg6ovfwGn+hHjaNE8gH3EPAgWQGzDkyi/8NNtozU5ojhhJrzgNrq7hZWLVxZPOf2Vr
XHasH4B0qPY6UzhLn6l5LWfmt/l+TE9iELaIacFj3Dav9BYZStFXUOe1LXpw21zwNDCZIF6Xe98t
3/+9wpFa8en0FWSpDHbD0vcHnewZZ9gzHRhBKZILmCAdEhAQgKVhSrvJ4N0+llHrZIX/C/K3eoUp
jqE2ykEneUx9siA4av0cmbLgDlL0VjL+PhqYZPdIeGgnZfDVOguOOBrpprMWUBaHYV69fFqWdNUJ
YuIB7W5khqg5krNt2dTEdoBpf3C3HQ6w13rq+Jg2pwuuWwYUHd5zQPdEkN3163AqU04EJpx9MXfb
9zyrVf41FNSCrYo7YZ26RiDtlWVtUv0zW5KfXsYPgvoHMvfkxG4OwCVmDc+lyosK/6+VoM8ZoKnQ
lk/hOxVzw4dt6lPTUGphM5IRHtHJJ+HC308EnBIkQYTIp7H1QoKKr1+H7LpnWJam0MUln7JPUDL5
TyPq8XxQHMXA73W/N5yJBlYQD4jUcQ3LvSj7COBZ/8rCnfNajnAf0ofVpZqsFu8hEayavfmoiUYC
dy9CLZY+Vc0+MDlQWxzIwGnSxssGq76/+x0IKcI8DuZhjYUed+PFNmzEFsG7JzsJvL9keCP4MY10
xurjxRHq6ffYOYwR9r+5/U+Bokp3XFkIyFxQCtzm7i5c3dlrRGYfbtFKMM/2rO/d6QGabe+G57in
L7l7NhAaKiwwxs30W1rmHKmqaaqcPOwH2NkC/EY5jnki/z9YVZLhmKFeqNPy66J5g9j5BvkKYQt+
JvvK90xUoFvrArrF87/YNuGiwtgwYAGSStldGN51De51K3AtYtyg7FQlJoMMTkb8gXEbXWw0QazL
59iahGXlE6Ekr70RQv5USbWzhhTZac3C03qVF4IaKo2NfODWTRpMr2OCEuTNksX6jF+zixmf4u0m
fnFwhUdHfyUZWDJZrlNvfw9fQS8ScFn9HNh4GrCe8mNq411jtsRPqGKT2tqT3o60wQV6TuNzM+50
OX3JdJSPunpbrcHgOzV3DKpWg+naSBlxidgsIdgCdWhQsYST/Bt8dq/dkOxagj7f/gVrw1kuKVEF
weF/hmsvODsv1RS8JT1SyRDwDKlqk7GxaFyk0IiyzhSBQgU+hNmWwIpm/97bBSFhdg0iOKc343Ym
AOQvMjKYhnbRj9u3kjeDj3YioxDT4EP+jB1LM4oxzmTujN4jOFx3AJCpMl3mGJe9nMMhois4t097
kvUlN0JS8RZq/Hn5sNq50YFA/rtomQG9kJ+S7N8/ptv+EkluSlYQ5twT0AMtjYcoTUS00l0XDk4K
wYxZKTTb9p1YnX9rUt610JErddkKIuEpOoKJtjVIJci3DbnrmtlVv9dJKtFvaSqtNyWND+sH6vnm
1UcDh1iTyaZKnAmDJRuUyqqVG8lJpJX2jDMreFanWD0C+SpEa1yrB86GnHxWKjB0aUgSD6PrEFOl
S1GB2VFTC0yVB8y1X105E+XeaOyE8mJCPXvipJXmgOEK4BAKSxgygnZGWJZuNILSImVNKho9LAoh
T4kgBnMfufXIiF1O/l2yfLTrFkz4t5qdGsdbCaA+SuHgqSw/0oXX8dw0oZoR85mAC8z4dWJwt+mf
Bc9l6cQfiYfTSKdaV+Zmk+k5j4Ip0lbCnO7en3WxT2AMz38mrTHKT/TVhryf1MP29kQipHbHlbTD
LIs7oaA7z9ZXCcgdPZxoNL9RRj4gx3cGD1be1t34r9zadQwyxiaFpXWiyujAPsOG4PIufEvUi1do
P+Y95KgaTqTF/qX9FvGm/36KufRgPlcOmzhtBfKD0OVSGvbhUY3ZFKvX0TV+v0FBj5X9q/AbWu3y
C12yTaCMMgkhN5PNosu26Y2sl6M00s3IO+HnFGOXBOcQ2qx1ivhST6Ri7HLav3zfDuV+zjBrxPVo
V95ZxHIOpivPn0pOTF/PEIaS/myMJYXbdzSBmG0urHWnkwAG5XUU5wIZVb2A+PzoSKqnMzof/++Y
D+1ScihFMtr0oU034PMH5txWRonzAnQDKjQQQyufzzszi7PVKARevyXWmHHaQHEx+MD0C1JK5LMU
XLPYleudXdpO2kpouKziBBWIWopoYPWCRB5IBVD8WpH0NEs3n9gIpPRyR8NWJ2ouGSH+w9vDuM4X
FIETi870bSkHnbp/6Hr03mCVgSMIrVsyhHK19PsHdeMiUU51Zu3KcOPgpT0O8g3Vp+mFGdfzpbLC
fY6M/twM8fhAtWtd2kApvLB208HTlRa+zqTDqbvBg4XqxjIPNopTc7cKN7raS0q7MuedAHBZnoK5
LZU8pSsdPS7m9w5EZ7Sv3k3h7NjKO1mxijAUI0A+fAtLJk+bP1w8BwLwsj+jBucZixMq4siNIIhG
SPOoBbjeM2Yv06nnYhoVynmjvOzSBYzOsvSTlvj9CDnRKs0M712dbHCEyU6es1zAiDAQMxlCT0Ih
rY40oPzFA4/nKtc98JLXqwShgVuDyQPwnpqnUvHhoDORfcSnOtExA/g0ciRQpgxjFuWKMgoN2ZU5
QPfVzpiDGQ2Syo/Rok5u+C6V8B2cKIMlr7nNecZSEKghcu2QNssrVPb4RcihD5gBTwkg9qhvOLrH
AoH7DXA08zcdXWPLkP7bkOVSGhy77vKZMxMlAk7N1J8G7UFc3rht9lMb9tiZCLCLd4qy86qx+Q5m
eZW36IDCV0YoMSwiAdMsKEAV0618uzs0q4yfg6q5fSILfYM9pKGxixH/98MVc3tLpvmnYXMxmdYB
H/HyqAX7cV668YRJkeooT2gUMn4DNKAtdMtbg4DGftF/TqfxbaarLDmB5PGLOmo2Iwq6Hlp/8/ux
ybQzMe9PY3fLN5AOAKW1u0PpuwefkWn0/WhY3zBp9sGJc/aJNEo3R3aisPy3Tum4E9LzCyLn4DoX
KnRJLWo0Vo7y4RG4l2g105n7ENlogjkR3mu3QFSp5wzXqxnnfXwXijcqPR4NGOKI6qpBsP4fbIZr
FInhvQuB2jqy69cz97MuKS+yfDan5ksamwjsN6zD3dGQEB8ZRVmLtI6FfZaYd95p3fJYA3AVGrrr
VofTunp+4QpzQSg4VslrWyN+zh0Zkqwcqf0ACA8Vq5b2OppwfMpVF62mXcefoYo4RdwvSaFinjbi
F7OKiNG66XSLmtLjkB5m0JPXgW8g4v3f5j7xQzhh8a0mKhU3XtEovLtFZ7/W56Gl0HlPFKybfNHV
52qToXaoo8JSWOz44CsyhVTnU0TBmV2oIeT2Mm68RDqtRZc1SCb/LULMqWFJB2uhFEhUTvEliai3
khKn9ExW+5SfMKe+sNrHcRybeGsw+KJzfBbBBtSKg/NjJb255ibCfo6xSsZGg1NmZHuPrZcwm/1R
hQLKGeD5a7xVddbftHkh8fYM0pgeF9BpZK0InjsWshPb1vTfTVg2Cj/poz2zNGzHgkSsEpdgJ8kk
JBScC5ndu97ajUlSxy61Fk5p5PkmAqVrzaNNjF0Kz9dImhewwHD52nYHHbequZcqBBk9bpQGiebl
exMBq8HcwA9N4szBz4I14lQivaxoLIPhh+XxHiUY/J3OehuGM+UML8pY/+P46s4AVILGAmO9wj5C
b+84AYFuk2H4eTQTDl+NCZVTC0wH+E+asKUcQDnHo5UYtaQlLELr7tAmb5x4zHd9OZM0YKZYCDCb
mWfHOZTvKFniRW2OBlAayjQuQ3dZfltNAFAzC2iC9Mis7Wa+kzW9bYYVR4XbSZXLOJ4Mx93XsW2S
tHKgeCaosearO1bxKJONc+Q0fwffc2ewFU3Bj1lLLvgIHr92V4FkE/eEiQNvtQot/EV6ulDgYpGe
j/xxZ722CbWmMPw3xshlMXkeObs9emQCU0E6gFT4tnO9wVI2bUU0pi/AruppdWnASpVKbLxoqCvg
n2qFVQN2ZVXzYxp3fV53nQuWZgeQJo8AfU2QT8h0iOJW++Rg5lxFEIfIOaFIOcz/eUET/5tddKt8
SQeaHBro4wyBlo5JY7jKJ7mDrB18WkzOTN+/gSH6w88j3qzKwsjFtZzErXOelfnMIddY6gfXioCp
Ekb/P673ni9/tiiellEazI3U6c5dZmvrqT22by52WNa5CLhcpMWDEbUxiShuz9+SKT8GaG/TYx4j
VeKh5wLyjEYrTGLJ7T0J/Xqr6+KQUHp2+tDbM+FUYPjSa9VXN3Y7UVzsad5VRuGanJVCb1L2/FlB
P5Vcl5rdfXfuGSWNJW0bV0+s6Q0L7EkN838GmVdKvwCrXfB3nCF1vrJODYXtDQbvO7zQE8pxI+p8
35RmConsi/3jMnUZVCUNjWv3uCartC6VHUeoNKw07SEAPyePdK8EY5AzlAeQvcJjfi3EGMKA8n4J
igMNDeTVgsXK1wyAq4lkgPnkU22Gd7b4OR3xoNiIIEENJER6WaHiTQAEOOPZ73eObqTVIQ3XagpQ
E+tPlnS2UL/tVMPksufH4picqKASizYdS2vZ3JmbTD9P2izNGeFamC1k3LFLUuN+JkFfM/l3uJ3X
93SIWTSCAas/YgPaGwjdpJVt+XpPyoto+Fwj+xrpztAQmkSaxTut0uJAK2USM5Y+MestUELaVToJ
8cOATeB3z8Hm3lZ0OuLP47mvM4A1Xq0Fw0OLAEkJbk2DWSuopLaL8Au37uMPib5UZB1ICCCYxyMu
21qV3CVMdbksuLe3gJ7DuAeXd4tmQ+ZNHjS1wK1KKaIac7r9Suf0TNsdGk1sS5fCAIMdhDtgPGKN
pkxEpFliwlgpxSdjLR2WF7BYeJ0prLlSQLFFBQBBfA8hbIHyctMF5RGUf7OhmCW/u8WcDVUoC/wL
xrdFGBcR1IqRjg9QJEH34Phgu5JtoJ2w4PLVLrrPcxUicdblLhsL0xLQj20L6f9Qcrnqq470V9fD
S9oo0TunYEE5JA029PPh5L14ZimJwDyvLwaLTbyOVf1Folu1gAYBA3ZG24J8uiDW7PjQCVC49Gd5
9U0zVV0OBhBiC1YphABnKT3XA8FdduWFVLGluWZewpzUBpZAQpDIr6txUBaiPDYaRMKtJO+DYrGS
zPBYMY0v97RHSsGYOlrNUz80kovbFh92KaKasuWh4jSFTR/lE2+J70CIZQvEOOIa2/WQeD/CrR0v
zdfbn/6ya1kCa5ivcWiz3B7xjrGsG8lyTFblOkrWjwZZKD7pZUysS2zzkWZLHMDf3WWSZjXJ6a24
Xtn0/AapMKKl/cRxmM+/VtTz+ZUfZroM+a2yahh6Ya0V18VCN4QC4w6gh4BVTMZlATEw+XBIF6yi
/tjOPqxUPMuzhUuVCVt0QBu4FhI1AqEbT6gptCH6fDXBCg2ikJeMIfp1mTPXRdytq+U6qa+U7SDG
SQL4/ciNycA+XzUwQuMB0QtKEDL9zdlvBchDWH6lhY3Nw5f/OE8K05Z6W+bEwH9Uh3NzTFUSJZAG
4cjQX3zEgiVVCtVVKuU5HdiSEkBMJXpiVzJSNRj3/ea4LB0g547wVCHsNath1xBBrZjpd8GEousm
3aysXVA42SXbWucLAhEChqkTCqhT2fiklpi+1auH+T7VmwUeyKezkV6RKnP6xCf1bCecUz/m+sqJ
yEjRZkL1wHk1Oew+BDOI0VdIUpdmmGEIURO766HJzQ3kv7Ssq6Y9IBuS7Vw9aaXtR9VkwhXgksDh
sQIcCaYVNEwtnfo1kVDdk3Ntm1BkWt45CzsG7bkGqp/gkj0sDi9+b7uy2k/cSmS5P9oyN3Cnbuon
PL82jpyDwEKOt9rMgMNxC5rqZNiTtvyWguuogF9MsLeNalIk/mJPCRNWa5Dm2nezUmc94Qn3mCVS
hSDbiVI8UX0893o9ye9IHCUI/ovZfv7YTy+xUWQT8M6eAJWtpawSwVxwnY+cCeAuKAvYxSsmAX+S
MwjT6wnBrDXjjE2b0/eAEYyHcLf+qQ6CqhDSaXX2MWXB6m1KXWZMaX2qLK3jyZc+zeSVzNlV2qI/
nwHFsQryREgWQkhFXhJi45zxgQZmq2nc3p/b9AuCwdJC0GuFztiG2VhIDnyiWhbuFEcdOmLHnjHs
rJANna4rZROtjklDN7DZXh1LXlHeFbDPLGxqe4Xa+CELUHiw6Kuntn7RJfF26+VMbhn2IMXVE2Mz
7d9/Vg8w95rLi8aGv1ONjvq+Cs+SV7DNShngw0zX/GfRih2kivqRqoLTjL0rg+F+xiTplovVF0Ca
yoItmPHjIu7E1kqFopVr9yVi0bRpu+x9925FgKfFkIvrW6lCQAGLdlHHufe6Lr9fEIQkVVs90k+h
fP2dsbiWe8Ueh2OHkPRZUFvrPO3Xkoytdl6jrzXV0CrScpV/H9K+fcFJfdHxUFjZ2np43GXPGtz1
4dpHeY0SuTCPGZ1IctPSeSJeFSSor9xuEmm+irX+gntCJbIdVWWJTVI+BSjLLJdaCfVIbjWoEeYu
D0ladjCSy+1ShtMfKqjVzV+uDp8l7acJGpGw2rHvXwdHFY/jrrUSh7nEb0EAEJ8g9g3nsbPESpqo
ULdPtyjhxKfaCYeJHBy5z47fgV+oDONVha8P/jrgMiVnxoAfkxaHmgxF0t4srUIRyk4CjHxDGMkA
Lq3eBWDkcvzVULTfJL8U8AfqjeejPAPj0Ljh8PGKcDQVML6G1NmD/SGQzfqsW9b+rGZjAUbMLF6e
by5Pax5oMoklpkLi0LfLapyBTJAJeq803Lju1rCIiJSoOCaqimzVQJZ9dQqBz9WCrmxsBH5x75Et
77OMJ2vRVE0+XYrkJ9vUuZ5TDWeDkfmg1WCFSbfONQ90tvOJm7G4vJZvN+Prqqh5ZHH+oUfHIQzJ
Tj1rgrbRIeGNTk/dNpnmT0Nl62O6DRGClUrS94+bJ1Z1/cLUHaSEf03y88xYOUZ6PLIJTduulcQU
+XVNIK29Ap9TXwKNeHYZNjsauTpOqta9uHHgLy5pr+fBl0kDf+XWvVclvRLo32wZX3vvb+PR70Mr
iNo0Vsd9VKg0MBXibx056UWbixOj0bcVLS5CtZm+yd5iOl1+SBwxqfo0/dU5p7AGYzWab/VNFupu
x/gmheUO6kzR+2UY9ZaHaqSEiucXz7P9eaoGe44ZTrpij2AAjFPdNsZcXCuPsqSw85Atf5anLt+g
/JgzKmgFnWxLQeGUl1rnWl6EivuIQg7ePqGJjmUaIFbOwnl8alItoqn9k9yWxOvk9fxkLFcKyGyZ
XbkbKzhlusSbk9oKmUMd39QhleT4L1cabIwebD3nivbD6+vlI/25BSaFVFEl+3SRMIyyLDcd2By5
Og2Xp7Egy2QtuXlLO/dP26HVLqkfgWljh/rItlTs2Q8/2einsL6RABTxRVsHuWlapsGpKqeOIl54
pnk9NbBQziKLCjMd+iqVY8UHwohM3fZvug8NaS50+gSbr5f2+a9XOqf3Z2SNt91b//Cl+NHFXkVx
L3i6pKzBi6CPNHtM/lO7u9WxEd2iunU5iDJQZuFQjajAqQFVLwQVrmdFe1GIfh+0IaDcIpat/R9f
bf6AJEFHAOet7AmlCMTqLkPWfCD6/SonAHxNdUSKZ42S1WUp2KP5Ud+W1yAorVA9JLWQEC+H/rgn
ra3OPwQAmFkmuDAg78pd2Ezr5GtYoiku+cDmvMY2g2TymWf156c3+KXjubxle1V84fCeXBaQCgRp
7d0QPg2kOfnoruj6SaC3ZsnJMD3GKFi9bl+G2r1ZfnCoVjmVcDRgG5f5Ol+rbSyiyx5DA3L5vpJF
fOoJwsw7TmElgGDhp2GnvVlivUyqWPjx+CcJC3V3QKup7ugV9wQxpsDa04A/ahh1t6W4DKlh1lWm
e6Bo3Dzr+jGiQJf+OTftL/9g/jOAlaf3POyY4Y0XFs+UTW00oKhca9rwXtfsNMx2T4ZgQQCndY5A
YZnR2UrwhVwOlY7FcCqYSEEBNeP49vaVWLPOY4Xk6bVjf6E7r8yM0KVBNKJA9o1O+AsPBdR8iDRQ
HtOz7Dh/Vf2dFuFra/HgBWd28bmf5Cj2urw6GSGSBREpO3u3SJirmBDpY9fvvWFlJcKhR+ULyQ2a
4+IzC2bCl+5vK/2d1EfwWJTdRm8fN3qN/tm0jQMPuGS9ioRZurqJAIIOw2l6maXCs1zla11RbvMl
FJuACv8ipSI1x+DcKRyWc4KfUkhx6fxVzhVvCiwmrnxSdaFg4eHq9R0OB/8uyfdnipcIY+fwrPRh
tBqpQfJoM4Wt/rcZBavFsi3c4l89KvDiohgEf3qHnhjNm4sU7RhFar+sz3in+N/LoNGzdkYeMlxa
pEjFnqK2Gy2BRHpw6NHpBSKSoiRLwHGVRFPPCQWl9N/9PVQMhCXPWUWtbDizySPoxCZ6u4veJVY5
ZkK2p6fpA7HfxQCYKbZQrRMi0bpHTdFqyl/9X7i8WQENPx3hspM2qF3DM9+Boctva2W7g4cv/JHW
XiAlECLYGKX6Pka64M5Oncuej77xtNlpiIXH2Ab96IsXY85Id77o2FzKgyc7b6BDKlKvrnyUs+Q9
r1PuyFt0KILaKCgVbHj+Sxa7HTDW8JHzwbopK2183vw8BhYInRipMQ21UwrR/HoVYq3mE90Za0sq
dXYmcRO36mkh/K/hb7kc8Tb5yvBbXydAKpQOruZKbWFFupXyPkrClrqq5zlcC+ZfR6JpWp/TzHzI
dVJHkUTHN99OdpKiXaHX3oFtaGCz2XLJVO4A8nq3zWFcNBZdb6W/yUs9k2sd1klZTzkJneWuU9Og
mlksQhAO7XSydJOtYgIptS8yfiSFuoqmrKJ1epwWoQaq9YfQIE3IuH+pBJHtf8g0qQ0dQojcdhh1
nhU4fQrYh3cbmzfIg5g9oEw5sb2nzHud25mmu7yKjzglcLTqvI2/5rQ7pQdWyvxLklADCw0npz+S
MVckeATuwopWQexbNmsxkptnMJnKKMMII69R/3R7DZ3gmIUhzjTE2/Qa5J6OeJ/+dGolsX7MREB8
JdLqb0xGuHbYgExwDuewd7fopyw3c+TO6+lrK34zeDs7QS9/inNZJeArRAriIrJCEv7VN47QWpTH
Pq6TTYsQc3JqsruKgwgGLtOZS/Q/ZAv03CidnNj6H+rFBnlK+AJXYlariAezR0qLdrfsWb8yONaf
wUXEimAaaSPiNAbnC2giO8yf6hZA8gxUWBZyp2sZvJRhSBeAJftwlKkhG8U4+eqXc1isH+1xHjW5
zinkd8GoZ+DNHMMdQw7Duy+MCUHuFwny3ZW6CCd7SBt2kczmtbk5ZcRIzu+rozzoG+6VxO3DjARI
ofNoyIYMEVFE3aIr0aT2hv3+g59H5veq6lpKfnuviaIZ7eN1fA3M5wYLNzOEvdWlsW/Rnk8aP+f/
4YBEmUL7VdxYJzHUtJ5dT2/m8qExkfC6PTwf9PL0G1yfNDepm5+b7vyuGnUhuDtqp3vK2ea/uPxb
K0TDAyUuGHDHcsYGqYFd72w6QLgfvdGfqOnBAXWwz0OBoYcpw00qH4Prn7nHHl0u+O9HVxq++SwP
AESWKqZjRZEucmmQwEhGwCusE9tqazX7J/KlVLZDABeXajD2DaKeZYulhOb0g8lIpBhm5yRHLWLJ
umosMZGpkUCs/6P05wBAeS4/1lwBoPQiS24O68+T45Me8tCor2PmnUst1cl742n3IwCNxW1Br4lv
USo+/OgUOk2eQNdtoPoNwM44svJVsgO8dDjpyDJHOkmjev9sLNsAIb0IK49QLmV2OZo4XoA+WMll
EJz582G672anTPlXYpBgOaxLcLS/h1Ow5W0T0PQ0nUMzGnzvyXxuJM2vNhoWFzYjAhvF9ItowajM
pofoLzWf0DU2SvtQywnzlxqwBw21SmBcu4JkBM7kuRoEhlmkP0gKgxxECh+oE6sB2DtwLAOw1SxK
54IzvghSNRq+Hmwdd1MeRO80c2juandAPbir8afFUjTmhK6SU+Y5CVcPePG11ZDlP1PAS2P3dnas
xRu55amCoZyb9XgA5SFDMJMjxfzq+B8VoAN96kKmwn75g9ooWKuOYPZ9tuW4UVdf+tnI3Qi8wOXZ
qH3euWKieowNHX1ADGU5ERp6vu+c27Jz7XxiLprZIa1okgWW9to4CHuyyBdcYDQcUrilYikEKDOp
18P0nPAI9kEVNB9UhUQvu2uMAxMOS3oT7QqnevmDzUEa7t9HCJ0MT5bhfj4LfJYzsERHfKt/Hyp7
ppB38kCnB0NElmyc/YnUWTNKAARifXjvoBliSHQAAHVg4UgY+YHAj7kY5gwK5FyRnD91AZvnLe/S
fRMGPFdmO4dWoCLpO6e7fHXLpl2XszIq1rSgWkIrVdGPZzLqI2eEkXCSfx3RONYpGZK7ZFik19Lp
/QCytRAXhKh2vZqAkbNRVXzzMv5o/upChouCzZbpkGBWC58+1N4ImdNB7Zmzuf8Sop+jSEkKnsIK
aPXpTf5v1GVO7VPSNXJzFNczjRONS8XEc+3yVO1Xz2cYcHyxwn4Iq/zg0rSNzqoOsd3TbM9C+AvY
63hzuDft2Hl/LnF5POyiffOGTbuFX62LGezFQA6VsAoe1j7f0smRhZ30CkvMbh32O6AqLFCCafVl
shCzu5PNIuHpPrBQW7p4OnAIdKRd50d6bIhv4QNyNSEJIIKL1FzxTWJ3Q3pV9Kb2uMaKqNT+PsUG
J04ybPs/JP0zWQ7dNKdJ60WhpSpIzVhIqY1YkPyEkGi8EB6S0pxJWlV3c6BrZ0JeW0JQD/nSIQKR
m+iXQ5i2hAFyF1QXa6x5RHyip7X13ZyFyOjH5+xaWzUb9PMjfqNXFs9q5idQ4cuKVfQ89gUTIvLt
8rL68SXmcdfxqXt4ZC6RKUNzHnfALOLVBl/z6F/VQJ9rCG+28S9Ja1B/JAzSQxIBr269fIRRvtpt
cndRvJlzeDvUROG3Nx2qFrbi5efUi4i6lnLY5c+SpfCxwo3NkZ/8neMB2CcIixGRN8bysIf8XvOw
tBQFgXE2vUPyyVEYvAEEsmdgsCGCeq2zgEuP5G+yRbDnuwq2BffdeVondMQs+8RFB//TqqdBXFPK
I6j/TfNfcwgz9AiFpKyJvE2DCpwGwRgW2dqfHv7emFJ1qTDz/Sosi1gEFcHgW/Nbp6raA6Sy8u4p
8Q3xZ/SDPR42GTzOOsNJDzdkGHOU8CbYM3Ly8WQK2uZsscUzhadmoy/owBL/E8pxpaQN7gZiVzF4
BdWd8OvxwBCq7NpjlUrV98cHUKI4tDxAOt3dPv97hrDf4eyyVZesc0CXtl9vo0ctQvths9wepuA2
bGpB7C+brlBZptQ5IBnBVcBxYBNAsn1L6uzc2CzWaXcD5SyLdGPsAqTq5bHr6DzEU1AwuELXueZb
U7Yz306NqFgg/od8mplcQKg7I5NFLJ+TotcVeQMv1BMfZa63Qfb/IMIjFRFzuYkE96u/4kNME9Bw
Pf95avrUHxCl/liQHWElvNqyGuIM//aJbZpMd5iORq6S/8lkxNS1sdBS7W0ShbFJjnCRagHqA2hi
m05Ala/PsOVcx3HdHHb73Bc5m2GUqcTT89iKPAuKS22KtrwNZ6ESwDNx+jEUUXEwWyvjs0PCl+mU
CJluYrJx71zAjONefBf/TqsjHIOEY161KDktDxjJgnDlEbXONQWqRa4WsoTXX4okFoDZIPwkX/O4
RZqcypHkkxWfwxPouHvS9B7KSsGPtO/zTvah2zJ/xzuY+lhclQlTi2sLUlpGjXeuHpLNPJSap/+P
IR8O0N/rAnzq1AQHxU+o3HCmgRiI0k8EN10ejwOQKQqe8poKR43BULEMQfFQtrD+sgP5i27onwzb
sQu88S7R/L24GqG6kWn2a4QKc1FFfZDN/JbDZY8eyiqgV59mwJUa5JYItF1tXC9oOzu3g7LJNi7I
9UBdaSfQjMd/tFRnb5BRMkIXxv57mKqibdoTSyFUxveprDak1wzxyeYktWGj4PYmcS6sH7c3g+wO
lkLZt64rRBh5i6KQEQ5jL3CzcntcKVHofbO88m9sdCWcMTAl6vUYrj9Upx8aLOXNQH6/JN/A38Mt
VIBI7Wowb6DLe8H4r23Zon5Nt25jxFTfBwGM93w3IX1+Nv/FaSIkkul/6sxUW7lOGkOi95AXc/I/
GcAFSmc9dRfiMGY+WNhV0+5F8b/JmauO4uvA1vHHVmeigU0by/pVfUUnCBLNmbHXUVBRN3g3PzwM
HWkuwqT6qgoKjfam+c7eAtkGfb8ou+QLTk0DNjMqsf3gZ6zMQHlrTesOOFVT8+BC57iBZ6+PWyIP
sC7QFkY0nZQNhhNQWuv7agKVnTLPi9lU1F0BL7FTHcGUzmXFRRKDrYzk3M+IAduZ+834b3b+YkCH
AqAWSSQM6Eo3Oy0FkguOnGyqDdHzouaPbHprqYUmJ7JRdqNMAjli7DTzI7vZV8go//6hdbfV/BEB
Kv3SfuctZR7RaoP7dDJLcJGnzgbVRtjRAfABLSAIp0Ig58L23gV8PcgZGz1N5WrOzEnEN8V1+j19
VyXD8z7LNKxE0T4xii5xkECi+/KnlFbZyDnucIAfOToMYHXlStM1uxkwxpw9/9TEHXWh8qzR92Af
GzC70Lqmxu1ts6wda4Wmw7te9dx8xaimFQZEBeB8QhOEYgR78ThewCLuOEXwtNFKhxx8aPo35HcB
NEZ2ExxWPWNSalHvI/xMotEtYM8+ppORO9hKsqRuWGMDpxwNL7yLdvtpq6ZpqH3+auzENuEruq+l
tNMM+bn+nK2vmFl7WOqfmIqKNvstqQItlxF9lt/r1t7lTIP5YPrGMr3wYFiRgXJ8tHOHu6gHqKBA
yeUC7b8qS9xhAvlEJPtiOU7yUD/8XaG0cRptgGL6Vo4fNXN/5HrJhSPPD+CcI2M1DWLwmVWy9wQb
74MTXSJJ262P6xs66NDMQV4R8xjO3timAIT4P3YoW3AVD5Jmz12bePULtcvSMZ8UiYNKbx70mF+I
p/b3HEI385hZ8Xnx+RS2y+VhIiev2rcIrMSTxtpIlBKGPlSXwMJBHgWzrPFRs5uyhNEeuVWBWCNx
xg2ld2qz9a77W+Nbqv0quBDIhdjVsQs/9BmsoyzSY6rwn3g8xfjjL40BpPmkYPBZXelxgs8L/S9/
wrgJVg092n+fERKsWoEX6nq7hLPwJQUcSW9sI0JfNNGn3fQGggYEEK31fxwn9y1w6phFNBPtyEf+
K1KS9s4jsBno34M+IXPFOQcReM/ZglciA3KDbYmcWY8aRGrfqUchK10uu2pC4vuNz0Tgixadh3DT
FusVEK1oXFi7Bh6l/xh9NgY6skPoRACx9QqH7FUr7MIua748pElOxmyHET5f4ZLRYxof4y++tAa1
LUxCrhTgeT26f/S5WZCwvsuz1ex9tLUlXC8hs4hRl6Zqps4v9y82W0fE3ScgDMg/Ifac4kNwviVS
Tdn2Nt+8UHsgpi7e28mCffUbrvXzr0XRYLs1+ULjNoQTr2BrD6HkSgFyRWaIhZYltdLRJYZ4u7BO
uq8tNaWUk+kBtv+ggxVwSvA7S54c0m+/4IUkQoHmrVwLVoky2GAuf4hruA5EJUoED5iO6/CWYC4Z
nFwch1jvxE3osjinrKttwffzB4k4UEaB/x0JldxBEz74JOnsfKaL3Guv9wP32jsdJMZJYgCF/wCm
9Ulbw/em8xT7vBrPcTKB2LNLYdsLgI/zNumqvalpdzicJtuHMWS0WleZ19srukWvRPcMj/9Uz8MR
s2T33ia3+ELYdVNN0c65hSBWK7Mq1ICUJaJg5H+nIJo3/9Ynd0/VOQID5Q0uRzWPiy8fJTxDQbX4
OUyO4DxWJLpax3AP7rGUO+u0zWWPaTxKyVqRyyfS3MWU1W32rrwaCfKhFOOwxL3TwLF1oGFNt0ke
XUNNw4Lj4UEbPbWlNEA75IslCnW+NE1LBXXwdv+s9Z8lSQW2fLiDKCovQsY/pFkU6H8pgITKSKHo
VLnLrE6YRshejPDRRWHKswJEZ2Xu582fOoNG0r99AE0hS16PM/26ptR/vMeOeic53VqfWOgXk49X
ilUUSMhmcaymn1V2a9fhO5swQbBeypBD8DfgfCnrJsh7+OZwivXjepefTYOoci5UU2m+M7cJGQBT
oRxQoQ//kLgBzuxjwzbnoR9PDX5naEcE7BY4G5ouULUKWQYs3agcKtPR6G6y4XDNo4zOgKrSYi95
dGF2xii3YXOKQmFwbYZY1qHLN0430f6E3Ks/VPwoBvqWnX8/duC3mhPH0tXT4rh90lfb9BbbAU51
Ke+s8L6fomp8pkH7deQa92z3P9Vl9jRAyTD8XGre3vvsl09KbNNiSfdeIIaQx1ctz5uE36OtQ9lo
b3Bz67ObsNIQtFH5Suc4jStNaEVFAh0V2wfMEFTV54eurHIvSlCmi8NcMe7bCpJhnePxtafAOlbb
9YFm4yOCCUvUvsmfgHJj6+Hvjy21Bs4/T6BLsv7W68fUYZ5O+Zov4fGSZCVUh3tLI6Z9hY7bTbUX
hSlmHPJ/yFJFXTbsXATC6YmZQ+2+JuDLtITMt8NXNQKO/45n6t9+3+sbPf6Dtw315VV1zt/aH7IG
RqsnvCeEWMXCc0QWwQuI0GMd1Ww6jl+Utbka1+afLMwRGpmUO22gD+jYTYrQkwZuYpuwAvSZInl8
+dFswfF7mIqsS2BsxU69HnytmQqojZvordAEZ4FDXCyJZad+8PLkseiCD3PThUkk2faTy7R3GObg
GcF8BXeE9wymdCx0sHqTFy6M5ujEUhajwzLeFzmjGZ7I0XqLFeIqjH2/ZCLR6SF/nZ0j9S+eUxgL
b/6uFL5oINxZ6uU09XUFMN43bt6yYhFO/s/o5fjgZL6MPGzs1roGzmSi560S0W5pbAGtZgQ2dybU
BEh7Z7qQAHQEOfeuVstID69gIv9VMyhVpJRH1PX9LJ16vvDcDxv2icqhLhfPwSVoUKzjlVSyoYe7
UPREl6jBn+fAuwyuIJ9uHAIyHq7bCmp0qnCVC9nQy+oE2bGXLMMbwAaD6U2D/xgzotGW6pgmJIMw
u5DQ6YsbbthQKxbzaAZUpAXmf0u00Ifb/eZwNUxEfSq5iHS/uA36B3cI1ae/Fx+9dWcRz8bBqj9B
ds4+7EWH9AJ2vKNJVFW/sPg2Hg10F/WBxvaHOYEZhn4gMwCA5Q+1Q6xs8Crsc4R6oOT05X7jDIli
IuMepJKM1Zo8iIwjH6cVXtnwDA+gpR5CV1ScIEtPzkS1tTEnCSG6OhttJk0PxxnVq9f2mQOw9IAH
+EuZ+CpDiXGrWJh4J+C8bLjnubSvEp/WzTLPXBlThejP8igb2FeyNNfk73lbZSM0I5JbsAHXtc+c
QaeSO7gy15zF/TNls5psn8WJh5AbSwbXjTGeYSBxO/oRNWKwK2C0+mVsMDKz9vBsTIxMCE9iM9PT
T1BgYbJkrBIuiXLIbzEnOYLrcp9cYsaNlOnbPCpcpmJuGe+E2QgAZiIBbldMaqTtDq5/BrXeV0cF
kfmZYVLp9q/uyoe7MYMC1FWz5ASCcCfz8qd8SQUC9LQ+yXmd27E9TRCujVew2ONXWG6YlYld+LPX
VbahZ794DxHmjZyCGzlPcqcEYkdkmmVNzZqsQrdPJJYfMuZqb1VlVG7RZmTXK52HDX/WLeA+yYWE
clFj3VPTjHAdL8VTaQaNhaYswNOYcvMpXhbpwTGMmfpIhj1b2irzC3gf795sJiUBsdD6bMF3JDZ8
g84HVhQaG6MdC8jSyzG6GK9bJfpQAsdY6CYrhMQyMmUVWGvgEjZlOM3Pz7Q6cYLcTzZf3OluVnxT
URAK53fEZ0tUu8vzk8rkuyIvor0fGAkvrnXxe/vRBAFS5WfgQNFQE4No9KI/w3Mk7S7CxMJhnTpB
ur5f8sTfVbYboZeFnVjDENSjSTM5LtO6XBuFb2zF+424pk0sZh2U7RwvpVGbH1rmZTLSuv5v1miK
xkglfn8hQ8tz7ljj+XejrGsrNHxOkwl8k0pLVoETOS1qH4iN8BfvJMexhBBBlLPiPeb2JA/xKzmC
IqqRKERlFtMT55eC3RcOyZpe3alQ4Yj8kvZVtTFtQaRZfcGBV0zVqtI0CueTFhDMatODvq6Lm1kx
UD294vMZ6EO0ULLMxPsPqsHWCxP0QhZaRqjMPhPyrOLgfA5FFEjtPnT92Sh35rbgrp+lAoamDPQU
uaJTJ6tlAEKxQQFgyfW1dqSOuP+VezikhJoAOI5jmpKkE36XqVyq/AT8yOiKjCvUxMk3wmULH2nR
gpMUF325kl767a9ee9XjkJrQ/1lIigBL+dWQARul0mcSXBR2xzirjqf4dyqUj0Mu81kyNgsXSjQH
kV82P5DhNu4N77EoWfaIu/aouI8U7ReQCJUZuuAVVGI0n5XMzAz6aNjKkcuYyNp2yGRUH3AQphkz
dtxQw1m+zKN+Z9ucbW6VZxjbESKdgUtuRtpWDdXqvML4YjcITEBLF0deWVdWgQyEoNGZCjL1IWVE
f0qyZdr5YMrKqOGixG6XpHwKM4ZJC5vOunnq0fO9qc2ZsZZWlaSCSzJ9YrMIKtwQo3PaoxgSQNXD
uG36S/rUI2tID2RqcsQ5WNESZFr/WLtCJiPU8EzZgiRPljStshpJ9L+YyI5m+xQZPF8ychlh4efq
lKsUWrnIzVP2pztJEJm5weOO+BWqO6Ll2Piz1zKMtJ8xltf50GeDWJzmaHl7+BU0L2OFwOnlZAs8
aayIIaN6dq/sic6dd4eM+VjOgpXMM41v8Girsv3FA0QeRmsgmeWLeCv8rt7qFrN2TsbsoAsrTFxk
6+wyqGxpHMvi9du6Q5JY22cj6vLm1a79Kpe1jaDMlacqX6RPByYEznieiiz9q/KehEQdNZVXWr/u
c/rnJ60uM9KPWF8vXWirz0WoGyArfH2CWr031i/USFDgm6fbhLqlC9jBAr+mltFxNE+5Tp/LOows
fcDyFwfvnf4ppx0Ekkbd1oolehzRtRNb+juGPCO2UFvmEqTubE2vt8FKNtkX1Ug92vDaM4w3e74N
ohDTrAHMF9QbqnTTAZz7tLRNxVUUge7/nFz7Wkf87AW504Hkr4fvhG8WEbEaOr23CQc6wGsrfhnf
oiHWBFd6ofLnV4gCnEvPWLEoddOM2Tzy8QI19qWG2IR9oXx34EaG2bogChqTQAZNFy9POS5BEFUi
Gt5WiCfhUKlIN+qj6eFS1hxajQgGA4bEjOzG3u2bJdIDh0Rez6DgrsgCpoBtyfw+pUY8DMpERYkv
ytqjPW4WY+EIkptMzHxemTTMvfTv9NMsVUM4i8NCtkZUzFAHm12nwypQl5Wo/Ch+RBuA6kIFAqbK
TYAlK1962Ql5zgcLK8eqMrZt6xckHge+ObtN8qY4/gmI4Ydk8LFZW5aBjqsw4jTHajQ0OQV7QhW+
NpdGBjcsrOF75XTY9OZJmqJx6ObmgymP7ui7AMMM3vUafHRH00s8ANO4TUYxuuPJdH26XvifX5gh
gwAyZuw8wNaU2vQ+SjiEeXmFDMOAqUx/ciSReWpgO57ym+LXXMSqV46AUd8TZI+Xqzt/Y4NzLzph
eL44NEpCvTNiM6mMZC1rlHHfwQC2TgdtIql/+oCWicgMvpRNyxMwsBBHhRXHQR/wEbmLw9Z/8+fj
O485Af2BLB94O7gHNN/suOoRbin+HAAEqHBBmrHk1OqEGsMhKjgF0rYZYvgKuv1xmK4PxZ5dFDfN
vX+9rVtyAXDY+ZHtrxWtwSvaU1l/p1wTgQqEmymRBDPyv4EZw/QbD0xttwUR/xJMXdTOVFWYDYiR
bjyU+HHnlrRFj5oNT901VSzJr+CJXxYRqsgIXlJeBEKm9IK34O6mVjQDMWsNKX/KQhiTfcgq+7ft
wqviyySGpvpcpalf4mbGEQULXZP0WKzpDh2g1kFWWsjmlK7FDraFONVTKB0LfdOwUbxzPyViOZiu
dUSOS1JrTveUMBN5s9BEirxjvdCO+oE4jHXoWIW9VpX+UUCKA2mTQGoqj7GoDT+pDtyB0m73x206
VSHQDmuev8DXyjvIIwi/UBOhSiY9RGmzZprpAR3vbQ/ouhzl3ngG8Tdjp2umV1D01z4REw22Eas1
G9he8yGLuVnEfJuvQ+sRpcnRjQxXS1viRzzgRiANC7uDHj67L+4CrQoCFi/eZAXUStQgjNIfBZ8w
IPpEoI7UvGFThTt1D5lCRyCt14Jlmzn6C5+TBRBfVCXSJSl/6o1/f45nMB4mGQHknjq5k5FIWz6h
C2KfRFz4GnlH5v4Vf71O1spfLK4M9JKRITPwnUvdpVOjeaRkrCN8EIerlA4/piNVfIwBSa9oS4Be
A1xVmVcWbNqSU3svP1xVVgMKFRW8k2MWMRUljE/O6ye2SgDKjTm2VCBqUhF+oBf9TxADVoCWrBJX
F/lB+HIx9of7AjfEbh26i4rpq9gZb76Lb1sMbeDT6XB8qRjKWV/5vBg7q9pneZ+h2h1tInbu3tx8
h3Mp0gI/grG/eOXsYCnUi34jny+ypLDIvCqmMIcc7bsfJwBgIADkudeSRdpQ7044XBSSfWz2QdC/
BN5FJbCDUnjV/UKyF3c4TXaV9gDP70w971KOE/TU7UUojBn7faPDmNkK/rDZSKV8TH7rM80nZXrB
CUt3Gcf3PxMbv8phSA/1YwSzSmuMa5B+qcTtJKi+KIBUeYjr1/Vb6RaeZFBeqYn83GCbfS4WvPfS
Itb7gNqxvqMGor5Pq55HKqe7uWkNaSsfBkWw6jrYVL00oevWMV2Ey3rIIEbOnhv4GzWJ7aMf4vOE
VroQNXSHQccsbkGJsM55KTqxzzGwWxK8Jn6cXu3y5SJN4BjY3VHYcXxtWLQHsedWTwMRTRCkPllg
N/J/hLIqjVKLPQ1aY9LwcZp3nypd4PvUoIHok4v/hUbaRknf55NZYCxzVvLRimBOvT7zKs9u2qmz
ccR0SacjRFmIOEuKyGRyQ9TvtkjbW5Fs565Uw8vHBQFTAyHNoLpT107Vn/djfcP0sSyvsHrZstas
SLyp0RVa6Sp5/5RNoV9im0K5u2R8GQsNw5I6B9nmC7XgZ0+oJFViEv59PmczhCt1iij1/5reHpgE
7dfxptoUpvnXNFuVQxpyb8P4psVWzb06xZlT4ysT0oVUXJzFdVMhvVvdzDzCtrFgoL8fBcuochM0
L+L0zrYxkVkyT0h7BlWF9aYQ/xWn8aIB50cgFpDFIrOb9K/lJlTb0Nj1DyVmh26Y3wOPO0JybR2g
U+BA9Kq8u5I1VqUE7dJEDSkk3N3eNkUVQPH544n1FYL6Oh9cHcOf1lhmRQ3/bTyXJc+ksHOggdMI
0yxr5qF7gXVkXJZ1k4T7/9KSCUWHlJplXogrKciU9kiPTSpcOqVCaJD6tFVPHFervvcKqkCQ43n3
vAKWOTxXdQXQvgGKZBr9ba+vk+17yLV4G196WT8zQMGo+yogrtpGa/1REPF5/Z4vvFxEd09FvHHn
40DBzKNy7sx2QMMmsMIQcQLAvFdnlkhd6FH0Sj13fXRkr+7mXt1x/SCTCw6E04dfs0o2qe42M2yV
cKvh7SOPyroDz2mlGPyT8gksFKYTG0kbdnSHCrl0/xZdqQwqCP8As9nMstgYgluiv+YIldq98atv
tl/UaMLqvEK/Kzco4Qo1NLmRqRd2oFprvuHZxWQRNALyyOWV9sxP2S69gqfwJ7rEUdIw6v6NUfNS
P2QU38UYi9Ne7QeYzqJXsuQjciI0UMNrw0t6hQ2qxwWRIJk6Alm/3wxNxkfJytIAd6O5UPfARiuc
U+pREADCmt9tJFEofJga2nkYKlWVwlzlUNMrQ5qJEWGXYbXJYXjj64Ri2dQ+ifOAOXvyzwFxqhCL
rR0lE3lL/rqsfjqMPwR6biNCpO9XKPXw0ppYBSnbW05ql/iMvNUrhiY19/WjuiYt4uVjRGHZnkSo
4mEd50uMdijyDE8e7MscZz1bC216DnbaDib5c6NjabU+ZsaI7POBoAjrE6J5e0zH06t8zKCdhehn
cJKxgW9Q5y4UxGeKTlFRF7H48LkavIBJq3NhDWE9/7gk2tbK/XWX7V2MKgc3nOtKNxZ7nRr11UPa
fPGTIualYaQpmqDUowJGEBtdTYsPs/Xt4r0XkQruO/ba26FT9dbgYRuYGHbfMC7futdCw4u44xjH
3JvCVsZYdapDJU0V2c6y7s2pWxO4EKN7olqGhkyC8bRCjANsYOZZnmo6FoeCKo6Obls5Aj0z18np
pB8a68qZBHrcl4ycuhriE83adWDOsjcd43SBrJc07MKIsjOtlp8ht+Y8TvSBJQO0/yjnuvO406qi
M+NJKRanKEsGv+vKo8OWV4BKFLXv8SeDPE/0eaDuLDNNNv1iFLglix4YbNh779NElgKXQEGnjpuJ
JNVzhTiyfglrhUHPmCNlUOfnA5Wf3x1eTbwHxdBuT2FBL/GBXJ7Y/W+CtzvPy35L3/b4tPy2jomY
4Z7NsDxB2BzEgLG3bx89skPn2eGXpg4feQpxTlMWRixEhelem6KOBxhPYLds9Kx0TyQpVbmPKlO2
QDBcS77UoEvmoe8Dhxkpsbp15jApbTC1YYI5X9tLU6u+m/rnbMKM1OncP8YazASsp29Xq/Ph/mFX
N7+VD0QrBHMfKgmpV6Oe7AI4Dc3vPNkFsBE4fU1vR8g0Ewm0haWv90cgQB543jB3QffaIrstdzwn
YPANZYA9waR255PNItTCU3Y7XPQ287Fd34g4ofbEJzuk8fKiTHtv37XE1ZGNnfXn/Q3uuQeV9DWg
IvQ3vT9KVLnt+QX0CiAfLHFA2VSsKJE19FM2Os9yTLRs6bUqVTVyN7WK55GGjGRjTcPLmjjgNrwo
eZRSLPl7p5JFEEdrt3HtxOxQh/WNH98UeMIXgFxoHd+LBMWCWtwGoNpjSEqVXkvXILtoLx0oAENB
cchhXEQdKoxl2ZuitQcCm99wgR7Qct9hvLalttOHpx2fyuycYMfpNLHKkJvCMyK1gZ5t29qrKZWo
wRI48LnVs/540XLgRvIAXjVi/uLnLXa5KLI59a4phTjKVSHUYKYeyHHxoEXqD+lLK5bVeKpoqAJB
4x2cSJC/QSAsbAbYTUwMuwT8ncexFc9i0XSMVtE2ZVQYc576rUr4ztodspNn7Y2uItPBO0RVozsL
qsMbcSF0y7Z26MCMsQ8BSj/WKNszv6DOEP5PAli4IyZwTaoqGYH2hR/n6Bp9jpj7wvlXDQZ5ccfn
TsbjClJI/D8Q0LYgFtOSTUT3hRjbGLioBvmRLnrAAT/zIdTkd+L84fr/04nkVV9Ec8BMyh761sg9
NIIDZ7pkJsptl+Zp9yQVp+6U/oWIBB3vuB4C0GzhkXpkmvlllHuup8dQmdM7w6m3rWnjbjhhk5LK
vxPSW/+2AvBbkCgC0iHpkV3E8g5mgjg+964PXLtPzVmJStEPLmzfMyOV5ci+FEEV7JtjBB+5Gfbi
sw/43BmcfdDnXwcagECb9/23PeDmI3mP/WGL/uIuLzguKKHTLcYMx69+5PTehQJwuBfnaLXvE7NT
c4+zxhInTp+30qzWMS9wUiwvSCTHIMIM3JbbzkN7bR6x2pCCzJdQLTToYto2aDcrXfEe5A/UcEaX
jGaC6lUWgBQeWEfOKqWMS1COsqDyr1jlDVzxOfSAKdAbGT7qJ7QxEjqCjW9IVIIKdhoWkP4CO1qk
BtygWP3vC2wWuGVGZnnwl/aY3mh4072/QOOPGLvSqQg5W3DDEN0PUaImbfhEm5HE6jdG6bnW9Xxw
G8MeM2Kt0ijRWSSCj18QomNTu+VqabfqT7QpgWATGJwQQ8R81wNMvCYneTZgw6MbDbwdYFGWV8xk
LCge5B/RxnhPaU/CqxPinS78Sk7WWMaHuc74sMkf/rd+HNKRyOIrb1R901t6EWDgKAUtzGi+WVtP
NiFiq0you0cegYolrZ935ZmxNasE7tlMbf+r7mY0Pz0orW4ywTixx+v/LmwhcOJhYvVeAuf5hWB8
PLkeo7OtAxlpy8N2LBhrigk0gVqi7kAOl1HRENAZyjJ6IIRYYgJ6UusFEuM1eNNuXH6DjC16Bmf+
EspVCowEnmZM0JKMJDPEeWbXIilEEgoVIL0SsqDN9GkoDcDnK3RFCU9Pi9nLwBJiy3Se2UCNRpz0
ZfzpPaZ/2aFOg7uPbhYQvI4tYCK6xZx5NZS+cgujT1qUibYX87RQXNqt/KUbfbbTaew1P+b6YcGp
Y3Lq6VEjdSEPq8Tfxbe+mkQerbNfJ154AeYC88amEMk2grqhPBw7XSDa8tlCp7C2ei2XHeom9Yih
TUC6B+nW0qlBrr1s2wlHuVoH6mecP0DZqlAvl9FVgfwatZbpQ9KkoZ4cnsKKP+h2+pOoi1yuGQwi
H/f6diL2wJxHMKfXudqpi0chOWXnsWTvcyONn2I4y7ujXc+zN3yoH1RDShNhKAlub6OEXxlbFRPS
S3pjStCK6k5exvOaiGioqUIl42QrnCjLkzwdYbQ1t0kauQVgKtRtqxsumw06G/PO6dvrPFi5FhXi
kXcLe9F3jTLb3MLRShSvx/GaLWOc/bHhiGiJ1N1Jt/UP7CZ8u7QhNwFXhvyGOZZtYUyXuyP0nV3e
VMejV72/uYeEd5gKJVY9a4qKv9eLQUo+j1dXUuOKlapWm628AbFBfjgRmFk5utNrDmY09Y91/U0P
aU0pOk9FP6B/dOwYrmO+UqkrP4pCfgJ81TKcO5BZrEpfSLWYuPckO9VRkFOPKYvuQsJ7PWHbcya9
Q2tJlrQ/4MgPsNeV3jfiY3aGcn2onWkscvifmvYKXD+99BY4PMRkeqAuy2NkrVxjCRLWuSIQSPnW
eXIPO1Z+6TXfzL5k+jziy4K5eW3YLanPOBWwHBLfI9BXZS7iAmktmWwyDXyEqtceRoh4StQ8xdwj
YfZg/3NLIdWB/HlIL0GVnVhiXuIBsLCFC0ZjZ/79+kvSoRZGB/olIH0ii6CAG62AuMZjSWgJzFRl
sqRrLnxcHYvA9Cr554MC4Qmn3KI6jqT0V19Cs/StT3ET1ywNXuVx8RNXwLuvr76rtooFTLaSrqWo
qlOLAMmLzWGskJECY65RvPRJzjnlstX6SPliC3tOawrXiFSAVh6d6ABcQblOma/NmqrlpOF6dOGS
3eT53C0oJ5SH0nRK7YF+L4xTmE6ghiwkqFSHZ0n+T/OrhMJn2m102ASTCs5mc2loSeSv4AwjVU6U
Nys1sTSIzPEoLTVYmcRxy4DVF27YZbCsXcIpauEuZHrmiuxhdQ3pBZ6v2kjoklsqLhak9f7nnpMO
kc6h1NaSx0XCIJ6t+Mc3SzDZBRqzulESG/UtXP8ZJHW3S/c7f7B8xXXTr9r35bYqomRnskDlPhjh
GXaTjXpABdSrUsMeYO1S4zNz4t/TJZVrU9Vh+HKgkfY9hbCSZ8yarXVBWMlLvBG1vsCCKpSTxlvE
gwTdutM3vwRNKnhtXLf7mdDUcufX3gDeKBT1RGfziGkfs4K8OGIHLJ1ZbxIIVBBA8uFIQP98tl8E
mz/KO2R4cFmfDSus5YGVY2ZvMVUTi6lPfplDYPOnDML1T9hYy7LEqYZuKZ8zLVVZcuVlTaxyfKmw
JkYnxYTPRulfo/vSImh/CaITSnm4sAR9uHqQk2Y7Kqj8aAa4L2zpt2DdKuvJeM2NFkDLreUptaAP
GAtbVpHBAkPPt4vF+9rQxyAdfFyK8ifmcSfwnkMvx3XZLzE1MQRGrkce0O7s+mqPDuA1YiN43iiy
/pPwmk02YKu10NBsN07neJbP0tJuAMlp79Ht78n+9plI9ecodYbUwelR/oYbE1UMLgz/yG4yEuIA
/I9HGgVBceumRUBBICuOhSJIC0GNi4UR9vcHIlKSwLBsbA7v9QxBtpx3/zmQsV9VYg0I9xafjUoC
1FO4gPZFo2qAqtSC/Iu0UOgaoYCmG4pTHRcWFIMIqgOK+VK48HjRFmslwS74JfnZ/XVqo905CNwD
KG5UrXgi8Ubx7/vUzETJ3i56lq9NCSF1n4PJvAhWlAGy2TDHM7s/6kGUhHskJ95geqsa4Ml7oPpd
YluPdRLf97IZiduCS3GB/eGa1YG5HucHch+NTj/rJAhmMGVFKZirXXEQ1rVtd79Bbpge9JJNB1VH
62s6ifT8fqcE5Uhk0rvv4aK5nNVYjsYP3yDyYzs/XeP64aNCzbqZbzDLXkhC7w+G16P56izo33fB
zCIdIS5m705v3BcswXcFvn5HQEN9rBt/inV5kShpeoVBuGamcadlQ8SUbKcLF+6zGu2V2S5M10fd
f/6sw2pLOMP/ZU4W5LSRG0cowyOKE1i4+cEcRjc5e7d5K+wEkaSC8LFznXvKSPE/WX9E4dkjaT0t
OF2VlRbRerlR4XQ/xIAqp74bM3fn2ObzfKoghe8oakr07fHQn9CIprmkCBrlQcItl4mXblY+AI/A
gWk1dHz9W+KZ+xZnNYJyAaeJES3JkgQC5RDtUdvXcTLwDcjw2oialrGhycU8eslROtbeuOGnLrjb
7X5WkLbYE+UwgedpRc9egjWWM17tWTjnkNtVzrDbGwfrQANcCclKsPfrDCPKe/VAoToTke1SplxW
Qs11hVmT61BqaLrS5jOxcEBQj2w1NOLhq7YmfvjvnZfJhaRLJipC4EtwSL++6YdICk+5l9dtjD6Q
1Lq+3CsRCtGNyMCw7NlykBJei+tSw5hK6alFz+t84PYjYNIXERFN+JCAjrWVtfU780hhXSgdZKuv
1t4B5T+QlQ62/T9kn69BKlHOdS5QJAcxO7y1xSPoobOShJN7fkEfStvn/4NshusUw7ljKstpvjDr
v6BaDLzN7Yo9Mr1r/7vhyUxGaywlTVDN0onkced49IxW3Zkbm+RVPsSP6GYltlxagRSmOKdgSYkM
eHa11+1atnWE1FDt6DkWcuS9bH6LYge4LVIi7N0humQHyY34JR6XJfvhNPEBsULOcQ7WRsEodxeT
21wiKs1icuMQ7b+XChzIkxVsbr6BOo3pDaArAIyvtCWA6pnoopBdeRL1QeJiAMHUjmnDfcIMm7Gv
frr3w/PUyUP7ntB5UDHtympzv4mJMXdAvs2qcHtXTVX2eaQtlshD4C4YGY7mVF0JWu56PlGYcywO
kLu8pHBzvGL8XeyYrVVqKkk1oj9Ctdu8ssH3/VuifhtqEZPBm4W7cWnEPErr5rEz+Ybe4nnX7jXF
EW2q+pDMFavhtLYqTTaN0d0cU4JLxa+NZwYYKEr3hiS0uhZ4tUPZHn/QnnUq0rwKSVHkH4M5Mpbv
EknGn8LqJ9gythaB+Fd+rofTgTRU5HFAycfERUSInPrgFpHAiBx8Cd4594B10YHyWIx66rU+47H4
j2MRsscEWvT1pBNIoZIT436HTuNWHuJv63V2q/rKJ3z8fKaCv+h+WjWn5pkaWBtGcKYum1/svDcC
KJ2R09CYRccE5ja1JPfuj2+gRCqQgls0XfgSLPdNagGB/Q4Zk7Jw97LeiOvLdmXwpUPlIT7wAeNS
1AsvuN1vXG2veGMGjjmMCx+sOWGbb766vXLUIfFNmT8S4hxWXSDKm0P3rcDmNSuX8YeJJjLnzhih
atMqDSTb38uWzqqmpUgzdv1KLM1jvCWdcoDb2eIwoHJdVQfSMfgWl9zrEM7orgIBoa99Cl5pqN3V
VflQR7ApoJi6Zwhde+FErV6DkqdzM7/wcea9BdFoTlNAr90AUg5Ro5iiFPGXz5Ud52BWMkWU35Zv
kjIYsVEl7nuexJvTXpUrzCFYTZ+EgxpEbhxEcxW4gYEMzAWJAoZONCiDjUK3CInVgEUZF1duwlPy
OvybWX7M5bqa4zgVPLriW3IvWpN5kBm/sFHKcz4PBSou3Jc9DyaBT/HWDRJ+szS5C8ZFI5zWW6lI
/nIQge4B8M1WZ4AAdkFazoV+/QWPST3637a0g+SP4lTy0cGfjiUtZ/l7lPHwHJ1Gf4anWvzaXh7/
9ws2MDkwkckqtz9w0vhZEaXXxharsV1NtaBgONKT9WOKVbHcAEuoJpndQWOh7tn8SLllin0/bjFY
jSU3Taflr0Xty2tNxSMSLRMDo1cMVDPPqw1DwcSXYPyOLtN0oR4e34sMX4Y67rz3wNijkEVQpccQ
kOy5kBQJRSEEKGufLGNNBpV6plOtk5rL+0j8L4KA8yfMcdaXDgeCD+skgy16M6HNlSGbSktCnnzK
H8uZ9RlLqyvZDrfiM2hhGjtdrU5V/JsnOXUdtQGGy6TiH8liJqqSM+wbrxCLaMDQAATA3Zw36UD3
CHru1lCy2nKHF5ycXltFnEk39vh1IgqmUxjNchugoQ+euPoomSw1nKI2aWWZgo1YVBI92N2anEbs
S3CtD/8000H3hgaL0IK3Vs74YMNe81kn82DlblmoVKsY5VbN8qfUKHMfOOrc52L/I4i7vEWWhrxJ
hidgzaqHN7p30zvpNtICH8oY4wXQWhUu8nMxYMUV+JJBUvWvZtFJWTUmSD6hV5zCXh+OZvd8QmXJ
4SpGqlW+LroKUqaL12A1Qj3EMfZvFjAthRJLtQ4/2tOH48Ybp2E3zxqeT+VYIUDqNtODeCIy6JEW
KdUDJZP0/5VdcZUuMX87QYBeksWqsLuPIPUcPjl+ki+JWKsA+sUH5CPpLY/lPj8EgWvME4RZ1qYj
YAzMZQ/VO4LBwRYfw99gdZXLW6xA1IVrVwTNyvgxnSlXVQHJXRW+N/kpteh/J7Rf1PIIlPe4/GqI
cSeSl742KDBpgW+Lk5gD8Rf8IA/FYHvahtAxQTsqCyTMLyPUAj5ShNX9uM3m0uyduhHwgMivB+pg
yWjzabYWbtEhY6OeOu2UUJXr/3kDpVnzjslkC5zRoAyg1SG9uCaq3VTNC6uMOvKliH/hdvtX/gxM
UR86hSPDVa8W+h5xvrGPKc/f5aGUgbzlzNW8Umd8D12RtWrmJA2sUqsvy6k788KojRI/53yBG0Jw
PcfdkGyyJ+JYmJ7+eA0oWVDJKavR2jrNMqrSiT2xSsSezy8z1h14Hbu/fvg9dckuC4xsDMFdBdnu
Z1CN0LkE5XLRJ2X6y+KVyKc9Qr93q2sio72lx/2cfSB4ZEOPEi/+yaybT4C0GyhlBe24KBTFzxKZ
GxDoVdA0nMvP9zq+29xD4JjwR/euJeFckkfndcVzboD8BpC+DAzCxuNIF6UnMVV+vN8VWZYtYQet
XXbAaCpDTt4RXhDFpOfa+i+uQv2x8g7Q4q1e8Zn2PEmIBiqOG9IhO5W8dgUJYg7o28AfixDiEusb
7Ev2qqxiW5GsQC95wcxcB9V0MfWYhb4DFMklHdfg8RuZ+jOU16a0QTHIqEWW/o33XPt+zMuTVkQi
CuEegn8XR6m9dKFFtgr+gXgop6mDN/wVE/lr0FuYLJhFBBgKWuRueaxarLHY+He428dPDgW7ADwy
Cw6WCu0N/HaPrDmO5TaBJ1G8PiZpIt8nTn4ajUY/gks4vAhWDeJMlCIW1XaGZt0ljsmdwABYgcQ2
nCm7aWYDkxP7OWwC82dhh9bSeIRIL0864dhPyEnLvw2B4HCc2mOhjTZFtEhNuYVk0/N2K8aUEv+9
gzVWbn5yHz88VLbvZ3qxDCldKFc5HsQ95m4EccIx2cRGMtHIyPSpC6wh4w+c5J5Bzom1mAW9P/fA
f02eOHazF3tkJJYp7AnsrL0HHaWM5SAYot5sXkh1eRG0MqerJtpCjKcmlVq7PZJ/g/oJncQ3YsBf
CRenjoCNKaZ15Dfhgx1M0N7DFHEAnzqyq82VCETpxoUCD8hs6kn28Wf18RJKwz7EuTvmow7Kh7BG
W7zQIk27WL3zOOtoYVhg28NdAh0vULIZPhJfsPtM3+Tx0qj+sIq/uMpxPnNL04Dk+9kv/A10s9zO
qX2C77PJ66oNeJauTJSOyFvSrjDcvbGK4TgQw5K9KSp5Ilmstq3JbYwiLeojIVshnA5wqvdhdnJ0
/DHie08WBRXrJ0q+i35MLy6Wc49Dkyz5BKjceYcFhGIkHL4GdkDSThLId2Gmdr8q+HlLqdZVQa5Q
tSSTS9TLsvu3BaoS1j3MVQrMp1HSkVsJth765RS8LVN4E/7Y8w2u66C8f1wkuhiofX+sRYedwmBP
ViltXq37PVYoZ8/WCNQJ7lv+nMiKfG3V+bMZdsEssgGb3fhwGwXbERxdRqeq84ARok0pmcQBIPNq
fNeftut8FDyj25xTSY2cza/QJSjBb+lq3xkgIe1kI2LtMcrcoCdHXOAH29Nl3ckKyCaxFvcthp5a
XqWR3PGCg9Gvyti36yt53QCrXponpcCOfZSaibXI64glPv8P2xMJhnwsjwKKZ+0trGRAfi+4Fq/x
Om+E9ruACne+LaGi+esZyTnrAhOznjrfAkLpFfmDBFfWzGpghJ5+k0BiuY3KlIBfq+DLHzlQTzTx
etYdIFEsQ+KmyZEB21TwUIpMK3ZbjY1emezgThZ6r/NkA/1rFrTsBZZtqBGcLTZag5XTV/CkCNvy
+yYpjPER6NXokHHTIoIP1tLBFaglMon+stDTwm2m/VD1QZp507uxG3zvqiirGu3jYaL9T0elru+h
ljNbLPIFNV623nxv+qiba4ZWyYu+3gLOf3syxkETOnfHaHHfNFzZ4evtlj4IRLYwfDVb2rRPj192
KmhLa1C2kY/nO1ac+LF05IEfqjinEPFDOy5/ToTyDMUYrHUtUrCe3/fZtRIi5EKK1ONEMpT9qDIa
UjGlYwhy1MT1G5UuZtxf1D6WDVlVl/Xold5kckasKXO1HaM6hzSvqt7jajWHvAs8TyFemiqO0lMX
/az9bhEOIraEShb1HTPsm0H702ZtiZCUVaE8vWYjPRJp+YYLOT1sXppNiOUWDRzt2eNu3oJ4zSfo
P4/KEBasAp4ke3Rq3Q5j6T2ORRU1TFRg2WPorMouEooXwtCHctTJeahzbSfMKZ4EjEz3qDyv7r5s
z7vNywdZ34eH2dip3NGSkaR1vM+UNth5xQFe2gVQCVlHpzFV9uZFvTK6mxubqouv05F3CwiUVc3H
c/4iSkUIRCsvELv+ebRclaX6q/cSJ6NkAgbmOayfSyMr6zuhtZyawn7of7S6k6yhnPgiD+N4c8M5
4tFEiKwo9y/sXELAGBF5DazTp5XH4KIGauTLRn3YEjcJKdq8T7Te7yWPdoQRLhKb/64ZSwSxUcaJ
pfrkfhBm9aHsIiW6IsSP7+/3xktuhkC8rXEfOszlsQBsTkFqJiUUh0G/5AKxbYcNlwLGbm6IlZeR
U5ACyUe6QCGRpYJudJEN199wK6cRQM1Jmp0J3WsZNittS7EgacXiPs7Ywy5hbDTpxwO9S+tfTF2h
Un2aGMfjkIIz3ont275cChInnMyUxmvBV1tBCOybLDV/PhGby0dMuoppqjxgQKbje72+h6YOOwlY
9I2TT/FwMx+EozQBDaZkMCc2ksyZqjaTGpCOWzec38s9UVD+VSFEJOtQfYXxlv6O7Sl4kD26A3JM
sAWvQNB021tiWRJBVHJsWPJUEAiCHY5mDN1JNke9rs1I14Q4/YFXHI7gpk2ozFVZ5inEofO0lHaM
Pz0rngsB5yem28gGp1n1PssyeLdw6u0YDDCr4j3fT2HJp/RNOibXijxKH4ImwJ4ROWtddASRtPlU
jpQyHf3BS7cSPDcc+8LC7RRGjRr026F9+3dj6VNQHS6iuNCLS7/IrYakIVk8DfZI4evfryKWukco
aw4lJJ1+gVAXZVs4CYngnQolXwCUoXHCB3WonmSjc7M30ypPu+iKHOaHXITFPGSKa97KhE8LU0aI
U2YJA6GcIXuQMwzB4YYTghMzxxeayFo4RhGTXVIFpfRSOOG9o8OxuVyNjdFMJj9mQ2gAwbbUSYTo
jzhd0k0qsPTWQMBRPEAQH91NvThdZGlXZtxblL+dgGXRZzeHS2txiIDQgHRZb+hJdPu4G962Jaew
EURL9c3l4kcXRl+kWeSAGf9UwnuBhO4/6cYgWPxyTZ+RA8u3VwieD0nlV3ZqraJXpmQqApYNI9YY
dB/0wo18mN8aD7PJ7LfiBt9RKODeLe101aqQTMpaEE4bB7L9FfdZpQCUdznYKTclqbR/OF1YnUwG
pXlBqC4DKbGpT5gPHMjBYXHV8doYwXL9rvWbf8CLDrPgOq6qYO0kBK8IYDv6q3CWqup+wsxRSMA8
UhVWyg8fbBDPiq5eHhtaXXviinLPp94B9VQJqmW1EbLW9pbV3rx0Wq2VnXWwWY0a2dqZFRBn6L5/
uWrHgTaMnYhlmmziKTjM7guIZa+ljkrwKdP63e2D4RfgEeD7CDMunB55J00XgZ4cdSBGzhYREQ87
CIYj8tCF6i1MfLJydajIkWgu2mUMymBWWKVvraQdN+YT9Qp9JaQLT46aYrDEM1sislVcIidJ6wUU
WTKJDJV5hMVgejKkLWYtoZnlsHmvhb8tRc5Zs6K4bMbtnedwMquoTo9zumABTQnNUSpINz+R7Olv
a8tmKs9OvR8kYuzmlJL6NHZMKB202woMhkqk/10B9NSTYGmn8l17s/oOILIh0MiTnCJeKRqF7NYy
bEVsO1qJmygNyyPiAdSg+1k//csH8dV5Er4CUuebJgCFp3ufDWNXLMWS0j5xQJ4DeFFKLkARUmV8
6X186AgNYQX63Zg5bVRh5Kr+Q5euI9lyMCvfwO9PDEUlLJ2OGML0+IYQSDUT2omvueXlyZwKBTM2
R4E+6717RCfeN7M0iMx5XAh/iwKbWTg0qa9o2crrqa7aM3xl1Z+zxANrka5MH/ITtfEf7c0gzpOP
J3NIMD65NljgqFpsJ0XUdBJ/D5ialPxyDJgi/7cl+S6gd4Gw/wqiXZcgXuxxG21+C+nudlPWgyxz
QgOIONeCAcgFuqsIrjUU+5KbzoOPuNl4aq8CXPotSD5Al+/8jMzPgz1d2N7Xfkk/ZgF4GYsWhCGi
kO4ZsAPc9UFf7yCIFC7YqOis2XTn6VSFNuzUt/ngW2KygEcTFULsxx1jiZBOtZRO6ITTbXwui0IH
6MqzXcMEXTrE9FZ3cwBZyn0tx9wzK0kYmBttciJC/7dGSb9u8ffVib6xVWkNAHzPeNwOpNeZp0Mv
0NmrlL1SPuNBgeGNvnmKrHrJeEn/Th1irKw0usA1OU4+5/qhHefKX/vLVOgDzA00PnpEwnpFPWSi
qq5buNT9fe3UeQMhhTwzW8y0a+QOYMknqU+Gcoe/tctSbczw9IhQZPeA6oUbBOKcHhBZsgvpxxas
wKQ/ogoV/hfcG4kkqxc0xUdQDniGzz/hn4wxQpX15uSEP2gKRrHJglWB5ayuSW5HqnmJifXemCsy
evkDWihs90jxvYiQVBr3PbTzji7X/a/ytVMN1jqfyvOGYc12eMJMjcIBG/Y9hDKqIGRHMU6y1Eh/
NVB7oyZeInWf2l1FqsIZb4XB3Ac2OliDGaD2dSd69BOGZA/0N2GgNcykc+qQ1Wqe6m/yWYO1QePr
MMzqQMxa8UxbxcwPKdkp9Ev2sZn7vTKZE+j8KMqGFF/Ypt7k51FaqVC5pslL0ehIQdnLpIz3fTTg
i4YLqfo1/wZhohNhi5K3N+fo3v8G51CyQymompXxYRoVn6TAQHUXJ7k/43lgpmm2IRrzEtSNU6FE
ZEd0avgRrNwb/ea0g1wDMuhvV0cxEm4kxXGVr+AfdfddcN4sLNaW1aafx1ewXaH43cq6/SorGqOn
49RawH6SfUHdyTHRLdW7BjQHgCU7EH4KCVZvnofCXna7ednh6JFaX9GM5UN724vM7IjhR8FQB2Rv
Wkk368Cd0Drw+rDcuJKDfw+JpMmC6YwL7vI1DsqZ2QhVtuG+a+iWg3+90u3Hkpalpg9wcxl98x9M
WuqD9qxFLzMWGVIGsxp4FQmwHxLUN8NlOn4y2YMMAJGfeCs/9W07J8KjyKNwjEAl1ZkFTWtAFqGy
y2/QCGIQzHLrjkWkxkZ3sDjoz5lHawyTPcOqDKInOt2KurcW/t6tOI0foqikFAwPTFo8pUDOz2os
zSw1HnzP75Xi/AiGrGJioEj/+LV31SPO0qq8MMb9Bn4dcLCRhyHUktR8IY7hzRhVyo7E7UxeZh+g
i7pJXA70fxtbOWZzIUTz+0rd8Knz45oAKuBYSjYi4aS4fdzilHXl+oCvmUJmH5erUYyOETSVFYdw
io1cBUk+5DhKNArzlBHeQeRXF8TjFbKztRuR5vIDBT1eO0R0mR2n364f0lk2i3pO9FKKmzpZjFbh
bahLGuRoLz1reikNZGd+qEXy1kMO3rkP5YJF9jaULFIgcsGA58HpXII8usbhcDvPWH3aqYPZRhth
oPtXkQHYxNB/QmFF+D3qYNzJc9sSGsKTjLpAnhLiuCCZJDtL00uXST8TZWww945PJuU/486ncSPR
ZvDDV9ATZusiSeCE77CpA5mKXSWvFdPsUUmkKASOJCxBaHPWE7PmXO1bHx3d1PYVtGCK2W68q3+x
eJi1L6uu16gH5mwf/tHG7KHfhEkrCDp/3iL1UNfnRtESduIAKC0OOZ+SW209zZ1Apmruqcqb0r4n
fqxSo3GZ1GDOD2mc8O7+ZowaOgjyLaxmII0eaN9fiXcncLt8kfTDHd06+6pfqVtfDLehW/gBEXrI
+sA55v3VEx91L1/aOp9ASIXlPMayz1G/5aoeGkcLhbOeVsLNlnKxK/oKNLJXXfBuE3SZu1S4pXbC
z6J7BcHP1v2MLHDERcEawvMb2jm4MQdU9ywCy/vCUlYaq4tVKqTOhbWq+zszSf/9naOQ82dCn9HM
wENjxDknnowQZc1Q30dwIksCSE4imGmOFhM+nPdb1MoIc0LMcvxTJ8ST1HZCvmNFnkOFRm87f/2t
WSCBNwAL2m+YECfzEPNkY3SinJqmeNLT2KJBW+pgL8r+tKKXblwVM37OK9xc7ROnAyEO1lTKUw7E
29Ehee7V7ViSCESD0TbysUYTaFXU1Q7zKHnY4akRE3di6XZbfMRC2Gl7NuRUoCRbBzHvnPcnqzYA
3lwvBDmL2F3g6K9qZuj0q50SyTAS57Dv7WLBmu5W2dsdtI9h1daEBsSWosFnDTkU28T8vLDu1Osw
ASxYopaZSq8MC/4X+gT1CQarckfDFyqyx151wcAlNVeJINJbrzaGZCmQhBhTh0HaAmLahaCFj3Wl
F4DwiuqM2mi+PDSbPTa0rkehJx/EviW1cmodlG/F+M1TLrn5u6YKtoDv1ODDBLXRdB6Mni8CazFp
MzPXXWituWPCnKlEIdJmVlwncTcXpB8tIwppeQun9rktSm8Im5tJ7F02XAPH/sClVeRa5TrTMvco
3Ez1Z1aXW7/+d4iObvgWhDt0FxD3cO8G1NezPF+ZSjpEu0Ah0yuMXNdaumwj3ngFD091sohEvB81
C7PvyBPKPG+Rj4SxRa49go5xJfOQ9lJ98YtFnokJUUCnefBXwwxc5RAlk/Ly2yfgCvGPBsdAJ8Sy
8eozMm/p1F5wTnDJ9gszy9Vkct6dfpYtqbstJ9mBUieqzwpPA8BGnhStBjpigDHAYyybup9jc3XN
IzMw4VA6/7S9vmL6kicPsz51Ap73zQnb558WKs1P0GHGqbTeiG4b4pqxn9yLDpZ23EF5g8ZF92d8
AGmNibNv3oRqqiZLi9jOQl2nbjl7NwHja5IxFgyWYxj2GDMcVafu0pO/a81sU0thjYgOKqOXqRcL
Z3nGkE7WzL4UyaIMNSP4M78lNR4nJO/AD4bPnpyBIQZZ2/5IE75Fv/Fmmj6EZlGiGGUPRVxJXEnx
QGyc3328ZDcSZyILTwIhmtzLaZ/QRsnpM2ohE7d1O6uExB7yWEHxXxdH3KfbM5i5C19qN8BKQzjG
6h0Dxy0xLwh0bqMDCCMG9anz3hKdqoxwcqb4RWgn8ykrwWNJ1Z2mYl2hGTJ2iCiKC3F50SsZrrax
KnIkENlFY2EzPNhucNOIk1E1aV/lkshtbQmMcF06rlbFbbAzT13dXHJCJxci+x4wSvOkouwgdR7+
UDbvA6tEyZZRXgcwu2Q+2DQ/sMATRnjcxa5UZA4OWgLXZGbj7+23vyxE6TGuz48H7lNYFs/reClC
xnCF4iiA26uZ5ScrkantVdoLrfuOg/UkqPq6tTsLE1oGpo0o7nP4XxGJpfuF+uxZejC28wQTONBB
jJWp6QGvW7CAVz56e/Ajkpht7JRphfumOXqUTT10v0mAvhPWBIpw5AltuKJd3CxRxdPbFMHi20jK
4E0Vf3LkzQe9vcdnGP1t5o1wOgt21WyImm4cLedEPsgStC5Sy7WpfYVbp9GwPzgYmbhi/vzvMw+o
Xgb6sGqVvWH/0DSNKp5COriFiIQRmD+gKzSEVfcC31cWVZoK852O9DmoyyJ/xLKbYjlfTNHweCCZ
WPWtH+MFigsGTrVaUkf/y0j7jDW0W1tr6jJfE1KYhaOkTBU5+wlo48pqUhLyF9bxlxsM9BkoTeu+
C8KpdriSDjGhNFbLm/jglBKra4P4py+tKwPrnOrmw/1/l+MaVO4NowEjR5LFa24N8Rxfnabh7fHt
maK94Aatnd8Wrjet1wpB49OEugfiPcOIEAQEezPpTsJeCa+ganyQo9glCH2//PnP9MfLzau5Wykp
4jy1DQfo+ikFTmJfkIaotvlAjrz7XVNwlpvaHeht3+Ob4fTS4T5Raff9b1fjnuERkigBBMnxbNXS
N2634ajWAa42yGouMqdPv8oviae8TvSKY6oglRzTTievTIaoHI6xJcyJKd9xWcfNVJ+XQFHcwQCn
fKEBDRL7eT06aaPKioCNXcMMIz1CaELbDTnJ3JTTyDmRwQeDYYXbTdCePo+1AwOWM5N6EU+BWsie
6O7AXacUifPL+Yx0aJbNF2NuOOfVxrXKhTPc1EXQ5y5bbquG1wU8oxOWk7awqT2N2wbdmvedCxC9
RrMzVytQqdtn/YqmTRhoR9JatxROFvrpTV3cGyjiOlo+yi/4C3QwtbWOw4Iihu6W3Xa49b5T2Scu
vM1V4tFQv7kC8o8Y3IYlbzqbxwMZjRJsfNucOSwK6SHKYjcxSzq5iHlvddWrz953tMMjXXYxYMY4
dRW+AsULCiqeF66ZdLIddgKeJQ7FS0ujOGH2nhB/sc6jMO3+6KiRdOwPmZLvNiO61Tsu4etq96Xb
dmnoUBeek34tePTGKvAdxUDsdVIu3KN16P/kO2IHSFLLaFVz1gQ42cAmCJOVX9tsYIrXYaZhtmX1
J+vkJD71v5XC3fK+nWEM05tUFuUwZBJx+K/A2hOy4pnEKha0hkKF7syru+rs4GjQUEB/RP/i2ius
9codydtnrJ2qnQfwhL2boywNB5eGGAsZ24jC8lXW9bK3TaL9vpp0paJrQFkJrA8HJi+Y0E3LRatO
B9EpDG1WSKyq54DxErIODMaFERai755IGNaLJUfPRMmkG3G6jSNO8ahdNtOfyJddDO72sLxegX4P
e6FGcJk2n7f0OFdwbyr+vO/WigFpkGOQTU7blv/nU89LZAQr0bmQhmpKiqLtpgrlkwnrp47uHNl6
qI9cK5cRg1CEC4C+j80K7l8o8pN2uYF7CLXFnvN9dQgoBIkXKjBSGHn02uu4g+CBm0E7jKvr4r8D
sne5pExGHH5Ke34DRfF7d5YIv3mMJABOwDXrOCC2MkqIikc7OTwRQejpwF6F1etvbAppJrDa6C2f
hX+fUVsjAs8PUbN1G9zQIhRrL79cgwydNjJvN6Ceoa2JKclHaSxYaRYhl/Nh295kA+2OoHjbI0jd
WHJbuUG+DTrb8qilB+DMKDm8vRxlTd9nuyGu6Ze02AEcKLF9AZRPXBmVaTR/AzwXAggJKs2BZs0a
C0xamMC8OAYMmmXhU7sf+Hhg6NocdeLNLw0njs8sbCNIWvL8tGsbi6w+KGdMnULrWwlS9PqYaWgV
U1XXPNY3HMdkh0A5D887g2zf5EFbeXM5vtdqWPDGZkssKmyPYm2dZMmM2jAwuBAzJzaylqef1rOU
4SexpqeHInz6WRVzx1rE0j0yGRr/5iaVaydkhnjjLvasWJls5Uc40hSsAsBbB+tcBVKNowE+d3qM
p432MQz9Nbdn/L725ImHb9eVqEgjq7fCGHFQKca21MpZE4G9CZp55hAVzYMc7mDlxl+MscX1BI8l
LrV5ORIQreRTXs+YLOFkCjKBF/hcqpvNk1Nf60gNINtemQU4V505CXk3AMgI1z/7+5nnYwJvmkka
xAKiv54r5HrO+jXI6/F4t8iEUfdXUHmxUdaTetvaPrMwUWS0i/bg7drXBdYtqA1B/TyHOXTo34/O
OCRMlkgStDBNopAL7OgHy2SxXr1PSVOQZt8LEyMyvp7Vw/qv3Mb/ly6MceygavO6QFtPyvir8Rv5
57irkz381zXWNRZidTw7CV6DzfgXPoDnpMxp0uN+QSqSuGktMP7RNQEtIQqZrbtCMHmfHn01KN+h
zpuASJtR8LRGhwQe8Dla1hrdcaMpTA390YZeHLYTDefn9d/17R/ntnnETieoRQYi5Y1eCMeDJ+yI
AQ4u1SpH7fqMC9h4f+TlH/mYA7N9IfdBcAT94dM51l+lU3jcJPR5Czm8vRjJ6Hbk23UC+50LOgqg
3ooeRjreYFLnFytgE3ayn+IoauYkjdHY8Y0IZDWQ2KsqpE2e9iQZ4/K769nwAeG2cnFBclR6J701
zVC+LY23bESeKQznSun5dj+zp3hL+myOUHPpL+HGUsbtZoEOQdUj72Nb/2z4tz6NWeRTR0vpPxOq
3gbYt7kXj1yltRNqT9a6KvQ9FTZeWpPGkU7Ym03RkPgC3GAQ+qlPPEvzAn8TLNJS8Q7eA7dvcMHz
BQsLLAgx0/rswZvpZnd8pWmsH+BN6UQcUUbB0ixsaIUAxdLaXW1t4s8R7M2kp41f92GsEkY5b6U4
f/jZO5aa7IEpJchWKvLqbLGaxhfcky8Se91IVogUV1OxJVfHh+aqc3wicZERaF0hfr6PTMIs/oM6
xnsNKv6T0huPq+lvCjwpvxWizZSj+4YSyurwfXrQQLoVdtzBideYu6w1KZU35DLq27VBXzbq1x4E
WcO2g/EBu3d7URri6iXbHH4hqI32NxQaNDz8TRR7mot8g5bBIjTX6D8mmqrkzc3b6S6nVP5SbaPC
e1yJysqWhgEF81aJUdTWn7UNjiW0Bbw5fSRuHR7WyFvGkB7BmDTmj6MDPhR+2njROOy6wcP5YtQv
2I+QLzhkZIC9pXTNuHtAGt/Jqv4idyYHEbUh+97ioZf+spTDG4GTr5sLRX4jZ5TUQfUHx/MvWz+c
GDuLhpxorKg/uMF6yDyGzfmwbEZ7GfRVVUWAcZaOQHMv5Md+1e9EJNSh1U6MhABjK8gbrWlkWpt1
qaWB9u5OuMj29zR9UqzHtxP58EXcZHFckQojgWneZfEPsrO61c7b5d0FcbewPUaTAJywYFNpS6Eg
HytDrCVsDhqDt/EVFBZG/OouTYuifmaL1EaaHIxhoKeN+17Ed/oRIcpKfWK3POWyDAUY2tx9zOzR
jCzXvgxzfPdoMqHzwzEeXc6MnxFZdN+lnGxJm1ZwtFoFBdNO7EltkQKSKlp+FubkT6Z+nHOAXXpd
zL+idhV9mFFSBgSaQ1xoyejCFE02JjwN18qO8zPLg0qV1lQqm2GTSZF+I6023xaYhIV49TcMYeUb
ut7XFQV6gA4+1JTflW/HjhjsRsSuUNRbA8wnEMf01TVJekdX8dzyQ02jwBHezQJnRQCdsG+ckAxo
h5SX21WkP/ks7TA8DmxnyNys3kk1+xEslCwRQKcm6NNZ/0z9YLdy6WJb3o/oxkXQmGJt3N8+OMc4
0YnMugUY6gfWQTcfyGcAiQgajOInn3di/WvIlqgZ7UfAOQdn5bkYHK3Nnwm0SaumSir9ZUB9YYr7
gTviSU1sUrmGQrxQUyUCbjRImga54Zw6oKb+FWu7onNN+l9/zcNitNzL2A3hrfY9c9LzxLtXJA0p
BgzN6qyh2lEUiSa8lOxh6XlOnyEWAdCKBsJtbZecEs4FGKxxZok3a4rYPy1pMvHvhawZnZX3FqvJ
MrIgm3hthJkRD6YWVQGaCHDu8a1gKn9dVrWV4r1jjqZjYz7seFSHrRRd0PJY7Et/CqwA+cFUQm/k
XzB2U72JZxpdryJmVCg3HrH+bvHXeGWuijAQUzagmOnk4zaADemqKCp6sYoRNFyusRxYSuR6WG89
Ip7m6BCOMJEbcKDnesgW2vcDLMx4L7FnK9TAQXO0D2NBPqoH8nHxpK/Kb4wEwNAPqUPwTdvHzPbI
nKfnMZjczuGCjcc+5V2p3zXGbOpl8+Ta+VONegqm6hSM5XYSsz0Im/RcNeYOrBJg+oMDsAS/TYPe
sxNFTQTBKGdJJOQ0HI7Kowbh4mdgPrbW63nOMMUSJv8fWlqxMbxsAqp/8MhfdktQGKAH4tL3zfyu
oDSmjNN3dA8VZ5O8u3dfi0VG4+oQZx4sZBT81rrCzhxStFOrdweCD3JNy8mlQz7GgaPZuU+aNw3p
K6EUMRL5dxMGuybOj/4v6RSefnCidXVG/UIgHZBt2uFc3SsSTddga268tsbG/XwJdu0ftOFl3Gtg
nRPQyM130HtUI2YB4jzL+cliwV9Grh2cszfzrI9xBskkzfpBOv3jZ/lpT2KRS6DXHAMqX30hTOa7
TxG7zxX6rIUvywRH0f0PNuRUo5n2it/sMAm3724c5+eaCTdoL3X8msp8EoH8vVbv1FIYzv15fHUJ
O0CAQYwVgc0PDokJ6tOSvkKRcpEpq0+JMDkKWz2crkfHzydIfNqyK+rBg1PCXbHHh04QBlZzLhTm
nHXbhjgrUNw8gKWIo90x+ujoUS67PW/+YsdTf+kOz2q+YszP1t0DwrnOq+1Y4xzhkXMRwsy53n3E
KioArwQZrEqw11dnu7PYNYrnp4dAfyYp/5W3AWKskoewzUqT/HvVkISqPMZMcgQ8UpE2LipGsABN
HOTtdTTho8jKGVht0v/WuaTyupYdDrfeS6rc/Mn18K99NZtmrEGRyYsTDD59fyzC61ziTh9nyyE0
7NbsTucgk+47/6zSsVQ/lPhUQnCi73O0hFVkZa9ohMLuKIsfth7ag1ObUNznLoZzExvxB7WyUyQy
pZ1mcnW6UghT0NPN/JdVu9TjQYbg+Jp72+HZlbTdAeL+E9ZLUzKHIUK0UF6dOnP+caMJG6pqpDlj
8odY8xf3Me6M+VUeKKeBeCkzxe8aScAUjUVpeEozbfSL5unnoThfptM0egJB9Z56sAQ6q6puwRcW
GAvV0PfiznH0DbNKOdR8sD7z/w2xRi5a9nxkq1wtY003Duwb2gv/FuSfPHRuIGebHPsee2zDLyVU
zPtaJEGhZTyc+7HNPyxaUUuRpDhC1M8apulHwtpRLjLo7SFhsjXu3AuhRMQ4viQ5A1hKmnLlGBBS
ES/K4tCCTO/QSbA7LOLWcoPu3XZD0pmtSoHboerYJiExNo1R7vKuKgE8JTNMgiFN8iWY4HAFZCOB
v0pPaQjEW0sP2Tq3aMRpDN4iL+2BmzSLyjjPxNn88mRoLyKztLhiIVuTxREq6EAOhf+cgn+jPXqf
0ZQedhYwxdmQWc8KLcKJ6n/hD7ili2xbhGnuv6OS6Pr/VRJDEbJXCPuSBEqIehdLgeJbezWJnM4v
hGgpSjSgIBFnvIN8BgPymZxlx8g5PRxDbbZ8rGbQEfA7rIYK3QVaSoMO/lFdQr5BcsBEMjVR+NC3
dUtJpDEaSTk7/V+nSY7ylNVLD/dDl2NmwtDQ38g+pI7l5pfINOVdtEA38M8wu0drtn/O26CsiQob
YxDPZcMLi/bd25M8VSqiIjpYM9PODqpWI/PHuJVB8QsjSJaC8K58Iq7Kw5i9tlWDZyk3XaY5ul5R
sSu4qf2a9ZtySYGjA/tiKBzfHLMLuq6m3gSxN5o2hmsDbq8BiThQgzOe3qiGFWIWls54KnGG4CY0
fdACgwBv0i4MlwY75db0b9+D04UybjeJdvgXE525rYXKpS5S9SNiwxd7TD25Zs6aOEPMMMro5BWL
tXmZr9YYBGMczN122dEVlQv5iNygPdQdDoQfn2CU0FQxqSqTVSUUxllTuqTulSVVP++HW8C4LzOP
70dZ6utwy1P2nKMoi6QsapJft2nfW1nshRcWPxCSg/sI53xqv74nrH5sfbfQph3TVpapbcQ7bMFY
sPOGdHl9wHhS31cGCUMIYy0psOqSbTzSKOZey5M3FwA4RTOgB8hAn+2yRdSe7rg/ywyH5KsLImuh
ugcN4vFyk5e2d6aJI3rRTYgH1cOUWmzCkj+fbefYP0BpKBdwUqt1ka/GwgEUAqARw1pO5aQr7c8e
NuGn7I/IU04bwpomolmeZaSeryb+q2X12yiMAY+As5CG1wAzTov5qSCJwASRZHtlFqXh2sVUz82B
g47ONBaSsjVJ6ZqxrCVEtkOFcTRrY3kjhUHUy/tALbcYBZJ4E10us25C2KLWUo42RElI9vm4LJKp
SKfnRT9a2+9D2uY55kfYsNbrN/D1wpGuvjBxxf2mxFE0ubgGwEyv7e6pcZVJMiCYvRigW/97VqpG
/KCMmEQu/KYBtQJ3f4XT03/2jZIKkS9FI3VSEseeNfXlWtPZJd5jqkDY3u0RjODKHzKIXMacobWw
OBu7YtU/2v4OgCeVyR4qXxHkzSOhAbKq+Uv1QZldTahiF05UimPgNixeQQ35qyc3LBo8rRvj4oM/
89PbZqqS+c8DdPE3lItMWE2qGXhPdqdhKKOIvRKzSHuMsZr7/69C0/K7OSOPHPQm6YmRwDMrROlD
jiH3ONN2meIgaJ+u3yy1nlR+B32GA0ROgksxsskXZpkJbTxd1ZXUC+ZV/eX+YzQipKxzZ5ohN7uQ
RAFcc/yGoCF6gYFUhsYch09ekAqCvVMPtZmW7WxISDxhymqvdgV2Wp2sms23cGAx0tWQugunMcx7
fVfa/0wkLtqngorwTDyaCqT9TyZhd1q3Nwsk/LYv2EkzXAoRN0TQrc5Ptzgnp3Z49qPceIGotYlg
nL6Mi1wpWPZOW6VOVNPJ8K9f2n/ZnwbwAvjEvvyPNvixPMmBOsKm8A3yfjzYMr3r4qMco2tzxXSN
0qiiI53JPi2jraoGIxfHYWzwzU9Pk/NorKLU759gtITYrn7Nw+dL0Y0I9NSs8qNa3zJYlsm1ASfm
Em2HmhuTs4vfouaYtYePCe+sqbvb+ILJ+ji9BzOdov7vKzgeXfOZgo1agfu9AARUqJLt+jto4Z5W
BTpF2GS7l06ux9MysUSbFN+dfroGRzprnTRZiuj+0zzjWvepFRgp3iOtMQF2SI47Xu6Cg9+pBOt5
lbCQjp4cR2cuHU5lkWbR1RiltCVOjqX1zRbi6Tw9FwNGs6dNWoR/P3IufBAug4mqM6bl+aoVO7pC
AySabq7QJzedltAd+cakpc90oc1QOLiM1FOIkAsfa3N9L/YHXL9sIdXYJHN8YAGJ3Jf4geeZdir0
zR0ypDhdSwrDyf4gwDXV5jXANtWafTfRzJvpvJbEPRuSh5hkArxe1qZ+a1cBSR0ZYrudLdBRyMJk
srr6mGB/Flh3PUBwtbaCzPOusgxEhQ2os04vW+PY1QUgIv2cNv0vtx0PUPP8B1mbjzMJbGvp7hZV
rdXdXxZjxEJGQe9h26EkPQeKDIJBjKfEPiSSf30JveM1570Js7AjPXJ53peNqdT4gPqwfkfRnjUc
TeiVSQijzSbO1to/vQalDmg2UxWcH1N9Oet4byhEYRv9t+gpvKq9S5zm6rZfUYUcJwMh8vqeMBOo
Fc6OrfT/McFkOdfnPRpYaNvq7CgqZblEgpqn3bKAsydd3ex/8JghgxCsgAILwyd/GOKJ9V9MBX9N
JOby76FQAARirtEbdF7msGxAl1ysOLdSakEmIfu3BngaR0Ze8RYr/Y6BhL8xYIt5p7ehNzq2JcL6
lYlC1fOhWOGoIVoVpxexhTa6xoxaIxMAYdRW+L7mRGF3Wjshf+bytI/30rudyXL55P8jx60Fmtdm
I5HMDHGAlkNqzUa2sVHkV7oyiUv/UNGlClDQoGvWArUztHwIuZXvGDqcM5DOLd61vAYi5Hw5DKpH
wLsDid/QJHrsD8+K5k3hX8Eq/2CkF6iuV4+5LWnvi+ibzCQ1E8NBFMKeTAEcYi19k81xClzEazL8
TkuDLQFyC10Zl97mbFWCox+dPBSVwQlqo+cI3GISaJl9XOUKEfGg5dXR6WfwxDhIcq2no6kFsI6z
IB/YvdNiIDUyHHg19M5zECRcGp3rUvMAPlraQ6seIiXScnmCWS/sDFU6ZNqvluYQgnDzKOotyDKv
Is2NyfWOfIC2JmjN2e0zwQ22OdWkdXPd5VA7c7g0M/dkCZSkRVzL2tCFYXVoELGvDHAM82V5R9qZ
u6b3smCGw/kzJxLTkeJR4uPdlVHtsf6H6r1rWUnGqPTBDbXL3LXpHDhAiMjjgXOZkwDfTsYvccEJ
NsT1vzG7pGoz/XoOfrJjem7JTXnpV+ZHdWVGWJzoeSaiNQOvZNtsjPfSSRG40VbD34L9sF+zo16w
awKEH+jq4D8c17o9fXEsuZCXhQdByOxLH2ZDFUMsL/L/whGgZYP1b1B9P8qSmPk/MD3CRaTuytUj
0ukExHXESyygKcyCxyKqOvdFA6crmy1aBzko57LyutSu3bEVlAHP+DFkhI08WQEDWN8xnSo2vsRn
2RsSx7pSO6fuzEQn34AKkGbDGuM/ehI8qxig4pZJZzyNlTz3GFgoV/R3T2SmaXGbi57LJv+/Zir3
3Bqa0MKb9xY1k4dwHa83Uye+vuHlNn7naF9SRt2+d71LEAQaMOYeQgLP2ZndtUKU4YHaf/1NLQsX
wYSvd3CA6xPlqKV/FHcA7aXhnKVr2X2Kkdy6tgMrHEnedR0yd5DtRNLWX6dJw4ps1e/Zw9m+KjUa
1uMhsiynINfGE20CYR1VZqTTCD8owJjSd7GKocFdvujXCIKofbDP/lHAfaHu9utY+0ZfnhRCZwC+
4MiqI2oWtnnWupm04SPpsEN8i6lbUZG8pgqjpFKq0B8KtBABQauNzIG61JB7t0H7TmhFurWX0PxB
9C8Ys89wTJmMsU0nBxZ721GFyjZxMiQk3rClhN9sSm5Kb9PUAoI2soa4wb2gaO8vg/RZIcE+LSav
X94Vv5bQyB+CwIRLL+HIZuZw6LelX8sMUWCB1Vqx8zjVnz/oE1qUI+0RVcZjQM3u99dBrTLIYuJJ
pA9s11V8nptt+BVn8KMpqKozWHau0ftrvu9KL7iNrHhPxOzGtfHN8MHVYlUWhlIkV974f4cgeyCF
+mYtKQoXDemPKq/mAGpfdl0LxWXK6WbR3PsOBgc+J8mCxRPeWVmITgcEBqCvisqu0as4FfrntDDx
l4608+VKP08my8NJn2krPE8cFj8Yg4YQl/lRajEKL1AXDfHpFToTij6rSrFXcZA3Gtg2+11tNm76
aDQUXvhS5/5plFhX8YnAV2BXBTRon0KIXfMC9rjMLkWmIpisFIX2OWHTgzJOKV+iBEuuzckga19j
6CoxcFWE/sK4INEqx0vEOnzjS8eTVOR7IRi4A/deOhxS8xs1TdINiqiEflt9w/fr7/ELsyA1FSPv
NTYafy1AdwWEnE4OZwrzzHJbWhcZzl5pzPjg5d4yq1NmUWD5yt3jAqQogxj4RXfUFp4TvR4NlU5m
C5DFck5NFRaQHr3Dpx9ysl1wS5g1PrzUMGYNvpDYKkNEYWagOKd2dQfQKBUBuaPQ3+i7ZdZC1HYi
CDrhIieEnjszQx2xNREQV3N6WPhkToNsSJ5G6o07HPlbE9JRi+K/10PxmGT4AVUrTOx00sQHzndf
kCRO4z6gsMkD9o31mYfpFfAPNT7KyDwe/WPcaNnXTA4F2XzB4SaDsMz3vrxnJFxqXc4K+cYLhh5V
+WNSpDrCmV1bFToZpD1ChDRUOyHEcgKq/7kGN5pErc+yA90OiZyacp3vjACDRM3dRhoQs0/ij+ZX
izz/rYaA1tqkCDi2SCBNOvWBrKCuU2HG1pieCHz+LQZ99GwyiZUAdKuiFVsxpmIF+W/U7bQeyNk3
1BxaXCK3hHgkakKfVXE7AMaVqJ+o20NwGRAjSUB5qgoFvM+YAi7YzXhkzBW33qrgnXKxlShjJLNG
AAq+PuQU9ZdEuvzCPG8g86vMKAecZ/1n4NQQM1FiAkK4ZQM5MqBifcIJ5YlL3JCjiLDMRlsV3VDr
GCT4LIWYXx5gl2sTYL8+8HKAWyPU7rX60Y45r+BSLn4kk1GKFAuSwdOZCNRF7EVPBXxGY+jOcpVI
fvze3fEAND5/J4qJ33qc9/S798fK3dUkUmGvhVdgGU0IYdhBPHTqX7wZfbgXli6nk/oTuJPRea3g
Uz5HG9Pva0/yDCbBQgfPmt0zbooKHcAz9rvxb3qV/8s5eCxS0ROduXiIpkGCqTLtPtRsjIlNGq1y
WdTyHtJi/AtoaKUGvtGLVN88Z45W6vKzRB9Arfyzi27xA0F8VkT7kzB6FNcij20Xr+8m1PRWX74e
MbO8qrWqkeb48Jl+aJoA15H12zN4RCU9ykuGfw+5q7l6AsJu3BwUJxDrx/hbNIS/bTnjz3eSBO9K
GlXKKf1EQwHU748+lodJ9TWCWqSaOgF1e3rpQMS3H8nnso09GgIk6c+3WK4iTrnjVsEb4B0H8JSL
JKtH405u4kPLXUKODLcKmQDY59WPg7Ip7wWiatg3F3OWoEwO816r+YINu17Fg5XEWs/ZMhNE4i/O
ja/4rC1TiNJhG8Kj7Idz/9hjA8H1SFe43blIyN+dGHYSssnhTf6BcvEarnM9QVgCGWX5fzsXICLy
CIa4y+BOaeKVAhluYTeOQMEAN5GBFXKIctIo0YqW6R69n987s3VAvlreM+RoMuqvBsgZqKUgnlS6
wKMLSTEzp1olxUgq42WiYNttky8at8Up7ZFcY9yglBRZFDZPnZjlSMNC78S22u8xHb9KaFO9d5Jt
XQP8mou6z2+fXfnhIqijaByeDewWrAdqkEltgtRS7WAJtJSBsOFNuBkKVhb+64bGHB+lI46tOupr
+dWf1qR5yTUTlXgyktCSsA3HXKrryfGydSg1nQ84ZJtDbrOehgKCpXr0z+c5G3KuCUuzlPUK4qvP
7fa9QXNSMb62Wn43cQ+3nATaWWg0RpOpSd6q1YOAFQxnMtsV7ID7of+9XCXUYm1dyKUKH2lirodB
UFsl+JFUsdYmW2AnW+qaG0uAHzbjTRemJu5jY7Zh5Q/86xlvvpI9oaD2ozr4eJ3Hlmet6duxrgNB
6vKiUA5DCcHBAD8vp1FL76I/42/FctDiCLEVHzTQHTnji05WZ2Twyove0w9qLt5gsyFbcJaiJ+/Z
uj4uFMUPiri7Hd8gQMxAgeAZB/Sk//AFLLg2oWk98nryjbZzQcKY7v1VB5Vq0BLEG2ykqrzluzn/
pzb2FGrA4CeyZQ55uXykcLjhakaxKLIeCfab2euaK+jhZ26dt42vc00Lh/U+BSugsEy8By3jZek4
mTu9KN59FHITRG6s0QS1KCwiOMwyO9yK4YhVhdDJk7kq+VyD6M3ZUV6UJjxFdJjN2pZg37Nw3TdC
hiRCixPqaRfZGJwAFhXWYlnw/K7M//VpjpF7FGef1i0nFutc3leWqgHH8uc/vSUlSpdhcpNvoeE+
kz5v+VVxLw0iRQlq3cvnvAoZy3sgfDzN8c8TLJjqUbAcNI1OVoBO6EqNahWghOXrpCYlDU/f5inX
HgLne9jjRKilvANN3ppc/sTzY2d9UOp6W6VL8RkLtq4AQ10sOs6nSB2luEDonhBAjSRznH+03E7F
vh+ickekMLosRlVv8n10WEQmGFHp5bAQvDjtGfZucwkWFNwxJtfSJYtmIvcW7rH6gOS71K4Q2swX
rHbOxdEXz85Tz/ya+3bsNZ5ZOFoHIdbJZRzXohNCIXqW2oBjTWUwhoHbDk473H5VzVu1Mds5C4Ds
XygFFFOLdkSeViuqY3tOo5f9UstLGkSlgm+3hgu1mxlKn88VNsTHkl2VXzF3HfN4VMXBoz1W934o
YB4l+G0ytW1pqZQJFBRtbPgTUEeeIIMFFztuqm8Dn45mH7SVn3sbCEL2qHLFZL2MxPMaEp29X0qU
woy6RbA8LtrElR5ikgHSb6Zi0ONRlDs4LofCHkPiyUPKspb1Fg4EnSLW2Bd/ARIq6sE0I8LKSMYL
qa3diicMC4TNi4s0SjXwZhxjuZIVqSQ1WObcwtpnLwiufcV4XbdtI1z6KONfbL6k5ohF4e4+JEwF
KYzk0ubZv26Bd19Ar2edkd+vBcazWq4tYEFqwhAgKQzQdRPL/znzR+AXrDeivjCN1W7tG+DHowE/
BHp4StW8+9/bV0SHgaowPx4fjgaLK7AhD0kAR27ly8uVo18BlMBE85Pwx9tN4iF9o4DNBS1Wp0UZ
oFWo9d/yp59VckzTi6LVjZa1vTJnD9Q2SQxQA0PEyasx198hY1eM1U00/CfXk7vVaEozCHVBY6wR
e6pnsia69Uo1IRP2Knr3+KtylPsMKvezUfyf60xC7Lw7p2gVoUnPGICI9STFiGkpaSQlDFCH/LtV
HV1RILVgm7MoQdjmZ8L+LCMYVmP6TjsRI1MyN0kQcO5x7ITI85UsjwU5U+wcuD9OodCWqQdGW6xJ
3Xy/H4izGvdTRjWc/Jhh7K7js6C+2gm3m5RvkQsWCAh49sWGma4XoYG3WbSictp0N8gREr9o0iTj
dndIB+dElX9ICmi4gXKBTlC1M89222Ie/QglLsqCQ85MhO1trm4bFkbkyJIgJLGzowmeEC4UNJet
6LJUZLyON4jqNQGFzDFOgsFC1aTfRmvD0r48fLaayDHlI18dkvcdvZmVKh72eNbmY8M98SsrcIwR
MAUD3lOhBUtJ6nIBJA909dGIgBNldGJateBlRFo1ng3UHI+k5/S/u9U8/oVv4RTl3irbK+ZvwOgC
FasxgR2hdrHlCiLKCWJRH8Xx8MeaoFJ99yhiqvlkgoOQ8rF0AmWJT2v9va9xzqmA/GR+yu3rr/9a
1dc72Yia5jO9Y/NLKebei0tFR4hFLA+dySMnqPIQC+LfucRAK+Kls/+Hkb66EUczCIr9DItEKJIc
sW7hBAHSy8gPAVAfMy7nsYD4snR+hFwcNi4L1vcW4OrTgbDpRPChDfJDBZH7IrOPXc23VvtKJNuv
kCh4hGp9BkQRH33RbBDz5+WwOX7Nu0OUDufPSb43Q8oRJmAvQeuNgP+jlnd2bl+zM/1UNoVxNgJq
OBxo4P4Tmbu5gN94LBlet4+STlO8SHL3iI4V2W4PcEr4rs0VCOh/rXVgXI2w1oKURfDBRHjQwaQN
GQpqam5Qske5SzerKg0kpqzfDhG+cL9roYvCyE5jk+oT9nL11o25SK107g+wMI83x0aS+OSpnFPC
eIlwpF3vsougmFhVRylsSTkVfC6T9Q9Uhr2j8EXwr8/fuYl3zY3BXD6x9WoRHFW3owS+tKsvQ1Ox
gZonixgfoSPgUasGliBPIRL0OENj5x8V2t9TrctUxK0JrIZSNsafGVqsSPJwHLUGK8aWDXwZXv7r
SQHeF8ZDurmaTdHpTxcYXEmqtRvDOBi4D7V96tRw/z0KwAtAMM/DWaR8N1BKdziMiKkKqZtiyUcG
QmLBzZN182T2P0UlU6J17K00bIx3jYTcG71SSs8yjCwHVvi7fCNEh82Frq73CXD4OS/XGeAo6YwO
XJ54kFXGpxx6ONYu1F1nrLWYNMiQIawvTiCHUwYMENhz3sNWbWVJKfAoTTEAuIW06snF8wRhzvxQ
5YF4cEFERzqOeTcJQsNhCO/sfpjZhTQ+RxeWoVDg2q+eUI73eaugujxpanBF7qqVs6hj2a2KZaKa
oTtS9hBy6R3i5kNVeGlTfehVasTTewYSWbar0QfB8qFyApdQrsTxrb/8LjkPIysj4Doj24kM1vY6
fTCrSGZMDxFpPKHxzuQH0wH5BYEZptL057b9+a2SY2zPfN5Y62VkKxR/LuU57pXBGLSkqkd5WZ+h
9mbNXs58O4xmmBoD1mvluDAIJh9/5agijxu7z8ag7bUDB86wsf+/6UROz6FJD0uReYz+I7NiVmx5
gwVsHJvtD5SKBgMYlz/zMAUm/LBoMtnHE8SHmWKdRYRGxMgxQ1RVOfPP9G8SHE8QjqItLQJ5Vunx
5xm+tlAZccKr+Brsh6K1S7oPlhsQ9D79sEj8QNjVPp2NBay6HBgESoBbl5lvJa2eOFfWFReo7kiF
1yBgxCm+d4WKSRqkyVzLudIf5AV/kKZPuxEagRFmyPZPKibfIaWuYgzJAdssfIDst4/taVCGsvKe
XobRGhZjWKmuKQYUEGVad7amfatSZkfvPbdWyTyyjQ7KBw3U8oLHdY9hbnMXMDNJ58ZsVHqICVbQ
bLn+uHWWTH8EymnCbDTckuY/jKLYtY80F9zBO3czVFDuePWwnbvRMlR/0PZFjxQaWy7x36UYksEV
FyHaIeIJbVekaK56Jyf1k5myD4MKRzYAZvGZBfHBImuf5H1ms+w49FQUYi11teDe6Km9+JYAnU36
dRCeBwVE9FM5kl31AB8iY5uwcFK5Nfr/tP2R574RinESUyp+jjheOtm6DATZu7tTX/v8fG9Rg059
h1nmyP5YnHCDryQKiA9jOGFDGYLVJ/zxozh+Xwer5Fg5zLHKW8LwQId1xq6uaIXek8/lHPHkr9mi
csVaDPREvcpqIStSiPreY1zzHmfN3FJoTRNGPbw9bqIdvH6Uraem4jW4G8dxRkqi8iTsVB60WU49
Eu6mrGlaEcHRRo6Dkgyzyb5Ya6moCHWL4M8p+fLZaopzhzZRGm7d4h1563Hu5RYQ0y38O/73QYVM
jm/15olQCkhkd1vugOsZAwGmRtnvssYpvp03+kMvZSOCzrzYwxkMIb/7gxbBREKgrfG3IxbJT9V0
w2UOQkufgjaavnkQEr44egTdVL8NXSwRJhwe4/4irgXJqZcQXPPMijXnMJ385PBlGBavfBIqTZl0
ab04SEOBMNezZdNpKZr/qdnMMVshErRoLSPTKYht1Gz0jR0VqtpORG0cDTMNu77fsJ58axLfl2SC
qSbdCEVF/tqBLS95bnZu/k1rDYh2BRjccgzl0h5/GcElzETHsqLARjRlzLPG9PDn9GZRlikCyx7B
lMHfSYJJ87XuAMr2eAgFjurhyJ2bniud0/mI5UvA0xwdMizBWolRwq80u5Gnqfa120FBfvoy+Nli
O2wehHSeZxj8dLMKKbGeVbFAJFCFKY4mdijrlPP01GuPYCc2F00WalATXCtVsvVQwXdHUz0qN56A
arUq/tLvmL0RrvS8Z3epMX3uMYGPGp5x3B2C5SM3eS+1AOKqMamHUC7TZf0KZEBkSn3W2iVxNP8p
e55uf6itTeCQ3ylmNXtVvvnNgcKC/ZQEgsXDtsV4OyFDBI6kg5ggPdsSDlwtynyOHiaaPoCerexU
JAeFPXQ2SXKLgOXCxgLSSn/PULHSeWGXiTyoQPNq9AaCKYO6CrcbJ96vpU+93JRu/Gv4bOwYTv6L
mj/6O01a9s5zZXqzjVl4ejy+EFj2itE/Soxpv46DZ6dsczfdCujim/Tt02P5jGFWdlOqWMV5sfVD
VuDzKliTWPh1nEq+FAso3kNDobzzMej98lbxRBfzCcmH8qkIDAQZy0unPCVLLDLJebXX6oSNP72P
g5C8Xxe3wTJDlnGwS+tax6fAIoiOelXSeu5yIaL5DPoCujpVrWKub+VaPrswQrNGR6rxvGA+c62I
Rb51XefO6qIbM+hqYDqaNEkfmGQpHMWHpb6Q2hCUS3I3JpcoJZSNqyrkf/inSoV3IzWvV1GOq/3u
ytBzQ/Z6S/YIz9wdKStmTIvg8hJiu5z6wqbgAW58BCFfnjbtOByyWSQswUGU7pp4Bdcg+MG9V5JX
JvEu95K90Csm+2Im2WPP0rEa1wtIFHFd84vem4R6S78Y4Gn2Qo2wkkZG05BCK0m+DlzTAr1ultxt
znoW17mtMNLPQAJRfWDXso5PLgPXBZ51NbdX2onZ1O3Yh3ZAZ/adkUYqOEM1Ne9hnUhJOWI+bBM8
DQpjliD8ijXofc94DzxdQ6zUGhDtgYMCDBjc0v1PHjbuSOrwRs7yQDk39AQOwgN6AixT/cfSX4jI
D5KGFD7DcJpx5HK2VTEv/N80WGoj9G6BSBCs5D8h/u4Oa9xpbsW8XaSf4N9bJDuxwBmPCFzhE0gn
W095XkwDrreSwcTb9fQNpQUHO8SGHeKMpF7usRKx1A3263l6c0kQSr4jhb9JNELodHzMMyVMRG74
9d5CSHcB/swBXQwAMh59KQ6b9WVhNQ5cP044t5LwOMoLuu9L9qShdOTz5doDOOCX6c+HNnt5WJ4D
2rpe7KWbJEcAovuIga8mJ91IhoU7cErI8rjjuToAojUwHeNBceY8BnuuItKFTxqfgwey6nMZd1Wq
ghB3uhijPUP65njpYFt2y6lKxSKVueHuvE3ik0Drw1BqGWvmc5OnyOw6W4nD85rwJgvVqczb107n
R74qTshxyw4gQ2Ccu1yT/oCXK+JE7JB3+CrIDDzXnxMUhBJ0vxmz3mNnqvONj7Ku1rmHFyQCMJRk
ZC6TCoedSLFo//OHKKm32oGlyFyjy9pKsq9vBwebWJ7O5TUwiraTygs50W8BwM/7B/ZKHLn+PV8x
MkAO7oVwTI7gK4x2uaoB/vm/qzCmyhl3WUUgsl+2Yd9CiZBu1vuz1oWVf5Z3JTrtSPRMnuAEhzbN
O+NX52KuLQiwTujkdhFt3YLakvqHiZbKBPwdp7D5d6KkAPq9dm4/Xe6IvS0lnTFeDcumnAY536sx
+vjppZhoruON77bGQ6OHiEl1nzAbYfaybAYMh58C6bTyTjGx5q4PJaOBji9DpF8DMSc91slnARah
m90dbMyg7R+oHd1ta+r8B5myGVri8vheIcjMV3J9r47DbJX95FKJIf7jzoLz6yVmXlDmis80q388
HmZJ31lZAJNkX8qq1zypR0Ys3y40+A7aaizcDC2et0SIt8F+8Wuoh+gUlrumQrLDLib2GfiDEQHP
WyhDkEbUWFc7k3RbgQBr1QkI9T8nV6rpjjSmMFvA+CANcFVMOlO8tl57Cm9d8wkMtXdRx1/5+k5I
xRQC9Iy3FD5CbpNBdMq34IC9D8xXUJVZIoVeZvsmQL762PIpkZKgO3fRYIx7oOV0lEdtgIiTBh7Y
BliMXqj1CijFPg6qPqYyEl0EGJht9VaonrDSVwu+IYdtT9t2FSNFEehaCxxBkYExaU40UeIA+FyH
tMLcRw7yOozOaLdY/ueAwUgOuPGpT0y06hubQyWkIbxecvULbZkWWL282/GslN20DK9CxiR2nsmx
PvPxJ+eD+DnsMN3aN4N0Oyf06I4h+KElfVEzwjG3IvHDTZ/nzMTLv2E/+l/RX8mGX3ML3UfXwEVF
ID1SPsuYaRLHM885Sd4Do7TbbHK5IH0iX/McAiveGZTlxlObd4qBT3Pjiu9JNTuUjltEcf+EjeAE
KvInGW6fwuek9GbP3pKShtyDpeYxlA1hDiirhWy04YYqPIZEvT+W+cHt7qjjEkwR0aRcOfBRDIfT
Yt6lpM2Z8ft0k5lNS/y9fttSYjGo1OxW/K/l5RrJdm8Bh4gXrNYVUnXrxDeed7RXeiSMZPKvYOnP
ekGgtvj9Jl3Fcfkt1unKL3+rtZGAWYSLAzEV2zH1vjwsxHjEjFKcyYJCZl0GzTIe1P7p03uoF498
Lr0VBUxzdyB8bw7dvxLn4GLW6kET9jsp3INmd5LuePawl6uxq9/rxoxS0/VUjyhZjGpLxQulxEde
XKcQpsLV/o7d+og8vyd5uWnu6RKODPi21RTf5d1T7sTiTYI1Q7GGIdUEHEkJM0Ao4tKvZtR3T+wO
KGjjej7A64m+BKYHFkb2UOtNwPurbYBPphTviBfC31wVcCJLXavTgMoB3WJqlKt1o+XWkQXE3AZ7
qfjRNEnmIcN+iiUe/8O//H3P7G6yGJqydAPpcbdK6+CC3ia25RgVD+K6BS0oNr9WzJs7oOP9qBA0
TaOAR1uz8ebh9omviZRIC9kFI2aTqiUoz13r1ENW9qL/u/mGRBkwih1I/B7QGdw5KzC1iFVmhAfG
4lS5p1Y6z2pfryjSfvPEqsEc2K1JsJQCpTlx10fPW3BDu/GW+zxmcO3phpuSihIEPlMP8lMMoeZO
nPmISp+TztU6IJdD4b+fDhSpgksR4pZyMgTI1hp1RGAvnY2GNK57uLqxle1pV3D63NRFwfX72e0E
KfjZs10KEYwZ/lIxYo82FIKyfVZaoaeV91KBx2ze2DncPr8gVvMagBJ1pS+CnATWJvU1eyjj3C1c
iTzTbM94BDTJ2yE1aqf+YS/vlgABhjoQRE4lJObBwrafTWajq6a+eAFVCkDc04v6aaiNtNmARgmM
JYqk4Kvy4JLqc7IN/Y/s71gslmiAzSejP9+j4cqMFF59rI+zsLfpgdJPxzj8kyOawwIJrrZeICLm
2FbhjDr2dkYXkRUfFROW0ugvV7I+sPtd3JtTsLXcE/XTaUx22Afj9K7RoQqIuGuS9CAYqkhoVzof
3cjI8OIdpyx4QL+7RU0ra6u3Yd/4Xn4/ldyv9agDiE8TVyxOErKd2hiyE+tBliRVfTZXuYq77z+9
RLr60YydEbL/Vo2ze8+YDUBY64VLNt3BNHTC77ITWAudq29mOX9UaZJPxpQAuPiJVo2BuqCSKI8y
rv23wefwT/TIUpbRoq8K1TPcN+2uZxT0I3B0S6NrShko7yYlRfx9FWLgVKwEQCrvOTbeH/R+aLoQ
U7P/AC65NBlk4vfT34/NZ+xeqvfASjjyg5jMohocf1z+IMv43rG0HiNUCgddKSpx56gVXKZOrk4I
lZhXdQzSTdLe2ELooxiSN47qf/bN0f+wdQRz09NIbmQCLh72CPgfIlEyk+evESUfTOY3fK8Bz/CM
EH181gAlG6WRf18sPyWNGIV8Qmu+KcZEk45+gK71rJHRj2mDJUc7fFwze4xUBbVEHJ4yNnph/6zk
1AtWB/gHFcX/Fj+wfsS9Wc0eKIvy+FU2g1N8IV8OVtYDVfGRrb9rfeYyBZmOgCt0vjS06Q+Qeabu
I3K4zH4TvWaKNXgiqjv/saSZA5K7VZKvB4ZC62tdXksTNJ10B2OgVpa3WurPNwz2uOEOUyw/vBhE
tlEV+7tzlstfn5u+vQSQX4v/eC38g1tgVwYgPIhdyEjULzLJ7UrGoRR4G8xWKEcQ5Wt7aJhoctlW
OqEK5oHvQAIXLKVZog9BL86jKAodCEZMV/1hZ33Cssi1k8uqfX2DK4tGAdbf12jGSm2Ln0GxJtX7
i9E51Xc9iEKFafzrjaan84ucNneqr+JN1vvMoJXEUXwEPkeK5N7Rpeb/sFsWcszr6VTT6LTIvfrl
GGG2Sj6ne6806xDbe5DAqvO9rdVozm3yfYRG0b8DNHfX9jqGHh0Hdv2bgup5qHD++gffgL1LD/FG
0Oz6sM3BLUOfEB8OE5uh680ZLF3ftchqYfxCXxp/9WRpCYx8zTFAMXaghyaULGcfWsegXnEhaI7+
LYyCm5X13/SHQiooDVsnIkHdRF9e91Z+Kd4VFYlUR0af2zPOFSOClV7qTuOK95IwFgykMPDvoGXl
vK5N5riobY/PtYhkvD8b8F6IcNHCHb3oGEvGf9jDHBag7U4FXxsfyJxr5s/7SrcCWEOLURO7uYSq
LWO+I2wmk+wS/nwAZEj1FXuaygBBukdyj8cAq4FoHkcByIB3SwPpZyIR4uXZ9u+wMXR+PFCkw3jY
5fXsl59pR7ddiOCnFFdiQTgvis085dpLEhUaCRJpWV3cMhjJFbtKrdk0mbfyObEX/I2utLMUNLDy
6GSM2yPceSo4g0dMCN0L3fC4jmxjQTmCNmS1lPWKnCeK0rs0ncAPSHmDJO3rR1mAwF6mjsmn27uU
u+mzf38+oC1vzW4So1wchzRgvfrz55AfYGljf7NSqVXi7AyU0zqexZkKBStkLH2MVBJsM1gyIrXR
IUJYXdqYJw9UNUBdVK5lqqb/DeP7q5TuW6Op8cjRxtubPRO5DLXwxZaugJ+QT99f3jq9fofF6jkj
pMvb3j7cO2ID/Dy/jy17CP4vcAucvAi2SlIK4ioUAd8oITFQSF3hOFIpBfrg5bTiKuJt+N16xuoB
UICld5GWhjGPQ0IcxstPa/1wGOrI/7Qu4GLy0yMtE6+3SPF8BArQ7/h2rtqaE4ZbZ80+383pliy1
s96dEtJ9sFT1hfDGXGtnygYqlAjEc9QXd9r8PFrn4qgQ0dlYeTVHKvRnlakHub8MeE5NtEV7yIKu
6AE1D/BPI0UCk+se9rTWBVnaG/UOVOPXKA0nYT9vkvNCRqD4+sHhh6QLQxZheWsGymVqzFPpKoPc
1dI7cFyVrzXJQj1IepMTusAnZVTTpL4LNzI8QwWZUW5hLNY8SzLzMY9sgmiZjyQ9NxYCC28JpXmq
9nveapOhGotVpQyFR/eQvB+rCqwJ9rz3eU37WftUpjV6fTrEfJxYibe6zCb509G0/w7JFQfv6Rkb
8ZniXm+qBMTPKMMb5gOm9WbVQSk9FymSPpnzyhuinv3vDjzdPnc0GWtFVpVMipI+nRJJ/JKkiJPN
iq+OD+7dHSEJBbHctxLTKnnBTGhjDDLngo5oxCv/JUzvAQOaoG8UzAqgHfgOHEa09pCH98BLQpxm
dstbLcMmCb3Ry2dK5b+WWoYZbdiCyfqZDFOMaJH9EVNVJAzPUuVjG1mYKaRK2ILk//8END49RhGk
q7LU7jBKak0lBawJeVBLB6AMUR1H80nNIIdrB/Zzr5W7ZnLo7wbrP/tsjwc1Sx5DX5btn+/vtXBb
cjFixupcGW+OYuFVpNDhRtkG6mjor2gr6nkB9O60NH9QSROAFN88Ev1eJetliE5xdhrBB1olOFhM
3jRPbeqDNhaiKyipK5igStJ3JEBfUJDPyzmPu2l4vAPEuDiiQH9vQs8EErPkZGj8SWIt07i9J43z
bu5VhG/WG+I9dje+MW+6ly2e1O9v08Khh6AzL6d0SyxVOFM13pnQieKxzCmqxg7Xr9/fDV4lMPvO
8/lVMx4N1rjZo55fTfVYUlpkqZopun1oaFbNO8OuUxq9NTRixo/P27xv79aDsF/AcyIWS/XPgHc+
J0tTxMEQaV1gBVqSHnmunw4kzgBAlAMw1jQYJBRcQqLnei11mKmmaTekI+qCp66VaySl3aJHYctZ
fRb4hlxt05ulfDv7414NsHH971RUXfnKSqLe4M2tQ/jm48kgscGVJCZC8InHtfHPzkABE+TxJwj9
UFtI2eUSg7Wg/7olpm49Bz+BPzwOVaASUduwAfC3BuPYxBktWN8S3ONATmDmVq+rOqg562ilzep9
Szfo7Nfrnct7ALdg/xH3rikB+bij8Oxy4fieoNUfk/sPC8N8budENku9Y3HUoHJQEXrABONvoUry
HKivMOXSbjUcJr1Cc5+ArEF6LFLWhyozA8RuVi/K4MS/HTMQ9q+ThF3t960rPJC9oFFf0BK/UBI4
X+mKFAtWA2TpQMj41yvvUQ0d0BPuoNd/1Ko5nVrZuVGbHyxY/oAZoCzkv6mtPZZQutptcq91g7/1
ijKwCAIuXox13SCW2evvUkHBs+DDlfEy0M5GAK3a2pFsqioJOgSp4sRDXHoUDMtg77ym3Zj/gvd1
SPezKD0xZoP9K9JNKIc+xsF3CqMfDS/NI+9RP6cSv7nys4Y4rNXRxsnL9Cuo9W5mjLynPueseIxz
Rvq7mcqCrvr7vcp3l0q0Hg123tJ7LGkV9CMDRNjTqrfB+IL5PRSyF26wWYF+rKSvaQtJ/U4+JLeu
wGbcv8ba8vO/KmC0QpeUJwRnnDgabVMt29MlKtjyVjFLfsz7HNtIcsaPXcwHo9ih3O3+v52cojoF
LAcpuLoPTmYmmY62r2IwzvAxnzdDth3mdQGEyLDYFSquUqN/cVkN33OzWWvKoLGBdLQq2AVCavcd
upvnYUFhl0tpCs2txQXrFsAdQgDu35r0hjnCmY1E+ltlYiJJ+8Y9xQ71ijVjXHVDipsdF4gbQMUz
E0lOt1VloabFcAEAUMtEz9Y5PjsV9/BUppxmPIaCrfxOTM0PraLeelHU/Tm2Jj09RECBgRX/y64V
05L9aMZxHXByQCRO93Eg2AHQD3+OAZERehvUg1SjAm7AgMOoUASw8JeK2Ps40K8ZnvTo1nSfAjqL
5LAhuNS1MV6iLGUeTb8XVhgJX+N7U4zZ4d4UPrC0+pjUqOdqY/uEmT/Os2Rmi+hhoX3B1AAWnm1D
MkyXhIJTDGdFmf5GhiYwN2S0nTBZ59xHUj9UASP4ZR/NiIduPxhiv40/jJ2ipI9Z8WCscQaj3N2i
JiU2/uPPhFGqz+uZa4H/1+4oFtI+kIWDyjEYC/quhHoTT+52stOsIzoF+vSwsjacDo4M/XlDjnkm
34tzh2ihosittrjydl6uHxR1QyomY3EFiHkoew90lK+YirSHQYgtgQX+B1XN8B+8IZIwxOaBsqD1
1C9Qr1CVig4GX27+5WKYtkvnA5I3zAT7DIhgDYvOIo669I893eH5DkuiurfPumaZGNhRMRiOl23L
ml/PMvzrjwnm1O6sKRdWhILiTg1oOWMCpqOYrYwOwoQ+GBPunosZmMzDNbhD3xQavhpoj0KUe5Pi
Wkm+NZ8Gg0dS0A0HbHYBzymtdULDf6bVpwL0LWOSbkArTFmWd/B1+pdOyNYKBwRM+hMEte3+8v+j
MmVM+eZItCwsBAXH3WkYCd3OyzwFxe/TKExNgU6hsb//q2ihzq5zpF5hVQaKV5WHuXYT3N2IsQNp
XngGXyyp4EFSY+ZWWdwSGbvocV2zAQPn0ZduwIttFcfaSv3Iz8eQghSSHuyh7xVjsqhG36uyN9sx
TDrze3Nrab/kjOGu0gqiJjyKBJUOvj6PFNoJ1XBF/o2lTw0IfVYUgdpQkJ4IFBv9Ha0GHOmBEhSR
ux7yYZSB5F701C06/lVkOygLvF2wXpCXMxAqwB1TwLNEyIoYcz/dyO53Gxcsp7Qz/xy4gZolBC5P
wVkAl/MDTWNzXapkGPe89raJFMDlz5/vtdYSjP09JsZdmJGZoPbdUOw8aIaoCGI0ZdXk8NGU+K9M
AGr/y8HFLYxBcWTBhZ9QLdNeF0+XrMeocAvxcksNh3tHsHX+V6TcYZGdzVFIlEKM2/KGvVWQLXkU
uJZQyVr4yf62IbdUzXZS7oaM6aCzgVHuYoorMzEwMKc9EzsefxMGD9tra9MY7dxBIaJx8KzwL7oY
oGNpixYa24srqL30ahL8pS8EPILzeoie33iVjfb9n1tNBDceVwedUhIHEaEgWbGpJdYVeJc+U5Ch
GV4XZXEN6Q9Y9LtdNhIWg4MrJucs/837TgJj0ypqFXtyPl61yIE/ZOwGYc5zfCw7QSyuFquGe/PV
7m/aaQ3EVJl7/cPcNAOPj6tLbulNoh6qn1OdXhSGLE3CjwpUhRf27v76uCeGIs2LCI3hV+8z3i2r
+VggkvNjuHuoWlYAZAaUtKRglsdAdv+0AMd7Vft9eMY1N3m2Mj1D8P4EPLKeDuehffuz2KcOABX8
z7Ql/gh4tGtM01g7t50V2zfEMhKXeA8YT3fM2BSgeO8jwQO30b0IVLo6jorUDdD3WECKZU+MfOhH
Ggs9g6crkOO9wcsDBzz3AwqgzJXtroGB3NoUuT3dBiRBBYoafSsLZMAQoFRekcDImOMTPwKkKW/B
Niod1ppbFT6eKnPP24esl6C6vdjLlARmkA4fGEhpeR+9J/0bsvbI5X5N7GSYAFUslhaCstPpe8G2
4n0sdeFTkLv61Lz2uXtl0a7lFOE6Q5GgqjOBdO+7HfdibEBTru20PNnn5N6Vne+HWFiOS0ya8RTu
CDeA+nu7FShXu9gZNVEytxSGosapAPsYmeEvC1/ihQWyjDJhJPXmU5vr3/zEjhWUWnVwToDT/9Ma
fKiXFQYn0PGNUKzOBbrcG0jFDOWZFSyCBYTI3Cl3G292RFY4XTpTLPK1b57zRO1Nurdd1h+teEth
iKsi3dpcsn/iEWVdtu1UvhsG+VppAMfgRQ8j8DoCzo8TEruMm1txz979ClCVdoYIUeEGbGkD7CTQ
soSM7KlZqD8LHUGkZUOTlOGRB4m+Ua4OKOcgMTHl0R9xeh6Bq1H/QrKZD8XaNnMojm6/jS/D4U7L
kwjTl2MweI1XtgMwoUpF8PGa5i+nVoyN5uOStW2u7wSH2zMtgSWs7zlvxAEQr8PkseoNbURqkF3D
Ku/CK5HlNk6ai1NwxxL5SKhqkoY/BkEsUeD+KCHAiBBHgp4NEO6CtBKnqfPyDE0tMfWDrIREknl8
SsR/qaIWbhaK3WbqmcfS+fEK4kB5SasbZmaZPvbwF/KygA2GqVRyvXxiMjZxdGJWGLPx17ZGe43K
JUMfDgwvhYR0RT/6pm4H2BZz3lgxwwFcd8pbISA9plwLTFOylO9fz2SJcdiIvSaUpXVr0lqrWTR4
uR+dKpMUJk6KzaXefozp0PQBjf8WsWMhJmogUyAujd+ekVV80zjsCxGuHORQMG+dC96USZysyKph
2VK1NYXtWLEqgMImKzqD+eYozB/+MyqgJl7I/KeL8Nv5Qk/a2Ge2a4P7yQr9f5ADjP/ErXDbJ6Rr
vQzgwMBuXpyHEEQeS4wb//VHMF15gxDmGtFolEONBecyGcORbREgNhcOAYtGXYcmDkMw8ZR/jFd8
X+A+K62d4VcGgan7D/qho2Ow1C1nLT9DT0kzAXlwWqLuV1zRy91WWk1HqGFHXsxwVCNqeZRR7gSV
HARKZRuTC5isIpKG2UhkLy+yTLxQhctLONxY/5u5G7QI70hbjRXVzxJG9KjmdHRp+2zTF6vX0UVC
odX2gFbbybEDrsceBQgoXpa3+iz9VEE+uF2iGelwRstLI+gn3+ibttiUHsh0lEzp6iXiHNczwQB7
HDtCpox7Xs4tYOHCMqctul80iKawOv2TlhiTxzpKPAs+6huGe3Mtt1n4lD3rhDoJUdkJKgBP2Ccb
93UnLPx1yUJ/eCYUiBpc+mclGh/2WJC3SaBRwHo3Tvok3bz+NcMx29U5zwRNyF1drh/rw1t4S1qR
62bIPNIzivtkrPpCbWxxuYlAkMwtOdWkdn4BHZ8c0omsdPlDmH8LQY2At1kSksWEBQncq/kfQfTa
TAsACCuJVH3JH0a7KyROUNsmdeiJG0yvd/rN8QaN/rM0HRg0xmTTpCFibFQRkwpiYCl/T6I0qPYm
dg4GrjbXGsmyXOdYUcFxiohu/9HIoRn0MGeYXE6bS+gFwkVHW5GPRNfhJbj8FdecUGrxv1ULkBII
+Z/ZPTu9GpFbkomIB8oMFMA1YFsHp/Hg3fXXDaidqiDdLZwWSDyJG65mb10D4aa0hOtIt/jlKGWu
LS2qhvDY0QAULca5b5FOY8Fd8taXaA9emFrJjKJho0kvNj1Ulo4PtzooFavnYjKUds9JMkQ0FV/k
IlV15g8KHpTWWqrJR0ZbEYUpMGRZm6lrgLLAT2yMnOe7xRB5WIzYjER6rHx7HfbliUH7970s2RPl
s0AEYJKorYfnwoqUBJx21aU6p3AmpmD9gKFkuDG2SFw2fEwnONOq7g0QIYKDOCFUY9vGuMgS/N0E
BF38TBwA45NijQUAxtZ8cvi3MbrtNyZ7D6Z2IgWg06Rlw/onwJQIEvy0NC9R8ho3wJcBz3+uYr69
LG/oFV34t+q5E2EUfwDbMJwrScnRO/MqzPsBhRQ7Xn7vKdtVgYtZ3APsuYa7+Jwim49ZKSGLwxHw
Ktypg9rBHCcfIMLP88+4QL7POjmdpnJd1z79DNa+NudWKDbBHNgsiGXr0xY6xRr95UvhoWK9EOHI
iaXcF1RsJTrnk4d/DIHl7BzV9xLCAJwRFZ+MQoTKFboJYM5HBGKxKqY/UBZhwKY/GiXkLSW23bfc
yUJlglFpAEtYPilc39hE6/wq6TO6vkNL8CSGDyLe6mNZXmQw4lrzHo6beeWj0TfvVkewhIL4K1/E
zC+VXKOoMV6tMGi3VPFL8/XMwaMvJr32OkrcMwWntp4NK74EGWRGbf5QFv9QhWcN1qybDjflUOAz
1XSOfXsUZ2TP9rr7cQrob5LrRtiI5u2zQgIOVvjgfqYw+WbTvQdjUJiIc73V+Lbnxh4+yX6LTOii
V9wY8i5I47xv0DujInQ4thAOGQ/7zwNWKZYk5XB4BALZPxG8oBnCbD5SCTdBeXK0CilMvVej/O2r
HxZDkWapR4r1xdFP0FbfHWbWTrBkkxSJZkQ1B/hf4GcRjcvgwvlcPCdPKKExA6WjiLpobj1OYGt5
i0N2RqOvdVeDymleEk+el5ig3Y/+yXvZX4TyqOTEsI4YYy7BWBHtcobAX6YdEr92dp2Y7cFX+TSq
zIlk5xVMcMr1cxmQuBqqIwUPhK/+x8AB025c/HHhCGxIkjH/h2avF6XmzWjSUkDniarIwFsth5Ix
NrKMoVNIzPiaD3s29go/TbbLT1WKIYglcuxQTfVnl7avlPCUjtSCyscirD/Dl58KcjHumNaL9KMe
g/kOclwcWe281WR60UazI31F4mqsyNqxkS97UCFfGujzdNQuS5dQjmkQMBGX7SED+nIWuuHFL+AJ
FhR+HuJJqEYBeZ391pCLl8weqcLfkigbd5uHFIV0W6EXE3KHJTydc3AUN58TC27VCrU3RvKCcSzu
/mFlPKzfGsfI2OWNImZkMB/xVeiv2zZdulVIva0eELw3prDbGzZHDnz1lWWr/pFB0g31UIp9rFl/
Ylnl7zlIeO42X1FvcMRahdDT4Y7nTw3wo/umHiJjEWNLLABZ1kctMCBaDdWPOg2qxvx52+w/eZVS
EQAaZORqk+T30MsOplBBmpB7iOu5gMUImr6UykUielUQkzW4lJCULW9oKvQD2RqMeUkSdy7Lu94K
hZBarqJRhDU8GnIfMHoAz9K/XBQ1hV/5PfUvgwpuwAtaGq03UoDzOhiVF7b5nWEf2gjFif5YyXXX
s7V9w8FxoDqkWZ2dYI5acjjP6lCAd91iM/WdidOfYvA9m6MoNV6nycxQQZrEICocK24jnrbtI/Zx
vZhw0JoK1rQGGNAAx2edJCI49lIA4+iHROjL+niNysy6EdfDYzB3WH9JXzPFTJm6GDBgp5DFF9fS
nFRDVcVLGS91WNxm5fjEEGJpcYn0o1Spgm0tViC4dR4rSs08F3lfEFtduw0Bbz2TFXeZsUX8JG/l
fJrAxqAt70KcO8Avpzi3w0VfNU45EY+q8I7V0/TE/6/LoSHVm3GQiXgS04nrWseWNPzS1fkRMSkN
fJsKjFx3JvLJjiI0X6dSgJEzL4jprxXKzfl4+m6Wj/9ZYoQE4ZBmjDTD4rleSMsYXRaRtL3rX2I+
vWKnYn9Dp4iPU4Y2d35uk+sm/UvngcKLGe2TJbHt6AowP4AhbXkmx3mIwBi3CQMjOTJNzwPHGNUq
PTdrtxnjybXgT0GG7njlhJ7GWltzVTYt1bkpf3pnqSPWTAiXuYNZScfV/zoS5Q3qDIz2rLpObgJ8
pJIiKSJKcYUXgbUA3pAoEJPBmlJASMoS9cdZ1ndOeWNL9A0bUv70KVZ7BZHkXrP3MTeIz758RwD7
UuNYwatMTqx+t1eiwvJduog3bI/lWvzyZlEp7qvx7qCUklzwuGjunQjv9W0Cya/WmUfUFt9s8vBg
W2nnuXkYvOz36NuJBaG8vJxfm6gniALkwW+tayoxoDOVZ4lSb0Nn3OKIMwHXHfifzqY6pUiu/to2
0ZGypL+C72tg1LVMXORBLmjYW+ow67HKDrHEMJ5RJ8Kx5pm1WT6y4a3o9G1NGGOYUJGU6nMquU7g
UvpZ1QYk6t1YvYOFR+tuIeeWuWrzchknGA3Ysg7Eu8LIbZGTjjKBaG+YU3bUX/o4G3WDTFwVf14o
HzPyAxLW7jZP3K+0IygZKSdPHvjxdx239QsB3vOdBe+hEngGAR2k4bKGNbO97mS5JdmdVjHPwvRx
LYVM3SYseyzGAx+0NAUGo794ClCCYDYnrmbbT3sVlSvyiX3WfU3BvC0xmh+ALadJDLcU+yHBiLde
kJm/yWC8PpvQmDLRoZqPDcRI3Y1z7AKU2wM5x823XLMjOmwYtppnnabLvfVXFMx2qJn6wvkP0lIG
tVHiqzWnTOQWznYT6lgUi41+wI2XJeb2C2FsdfhaXZ6SYltvFPrfkf5nwgbZ1qoKsXLEDSI7WlAw
JIOodVy4GF7M9UDFCU9VcIoGTGwg2nRAKzCSvB6dWIRL7Wgb91zWA7MP9FtIedYIQZVKd/SXindW
KFJW2L8RDYDZQqQwNpsH4MsELE1kxEFk+mUwVICHvxemS9Du2qlS3+r+8+kB2GeBmufwHxQS+Je/
0qTXVYyLReQpySB0SFs2PLFxB830+OaFazHw5+cLzsUVMe0QGHDAIC9GTr/kNO10uvraNDkujtte
c93/BpyDpYtB1AEbXwfMr4TPruvwX30v668fnhvDWBwFYvwohVdwOT7DERon0J422L5vRGJWER07
NBOgqVd0WZKtPDd6zlrUdB+ndRPUuzw5AtflMPsCe0DS/YW3vu8wsD4TeItczM0F6HAfTi2pVVUK
vFhY6H2M8NlDzy35RTUiuugpQDDKSeMbyR8Egbd5B4LDhERv9S3DLpTEjylhugKk60wFuI6U/WYU
qTLkE3WcaoA6EUoOWJgtIWHJpHPbaRUNysjIaqsT5HTtayiYsOs4rrG8j4cnR56QtIt9t1c4+rPd
5+k4BRtXAdp3vjyj2sAGi2RgVF1i3ZGEMIX1jWknzIxozZWoAd92wuZIG/lTHqLAtv7KN+EYHemh
VsEVh3ikMGdByPNHxdVhbUd7Ldtz1k/nZYeFNwBT7BsSEWiqjCgatNUt3eJSDVNTbYOnSRj0rrnq
P4e8hoNdG0j0iDWYRxBB80VF99XeZQiRT+XQFjvJ/rxWKIgJDvl55qgSY1K/cT9ao3ltyJH0oc8x
VK7dQOf55cqWjcaOLxqLyZnLBieIw9aBSiX9Q9Vz7vEpAgNF4y//dovxsQJqMxeJMR8n9JxzHXJf
H91BT7p8YA+vuxZEMA1T3NvXQFKZj0GN5CM2uKjRW62nvuvGtSvjWJ2N+3cGfF76mUfnzHkWICgM
IjHwRCbDWWAEImR4S9wfe2gfFWkei9pLHHLfm4CQO6l+RfOp/v7TPA/J2DH87nAANFI0sv2/aYhO
50OmD2lXPDM/NQJo4Kwx40BjLXZmq2uNsjUtUwjpOf48S0ey2/elGpXqbAbKFkXHDZyjIw/oFEPv
ylwmt2ILTazGAJFiZLcVa/7hM3621QTYOMriYx/tcH/OVnt4gg7OVjBWx1T+lFv2fnLLKIS2kW1a
xCr+vPnw1rDt5zLLkk2LGsXqCay+F3hFU3uMpBR+f1IT0l40c6T0brXgFoR+LcyIEQUPFTZ+GOTF
W5ss44L7ObBPHB6K9KUOI0NjUQwMwGPkYGqPsFXVjF9oOXlbe+DFEBHlXBm0epJnPiXLu/ijfQ7L
g0u1fMN260l6X3R+52SkJ42cC1u5nb3sWNKXUp+GBBPffFI6jqMTNsHvep3vsCgEgfMewe3k/YYW
B8Mx3Cw/YA/No37X0kx1q2XNGRF+xbVFvIN3q5Beq9lSBqnr7ahMPAw+tj8BB/szlaVLLKzmbg5L
2ExIbAFtZtQ6v1k/WewDNIgwGQspn9HLz1slWZmXFTM4eHaMwuK/pccSaeTsUSdUI7Jewog3eSQt
RlY9JMd/pSQUu5MjIyPpZ+QgeI66Srkckdg7WxESXd1mek1/G6LSwDBZRJtWkWS9IfEV//Eg72iC
8B9ULwLZRI1NNH3S7sZk0i+SantlHCCIMcAL73/dDjdZtxOhdbxaq5W8JPefp2EH1Q/yvxXwaMoT
L6izHEsOr8zb2DV0naPneaGnP03/yVj/VHdxyoU7OGcyO8OGBHXTH5hFZs9GcsYxGKIlcaTq73Ue
mPAh0+5S1VlQM1lncCyWn38Dasu85Mbr4Qh1ScaO4GH//maILSZI10/Nc1gx+zcH7Eh7UOuaG0yw
JLcyzV5hfss8liT9lZeaK9rRG3TZ3+jBaILBwkgQuFTlUGOXu7r0QNvD0VoqZt9wDcL7xDvvJE+a
L6Mwa0VDkxEDtC2liA1kXeL/u3lzYMa2Wry3XiIbb8aTEdsoWYX4sU4jjL8/4106Z9dIv8EZ8A1D
lDCZCPpFes3lCuW3CmaT4KexDYkmh+8++ohNqDNvlMijT86Ue1JacYM7FK2rXeoIbK7igxbI97Cg
1A/Be4dp6e5AezVMvudrXS2nPy8hd9MQZN4LuleKv0P0AsT+M8SYV53MmuN5ZHdYVz1rIG8y5MwN
ZvY7TxfEWBv5XW79RtOEZnpKpRO6od6Nx/k/fUWbyBu9Rcq/exna7Sc/Kq86MvCHiFntlqvpqoQ3
tK+REZnuXGoZhxwLoi4mjwguQOdltpx7Zq0kc7fP83dMrwqh+amG3BMZm/ntjch091VAHxDIUteG
AHBC23YAxgpPFyNdbK7eGf9GHDnwP2/wFZFA2lsoFeHiWFgVeqk3Vsu6f91gctqDP/U4iN2OMM9a
llJB7X6oqbq8kGhbZB9AZsUcFLjwZM8BSaqZbVkLuJdA5dO8CLejo9tneDP7Rs2QLu4Z3cqXrgLx
arEKCKcJkbzliN0zVIhvoJBxXLkNUekrek7RctvREx9RJnQdkNo6Mk5TTZsMtsXJ5GYKvdA/B8AO
tef/0Meat2xFBgZlsQQTVoQfAzFAjOBGjz3M8C4tkMETfd5QdlX3W46D3VGBg5szD6BzMWN16bh6
dYiXPs6gLI4Nbkz+hrLY5xVteRFoveThgCpNE4fGzZlPhyODp9aNzy7TMp74d9pjNreLObGzrN/2
DhHK/83Iu4tMiGvUD/3BttVENVrL4RHD2DPWBmK1nGUet+fds1G2FmkaI5DSFHR7TM+AJLv9i/ks
XQojealUfQ2Vodax/Zmrgkuk4y2Uw26/7tztvnJLIvxI8C0rhj5OfI/IKj3r0FRNf2Kh4V3WhjdM
4QMmxOm15Qpbj7dqiExVP7TcWtpbg/NfdOQyIUIoE9GhEq0AZsuTSzRfYvgEPN7Il5DsgyLcLEuf
FZLixoRBMKjnlPj+fZPR9cYSWCo+64kN8YS9+lfdcXeTQpZRkTMBXKt0ljiPNNLcdygEVJKkah3u
YFY/VWmOmDzCZAND4fYS/SY0wAZd0ExeTvzAUA8UKIn82yyZEuNi5emVosqn+J5FP1bwkjwZbAjg
3xAqU2bZVVVnXXttd1gL7d3QY8T+3tkvrmF2cho6LBDkB5h8kJ3mC/huTV3UpRHV2HBJUITbxKsU
Dz39UHX+j3G50oxVlScbaXGLEjuxOf9euzhcYKCqf+MWbOnzBXNuKQIikQl+chSt1+X0/jiG++4z
2WSdPIjF5375dpMkos5qyYUPp0NG1c4Ln6zou7Ov5SxM82cK9fm25/qCozeNR3z/6Ceyb48aVFMs
2qdFzm/qQMXhWLFR33EO5gA3QSH9vzQvVdcc0FN+n9rWa8FA1n6FLScOyPrHDa0bhLeE/AvxS7s4
6JO0dUZtFdznV8NDZc1MDsiWXuv9+SfZ4BPpnM/kQ7SCt5zKCNzqdeCwb1lMRlWHsO2R9l4s5sbP
cUhEu7kzS9Io99nF/R2nQkucQrlthRb+TyLU/668JWRo3Id8amEPpKRHgk9YRHUW6GbXOrBAgCJu
eQzqtGC16LSS4OjZOoouF9GoMdiAmx0FNNx594WMWNEWkKiJ1MWENYJ2rZ83/q30H/8UQ1JaHDfS
83bXyFZVSUaLGGjZ1+SV5otjABxiGY3zIF+esNcFNNW63yA0xqVRyVBZT+1QNQj7qkm+uMVU2fH1
pa6LfVTILOhaPNzpStkrtgHEP1k37XSKkgsdDzNjyhqFf7K2/9DZ1plmwA4Jez0cMc2mdiviey0K
X5kx+uQPjMtxMYL+C3g0sjjSYjf+nIusyW01tv1OUrh/LB10jwrsELorxHCl54yrlfJLqNxUG9QE
JX1rigMy2wTbFAOPfqJU5XHns1PWanv+0TTwV0TRnCcZ7UeOuvZvO0FZdVEg3QV5HA9T4XUsuXRF
kPYR8zQgK9cgREanS+p88+cMKQYH0itVsnbEreu3rbKd5FKGLD+WnWO1CajEHItXkh/j5ZdGnoxo
gcrYhRy6AxtNFkaCzJ0WR4An0SQbSXRKPRbfQlPth0I+lN0UI1AP0QyW1E6cETwdHbilJeb62rq1
LWYuwayNkUu4imgEZuwLz2V+v3l+Sc2tHLmCJ1I0tbHcC0CUbxqy1gzxWoedog0Gr4jtNd2r0ZLX
LzmBd8MgHrFZYC+3QfSiOpzGDl5X1mMg6r+sE3iTsX9f3XtL3ahsIRUxcpY1VB6tSZ8BEkUz4Vaz
lYWRuMY8fYYVsDp2iPe/xSZ3cKnF/L5bdVHrO44a9KqdsFjO7Y9nOTvD7tr8L1aWAtWmbt3CXSXd
K+hZwychn+kq8dnbUNHWj7Pj1r0kVhuSWoEVsP7Ubmr2YrGNRq+DzQSn3B+8P8u6drEHMPJZXIMv
fqcnWSSS74kXK9HtdoqAhUDcGw+dr+QF/PIdjR3KdR+uA7STxNXQR9xpdDb+h7b2ZYEgaJGAKIXy
hNYttBVQkGVT8PneCfKyb7oe0Mf1MZCK+0QWOneA4y7fFkMIIKEy9tkf3KBg+5YRptpexmRuoaGb
CXfg3/JD+vevsmiiLWGhwSKW9jXai8TQyRTvETNO4tTb3BdMwsKAGfucxFaBQ3D+u8Q715f1ySzI
DfbWWQV4nu9xSDOnFR9+GM7GvRjlbid2UZ3woNt2mgm9uI5zFwFS9P0UvvrJ5H/k0jrOYzxLswTi
xMPfUb0b3ZUf5Oa4H1Nc2ObhjqdvvQrBwE2wB8JZv07iYYuUPP5WZ++B+coq+5pwDKsX4R76v/Cr
znj2hBV9kRcy2sKU+YXiHx1d4qJ3bWtK6HChigMsdnsUiW8bwfKMuAxzXfwOdqp/wKuvWRql+eCV
XwLgRtiZix0Z716FqsSw0TDN0VHyQDxfl0wMz1Mt58604FIMfi7jr9q6moyPsWjIOT0D+xcRkEIp
SLKwTl4JzExAmw9LgTvp/N90Ri7oN8sk15bkqQRWY3jCs8DzC5Ywzda+5lhiOflWym9YunVUCeIa
q2hjb7S+3wwWpd29RSfvA23dsuHieWSIt5jmna/+b0qvnPsyM2q42QR5ZWJk+PdALsAFCXpjhuO8
SpS9XvCcjZG2FsJjbfV/MRhhOGoyIZr9X+CPr3bchLYN8Ir7DdFA/Bg7sqXUVN+W70gE1nKjO5K+
p+Fd8FWh/ZbvB3r71/R+U1/qHOQqbMtdwyrAIxcWhrjY8PRcrX1P5PqGrrO0XuQeg9O6XK5aKdfW
eRu4ngyxOoVNRgpdyeV77pbXpHaNl5IVO91phfDHIK3+ej49Eol7odBXHIHX0w4s2PitxYRnGthQ
n/fXZjY1m+Z6IzGJ6mP3daYsaOVzPf2lDPGKuzSkhk6GfOpHZ7LO74a00sti7WtFmjFC+MMFbZ/t
TCqo8XWuBoCdzYrUBplmVwMw+pnRgASDfp8SRALGSU8q+ZIIUeUUJkaalHCB4wQbhJR4hU24iKbm
fp7bSXxk2jEaRuVuqT9DCgOAOywkBjNye4F5n0yMnA8FAttG0fQzJ9LotRqunpN6/TQy5Y+Ys7fL
kNo7mDvlbvIQLBLmqG68iigri8RCdKFJMKUtHSwc42i/cs1OMKtkXskGMajI7aXSzx9dvT26Qkba
NbO7Md2hH0AWI8bR6qzIjG6s/4CcLMOz47TQODK+VJGSp/23qpbya47j/5uIM/g3+MBb59jfnfBP
WVFAVLLhRuHEWetf/i4idopRvx64xlxkRit6mt2IrX7KpxV98aUbevWChfL/9NN983TpmZUZcRwV
nhQSHY4KqmV5/pdYODiZK9ItXLCHwqiqezfo4atdTlUF/BVG2S1Z9BV6pqygwLJR8P5ubT32hmYX
2/F8tsWdXx4lgoxJUfPGnGXHWGG5mtxAQAY3v2zEC1DShB6JCrEQEPZFe2GPeTPh22okuNTiKZaj
swvW7C5VKsB0FhKrcYFwEdqW4Qj2uFcePHlT31xnBiAECZzB68QNfWLj2GAPFkrqLEvoUfVBjJSA
SD/IZ17hub0NxOz409DxGUNmucA/VzTIhBUdal9PmSgBI2Ai1w+c7PLl39V/hQFad7mPqojRr+OJ
Y0QVBItQQR+zvuhm+UuMz0ydi4TlC7bpaA5wkwys3FbiNBXe5cVG8b4arUU5B853jjysFDGVDzB4
MYmSkggTxuTXHKEQQeT8YQtXOqPIJALOcblyosy2CoozRflPeZ479ffcCtyC+TBwF2MZ8ut9VtWu
jVN82a3l3/r8Lwzfz+Dz1OVfH4feP2XTqRDxnm+/VpIGkwXE/GMO6cOgsFqjfthdGXZQ4pnaaVqG
Qa3mwSfWV+FX9LmQT1tOKlKxBIrsKPdOJ8qLjiCV9qxkRrUf/RDGjWXE8RF2161sqUn3w4sGLvH1
7quHmUC4//i4EAx5yxWTqCzcmc0B6Aj1waJa35ZiQYiVOF8uT9SESZVTOkOKvfeR+YaFCdwknl8P
dfa4j9Vu0BWgZYVC1jYE1hJEgQdl6LhwXA5DhkR/fTrzqc64ZEwarORv8o7nl77cC/1KvOGUKd2m
HDSqdorg95Ms95Hs+XTTzIMLi0P6cy0SVQEKar0ro51k60n3MzmUsnlwf8+BmG1N2HjrGUvysR6L
ves2v2fcxYGsikmudC9nEjwxL2iuHZxVVY527Pkb3cytLF+LdVy/ymlC8N1JXUl882ag1RZkZazM
DdhjynvFzIVRlgvTyc3/B/R+54uNauxi5jdTCKHPKEnp8gLXuut8jdkkE27ZvJAC6NAB5t/guTir
R1fbtnW3o4+lqGr7HngmxE4zpPXJ65aWe0wJNAh4w5OqIL7wobocuQvIHdoi1yEBSE3T5Z9/yHIu
kO0YokcT7Z/Set966jrBXBtOZOhQUlRWURmnz8f0Npd+fliJbMmOTO/clT0w8PpwyFzQ26LpUDq/
xDP8uCmoNSq/TKgpxnp5k40etH73McHFfsitzmlxst737tsusySq9C/6yNp+Kd1xY3lVS7iY8eQ9
H6yOgklq25ZcOezmHXfmdw7+9zP2Pvefm6DW5xt62jsYvuCsVnKNw4f6a0mEeuAl6uts/5CtkP+0
eokXo/KbVVCf8o6qxiOiAQzWsUsii0ud+of2f3T+Z6ZPEnnVgyYwiVilUwhAAIWPsCnn3u3x+WaU
SNcwGYzlFQKs3OR2xm/WBSUhnQ45FSaIMjn2Z4JeqUybqOnCKVm8EZgFNVPswU/Um5QSnRPvEtSy
/rxUTGJuOZQNpcNYs09KADZwa+Jwf1xEz3qnfy1QtvjEp8pydb1g7JxoyPuZNJnrCAcFsJuM6Qla
av0jeoLmXTDJ1DWGg1UcoOKpmaNEGmez7s7SyIpY6mVnUNofTpMeBOhQjWzbHfE810MxrHJE3TfN
YKsWjqfFuZ6Nt3NLnrKv34v6bysHajzNL6xuUxT8z59JAa9CkMulnSUghZbstCy6RB2sFbXksjXx
xRNwzGBZXIOs4lFl9hoKfjv6KIgy6i2OmgYYGD/rDkUSaIZ5ZiSHqurdX8jJbWDG62iOLmkaMB2m
ZuJqgJYGBIZxF+2j+TUAq9DUIGDGXymMclHCP4xnN8L2/ogftpSaBdtPwSESNTVpWejOo/xVf/+/
/sMOZ5zxqDikn0xeewI2L657KPHjFpGUKMxvpQMCHeLl5+I95hS9+zzWElXwGt7fbtdZ5RhrcllQ
zStnh3YdsOzidxNEzNdpuMibqO2+3Cff0MxrWUeTyYZVgRvlCct+34+kz8upXMONKEDm1wlj/oRe
n0pP+8vi63dl2DTYPA7gNOCD6iDN36vkd+3hnC0mNFfNDMojchmxtLaiya3nXR7OEflILSdEAC6L
cMds4q12/+PdpkZ6fbBAiy/MZR5mF5+1i0QWeSX6h0vN+V3qCfRIzQT44e9jehIYkn97vrXXD1lw
eqgBOpOHVV+vsyuoYjIA4g+KODOMGC/ujpSdD5MK/PkO2cceYaCRDpQK/zJBZG5G0Ae7SBJ2j/2K
9SD+tppQvTXZEwrRRiwhU/BoD4zXnkp6GGfG+hjMahTa2rB97mWW+B0PNZ42vESShZpGcUYYrLeq
Qyj0GmDIwhFJZQD7j2/RNaprPBoirpMxmsbpsIHlMoKSsWUKx58x/d8adDkiV02cOEEnmOQMWSeu
8zb2RND26pThkBu3zaiwWq570LslcVe0RhF7RcErR6AgvQsCXLk0N23g4EfEbPNELq9Fal4vV3Q9
omCNky2uR36yRSaqDnXakThH+NtxqNa/fhzsVsvByKLK88S0sbHCE6JV7Le5gyw7ODIFxdyDrkO3
Jq10uYU4GcbOoPL9zwXjZ/Yv5qyMra69hugZPKDEbW4Xiu9uSxp1L3ByfYClIN/bRSTWnGLbeaAW
4boRjweFhG+S3kqMzS+eU4SxppwZRZCeZP071ab7Uym68J1WC6HfPk9pdhbgEll5b6u8yVMYiCHC
sUV0PDElLAAtj6aOiqXeAoEHFw3j8irlEgAPCjtSjKO5q6m7XTCgNeYIvlan86+eOzPuceZyNBHF
aUHeQhdB14TLI7xAhJpBalZ5jZrJvzBWeDiPQzSmB+JlNxe88d1s2hsO4dAjXgv0iyLbEPRFpgkS
lGEPIiMpO9ESaFHoOcNi2VFsXnITGUEzizxuyFh9WQDzkxrttW+oyYEwURwYKE4B6mqHtmPASzaK
Q23Fuh7EMGypWSfukf20RyJVl+4NbLRjW43vTFMOSEPqS7DfZ8QooDycRcWZnSN1g2pPJwq+Bxib
GuS05i31cyRGofZ3z7Ss1Ocp4sOU9mPllaNy9tZauP0YAlIiJGhNzC3exH2eEson23r9SGgk0H71
ZwecfDoWQK5DJjOu2O0qfQeNBITQlBKCChum51uB7rQhlBc0e00TKZmdeyDbbzSmP9IjttnclbRK
PbA09u0T6a7O7oiuGuOEbEcHHdkSGASM8jQiKeloABf9ka5iEY3sc9iVwFAHzXIjpRCFCXrYkkRm
62saM4UM84h1Kfz+wEs5QBI6DQqPLecaGDrTe7ZyCkBf+94pJPQQDtwoIqylZIEkd5L08KRt6m+J
fx5SDOWafsr50q66KpHrLUsZtiMjW1s0ocvh/UnueqFiCQZrzziICd8GAgWIvmeCEw9GcHRYk/1B
2ztZQN/Kn5nyX1a8o4ikiJj2kMaD/l8T6Wjw9goSbBDKu1RvXkuYHqo7Xp6lRzRqw+Z1Y/2e5T+M
5coF1318/OOMpekrR/3J6cvupSKxtGyj9otYPFUZXLVKueetNXLyIVVmBufTCWwj+nThVKJUKhZF
0LDS7w3alIlPolTcgMI8mjkqrhVHiKmq2HxrmV/Z6AjOArMSf4NF6zrqpBPhyP5q10D4WHrY98UM
ITlEc6UJA+0Ao+nVMcnSxmKqZx0TvLCS1P0cXWRb492KM5X1c8dhmA8xVgND4atRiVJugEZbKyMm
KS9o8LnO+AWt2Y0xdssDzEv97MMNLiHed3vmZI6Kt6Qx9s/o8zC4kQ/0hWNQgJHWsjx2640TVpCp
+qQ/SDCqpeaQ0cTDfl6ahLH78FjtrSHqr4UJWZE+PdZ4lzXHscNbyElnLF0ifHRwv2wYeLm7mSNy
NsT+pZm+5kPamVL/L0vwMQd/riAAMCZnI169wazNmx8diR0RRDy+aNVpj6i9FIBv4glSlHg3Alzi
9nCqWqFmRhZS+0ir2S3aHX2ha9fjU0Z62YaeirQNB5YgsKO57FIT+Qym3KXDTrc3IGBY1bu5dJRb
8HoDbyaxX3ZnSny8F+OGE6J2V0oqU3ESIjT37PcdLt0aXTbnLZe7pw/q65ZH55JISuS6bNqvXVQp
sl77LT4FoBTT/LrVwU6PFhzii4lpeF09MgF2vEQCdwqnGPMQ4zIrpIc13IguV5AobSZ8hHqukoaZ
kyvz6U8UBp0s99OI3Xf1ga44ZrloTQakChTtzcqzC0blR1VuO9nqdIWqSpNI46Q6fnYrB4Zw2g/q
Cwe24gGORSnBiD9RZBsZ90EyCgc7z0qlMlBWd0XqxWgP16cqHe8/yR5loLYLKLdhTtD+0DzWuJ5p
bkp0LuLAdFuSX6FP0YONw4x+C/sUhDGlNSx7eo64goZpUZilvNs+EGnt0ZIvXDUG1dvKBSsIkRnn
at4rxD747QGHIJYlERKCNAFpVp64UHd2xQ4gPSkyM+Si6Get1/FKVdvHEekP0vToaQEA4jiSqFj2
ZIObL76RC+Buva7Z1axoUB3xQrBFhZi+otsSA4rTW1o6H5ClQZ9xMKombsJTJfA/NEt8Jpo5KD5Q
HWCEn7HQIY1Fjgp3/Ok7FY3itEnZ54LcaoE4Jw+dA19h2HbsQ0m+EH9qThZf343ABV1J0A8j/3PU
vdh8MuiQ9rEQpEUC4BiJSb95dQn4wbuGReyowYtA8KeeM9E/c/DEPPTCEztwglG74Jr/DcxABkKL
thsLEEzvr08AN+ABKoMgsa/bmHwbJBj1dUbEOcAO7ogiv+B2srkN/E+Fwgm7ma/0Wvv4vLKGXXqb
R3H0aThOuxT5ONx4DnpXtI2d45+awSDvxyEE1R4NY8rV7WOyMmzx92rCzGVmxoE/EDcbgmUXEglv
bX4W2D7VJGj6x6kmmcFAZcCYSrgLsrTMXRe/ll5lAZ+r+gfnbcCCVRRNLWctTS1xsp1SbjfKnJOk
xbxV2bqc2nT83AmzoimRjHQH5PFYQM4AvFE5hOeO/+JIMeG344LBaYUdjcqgK2UcCnzZgq+3GIdd
w5RCAma300JNCzBe1I74MADeAHxuq7ZJAvFZbn5vWogkKgwJeSO+vQ4Y0C1ES4E3SqO+1Qheexu6
Gn0LdblfOTB66016f9YTbkC0r5In0Zy9/vn6ufBQpm4tWtDHnM7UQK1y6WXndfmELfAYyipkxcWC
EwJ6vkfWv9ukb7W6xyduVcZ8HP5MJMdlmzRzhKK0pTgV1MQ2sPbzzjlxZd9qTgUfMBPMzxnzYMYO
iwMLrrDmmtP6UCzNwiqZowWaVhP+3i1dXg6/v4/0CZaEbgCA3PltuWjEMN8mI0vcc/q9M6XSho8M
4XXHgBhH8qNCQFjsPbXzgaU3Eg/XivSm0UIIpnP7VuRlNmdC5XsdYQdu4aq/SyTJevPq7h5FAayA
d85u+4rGHSXQ7JstqMCVMB/1o6b3gEHr3VyVIJLGHnZm1iGSrWwcJ/e21zsv0PI/wulLquVhax8F
AJCdzpUauFy9DJ2BSxJiaqmQ6+EeE45zFjfJhNB7HWIzjPtdlTjrrrI5g2Q8mg+dhkUDV7sodySb
YMwk2iin4VZKHxT5ujUahCUmkU9WNh7dPkPpt7pYw+hRWFJ8TIeec1PbELLVMPCQEvjuDrrCIm5c
hGefNwg+FCLcASQ1Ckstw54xjZx4nAy7gbAIXudfsKjIylgBf0dvVjstP5wKoYh4NV1p/zCL9xX4
KylNpG2OuZvmvHYJBd5gbsDDhVCy9uxevcTI5o56Gnw66GLmc6h9J3UO6rBbcmkMIefK+INV5Pp1
J9n1/PjzVWLGGtpLeeiQwPeT/P4//FLPQwAjSScBLrLk4gyk6esw12TJ4+Fcq4q+4EHYOaY++ynk
yP3goUyp0uMjaPA7kPM1NiFEnB6eCHkkIbMiNVfFKivTfQQ0QtosuQLPixcZ8QTHmy07gzcu8McJ
uxfjNw9E2nijwa4bHVLVb3q2k4Od3s6CCHa1smUDSqJKMGDjnXVQlqQvroiulFhxCdjRAAkosFlS
zuJIf7iQayLivswv5sV99Od+zIrtHXZy9Ouw6v/ZvoRiEc6/k+2sSxOX3etkL7cAojesslN+7+r9
LMWauAClRt6ZqV+/UJFxIcn0woJ6VMqx6BxKji53fCG4O2DnYA1CfW1+DGMC9Yu1MWFZ1HQiT+1n
YsdDy+MobVglJ3AFxYBygf0H0gUvKizfxdUg709NJT/sNVtFBCEpM8ujouvjlYHdl4Z+W0g9+R79
DT9BgqBR29cZD1Htat3ciNkl4dxobkOCNRMq3EaTdysGbqxsKDF9S6pC28+fg9UBBk30Q8NUrPvZ
ZlLhec3f8UvgZvKgBABdLfZV71FfYddFWC1e4y9I3qKd1epphqanQ4pVgXlFGZy3353r6Btcj2Hn
oF6G8NO44WU/czJeN1vX45DBawmmo1mMBB/mSdQEbvN/t34SFS3jbXNtia52l3M2f0Xv8Y1UrzVb
WhYBsVxiHbNhxUz1EtvkrkUmn5WmSfZ9fX7cV8LMXfMeKI9KQUJr84X9B0sqdrCZQH364vjMZV74
ECmoMd5lwRq5dATFX/5KUSGfyVLYri8Qveq5CbkDC3OHDnlg/NJtc293B1VbW3887cljrmhede+7
dqN+WxqFufrVcEeFcXSCrI6m+wA7aeWCQzG1Qf461Df4iDNGw8Rlw1R0CMnNQPbqyfj0ntEJ02Rt
FXG4zwSxXSysEFrNdwLX4EHdycpoSCw8+aV1H0+4mHPzN7dH3uJHXLx8eAXWGbto83SzzYpJZg5e
r46JbRWMruyZ7uB+kgjSdFnym8DAgnvbc9DlxfWjldvwWeOXa51l/v7aZMjX
`protect end_protected
