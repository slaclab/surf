-------------------------------------------------------------------------------
-- Title      : 
-------------------------------------------------------------------------------
-- File       : Arbiter.vhd
-- Author     : Benjamin Reese  <bareese@slac.stanford.edu>
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2013-04-30
-- Last update: 2013-09-25
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2013 SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

use work.StdRtlPkg.all;
use work.ArbiterPkg.all;

entity Arbiter is
   generic (
      TPD_G          : time     := 1 ns;
      RST_POLARITY_G : sl       := '1';  -- '1' for active high rst, '0' for active low
      RST_ASYNC_G    : boolean  := false;  -- Reset is asynchronous
      REQ_SIZE_G     : positive := 16);
   port (
      clk : in sl;
      rst : in sl := not RST_POLARITY_G;   -- Optional reset

      req      : in  slv(REQ_SIZE_G-1 downto 0);
      selected : out slv(bitSize(REQ_SIZE_G)-1 downto 0);
      valid    : out sl;
      ack      : out slv(REQ_SIZE_G-1 downto 0));
end entity Arbiter;

architecture rtl of Arbiter is

   constant SELECTED_SIZE_C : integer := bitSize(REQ_SIZE_G);

   type RegType is record
      lastSelected : slv(SELECTED_SIZE_C-1 downto 0);
      valid        : sl;
      ack          : slv(REQ_SIZE_G-1 downto 0);
   end record RegType;

   constant REG_RESET_C : RegType :=
      (lastSelected => (others => '0'), valid => '0', ack => (others => '0'));

   signal r   : RegType := REG_RESET_C;
   signal rin : RegType;
   
begin

   comb : process (r, req, rst) is
      variable v    : RegType;
   begin
      v    := r;

      if (req(conv_integer(r.lastSelected)) = '0' or r.valid = '0') then
         arbitrate(req, r.lastSelected, v.lastSelected, v.valid, v.ack);
      end if;

      if (RST_ASYNC_G = false and rst = RST_POLARITY_G) then
         v := REG_RESET_C;
      end if;

      rin      <= v;
      ack      <= r.ack;
      valid    <= r.valid;
      selected <= slv(r.lastSelected);
      
   end process comb;

   seq : process (clk, rst) is
   begin
      if (rising_edge(clk)) then
         r <= rin after TPD_G;
      end if;
      if (RST_ASYNC_G and rst = RST_POLARITY_G) then
         r <= REG_RESET_C after TPD_G;
      end if;
   end process seq;

end architecture rtl;
