/*
 * -------------------------------------------------------------------
 * This Verilog file has been automatically generated from a core originally written
 * in Bluespec SystemVerilog (BSV). The original source code can be found at:
 *
 * Repository: https://github.com/datenlord/blue-crc
 * Author: DatenLord (https://datenlord.github.io/)
 * -------------------------------------------------------------------
 */
//
// Generated by Bluespec Compiler, version 2023.01 (build 52adafa)
//
// On Wed Sep 11 15:19:11 CEST 2024
//
//
// Ports:
// Name                         I/O  size props
// s_axis_tready                  O     1 reg
// m_crc_stream_data              O    32 reg
// m_crc_stream_valid             O     1 reg
// CLK                            I     1 clock
// RST_N                          I     1 reset
// s_axis_tvalid                  I     1
// s_axis_tdata                   I   256 reg
// s_axis_tkeep                   I    32 reg
// s_axis_tlast                   I     1 reg
// s_axis_tuser                   I     1 reg
// m_crc_stream_ready             I     1
//
// No combinational paths from inputs to outputs
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkCrcRawAxiStreamCustomSend(CLK,
			       RST_N,

			       s_axis_tvalid,
			       s_axis_tdata,
			       s_axis_tkeep,
			       s_axis_tlast,
			       s_axis_tuser,

			       s_axis_tready,

			       m_crc_stream_data,

			       m_crc_stream_valid,

			       m_crc_stream_ready);
  input  CLK;
  input  RST_N;

  // action method rawCrcReq_tValid
  input  s_axis_tvalid;
  input  [255 : 0] s_axis_tdata;
  input  [31 : 0] s_axis_tkeep;
  input  s_axis_tlast;
  input  s_axis_tuser;

  // value method rawCrcReq_tReady
  output s_axis_tready;

  // value method rawCrcResp_data
  output [31 : 0] m_crc_stream_data;

  // value method rawCrcResp_valid
  output m_crc_stream_valid;

  // action method rawCrcResp_ready
  input  m_crc_stream_ready;

  // signals for module outputs
  wire [31 : 0] m_crc_stream_data;
  wire m_crc_stream_valid, s_axis_tready;

  // inlined wires
  wire [289 : 0] crc_rawAxiStreamSlave_rawBus_rawBus_dataW_wget;

  // register crc_crcAxiStream_crcRespFifoOut_interCrcRes
  reg [31 : 0] crc_crcAxiStream_crcRespFifoOut_interCrcRes;
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_interCrcRes_D_IN;
  wire crc_crcAxiStream_crcRespFifoOut_interCrcRes_EN;

  // register crc_crcAxiStream_crcRespFifoOut_isFirstFlag
  reg crc_crcAxiStream_crcRespFifoOut_isFirstFlag;
  wire crc_crcAxiStream_crcRespFifoOut_isFirstFlag_D_IN,
       crc_crcAxiStream_crcRespFifoOut_isFirstFlag_EN;

  // ports of submodule crc_crcAxiStream_crcReqBuf
  wire [289 : 0] crc_crcAxiStream_crcReqBuf_D_IN,
		 crc_crcAxiStream_crcReqBuf_D_OUT;
  wire crc_crcAxiStream_crcReqBuf_CLR,
       crc_crcAxiStream_crcReqBuf_DEQ,
       crc_crcAxiStream_crcReqBuf_EMPTY_N,
       crc_crcAxiStream_crcReqBuf_ENQ,
       crc_crcAxiStream_crcReqBuf_FULL_N;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf
  wire [71 : 0] crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_IN,
		crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT;
  wire crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_CLR,
       crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_DEQ,
       crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_EMPTY_N,
       crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_ENQ,
       crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_FULL_N;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_D_OUT_2,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_D_OUT_2,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_D_OUT_2,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_D_OUT_2,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_D_OUT_1,
		crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_D_OUT_3;
  wire [7 : 0] crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_2,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_4,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_5;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf
  wire [31 : 0] crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_D_IN,
		crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_D_OUT;
  wire crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_CLR,
       crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_DEQ,
       crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_EMPTY_N,
       crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_ENQ,
       crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_FULL_N;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_preProcessResBuf
  wire [263 : 0] crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_IN,
		 crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT;
  wire crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_CLR,
       crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_DEQ,
       crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_EMPTY_N,
       crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_ENQ,
       crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_FULL_N;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf
  wire [1031 : 0] crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_IN,
		  crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT;
  wire crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_CLR,
       crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_DEQ,
       crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_EMPTY_N,
       crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_ENQ,
       crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_FULL_N;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf
  wire [1183 : 0] crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_IN,
		  crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT;
  wire crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_CLR,
       crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_DEQ,
       crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_EMPTY_N,
       crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_ENQ,
       crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_FULL_N;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf
  wire [39 : 0] crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_IN,
		crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_OUT;
  wire crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_CLR,
       crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_DEQ,
       crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_EMPTY_N,
       crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_ENQ,
       crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_FULL_N;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf
  wire [263 : 0] crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_IN,
		 crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT;
  wire crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_CLR,
       crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_DEQ,
       crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_EMPTY_N,
       crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_ENQ,
       crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_FULL_N;

  // ports of submodule crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf
  wire [319 : 0] crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_IN,
		 crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT;
  wire crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_CLR,
       crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_DEQ,
       crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_EMPTY_N,
       crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_ENQ,
       crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_FULL_N;

  // ports of submodule crc_rawAxiStreamSlave_rawBus_fifo
  wire [289 : 0] crc_rawAxiStreamSlave_rawBus_fifo_D_IN,
		 crc_rawAxiStreamSlave_rawBus_fifo_D_OUT;
  wire crc_rawAxiStreamSlave_rawBus_fifo_CLR,
       crc_rawAxiStreamSlave_rawBus_fifo_DEQ,
       crc_rawAxiStreamSlave_rawBus_fifo_EMPTY_N,
       crc_rawAxiStreamSlave_rawBus_fifo_ENQ,
       crc_rawAxiStreamSlave_rawBus_fifo_FULL_N;

  // ports of submodule crc_rawBusMaster_fifo
  wire [31 : 0] crc_rawBusMaster_fifo_D_IN, crc_rawBusMaster_fifo_D_OUT;
  wire crc_rawBusMaster_fifo_CLR,
       crc_rawBusMaster_fifo_DEQ,
       crc_rawBusMaster_fifo_EMPTY_N,
       crc_rawBusMaster_fifo_ENQ,
       crc_rawBusMaster_fifo_FULL_N;

  // remaining internal signals
  reg [7 : 0] CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q1,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q2,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q3,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q4,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q5,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q6,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8,
	      CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q43,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q44,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q45,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q46,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q47,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q48,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q49,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q50,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q51,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q52,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q53,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q54,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q55,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q56,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q57,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q58,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q59,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q60,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q61,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q62,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q63,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q64,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q65,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q66,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q67,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q68,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_c_ETC__q42,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_crc_c_ETC__q41,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_crc_crcAx_ETC__q40,
	      CASE_shiftAmt69932_0_0_1_0_2_0_3_crc_crcAxiStr_ETC__q39,
	      CASE_shiftAmt69932_0_0_1_0_2_crc_crcAxiStream__ETC__q38,
	      CASE_shiftAmt69932_0_0_1_crc_crcAxiStream_crcR_ETC__q37,
	      CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q33,
	      CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q34,
	      CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q35,
	      CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q36;
  wire [287 : 0] interCrc__h169911;
  wire [255 : 0] IF_crc_crcAxiStream_crcReqBufD_OUT_BIT_2_THEN_ETC__q69,
		 crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139,
		 preProcessRes_data__h13182,
		 x_data__h64227;
  wire [31 : 0] crcRes__h159813,
		crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132,
		firstHalfRes__h159836,
		firstHalfRes__h159845,
		firstHalfRes__h159854,
		firstHalfRes__h159863,
		firstHalfRes__h162198,
		firstHalfRes__h162982,
		firstHalfRes__h162991,
		firstHalfRes__h164072,
		firstHalfRes__h164856,
		firstHalfRes__h164865,
		firstHalfRes__h164874,
		firstHalfRes__h166516,
		firstHalfRes__h167300,
		firstHalfRes__h167309,
		firstHalfRes__h168390,
		firstHalfRes__h169316,
		firstHalfRes__h287806,
		firstHalfRes__h287815,
		firstHalfRes__h287824,
		firstHalfRes__h287833,
		firstHalfRes__h287842,
		firstHalfRes__h290740,
		firstHalfRes__h291524,
		firstHalfRes__h291533,
		firstHalfRes__h291542,
		firstHalfRes__h293036,
		firstHalfRes__h293820,
		firstHalfRes__h293829,
		firstHalfRes__h293838,
		firstHalfRes__h293847,
		firstHalfRes__h295968,
		firstHalfRes__h296752,
		firstHalfRes__h296761,
		firstHalfRes__h296770,
		firstHalfRes__h298264,
		interCrc__h287463,
		nextInterCrc__h169222,
		nextInterCrc__h169223,
		secondHalfRes__h159837,
		secondHalfRes__h159846,
		secondHalfRes__h159855,
		secondHalfRes__h159864,
		secondHalfRes__h162199,
		secondHalfRes__h162983,
		secondHalfRes__h162992,
		secondHalfRes__h164073,
		secondHalfRes__h164857,
		secondHalfRes__h164866,
		secondHalfRes__h164875,
		secondHalfRes__h166517,
		secondHalfRes__h167301,
		secondHalfRes__h167310,
		secondHalfRes__h168391,
		secondHalfRes__h169317,
		secondHalfRes__h287807,
		secondHalfRes__h287816,
		secondHalfRes__h287825,
		secondHalfRes__h287834,
		secondHalfRes__h290741,
		secondHalfRes__h291525,
		secondHalfRes__h291534,
		secondHalfRes__h293037,
		secondHalfRes__h293821,
		secondHalfRes__h293830,
		secondHalfRes__h293839,
		secondHalfRes__h295969,
		secondHalfRes__h296753,
		secondHalfRes__h296762,
		secondHalfRes__h298265;
  wire [6 : 0] shiftAmt__h169932;
  wire [5 : 0] ctrlSig_shiftAmt__h59003;

  // value method rawCrcReq_tReady
  assign s_axis_tready = crc_rawAxiStreamSlave_rawBus_fifo_FULL_N ;

  // value method rawCrcResp_data
  assign m_crc_stream_data = crc_rawBusMaster_fifo_D_OUT ;

  // value method rawCrcResp_valid
  assign m_crc_stream_valid = crc_rawBusMaster_fifo_EMPTY_N ;

  // submodule crc_crcAxiStream_crcReqBuf
  BluespecFifo2 #(.width(32'd290),
	  .guarded(1'd1)) crc_crcAxiStream_crcReqBuf(.RST(RST_N),
						     .CLK(CLK),
						     .D_IN(crc_crcAxiStream_crcReqBuf_D_IN),
						     .ENQ(crc_crcAxiStream_crcReqBuf_ENQ),
						     .DEQ(crc_crcAxiStream_crcReqBuf_DEQ),
						     .CLR(crc_crcAxiStream_crcReqBuf_CLR),
						     .D_OUT(crc_crcAxiStream_crcReqBuf_D_OUT),
						     .FULL_N(crc_crcAxiStream_crcReqBuf_FULL_N),
						     .EMPTY_N(crc_crcAxiStream_crcReqBuf_EMPTY_N));

  // submodule crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf
  BluespecFifo2 #(.width(32'd72),
	  .guarded(1'd1)) crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf(.RST(RST_N),
									.CLK(CLK),
									.D_IN(crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_IN),
									.ENQ(crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_ENQ),
									.DEQ(crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_DEQ),
									.CLR(crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_CLR),
									.D_OUT(crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT),
									.FULL_N(crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_FULL_N),
									.EMPTY_N(crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_EMPTY_N));

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_0.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable(.CLK(CLK),
													.ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_1),
													.ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_2),
													.ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_3),
													.ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_4),
													.ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_5),
													.D_OUT_1(),
													.D_OUT_2(),
													.D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_D_OUT_3),
													.D_OUT_4(),
													.D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_10.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_11.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_12.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_13.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_14.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_15.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_16.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_17.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_18.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_19.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_1.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable(.CLK(CLK),
													.ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_1),
													.ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_2),
													.ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_3),
													.ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_4),
													.ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_5),
													.D_OUT_1(),
													.D_OUT_2(),
													.D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_D_OUT_3),
													.D_OUT_4(),
													.D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_20.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_21.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_22.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_23.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_24.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_25.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_26.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_27.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_28.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_29.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_2.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable(.CLK(CLK),
													.ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_1),
													.ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_2),
													.ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_3),
													.ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_4),
													.ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_5),
													.D_OUT_1(),
													.D_OUT_2(),
													.D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_D_OUT_3),
													.D_OUT_4(),
													.D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_30.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_31.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_32.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_D_OUT_2),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_33.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_D_OUT_2),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_34.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_D_OUT_2),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_35.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable(.CLK(CLK),
													 .ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_1),
													 .ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_2),
													 .ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_3),
													 .ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_4),
													 .ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_5),
													 .D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_D_OUT_1),
													 .D_OUT_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_D_OUT_2),
													 .D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_D_OUT_3),
													 .D_OUT_4(),
													 .D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_3.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable(.CLK(CLK),
													.ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_1),
													.ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_2),
													.ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_3),
													.ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_4),
													.ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_5),
													.D_OUT_1(),
													.D_OUT_2(),
													.D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_D_OUT_3),
													.D_OUT_4(),
													.D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_4.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable(.CLK(CLK),
													.ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_1),
													.ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_2),
													.ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_3),
													.ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_4),
													.ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_5),
													.D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_D_OUT_1),
													.D_OUT_2(),
													.D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_D_OUT_3),
													.D_OUT_4(),
													.D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_5.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable(.CLK(CLK),
													.ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_1),
													.ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_2),
													.ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_3),
													.ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_4),
													.ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_5),
													.D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_D_OUT_1),
													.D_OUT_2(),
													.D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_D_OUT_3),
													.D_OUT_4(),
													.D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_6.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable(.CLK(CLK),
													.ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_1),
													.ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_2),
													.ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_3),
													.ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_4),
													.ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_5),
													.D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_D_OUT_1),
													.D_OUT_2(),
													.D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_D_OUT_3),
													.D_OUT_4(),
													.D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_7.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable(.CLK(CLK),
													.ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_1),
													.ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_2),
													.ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_3),
													.ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_4),
													.ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_5),
													.D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_D_OUT_1),
													.D_OUT_2(),
													.D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_D_OUT_3),
													.D_OUT_4(),
													.D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_8.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable(.CLK(CLK),
													.ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_1),
													.ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_2),
													.ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_3),
													.ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_4),
													.ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_5),
													.D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_D_OUT_1),
													.D_OUT_2(),
													.D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_D_OUT_3),
													.D_OUT_4(),
													.D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable
  LookupTableLoadSend #(.file("crc_tab_9.mem"),
		    .addr_width(32'd8),
		    .data_width(32'd32),
		    .lo(32'd0),
		    .hi(32'd255),
		    .binary(32'd0)) crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable(.CLK(CLK),
													.ADDR_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_1),
													.ADDR_2(crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_2),
													.ADDR_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_3),
													.ADDR_4(crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_4),
													.ADDR_5(crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_5),
													.D_OUT_1(crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_D_OUT_1),
													.D_OUT_2(),
													.D_OUT_3(crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_D_OUT_3),
													.D_OUT_4(),
													.D_OUT_5());

  // submodule crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf
  BluespecFifo2 #(.width(32'd32),
	  .guarded(1'd1)) crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf(.RST(RST_N),
									 .CLK(CLK),
									 .D_IN(crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_D_IN),
									 .ENQ(crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_ENQ),
									 .DEQ(crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_DEQ),
									 .CLR(crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_CLR),
									 .D_OUT(crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_D_OUT),
									 .FULL_N(crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_FULL_N),
									 .EMPTY_N(crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_EMPTY_N));

  // submodule crc_crcAxiStream_crcRespFifoOut_preProcessResBuf
  BluespecFifo2 #(.width(32'd264),
	  .guarded(1'd1)) crc_crcAxiStream_crcRespFifoOut_preProcessResBuf(.RST(RST_N),
									   .CLK(CLK),
									   .D_IN(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_IN),
									   .ENQ(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_ENQ),
									   .DEQ(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_DEQ),
									   .CLR(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_CLR),
									   .D_OUT(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT),
									   .FULL_N(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_FULL_N),
									   .EMPTY_N(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_EMPTY_N));

  // submodule crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf
  BluespecFifo2 #(.width(32'd1032),
	  .guarded(1'd1)) crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf(.RST(RST_N),
									   .CLK(CLK),
									   .D_IN(crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_IN),
									   .ENQ(crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_ENQ),
									   .DEQ(crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_DEQ),
									   .CLR(crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_CLR),
									   .D_OUT(crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT),
									   .FULL_N(crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_FULL_N),
									   .EMPTY_N(crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_EMPTY_N));

  // submodule crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf
  BluespecFifo2 #(.width(32'd1184),
	  .guarded(1'd1)) crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf(.RST(RST_N),
										.CLK(CLK),
										.D_IN(crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_IN),
										.ENQ(crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_ENQ),
										.DEQ(crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_DEQ),
										.CLR(crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_CLR),
										.D_OUT(crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT),
										.FULL_N(crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_FULL_N),
										.EMPTY_N(crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_EMPTY_N));

  // submodule crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf
  BluespecFifo2 #(.width(32'd40),
	  .guarded(1'd1)) crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf(.RST(RST_N),
									  .CLK(CLK),
									  .D_IN(crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_IN),
									  .ENQ(crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_ENQ),
									  .DEQ(crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_DEQ),
									  .CLR(crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_CLR),
									  .D_OUT(crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_OUT),
									  .FULL_N(crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_FULL_N),
									  .EMPTY_N(crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_EMPTY_N));

  // submodule crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf
  BluespecFifo2 #(.width(32'd264),
	  .guarded(1'd1)) crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf(.RST(RST_N),
									   .CLK(CLK),
									   .D_IN(crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_IN),
									   .ENQ(crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_ENQ),
									   .DEQ(crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_DEQ),
									   .CLR(crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_CLR),
									   .D_OUT(crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT),
									   .FULL_N(crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_FULL_N),
									   .EMPTY_N(crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_EMPTY_N));

  // submodule crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf
  BluespecFifo2 #(.width(32'd320),
	  .guarded(1'd1)) crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf(.RST(RST_N),
									      .CLK(CLK),
									      .D_IN(crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_IN),
									      .ENQ(crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_ENQ),
									      .DEQ(crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_DEQ),
									      .CLR(crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_CLR),
									      .D_OUT(crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT),
									      .FULL_N(crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_FULL_N),
									      .EMPTY_N(crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_EMPTY_N));

  // submodule crc_rawAxiStreamSlave_rawBus_fifo
  BluespecFifo2 #(.width(32'd290),
	  .guarded(1'd1)) crc_rawAxiStreamSlave_rawBus_fifo(.RST(RST_N),
							    .CLK(CLK),
							    .D_IN(crc_rawAxiStreamSlave_rawBus_fifo_D_IN),
							    .ENQ(crc_rawAxiStreamSlave_rawBus_fifo_ENQ),
							    .DEQ(crc_rawAxiStreamSlave_rawBus_fifo_DEQ),
							    .CLR(crc_rawAxiStreamSlave_rawBus_fifo_CLR),
							    .D_OUT(crc_rawAxiStreamSlave_rawBus_fifo_D_OUT),
							    .FULL_N(crc_rawAxiStreamSlave_rawBus_fifo_FULL_N),
							    .EMPTY_N(crc_rawAxiStreamSlave_rawBus_fifo_EMPTY_N));

  // submodule crc_rawBusMaster_fifo
  BluespecFifo2 #(.width(32'd32), .guarded(1'd1)) crc_rawBusMaster_fifo(.RST(RST_N),
								.CLK(CLK),
								.D_IN(crc_rawBusMaster_fifo_D_IN),
								.ENQ(crc_rawBusMaster_fifo_ENQ),
								.DEQ(crc_rawBusMaster_fifo_DEQ),
								.CLR(crc_rawBusMaster_fifo_CLR),
								.D_OUT(crc_rawBusMaster_fifo_D_OUT),
								.FULL_N(crc_rawBusMaster_fifo_FULL_N),
								.EMPTY_N(crc_rawBusMaster_fifo_EMPTY_N));

  // inlined wires
  assign crc_rawAxiStreamSlave_rawBus_rawBus_dataW_wget =
	     { s_axis_tdata, s_axis_tkeep, s_axis_tlast, s_axis_tuser } ;

  // register crc_crcAxiStream_crcRespFifoOut_interCrcRes
  assign crc_crcAxiStream_crcRespFifoOut_interCrcRes_D_IN =
	     crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_OUT[7] ?
	       32'hFFFFFFFF :
	       nextInterCrc__h169223 ;
  assign crc_crcAxiStream_crcRespFifoOut_interCrcRes_EN =
	     crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_EMPTY_N &&
	     (!crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_OUT[7] ||
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_FULL_N) ;

  // register crc_crcAxiStream_crcRespFifoOut_isFirstFlag
  assign crc_crcAxiStream_crcRespFifoOut_isFirstFlag_D_IN =
	     crc_crcAxiStream_crcReqBuf_D_OUT[1] ;
  assign crc_crcAxiStream_crcRespFifoOut_isFirstFlag_EN =
	     crc_crcAxiStream_crcReqBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_FULL_N ;

  // submodule crc_crcAxiStream_crcReqBuf
  assign crc_crcAxiStream_crcReqBuf_D_IN =
	     crc_rawAxiStreamSlave_rawBus_fifo_D_OUT ;
  assign crc_crcAxiStream_crcReqBuf_ENQ =
	     crc_rawAxiStreamSlave_rawBus_fifo_EMPTY_N &&
	     crc_crcAxiStream_crcReqBuf_FULL_N ;
  assign crc_crcAxiStream_crcReqBuf_DEQ =
	     crc_crcAxiStream_crcReqBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_FULL_N ;
  assign crc_crcAxiStream_crcReqBuf_CLR = 1'b0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf
  assign crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_IN =
	     { crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_OUT[39:8],
	       crc_crcAxiStream_crcRespFifoOut_interCrcRes,
	       crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_OUT[7:0] } ;
  assign crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_ENQ =
	     crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_EMPTY_N &&
	     (!crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_OUT[7] ||
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_FULL_N) &&
	     crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_OUT[7] ;
  assign crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_DEQ =
	     crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_CLR = 1'b0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_1 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[7:0] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[63:56] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[87:80] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[71:64] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[95:88] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[79:72] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[103:96] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[87:80] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[111:104] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[95:88] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[119:112] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[103:96] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[127:120] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[111:104] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[135:128] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[119:112] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[143:136] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[127:120] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[151:144] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[135:128] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[159:152] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_1 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[15:8] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[143:136] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[167:160] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[151:144] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[175:168] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[159:152] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[183:176] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[167:160] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[191:184] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[175:168] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[199:192] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[183:176] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[207:200] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[191:184] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[215:208] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[199:192] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[223:216] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[207:200] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[231:224] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[215:208] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[239:232] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_1 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[23:16] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[223:216] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[247:240] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[231:224] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[255:248] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[239:232] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_2 =
	     crc_crcAxiStream_crcRespFifoOut_interCrcRes[7:0] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[263:256] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[247:240] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_2 =
	     crc_crcAxiStream_crcRespFifoOut_interCrcRes[15:8] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[271:264] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[255:248] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_2 =
	     crc_crcAxiStream_crcRespFifoOut_interCrcRes[23:16] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[279:272] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[263:256] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_2 =
	     crc_crcAxiStream_crcRespFifoOut_interCrcRes[31:24] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[287:280] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_1 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[31:24] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[15:8] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[39:32] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[23:16] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[47:40] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[31:24] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[55:48] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[39:32] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[63:56] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[47:40] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[71:64] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_1 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[55:48] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_2 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_3 =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[79:72] ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_4 =
	     8'h0 ;
  assign crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_ADDR_5 =
	     8'h0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf
  assign crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_D_IN =
	     { ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[0],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[1],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[2],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[3],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[4],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[5],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[6],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[7],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[8],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[9],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[10],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[11],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[12],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[13],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[14],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[15],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[16],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[17],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[18],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[19],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[20],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[21],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[22],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[23],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[24],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[25],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[26],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[27],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[28],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[29],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[30],
	       ~crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132[31] } ;
  assign crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_ENQ =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_DEQ =
	     crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_EMPTY_N &&
	     crc_rawBusMaster_fifo_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_CLR = 1'b0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_preProcessResBuf
  assign crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_IN =
	     { preProcessRes_data__h13182,
	       crc_crcAxiStream_crcReqBuf_D_OUT[1],
	       crc_crcAxiStream_crcRespFifoOut_isFirstFlag,
	       ctrlSig_shiftAmt__h59003 } ;
  assign crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_ENQ =
	     crc_crcAxiStream_crcReqBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_DEQ =
	     crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_CLR = 1'b0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf
  assign crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_IN =
	     { crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_D_OUT_1,
	       crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_OUT[7:0] } ;
  assign crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_ENQ =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_DEQ =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_CLR = 1'b0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf
  assign crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_IN =
	     { crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_31_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_30_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_29_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_28_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_27_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_26_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_25_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_24_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_23_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_22_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_21_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_20_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_19_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_18_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_17_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_16_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_15_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_14_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_13_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_12_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_11_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_10_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_9_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_8_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_7_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_6_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_5_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_4_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_3_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_2_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_1_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_crcTabVec_0_lookupTable_lookupTable_D_OUT_3,
	       crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_OUT[319:288] } ;
  assign crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_ENQ =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_DEQ =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_CLR = 1'b0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf
  assign crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_IN =
	     { crcRes__h159813,
	       crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[7:0] } ;
  assign crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_ENQ =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_DEQ =
	     crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_EMPTY_N &&
	     (!crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_OUT[7] ||
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_FULL_N) ;
  assign crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_CLR = 1'b0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf
  assign crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_D_IN =
	     { x_data__h64227,
	       crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[7:0] } ;
  assign crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_ENQ =
	     crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_DEQ =
	     crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_shiftInputResBuf_CLR = 1'b0 ;

  // submodule crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf
  assign crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_D_IN =
	     { crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[71:40],
	       interCrc__h169911 } ;
  assign crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_ENQ =
	     crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_DEQ =
	     crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_EMPTY_N &&
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_FULL_N ;
  assign crc_crcAxiStream_crcRespFifoOut_shiftInterCrcResBuf_CLR = 1'b0 ;

  // submodule crc_rawAxiStreamSlave_rawBus_fifo
  assign crc_rawAxiStreamSlave_rawBus_fifo_D_IN =
	     crc_rawAxiStreamSlave_rawBus_rawBus_dataW_wget ;
  assign crc_rawAxiStreamSlave_rawBus_fifo_ENQ =
	     crc_rawAxiStreamSlave_rawBus_fifo_FULL_N && s_axis_tvalid ;
  assign crc_rawAxiStreamSlave_rawBus_fifo_DEQ =
	     crc_rawAxiStreamSlave_rawBus_fifo_EMPTY_N &&
	     crc_crcAxiStream_crcReqBuf_FULL_N ;
  assign crc_rawAxiStreamSlave_rawBus_fifo_CLR = 1'b0 ;

  // submodule crc_rawBusMaster_fifo
  assign crc_rawBusMaster_fifo_D_IN =
	     crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_D_OUT ;
  assign crc_rawBusMaster_fifo_ENQ =
	     crc_crcAxiStream_crcRespFifoOut_finalCrcResBuf_EMPTY_N &&
	     crc_rawBusMaster_fifo_FULL_N ;
  assign crc_rawBusMaster_fifo_DEQ =
	     crc_rawBusMaster_fifo_EMPTY_N && m_crc_stream_ready ;
  assign crc_rawBusMaster_fifo_CLR = 1'b0 ;

  // remaining internal signals
  assign IF_crc_crcAxiStream_crcReqBufD_OUT_BIT_2_THEN_ETC__q69 =
	     crc_crcAxiStream_crcReqBuf_D_OUT[2] ? 256'd1 : 256'd0 ;
  assign crcRes__h159813 = firstHalfRes__h159836 ^ secondHalfRes__h159837 ;
  assign crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139 =
	     { crc_crcAxiStream_crcReqBuf_D_OUT[33],
	       crc_crcAxiStream_crcReqBuf_D_OUT[33],
	       crc_crcAxiStream_crcReqBuf_D_OUT[33],
	       crc_crcAxiStream_crcReqBuf_D_OUT[33],
	       crc_crcAxiStream_crcReqBuf_D_OUT[33],
	       crc_crcAxiStream_crcReqBuf_D_OUT[33],
	       crc_crcAxiStream_crcReqBuf_D_OUT[33],
	       crc_crcAxiStream_crcReqBuf_D_OUT[33:32],
	       crc_crcAxiStream_crcReqBuf_D_OUT[32],
	       crc_crcAxiStream_crcReqBuf_D_OUT[32],
	       crc_crcAxiStream_crcReqBuf_D_OUT[32],
	       crc_crcAxiStream_crcReqBuf_D_OUT[32],
	       crc_crcAxiStream_crcReqBuf_D_OUT[32],
	       crc_crcAxiStream_crcReqBuf_D_OUT[32],
	       crc_crcAxiStream_crcReqBuf_D_OUT[32:31],
	       crc_crcAxiStream_crcReqBuf_D_OUT[31],
	       crc_crcAxiStream_crcReqBuf_D_OUT[31],
	       crc_crcAxiStream_crcReqBuf_D_OUT[31],
	       crc_crcAxiStream_crcReqBuf_D_OUT[31],
	       crc_crcAxiStream_crcReqBuf_D_OUT[31],
	       crc_crcAxiStream_crcReqBuf_D_OUT[31],
	       crc_crcAxiStream_crcReqBuf_D_OUT[31:30],
	       crc_crcAxiStream_crcReqBuf_D_OUT[30],
	       crc_crcAxiStream_crcReqBuf_D_OUT[30],
	       crc_crcAxiStream_crcReqBuf_D_OUT[30],
	       crc_crcAxiStream_crcReqBuf_D_OUT[30],
	       crc_crcAxiStream_crcReqBuf_D_OUT[30],
	       crc_crcAxiStream_crcReqBuf_D_OUT[30],
	       crc_crcAxiStream_crcReqBuf_D_OUT[30:29],
	       crc_crcAxiStream_crcReqBuf_D_OUT[29],
	       crc_crcAxiStream_crcReqBuf_D_OUT[29],
	       crc_crcAxiStream_crcReqBuf_D_OUT[29],
	       crc_crcAxiStream_crcReqBuf_D_OUT[29],
	       crc_crcAxiStream_crcReqBuf_D_OUT[29],
	       crc_crcAxiStream_crcReqBuf_D_OUT[29],
	       crc_crcAxiStream_crcReqBuf_D_OUT[29:28],
	       crc_crcAxiStream_crcReqBuf_D_OUT[28],
	       crc_crcAxiStream_crcReqBuf_D_OUT[28],
	       crc_crcAxiStream_crcReqBuf_D_OUT[28],
	       crc_crcAxiStream_crcReqBuf_D_OUT[28],
	       crc_crcAxiStream_crcReqBuf_D_OUT[28],
	       crc_crcAxiStream_crcReqBuf_D_OUT[28],
	       crc_crcAxiStream_crcReqBuf_D_OUT[28:27],
	       crc_crcAxiStream_crcReqBuf_D_OUT[27],
	       crc_crcAxiStream_crcReqBuf_D_OUT[27],
	       crc_crcAxiStream_crcReqBuf_D_OUT[27],
	       crc_crcAxiStream_crcReqBuf_D_OUT[27],
	       crc_crcAxiStream_crcReqBuf_D_OUT[27],
	       crc_crcAxiStream_crcReqBuf_D_OUT[27],
	       crc_crcAxiStream_crcReqBuf_D_OUT[27:26],
	       crc_crcAxiStream_crcReqBuf_D_OUT[26],
	       crc_crcAxiStream_crcReqBuf_D_OUT[26],
	       crc_crcAxiStream_crcReqBuf_D_OUT[26],
	       crc_crcAxiStream_crcReqBuf_D_OUT[26],
	       crc_crcAxiStream_crcReqBuf_D_OUT[26],
	       crc_crcAxiStream_crcReqBuf_D_OUT[26],
	       crc_crcAxiStream_crcReqBuf_D_OUT[26:25],
	       crc_crcAxiStream_crcReqBuf_D_OUT[25],
	       crc_crcAxiStream_crcReqBuf_D_OUT[25],
	       crc_crcAxiStream_crcReqBuf_D_OUT[25],
	       crc_crcAxiStream_crcReqBuf_D_OUT[25],
	       crc_crcAxiStream_crcReqBuf_D_OUT[25],
	       crc_crcAxiStream_crcReqBuf_D_OUT[25],
	       crc_crcAxiStream_crcReqBuf_D_OUT[25:24],
	       crc_crcAxiStream_crcReqBuf_D_OUT[24],
	       crc_crcAxiStream_crcReqBuf_D_OUT[24],
	       crc_crcAxiStream_crcReqBuf_D_OUT[24],
	       crc_crcAxiStream_crcReqBuf_D_OUT[24],
	       crc_crcAxiStream_crcReqBuf_D_OUT[24],
	       crc_crcAxiStream_crcReqBuf_D_OUT[24],
	       crc_crcAxiStream_crcReqBuf_D_OUT[24:23],
	       crc_crcAxiStream_crcReqBuf_D_OUT[23],
	       crc_crcAxiStream_crcReqBuf_D_OUT[23],
	       crc_crcAxiStream_crcReqBuf_D_OUT[23],
	       crc_crcAxiStream_crcReqBuf_D_OUT[23],
	       crc_crcAxiStream_crcReqBuf_D_OUT[23],
	       crc_crcAxiStream_crcReqBuf_D_OUT[23],
	       crc_crcAxiStream_crcReqBuf_D_OUT[23:22],
	       crc_crcAxiStream_crcReqBuf_D_OUT[22],
	       crc_crcAxiStream_crcReqBuf_D_OUT[22],
	       crc_crcAxiStream_crcReqBuf_D_OUT[22],
	       crc_crcAxiStream_crcReqBuf_D_OUT[22],
	       crc_crcAxiStream_crcReqBuf_D_OUT[22],
	       crc_crcAxiStream_crcReqBuf_D_OUT[22],
	       crc_crcAxiStream_crcReqBuf_D_OUT[22:21],
	       crc_crcAxiStream_crcReqBuf_D_OUT[21],
	       crc_crcAxiStream_crcReqBuf_D_OUT[21],
	       crc_crcAxiStream_crcReqBuf_D_OUT[21],
	       crc_crcAxiStream_crcReqBuf_D_OUT[21],
	       crc_crcAxiStream_crcReqBuf_D_OUT[21],
	       crc_crcAxiStream_crcReqBuf_D_OUT[21],
	       crc_crcAxiStream_crcReqBuf_D_OUT[21:20],
	       crc_crcAxiStream_crcReqBuf_D_OUT[20],
	       crc_crcAxiStream_crcReqBuf_D_OUT[20],
	       crc_crcAxiStream_crcReqBuf_D_OUT[20],
	       crc_crcAxiStream_crcReqBuf_D_OUT[20],
	       crc_crcAxiStream_crcReqBuf_D_OUT[20],
	       crc_crcAxiStream_crcReqBuf_D_OUT[20],
	       crc_crcAxiStream_crcReqBuf_D_OUT[20:19],
	       crc_crcAxiStream_crcReqBuf_D_OUT[19],
	       crc_crcAxiStream_crcReqBuf_D_OUT[19],
	       crc_crcAxiStream_crcReqBuf_D_OUT[19],
	       crc_crcAxiStream_crcReqBuf_D_OUT[19],
	       crc_crcAxiStream_crcReqBuf_D_OUT[19],
	       crc_crcAxiStream_crcReqBuf_D_OUT[19],
	       crc_crcAxiStream_crcReqBuf_D_OUT[19:18],
	       crc_crcAxiStream_crcReqBuf_D_OUT[18],
	       crc_crcAxiStream_crcReqBuf_D_OUT[18],
	       crc_crcAxiStream_crcReqBuf_D_OUT[18],
	       crc_crcAxiStream_crcReqBuf_D_OUT[18],
	       crc_crcAxiStream_crcReqBuf_D_OUT[18],
	       crc_crcAxiStream_crcReqBuf_D_OUT[18],
	       crc_crcAxiStream_crcReqBuf_D_OUT[18:17],
	       crc_crcAxiStream_crcReqBuf_D_OUT[17],
	       crc_crcAxiStream_crcReqBuf_D_OUT[17],
	       crc_crcAxiStream_crcReqBuf_D_OUT[17],
	       crc_crcAxiStream_crcReqBuf_D_OUT[17],
	       crc_crcAxiStream_crcReqBuf_D_OUT[17],
	       crc_crcAxiStream_crcReqBuf_D_OUT[17],
	       crc_crcAxiStream_crcReqBuf_D_OUT[17:16],
	       crc_crcAxiStream_crcReqBuf_D_OUT[16],
	       crc_crcAxiStream_crcReqBuf_D_OUT[16],
	       crc_crcAxiStream_crcReqBuf_D_OUT[16],
	       crc_crcAxiStream_crcReqBuf_D_OUT[16],
	       crc_crcAxiStream_crcReqBuf_D_OUT[16],
	       crc_crcAxiStream_crcReqBuf_D_OUT[16],
	       crc_crcAxiStream_crcReqBuf_D_OUT[16:15],
	       crc_crcAxiStream_crcReqBuf_D_OUT[15],
	       crc_crcAxiStream_crcReqBuf_D_OUT[15],
	       crc_crcAxiStream_crcReqBuf_D_OUT[15],
	       crc_crcAxiStream_crcReqBuf_D_OUT[15],
	       crc_crcAxiStream_crcReqBuf_D_OUT[15],
	       crc_crcAxiStream_crcReqBuf_D_OUT[15],
	       crc_crcAxiStream_crcReqBuf_D_OUT[15:14],
	       crc_crcAxiStream_crcReqBuf_D_OUT[14],
	       crc_crcAxiStream_crcReqBuf_D_OUT[14],
	       crc_crcAxiStream_crcReqBuf_D_OUT[14],
	       crc_crcAxiStream_crcReqBuf_D_OUT[14],
	       crc_crcAxiStream_crcReqBuf_D_OUT[14],
	       crc_crcAxiStream_crcReqBuf_D_OUT[14],
	       crc_crcAxiStream_crcReqBuf_D_OUT[14:13],
	       crc_crcAxiStream_crcReqBuf_D_OUT[13],
	       crc_crcAxiStream_crcReqBuf_D_OUT[13],
	       crc_crcAxiStream_crcReqBuf_D_OUT[13],
	       crc_crcAxiStream_crcReqBuf_D_OUT[13],
	       crc_crcAxiStream_crcReqBuf_D_OUT[13],
	       crc_crcAxiStream_crcReqBuf_D_OUT[13],
	       crc_crcAxiStream_crcReqBuf_D_OUT[13:12],
	       crc_crcAxiStream_crcReqBuf_D_OUT[12],
	       crc_crcAxiStream_crcReqBuf_D_OUT[12],
	       crc_crcAxiStream_crcReqBuf_D_OUT[12],
	       crc_crcAxiStream_crcReqBuf_D_OUT[12],
	       crc_crcAxiStream_crcReqBuf_D_OUT[12],
	       crc_crcAxiStream_crcReqBuf_D_OUT[12],
	       crc_crcAxiStream_crcReqBuf_D_OUT[12:11],
	       crc_crcAxiStream_crcReqBuf_D_OUT[11],
	       crc_crcAxiStream_crcReqBuf_D_OUT[11],
	       crc_crcAxiStream_crcReqBuf_D_OUT[11],
	       crc_crcAxiStream_crcReqBuf_D_OUT[11],
	       crc_crcAxiStream_crcReqBuf_D_OUT[11],
	       crc_crcAxiStream_crcReqBuf_D_OUT[11],
	       crc_crcAxiStream_crcReqBuf_D_OUT[11:10],
	       crc_crcAxiStream_crcReqBuf_D_OUT[10],
	       crc_crcAxiStream_crcReqBuf_D_OUT[10],
	       crc_crcAxiStream_crcReqBuf_D_OUT[10],
	       crc_crcAxiStream_crcReqBuf_D_OUT[10],
	       crc_crcAxiStream_crcReqBuf_D_OUT[10],
	       crc_crcAxiStream_crcReqBuf_D_OUT[10],
	       crc_crcAxiStream_crcReqBuf_D_OUT[10:9],
	       crc_crcAxiStream_crcReqBuf_D_OUT[9],
	       crc_crcAxiStream_crcReqBuf_D_OUT[9],
	       crc_crcAxiStream_crcReqBuf_D_OUT[9],
	       crc_crcAxiStream_crcReqBuf_D_OUT[9],
	       crc_crcAxiStream_crcReqBuf_D_OUT[9],
	       crc_crcAxiStream_crcReqBuf_D_OUT[9],
	       crc_crcAxiStream_crcReqBuf_D_OUT[9:8],
	       crc_crcAxiStream_crcReqBuf_D_OUT[8],
	       crc_crcAxiStream_crcReqBuf_D_OUT[8],
	       crc_crcAxiStream_crcReqBuf_D_OUT[8],
	       crc_crcAxiStream_crcReqBuf_D_OUT[8],
	       crc_crcAxiStream_crcReqBuf_D_OUT[8],
	       crc_crcAxiStream_crcReqBuf_D_OUT[8],
	       crc_crcAxiStream_crcReqBuf_D_OUT[8:7],
	       crc_crcAxiStream_crcReqBuf_D_OUT[7],
	       crc_crcAxiStream_crcReqBuf_D_OUT[7],
	       crc_crcAxiStream_crcReqBuf_D_OUT[7],
	       crc_crcAxiStream_crcReqBuf_D_OUT[7],
	       crc_crcAxiStream_crcReqBuf_D_OUT[7],
	       crc_crcAxiStream_crcReqBuf_D_OUT[7],
	       crc_crcAxiStream_crcReqBuf_D_OUT[7:6],
	       crc_crcAxiStream_crcReqBuf_D_OUT[6],
	       crc_crcAxiStream_crcReqBuf_D_OUT[6],
	       crc_crcAxiStream_crcReqBuf_D_OUT[6],
	       crc_crcAxiStream_crcReqBuf_D_OUT[6],
	       crc_crcAxiStream_crcReqBuf_D_OUT[6],
	       crc_crcAxiStream_crcReqBuf_D_OUT[6],
	       crc_crcAxiStream_crcReqBuf_D_OUT[6:5],
	       crc_crcAxiStream_crcReqBuf_D_OUT[5],
	       crc_crcAxiStream_crcReqBuf_D_OUT[5],
	       crc_crcAxiStream_crcReqBuf_D_OUT[5],
	       crc_crcAxiStream_crcReqBuf_D_OUT[5],
	       crc_crcAxiStream_crcReqBuf_D_OUT[5],
	       crc_crcAxiStream_crcReqBuf_D_OUT[5],
	       crc_crcAxiStream_crcReqBuf_D_OUT[5:4],
	       crc_crcAxiStream_crcReqBuf_D_OUT[4],
	       crc_crcAxiStream_crcReqBuf_D_OUT[4],
	       crc_crcAxiStream_crcReqBuf_D_OUT[4],
	       crc_crcAxiStream_crcReqBuf_D_OUT[4],
	       crc_crcAxiStream_crcReqBuf_D_OUT[4],
	       crc_crcAxiStream_crcReqBuf_D_OUT[4],
	       crc_crcAxiStream_crcReqBuf_D_OUT[4:3],
	       crc_crcAxiStream_crcReqBuf_D_OUT[3],
	       crc_crcAxiStream_crcReqBuf_D_OUT[3],
	       crc_crcAxiStream_crcReqBuf_D_OUT[3],
	       crc_crcAxiStream_crcReqBuf_D_OUT[3],
	       crc_crcAxiStream_crcReqBuf_D_OUT[3],
	       crc_crcAxiStream_crcReqBuf_D_OUT[3],
	       crc_crcAxiStream_crcReqBuf_D_OUT[3:2],
	       crc_crcAxiStream_crcReqBuf_D_OUT[2],
	       crc_crcAxiStream_crcReqBuf_D_OUT[2],
	       crc_crcAxiStream_crcReqBuf_D_OUT[2],
	       crc_crcAxiStream_crcReqBuf_D_OUT[2],
	       crc_crcAxiStream_crcReqBuf_D_OUT[2],
	       crc_crcAxiStream_crcReqBuf_D_OUT[2],
	       IF_crc_crcAxiStream_crcReqBufD_OUT_BIT_2_THEN_ETC__q69[0] } &
	     crc_crcAxiStream_crcReqBuf_D_OUT[289:34] ;
  assign crc_crcAxiStream_crcRespFifoOut_readInterCrcTa_ETC___d1132 =
	     interCrc__h287463 ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[31:0] ;
  assign ctrlSig_shiftAmt__h59003 =
	     crc_crcAxiStream_crcReqBuf_D_OUT[33] ?
	       6'd0 :
	       (crc_crcAxiStream_crcReqBuf_D_OUT[32] ?
		  6'd1 :
		  (crc_crcAxiStream_crcReqBuf_D_OUT[31] ?
		     6'd2 :
		     (crc_crcAxiStream_crcReqBuf_D_OUT[30] ?
			6'd3 :
			(crc_crcAxiStream_crcReqBuf_D_OUT[29] ?
			   6'd4 :
			   (crc_crcAxiStream_crcReqBuf_D_OUT[28] ?
			      6'd5 :
			      (crc_crcAxiStream_crcReqBuf_D_OUT[27] ?
				 6'd6 :
				 (crc_crcAxiStream_crcReqBuf_D_OUT[26] ?
				    6'd7 :
				    (crc_crcAxiStream_crcReqBuf_D_OUT[25] ?
				       6'd8 :
				       (crc_crcAxiStream_crcReqBuf_D_OUT[24] ?
					  6'd9 :
					  (crc_crcAxiStream_crcReqBuf_D_OUT[23] ?
					     6'd10 :
					     (crc_crcAxiStream_crcReqBuf_D_OUT[22] ?
						6'd11 :
						(crc_crcAxiStream_crcReqBuf_D_OUT[21] ?
						   6'd12 :
						   (crc_crcAxiStream_crcReqBuf_D_OUT[20] ?
						      6'd13 :
						      (crc_crcAxiStream_crcReqBuf_D_OUT[19] ?
							 6'd14 :
							 (crc_crcAxiStream_crcReqBuf_D_OUT[18] ?
							    6'd15 :
							    (crc_crcAxiStream_crcReqBuf_D_OUT[17] ?
							       6'd16 :
							       (crc_crcAxiStream_crcReqBuf_D_OUT[16] ?
								  6'd17 :
								  (crc_crcAxiStream_crcReqBuf_D_OUT[15] ?
								     6'd18 :
								     (crc_crcAxiStream_crcReqBuf_D_OUT[14] ?
									6'd19 :
									(crc_crcAxiStream_crcReqBuf_D_OUT[13] ?
									   6'd20 :
									   (crc_crcAxiStream_crcReqBuf_D_OUT[12] ?
									      6'd21 :
									      (crc_crcAxiStream_crcReqBuf_D_OUT[11] ?
										 6'd22 :
										 (crc_crcAxiStream_crcReqBuf_D_OUT[10] ?
										    6'd23 :
										    (crc_crcAxiStream_crcReqBuf_D_OUT[9] ?
										       6'd24 :
										       (crc_crcAxiStream_crcReqBuf_D_OUT[8] ?
											  6'd25 :
											  (crc_crcAxiStream_crcReqBuf_D_OUT[7] ?
											     6'd26 :
											     (crc_crcAxiStream_crcReqBuf_D_OUT[6] ?
												6'd27 :
												(crc_crcAxiStream_crcReqBuf_D_OUT[5] ?
												   6'd28 :
												   (crc_crcAxiStream_crcReqBuf_D_OUT[4] ?
												      6'd29 :
												      (crc_crcAxiStream_crcReqBuf_D_OUT[3] ?
													 6'd30 :
													 (crc_crcAxiStream_crcReqBuf_D_OUT[2] ?
													    6'd31 :
													    6'd32))))))))))))))))))))))))))))))) ;
  assign firstHalfRes__h159836 =
	     firstHalfRes__h159845 ^ secondHalfRes__h159846 ;
  assign firstHalfRes__h159845 =
	     firstHalfRes__h159854 ^ secondHalfRes__h159855 ;
  assign firstHalfRes__h159854 =
	     firstHalfRes__h159863 ^ secondHalfRes__h159864 ;
  assign firstHalfRes__h159863 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[39:8] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[71:40] ;
  assign firstHalfRes__h162198 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[167:136] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[199:168] ;
  assign firstHalfRes__h162982 =
	     firstHalfRes__h162991 ^ secondHalfRes__h162992 ;
  assign firstHalfRes__h162991 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[295:264] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[327:296] ;
  assign firstHalfRes__h164072 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[423:392] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[455:424] ;
  assign firstHalfRes__h164856 =
	     firstHalfRes__h164865 ^ secondHalfRes__h164866 ;
  assign firstHalfRes__h164865 =
	     firstHalfRes__h164874 ^ secondHalfRes__h164875 ;
  assign firstHalfRes__h164874 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[551:520] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[583:552] ;
  assign firstHalfRes__h166516 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[679:648] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[711:680] ;
  assign firstHalfRes__h167300 =
	     firstHalfRes__h167309 ^ secondHalfRes__h167310 ;
  assign firstHalfRes__h167309 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[807:776] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[839:808] ;
  assign firstHalfRes__h168390 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[935:904] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[967:936] ;
  assign firstHalfRes__h169316 =
	     crc_crcAxiStream_crcRespFifoOut_crcTabVec_32_lookupTable_lookupTable_D_OUT_2 ^
	     crc_crcAxiStream_crcRespFifoOut_crcTabVec_33_lookupTable_lookupTable_D_OUT_2 ;
  assign firstHalfRes__h287806 =
	     firstHalfRes__h287815 ^ secondHalfRes__h287816 ;
  assign firstHalfRes__h287815 =
	     firstHalfRes__h287824 ^ secondHalfRes__h287825 ;
  assign firstHalfRes__h287824 =
	     firstHalfRes__h287833 ^ secondHalfRes__h287834 ;
  assign firstHalfRes__h287833 =
	     firstHalfRes__h287842 ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[127:96] ;
  assign firstHalfRes__h287842 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[63:32] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[95:64] ;
  assign firstHalfRes__h290740 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[223:192] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[255:224] ;
  assign firstHalfRes__h291524 =
	     firstHalfRes__h291533 ^ secondHalfRes__h291534 ;
  assign firstHalfRes__h291533 =
	     firstHalfRes__h291542 ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[415:384] ;
  assign firstHalfRes__h291542 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[351:320] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[383:352] ;
  assign firstHalfRes__h293036 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[511:480] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[543:512] ;
  assign firstHalfRes__h293820 =
	     firstHalfRes__h293829 ^ secondHalfRes__h293830 ;
  assign firstHalfRes__h293829 =
	     firstHalfRes__h293838 ^ secondHalfRes__h293839 ;
  assign firstHalfRes__h293838 =
	     firstHalfRes__h293847 ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[703:672] ;
  assign firstHalfRes__h293847 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[639:608] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[671:640] ;
  assign firstHalfRes__h295968 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[799:768] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[831:800] ;
  assign firstHalfRes__h296752 =
	     firstHalfRes__h296761 ^ secondHalfRes__h296762 ;
  assign firstHalfRes__h296761 =
	     firstHalfRes__h296770 ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[991:960] ;
  assign firstHalfRes__h296770 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[927:896] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[959:928] ;
  assign firstHalfRes__h298264 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[1087:1056] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[1119:1088] ;
  assign interCrc__h169911 =
	     (shiftAmt__h169932 <= 7'd36) ?
	       { CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q33,
		 CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q34,
		 CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q35,
		 CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q36,
		 CASE_shiftAmt69932_0_0_1_crc_crcAxiStream_crcR_ETC__q37,
		 CASE_shiftAmt69932_0_0_1_0_2_crc_crcAxiStream__ETC__q38,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_crc_crcAxiStr_ETC__q39,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_crc_crcAx_ETC__q40,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_crc_c_ETC__q41,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_c_ETC__q42,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q43,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q44,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q45,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q46,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q47,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q48,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q49,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q50,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q51,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q52,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q53,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q54,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q55,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q56,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q57,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q58,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q59,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q60,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q61,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q62,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q63,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q64,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q65,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q66,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q67,
		 CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q68 } :
	       288'd0 ;
  assign interCrc__h287463 = firstHalfRes__h287806 ^ secondHalfRes__h287807 ;
  assign nextInterCrc__h169222 =
	     firstHalfRes__h169316 ^ secondHalfRes__h169317 ;
  assign nextInterCrc__h169223 =
	     nextInterCrc__h169222 ^
	     crc_crcAxiStream_crcRespFifoOut_reduceCrcResBuf_D_OUT[39:8] ;
  assign preProcessRes_data__h13182 =
	     { crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[0],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[1],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[2],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[3],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[4],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[5],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[6],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[7],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[8],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[9],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[10],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[11],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[12],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[13],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[14],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[15],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[16],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[17],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[18],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[19],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[20],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[21],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[22],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[23],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[24],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[25],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[26],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[27],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[28],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[29],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[30],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[31],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[32],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[33],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[34],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[35],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[36],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[37],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[38],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[39],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[40],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[41],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[42],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[43],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[44],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[45],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[46],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[47],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[48],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[49],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[50],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[51],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[52],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[53],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[54],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[55],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[56],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[57],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[58],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[59],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[60],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[61],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[62],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[63],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[64],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[65],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[66],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[67],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[68],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[69],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[70],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[71],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[72],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[73],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[74],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[75],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[76],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[77],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[78],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[79],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[80],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[81],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[82],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[83],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[84],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[85],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[86],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[87],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[88],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[89],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[90],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[91],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[92],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[93],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[94],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[95],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[96],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[97],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[98],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[99],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[100],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[101],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[102],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[103],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[104],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[105],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[106],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[107],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[108],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[109],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[110],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[111],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[112],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[113],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[114],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[115],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[116],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[117],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[118],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[119],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[120],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[121],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[122],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[123],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[124],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[125],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[126],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[127],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[128],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[129],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[130],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[131],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[132],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[133],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[134],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[135],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[136],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[137],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[138],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[139],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[140],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[141],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[142],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[143],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[144],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[145],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[146],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[147],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[148],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[149],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[150],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[151],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[152],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[153],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[154],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[155],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[156],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[157],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[158],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[159],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[160],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[161],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[162],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[163],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[164],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[165],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[166],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[167],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[168],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[169],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[170],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[171],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[172],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[173],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[174],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[175],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[176],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[177],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[178],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[179],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[180],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[181],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[182],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[183],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[184],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[185],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[186],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[187],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[188],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[189],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[190],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[191],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[192],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[193],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[194],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[195],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[196],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[197],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[198],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[199],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[200],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[201],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[202],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[203],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[204],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[205],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[206],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[207],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[208],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[209],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[210],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[211],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[212],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[213],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[214],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[215],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[216],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[217],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[218],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[219],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[220],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[221],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[222],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[223],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[224],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[225],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[226],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[227],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[228],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[229],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[230],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[231],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[232],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[233],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[234],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[235],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[236],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[237],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[238],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[239],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[240],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[241],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[242],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[243],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[244],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[245],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[246],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[247],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[248],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[249],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[250],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[251],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[252],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[253],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[254],
	       crc_crcAxiStream_crcReqBuf_first_BIT_33_CONCAT_ETC___d139[255] } ;
  assign secondHalfRes__h159837 =
	     firstHalfRes__h164856 ^ secondHalfRes__h164857 ;
  assign secondHalfRes__h159846 =
	     firstHalfRes__h162982 ^ secondHalfRes__h162983 ;
  assign secondHalfRes__h159855 =
	     firstHalfRes__h162198 ^ secondHalfRes__h162199 ;
  assign secondHalfRes__h159864 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[103:72] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[135:104] ;
  assign secondHalfRes__h162199 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[231:200] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[263:232] ;
  assign secondHalfRes__h162983 =
	     firstHalfRes__h164072 ^ secondHalfRes__h164073 ;
  assign secondHalfRes__h162992 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[359:328] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[391:360] ;
  assign secondHalfRes__h164073 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[487:456] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[519:488] ;
  assign secondHalfRes__h164857 =
	     firstHalfRes__h167300 ^ secondHalfRes__h167301 ;
  assign secondHalfRes__h164866 =
	     firstHalfRes__h166516 ^ secondHalfRes__h166517 ;
  assign secondHalfRes__h164875 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[615:584] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[647:616] ;
  assign secondHalfRes__h166517 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[743:712] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[775:744] ;
  assign secondHalfRes__h167301 =
	     firstHalfRes__h168390 ^ secondHalfRes__h168391 ;
  assign secondHalfRes__h167310 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[871:840] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[903:872] ;
  assign secondHalfRes__h168391 =
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[999:968] ^
	     crc_crcAxiStream_crcRespFifoOut_readCrcTabResBuf_D_OUT[1031:1000] ;
  assign secondHalfRes__h169317 =
	     crc_crcAxiStream_crcRespFifoOut_crcTabVec_34_lookupTable_lookupTable_D_OUT_2 ^
	     crc_crcAxiStream_crcRespFifoOut_crcTabVec_35_lookupTable_lookupTable_D_OUT_2 ;
  assign secondHalfRes__h287807 =
	     firstHalfRes__h293820 ^ secondHalfRes__h293821 ;
  assign secondHalfRes__h287816 =
	     firstHalfRes__h291524 ^ secondHalfRes__h291525 ;
  assign secondHalfRes__h287825 =
	     firstHalfRes__h290740 ^ secondHalfRes__h290741 ;
  assign secondHalfRes__h287834 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[159:128] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[191:160] ;
  assign secondHalfRes__h290741 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[287:256] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[319:288] ;
  assign secondHalfRes__h291525 =
	     firstHalfRes__h293036 ^ secondHalfRes__h293037 ;
  assign secondHalfRes__h291534 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[447:416] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[479:448] ;
  assign secondHalfRes__h293037 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[575:544] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[607:576] ;
  assign secondHalfRes__h293821 =
	     firstHalfRes__h296752 ^ secondHalfRes__h296753 ;
  assign secondHalfRes__h293830 =
	     firstHalfRes__h295968 ^ secondHalfRes__h295969 ;
  assign secondHalfRes__h293839 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[735:704] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[767:736] ;
  assign secondHalfRes__h295969 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[863:832] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[895:864] ;
  assign secondHalfRes__h296753 =
	     firstHalfRes__h298264 ^ secondHalfRes__h298265 ;
  assign secondHalfRes__h296762 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[1023:992] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[1055:1024] ;
  assign secondHalfRes__h298265 =
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[1151:1120] ^
	     crc_crcAxiStream_crcRespFifoOut_readInterCrcTabResBuf_D_OUT[1183:1152] ;
  assign shiftAmt__h169932 =
	     { 1'd0,
	       crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[5:0] } ;
  assign x_data__h64227 =
	     (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0] <=
	      6'd32) ?
	       { CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q1,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q2,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q3,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q4,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q5,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q6,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31,
		 CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 } :
	       256'd0 ;
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q1 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd1,
      6'd2,
      6'd3,
      6'd4,
      6'd5,
      6'd6,
      6'd7,
      6'd8,
      6'd9,
      6'd10,
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q1 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q1 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q2 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q2 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd2,
      6'd3,
      6'd4,
      6'd5,
      6'd6,
      6'd7,
      6'd8,
      6'd9,
      6'd10,
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q2 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q2 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q3 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q3 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q3 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd3,
      6'd4,
      6'd5,
      6'd6,
      6'd7,
      6'd8,
      6'd9,
      6'd10,
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q3 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q3 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q4 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q4 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q4 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q4 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd4,
      6'd5,
      6'd6,
      6'd7,
      6'd8,
      6'd9,
      6'd10,
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q4 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q4 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q5 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q5 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q5 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q5 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q5 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd5,
      6'd6,
      6'd7,
      6'd8,
      6'd9,
      6'd10,
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q5 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q5 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q6 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q6 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q6 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q6 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q6 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q6 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd6,
      6'd7,
      6'd8,
      6'd9,
      6'd10,
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q6 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q6 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd7,
      6'd8,
      6'd9,
      6'd10,
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q7 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd8,
      6'd9,
      6'd10,
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q8 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd9,
      6'd10,
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q9 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd10,
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q10 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd11,
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q11 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd12,
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q12 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd13,
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q13 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd14,
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q14 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd15,
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q15 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd16,
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q16 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd17,
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q17 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd18,
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q18 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd19,
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q19 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd20,
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q20 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd21,
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q21 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd22,
      6'd23,
      6'd24,
      6'd25,
      6'd26,
      6'd27,
      6'd28,
      6'd29,
      6'd30,
      6'd31,
      6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q22 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[87:80];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd22:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd23, 6'd24, 6'd25, 6'd26, 6'd27, 6'd28, 6'd29, 6'd30, 6'd31, 6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q23 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[79:72];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[87:80];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd22:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd23:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd24, 6'd25, 6'd26, 6'd27, 6'd28, 6'd29, 6'd30, 6'd31, 6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q24 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[71:64];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[79:72];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[87:80];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd22:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd23:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd24:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd25, 6'd26, 6'd27, 6'd28, 6'd29, 6'd30, 6'd31, 6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q25 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[63:56];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[71:64];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[79:72];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[87:80];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd22:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd23:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd24:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd25:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd26, 6'd27, 6'd28, 6'd29, 6'd30, 6'd31, 6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q26 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[55:48];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[63:56];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[71:64];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[79:72];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[87:80];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd22:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd23:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd24:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd25:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd26:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd27, 6'd28, 6'd29, 6'd30, 6'd31, 6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q27 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[47:40];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[55:48];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[63:56];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[71:64];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[79:72];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[87:80];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd22:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd23:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd24:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd25:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd26:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd27:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd28, 6'd29, 6'd30, 6'd31, 6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q28 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[39:32];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[47:40];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[55:48];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[63:56];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[71:64];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[79:72];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[87:80];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd22:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd23:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd24:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd25:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd26:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd27:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd28:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd29, 6'd30, 6'd31, 6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q29 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[31:24];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[39:32];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[47:40];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[55:48];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[63:56];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[71:64];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[79:72];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[87:80];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd22:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd23:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd24:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd25:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd26:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd27:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd28:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd29:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd30, 6'd31, 6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q30 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[23:16];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[31:24];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[39:32];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[47:40];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[55:48];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[63:56];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[71:64];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[79:72];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[87:80];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd22:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd23:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd24:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd25:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd26:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd27:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd28:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd29:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd30:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd31, 6'd32:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q31 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT)
  begin
    case (crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[5:0])
      6'd0:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[15:8];
      6'd1:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[23:16];
      6'd2:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[31:24];
      6'd3:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[39:32];
      6'd4:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[47:40];
      6'd5:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[55:48];
      6'd6:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[63:56];
      6'd7:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[71:64];
      6'd8:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[79:72];
      6'd9:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[87:80];
      6'd10:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[95:88];
      6'd11:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[103:96];
      6'd12:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[111:104];
      6'd13:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[119:112];
      6'd14:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[127:120];
      6'd15:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[135:128];
      6'd16:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[143:136];
      6'd17:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[151:144];
      6'd18:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[159:152];
      6'd19:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[167:160];
      6'd20:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[175:168];
      6'd21:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[183:176];
      6'd22:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[191:184];
      6'd23:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[199:192];
      6'd24:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[207:200];
      6'd25:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[215:208];
      6'd26:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[223:216];
      6'd27:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[231:224];
      6'd28:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[239:232];
      6'd29:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[247:240];
      6'd30:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[255:248];
      6'd31:
	  CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
	      crc_crcAxiStream_crcRespFifoOut_preProcessResBuf_D_OUT[263:256];
      6'd32: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 = 8'd0;
      default: CASE_crc_crcAxiStream_crcRespFifoOut_preProces_ETC__q32 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q33 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q33 = 8'd0;
      default: CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q33 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q34 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd1:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q34 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q34 = 8'd0;
      default: CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q34 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q35 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd1:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q35 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd2:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q35 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q35 = 8'd0;
      default: CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q35 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q36 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd1:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q36 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd2:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q36 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd3:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q36 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q36 = 8'd0;
      default: CASE_shiftAmt69932_0_crc_crcAxiStream_crcRespF_ETC__q36 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_crc_crcAxiStream_crcR_ETC__q37 = 8'd0;
      7'd1:
	  CASE_shiftAmt69932_0_0_1_crc_crcAxiStream_crcR_ETC__q37 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd2:
	  CASE_shiftAmt69932_0_0_1_crc_crcAxiStream_crcR_ETC__q37 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd3:
	  CASE_shiftAmt69932_0_0_1_crc_crcAxiStream_crcR_ETC__q37 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd4:
	  CASE_shiftAmt69932_0_0_1_crc_crcAxiStream_crcR_ETC__q37 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_crc_crcAxiStream_crcR_ETC__q37 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_crc_crcAxiStream__ETC__q38 = 8'd0;
      7'd2:
	  CASE_shiftAmt69932_0_0_1_0_2_crc_crcAxiStream__ETC__q38 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd3:
	  CASE_shiftAmt69932_0_0_1_0_2_crc_crcAxiStream__ETC__q38 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd4:
	  CASE_shiftAmt69932_0_0_1_0_2_crc_crcAxiStream__ETC__q38 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd5:
	  CASE_shiftAmt69932_0_0_1_0_2_crc_crcAxiStream__ETC__q38 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_crc_crcAxiStream__ETC__q38 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_crc_crcAxiStr_ETC__q39 = 8'd0;
      7'd3:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_crc_crcAxiStr_ETC__q39 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd4:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_crc_crcAxiStr_ETC__q39 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd5:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_crc_crcAxiStr_ETC__q39 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd6:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_crc_crcAxiStr_ETC__q39 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_crc_crcAxiStr_ETC__q39 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_crc_crcAx_ETC__q40 = 8'd0;
      7'd4:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_crc_crcAx_ETC__q40 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd5:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_crc_crcAx_ETC__q40 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd6:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_crc_crcAx_ETC__q40 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd7:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_crc_crcAx_ETC__q40 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_crc_crcAx_ETC__q40 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_crc_c_ETC__q41 = 8'd0;
      7'd5:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_crc_c_ETC__q41 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd6:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_crc_c_ETC__q41 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd7:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_crc_c_ETC__q41 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd8:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_crc_c_ETC__q41 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_crc_c_ETC__q41 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_c_ETC__q42 = 8'd0;
      7'd6:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_c_ETC__q42 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd7:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_c_ETC__q42 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd8:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_c_ETC__q42 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd9:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_c_ETC__q42 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_c_ETC__q42 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q43 = 8'd0;
      7'd7:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q43 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd8:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q43 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd9:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q43 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd10:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q43 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q43 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q44 = 8'd0;
      7'd8:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q44 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd9:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q44 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd10:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q44 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd11:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q44 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q44 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q45 = 8'd0;
      7'd9:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q45 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd10:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q45 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd11:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q45 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd12:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q45 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q45 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q46 = 8'd0;
      7'd10:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q46 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd11:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q46 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd12:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q46 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd13:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q46 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q46 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q47 = 8'd0;
      7'd11:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q47 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd12:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q47 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd13:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q47 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd14:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q47 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q47 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q48 = 8'd0;
      7'd12:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q48 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd13:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q48 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd14:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q48 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd15:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q48 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q48 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q49 = 8'd0;
      7'd13:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q49 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd14:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q49 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd15:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q49 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd16:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q49 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q49 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q50 = 8'd0;
      7'd14:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q50 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd15:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q50 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd16:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q50 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd17:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q50 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q50 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q51 = 8'd0;
      7'd15:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q51 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd16:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q51 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd17:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q51 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd18:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q51 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q51 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q52 = 8'd0;
      7'd16:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q52 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd17:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q52 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd18:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q52 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd19:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q52 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q52 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q53 = 8'd0;
      7'd17:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q53 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd18:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q53 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd19:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q53 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd20:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q53 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q53 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q54 = 8'd0;
      7'd18:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q54 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd19:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q54 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd20:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q54 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd21:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q54 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q54 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q55 = 8'd0;
      7'd19:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q55 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd20:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q55 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd21:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q55 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd22:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q55 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q55 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q56 = 8'd0;
      7'd20:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q56 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd21:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q56 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd22:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q56 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd23:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q56 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q56 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q57 = 8'd0;
      7'd21:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q57 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd22:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q57 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd23:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q57 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd24:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q57 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q57 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q58 = 8'd0;
      7'd22:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q58 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd23:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q58 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd24:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q58 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd25:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q58 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q58 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q59 = 8'd0;
      7'd23:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q59 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd24:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q59 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd25:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q59 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd26:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q59 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q59 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q60 = 8'd0;
      7'd24:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q60 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd25:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q60 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd26:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q60 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd27:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q60 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q60 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd29,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q61 = 8'd0;
      7'd25:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q61 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd26:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q61 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd27:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q61 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd28:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q61 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q61 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd30,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q62 = 8'd0;
      7'd26:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q62 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd27:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q62 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd28:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q62 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd29:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q62 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q62 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd31,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q63 = 8'd0;
      7'd27:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q63 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd28:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q63 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd29:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q63 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd30:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q63 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q63 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd32,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q64 = 8'd0;
      7'd28:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q64 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd29:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q64 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd30:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q64 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd31:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q64 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q64 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd33,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q65 = 8'd0;
      7'd29:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q65 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd30:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q65 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd31:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q65 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd32:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q65 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q65 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd34,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q66 = 8'd0;
      7'd30:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q66 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd31:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q66 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd32:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q66 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd33:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q66 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q66 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd35,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q67 = 8'd0;
      7'd31:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q67 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd32:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q67 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd33:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q67 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd34:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q67 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q67 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end
  always@(shiftAmt__h169932 or
	  crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT)
  begin
    case (shiftAmt__h169932)
      7'd0,
      7'd1,
      7'd2,
      7'd3,
      7'd4,
      7'd5,
      7'd6,
      7'd7,
      7'd8,
      7'd9,
      7'd10,
      7'd11,
      7'd12,
      7'd13,
      7'd14,
      7'd15,
      7'd16,
      7'd17,
      7'd18,
      7'd19,
      7'd20,
      7'd21,
      7'd22,
      7'd23,
      7'd24,
      7'd25,
      7'd26,
      7'd27,
      7'd28,
      7'd29,
      7'd30,
      7'd31,
      7'd36:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q68 = 8'd0;
      7'd32:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q68 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[15:8];
      7'd33:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q68 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[23:16];
      7'd34:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q68 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[31:24];
      7'd35:
	  CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q68 =
	      crc_crcAxiStream_crcRespFifoOut_accuCrcResBuf_D_OUT[39:32];
      default: CASE_shiftAmt69932_0_0_1_0_2_0_3_0_4_0_5_0_6_0_ETC__q68 =
		   8'b10101010 /* unspecified value */ ;
    endcase
  end

  // handling of inlined registers

  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        crc_crcAxiStream_crcRespFifoOut_interCrcRes <= `BSV_ASSIGNMENT_DELAY
	    32'hFFFFFFFF;
	crc_crcAxiStream_crcRespFifoOut_isFirstFlag <= `BSV_ASSIGNMENT_DELAY
	    1'd1;
      end
    else
      begin
        if (crc_crcAxiStream_crcRespFifoOut_interCrcRes_EN)
	  crc_crcAxiStream_crcRespFifoOut_interCrcRes <= `BSV_ASSIGNMENT_DELAY
	      crc_crcAxiStream_crcRespFifoOut_interCrcRes_D_IN;
	if (crc_crcAxiStream_crcRespFifoOut_isFirstFlag_EN)
	  crc_crcAxiStream_crcRespFifoOut_isFirstFlag <= `BSV_ASSIGNMENT_DELAY
	      crc_crcAxiStream_crcRespFifoOut_isFirstFlag_D_IN;
      end
  end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    crc_crcAxiStream_crcRespFifoOut_interCrcRes = 32'hAAAAAAAA;
    crc_crcAxiStream_crcRespFifoOut_isFirstFlag = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
endmodule  // mkCrcRawAxiStreamCustomSend


`ifdef  BSV_WARN_REGFILE_ADDR_RANGE
`else
`define BSV_WARN_REGFILE_ADDR_RANGE 0
`endif

`ifdef BSV_ASSIGNMENT_DELAY
`else
`define BSV_ASSIGNMENT_DELAY
`endif


// Multi-ported Lookup Table(ROM) -- initializable from a file.
module LookupTableLoadSend(
    CLK,
    ADDR_1, D_OUT_1,
    ADDR_2, D_OUT_2,
    ADDR_3, D_OUT_3,
    ADDR_4, D_OUT_4,
    ADDR_5, D_OUT_5
);
   parameter                   file = "";
   parameter                   addr_width = 1;
   parameter                   data_width = 1;
   parameter                   lo = 0;
   parameter                   hi = 1;
   parameter                   binary = 0;

   input CLK;

   input [addr_width - 1 : 0]  ADDR_1;
   output [data_width - 1 : 0] D_OUT_1;

   input [addr_width - 1 : 0]  ADDR_2;
   output [data_width - 1 : 0] D_OUT_2;

   input [addr_width - 1 : 0]  ADDR_3;
   output [data_width - 1 : 0] D_OUT_3;

   input [addr_width - 1 : 0]  ADDR_4;
   output [data_width - 1 : 0] D_OUT_4;

   input [addr_width - 1 : 0]  ADDR_5;
   output [data_width - 1 : 0] D_OUT_5;

   reg [data_width - 1 : 0]    arr[lo:hi];


   initial
     begin : init_rom_block
	if (binary)
           $readmemb(file, arr, lo, hi);
        else
           $readmemh(file, arr, lo, hi);
     end // initial begin

   assign D_OUT_1 = arr[ADDR_1];
   assign D_OUT_2 = arr[ADDR_2];
   assign D_OUT_3 = arr[ADDR_3];
   assign D_OUT_4 = arr[ADDR_4];
   assign D_OUT_5 = arr[ADDR_5];

endmodule
