`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kk6QOGARuCrtK8kxtvLewRDnP2y0lX8/vax5+XVdBM6F2koyeujy1orVf35VyXQDN6qen3foHDQ4
XLEYnTkbWw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FVV4fU6gWgJJqZLS+kQi0iENeMRNSz34w2syv2Te0541rlZC94IhkHhyY2tRqoSmeimAY/l6Er5q
UVkxANvR8DRctD7sTAqTvkxNsAwzFhACn9xUQ8/2zRoCANferYpZHpsMAml3Sn0bJI8TXTagmIDl
Y3vY79giVRkJ+XvihTg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
i9GiLkhLA42oyRhEFvJEHkRlvKieUcRabry06xv4HPNgtBFZbcwWIgZ0EnpBsd6+lHjJV2SMtJ28
+3ZTA5Dks0Jq0+hjQHunWlJlAPNzpKIgZ3YZehJaW6vLNeVyRaVBl60L7H+Y6ZQLjy0noQTqWbGT
uM2fkQdf/F/eg3yNALAxDRH1wHufH2JBp3QkIqkWjS4EnDfimPbKB7JRGAE2ryxuZEghVm95UPrm
1j6N5Nt/xC2w1VQbSGzpG+uggoJ6sN4eobfLzBO77u5Pdv4y3ezF0V4umvofiAxc+gJrMJ86gAFH
3jMr7/EiyxewNTe3lp+ivrJojVvrJ3hyDGcp6Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LfjTTzedznHN5bMzyZVOlLXfI5jIQZKUE4BXpOAUoOWn4J30tk1i68Vxqc7QbZhnP6SFgdCEh0F3
h+o/0cR6W6bcxZK1Nb/p0ODnDSw55jgGwevS3UShX0vm2zAHSYefA7y5frnjbOzFqF10xbjI3tjT
Ncxj70v2MzGxZrZks54=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f3cKiigd59k5rgd4tb0lRkloMU6taFXzm9bsiDEReJrtypI2nsiWWi7WHsYCR/47ZYKqSS0njzA0
Ci6vFXAOOWJxmZugxRmk2f7HB+4BTLFM0CQTTs9YCF1Hi7v2TjIBAJ3dT4PsaCBot5WQJ20p153s
VK0ABahSCkD1kJQfNAEv1E/H7oQRZGVXPRa/EeT2Cww7TkbdtVC9B3pw09jIIKv96COmpW50nMOb
jLT+uUaGJ9iculQoRCjjaRoP1AXVYDnS4FbtwkGNp8S9knLOv55RsQXCV5v+M4Qn3Jzr7yzvk2I9
3xKvXTIczHQU5Uo0iQYZExNXobmv6ekwY+zsFg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 211040)
`protect data_block
TlF5IiFWaRGnVlp8/K/DyqeM2L5qgnFxykT5KQeQUV6dy0zxdLkvKnSESf24Nn0GdKj5bNpypsxI
r2zyutG4NCmefTiD/78bPpCyiPdI78B2IQMwVNPy4cJh6NO8sLBw5kPL87yPdjcQNnW5E3LBowY8
P1FtpGT6NpnOK6iKskg7QDUvrKkBZeeSx68UcR0J7dgCuN7vrN6O8r2iK225jb8bfs4cxSi8m6Ro
4gF0FOvCYuD7zbajI1k4WiXGCulB4dFTxQ4vZLtUkb3PL15Zgbz+Mec7Oq1zEBg7qlJnLkfNLELo
NuGHsgInGQ2vn5BR4AM341s3p05IiySnvl9RZeirFuECR2c8oGkY56Mb3RVaqf+n/38MczbYZak4
SnTC6SwcBmi2aXN2uysW2ucYGSh+G/4DvBMCwU/fmw3su7u4CI4Ai16A8l3933mgDu5yyK3RYz1k
st+aTsMBrs+QYMqdnicIWI8CbeaJMqxa+eu9Se4OcW/c5VN91bHKS3JnqpJSAENMTYr1ESSEj/9B
o+yrqC3VvO/TmO53EWD8mnZBx1G45XnK2ryYA7+cf6zumrFGQgrcM8tfcPgpNrIaG7jsjLScKRRd
Dpg/iHIMGglVwbOVhjONMiw800GCE+nUY1/KmsYh+gqfpwqHX3lVkNFff4KqvehzjnszHPoGaf7x
Mjv0f7i86+0zUQ46suPM10Fd2CS+vaM5k5EAnDOjhMJUGYKUVNhPe4muqziMTeGYk9JC8vPgKtab
X7Qgdl8Q9nvPQpaI8Egy4MtQl22FlOGZZeiaRwjJ9v3m5ZsV482pSCW9w89Th4J1dOi52v0BQCFH
kcFsR9rgw08pyPwNVjE0dqsfyG1FjC5bHujLlkcieNI70+8XJRuoLqGzjOr2Hatpmuz0akOUAgtc
Aq/MD95D6oxmetflsEsgfWmaTKjRqDJVtD57qyPbCZmlZzTf9VHLm6NAe7/ktRo70L9U/RZZy8yi
a7k4wny095a6jd1zL91LbdVGPHwnTv7k7IXZGWCWG7zqADQm/Acj12/dvmmUzGeZYD6GmlEA5fHF
0dDFISXT6eETeUrNb+XBqowU3qEpHsLPNAxAnjzXdT2X/IKCHRHJ0fVqmutPzxUnrlcfxKX3bMS2
kVVaPEYZvKKjV6YbxjjOb22I3untOtrEsNxHIMSeLht7jwsK0NXoDZVCX2waROZ285/0OB/4Cv/Y
m6/7iVOPuL0ESyiSYoPuUpSolUDkanHSEwe7TGowZsYdRYgZoIJKVs5UUYRT/jwefdq7I+muFMsZ
rJdh6nZBWzuiIFF7xzv3tlfOSSpxXt4KI6VL6r3mEUNIj9Oc3KIol5mM8y0K4OTva9Ctqsn9stSe
nu9MqrsXTQlEiMcXEnUfqfWS1qsVaIS9p1NqP2cmidECTXxUbspY0wKHz+ngYL8Oc7m+ichES4TW
BcWwLzMnOBVvdLhr0vun8Nz4UItKyWXc14/09+Gcc+ngZ5wod1aspjjHKCKOUGUouk67ONC2CPzE
wbhbbCIhzOJFnnfZW0lmKVZsQFZu6XbeNKdSop2dfmrLKE9vsvrdcGDKTbY8U8Yiw7OJn8cMEfbX
CISsgjTF6DcYpo2g4FfTFaU9U60I8TwzgbFSdEpHLe9+gniKvoFKSco3814lpnGgJjw1LyEC+JPY
N+NX+wgKsMMnsP2v3f3Kx3v/ISelcIquZAP27pCvaSu1LAYmNdwZO77I5i7QehTEqi711Gv4cDK4
L9gmcqf26Orn9zMkrRS6Md0jCMhugdiaxlv8diU1aCAX6uJqcQVE8Xu3m/QrLyJ1sA8R/6qkzPyg
QXR/wjXmw36GjdpTSbiU+iWwzPriTwl/DpIpaGsD/mlmK40IHdZjnq250E9LgwCljHDRVu8UkW80
XesjsftFSwbiaXUGNjYwyrKgg8XQ8SHC4wfTKSXBDJUjrf6XGNVIBcc6Ug+0BIRAX22hGT8Uq+Mv
0FlKRrzGWa8pgk719xZ5+vTjxhZECd78zW6/NTDpl2iF4p9rvkvV7RKxuiljc/NQMwzwG9AJvEfx
8t4XHF2rXORotLbNixvctoxUCCsfA1gCl/8ct3ig22LnrrDywi/0dFifnk24HFqldqf0hCUHUa7c
SwQZI+yHYPNRRBMITU0IwP5Kx+94lzF/0Scy8zXVQOz37RthYy/e7Ny5yxxqbn8jEEbWZT5G9ZRX
ItfrBvY//ZEvUGdu4f8FBDku8TRMA019Av3zrUp98sKD9KCbR0ako1D/RQiWsIQ5J+yhdb4MIySb
mvR11p33la3e9k0mFFOjLMpbuCMn2tWx2nJL6ByWag7fkuFv7nrjccoLFhP2B0hUDWajoUbuvLJ+
BDlTGWNrvBWj6VM5fTgU/SF5hk7BcG9LCI2GA3+RbtE9+SLzGdrXRoYUeE4Bxyot9FwLjRlQ8wQV
O83LeCKwBaNq0oftlEtxr2g7La6OUpUTsL7/Sw2+C/PY4ySTq+UXC62IZCA0zbxP+cv6X1Z5NSeZ
tdbn3oRvPlMctobL9O3SUmIFDi4gn62W3+GQlvKMkoR8SO97JN4GLfzBlTo4AE7UBr1qd4A0PXTi
3hOCjXXGTqvZbTtK+N/b4951ScwDeM/H6PSCJJiY7E/Wmu0dC5LArMYyS9Zyt8yL8FlG83S6V565
xK4QtQiUELTJ9FSSTAPFU9yLfURGedY8WBf8WOrBtGWzCoPlc5NcrNW+dvaaYbBjMl4e/G2EmIcA
7u8Mge7uOIHCjWdH75vCj5gKXr0gHaDC/jqAhydT9wPVhC6PAAqm7zQJH9yPa5gQbYRENTO7W+kR
EZE+TGDdu6DL7DQf5S2PWrNwxcDAtjj6Yy2+3FRROKLjhdBfVGY3bD+NAk1ct/MtMoSG3PECGuXE
a+159I7oQ9n2nbg1EjYR21ohyO99SbyKDM/30iYipAwP4oqQthlbD6/Knn9hU9lgy+dg3St9v1Hj
cI1KIbqoNuRTeG3qAUZ5T1KNgoOxMcaWnP3O/ElLpmv6FtzreR2gUmkQbn/MCOra76KYY2H5Sv7M
WmV5Hti+aVYG6JpmMj940NzXC/1ADz5Ygiy8TvoeYpxcM5pCU5zNxJ0+80/kOI9pt15Nk1yahdMW
ptlQ3Z6JXSSKhgtQRQxH+Ej0zXxIsPFPkHO/zoAv0s00w3uMbvOZR44C3NsQfDzP6woAali8FIl7
kQ/fcnrrt9XuuLDO0+ggb2SH7Il4hDFjnTa9oj20hh7PM68eygS+PLwFFKmc/ycfFUna3pMUE+F7
l4IQmPgAvHai5FqdA03PJK5etcr+l9U4WwAftyCB84TR3S6ot+knWZ1CGPDT5Nw1j13Dvs6xhB7j
QUGPmWKTcyQUgMehgwZZvC2J8xZSa43+Eqg2aW/EHENul0ocpS6M3AEXUsyxHGtuSrGBKB+mNzXc
GRyMdwFLvl/rKbovJ0GuxzpgVv80fOQjgI/i/rS5cotZQj+0qTCqbT0xsxsEWvg0kiqoWNgzY7Hd
EEzutsOoi2IepVSh5ZVUhSFSNFODJ6A1WcVnzzdo1XhswSXsFx63CBn5c5LuTm/njaVYR9v4hNT9
UiIjwJTvHtX3SFag9kXlTPEkflj3Sm1PQuJoeKgA44uW/cZP5BL49oRagxDWZgdwb/eZDvJEObb4
K4Zka6/6wh9yTFadA6JIXYk9CZ+jWqeBiUWngXFUCmFKRovxOV36qqrVHBcsB+TRHhIZvMefsTJo
qJIGvo9R/hP9sVlGuiD59aKkjzQfDNxfIZp7mivlFj4rXoS277B583FxO+ouBvRzfwW2cdBKEdTf
3g5932DVdaFPeJ78v3PFDJ4AxKf1mZ306acc1VjdvYM+zdZ4GrfIRaTZtqLIKi+/sPv3dxfKA/FA
rrRV5fCIY2H57QC2XcsW/0CG8fKMBW4bGAhrgKxxeOVu0/UFWrQtFDm3oLI3Yq6uf577HqXOmufK
lUsv4VFGIqRTI5ifVsZhANy1iauxe7ov8d8vxdfa047/iivHs463R913Fycrfg3szgV2t9n+b5tn
mYSQWui1YZNj89QLjZCUp0lLs8pweAsx4Z7vVu2kxTyvhdnNJAtWqWakudn1Rk58H1GGyps/74Jw
ZAX5GblGBRpjSL9CmQp2LomQSu/QGXrLS1uN6S8nKB7b0ojYKyxurpjcKYo+yrRBVIZZ5qglParP
o5CixDwT1gw0VTQu6COqNGgrB88p5EkYTiRhHo8aGZBdoeW5lauk4OqgBoxutMt6LDdht5IYs7cg
weEgNw8nyhY6CV5XXVXYw+2LQUwfnjeqVDcYgO35IH/N1U7N7fD45uMOMIAcrHfHiFw844lPYGVR
5NawtYZ6kicm5JFf2BBfhEiDhUvbDzRdN7JqjJ+V2ynm2EExjFlE6wUNmqyp7hQEYhxjevJ62Zm9
mOBWAxsct3l1d+rFgcZpBlaQBuuIZZay2RIVoDdfv3q1b8wHLf75R3Bc2gOR+OaPOO2gcfP1atPg
KWTginzLjaZC1up0HaJ9iP3UNSRsGVq98FVMtPyQkxCMzqOCzxE5aWei5i/4WZPfgPMvT6tqJf3v
i4eR1IwmzZIot4pRKSNKe4Bd/o99bVBGWRm2G7LLi40g0Dr6sLJbxZg2um+uCgPKd2ACqZNX6Xlg
6Yfgw7Jb8A6RKjeZktBD2Ix2uc4Sjn7Kk4FtaQvagYEDy/ktZ2ElApnKtgaEHO8N7SL1tMDJF0vh
lq1f2nJGFxI9AaoZKYb92rW3oKO9/SlDK6NFHCWyMiBkJpmz6F8Q9TQ8Z1ru0jDZoApMPBRd2LuK
r9GiF8okBqwvMdQWkqgHIQsCPzQXkzs+7X6JFDPw9EXnKsLnWq7YtmDKheOPle9tulQwqkuBJuSY
jdcnMwrjRKVkDIpX64ECuZR36DIw/DETLTMZ/wln0RQpkTmJZ/xc7OAXdcy745bYiM7f0G3w3MGu
7TLDg0xFIJdE4wwbTVIKGnuTuggmiNojS8fr3M8KrMzMIPoZ/7ODedK3pxjw3DJ6Cg+RVTFPgGZ0
pjI0JyIsMZj4i1dKcCrHPujS7Bc5ffwQYcW/N6haY5UbXE25LpzuEgDZst84FPSHzEAGWNr7KjD0
+4OKJRs077vSXkoEk83rp27FdJONg/oVxLHGtY8X+1v30AzX5bnJapS4xq7L0eJ1W8wg0d8dVw9N
3drN2qJ6eMvuXzGzBObACLnvDzLynUD4Q4JAlxSmvE9BAToLh1BH3PWa3182oub31e8A5jQwa1v8
ftB8tPiBWxvAS0od3ONgAzBBYTSP3N25DlGKJAgU9IMg7WdysZ63KqWX0t1AcsuvBpV4stNUX4XL
TVGh3dm69AHqO1VuQHn//EeJLSfdxrL85TZyZ1D+nrNJjDqBja11kRLPNVVGFKrCAyle1dz9op9X
e5/qdv79VJzlhn5NAKDBC8fLN961RmJRgA9KtASsaq0iwP1uuGW1lsfPpXFivrZEluVN1vzPa9R4
/op8i69Scpj3zTq6b6E/g3GMfkIFXO+S3CwonAFl6OCelcyr9aZddsjCrqxT0LlYDxJREb+n/1kL
crwkDVvZGvGmr8wrqLK7t0BrAak86imu8b4rHCY3ei+VZ1m/VSkZGXM08yl82rx4N16mqGPv6r31
rzqIhQStul1v7pD39n+RP0BPjOZQQvAV8BngJmY/57LcXhSvhoa39NJb/dlywRA0dUFRCJmi7I8s
1+GKTH0TRk07yJvoSLhXBNoREabSAAykb4/J08Vic0v7oTu2XyI58jx86ycZ4BE2cARZVZ8JxoHd
vBZrzqz3mFUJRqzI7R0SB59dMoA0v2kHZZlLYariviiRPppcpPkQqRRymHOp3QzG30FHfKEO1yYw
yEfXY1KlSkvTn6mati3xq+S5IS2Av0kv2cMCNX7p2WB28vWKBYCMGCuo+11GdhmRUYXwPbG2pB/w
XaWyGBu22kRXJKY25ngPW/9veSViCjF4+VPGRnsOzti+YQQiYjKMf/dY+ttwRW5cuXQSnOPdSwCr
95/0TgO6cG8Mp//+rB+yXJSAAWWU/IGExKzZ071D2xuO4lOxychQaSbKibch8FPpwFU15epznZhn
Y7fN0hriwh0lsBSPaLV7z92LKdz7Bso0bHO+f0d21qokaGpHMMcp4SD2zmxoaPxZmo684l2eIR67
EhcmFHsOtlxRkfw7vYCDHgi7usJnN12NRyq0c5JYJmUpJ/WhpnV8tHK87lD0ZZVmnAZtcIa+qEr8
hZZbBoHAo/N7AM0GoeSQvynhyQTeQLAyys0JEujrbYRVsV+iAzsYKzkNf18NsJ0kb3Z5n/hDwbFo
BnflTTx63oGF/jZcqAABBR0bYnxfmqNY2Hf90XIpwl/kex72KOuEQzBi1028j+cTH8HxSBCT4xLW
OgT3jBgq1FtmvhFtXAOxUTjakbRagf37n8vmAN1JCP/gRXM33AslIQoiIcqFbCFiUxMTXNqHfs8O
fUlOjpdbAktg9HmYF931e+4XfgIULvpO495yd+w4wI6nNoDE5YKf8AVSQxt0S8J2Zx0nuMvsUJrC
HRBm1h+xi0tFMRgPf5NoAX/wL3c75Hz8TWKR4HfOgFDnlDdQOyGTdVcAio8yJTnb4Ih+A9Pap+OQ
7DPBAX5F4IvGX2TxpVIlUNCpoIy9KJT41D3H54gEt2zmCNpji/Rfw64iiXo1hR+52YGUPnlJIWlj
4f5M0cuN1R6162eN6agl9AIE3DnDi7dBjfqWNn+/9AsOEeJWcNwSzXshUiwTsIfwybeDLdSjM6Xc
hC6Sycr/ve4zuhQ4ZMd/SpLwy8yo5PVpPmIx7sQRgusnQAVwl8Jo7lutTavX3JTqQYTJ0/HX0XuF
08m/KNYaSLGzIXfcFDGGOZ/hPTdSLOHcmbdcHY3JCEeRGL3bW65iLh9lLsk7oGvczIBEtd2T49KG
VwcO+D4PNUuikAFEC5By+SyIN8nNG8e/IOr38coUbUL9aMgOYMAC868SwoE6ouaa9hfC84dXySvF
ccoizmCERzm43la74RRfW5z6BtsjkoEMIlR1Qozcn6aSpthtQVi0y/wEhYCUMiqOK92mo+GtD1KZ
Ts+Jo+PE1Zj7yIGQDAzEbtzNoB4jF5c2T+3b0I3MROoKSeWlu7GvQ4XV+XMMF4SujdiiklGDI9j9
6OKHRxLTL/NIgjgQpUABdrSoN+0g2yGii9S7/g0QLDgKISKF0U8vCEgsKgYH93EHfT8MBygv1YQd
xZpV1+pwxKmc1723dBSeT2aQPbzw2UIelKB74H5mOBdKg08pGihxPFvOfhhjbn7+Fc77OrRVme5A
4JB+GdnCe8nD260xKi+EPwOqfH/dL2AHBYIb++atWSXpreaA3qj3M+joDIWUwz/fhd3iOt2Dr+tL
02msUZP2KhkrrJ0Rn/2M+sXPfcuYZhecmI6pTaQSyMu4qVVwQ4I4B9++ZgyMgeJQrKohkOTHEQ3e
iL05zcLPUaks90jJFqVxzc+XplMFBfcJlAZsOJIvRHAvDhQ5g5oyYGeNYZPFZyJBg9kkyDL3A/gy
+p/k6RnPZEsIVkid4XH1wF7CnHVsZNXTRpCmZXnojCfMUUA0Ooz+UgQ2xrpMSRertxpfXuZIrA/j
X8yU1HtFf/HI31oifk5M7z7RHiSpBMtQsyqNZZ8/Z0JQnwmTR8TbRPcCPmv8flVGhD1BIkYNlmQ0
/9QRT5CzqJyX4/P5997Pp5nYyHQ5i0IdGvO42l2bzqZgP0jrOzQ2StGjgKEt2o4+3CYnkLZaoExy
oCNnP5K+hQxcJtDUchLIe28Ji1plPrAYXEDetZCiOXFIoEkWGX6NERf48W0twivre+oAF41EZdVj
pEXxvNKTujrmqPQj+IKyrMgS8uOQwU3aFFXs8g2Gx9rIcu149TH5XkEn40Mx/hK2d18mg3uyF+IX
kNYhez6I85baJk+0jD4dgB203LozopH0k63fXZbU9+Ep+Ej1w7SO3D+msatGgzyPC0ibKcm9tuQZ
yEQQGBGY0JxltFEjAKxJeKx8X1vBxZuooYjg3jpKBb58EE2HuyWbvDpCFesGXA7BQVZ8PGAVESZ+
DUWzTXggcmiK9wIAc5wFEvKQ3rZjEh+v8o3AZIyf0bPneEIncK7feFxd49bY73gA7KJ6pBt/BRyg
p3hyPZo7xroF7woKHnDOEQ4ptI/MuVZQIlIoYXo/UOKQ2pCBmVHX/D54dZsk68sZTXdm6f0SvD5f
HtGZDc2nSnCn3w+OFr6OCGaZwF1EveVn2Sywxo7FxEGY+IgzIHp4e1H8De+KL+m6QraDGn3X8+ot
Q/4XQmCBMwwkm4SmlN5QzO54ijSfEwm9NO5qbM4bbt5PovaUJSBLHgncYaOwNEsZpKGS6Y3j877K
xMTHOxvA3Wy9T3vypWC+WPjWjEdVZ78rCQgoHXGefTjbjM2JBkqm9wUz4UQ+SmRfD5jAH5Qh812z
8DJ3cJJwC9pYvItENmJ2PT6N2pTfFLVo61MkEw+phW0aqRSjKlMqxbKuqgzgxooMrNQk9IFTIAzt
yOFK580xwWYdEB8PgM18gbkvdjb2DWugrXr0q5khig/fU2YTDn6HIa3DrtLzxxOChrRTefPrgBu+
Fxn4YtVdl4hQzFzYFh/ccoQ1EmiS1zyxu9XZTgZ8GJGhsRqYpxAjTfmwwNA9lnVM9AbDv/RhZIMf
ynl02XLX8m4yCjKtXWUScq0IVqHs7uV/jnKwlcKVRBYdIqI80yXp/OSB+UEwJnA+GF77/wCoGUYZ
UeapSxkCFLRAspqsf1TPlb0j91rWRHs95NPd2fkOr6dRp20l5/YIJIQGzS6ay2GaofrXS7LR3+6P
EODREzbIn8RVnOJ9UiDRbyaFRKUC7wHUUlsYTD7Op8q0N6CGQnOPm/RbfP55GLBifrLT0fslkQpw
kF6+mbFped7TCu7JHu5x3SAZhsYJjHoePQFBP+dhx8wt/OSIfCmLytkr26QIe4cn7PLLdaISl2QB
n86mDbQUfb9iony/oD19wtQBsWVauWyCPMiCyIAyCYVtdrWYRuAHgsxa5hnkVXu95WbnKIGTI5TW
3Y5K6yDDSEuIlPEqS6rW+Xa1p4u22GbOBWoIWr9QD7BtNBCZZYQ20yAxOhw2jF+lgPVrAehNWkyK
uNq+q8tmXDoNFXezTBdSdnfJUX++/SW41/ZRxrP7fe7493yXjBeCTZYvCnztBmqVdVDOezawa73k
Zu8Vxi+FtYEXGcJll/Za5PtRK4GycFGnyLy31m5sIr7V5NqpiNpK9/HFkDKaD1YDEofe1Y61Vtx3
u2pE0r5qqmK4j6DdtwZxZc34sDXp9RoJ7Mw36gvvKnwjhfSVJ1lQLU0uTQaTCL0ORDv103WaVav7
H7PqckU9/t2Nlg6GIzu7p7DGNDxjji5+pmkdbeMWdrdkHo21fptExgIs0+WFOq7TTui4xfdC+A/q
h+kXVGs606iq8mJ+84JERAQxaC+MMGuuQYPXqWlS0ZVz5w/fDDjphFY7VWkk5l2FxHS+1XrqHHg7
JYmswFGgv6mHsgPg60Eo2aYe5e27mZupLXO8ZP5/nohA4T4mDe4qnDAyl+aABksqDuAS0VyW9unq
+CYNa0ZyKvTKosoST0l+x2isZ117nkZ628RlGYnvXDS17TahfMS8fysm9zxPvKwqeZWiJH/Iu527
8ZatFdEPzWDPHukkTce71gQkpx3n2HFAFZi6uS1Q/AvfB2FcDDKUKvQ5jnusfLsy4JOAKG9/E6Nv
mVYVBYLz4kaepIeJRxc43RfduHwmoPDQnMFHC0G4ygpG0gG2cQJle3aBhFcvj8FCGv718Csgjbqz
BDICVfdr2FIKh18/7j0LY+tQyXNwwEryBtDIU0IX3e5jbFupkiz2dehoEiq4y/OUNfrLbTWI2Ukm
n6xXFHCDLFYd2lxsyhfSq1FeC5yniz+8IP0ZZ8KLgrMsJUbBpOzVauUlwKmHqO5ZXsYAzkgGFgNl
rLdgbCB60mTlBM1zHVx6AHzFq7wNJaMHtM9M+k+4kHQEUDvdqmvXLkFcymbwnnknOER9yYUA/JGz
lAINU/qmz9gNWDOEKxcj779rM4nwEFiieyXxoAiIEhTiRShwNq7svzmd3HrpHy14epf86h6PZKZY
s95LSxkIELn1wbrHm/Q0nowoJmdrq0JRFNIrH0CP3JF4Jft6ZHvtSIlhIg3fMG55V22mwplER0Li
cNffcV8TUNVn/E/oJwJ3T6I0WypChFIQskNz0xe4pK03tDNAqR8r1K2zfnMV62Lo2ugNUKQwMBSu
nkXYFkjH1iUDMYqWM+38iDgM7DycZKX6FuDDyMKzkUL6YVLi/yAGNT5e9LmCsbpccWzetKb3TU+L
sj89Yj4yzH8nyM88eNRgIeKbE+/6KITSNuf+JnUGUcPLQI07EK9nLPXLwv0+5fBK7FvyOZiu8Mkl
9SodvAPKMQ36wDneDWKnsDi7AawEjIFWWJVxlJy5OAxYchQzD4Dpd1NqxoUk08cHa3IVOIM+OEEf
S20xGg8NzjMcOKCCkoGaZdSqRKDgSzKWDWffvXNl+o1tWjvIzV5HlkFhlObQX4OefP7MH7Yi5V3X
5gPy0kPuDwRSjh61xfUgNpwI4Kda9oY2DOavwtX+24qMNFfnQ63WU48ZQI155FbQtwTpmfmYM5xH
7ql1QYJA1bWXJ323Y7Yt2SXIw1yQSdAdwwv6Lt0Kixf0UzUJHLV+J2fzsO6hucwbeGhWpYP9pmQf
+5cQQb/XfRBJO7BUEKSQCmyctv8irLi6jedeL5USsOz7IW2S+weleawwpD+SHzvRoi85fb2VkFc1
lUrOYkTv/H8XSWTQVkB6p+SHiBZjA1g8BzIh+lZryU15OKJGKjY66BOM1XogD15qJrSSiaWlvnXv
Fq6HMU9G91vTJDoa/1/S9fDHJ8CDM23H5EtsZD1GKuNfU5OEy9IHrINBo0G5TXdX9pOrandrdZNe
xXIBvjWSVFWBlocbupSXKMK280xoe6lkQSLvpZAnE9sMHbrA6AYxlJGDd9KL5/SfbwvGZ8BbOCx2
Mx2C4JSqwrylZoSCQLwnPoo3uvLqOX8m8pBoMC/zlU7l2WwnzyZIr/JV8VqMBsLOFgkmUPKIQODJ
q685wUA2mwY84yLysjAplhu1ccJaEnkUMQPo6i3JmrMXszlNxFgooXQ+TgDTHqBaDkyYu6H8TYsn
fqvUMcq/0JC7j74YaakZRfP5hY2DMUjqJu03CGTRAE3GaY5zdLciwX+zKB7Gmiu4xY1FVhuclQ6Z
Z4Mvw7hL+qRYwL3+aJ9+ttEWOHS4ruPUGe+R2+sSLFnJjEbOQB3oe0XREdFkcZEK/rhPKsStqyRL
HOFhLtSDeZNEwBWnZmYOYQmgFldcSIFjlHBKhyGGLBVJcSbXcl4W0KXDJXInwUsh+6hNMtBPLndV
NRUUYXwVdOKdeRi0uT5ke4AQwbhR16HrzaHTbO2cQuM//sn9p+kDxCww/OtpLKXDdBwYS+HR1Z6W
DDhWrOSCSVRsPmVOVD2ll9oAePxCB40HxbnPm801BVlrKY9RLlQIKT0n/9vf9621Tyo0jCSjxokn
0Bnl2xFHpmOl4g9nS1JiZlaFplT4Fanki7/JOZ1SX27ZuA3DGrbuP5/uZl93MLjVaYD7OuxBPn1N
wft0rcM3QuvfZlOPmJop1zgQ5U6bHk71sMEE++IDhJpqH8PrnQtWu7/VWdu0qDc+bOIrGRc6aEzJ
r8B9xcY6dLwtlnFjlHck9MOOV0Uy/zux2NWaKzeBTelOYvkMPuQZ3DSnFE26+NZUv1+xEw1aI+3H
27lvzu9E9lspwcYMCgUPNYHfV7ZnHdHZl0MWoyBzu92WmTKOW3OkUav1FujaWKRNxcQUhHyCozeT
sF4OjHyVE4bx/0CSt2+lKNwVNfr7vbztcUJfca81jS/TjYX8dUiUSsX2PrSUsz8wwLZjHgtl9JN6
oyuwlLTQlOA4KcuRsSPHe15WY4vMH0BP5jMCB7FlEf9DEcb7Dwr4Pm0D06UCPYd9fL1yJY/8jIB2
TWdRswBS+L0adOrDo8fn0wWuvmajhzpERW+6tBtAt/OUL/nKtcCU/3ZRJddluQ6YArLk45qiBelP
sgI6XdiukCw5wOHnYkWMtveSncKghRHZN6LB10hOi/EcdMi5aHAHuRH+CmET7cpzDHI8xSBnIKj0
uPldEjS1ZaSf7X5m//1oWBcKqDKhG0LCMuQB+cTLDtLQC6QWNvBPIhYtFy0T+zdpvoYAlScKW+lS
BP7VUS+6OeAWA+rFs3OP5DvAgs5Ui36SgnIyMzeAM88Q3hs1zhmJhHbjqrNwENKRHPGpzXcgL4kk
heuOBxvIu8/zA2lEw9pOzbayrt/Ycao2d0vYOjEfy1RqYWACkcakJOLv/m88MCfxFmNFt0y3AWZ5
RJnW+Ewt+JOnGB1naWiUVRHmFWxmZJxhZ0Ulq3ILuYu+GFLQftjipUSoQwEos3xmP8U/U3PO9VDd
fOYWCoxAmn8OFHo45T1exqOYsaPWelbQwGpu3ixdmr6UIDwpeOX2EzQbKfghhpdZx7y9WLR8+28x
TJgeZTzSa+bNb0BhvYi7iJiyrRO7yGtIhs27weClJrvnXSWYPPXVOcDuMNQA6XxCJcxwxmsy0HJz
YmjmBAjRVw5d7chuM8A2Ge6SuVIADbdYojWlUd33KtfA1zBEn2fmq5tqNxENPFHQv8U1CuWbmXpA
Sz+iI2NKH/RSs98Jc/NI9wixN6U4wZL1nV4rbXy6WVlzHbpuw8IJOiEbJ1uIPYDXMRR2WoLryKqF
hYKp5KfLBthbaCaZ2GVbXvmJj8O0Ux4IC6hxgElAcsZC27VUto8IEPQQmqVJp93SmQ4BKBwFg5K/
N81FSpsqqijzA1G+DIldqgWERzF8MD5P2avfyILjbojNSkRoV5lrqnVTWSWQhHit31lDc0ol5LtT
j5KuNrTdNYI5pzEFLLxX7AdpYUtW2aH/OnYGX19ibtDCmMlaMKWHs/nxYlArCNDj9P7vff9nUKmS
zCYfhw6YF62bObl/UXtyGew/DekhBuRtiIXfW1Xs2SV0bryTgrPwmdDTwBGAwnC6lxJxGuhUhmE9
1BmWiNqL2jIRnlaR21Zn8yevcWBQ+ebvMRSDAzq1DGlGKUcAtbqRBnsooqcvKXdKsrcJ79SBZVQr
9X1TDoCH9cUSaN8bI/Xx8nZ872gjNXyMoEaB9q4x0yNvxxCMsMFu1KwSFuxAuFm9vqEka1QKyi0q
dCUnEBKNmijg0IzOYOPF5SoayNzdBRwiswdxMJKimRvYOF9Ub4Ps4qN6GR8tEtqYoTw+sZ/FSclv
wqmTITRiGjv+YyyYtiSxaZhkPnoUGUysdDhZsa5WTp+HEdHgl0KbVWVxn3+cpFHJZTqwt4a0all8
Xh1xv9DWNq/bc7NosVXfYzFUYhE1+khIExD4hSTdg7KafhEhrcVTDE8ONT4t8clyRD0fEDwo+MLM
Ga3SLzzzLARm1oa38vJnG1iU40xmVmqcbI+AjTj61RhVpk19GGrHLmypWLkDRR88Z/8xV0pjz2wp
aKq/dzJW4hRG27QtlAEw1sbvytHDts8DGqkqWZS9qkoQbcl3bib1PgVgBKthnywU9SU17714JnR2
s38OSQPHLgMTLFdZ5EpWWSRjZDe8i0qeItYPg082Htg/HmqGuDbw+QdQRG0LdRcZz5q/9GvswTKc
hJzprfgpbwOsOJpM7xjkjOimpW8Zt7ktB5oNjKqP4l0ZzEC6uHLYzIJWbgWBO09pu10QtfD3TEMF
vT+Oy/HH5HuBy2WbyD2+FiZolWRr3ahgjE2vqpMi1CjdVlhth5VwzqN67pJPKhXvB/6zN96o/NWm
/raohfDZEc7dBkF8tCi23Mco8yB9IJDkwURqXCTxEiNbIS4zA5f+GRnRGMt3jAz6OD3WW6lrFZiJ
Z1iISELFx3GERUykK43LpcvpN5piDjdyeIvMLZQx1XQKv+317wY2MbTxLt/AJyV1Zle9GXdl8T0z
49ZGWqm/wvWp01uExJvpA39pxZUfisgo9luigQxQMfVahVQ2jWqwIx5Oc3mymgd0CelTZpBBObVq
6GMWPaHVedSJKJ9QIJBV8XyDaZywRnWt/6R2tr3fKxfv8Z2CUkXpfTA1WjcuhP1o7ZcsQZg9ALwK
OCu5jiVLcl4ooBDxwbR8rOJq1J7VDm4mK35PZQfriVeGDam37q3adolhf4PiXtwIygKjmoCon1OM
T75aoO6JXNVl7CsXhPxRe1ocpvl+F3OYOCUZ1S0oxJfetC986bj7oYOQIMIabLhGVLX6oap7RnQo
/qx27LBunzZtP27d5d27fTLqmg9vjLUx6s5dRAMySI6XCobmAPPYYbKQXhMGroTnlxOAh+s+u2+e
NcjOI9rTtu7PjVeWsnsI4Yd+U7IMdE+IDb41vNfCrYKpw91wEYXQj7tcqBmZLVY+DH9woKgVyCb+
9hAjA8pKSyRzb4GqjtqTs4XR3QrD9IQeNOPKM/FP/vzJ4wqNdUsAX956/E/WADSKXMYz5l/eq/46
fAudbQKVKIF7ExdHLe6GThLn3QlLjkgVC3epKj++ETlnkRTivPXd7uF7KSuEsi7c3anb2OXFJFxt
WvCE9ZnOhxxUUDRAntX2wEPALW6Z9dH8r/jQ8r+1dXpaEp7X5I415g17RpyK7KP5bRIjl9FNM96c
vYKaALjyDYICH9LHuEDIlT72JRxLoaMw8TsHgFAgBUmR1pt7+NGzB2yGzsgYRM/eqYTD6DSnPdDM
F9JeWktfcDwznLQlbcK6uQv81FaXvKkesril0Dkbbh3+SLkcKNPCnE7cca4we2IOLh0detYfZ6FZ
V/uNX/mqbVlZfeIUJ5TZt6+cqMsESB9L3Tn3MmDUHZPOfcMwa5nPBSXwNYiajeQVlQAsTKzb58LP
Dco3VT3ps29WDVQStUNhrOkF+vkYPDQlfe5x1YBhtwqqs+YaBPKUHuvROMTRMUSMmBA8PodpCwgy
JchNsx0Ga2+8IuMEhQ/mA6uQ+4pOGJqD9CU4cc0otcBpNzQi/FvrmawJC/9ySuWfDDHiIwc760vT
j0vbASzd7ajkOPeZnHVbT4waVAKOpRYMQFjdN/R5uqQ46MAPeBqTV7R9XVlDmTfNvkWOWQinHKYK
QZiBEko5TYpW1Iy8ndEqYexKcN1oBH9++DsVfoArP/TXl/13TzAO3BMUshUUb781sHRfT5vnADFC
HwJFxaqEAoroG6gbrVyd8ZHIvrCBD/6gzP87Uvx2NtXI5yPQu6EtQG2MgtCNfqr+i75XbNzez20z
20j1fZnKDq+QMf+1xZb4fx+/dZemGjX1/TnjXzf3rfuJMm1nW0f+F//0vJZgpQQq5cUWrH0Mhg+b
fFAoG0QvKMePxhOcL8IvbwaKRI7+XNS1CPX0M173T99D/4bcW/6v7d/84o6RuW3/rDI0ewMGl9DZ
80LPtRslxm9kO8PAsiGCSKLAcC+0skhKdPnF6liYeZ93WyeDV7WsTOBTJ2UXDyL8dQmVQ8LQXI1m
YT2cHxO0h8sv0VoLS+25RSQkEEtPerehjIZsa0+DFU7jlMU7XaVddHY7I6sTMOya4CDRB2VhFxPM
ZMT19AZEve3shIov2j83ddZRV9OwJdxIWXCpqcHHT09os5CB9zt+Vnf5SCfY5i9Xhz4q8hsb7Q5W
QfesAXb8nW5ioOJRw/ENyWlNrME7KI2NavdqJ2mIwnGHzv7WhiPbiEMPrBmi9csRv+dbY5613ROd
jJOyN84oVNvTL/SUjxroRnTC5Cd37qjTu0MKH6sLIFAr14Fca8/RzxuRAIKUo/7KRbnkH9wA2XC3
A3m4owgvrUmgAOTPoeahDGu57WEv++pst3i1/u4YpYFQwQEtUWurP0py2JaPVYkci4HhVoX+X2iX
o2JCrz2ce5aVlF8cnG89Kq/GMD0iznqZdREaBrK3UUpEe32gkaZ0kj2Qr5hZ0xeRUhi6m3S28bgP
ChjoZ4o1cIGW1QJaf+gG9I3qMoXjzurA5Sx8a1jqwt7fyANw2MIB7+pUnANvnvCDfQoutpCzgs+q
jq7JSIKfyV1GEycytgGUAm31ZWVPkvNjcgyMjmhXAJ+y+ZbFAd8wrmLcMuIe1Lvg7HcpezZUU82G
dHOwcSQVrv/KOr8bZKZi4b5W3ETH0CgS4LfdL11fYUWh9r/hiRS7dMylh6g4n3AUPGEwpXerkDOR
8NmcRLrouAbs8H7vgNZ1KeDH2AMMVT7CAqlKls8323KnUWTN2c8T509RZLly6rZO4aTPipYoSEC2
fikr9zczd85oJY6OARVSvlxccD37ERzIijmbUc4Fv8ma86sBSodkjWsfGJZfjGuyaPC1avkFxkh7
6RjFYnYLln+26xaXTvPwEtndxIPfP5kIKbgpiRjJTmS2YZvq3fTRvQtoAk9/R2fuQ2hu24hmdK5Y
KoXzODBrIzrXwEMkXfLIgl3zqr9UjIadsH+zTP3/ynlN8sXeBZwmmU0UNN798Y10/S2L89yKioRS
k3MDKmyQktp04bPgbFkTQoxFDi17kmxRuypxPE+rgXEvssawIRDUU5JwVnKxtPx2bPfURzePTVXt
KNetq2SGGJban6hOcPIWXqvQVXnzGychzsHMdnD9Srqa6XZVvwdsLMuKScAgKJlZ1DSr0JIrZ24/
x62dwN++8vJ29l4L3Poxrd0QHeRGZUjUl2+8kBn0emxOf6ABLr81Su6HI8/OQFbA+ACP0lyyYXT1
1v2+/FDzYL1pgScwFVqrZeUxAD0JlOyH96/IruKJRg6ADPXvbYNgTOfYqwiZ4ggOTlO8Slr+5n21
Ey5d2U3w7bGRDZUUTA55S6vMGrgaxO+3L6bJFhjUvFajf+vPFenOEzpGTpSUhAPPzuE/TXyDKpeS
X96X+l7ADJaYdhudWisZk38LzOcAThKpsyctNSM8hNJDfREjqpOx6A0gzfhULC3rZ8bgo6f5MBU0
t1/AEYTx9zMYpzuIkAKYqpsftyR9peyK9psa0Bzy3vwPj2vC+1jJsMJuHazoEkRN36mpc/yTfAz1
P9sXLOmzidP4jdePe6h2UYjwHuU/rBbII4JZlm680+IYMDfTXsDeATvO5qgXFjxv7TZa0yX/YZ1F
8UMlw+bJYLalko6zpcOfKb/cWw8AfrY0Hb25mf6qaAYkKCP1hDhN2nypVGH1pYoX2MscqjcyvsUH
SJswZL4TEip+lC+sv1NOAtecylerpZCa3mMk6XocHMi59C38pEDM8wwghBTTOh6yJy4nQhm4dsVN
h+SCFKq0zTrdmsBuOT3H2A+C8C7Reses0WXG3LB9HY6jDcyMyOShENVAcEOulhlX7cOpCB4s2Wdc
bsR8/Tm0r4rsGnC/TjhdpSdlRn2vstYVBF7Xk+KE2ErT+JKAkTjcs7m1FCWiLvTUaLGfjVMxS18z
/KLrDNRC/TQnhCH7H39SHVsi5f1tl29vJuqAoTQm0gDQJbA4NlA2lE61kh10QfuRJ7usmSVnAP/F
sZGaHHsuESJi4bax1Ws1NHSs4LvgZ6TEZIQOyE/Cil1ODt836jfvsrtKLZxWY+lCin7hW+4QrVBN
WixDnFpHKyBZz9WSFFQfvs1Gn1erC72TdrRY98J4EZuHzuz5Mvu65Uk5AgnPbSOTBXl2RP1pgRO6
u1ffubx9qlUfR4dVnHoT0Vg0+8aFxdwRN9WXe+vquaUx1XbqNAPdtlY2jMMJmdKd6nC3aMNn48NA
j4K2MdQrota+HIba108V1GuZz6dTaVjvLxOgRer2GGHIG+WD+FjQ5SbwqynCWzov2RcJp4ycWLxz
bMek5pTwve97+X+ZlGFXpfZORTcYzTYmrghIEW9U8sfcBMQ1p+DjSKoyWiGtCS8SJ3xFMRlDyYXx
LFd6/YWEQeYAwGtAHHiHCxDUtTU51ki0f3mFE9JeJJ9+sreADQFhZ44VKJ3JWmZH46flthtoNEjx
3xAQ4QBJqv8zm/4xIp2fswmMHUOlvWGrCC3rV2X9WcRzw91PP1U6TwdSS3i6ZJi5euzUvMqiVurK
TiDHcFHIRTusB9jGm3S5R+rwQLcFE/e152grc77udDloPBe8jhyOMVxwfXj+s0c5KHB19KAQx6pS
zSrK0OEtSnLVDFol5kO2JbtlufaoS6WH1AQg5tUP357boSFJTluFjm6+TaYxptblfR+jL50B4KfL
4B7ooZe2Idi7GOi9hdZ5VFcVXPoL81zv+IMIseXM5yR00mw+arEpMFZlpbZD/mmdHyXjS+2zwoN9
iZq1+8CFJkNBkmEf6Vb5S9W8YTAu0ePxlA58aZzgHqiJZipSqo9rlJg08X9Kku9MM2dfkZgcNiN1
ggI5QpVu96MOusTgxXuEvKhY+JCrMYA4+kfDrTzcwp3UuQJUtJsj7orJdhiowHJNmok4ox0MY5wd
8yDb7ffX6bKPKPe/yVzzDatOgnh+4nLQhuNGECiM0c285DtWipcUrNHhIefOxaksf0dSN4dQSCfJ
y3S3GdbuUss9zxA4TAA0jDxPSarWMDk0cU9tICphnPeaVo3/JSqqaz0lfh2dfGqBzfWBGs78bgaO
bGXyrvWMNrG6jVzmHA99WgfXxKw38mLhAIfe3Q7dBV3LzDEpQR3nB7DEr7VAaF025mmTcPANzWLH
H3AhCbHl5pXDZxNlaCc4tALW+hSyitNfSq5affJ7XuiqlAjP8xei+6UOUQpWCUNWOsnNvnN/J0/w
qknno97Jw8RFJKmGbkABtw68A6E5eLc0dFGJ046hguRg4hPbWWIzDihcuPUGipcfC6ppCKbhsWz1
fK+mNa5v1izibLeX1IfA1f+2Gs8o/8L0pcOT4MbhJi/lHXhbrbLNr9nXtHJV+Gsqmr6PfosmOsl7
WytzzYkzhxQdiToRv4PBzJulUMyG3ssg5XKr9r25yTpHWqMETE3/NpDnNDnfmzCGOOqf9D49Kuaa
faU74Sd3Hh5cNKVnKq+T8Y8CKoj8EiPuYzGDFZl4cQs7pkX1WWlji579BlUVs4bE78Q9kSp0eT7V
/S6QL8uV06073VTegj8JAJgrel9rzEVmWAKxQGISSeBBKzDwdSaWsP2fmBW4uVpNp4RRFdBtuVIc
1UOSzmDzlSLSZY+SuuTkAMmjpGhve9jdNfUPNxgSreF/7pn9U52Ru7i8LAk/kZfugNDqBsdRj5N1
PeMW2WE9fKYUDAwUirjZs0zvBqCqKzTrDemnP3higIbo6rf9sPFD2p91DH/Gg3giVtt8y59DZO7o
Cl9YRiAs53Y7wify6t7a0w7hYlU6FnkmQWOeDGBWLfoS7WIWNWPvTBqPcU8bujGrJ9zvjEUUL6qE
RbItTavv/rQTZp8eYCKEUFFZn1kgnvW63nu0mqWcwL7ptp8fYk6g/ZGUUx6y1A0mYd8tAhAmuLcB
cTlQlCSXe9AHo1gHiT/VQGvwi2OWdTAEhIGiQHvZ6EyZ5IydAjAYnNa7Ar1kr6pNPMaD4yTKfuqY
/pYbMlRHIedQnW5HiNf3HiDmubtyv3VU8Bti/lxagsNpnBmVccvEfPdx4As4J1fZZI6r24yXFcir
1oYt85UkDOIQB3BAMV1wF7AdUru+vYYCNirsbIWttEVjYFu3do6SM4NPBWw+iP6xHNL4jZn++Y3+
HgozLf+8RKyELbEEmoItKc/bscstWLn8Kpt9dX0oePULlablb34Tci0mni1Mj5L4nYubPSJJtKoE
p6tDWFiq2QjKQu5MaXPMRq6KbCdDYpovJleddFQANMLanxSee0f7eukp3v7wIEVI9rOXDhurizCK
/JOhO9a+AENS+21pCCsRhPiv4bNZLEu3wpUfgMnzHj2CZgbA+42/xslxkX7KxUcRxVLqZXgwtV0A
qXnbA52h6coprOyrDc7VoF3ttXYVmZ9zGsGw4PGIxh8HWukzEPFy0W2xqRSD6wkIyR4fWUytlH2s
z8JiCB0QeiPnljeggSDwxbTfPGkrctWhCWEP9see0U4prT1jyVvxcIJOb0TkZQX3pNejonORr16q
pHhUqUtYY3e6Ur9a7+zgnbkOYcG+6v6zVb4uxcQ17OwvqExBnzsN9q92NMCI2+zO0pe0A7X14p4v
WTOMlS+sEdS3KqA4IXbJaanadBYqtPhLJvj13qJOqkx/V/1pg+76x9kVlSvg5lLjZAQuCH/IBZ3F
7PoIKZYefnRZy+zxPcI3UtSXxtrum4j3s0d0wVlS/zr7+asvR0QXuxHA69VJmVQJYa9Q0mdGN3Ds
0ybbwJzMMRcF8TW1ETlBpL4wcc69Hj5mohdc3MmumXT0stuJjB1W+ApcVA/s/LeWUwxbS5vWgPuj
bIpBqhB7NLNPtPrbUY0Q0o9/i+BVyRpG6YiNjaETEvZKp7YSjaEgD9oD/wwNfZwFJtM0HIR6Xw/H
asdH7oI51p0fCNzK1/IB2M1S5j5GzJgleTE+3htZY5zKkLWtV6GqJmqT3Y5Wa5DTsKuLNuZac+q6
uS+4idVZ10724R9ur8BdLI6kwmcYJ0SBkkntClUwLFUh0MmUcQjxoENIrIXA7QVlfDrrmHWYxPtk
OylI9/Jdi8hk7C/kaSdk5aiHZxyg8hVC4F3XRdWElEc1c6RxicHoFD1Wl2D/r4a5wgxCKqBOp5Iu
aJHwFqPLilbMWWpRCeyxarH38oZb42EMMZZvda7FH4hsfnrjIfu2Veo+QX596e2RW1aEKNq5tyHa
6Qtjp/gbHa1rp0pMP28EP48SHIx54aWjqJcT+uhgYPOQ+2hI6eY/VRH4WMXck20xhtv5QJa1tanv
9QrZxeKizxZ7WhhoKKrIqqoVUN8+8+p0tgWuLwv20zIBWj5R1ONKqWChBY/Ra01qQ8V8gXIUkldN
3N85QuaRdWawxtrG4wrpFLfOjgk10L7JJbIyh0mQCIC93CCOv/BL427JlY30p4S+JG8PGOMFKSYx
ApR2MU7w6BK1JYugK0L9zAocMXx989MM4KWLcYUhZSQweJiZxz/X+mYfPuzbtX9W+fohiDjOyCiB
yYWa3wsaFSzpBF1wKjZk1HpYdf2LG+RleQ0ekNR3ETGuAdzeV7FrUf/HsI85fHQ4W7JQnusXF5kk
+0KmM3Yg9KrJlMD5XheZSFXQCO292FtHg0B8i1eiIFjq7gcNMQR+AdDF9v0+a0sqaUGVdhHwV9e9
k0oODEtofYqumoCxqGJbVRIgN7AeVQI2sR6Tak2SYuAPH2ZqVpJjpp5QHeGIx+oHM2aHCj1N+cJA
TqpdL/GEMfg++sSKZOtiycF2Mnlrihc7L00r4vU+SXuDI0hAA+rUfPC3oYMkMIJW4844bW/Yvlqh
j4/0uoKaydSuY0/QgW95SFODO7n+0o+3ePEzUwygZ8ls1dWMUitYTmpz2gS4NAccuY9JxMKrhGcT
iShGI42ZxF9ZY38qi5q9Kr+Wfsvu4fuXGZX3e5CmIYIQXfLpt2N+lYZ7jWf2M/6d3dOsKtCWTa+z
JyWoWrxkNBlxDd6qeDqhjqxn8gtjXp+1DSGWeTH+UdmTzfrgd7CJKjDwxd+7VDJyZigX4xj45FSA
bewrUNGtupWD1/1nvQjm/4DazEhR8pDLX60zuNWL9Z/254SvOIIai86vbUDbN64zM8JCdRSxg6dd
MGaHhz6jOp/1/bPDvvM4jPFgWZyZH/2LXedN4mPzYpEVxHigHa8FHpiIr0gwMOlg7dUcHwmOayU7
ufmiK2nQWEu+YZczLT5+99HQWizf/Jqvy0izj+K/hn+xTlt9jVvEAmYchwauWbDi5K+aDzMPEpI9
cS1XEE66s1JFRFIgDsa4NE/CkTPxhjuyjB/i06ihiUL+s9B3ry17DNYCa8VRcv+5HcKXzGEKfxem
Llt1ZOuYC7Fg63zXp61XZJzX/ZxIZYwgWzMVcVGTOiSgemmok/BY9lNj0rXPiZrHdF0QGFFvhjDc
XuvSXoAloKqDYLHfz5HwwDCBUev2tn02g1jT/Lq3u/yLFWV6/vB43fraPToMoluOYaBV6vCsOSXC
QdXglaEesminFZNDKWttbOOTjcDZxD+6fkJMwllJeUYB8YuU2wdLjuhDxjfJXvknyMVGsmPdBFFE
zuJqP4IOqv1SrCWMkZP6puqRrj6YZFvk2OpIYgm5siwdaoUpTiNp4BsY/IRF4++D+vs0NEUnf0Mn
SrhJQ8HTKis/tiI/xaNBH2iw+nmv9lKa3iP4IIMyeyOvZVELI2Bkk4f3C1TvScMK1xhTjzqz/NfQ
xJc3mkB0LhXLy79h1f6CmUKFTwZ+KBv/TyiZkjPORlGxaR4JPNFGhH8p/zqhKcVgUL9lD1xtVzw/
124gJAIM5osaIIgwVgYjJ7+C5awRAeE9oinNk3LsM2dicoTbz7TGqMdkfaco6i4EjALsEzxSOcYU
1KDZVQWV8TxOUsqpQMtMLdM+zemggdFTMQ3+IX7v7TQnouwGblGXiIIwN6Grec+YDI+Lwt2DNyU7
gUCkRDo3O7zVuTVN/lBnL6ed/rGhnJL3DgGH4MRfeUccqo1Jjj11RATj7ORVJsf2Epl+HZyTPHWz
fG/XswaAXg7hsxVL1dZbbviPHS3QGfbvnn+aPwDuB65g/rocR0QM6I1pAju1PDADtORNMhZOB2wW
jm7sikhNwLJcdon75FWPoCseqMnwUKzpcrMaVUuPyKuiEebGDXGPgneIjG1pQeYKmTmGc5S07IS6
HYfLcp8mvijPbtjVZFA4zTqsLXlm0Li0MetWPBzlkBlHCbIZ+ssqTNLFR2H1Cd6IYV6KuhWWD1bg
dC0mOMQD2aGNeMMAOsEURsXR/utelaJtvl4sVLLeWOzN77UIP4IUbPmWglow5m93OXdsXbBOjtwd
C4Tqs0JTJ/0JsNqZI4RoNDHIp1rQ7drrlXq7cCNdXghBvqA87s7FU+tfKudS90vjDkhv1aRg5zZJ
uBRXkboVXT8BCfejPaDESNNSKR+jBjvfj453mbAkp3aCMSir+d1xyhRGgqJPyfvPdLyxCzO7KBNh
5OecSDhLTOiGxty1/gkHB8rTQ4fozIhwSGtjnhEBs06XOgUotknp9ICc/klDfbTC42ylr6XWChLL
8puZZ94A4avYKAblp6UGta5UWMi+CpvtN/ROVGHLleGMMbBf7n20g8ISlRwV2TRvaIuvncfeVSnh
Et6Q+fugEI+rgCyyYNa/wfmKlmNa6/QSxPoV/eau8GQPgnAoa+KmfkZ71eHTUgcMqpwT9pCM0Y7E
flBRsVUc3ufy0FYekVJcvnvsoSA9xOS4kfHSVihD1zBUEmv5GDsr30vjcEelSstX78G3ax3cuIE9
0BalSBlNqQ7S/sfVNWn1j6TrqaEdZqMP8cJxvl263NjRJaAKp7HfJOLU0DsWtjcYYQvvlx7a50o5
1K4DZaRRIm7mHhe8q6am9zVR0hKgIZgeHPNk4PdFxlWCGflo2lR7faXyDqQDCdaj4JIdbln4LtJy
/R84ZfX/BSXtu03b+Gkv2PrtdXXSOZ5L/xog4PGQ1ULztE7N+xLaZaFiPHjxjKIpF93ZiUooQTdZ
5r1tg5JVVxdX5PNfRRx2fUCrqnGX/YpVdjAauuv3cfXurr4S1r1Dq2TvDL6nFy0evopXe3kA7xr3
z0qVc/0u/+gMd+PBBuARXRiI3eq656dSy36xBpR7tF7QsDkUowOKhkxW9uDrFqTv/1r2WnwGaq8/
4DTxLAu+OnEFY4ImMl41ky/S5DFrlMieXufsGZ3IR9dBp6b/XnzkNxiH9nv11Sz0RhGiMadXlX0G
dL03Pjh81gHNVhhrMvCF7jj4kXZqCq+lh9ApqSTp4WLoVVvl66cxqsDxLjpaiH/XPBuBqGOoX35D
Do6hnyP9oNioD0A8fxlpXpnZHdo97T5Ol64wTHGsuK/rq0Z3dMTRiPcidlcVpL1UgAbI0pbQOAgF
JiCkx0ejRFBJjSHHpz+pCT/5wmkfvMBhnpwSxfySSiAxGAWfesoZBmV1W4DGUasyyAFe+3Int5GL
k3PPjYXX+esffSe3Xn/YyVULdyW1ui7Jjgk4kuxhloWhnM91IOX33SG8hSPyKEmF+9bvoSC8vv/3
J4MLkWBWOEu0ua0hHmzTH8GblDC6Xsc2LdWXMriGqP87AK9f+/YvW3RX4ygmQ1WhKK2dIzm40G/r
X1fA8AXfYRi/+Ytl7XJKuBaexzVvz2FCRdM5AiHwb7QZiOOsu/RBixaXuSpKL7vcwxITL2jjgH+5
tMDzAxKNGOYW1stujobKCunDhVqy3mJzS/3Q2N7lDB5rWiR3IA/U0CrxRBTD5o2OB5TcD7/vIwFw
JzGeRjl6fTcUKglmS4Yk1LiaOtpdZ6ClmD0CYQZ7Svlwh5UZHmG7VjRhxgb1Z//J2OseoiLaca52
oGt8liq6m5jeBlV+6J0B2nnlcIHO8qA8lcgG30JF3Ej48N1Ri8VzB5FQ7Z6uRvl5mobeNEfoOTgQ
GfTejGQv4iztWeoC4qpddq7qsjH4U/RrSpa6RISR82kUpaH0OHPzH5oHuUTZY+UWNhGZPnTFX6qw
FvhWuEdUBTaTL/JKHH4kV+xMNZm8oQSvVbf63/kRBXbPCLOMaWRbZTACAQW68iw0B2qCpMNHiP2u
4s+pfIc2+9IQhXtnqK/wBdLVPaF9gzZcscVvMEdAf+ykH9EeyMEUITh3NlF18+JsNiYb58d6pAhI
a80mD7ISG7chPHPQfAEnkbgMJlMYVFcWqOsiCKMXSSD9TQA+twdgEF+y4floN2QBRpuzecvgFFS3
NNAbNUb4YtWSiP7kYkIqqfVov0R01psvd1EPcNXBX3EspIqk58ZwCF/km8KmJukfBe5sPrk/kRs3
OXmHHfH+ORK2mJZKvXqGSvIVT3NUCbFgJ7L2i6eHgsyqtkWHyht/btPVs30scvB77kZa7EjzFx4d
5LvDUOF8nNOVPAcfPpFDvRf4E9YpoC+lviNs7hL+vEKcNzB3ExjuQ8ZupObDq0h9B6R98o94DfX4
iv7TDTJq66tjSS0vQXmAN2goQZdANya2+TIzLbTOFnlR76u6QqNS2iK9OtmDppil1KNbLcBaQkjq
irgdZm+brMfM/FPeSt6wn2Z3XTNNdD6zXA6JRjkotNRvWjBgPGYUPrwlgpvM/YgHkrv+9WTES/hl
/OfYbfcaG4qY4o/2VBIVsEG7Y1K8iIEMsAdo0waPQAtRNbBfB+//NJ8d87kbRku4IsXeBGXTGEyH
DQuqBle8MWd2GmjQyVMslZnlPKU+0wJvn/+B8v0i84eqD105aTnID3iA1ERAolW3LoTS9WaHK9xp
QAzvqBFSqVymL68rIpsXmy9cbApS3k2mHy0tILp0wVnKj58/hotdctAv5yZWNkHOwwlJ2gDoLu0M
Xf7H9prLS4x+kEtI5Y/nWAs1yaauBHJEHwgZ2qSxaoItyTATiDAgrVyeCoA2UYK02YDIgp568jsJ
HFU8UK1a6wK+O5yr7r94u22VeLxUw+V1w8Wsk8sl5SJXVIXp/xbRm/rLyk6lADr2qV4IATF1CuuP
w4CZf3wBXUL9t9qTQ8L3N5j4CUkDSyJxbqkaRDG3Zyu4CH5jjEIqRHDcaMX+5grizyiUYK1VifSN
GIJTT8WRCMo2Auw97pVhAmXaGngCFpcu4V8PSkB6pSXIvKhYflJsQKoLZVgSsSEBjIVK+jiKPQF0
zXXKrFSJTKlvy8GBG47ovc0WIkAzn81KnRqIpwCoM3Iq7vo85AVz/oZ0nuCRAishbbTbmk3CrNoL
QboKZwjEul1skgF0tdXA+lcWn6Leqo5KRpRIXpHBFql/ZGMyY4POFgsmktr2CUIy3Ers7j0YpWyd
aWIl4HQ/E+Nu73Qd3DFQwi8eZHbyKPH/BTacy3owW5qMS6eixkccWIQGhHU+UNf4WiK9pDtThZqQ
Ve/rshqf0nNQErpgYmriC+DAU8ushjpIxaMlhbTwtINeKJoo8MS4Wiegb+1AebW/AYoM/izLvaRq
sUvHoyEhKL7geeJfWlsEYa2A25mRvfQN1rZ/f2I7TtqKGuGRxSxluokbyJlUoYickixTBq9b+Urk
vCUchTjRFYDEghtIofSnHkXlx+Lxow+aLZCP5vFM6MFrmsG1A+2Krrs4xNRGtMEEXNSlrkjdiMTd
qKqIVvJFuxajcJ0/JeNu7jwB4EQZoj7M6lJsm+PgngzTB1M9647byADFRR7YuwKQxx6pqt192sA5
Ci+Ff81wkfS9S7X8D3si+g/6vwQT0n8wRjubUa4qNWyK8MD6PBFnNXVeMJeF1P5J1Kfs3joEaBCK
v2af42mDvyTXbaaRkY3IiC6LrfWa/CkqXDT+u4e5oz+nuo9+Fel4jZbrsLtolBXGKXjG3F06LwQN
lkk97cbzKLreKrVfFoq6LHDc6CJnqAG/T8iBCQrLdygcUFxZHLq/qGnxS8XBHEuC23q30DUyP/VA
0g4e7QwDNvkHKZFi9Cstx5u3HtavX53KW+PiDiFmHJ/Ls8dpMsPzRyGUpmIb7RteZQsf2hrYzaAi
ND1eAb1JyBQrQUIrS6OVmU2j8Sv5E9sAggNW1InMd3jWc+7ODMK4UWCLw1IUhfZIjClEFjXhRK3U
9ZkjhDl0/7TiRX36brWzzXUPXp4sXf+kBJ9Eu5Bhy95IWfPLmFDNUoYomE9NT5L7+N4KlQr4dqTD
Jb29DbaaNQWQKkMDNOPwSTzuUYExoswFbraakf15xmfRnyI7Ekh3b46bwFCuTg8iGJuDZcUFgDg6
FugaHT4HfEkJRfIg44m0aD/auKaFUlWlwdYwyrTxpXyPgouQKb+h3mUwfB7/3RQ3Pl2Snk/yZK0H
Snt3YzDqyJMSaBCaa3MBwKi53tpYlzwY7eQ/G2CCnpC3dodf7vWfjCyx9jrFMwC35jDJJ15VOrcE
ez2yz8PtrRDKtRH87h0Ifw+y4fHIVLxx12beqT/TEAbhxJrMrbSrtOFJpb2yBNmufRduMcA1Ynlj
kR6kaKA261MpZPngEbGltufrsEyAc+r/GdZgDbQAgzyngnLRLiVxO0SKsCmjlD3asrUTHhWRrAC9
zf593Kh8yo293uC19YuuFkhlziZhC+TDYL42EBWnEvHeKNG4RWLmBseCXQfAiSomzHDw8qbBzMMN
m06p0GGbUVdFAotk9QYKctjZ9AR181KsM7Qul2rwvcOsIaPTiL6kB94AKHHr7H5nKb0XtJlvAol4
rBYVd/Xpe2cjKhsHrkaVZS3/gX+O3USVPBpNA1AwodU9olcC2anGEECQF2GQDisE0iwPyr6Xag9Y
Oehv/8bCNvKf3FHV9b2zu4KS175nXzeZJSc7H2+4X1/1GRIDlVdYJ3ad1uJgJiC/KY79xnpC4c6n
HhywoOiH82petE5AXhW+9NO7piOCjJCCfSRNC9/QksYrvK7iu3Za9eE/Y6Zkzx1uT8eKThBw7Ddr
jPCQ145YjZiS43p9ywYzdO6O7060Toiav17I7otGJVPYulJQ8UqeKEp/du0BfrjJBt9P1vSRYTut
XgDbFSGSn5U7BJa3+e1r/YNxE4TXf3oZbTm1ZG3uE7uSN7whGdGgQH4y7nSo0VZbjdPF/StBfqXz
IwDwIoOBkgg582amtAKSUtYvreiYg8D+fQT3cqCbG8Yk3fPFx+2CWHOuwlGWHuLmce6jKb8pHmSk
2ipK9Q2q5p6vE/zCn/07FylzuVIe4A17eUZCGDfszpapavvTA58SrpOPyJ5Dl4F5Hh7LE5Lq3L/K
IucJnEE+C9nGvWoejixJ4T0fUHiveQHiOa4VxbdD0Ne++6hwu1+wqpa8UjkYxBpIJshVND4zrw85
38BpUCAibC2PmGRBc/oF9LbcpBSOnnsHD0XQsDNPlU99MQ+AdMOoMdjHKFtjEySK/U0rjhNMU5DH
ZtAju7DJcinFrjxDz4w/xojBRMjCN5YHP8QJHkZSoipQx4EwMyNwjh6DtU7oAmcki/z2kTDr52yg
3c4JgcscXJOxfFL0mlSP5eIBmlUxHoj0H1wPkyCZ2cJ6DTMkCNvJk5bYpzXPnx2FaoU8wkAPJtXD
8tWSxOkrw1tuP/jYWHuS0NE7Iem9QzMWepomVecLvlSZ5ppGYb5ftiVRi/itnHFwB8N1Z9DrvgzA
o+CiPVLuR0GrkHdrJpCsGlZ5Ilpt1vVq33F3K3ZhcVprvdWfcNJZ7Uyr670p2bvEjQi0fd8mruK/
UhjzCnXvyQdYn4fi3WMyMfIHik6A/jV1ArYT65RtnqVzexMGP7+/HoltxJpV9bH8abouqpHsnWNo
dEsBoIijZEiWiVxhSUIgO9A0zStHcH3aQ5dLHNzGu9mRTnmAL7Yx+slpdbtMCrTV0Sb/4Neo4bSJ
sgUnsST0vNcEMjm8cfeRt39/ddZdD611GZ3kUJFfMyVLpVE9mltWD+pA49uCuoq7H2/xing8PH4S
PwvYNQf2YDOlYRpDrmhXV0uQ46Id4nbgqy0PR8Eqdynv+HkD1zvFViidIQb0ql3IATthTJz5kzu2
IuuSEihIpbEGM2z3I96toDM8/K2y+GqGOgBQMcMvd4qri07bqI+XOsz1x90mAf6hUNgb0MsJpYE1
O5od2dw5Tv8ITUMvdH9N4l7Iia/oTFjrsIUy6QQ+yQttFomaqirT98Z+/+aqA78XuifMFHaEuRs3
Lq585MHimmFHIc7MIjx283JV/vNKtTSpRVDMEPXW8/HwKsb5Va3WCyj16uv/mOQ109iAMA4H3Or3
RJu9o9kt7zJhzvqqGL+TtWbQIGTUhk6Ah/Xumjz8eGMGVLBirmeudUTFCUkJMyoXHYJUJhk2siCC
0801sbywkS4OUJ/xsj64BJISGbX44QkKVcrS98/E1oiPcccyD+chSn42abHA5tFkYhtpet2IigXB
TzeHYRlC0d5FfpWJpcbIEj6TYW9K/vwzZ7bTg4IQWIheVHx9JgdVrnnOXg6VXsiPHH+915Uw1eEZ
hj5SKUADmwMrB4v1gLT8ZWmF2v+DMnPKWmtRvuBlHmvOMm421BF+MuvPkoobcjk+b65MVHrJZzMa
ojBXkz01Xd5Cx0/Ul9SnqQFNVUj5sY8jibo4QufGxPhdUKiwNHC2hF6ghGwm5wO5piyjnlBApQUz
DvpxdMuu6w6NoroTe6wY4nXGQtqgzTiAGByJrg0+gRKJNUmaYMdwl++Ldzhki4zpfX4aZ0okMHcN
alkcu45GUGzE4daws9B7BiFkELf8H3ZNx2AeWLi7coZK3ehR00JbWFMypNKpHvG7g2m7fN4co83o
lJCQ96xbxXknYbeLsHtArirhSS/2juFoL27oJ0s19vFViDGXJ3u21gELoBUs7qwJM2AxuOx8evoB
ngBThPeUzdLTf3W1XUxGTdHgjNBpW8Id2s67VVZ3xOksulAsBBj2IvMOqti6pIBbz98sYdyMSb4L
JYkYPFzQXh822N2pWm2luzTi0Ziku88Nq5tCgOwzr4XqjKo6Hk8MFO89OEydYVqAfiPfY1L8IsO0
ghi4PPvCzXzAtd2T52DA8yvgxe3GbplzrFpcyFVFWysq3UUuWtANXTuBCr2Mp8mQSqzNiLaMp9QC
mPNJ6ufALJtFIflayYEpIVO0IDAek975lLjOdxSSJuwNnl/wPGH3fsTOgmFbl6qDTxLt8U3PHte6
cxtWbR/FvEVgndxHFKbzJ4XDhbTu2Gpa+kS5teOkdQdm6XfKXuBvTxLSJ7iu/gzUV9mU5NEjrI/Q
7FwFmxmhPeLj2WCNRycS1w/3qgNgvDmj2stTAO7K/wUx2m9zQ6HIO2jBLCKuhBcZtyT3pG7fkgAr
9yvMUgG42kwN7gnxWr75ElwP9tCOz1UOb/9Oa7Z+m0kdl8vol/VFSZuYMrua6mJsIWERM612UtbY
6xPABHqN+KY8Oyjucp3jlYXXs0Wpj6U1BgrfiDKHAjgI9kk5Rm3u3PAwgjIqV1rcqkGLO8+WvcOI
TFo2g/TMB5Xk1YMFVjseXGZBNkhX3Vqy9YNbEvuBYBLrRcgMIv9DbiimxPnb4VGqeK5mTN6bQ9L8
4Hft+FRtDbBSJomFDtDAtiApY9PwWxqX1lUmVGtbC8d/WBTPacCjWPcJY0V3qtqgbF8w4fwPvNzs
PLl86dC0XHNhSVpQKhWjDPB/1saKl3QJPy+vDSscr4r9zZiiM7fxedE2iIADE4ffSfsP0v7uLGXw
DJBazSg7Bikb9rVwlx+UfvY5j1c7yb7zNwAtUeXaBVmd1gCnTVn+QYqxmjpnjhBAUNtzBJARbZBB
68qKBdnzD/VSWaThCqLokx/0o5dGI42CjS9fgv3Az0dfGOCbDlPJnmOhmGucg3s0YMv55KhgTD3W
uMIHC0QXUqNJ1hCxlT7S6z+ZMVVxmFdW4k7WNg7uO6gjh7R4Sj6bY0Zy78412IHbxWjs/+tdMVbK
+pdTPVknSpLJI+dIp3QSUXSFdgRn0dxOY2P1r9lRO6BrOYXNTT6a9JALaCoA6hUMi/90U5pYmZXC
KWsfPveBT0497WCB69xlepAhsnqA6grzufHS3Z2O1IsIYVGOAGC2Ad/RnsI1MtKzVSONAQ3KgWZl
LvRepIGPZFjm7t5loMYcUFVedhe8B6oP11Ffb2jFvP+Qwu3k7ll6QMMlcp7/fqWKS2kjEgVlM1jw
3w+ATtx8y2QHZAUF1erYMJWohhc/1ZQ4KEd/eFtMMu2wbKvcyxlQpHXRAcDiVKQifnux31PehaTP
QRBuK8gCa0HnxpFj7ghDhQwDXLwiOXf9+DZYS8BGp4sE3aZmjo5pfXhiXAphEq6mEqq9KcVQmBb9
Wz1M1eQs9olpNFWGxdxBnqUXpNtIvbcL3x5h4DBQ6vlYLqp30XNwmRq+SXEU54QtKuv7JKyShR9U
WguaoAmKtnSGc6xHkzdvWbx68jDELz2oU/M0zULClrxsplcI3A9lpbz/c6iv+tQt3E+EttaXxYRK
fX3Ps5kN9dBxACJuFovbqORSVDpN7vfazrufk3CsXI+cQctDXEC1psvZp2J0l+SsDmrDP8/fyfEx
muj41sErPb5Il41NX11R63Vmp6tGzEru3r/3TudgJxiaIqI94Pk2DbDMLS95QCYgW3b4LU8W6CPi
8U+Swka2sd33HCZpvvQjWQY1m+mEo5IE8xBVD+4gpleMFAGzzX0lifg0CP7vD7CYW1C1ML7ZcZg+
t/V2B6QVyaTmeO9tNg95NqaRsOiK3X7UN0DxJFPYo4Wj0bbDMw/m0D/RPrvdj4xzWMlJYwhcedG8
zDqwOyanmiE8ND808RMJEl3CClKYkSqN0YjxirRvxvhWvSOFRAA5pC79d4lAu+YTQplWYYtFdsLZ
hjMBqVM0QJhff+FewUDeY+SUfN7fe6dhJ4boFuINSxGUhg+5EVKTjWNAUNgXQMYKJngS5K2np2G2
+OdU/4cS18uOAdi07bxVvKhXCIiKdYOVy3CJuRgsKCO9Pyj1e9HxyrHMQ0VgFgCtRWo1muljmnQf
ej8R+uen7UBWPsB7HRAuaBsNK8pEodn2tM+LqNWyHAYod5u+6lPFGOaqLmSF7wEyaOlT4LYBLNPp
3NWBSO5WApoYxjShIQKCP8nCq6fPRYlYM1klt6FzadXVIrngfku5el9jE0q6yzgrik3kPZmbPCtc
gu4Q1upbx6JLh1uoEJmgxbMQ0gLSrGDdm4wvogOXdRdF9Sa0ZkkXVLBR5j/z14O/RkFHspN+pIgw
R4kIdkJz2K+NzXmBX7C9JaDLxQYOZ/WRDDaOlLaFeFkPd6WQpl/21JytxXOMQUSOhcgXb0wvJ2N8
UM3Eu5zSjP9ToHF0ZntCjEx6CJsUrGgAYyMttvMq9CyVjTGC2Ms2+dvWT8qARrDlncFoUfBazpFZ
SZmh9dtkQ4v/iMbkQWTx2/Zk7V7LlhB8+NaSscKgwOK6Euyf3bGeO6gpH4FoFg0qo9s8BS54Ax1Z
A6LXegpdnm03J6AJ+ddwaQzOKT5ARXRxeAi9tFvafhZCXl1B9zsVcM5EDMAPaBgUVQmfR5zrDc8s
NGOXVuCM1jI7BPF52twnKKho6KmDLONVMxRMIcuk9AT0LgBs7k2mOIjQO/xapmRJYOVvMwQ/Zy4J
bC+KLwg/tUFXGo9B7orNp2fwvwUkYHUaLItQxjlKF0LZE3xanm1WlRnf7sfZi/w2j4+ox34R47of
jId/2MW0LO++wKlSiAwkH3iQJA08X44nrzdnuvihDuGxqfZT9behw83cgrixwxVXN7mhUxwLV1HE
Qix2b0UrhQJp2ilul8VlQNS8G1Zyz1q9k/xdt8Ovno7lEq2bjkKwwiIHaLG46Ndeiwz9F5d6GyFG
TtWvEBTTf+BUQnT2XPavydZH+Nkp7AdcI4/KigIoz32HJhee2E0dTN7pGv1UDRjDq25GP707gg6Q
oxqHZcG800ctOc/mEqBCftH0pz6V+IGPpmXMB9BwlGkD2+1SezaGvhhBJ+yoV/5nmt2kx11OiyIA
4N5Rt4gASknHxHgI50lz/T3dNiSFc28ly6yxsW4sU+aoekTKNu+qcfw/PnaFGPLvwYDQVW4avae/
EsqeDOyr6fBWxzXd6GZew9cBPW52xAyQDG9iuerzGnJnaqXoiKueQGedHH1lLf4rKjRqAJQcagJX
P6iPJQMaNPbsOK62Q+v3+FCnx2mE41dyRP9cmD9wT+uLXMtt1jvJY8/wVkfnWmtJk5m0orqc3l/s
7oS/eaJpIqjtSIjpwW7H4d6jfq9FSdvkycNVw+Q3U/sYVaMIR2JYZ9R+jdtvww7jbsPv0o3XkCCw
Odoimq66/d23f9JdJYAB6YlcrzA1sPLBR/IKPiToTqAOpm2cF5wxwAx43paTlC9aPo//sFOzbQ3M
VILXt6QHG1DREN1FtA96deZZkUOPuZfnsumEWVSjXPfGptX2wyV+VTyps36Zg364Iwb/cM8QISXv
YX/fOt2RvrCqEslHC76KH/YzacH4urvGQCEbZNgruM2YiwKcKBbH4Fh5jlsF41/fm3Ftvm4LLZKE
YPkPlRosAlnDiczW4nXfl2riz6KmcB18rmMBOS9uv+anZkNHHiJAJm2gBMYAnEkLPAk9WUypl/CJ
uvdoYXquasv4TE97CVkmOohMMFmpwenS/iLw0vM3GXWNp+TqQeJymHgu4gujr1+a9d0og/iaU/ks
gaWrrxVu4Bin6ERPhcIBbJAxCPVsGZD9zPefKXroUfcKzrjnQsu3epMPRjxi8lXLhOgncVhObI6q
DSYgTVf9kL93jlQdSRn1kwC2El1NpBHPGd/+pzF5g8k+B+sGq/eolX3PHvA+VVIVeaU98UFdG6hC
GqKe+G7VIyhBaJ5HwCsmv6oZ9SrqMwbvM0nlDhbwD7kAXcNtpkX8ONPoOLrksL3DIOjxAgUjwoZ6
gzuSJd5EItsG05AkpZl37wE/giU03U7IEKqfLlwZJBG6pT7ravB6BE2mP0nMt/7MGGdyQg/3F1Qf
orbjnfK4sZOQS0FRR2oZnFoGor9n7RNpWuSXRJ8/cfg/4/pdhkN2Lv7tPskVx/7QlMdjbzc+b51s
ZtoeyrCCIJMuL8Pc6m1aLwhKxoHlqKylN3ZZRacV0etEojmZa+ZCwiYnSe/K3Xk8ly0QXJQgHgYT
VkiJPiAe/JKLg7CAss+wEk7GaM9d47FmQ7g6+Aees+Teas2YIuOBrhc03W4N05lOxEm0qL2gOUaE
grPG0Alt2CfIwsM8JRB3W89MhNfSIF/5Ni95efOW6rOzHYTD/27UR3OHOjiqHDnPEoVVzh6tL/Fx
jWlP7y4jikjYXN0Np05HM3YDei+1YuNclGXl7+Q+JAQoHCIfQ7ntiBkmioLCIGNbtST/e3YkySuF
IIe9UdKS1QDmyxmmE2sPMmuVBhd09JLPXxIAnid/Xtxp5uLTXyMLsM43ztYoF+rdcNjZyHg0gavV
aXTfLJNwZ1gya13jpW1tNBO+YiLgYBZ0oLQuL5yLr8u7mCSmpDpACsSGn+BVgYpHBjKDuIlgqpAr
gwgo8AyB5n690s3/39DscsB+MbI+UPLZyYMKR+t0mltWTzSDVeFGlz5gAXvUUBDs1QTr04EGeqOu
OBvjAuSdhI61khwjIF+V1QxWhnMRdxcSpKX4RpGkNJd7MBcDBfggY6KrLZKcOcfQKciODBcgHnpt
gwCfca5Gj8dGBKDnlUVeU0/m/H0XdVwtoyvihHFNozGFXSc71gdGhdnC2ZuVJFbVKavCxhSL/AEX
KeiJm8Zz0Ra229JrVXlRLGuadF1Q9GKoxwXOA8ui7XAx/2U6dNvvBTrF3ammIhryA0nvGvrb2S++
oHmBTtxXw8Qpmrzcs5urJIJGOknwTsYTNfBWl4fWYq38WmYVunn9L9Jr7HllRnScU0z3tcoMUIb7
Q8qMfPQ3m56etq3/5MzFLhhjzbBO/fifGKcAxHDi/L4m2QdWP9LfZT/t6DoVRZveg/bnZL9RAWT4
Dhj5QsysjwXLDRp7lRtbmRTxCoZT+B1Y1jJDlrXmEIT4tphvK5Enf5GUu4uFafpEBbIk1kzRVW8y
R3paNcmnWoVfx3Zf4FHS+PFjA0F77F2UPREEaOVB1lVMer8ChzY/68wjo+aVy1zvl6JCT5EGcawV
66SdZtRgFiOvIGxt22UWoAOtqfr256d3cH6uvrcoVVGKVvWjTENDtr1rZN17Q+ggTq2W3TIBbXk7
ysK3F7m3OTpLoF/O1yuPPCNLrtfCmiTgRHm/jtHcxEhezLrtnzI9YSO6k+3i2B3CzDUlC+20eexk
kHOOcAh3u2jMsUvcwlV0zrqL7W1pt+EXFvxO0xk+R7fsVJIaOea/y758uGzxDbwMbkXO0db7qR6I
HEFK9K+6sNFr2xRtCXenSnEmDRp5Nous6J7SusvzzfpNAMWMgcCjGyezH3WcpwFpYvdF0OPZqN6b
W92T0KgNvb/Jr+JosvJ6cRMPLAvjdHJm40vn3BbASDfS0uzb3fR7Qv86Rv8I2D3TqbKQSeJWr5RJ
8v7AA6o6hRp8XaP78T2iGtLjdvnnxxHYWl3JFGdhJzLI5jZ3EFLOReP8gZjh5r9nGZWCSU+gu1jF
J7gnDN+63d7R2/wQT0qnaFMabhna/jLLXChT0oSSmEqRhs4pmH6PVd5gGa3czENQLaP3MMAXSPu6
h4vjs3bpWDpGGICmdcR4Jv+Ow6U73qdHzsI0soe3S70N+6ujakeIl69wonHbjLIrE5Vsg9hS42Ab
wWRob8f1ic9vrwkv11mdkIE2QRkmuITpJcYosdn2Rki2JpdvlARDXNsi4/ea0qYJboa9DqYmX3Qp
SG1C8aZcO3PjLxWGNkZKwyJNLb/wFInpCqLWs4YR84AobD9+T9nNrmLJpSV/4vOdwwbH3emYDIi8
hpYkoABwi4Yog1wCW2wLAlGmJnelaVnI+7v38U/nAYsCzt2mRrvibrqzIR66d5y8Wlb1RVfeEroz
Zr8iYpB/vnFis5Wwzc92OUAnQ42UJPoH/a2njUl7hQTQunaEwDgDRq9G5IF5tadNpnJ+VOhSA9Pa
UwVxzEJof7yM+yI1jvCW5OBB3LVQE8SUWsQ2sXVmb0H/TLRSKTLbq3DpOYeBknMkviDlsi9XyeZd
Dj4noaFd9WWIxHuhVZXnJHLgiMBRB0tha7Tv1ZEXYN1dac3qw6+KumVU6tFXHNaXOxAz+ZqlKcHg
4s36/bd7l/Sp4Hyfs6hEjZHMehsGr1mFj0GWvPBaUnZzt8uV+KhOBY7olF714xHgoFfwtZ7grxa8
AOMQ2plwojrDzMjlvHy4vTv00dCePqTMRQAJtOu9IjF/5ILGODJmGv41gWIlrceEiuZeS6L40i+F
ZIlDAkjbE2k8B0bsurxNO2om97Wfn3bA6FRGZxfFhGaMiNoztKkX+JhdZPTeYbW3n8RB9Y9UFOzR
Lv82ZbQsbOpZsV6a7WFucuZwY70KKYWj5vM85y2xCON3yUqQR6FOGcKqY7PBSG8J5ZK15qQonQ6V
2LyWNrPQX/7Dj4wD/bK+RsxmxJqPhHw+YZO0LQryvX9OTKrm7EVBvv8dQDQElBaNO5NswzqzQa8D
YuuCihHJbubH5wLielYR5s5Js3OSDzpH18ubK0nGOsgpKxFkgy0z8HZgqvRUM6NK319dqPOTXaLK
poWiLx5r0z0+puWSjFKk0jZGWFNKwyqwIqqpUJZqDOaeZasganILGghQ8dUNfQZvQazhhzyClZtO
JGkz5Z5lX/FV64yKzG+dsj5FFdy+XS5IW3Q9kEWEJnzgOH+zOR0TOIn5JVTu42+hjI/VVEYe95tS
sI3UHcYLbcvkO3FcHyKg5uKQfOuh9hlXTxmX6RAQONCBGEpZ/gNkuR8v3d88NZvjmFy1BQo2sOJv
hbujo98PQTWAsz0cb6o7bE6lNEK7Ti5TunGdtMgOWZzhojDTMplC5Yf4be9P6Wo4Omz2+JjTSkBe
ndoLMLEwpKs0Cq+AzPpPlLr7TJbt8hE1ihIMxkEXwK7Pd0LyR48Tt70RflRiAqD4d20FnN1+W+qv
oc+PXDTw0QfkQhOIwbEk3ROq+0l3VV1mwS32Rh/xKe1W3F6XQhFLreGprHz1xfE2oZS40lS9nGNL
ijPbg9oqq1QnqbpPy+Xgo4ZMtW4M4ld4HfXb3H3fUe3404WLv2px7jNdsLoWWLm9Wr3MRpKTk58O
0s2zc9bEkryrQGiQyGkqTDNWuYhMDDvL3vLKS/i2e9xamI4iANO+lu8ZZDqHjRnpeBagv6DiPfR7
UbASfEjgpaCWoS1vdhZinFIfk9i624+nCXzXctzBM0SwAdKyfeoAou8YZPmZshcAcy4iHSOybBMq
12GVHWRSsey/pRHoJ0+6kgcZVIl/uV7htT4RyJ0AiStAuCUL3AaeZGgSLeDEpYlXytwl8g+zEJ+i
rwsvlBVaQSA+DTyj3Ly46prYipxqBx/CjQhMA1niqKU9XgvpN3M2zl1/iHNFTmiMe4Wbjj3RDOK0
T3G84fqgdbr6W9og+8OnkWjvWBgF2b3v1d4kKf5dM2Cp1DpBCGnXRd4QmJYPBuc2dAQ9pHUTRmMX
J8MugRgvtTfTKvhiRMjqHyumtl9c9kGAyCCQUOABud5K/FFUtd7Ts6BoyDhWmeg35OseE+sN7HeN
/9/9U6OcW0pIcuACXZ3F1hxF/GoxpprDwOPlgld8qdMK0iZ0nt1AKbL5nq5EOJYflTle24UwR3WJ
ieMtYJly8U+XlUltONrLpMFF6gwPKlPYMnKnFGF/4t3pvv2yiJQ/4cmf2/wBKuzj/jofPhgVWOgu
AIunM+kHvKHdfi+ZWGyfnejYadzLOcTmau3bUPeL9BIBkIvLuvw5HvngB9kzXSHcelI6AJd07G+r
r/DL7IRFaUCgrMj0M6gKcmJWS7pRDxlCgoeAfpOjrO1dP+VljvCrEl1pGk6iSiFpwkAIo787Oy2C
NVWjbnr1hE56MQBiLiiIhmVzQHDZG2MctfyDSnCqIXsRKCUKbk/g7FAFpJ0bZEY6tPng/6xuBR6R
KcMW7xow7o6k5FTjWvogBJbKAc4FsJLasNUCS/NTAI8RLNSWR2/37MwOsVbZpn1B0deUHmEOOdCt
IVayagTU3tHdXvSCKTJKnQ41eFK+77sc5wj5+nmJs2avjILDTLixKXsF6zSy4059uvdc7nLA+0nO
ZUu6T23E56Vo0lHw5eApgLYDy5FY3ncoVr0T3pWIBBHO9jtfhOPYlx1Q9UNajmt+U4m4NU4RJpCA
lh/YpFfNNcDcbQeUS1rVZ9VIfXlRn6PWRNzyjOQcp4yMTJh+hpidkLQdrkYzbeEUkK1TqV/6VG9Q
sGBjbU/P5ze/KdqOa+j27i0bKHnm0zEBkTBrRyOOZKdmb0+lkw0EZJu4vrhxRSpffetEQqoCpMUz
8MTEVUmMpTK/9bfgYi4BBn9j0K/7KzexWYAZwZQXu6EZ2WFJMPWJN6w2YH7mF+g4QQ2l3X7e5VFn
oUGGZ0YhWBzzgj2PH/G/z3FcgCYbUD3dh/UBf4Mx8A6fnkvMvdBPK3kcn/fLsaJ+sj9sgoqYMiLg
PeyZmyLe7o66hGtwr+oLZww3MKorPerFLwNZe5OU7SjaN+KET2LwcYxyb6BluR1QzhS/j8fvJ3Wh
T6vC1UMSST/zbmtDCwZwQD1YP1UbhyZPDyLonrronrQN8XcpCKp0tuFc28xKsXegTrJ24Rpkizbj
mLmBM1jfbdnNeqSSGJeWorbxKTensykzUgYZ0khpwE3DCrmHLw0QBtweaYWFOhcVXz0O4qxXN2UJ
vmDv0iEgwmFfw7j9An5Rr2y3iIS64Od0xP/xjhGJ9TZdpd6QRrSf7TZhQMTjMWW0znx6kj6QwvIR
aBzU7bOll3OJTtu77mA2+gkBD1P3iVdnbutFB11BILdmI1GcTELAXISf3TMlQCOyHVCnxiBBUdnt
5Hx62rqEFNLE8IydEjBNYZTxdxKDRKyWcIG5VuHAZWh12MEvc2H5lj7urFfXVA4TDimFbQj3FKu0
RHzD/EB9oS78+W5Uy+y6YrAdFlweso3oVgmlfUBu50jrdBi6GSFq7u9SxYSWZRSbL53xnW/+9N4N
Dl7V856Ec4AJiVTEnhFmEl0gtA0I1Q5a3RdmAu0hVBuRjO5ezOKh31DzyCQBgc7usLSG4vxjCBXP
rpdO0641ZzSJNqNVxhk7bDChQ/E+2JdFu4gC6A5YkZ4XfyXv9B49MOa1jlhl5BmnNLmVWcDlfzsf
YkSt0o9TF+bd8sBCXt5Ds3NfNH5swP3TH/J8/6dAwY3C/bbdeMWO1LDRj/ehXNu5XjKamQonyusZ
tT+e7h8AzgJL7AWbrD1pOG13rV2XEW0F6UqAEs4lLK2sOZXe0B1XH6oa6TmyixqKVkTm2IXHnGO4
c6gJzS1TRITK/g/LahFXCjy99JPn2zeMi+qj2QCkt7Wga5tyTEDKfZ7ld9ugammKZsv6aqaF0OPw
xWhhFsToXHNWNxubl/juoB+vikXpXxeycn17nzeL9Mygoax6vcL7FrBifw1a1EPdN+tbwxKb1HKe
9Xq9g801UuCxlHOxW88PWzyRHj8rAebClVN8Xdh4YAvGs8YEIyXuQfQXSW8yKVYX+wWm7rcB74e9
5mgp/CeegWncaaTP6zNdD2BWRjM0bA1q/zAAhkM5xdTTw3UN+Z5xpOmlB1rDJe2BLXHoB/464ndz
FbM0NBjGvKcFjveQdaK3X8Jly8tXUDm/U/F1TSRBpiICTvpQ2fz052BluKWoV413Bdbt9Nucpl4I
5NQmRmyOqfSaNxWE0DQdkZOIfUGXkZ7ksFjtMEU5sKMC77Cd1ebmfNxXqZYS7pPAo3Eq9uiwuIua
l2wO3sJafhjsK3Mlmf2pcVT1XmGmCtsx0KTxx3IcFGi8W+5BhIZhr8owJ9mwL83GzBkYcJVHsg3V
h65dlEUAXHgcDtdE/pehsOvY9j0Ntew6Lsg/XVSSXQ8RAtD/WhEFihFIx2SLS+H6eTMxu/POr/uh
BOGM7q7UhhdHPgWFdgLW7wh94IfirA9JVGTHWmGW8S9p0q+qnleE1iAi3k23Nc6SZu+QojhoGA4m
s/6dT0I1qwOmO1vVTGau0ZZhLMKc8Bd/sSAWAE2APSHXyW0WKxbO9Deq1BDSvZ3WsxZuVloDZzw1
/LUDm4F1qrbAeXG7G0yfsVPPoT3s75kEndNQkkuxVgoM/6VcfCOvfIMBBDrUWeXYTrWl3eMkhasD
XgKZQSRggTXMPz9Z6rYECR3fQRRdrsGRFT2SSFoPMTHHbN+ZLMC3tCFNRyXEpZdEgh6LcIEMTQZW
jVeU718kL/pYrtR/4KIeLHZCjEmd3DQprsiZCdi142ckA3bAKGnbp1jOJReLy0rGzNZvf8PCU5ag
bdOznv5mTTx74nThSCDpHqnJP0kQiQf2ICxl9spVIizrx1sHcBw5V5e7q/l0Ci1LcYIPJ7+hdIoB
NUb8iPlVxF3Ch8ga6pHk0A5FfJ8bREvSvhuSO2CtEHEPJz0+F6vAIPkU0WZnNFRRDDKLSS5KWgeA
DOpFI3Wj7xOb8aKv0RSbOBAQIS6st1GYr+U4K7S2/2NMp9k6rJQqwus3uutnNXI9J2ZkFWMLpl0h
nRrCeKYiYCp41kSRCb40f4DuVsjsTSiRTg3ZttFcmkzuvFT6CBTWLMyAXp54CHsNMhrV1CgHt00A
Y7ypX8inLLWB/k+1OfqYD5Ikz4cyyJRVtPMBJc1q8EE5+RedvMoYnIW9FMPExxopegKPnjwoqIoL
hvTfjh5ViAlRbss1O04oJO08Ebt6zGKGuDk6kTatYxGtXJWEULkY6bXoyWkerXrq0w59MZDrj1UC
YrKELiE6OmRgn5L/EhDvF8YedCi1sxYp3mPSjMS76LM3baXXarjLn74TLjXeuQkpVVvBcVaAQai2
MHsDCUTdYT2Efa4rIQ7d9iXYdhGr4q9Wm9HF26u/51eZ+rww9nITjMk51VTtxD8hocGJBU2iTWF2
BLIJAEfTPSl123Ps+t/zyrvFSzcfukeo4pAwTX5O/a9aFpH+TxfcAoxQ01CAP12IDnLOhoCciQlz
mP+bzhjg2v1EawLFJKo9N8Y1p+QBaDZCkLehvfvNbxlC+6STIPTkgMBbuwFihKfsty/eg4HoclPc
sZiGh1G0vJza5WVFHCftDc6qoIpytlXL8TgI0bOrQB9HeBraQKPsZpcShDXMEUMoJg91LlnMcf71
eKQAZlDysyXqWRhI+0vDeNHbdJw0PU83iQNKc4GPIk0QrZtLvl4Y8bJbUOYwE9kv4L6kHl4+D8Bc
XF/dlU0s0rxlKlz2GoHi9KtiH7ew2d6gNo0SK2rRdVt3FEGkL1kIAH3QEebgOWtNsu3BnrLhnzXu
vyDTEo9K8ggLYSKvWYI5AyyIyCKPXhIBt9cdXUTKbUI3CBkBWFqGnWB891Fsfbyz72Qbl97BnxeZ
sdaSFD6sqeLh+GbtU+gkMDfQREligDWHEFQD7l+WmYzMwPHp2ss8C8+FmHKGQ6AhBSWHTM+dPzeD
Ev7lRWLoHUBM+QRAHkhqT8ZDpk+YewFDkvGgtw+T0KWgQXVjJP7jrWbOmyBPe4mEiZt5aiot4Dgi
zAjBWXrizwLdpnNMB5ELYI7MVsffdrf1A6Om1gCT3vXFo/8MWZdMTp/1OGNKuGWqHD/ye45+ccD9
MjPKS3cxRBFfzywZcsr/t1xkV8b5amhPm4RiFzjc2qIg21ufETh2+6N0X3eBGURdbvcGVF347Ui2
FRdv6FgW57LyATcirzkX181tPXggRemxBDfs9X73X6qVWdS3lM/b/r49LHZFhmsW1IonkioF7nqP
Ti8NcPxS7tY91K1q3As3I4EnAfNKd5/sKC27tM/xWLzx2bPEjPt7Fb+TJ3Njrt18Q8fJLON+qKqT
HOiA+WTjlr4VMAgld/ZxF5BC85Fpllk7xovxSdyEbgHOBz2fMtmGc5lwNuZMldOTJZ5UdG+7a0HZ
x9pw+eHm5hj3UCYU0VLiRWQ7X0y6j0XaVwhBLL3I63dk+0120vZw9Tlmjrq+bWAFxzgGmtbPvmUM
zaOLfF3FplQ7i7QJ1uymmclWzuHQNuOQfCEkVL14chZ0EosdNjl7P0xGWYzZ2IDdvOiAUFrZxk/9
F3sX+1U5YZWVHcddyqeabYC6RWa7Gar4cYJ1nniGQYFe3GNn8fkXmiPyrD5TuKgQ6QhSIHMeyTUC
3AEBKXg7yH6rwJO+MTgYwRCYfP8jaqIlO1UOGpKFl/TLa7+vd2NtFuktGZJNoAvphqQY2bH3+nxz
8A8vNr8JtMafvBPsaaFOXxJBPVp2xqM0HCfE0AKAOkxyZV9vcRveNhqa++v0x0MRVe7QMcPjzfqx
3l0PFHIMc6uaO0nMniT6AGfxx7MX8WqWmGAvtixaKdp1IWDNh2uRWoATV+tco/KHc/khkdBo96sj
wNwuRDCeCd+KL1Ydiw1eoY5WAKXv4miJ2X6BLGy9gQkQvWC9KehBHgmVP9DutDIx+Z5xjJJYLSip
VxRKqLkhEPpgrbq6nQhfMOWVN4mkz2c3jIerSOc/qde/VoK2cbwmCYHNkIDWAQSyUAQ5CETP+S8x
ef1Ys6h/7nf5JfJoBYQEwUJZIlgZwaTcPLfVG3RXLYDE9mjFTN8BiM2ViHaOpb75OzsnwWAhMPTQ
KffAa8U1/SGjF2SLuj5pD1kbmSo024kA57AfkE4P+d/JP71IQBlUMF37TXgKvufVhsQsMpk+ftWW
2NQYF6dnb2SUSz7mzkPKDEqq6BmNn+Gyf61uAlj0TRAo+nSAPeiNmXyUIeq9ZP9jf27pPoQDNUl9
MaEWBOEfi/ve7W/2J4tzjeff5TZc+IygnUKlhwZZFsGa8chMIwDcEwkNXNiiRe6y3rSQ4wuEzvSW
TsPL+LVoORKFjN8i5kaQAz3HcjKJMATCxMX73arYKV2MnkYNpV0utQ+qxAAvcD/xIjt/jbl3xayw
Lht9hvw1Znsc8gc1vHY/Fw/FuXhu/8JTzGmyZ0PxnUw+ZcvrbSfEZjn3tOv9VmK8d2o5UbOr6ql1
sqYW4wicBP3N++dkZknnooNFAGCmWqfbyeytJNldHeTzAF+/RTrGrDjxb0sKlPZ2bs4As42OPUVP
qz04Y2XnyZmPcd5QWPLx9v7/OmuVF0CWIXo/cLiueDRVBc0B/xDnM73uZTepQ77uvW7WRVaZ56q3
7BFDSfdVI60xyhQW2TaQrPeO/sn2GW38D1xY9Ofzv0Hy+dpQEvQGjXpvjU8kOvl+X1hkmUc7NImX
iD/oLEm8AFp+2LwovfFSpqzOmHWRRkNPGGLRE7pis/Hki+90Akva+H4d05kZoFlpDIcXtdmU7v1H
KfXXYzKet1/3PKLTqPUsTpcI0IjARu//+G8Orv0znDoVFCoUDhHVw0eYlk5f90roERYl+5CLqN9z
AaYb4zW99etxWXYRxNvofzkl8BMNwS6z2YxEatUmC0hdrxISbyf4tQMDJEkcFNKMokFicUz+h18l
s94zjcfNaVbZ1drb6QeXvOPLqsHbDLB+hBuSv/KE+JRGt2HciCPHG7NkEzDhNs0EQohjl+X2x6Nd
sq2SURAHtFWM3rvqhQxQMew12+83jV7KukNifv/qLhtUOLwFZHaZZLpKicHDS8lZQ2SmZgsCdUPW
oVrmj18VuReKI8zJoHILpuyhQykRNC+gyAO2KdGyQfOP2IwEtw1BqP93VRiG8G/cGdQWZPpBotur
A5PhmPVqtR/7+VGt976E9MOhUod8nmel4ajeoL82L+KF49SUTwh9zxS8wCxIAtfZCqWO6RsNSL1n
GUX0PmcuvX/8N9reu3QglfMvORhnMNLVIz2v7+0LsmX0IlxsmfXlvuRQrKOMTyDTWF1CHA5ckxD2
PbvIyq6jt8ISeZ3hrd9twrHn6ztFzBA/3FfCai8A64sWX6OSVjP6vcnbViBvCH16reKMd1aZi+v0
9EhSSWLoQtuWVOyPrUJ9OAsSPfl7fWwBnHy+WFxPp0LQRWT4Zrt93TJKSc5qEfHXEk8m+JKmhsaF
MO30wKNyyHeEpHTJt5ud0JiOlk6sf3Op1+AAtBWHKOnXPLEXwP1lhRDDEJeb/L0stjT3pRPRdMgO
qHUoZKjYYhsmlRYe4CnidU5+ZtOUeZX47Qk2Hk6o6o9GtTQ1npjrgf6+pdF3xBGjC1hrAIqCtNjK
Q0cOixoDkfAjfB13N6UtPvRma65ckhcxUyoFeDTSI9XW0yBmvUW4MEg/x3kvZ5O3fdDsUt5kWkIP
XPfbg90NyuqttCB2IRuNXrnI2mOFUOtyCTUnIrRheS1w+zPPW49NTRKkkaPn3y9tkp7uqRUxSiKe
TAPVhpWV/PEciTCduzaulpUwjbaxRdMAIznJE8/cSlj1y83Ht+JjmR8c+cHYfMTIcTBBg9+5YzEQ
YWTI9dS31PCCoR4tp1ilc20lb2y0xScj7OS/CmpjW5NIerTksUaBQdmc4qUHL/KvXhHeztjFyYr5
AtCpLGJlvHEZ9pmEr56ZNOrMeN6cASoXbm6YSJ3NELdtpyPUNYDMQlhw0+D7+ekzfDk6edDUSg8E
zGuZwWEySyCKQV48GUWPvTHuMsfFVa0wqRyB2N033nXvK8wUjJeFRLqlh3PC4equGvVWYhQbcR4W
O8vXmh3y2EbcMpydJnREX3iIZLc985y1S8fTJ6Iy1hoiCaXezLBgEbZeRWthwhZnJG7uF+u+PLNL
EdxhgLTTUVqBTkmS4AxcNcaRdpkI4WeddNyUxvYIJ0rXGkGhD8ttOX9coodRVuYW5bf8CWBwz93T
2rDOHDFvyjkt7f3Q0nUw4VSf+dvwEsKFxmqnvgkoNxr5twt4DyKmIKMbpznKtDh9mzEIGWH2MCUp
cJH9jedL4ZxPo5Rf9BfyTQ3yjoRDc/nJ13Ax0IUTaocYIYOFPpMRpfa5fGhS8Ixc3nPhgZOZukKZ
TF3Rr3afYaajO4K5YF6yJjmu33D8kwATTd4pfJ54E2MLE32pC+TJxXJiY6bpMzzEzqFpvOF1LWbo
Ou6Mhv3HdbwyBpBVf7AAyOX62KeAKbescm9tJvrVRV0Se2T3OeGaLnTdbsYtUoD+JsuZqpamVdDy
2efw9B+Vx+Q2An83Ww7NoL0dF4rPa+yV6D4GO32RydwoVuzqF/ieEnwIdTDZuMO7GPPqqr69mYCo
kOWKp3dSlaZ9cYmLOEiRicKi4CcgYpSxECDXzuBRxOaq57gluxCDiMNUcW64Vpvan7uISK3cUGsY
lpyts55nHuI9n8NcJL83Wb95M/iv0dm56HoHk9BrmSCD6vEMmS//INhDyumSLuFDpI0bDd3sfPdZ
ehZJZp9ZRKRF2qZZIjFeFRoI8+164v5h9XkaPBVG0oo+a8Y9mK1NPpa4jK2+yA4HNiETxWaHhzge
g0/vh3+mnl3+RQ0c5Uner2ywhHGG8C7UKJUcQ8AhMM9qIRi9m8vxvhNLQfbii7PkCq6vpK5y0LJb
5BRWPDZ4/uSowcUJkqE7hlq+2pMJ50iKXDKfu2JD90MMBnlyTRXeAZNwFk8FbIEvgZgSUpMPzMEc
gyX0QaXiV7c9DApoy6mL5Xo32BiGWZM8foJqslbgL+rAuqkoaj5cbUXIDLzMwODgTCHr0vaW6C7g
iuC2rQICQPJNj81lg9eCZzAO4HlLjk1hAWShG7Iz/Xz2Ncwof1WCRqTfuA0Rldpclzq81nLJ8/nQ
kMXEbauBwxTgRGoWk43Qx7YyfRZUzuE1iLfA0l+bm0gXh9ql7TzOcJF0tcgk3hqOUcscizyooHQH
8therJIQBmtZLSqI61hSvVN2WkDg6zOI8lA3nGp/gIUII5wXaFauFtkOUedfuJxWAqZHpdr2Vgjo
qz4sB3N8ZTQ2Q3F6CUiUfjs5+kMeqIEv0c3SbXuKzpKHv4CLj0zarwJ5g7hDeQFdDct4VwTD/VEh
ewwL/lh6OMhTMsyPOVcEiKZC4k/Bvv+eEVlGiUThMQI82ao8xXTr40qHwnsyeeSR9oybbZuxheuv
FiGrJIFCTFHyNCzobJgL5NiX0L0k/Cob/vBCHvX3406bZ7Q3Q4kpEObcdyO58SrSTv7a6XoXwa/c
CBEaJkcETGTHbUmmorRYPgdNOyqG6C9ANiU8RBfb22/rsBFJX1rOhZwFsxgdyKT8fehfZ/wezosJ
3fHUAUusp7PRL3jyeqYXu3duKwaUs7m29KmRO4Ngja6YU68mx/osoSj4tcJ9gXNnEJe7scskTyb1
/9VmEc2N4m3J3WV436GjdtXgKAZgN/C/mNqSXoMK1ZkWi1fJmMtZzScEea9QGWp6YAAIych/9H4Q
KZ9IpbdnQYPGV33HhfJb0aOG2WpN88foA8Tc9EqWEj9B9EmRaXRKTOa7C9cAUXbu1HrRFydXn4e6
AZZ3bChiQAn5fgDv4QBrYFH6GVZrskhcRyMRKAFTJ+qPBAx4suRSoPumANRf6LWfq92ZmNDj8KVo
OmSmWzAQGOSsdiFZE0784acjkFZDUOG/vGPjVcimcSZ920tZxfGarP5MP5oFfsMyvZ2iWMJq5vDp
nmPx3MW82++OLfVJB3SZ6+fsUng8u8aDEdTRf+7ooN0DkMb1svo0EtQynEkNOLG+ImbuOVYzUetT
iV/Xrsr6828nixzZMULhiHnqauQy/dvkwpvSwVeXKTn+dGlHKHCxZpudoNWLlIPy05S4Tz1EElNP
Pe3IU50lBZLHeV1kAWon1mHQPQfebnFo5B95eUFKogk5N9bC7piLfK0bO0541ItU+MQhB2ArYuWB
mCGTUb2v3GA6sj4C+uwczE05Brsh+WGZ3uQ4Ax4nXaHjpWUY1peUiNtS25Mqx0/Gwk8MQ/wxhsTO
Axi508WUiYGymBFK8t5uIaVanRJZDY5x7USrnqCsOOWW1XrDuhJIsD7778c2D957TJ4yEwOTzaKl
peonPJNgTy8pdFTVhgTVbq/ERNu1FdU4eJpZQtqcpajtWQvGNM30s5fetmOG+L4Z+/bz80Zhziru
Lm/xCR7qwm9Z1PwNNWpWlaU8QRoqExbtmgRus5/6iNf6oKmcdyd+5RsBLvf3qHUII/i6gquPMbVM
PWPRnuhb/5tPL0uFVDbu1q0PzQTKSSSVwZDWGll2yDSjxJJLnNLMDMjJAyS52ARphHstxfZwRuUK
Kc8Tr+KJOyKCZyMgIL7scw1N+Q2o+JPQBrAkfWPTxfCX+2SVFLWeHf1wz/soYg2Ozwb0ndsgJKv4
ZuCxStXpPO422fkxp8hfGH5O04mFe/zAfIc4xIevNE+edHor/9+fmUHcjcGKcx8JivVleOTRUGYF
NJrBStO+LnKzvh0p6d2qbi26vyhDEuE1k/aXRycymepB82Xuuo9h4xLL1snmawjY5R3PM1ru6yk6
eewlIQYs5tXEd75SPn4IZ/HHiZnr5z9wL/jXAkBd4Jsd6qQzkzTZc1frx1kaZLhW7uVShnSZ3o2E
8EjkYLCZFTx433Cf+Ua56oeVjb3fbDHlA3ZqlmeBLR7OiTErEztTsam2rbW035K6Q5YAtFXMSK+i
xKxLvULj8XeYe2TTVA5NhGPfSjuIb/uFGL2GC6+eJm5BwTD4J3C0mFIOTnmcBXHBNi/jIkT8oymq
dlyR+U37OB1g/uZjSRapaNHfOVPCVnf6u67gbzAJeLCiwfJDeFmUMqc4Be8nXkGPY8UelAvUXWJw
SxABeRpJQ7RbxujVrrESImfvrrqCOLeneFxWx6ogasZjZsP43FXJcQmF1+iB85ONi31rEiwv8sYz
WDEiJdJlTPC9r/EqZVEtMfQLzNWR9qa90ULCldJ/Ci2Z0QuPGrvlstOgpqTf/HdOhhHKbG/l5S3z
g02CNj/Y1zpumXuqzJCpfGwszdRlESH1rqDIPcfzSWbF/HKwRxXKEuojs+lTTSFCb/49WZKnA1Ox
G2/CHs/rBSLIfkAEQIY0cdog30OvxzqFTd3KgUoOrkYdKrq3SJ7vbdcylADuUQ7IB7Haa5FADhyn
oW9y9PbJmWiNO/hrpfHU1Tvo9dGLWdczBVmh5zGzwu0R1Z/oCbwS7HXfqpJUraImBszE2Kycdt4W
GLDQc+EfUszeYQoAyLLi4Fagd7FxSrYO7QvpHojv6/7RNUK+Oa5F2YHco4AH/eeL+rzfAn8YcXd2
13l0dSR8YUpGTog7+7dOFi+shW5AtjO8ex1i0z/R5iy89MOkUXqvBOpWzNafTNDFJyyTm85WeZkt
ytRDCdQS4v1u0VqqsztPUz2LECHB8G8ZJKsW6gayuS9CawPkdtMtlNBGyamfvuRLB0kYzuDEXTQA
+v0s08mH34lYzmqCodEGxCPXazMY9DmY7DpRCj6/khd8ytDJzB8iwYc41wIa1cfNwJ+m+xE6u3Gg
xanGoV3d/FNJjJUW44fgAIwA2ej+cKdn5QcSH/7T97eEeXWyeZ6kwDwuzUwx/vhtESPPWHPxBJ/w
BeGnR4Vfh83eAF3nfDFsksybqmeCAjIfqaQdX7b8NgZszjW6/DrzAoagblfwfbOppH3sr/nGTTnA
w1EuD1TER3RGgjVu+ow2Qjo4Y4dMllLlrmg36pXKp+xr67p+lPoCGj4SRmwV7Y5lqVMWc6ukqTvB
3c8bXcJPQxGifDxbQUBin6NFaPLMYS0s0ienHSScvTWZWo0KGMBu6QDf2gR9T+GsEkfNs21C3cF+
A7Y4M7U3pIJ5VwmV8y5V1dglQX/5Rhc7gqbOoz2xj/XsXjlIsWhL22qdv53i1WrKvpqOwILRqA+v
Y89ZmCwINbmKiZrf1gL+uzgFzSc1DCNMO0f526EbMVmpVvraCGxs1IzKdIqPSlzn8WAEZeLcck2P
a0bCkVzuCz1+wbiTB4U1Iu3S+9TGxDtveIxo2YsGYyclLUwzBQaHwSYz8QilThVzQXf993/8wnYE
Iuw0AFmWSVAVkSXpBDtep5Lfv5mDYMwxkRULYAb7oLjKGR9r4scows4blSOvfCNCRgh/1WFZQ19x
3h4vOn5cP4uU9Hh8IVfIy56Biw2vS+OZzgroFPab/LD76TmM0+z4trzK61yh5kRrHQP2Xk37OVJy
0UMYp208uA7wueM2pzkZrb7+t/gcVfNDpp91IkRcvQ8ufhWHCznVARjX0viA3kV97a8Neod+Tn0w
PGObpbBz9DB9xoGW5/IqXvwcUEYJ85A8Sai5FKQZTEJVfxizj7wQ0ssg05edV27EQ+fI1PSpE9pm
qDq/8j5S7GN1ICR/ml5TOagi6EF3YxBgAQwdkQP7iHkVB+o8iLM+ra7iMAkuZOyem9Fve1cO3bFR
sF0ag9+AvBI1jUIy6lJenwms3gTI/7qo4I35DZ8htI0D7OQ4J6qKhl4JuWkbwEid0GTCYGwsKTB5
6GvSbSOECLazQrYM721g59cr1dImbnzEoKOmOXqsleBJKIY1ASYaLsu7d6GvipSk+wR2ZCZGIK4j
+4Vqu4SWHDNjqFSQFYvxP6y5yTDOe2YxHNgZ0ybhTW9fHG/XV7j5lzfZ/xQ2c4A3mEiygWKGfOMC
8W4YunLv552iW8F8KWK2gcF4H0EKNNRR2wTDv8yHRflVhfdjGzlp67KIc2G2mMg7qN2U2HUesNta
AI12bkqDDUBopGsFIy7EZh41Zu5kROi9yHe8VzGrlx3h3smKB793YhDCU10hPR33/dd/YBzNcWkA
RqZAUMNEWaI9sv0M4bh+YjqxXkheYsa1hR+mCK7o/A7yqNDCV7oce3KsomSrQ5ezWtZQpiz6kKsU
DIOIlGHW+3slzhS7LlbU3hlBTTjFHgA/WDYBK/YkrAdBYkkiWUTRsz8hq7FM5hRSbYIo8afI/idb
NjPv2dOSgk10pgaKvBl1aOUmWNm76ub6rCTv9em3BsCopAdPczQvoqmFy3iYpEfAxoxV6KmqdO8+
u/V8q+cWmYeYL6oPITCCUEyEt6v2N+H3YXXP9B5Ohwz4UmjwuNnMNbetjpMXPqO2UCS768T4gh51
VTMRIUEMtdvYiOuzYJj1s3J43L3Z9H/KcbdfNpqks7cXrmNMrvgGxq1UAxJYOahVDDQZHjdVlUVZ
TwW2w4+QshM+5pVoAAPlu/DhjrXnfY0QhkMzq29gjbVw3O6R14D7dD3Y9EV4TwGdHexpamMFaZDJ
9gjijc7xqhUKPeu26Zc0uW0mmp8g0/Z2kN2eUhSedOW3Y9S6gsa7bXEOvdFSE5Ml9jsyB3RuPRap
6nSE9RKpW8UuIpdFkEbZ36a9sIz7EsIqVfOqq0pUfAv1/8Tcv6GepUruaKenuCo70o5GcCEEER/Q
hfDMJoWN+z381ZI9ll6nCHI5J+hK9ox/vSZgdG0TxyWmfdl4RzYwMYTz7FP0I5h5P0vBZHUtnwsG
Em/cQCSK2BUZA45gepa7I61zcAFBAhwPb45OK10cdPEKiHszUHZr+pC2x7niS+fw8qSVfORa79qk
+jib71kd2VFvoScvnxzLvg5P9cSq5zzIz9k8zIc2ZSdouqJU0mZnTVLpMTr6eqPr9r7WwnlxIMyX
bPzpzzvcGLCGpQJjSYv+yDXCTAivT4rxu07KIypvk7hUSbBtkvz6hHRcmbYLRkWLBSYedieonlPH
F7a0cCFnN5NsVwnWlj+m4Bi2pnCa8mWKy6q3fy9OIXN4Gb9drJRC4AMHFhEG2xEmaw8+bjJnn91K
KKLMcFCPJzknRY5GPMEocblY7YubksqAofDddJka0DYtQtbv6mcNLvebYarM+0Ob2BcYORrCBnMV
gWGgAakgZEXEs+jUokRKhPVzxS82oTcjbrpYi3r+Gl579iP7jV59c4Nwcy4sstAmOJhUpmSI8MVp
JstNlKO191VAUSOyctv5peqU8KWygm16pLX9k9SC/KFkI1oWb/FHmxbEfzIfVgFT+OS8bwvHDFDw
I4IkhDkhuCfiluAnwQG8N8SgoZzSH7tIgT/iku7aBr+mV+ZE35x77MH1nReyCTh5TtTk6WNnd7ul
3VZzP1D3UTd7dzKjAf/LC5XhZ/9jzvyJ7OU/5abdy5zWAymiM9UnlqqcaKj4qIa6MxMuil7zyVyw
wTOyMXcXmjIzwNaxDA8hu4X47WCvtLTF5zgilhOWK8siKyF9KCA/PEbIgyj5Nrfn8Q0/8VuQEHSk
IacKeZapbCvDg4i3PPJ91MZ4DV2Og/LzWbWryTkpWVh1OSFiUQomLNi0h9gomWSjtyxPs51SMJ33
a4th0B0d0kANXo9PmQONP/vblzNENwu3R+vcelw/SAgXpIc24qwLrjX1Y59N18QZ/rz7cVbkxsu/
R0Bp2ym8e08sNj/iHWarZOs9bPf2FeCWfG4CIR58K6Bmj/vqC5eWm6aetINwlmSTMkBTCyaxmiFU
K8LHftQ+6MF1KuMm4X6PISXije7+XfNHUHGG2nTaz+etfu3h9Jg6O0wqmK54JTXT8TMADJgG8KrH
hBPFT4EOnBIZJW1T9Idwqu+Qd3z/Vpg13s1LLR63DN5LCbwXsFRh/Pyn4uU86VVOec1Jxixwlic0
3TiHU9jgvGh1JU7k7jcYVXtpwgEx5wqG4MvG9PA+TQJAOFCqhIF/N/kccagTokQhHeKV/PegBVDk
OhVgE3rZtfTtq/0oEPqq392cpJLjgQwVeJc9Q0xWgzgt5+XBr8ke4vd1IQ95v9/ZLATuaSsTvylV
k7ymuvhR/ktXzubvc5SdpEN58+UfKmdWIC7U5F7r7RwHctZumbgGAhympcWGQ4+0WtB14jAmqEsM
3iNodntsLOiytvgVohO86nSlU9ENbUgJ/4EA7ujZfUsZAZbeUHHnKizdxiN6JRGEv7tmlZSmCbUo
LSWGqjdFI9NN+fWzTEwkSf9wCAFbYLZgcDltoS4+7i3A9rjJmcCIAEG38Uy5cd0Pw5WYgC76A9ye
7NTm1CSBb6n0MgMSe2boc95tDfyEw2mgz21DIkyJoYiCLZOzKidn4xgxBmAnIwF8Ikii+HVJyiYK
v0O0aYv0S8K4zv0Jhsyk2vSmExyUGLP1tBUX2QNukPnPDBLI4haEg7xg/Fv/JY5JmwzCer9M89fG
HAh7Ed/mJKp0wkI4oTw6mr1UI6K78mWDgc3j5hkoRcl+4FhRAHGySd/7/d2sMnavFqhQltnfMrW8
/yvkciSb1w8remRZ/094oQnhk0d9rRc+Dn5j7E1mENpPsY+MiCvPsJol7E45xedBNKae4nP6+FZb
Mvkvl2/UXkookjT9MMNvqmiaFzQZDyhoPf7Z+R4wYeBHF3d7DGSfhd+Jq8q2/deN5OT/rMt5a3Dq
nUtuMes1boPQL43KJxUsYE7WM8ovxkuJwbCo8pd/P4C0F6wDfAGzrlhLL0Y3+EqBukpVgLPRoyXv
P1JJoTSWvtUnk8fmplLnIYggyuoC3dp5zKF6AwkGkakIbBolQ0atB8Shx+3LYbC7Dh6VCj1oy838
GC6vA6CPa/GIo97hv8gZLp/Sd3B2EVdmfmyClTY3C1ItftJfKFLdNT//43BTaDEVmymuVj0LeVsy
mO7ycliPluWMKaupYDSQqLWImQpNqvSg6Wvf+SKT0bEhbY6uB7GJFAnNWOOg9TqLLg+vAwAZslqj
txok6S5f3FosgX2pm/unvRtFVAhOFwa0J/8iANHoPH9mUbhsQ4PRwMveiL8D77NUnsTPlPpIj0vh
CXlAM60Dfg4EofeRpzuKXdi7zfaoLmc2ueITCntV3oRZE5xj11fCKZih9FIZO2HVuUeikPByqgpB
+wUOQFsPxjhPJCOx7NJXBFKOfwZs5hTCEMtVidmIggLyLEm/UUuUySV/ew8ttSPZg6I74BtSRxeI
xIlNEx3pwtPOAaX7Us4TRuqwczBHMf2LfMh3g9ncSxPYbna5UhWbSK/UHmEe4xKO59+nhlntk5B6
bGH/HcMXHoqOM4PEm0ow9YReSQqzLbB7rBnRMXec97UNY8mcPjMlJBqUf5IOJZSAq8sigx7069JX
kCiyvQjKTWMZQyISpQMjab8JC59k4Q7xkaHBg14g7eRuqK5HfsJfT79dLgdd1yXh/RRhC0YejBj8
V/XCorMZqimGXZ4LzTvt5V3O6IKIF1KzkTBFCT3dbjXlOE6HvbjFj/GX9S4PK8MDitNq8Lw7AojQ
e4Qni4WNkWVlcSY5QSDfISheona09GtPy0zptG7uBgudd8q4VK0dhgmp8DtoKNiCbzx9cp/kDanC
Rq9lbFk8qvdmsLVMyR1JuI0fLbQuP+8ByI/GfMR2AW5iv05Velz3naddJemm4URdhS9D9BL+ce0B
hioWuLnUJXZ7GLFFv3yt8beLdTONgqodF2Pi755G5ktvrH9E7sEGZpV0+lSxuGQGObkcuJJJ3NOa
KF7EjDRi1lrBl/uzYWWAw+TqERNH/jO60xURO0czdUQW3Jf5x+b0EYiRWbeONNZeUalj3H9Zc5Fv
hzOmZoC1od00faZIPxGeXgZ/NNHZHa/Hn+E5M7N0ty11+P7Fq/0s2lxLbalXiOFPHjTxG1g4y8de
f8qEkeS5MZyXqTj6LUbKuckPfibIPISJ9BpTPvWGMtrioU4SLzZROqcOJfZCSV1lcUW/LsLJk7j3
2LuOSWIjsXmyBQK1+/Dgcj7gVfGu+s1DzGO3Ijv/V6pGriDt7cvMMWSUO/Gqr8mLV0JwzyzE5VlW
AABA0sEMJJ5sOzXV74Q1Ho6J8mUKhxphbspmZ77rQs1fp3WUdxsiIHFMlqtvtEX/WJOcFhPu9T9p
gcoS8+1OsKQ78PwfRRe8+j58GyjrGFsGSsHbNfW2E2qYhPLYQKQP27MTgiqg2GMXLVUFRvTfP7t/
fmZjbX8E2vjIHkQ5Vf52ukxy8FUQLomU23li4Ncwk84SipZ6bF1IkoPSXlj27aMk6D+OpSB6qP/8
iMhfZ70kZV53AW09RuVNl0kUEf6qEtAZ1oJ1uTdPyxAvgbb0Ovi7hw2gfmpypcX+CAByA1LN9THR
kXqu+nEpskZXZkWszM8E+QMsGaolGXsfZ0eXEJEITgYD4ifHNoCoScRKjdN/yJlTE2HBpmU7pczv
GiBP0waSunarDOFl31IYvmj1qbyFzQUd+cAUwi8BzXe92Ga2D23OtqHPFpfSLObyKnb9Zftv3VNS
HNDFFBih7VAcGTcfFdqIdrfUj/nu6fOXmuPq5v2HSAJ44m3bsVjfmOcN6q3hbcFJZNV0KWibUlpV
LcO2WWOjJVm7LBOcYXLCJf9Rir3V1Ip2YAoFYdh+Pl2R9hd04H3euYZSQv9xe9m5/75SiaFjgSRU
ICUoznlTYefBGIo/YMKPWrT7zECaLj5eXY38rOBOEqzZBBIV/Stq8Zu2DXgL0MJKGUtt16DyrK3m
ZzM2S4d1sz6C/j2X5QJzkjbb3+gevQ0RTyg1IcnrZmIevuwhhVZG/j/EjaBgdT9g9nuFnBr9BmJh
/avLNH/JkWoaqzXo5NlnJ8HYasltVXU5Nf7j/6F4r5Sz8XlmdoWf1KfXqzlAvOy3sn58vIIH0m7n
s7XlQH1ZT8Py+wpblRnBe1wBS1xtjsNgCkJEwY5S33GE4NyUDsEajX3rYZAuXzhVyxwD1c1x4x7z
Ukc0XP9woEvA/Wj6X3OFWvOiB82efmdlJN+92U0uJ/e8sXU4HMGNhsq3GpGbhjdyPTA4G6MiWUj1
8hyhwGbaOmAF+iPjlfPOLnv4LW0iNLxuFsj+E7aHh0vyVA1/OFLyLZdmDCEf403WFiiiTqd4RlL0
KdLEjmSxA2NgL50i/aGAb7mSKwrM7eVNOtr4IlPRNM7DEdbt5rgKEB1voiWsVMA0odxdY65wpVp/
C3IyqjpNS0yONSITfwS2r760ebOVUdu5tQ5i16JelKlAEdMSRMFsDNXYj7+Xcu8kptbhkWOrDq+S
RQkzl7esjTbZ1hGlFVJgtmTIYyzznPVZs8ON/f2oOyxkp7Or32qY7ZKnZ3J1RsQ2dKfR1jiYLRu5
onaBtEnF1ynCPQt5W3KiSC3l9PidGMaU0kiY8ndawSkaFaIWCCBS1n7te29zQihaokIx5shjEz/C
8B/EnoRc7eEZSLi/VB63Q1c4KWjJxylBpNrxS/v9nSz8cCgGeIp8alLurpMp7ywn21HaDnngc/4t
nncZbs5uZ46sO6KhFSxiMaTNz1w7C+6EXcBO6uyRhvk+D6X06OfEAWPzQ3amA8HOp2KWjn0OiL/1
Hi9zF8Nsffz+0NxOTxu1t7kRPin0jJOojvesnNdYe651QzasECgqUGjdLKwkXXBIVjp5/gSsKzKS
P2LWKIrwXuXRMz226IHFT56wLg++u2GZxDgtbUGkFBqbBhnxFuDiXRMuaNJKmpJondE5Dtrk3msF
qhTcp1NwmDgOZIKy+MP67QV+b54ah7eZqlsPsBhHQrvY9sqVdokJYwwqMpNDtz2HohQiyWea2VPj
0m12qEonX6Qt5tG96rWL187Ksq2NHsz0ivvMgdK018ATt5I5gDiWn3fGiZfqIIEtZ7vE8adu6o6p
fO9/QU1iXfuC/vGNEfJGvxSGTSHton1Yj1GhZLN75B1ShBjDTIJ+C0v1jHBLKHZNhnnkUegzC8YL
hC7yLfX7J5wDjdByKBGNEFxo04Op87367rSLZn9hD4h9+l7djmRqrsArimyt+BX1qhuEea7tiNI9
0o3EczBIlJYg9Wmw7HFBLazYupNqbsPnG9Ismx5uCxXWbL/lx/vezramB50b/NUSOWAOCixGeums
2sxp2xAogKdEtF6vCRLZ1Vd42bU6431UTUwV2Jqg8AIbBhereyi68qhpXKNQgS6wmrC1Hw8pS6jg
oLbR2MF3wtY6zmGifWY4Y7rq8v69mQqeBQSlCDgYv3YnyfnHUm20kW3e71fcM5B3e9nf0hFJrMaa
z0ZMGnhGrStUzyPbgVYjVItmMhgOsTefpjX6hO4ibrgxZfH27D9qwlOBFGXVCF+FoVK0KrRMWKWJ
hpKcRwWzRt7BNmOaRfTwwd4+2oAqHvbHu11ClL/UHe99UG+JslVGXLBstB3cP2iko7HwvTVWvw/b
hs2g/gc7IMKDVsMlvmmzJdhyg0PCMBiGdsyuNuoPkvIRBfsHgAE5y3e6z6CFE4zxVeA0sPSrjc/w
FBLQEEK4mFKLpnNN15/gdMTs9OAflNhLAPJWIvWtmKj4lHw0an8MajTywvvQhthkEVmrGiXhbmv/
WqD6+9DzdjgfVKpzwxhPKBVjMLlvkr55ecaEFIm5+H6iQvqIUqHI7cQVvwIXjq3uKPDpBbDdv/bB
aV/bXSK7M6jp6zd75gUoYzaGgDjEQ56DuxDFC8mKY+rhBbfxbpVxP1y4GZoM5i4WOPhAviXBUnDT
zn5KXh1yR3YJiMvCUCXb11W1UaiJ88gMVBXYx6uVKG7QK8DURpVPfeIKc1cHgNakFYiF5FiZScNn
WukJrOx4xl1JjUE3W/l5ugJXuhD50Myj/gcnwdkOCZDsy9TV6f/gzhU4QFZgGMlA7T/9fMhwJVbd
CYj5e29BrbZkNWbFjfse1h8X4i9xtnNrO9ydA/k9sN33HNnPr0ZvViLZ03E3QSt5X7GNh28Z+3rX
tBOnjTYzFZK65NLw4+4xNqFE3sal2CEtSGXqya6I+L7NfK0xnEQNgMqfOyaDMNhfYyBTLfp62lsG
iLjkWQ7xYlv9X/IHIwBbUv9UQ+dvFaBTE/t679Xqcn6IQmWWoNUqN1zxk/LfQyxx6+Za72UMVSm/
PO/+jH25hXtOxOvjwsEom6fHrUSIi8r7iiOULYuuTCZGR0Z72t/dE8CY6/BTkyBxJIaDEC5OpbAq
T63iHNqt0uBforGrdbIV06Ck1dKcpMYxDsyxlQD1TuIYKcfBp8ff4DvZPFaNartVomelSFOQSzQ1
os3bMomF/ug9pqkIzySVAuceMkT2e4MsM2a6Kqg51TTFylKIWszIS//SKgHciPcjnJIWrXVnLhf/
ddobIpbo5hISIkMya/Ks8SZ0+tq0F0WaSQZPgmBQqo5tYmP+DKN0QGBJFlaqfk8OrPcnHCqhKt9R
Go5w9r2V11pchSmz19tjc4kTa4EmQoe3IPuT+Jmv/La61XsNCYxpR4IapkEkuGGN6zYcrf1VnfFW
x9MJNCoCFhJt9NWqrb7whkx3ATADrltqfCN0j5rXZPiBF6PHx78HMI8laq25Q9yidgWzooq/hC7w
Vnc08VZnc8N9YxRAewNKLnSRFDxf2z4Kr/5O0fx2x8MAfI610AZLhbwFoh4ub93/9Sv6xtzfoMtA
9g+CBM/kFURgkhx1bWUGN6cIxWgRGWskcZDnAHCyP7hfce6PjwRimqLQf/MdQ49lHMG+erEOpob4
W1Pidr0kdQX2c1PQ3PuyC+yo5gPaSd3WAYJiCF2P6Kw2IrhhS1EGv9ZUClfY2Rvn+Gwy84LJ+cAW
B5rRa2fWQ4CrJHeyGm1bQECg5H8iRprFcO6ijFHafNdDkyIOkXywIYj/U+VNRSjpVLT4t8w0VTqm
oY16bvf7BN/au9KZrjIq9s1VrgLeOXYI05z+QJgoFGns67oEsFUnK0MKTh5tgWKLl6srElOhuZc0
lpR+i4W6hQHdTV1PyrLK1LSVjjawqMslIkDg5cqaYFPF/Fd7ZJiHn8BWnQkZr+ZLO5NemJEvN74X
1fZoiQyW8HAPkniAytlGGCbWr/bAeUzEgl2GFK15GXIrz6e9A6JTsJb7HDl7x3faGNPIzykwLmuD
R3mGmwIjeLR0oiWck6yUX3q3R998EhAh5A3Q+5/zm7CbaK8bYY/QUBVv2jxmv9YGHFnVbifviTVa
0/l+rNfsKs7n67S7GMMnHCzNHPd66j8oH2RqZGAuGh2jwg28tNPXq0FgKel5F9ztNNQzE61BnStr
gO91lJou2grLb1bJ4q9d04buDu1Ncftv07lWZKeMjBSgBify7PyI/IZmct+4+FYoYA/aYy3JDY3n
emzHvI6JEaisBc0KyUOBMlBpGDS6kE0JYySeWX6vrLwaWtV3o3YTZ+NGwz2vdV0jwdgFnwbrWh6E
LKkFdiyy8KBdZgJ8Nvsq3W9fJaugRAAls2VrZ1uitU7+C/TVz2IaigmVTtQ3J+6EzsoFpGHxRJYq
jazPu8+08wjgUBF/I+/YE1uSRppZwnx7pPmUI2qq1ICwa78M2V+z6jEC1eA3eIk3GRlBqv0vw7Gr
1kvnukR0o7CTUg5/6Ykck1f0XMPUUi0y9inF+5BJzRsY+et7sBv3Wfc3eZRxkJVnDitkmVMKUOAm
6E1w9qzayRPZLSU5MAtIU0XC6avHiyJ4QuyvD4rWRgGKAMtg6gjEOWwTvagbmDdeWBZU19tlNuaN
mEQmGh38wqRRRzOcFWvc9AWH4Nb3kegYAZhP+vuj9nd+c20zMtry6VjYIkmZaDqAdS4vZIOpGPYl
GSBtTuQ5DRXLj6CPzjxirdEOClC31YlPV1xPX0liAcVLYrnt+iGYj/yrMdMlp3c8r5ma2M1yBDgA
LgkgD0Hp4U1/MRrVUF/8heU2VBC67R2H6eOliPRFHZdlG+7ZWlv7o+GVIzjwmq2DRWFAaLgDEggL
HLVoYoQLlg37illqzCyNkwp3dY4sz++qc7N0uzb6EEzl/SgqrlVS+RvID8cMXhpdzK70HdjiUIgn
OmeEQ1SIQmgoJkJrl55/UENjmLLUn9VaQlOybKKOW4RxcPe9nwsUNIHZXOJBfHJOKYsVzaiFO9ku
nS+UFN1Eb5mdtNwychNONNjz2SjaEUjHFyyiTC69OS8J5y+DpUhynJSO+aNs7Oe6NQKqCLfWpVvn
sdjbrK0Qaa3VGGyUlGjVcRBwmVCz7YIN6VxjBY8u74EPTj6m8wn/d8oP45s29Mi20HsacZYzlPu2
9K6NSlLnuZW5osZCJw8zan5T/z4ZonVEYaxCX9BTed9yOCAswHL3sYjRaWOlURJjZ9WOarh/a7++
Oiw3gZW5iykZ4RAntFhmSkQHdZzyEiuDkWW8yEsx0OVQZeKyeZqxu9CrTOGIfvTi1UkVzdvUBBP5
cDFPTEIu6TIuOJtu3vmBxzKYtUYs4trmc5ugozO9CaKHVpNKM/fatOBK9uik4pPhddd+F1oda0cn
hnEI0J9aLW4KDa5M1QqYVYl+R2xT4pQN4nJAP5e/ROyCXDfIC/FxI0n+K7mFiv21NuRmSfxuQqWS
ftrSKPqG23o71RHUBl1PRz81Ii5g654jjj5MBnZn5oB4TtnHahGB3Eq0FbXgZUKwbGftAHMcI84D
1rjeuWYlRk4RnVTCYZJczyzG9vvVB0inuw3K0WbS2bXkZSWS/PdSuanwuEdofSJkWfxIZPqit/wM
TXlgHktjXjUiVAhSwbqq+5iasLLmXhkIU1JuShI65TtiMmetosMUc0SWsxP4qjF9m4voLUESPjI0
5McYCQE5lGbefqgAjfmNvamD+L4BnvPmYqAdslAlQ12xvE3vKNUxVm0iPR2io+Ro5ZBnq2/ZkzbX
r5gvVAoZQhrEN998rkMVAaXPuxBNoYuqePph9C6TX6cgStILRRFZrx+1rM2inEaK0GWjC3WYkiN7
XHjXCxHz8sz7rE+XEOQ3MWkUaNgNH4FBIPtNmmtNbicBOzpMmQ18BjhscMNCFJCfBKBLfM3EApAT
Bg1BgnHoiNNoJkclLx77OxumRXFx7aKVrxyR2YkTUhCxchcDYsk/AhZiBkYdIK/TD/IzYzJXI8kX
1J7QdVHvqITy7sQ8k+zc5FLWtghkxEpxTO4M6v5uRjLN4K2H7ABRDGNyvMR031A8SBitJOL7XtLf
iLx0BQILnt3CXaF5QYVIuNZE0342LgrXHgNITWV5IRFbnEmnmTHa+buipNsYJQWwBCjwkDwTSqpu
cymWJ1IFva2lw6HXDyfSkrsCBS9wqZxfVvAJpeRK01c7GZFQAWVfjWkh2NVyaG0eE1vbVEy6P4OA
IBO4Wosg0B95m65IU+4l8W605O3MiRPDg/hfCDLimJUDotdcOOHVQB3fCcIVlXSqeETkMdoxCAu+
uZKMSsDr7d55cQJiCXTpNPP/9NgY2QZa4J18uwpTSfZpNEG8y1zNnMGsvRQOhpUkAealKknw+kvz
j1gOUc9j0l5uJC230yxwrdDK16/CQR94USa9hPcigCT9TREKnL922IDm3w2FiCLaZRRuX2cczqGO
QCEUBeDW69QUuzPA24cx8p11ZnF/d5p4oGY94I2RlY8Rsh8gmT0t6tQ/7EigQ/POqA2QW19h45zL
0B/VjOMadaZ89SkV5NghHbrzLFGY+bFM4T7KwkEa5ZtO8oVszqTephEvtBUSePRimd1oi4xDRNtg
LGuL4Fwf3puMcBRlTKHdB+W+cvFU0+RQvRJaRsgCSDY86/evoqNdh6gJN1jnYWhCPYq7hB0IelPp
pj3TMRDnqvFWxDKmPOWkhq4fkWZdwwqg652oJe+DOlzPsDuY37xc6C7ue1lNS/xx60hePbxIAeJQ
k9spkv5CozMY7YJxG5Ag1Wu6rS1XhOOdk4IkOtb3MKLFR6q8Qspc4mKHqPaRHoYpdrioAIiKuWji
m6luF4QE62I3JcQUTzXdxXUz6qFyLQYkgvwXIvAjWvPreNSM/EQPxL1u2yRhN+cpnTMGpBsK5xLQ
oTT2iXJXcCxC1OORNoHZ4xPiERWRQUqJQlv49NX4mdz4xgLOao7hMwV66vT6Kw1vCcHJgdj/lhlJ
tm5j8rbp6tA0pw4iJdJXjC1v5VF2diJeyHiIDVe1ttQmziuNoyscnfNiXy/oOvKF3oYLQrH+C2bk
98k4oNdjBjEspSxrYqeIHNLN+AFqIfIF2v/9gYTwO34/t6Rb0qXfMepq50O/fYRL2wCih/VXt++4
z/BgBpsEvKtCSIg6RvOvxwGx2zcTDKkq94O6OqhQEvmD982fwYpDPn2wXUmrKs14x87fMPST8fVS
pKZXmPsX5sscYoOzxnGpEe3Qn6Ubjc6gU/yVubbEmi06QTwdQoBbS9H0wAhKVMwujAMmzcDdEFr7
9nV/mmv3rmnz6Zs/Q3dAh4KmzVmIYhqPXZXBuwib80KcGWVi7hNxmc2eGF3ZqUnGirrQ17L5WM/C
XbMHblwAhG8zYNZsyGTDksgej5oZTIk+x0l3ae5DEdTattmd6wa93RyCWaCkTk3CS2inhUZcVNLO
vNPNrloRZG/3WaCuOZQhA9xsa3fKV9R1JMgPWBJx14SXdKplw6J7zDDXFymq2XMAJ9qfSix2XMqD
M2P08Eo4P0iBBuYN1WTDt4FIeLY3xYXiRbXQaRpS6foV0O867ikdQ59GXRbbLOwYAAfFTMzmyHY6
QL0VssCUvzgWYa7YvuyPBaDTrfnQib7S6V5eptZ7HGconlDExN3YT5VoSdteNQUtYnBSJb/uS+3+
47HeL2KjOH1xei+Rm5dIfJIjhTjHgBIn1rgQxriiV2Sv/C6lpQQdkmIEbk4x8FZz/Tkmk23Q3FR7
CcUjXjJ/woOgSDkCRRnlrKbG2m7saArJh5zoHnbde4y3zZ21z534UtDWGmf8carQ/DSy8ZJU6+lI
h/w0s9djcgxM/TPANyPW01jBdcLuwYfqIzEYrHJFqbDdb5OoRyHSF083DNVMXedMAA2tQFx007WB
4gGqG//fGuO0tgL6W9LaX358mTtZGRrzILslS2BDtMAGtgLnHtcWUf+YSzA10OT0NAThNIltTJOB
Qi5Zkz5xg/zG800klkyYHL4JWBJhTzsRlWJpqSneR7LtdAIY5uzfC2X3DrUj/hlqnLd498bjKpkF
lBAHS5DaL0SXw2jW6zFZKovF4zLgUKVKCcAq/93ay/WGbmM4ZzMGuMaIXVPJGJuar/f/ywqFmLyu
oTwAeV6oTOt+VJKWiWR5dVTdGKLaN906ormPD9b78EZA05W6B5QEB1YDzABOIig79nKlEqh5w9th
ztE29ig8Ny4TIM3PVVEcbdUqAYdM9YUZ211ZDC2KcGJ6rVTc5Fg1mkPibHJrI6r+OooYbbaofaS7
vOBOEIyNyKMnB3g9yf0BF5fctGijhQ1fHZ4wy52iBgmTbZx+3TT1q5HEax16NMc51Hp93GbwGc1+
swE00id1zNpMylLe+QP4WISmKQ9xK8zr/fiSOJEn7E6AcrVjLni5NdNoToupgrKrKpfbB/r7DVKn
s7+6AoIzoSzZuHylTeZVI6+3jjdyP8I4EFMYR7FVqYFmK/+19xJsQ7Jdmtz14oJaVqt6X6naj3xj
HB6W2WVHltny8Eqv8gcAKuVOSQoiNsH1Z0hk4zZ/AcmOohUiU+/y6SIsV5+fDeA9kMShfeCSv/fw
9LnJ/g8Xmd6g4hYsFnqEeodnzI62IiHu3wrfkokQUbsL2w1YI6S9xh0b9352l78KXDurRauIRfXW
tQo99JDuLSgcjRpxPnV/ElcQA58uMz9/U6gSB+cYhDY4iZzP2Rk9+e2vo0S0Ct6JAz2T7dihaE2v
+V1vc/gzIwaMuRhbBHwqMU6Ral2DUK0V3QRYjO74Yhvju7XUq4HtZGNh5EkxEob3ZZR99eQF36Bw
XLUy54thfTEG9W4Y5IXp8QnGvg1a4l86UHerJC9jgS1hXly86+jQqoI+GbE/lL0tWEVJeE8H1sOo
b3HJBYgciDc9z/4J0jN8K/fhsfIEgr1ZJCnBuuS2DrHZAbQ6jj3I7FnDxuPWpuv6ebBmej/1FtsH
tHCGwfkqfeOVzYqHamEWGskk1PuXhf24iYMtXcI1AYO68mFDI9gtK+AIGIvSvJ/Wg8Av7puQDjzu
T9ZnnAIpcOFECisdNxcQyLKnGtI5HmGuRDTpUt7n2K+ogkVgVL9xyomECKdOW7DUFreISoF3UWht
GH0MxwsCfWyAhiHFcQT/0PTgEet7s9VvnYJwuBa5T4FxI9OZ5ixWs7khD0DvnIjigLfEjFd0eRdc
56UzKZWE+Rb61rM/QpVnPQGoErPYznXEKS2u0QXTrl9pMiVyNvxk1U1k35xmW43y9gHSar5IksvO
RF2YhWqYBhL5aGS6glxHLgLnTx/omX7DMgEKze6fVwkhNHAyioENW7A+WYvK76NBsyW4AoGT9e06
L4QDajPwM8TSgfFXRGuQehgoMTqPoXCQCmsffzFIjDxU7Qm7qNyBnTCso+0lVA1lSGdNmR6zilF+
OIVrQdHSKOUELcQT1y/PL3QyIi63kp6xQSR6xUIwti7lxHa6vK3XvybwlRsepxuMK1a3yc5nGqjP
nYUDS09hb+5YjqweuczOqzV4VrC8eocJhiak0LhdkIGdDhtrW7PcQ2xOmFrMDw7KiB55C4T6rXQi
H8suL4TtrkBgEuVWiEKvplmxzZTQ1YO0c3SWh4F0HK/aBhxEycwF9Ssx70PFXyFHyPIRxrakFgqT
FSqBY3Df2uP56puwOEEq/jZW0eAo8EZKZBKixcTWjpqglo2m6OvB/OaWuOg3ZsCTJk1ur08/wO7k
Rfd7GzNkj5ObW4Im/cpLHlSBazwb4KGx28fuEFwusS7cc1qui6kf0u/mZm1Uax5okUavfPp7MskC
iuEaZmXJAe6UW4/TFYxbBdsuALmxbCPda9gMLLYCNOjLKppSchfOC5+tze173sN3UP2r0f9hDEtd
ovN4pyh/WVfylNoF+d+xhzZnqt9cs50y4UwVbSgrrDczuyepbT83IzcZYc6I3MwSVQZmXsNld6Qt
dYwxZePPMy18NgdYxyKbVlUHhbbMIp2D9eIs3MB9dpxPwNte0Epp+i5QLZD82VmPDW3wynDZZQw/
wT3+NU+ExmrCBlgFFjo/u67R/H38xxNYJFQWgtGBy3bJTqgwUr8uPqpficuiIFlFMISX5wqq5sY5
7CklAeP12g6u3jhrIbTBeVyeL7p5SWfyew8p9+/6M1zX7LE74Gege4DQ9cr5+oiN1aLzLDRsza6R
RWzv0Yqm3rXM2/ffbaLHy9FnSqyJAj/iKBa4b1rNhQfqIalaZzvnewEO8x57+itQt6wQpAmKO/S7
2qyElMI+H0znwoIH8uocZPTZyjDHzl140PUhLIu2KYK/hkBylXnwWJaw0LnJ4DHsPMyxf0Q7f6PI
Kuwv9IM5WC3NxbwFP30PzVVmriZNIMfcFlGIhNFcBEWF+BPSIspbrIA4LXVIsA6OhdpVvQ+u4tn6
edgn8wRuMkdSi27dEZpKiSRyZEEZvRBoPEWDRHxC3u7l7F3TC/WMbBhj/Zqfnm1GueLIo/C1ZWHt
SDDOz6KfBXCYJIQpuv9DrLxD2yixIc5KZKIJxIwB195WQd5BYST7CDjl75Raq2Hr+qrxMCpLKPM9
oDH1BgfjJp+RM+F5DiFyS1ITA4UZQgGWwLi2n8U+6KKYtiHl+ygD54lrGYGodWe8KOOh/H54pvB1
8z/0wojExBr75vau8sE6MK5m24Sr2a7F4BC+e/WmmwOtXGk+0yhIilCFEXur2mIJpxWMDpXKyQ70
95udVB6u2KpWEQXan1kk+mCrd3F/P8aJ6JCwJPUQFPTPK0jUzBhOnnU3x4FSaEMK3GAHd/Bsk6Uo
fNYrnPiL9f6+8CccVVNe4SS4DCHXxK5ocMUbTT4mFlnPXAUCMDuwT6mhQSr29q5Zuyerw1VnND7P
FD23/a50mtHhjigeRiYOCIOKtt5NRJyXtC0RkU7cb3O6wIUuu3UNvNI04CCmEwlw+eSQOcHzb+22
UJqYfqKy6lbOalLjxazmk6MmL2CUgTFMRSA19tJzwV4HQovkZOrthik/deKVA2MoMYs5A/H429DX
Zyo6zWbZJNORlFk6YX2+EohEk6acP2u2LotjyDUupfq20HVHgGhICLsF5u5vvcXfdCP3cqADxBjP
q2dryzSs46wrEAQGrWc+psxzFO13l9gEzDY8GYKBNGWL6w3Gycn/DUODxJ90mGlPSDJpAcsg8wQr
SMRZT66ROa6RLXmNPwAxkDv3MjQ/JY0kj5khCmBG2HSaMII/W2qIOebhoWxtZyEdHaLzhSFvuQJK
QTtaQ4l1wEpLKBCTUd0scUTK5gyPKQYtN8nrV4ezLY7/EPp9jANaBFkv6Yv4o5x081a6j1OJiF2N
85/pIiRoFeQCEgn9BCzxVBPiJRVbsk8TWv2MiVvssaqHrJqpQyNOJN3Z5OdQV/DSA2kGUk1H5Tpc
6yv8MxKjJjRWuUKVWMTEf4ZSniRTH7dotpJUBwWLfawDSw9EZUkfFlXXd34Vjc6GxeWG/ejbWvU+
GOEg7NjDAXLYdNtEDEKWAJcNeGWSjpJQ/H6Zhw7VWqrLo7xeitGsOt0N1No6Jj1tVa9wLLRdTIa+
+RBA4JrbyTwxGw31vqStFxDS6SKp4Zum6t4X5ah5La8kSD15dwS6s+7J3U+z1wsSv9z1jcZcKbQ7
ZZLKBXYhSAq9Chv/EBpMiVqrp043omH9g7vCN6BCMND4drq3VNgC4M+eVXSmXydZ9CTvThyiEnxN
m8UfpScNAK8b3PMDN+z6e/zF5LWOxO76Ae3ieOK3A6dmererWuIicOcj9QHBHsb7apZ5yGZCqkkW
dErmLz1EAI4ethXOzHjPPrm7IwDmFpx/xyeXAlsX/1bpR7WE5UlebdMq8z2osriTfVw8cpj5xTyk
WEX0mV5NvU0cKaib0DBvVSauCBEDDfangf40oZG4qXFg6/AISCmvA2KFjEYe3TUjO7pR59PBDtKs
MZ9d6geRDyozRpMEzslizp3j7h4Oja2bqaR7DQ4aWkNOQM/QTpNt1KpcSQP/1QrCvA6KE27zn2CN
veJ6NJuvdaNA3Ywn0DFFm+Q1k7mZrAyCZ5dHmAPPJSvW+k0Y2m3Uou3RdKHjgr9Se9qnlqY2B7yo
KRaldNI2D6kndhSzTiqNr/s2ItI7aetTMKJkHAsRb2rpQhx9TVAFcteD2tjHR7Nw9+PGkSn9Ct9b
HPhwXoJ8uA2UdH0W4jjFZMnL4N8xVR120abBGM8m+KoM9wgsd67qXJwjKmU/eZqXfT2SgoUU83xQ
MjsUez/ImzcjrwPlQx8XlvGEhncTSgvdGYVRcG46zbUrTnCwSncTR1YMmnhsitF8ZPqekRngWvim
arQd5r4da2P+4hPJoAMCn+WkkjRWjsBUyCMHonw7y1Z5VBFgFBVEH93EWXx6E4ugEAb0OqL/FPTC
WkRsVbCHPvgW1JCj7JFnqvWL1nEaCSMU+w37rr29bB18VidovvlI0iApETt1vZnGb7I3pbD1IvR3
INwpEtDULrh35XcAU7dMntKzVc0eCo8ld3r++ayeOi/gWKgLkO4PLtxq6jeqimOZJPcTNmYvF78T
tRAXIEzhj7KjRL2EdF+b6aBgr9RtBh7LtCR1cYnfGg3f1P2CAtvhQH4eyOcaCviRct17PV/CN+pe
W6vhjr2eJacPimIfCWt2hKd+zugh+3oXVynLj3PU4/CIXmKNH7WqbW68SOc7ljPuMh04JpHgOT06
+I+lXxP8tTpZCESe7tLBNo6dDiQDv037lzSCapabivBwJtgD9cfY48ZA3VimRTe1kdFQ7/r391qp
9CSNoY4uttDqG77gekEIrhpqp8llRoo5U8Z38OzkgMwOIZqX8Nr+QVVcPuB+RuLIlvROl7apAV9m
426G68SLK1ueUbn4fHndTOR6YAlpu0h5REtfZVAcCkQAz79DS0ZZZ72fwESHjmy8PI9Na+NMSfAi
qMk7ZpKwkLXUwYjwC6ItDmOj24W40PQpXKCsKC/vDs8eWcZgN9koChLIT7eZMKxsvcu4QNW00SLR
pi77EFjGBwoXsK6xE4AJZSdbp+aHjshifEMGRQUs9rpOY2lC+dbqtddEF3g+Ehv3ZLGAuoNFW40O
g2m6uxKzp64vXVekXl/fDO72KT0lwckX1nJ+TYN5z4GjIROR+KdcGitYVNBq8wpShD2QpjwxZRIq
XSNHgtSkz90/FZck7FfusANgmOY6BwiQZxNABKhhNzla6HqFUWkFezvGsmyRQp3KmMoINFH4BTP1
tHcjGu+nxhVLjuTOQmHM6PmA/wheE8Qn1AH7Yw85Jy8BtEj9UnxvNLQqk0x7IUPhJoO/GTHdbp9i
8ZXpQDvZ9i32DhtCmd3/LZ9EUuh79jtEGp3JYusFmjEccqdlqnHfFtyxvJV81o2t/Rsd9M7wlqLH
oIiFtFXOIRqKNKcyXTRoEw5SsnJOfjhRPk2HmpjAVLDHgDsiC1RzPypFVwAV4IcTeO90powkR9gR
ouws+10ruZQXAC7+qMau56tiXyKlgG4bbrrXvfHjXOHuhretI/pJkdZgTwwTznNFDY8t5hMm4V5U
VohXBpQaqaH9bC3vZ7JthgyZls4zHsrfM6U9lJiC8gCOBEsy8EGoi2O3NTnCBZIzRXYwTefic89D
QrYN+V010Ppudi+OwSGo03EkkqVHQjLmViTF9lndbMWbtCbm6I31Ij+92hiHCcuMgRTFTXZW/DUc
4Q2z1l8k32kAaBxPhQpMB/Ij0BXMdR2jb1zJOym6o9PkZbnJmFHlUQwv74DCPLaEnBljJk2FJysy
4d1MBySR03Xf7U9XxMJbOtlTO85px670N0QzhbyqlBhzYjf1rnjcav77DYA7unZzE5Khzf2dGB0B
IaGGDVUQFJ/z8PwiHJFywT91HRR8YWBlzmxQ3VIrUM8eVMFED7SL7tedf3L4lLw8OYyC42ub63Ex
ch1SmaDDd1CGnFgSq1QOmCvzQ8+dfVmP3o8FUrp/V9iIDLCFP8MLYxdFkqjiNHk5buMx20q0I45a
znzUjXMQi9kKFgyfuwiGMLq6RIx5M5xXavio3oaUmKqkfZaIxklLtGIs17vsTN+ii/dcYivSQvln
PY/CM53EXBnKCcLx+8E47fv7CnifW2pLmjNpp83Exe5TFI9g4CRf2/gs5XmpU6z+ho/Mp1VuI/VW
yoHAnh0rQOSNWwV99elm2E96kUiH3X78TsjzOrIjLtLRJ7SF9kN8FK20WoTRePNjMVdmjtNAjgsw
j/xcQ1wspp/Q1xkqKaoK0xAfk20lCM19d/Vi8mQXg8sRMkmnHdDo/HGn5/qtKuX938XgZQhkbVVA
8YHJo6UoyINoOS+ldNCJtPzF1wuScu/U+bwlNq3fmFdCkiTO7UBB7p2mOmon2cHpHFZ8iEl8F/YH
nFwnlhGBtTacsW6URdY/HJ/PFAQ8D8To0dW4TDANVqL31IG/pUF6MUqrvnRkjnrj4N272fAN08Sw
EUip6o6O2mmWnYiHEi5Wepcmb7JUFrjtmW/pOFa1yHemi5LtIXLDOWqCHF0D4kCt/mlXANj7GCG4
Xuc6RYa+V0AlkvyIx4tKsTBmUaCSISjhxVRyszCQfPig+5PYdW9imj6LLT5p0nubssLhXwSdYE5r
k0lzL38AiGDZRcIJNokRWEicakoWrjgRHXQhZeXlh5Oe6cgBpHkBm1fE+A2tp9MXiAzS0/UUznUm
fbFyRJUK1lV7Xb5+G8voLJPPIu83kc34d7v7BkneKxQf1zDZZi+yuh5j35q6GJxVIRqMYCC/ItQd
IyrumrKixR7wQvq5jwHGCu8GTi8imqHYAzePdbZ4ewC31GkC6VeAA74+wfuQbC7zcbyYO33KQz/x
ZoxH70bwze/OTeDTw8LsRiqVjNMkZ+dykVo7QqBVq4ks3ag44F/cvYkuYinvDzU6ydnQzSdbO48Q
LTxsbUtFDGL+9xHMljcTPjTo3okOrqVp9IR8Ev4XZvHldeuwp+DV/wJQkvCWEL81NWgiRHtis+Qs
KlgAqvrBdnVO41UEKs6lqvTfhSwS6I/W+cT3/s0x6DedMrtF0YNpVtLbbqU5tOZ86dU0kwafjboQ
D8+MFDl26XEuw9/hU4s3k2h2gT0dGCdiAM+dz+DMRhUH2nSGyIr9/kaW0PcGFJ60YmBfb6l5pihy
q7NFPwuZlJdbIBk1AhYwbCt2PqoQP4kJPbNvTNrTwqISz3zBHJiv0GQ4jd1/lQqeS2hMqR4EPkV/
yPV80dmL3T05LhbjKE0kySwH19XhVt/szd7rR9SoroUJm8/L45SXSCBPM/FT0upyJVgXtS9cojkN
6K2WYbA80AUHsW6FaOOgn/MbXdeQeJMxbsyZVuZ1yQpLZLXR5ISQlWJ11DGoCD/v0NAJhrv7zZOq
uvtzY7pkk5RqDM37TFnTB8cHBq7TJGoVgyMkpbT4ZcWSfZTmFNz7uqN86botEZ94uVkVtt67h+IE
ZhNWR+oVN1lLamrtSWnpibKnK21+l8Sb8l2fU0ttODI1EWpA5pPRM1WO62LGKs2upH+IiBeK1Fjq
5EZjGPsb7fIOWRjuPOVdov1+wcBiABCqizB3pBpc2/RKS5eL5pcnVEDQPg9zOcSlM26kPq4Kp0HY
9m0qyZ7OPtsLPHd9tP6RimqBaV4JKWwKrZ2iEgHmpvX4LrjnLRkZi+U/7wNQ7HieOgkPMKbx577+
iRyJ+/Hcbupqn41MEZvc7N4o9TwgtbYqXW8MLYZge3nib+L34vIg1Byy4CtAiI5g62p59/NT4BNz
Chc+Pjd4Vo/ccUPHseAJBGemO7HBAyYCqhKb/OnPLQh8dxqWlTBg91/3cJXB/DBXbEyotxqy4JsD
iuIa2DiJURSbubL5Upwr2nVn0dYDmE2+QiVQjtxt66ELalIpxkCnE2XAUi9bez7iZCZD+B8/59QK
y9kaUS5XH0fTld05HHrX1aQpuO304MWG5X6KCqWpbJ8T5DF6Bw+ZNVLL+/HbnuLaDk/pdhH59KwQ
Fa0G3bqBIAN4ZT6IC54/kwk/vFlH+5fugGIlzhC96K8LgRb16c/8Nv8nn1ygDkckGlC6Kw1EoXC3
D2qMXynVkK9ghYxTGpDuolPjRFbP9TgqSoxZRjsKadWwEDmOy0ol+R6Urv2JaEDHm/SwY1MzdHfJ
L9NyK/+GiZO4LQIU7ujKiFYs7GB7eFtws3TrbG0RBxVIo9QjqymSbvwULhOJeXQTNijbjbcRAWW8
CNe02BQtTULe/WCphi3Cat0O6zC7vAOz2yjraWoRkfxfXgH11AsEYZB/vD214d9eVj8xQHAROxhy
t2vSLj/fm1PsR8Wjn7/BVg2xHEkLRdXK+BpT7NgnivwfABGDg8HLkQq6rF0856eqdT5MqBoQd9Kr
F7adAwkrRvRug3DGW2vf8WDizRsOLFS8G+JKVrDmzTbcswJbgd4gSBrDvNSmcTSXlCeHw2lXBv4J
Q2tKQrvcdhgsJgKyX+0KyoNk371eaR9xq4JDQamxlKHGZMP7M4+d3fgR2j5jg5ol64XoAQXKQWyk
qJYoqERyljMQgS7cbIv7cuVwIchymsmh5Rb5Wq7Ccs0Em9UknPjhPk35Xea6jb7BMm2AXeW/sdGy
uAz/wiV9VwB/tl4w0RXWdWk8J9JZJTa5V7zfwhUeCSBstoXwINXdFX+NKdHbnCViPLyULaSGHBBo
r5/S1LvcmPL7lrwEH9ysVIUDHIbkLuD2C9fSlJeGhUD4Zgq6trDSNUU7qiUNF4sVG4Kk7bGNI7hf
ifn4Qgvb5FX+0noKK8s/QUZwpXXYGkaz/XOeDvFOqXrgnCQNudsNhKdUpwZJQDKGt4py7CIs4si9
dZ7WBl6moAzY0VXN4+05HZ+o2zX/OXdSDm2otoHUMP0LtOjc1lw2aLrFENtHfyC6TtVCBk/JpNMw
zxCTvQucDkhS3T+HZDVTSv6xOarGnUH5JBzP2TimdAC8xEYYA7qsDh0m05jahIFCb6laHUJ2aNKh
d+c0A4ccqoBOqBqTkcOzBSUUP5r5C7rjS3KgLq1LwhfjuIDcospGh31FnolmxW9BSn4t+KcuNj0y
iszpx0DmfEyt0TVuMGgNEZgm0n+Wb/ty+C/C9iiuvNP8D2/SD2AK9T8/VuKFZjbfOTAzOacUq4Va
pbrYqZoSPzvLnsIjP3QmvPryfmoHT1nGww1XzVOXnqhKZbiOjwyZKnKiYNkk1CJoxliD7Fq5PR61
bR6qH3DxHS4bqcvYgBET8mVspHLRAaMQjgOCWCHe8srwOL7gsqlYrq7OOIn8hqjMQCUepB1Oi+m5
pDx1XT9pzKInEsUE1qaWJv3EAUcb2ESVGaHXb3AIy4i7YvPqOmiQQM7w6Lsi4MGMEovEl1LFRWbG
F07DjEIRlB9g88OpFoi+7IfPBGWb7VyK89Ym43u7yCrb/1UnyUBb0rMpUfwtBu6e/UtzkM7cKONS
L+Sgw5DNAwvo1dY+jr5r8j4H/fsxtJSyonB55wclkgoabei7Ig6Rj0ROBuWxkswmTWXoiXaXPeWv
TdXT6xYrqGFNt5cmD33bDt5f0b7NYMtSiNAHqUSUjJ3/FVZc70qlxoXbD7JzbEDOO1J7ecE9ySRM
dvPkRpRIqkSeWMSOPxX235PjvdUxjjTvSUkrwxybP94iSJCQHjmJcOKgHewkoa75k04AFbRQEPfM
gxTM94qWDScSaxYl5LOjD7Z89dUwV1YUACV/Av7CRTyvYjQhE3kSe0m2rJhJeQT1fCGfYWlJ4A34
3w0k/X/f+XO1TxSINr8dH73I4HvbuP598IVeHux7u7ge3hQeMJJXeD6MC5mUbfotGefiZM4j80YT
kAdujS9x8XLzjvCAy3yJM8osIk8KwDzEB070rh/rJQVJnkAN9DG+w6wtGA3FuYqtZekaLIWawIGz
wxZeBfKCZDVCnG3DfcxXdtM+AgizHQJ1K/aT2n2WmlOZsH1jhS4bEgedzEsux5u2YO+A8h2QfHeW
w2N2PFGu/l9EBBXwdX3Yiu8u21EIRxcswQ40H6uT3dR/mP/Nu8QIHyXRrVUM2P1s0O6ayVKv1BQT
I1ZiSJI4pDIlb7rqZFlOq1WItbPec0WRrSBuea/CJJi1FzSKyW4brjNwLpYFTc+Pg9RBdYGPx1qA
FCM4LBYRWHkMSIf03ghWDlX2/LwqW6rpBMueiHlu/iPanw0fXh2BVoI5OKnLYpGj5UAJDV/ny4R0
MeZjSlnDZglxPfH7F+8ndSVJCWiXChBwuD0Hkf+9NmcczvsjvFXyj8ettFTWh+9BAjAaYisUSfpw
NORg/fN0yhN7UWLulDMTIiNjmR1EGt9Buzo4eh2gbW5Lxi0P/kX1SQgVyT1mojnKa8O6hmBQtNJi
M/VxMGxQ4n8SIFj8DVR9cpF4d1TukLIMtmzC/d3WRgDXVoVAo3Gomlbds4NRHJ7ZqkWY5WNELxnv
H+jDauixOEVnmHmtCrN9S+pQ0hZScmduWmMighe/1tYeGHHJ78dwZMWaWoneCIqqfI/A9KVZw9f6
m0wfuzXXNpFPlulJFaQbAvMjZ6BnMSBWmESiY72Vo0AfrEf4aGSZcriPKELFGpQVG1z7toARWVlg
Gx7U3rcOuU8NxLOj2s5aO54yvJ7DpAgQxsXkdo8g9I5/oqDYH/xYSe0yAIhi0+KqmQxNuciPizJY
u2wUyRrDPD6LlP5n1cwUUmVRMYFsOOU8pssLY8tw4O/Lmp3nhzd3H5HAjwQ6KD4sXWG6D2c1PuP6
EGNDwIGQDU8PZQ+szCbROpEwZyp4O7NYBkKOGnoJ+pRIeij9YrXbtW1amIIYYczmW2HdMyKa/6fL
7sSvYNcYyznIELa920nQSMgvclmc7h5HsmzCmMe/5Jbut+Kwxc5Rx0FwS808gpRjmlaWuBlRYFJ+
GQx/P8wGsczNWHbq166uKx4vsHAvn4ZjAVFKWSq8Rio5LnvcMiqHFZhyd+iLm2ks7sHmAomZvmck
dP3vp+dJmw1XxSo4MOB924LHPKXhwbjW3bnFMWFaAxmSs5yVC8bmv4BAcq9wvJwOytPUy0p4MGmE
8xSiWDWqS7WWfunTiVFe1lIR3ZcAff8YUmF2If8jnfC2/lGXi549hzKLtuDxKonzn2ecu5P5Rra6
dk3CBVbn9PAMxBk03x7dqFhyfvhpydBAcec6Y2FCK9aJPh8488g2XZ4rKm2muWDOxMS88H0W2LzV
pBkh7kBGZi2XCTptN4j74FG+zyR5j+TWxDZe7e6neftdKo/Nl+XDsQUveEpKufBwgq0DtYjNwgrI
DTZZhIJ8haevdGALbmYgwY1EF7GtxffXAOJQNmabWdHlcX6QCYTGsNxl2MZod+W1uJhkEbUYmP9r
vJPFxyYpI+UMAnm1AlY5vY6GiCEcCLbSFp8RWl9glNOxR7PEhY24QVidxhB5iY+7dT1pVju4ZrKH
HI3MSHyJNXgXLsbTwcK99gaQMiTkbh61+uWvC8IDBDwyDBiJCwlIv3tFry/evVazG3VaRl7sUMVF
bC57bO7bp9ixM6FOBbkVnQ17VQ7KbuMf2NH1871JNgNd5l61Yq41yp/Av0O4BlWitX5yR4flxDTB
iuqLfFCt0fLNsiL6/8Bz6LGv1PRwyHCI4zwZ8lpEthn0RnX1ooyuq/2e+0qVPcc2U35MMW9AxJI+
/Q5RC+LCsYOeYQLo9+2D0RtdYqpi3OmyyZf5LkErZM0UXIWM7OSsglBRXTF8J4/j7rPzgdQetxBR
zOX1n7uJM5mni0S5iBS4a3kdsbfbeYjFApUlPCsBvMrWUUTu75hUOm4aslIk05xMBv/6SW4cX/mx
7QOwpqoW60a61z59u42EC4ZN2nGcdKnsy/8UuYHUaEVXu8KBAmuj+/xwDr++E67WXW8QSQHqelOG
UklFDJvWOYCy9bhEK5UNZBbRaULn99CNdXh3hB3fWiDkTrqxPfG7Kg0rhpRV58VUoAP+6t5EbNnp
Wg9l/vkRkGiCQ/mwDLN/IToVyELf7btH+SeoppJK99qNeSVj0LeOBmoC/Qkc+RLaHqF5FjAvBFYX
eyoCj8EZs9TPfT2UKPql9yQChWJ8m7KYr0cT1Ev9eHU0qXEmpRWBMsXAiwsnUrXmZRMEHL2HNwmb
E53Qyj6/K2VFfXl6qCJPiT+1D29Cubza2qX4Uc4iS861pPk3GngZGm94VBxVZrSBc1WapsmzWgnF
iY26oys/SusD0GOKjGpOgaMiBHTNWhe56+Nut3NEbi1QATFnryohZEAN17oKhP3VALzIhZAmFj72
URDrOxYw7peQTrhNQ0+F4JrtUL9JAloM0QS/qZcmgKP0xvR1ejJj5V6gndnID/NjoL5Xa5c9pbR/
7MFBZTCrrtf/bpzpt7D3NaRNR3qMKVXiVbTGJ7eGk3HpArVKWHkLn7B9nYDIDLcB5Y+2+nPAzjYx
au711efPfjj5GZUNFAkRCgkZdXYjfk/tsfFF06fDNdLbPs12+kfOcdUmegChokIfEwvCyeq4WWnH
Ot+ZP54I0dT2lk6okXZRvXDfOVEXB++P7Hbs6UMO2l+RflxZnD8HR2kqJtlM8s9P35vae3+vNpCQ
6lIYrWt4XDEyJpym5kBfIzPtHC+jCFf5P51aoNY3gehOVQy1f4ufzRrO6FVYPK96nLkFsUrQ1KYr
/6qp4d4M7DMuE1N1k4hBYQp6xWlrIBJL2j61cIVuXSuxLreLhxe1x67dnC9MY7Y5pLtwsxccD8Db
FLcSlQwRAJrOrU1wBH1SSec0xRvEeUigAocbt8kWxZx69xl5x1CTrXj0V5Udpf5WR6NKr5rtVAFI
Z1e+p7tJjd8gCNGcAjkUU/3TZNn2bYMAQa0EF3HZpQQ5TiaHe0TAOLkmi0+jF+x+Po1L+XWUMqic
/euDZc4nn6uxHxyV1+hEGwhIi/VE1gHhamodF0vVJDwWwAxVSYXWFY9MWOn1xiNo8ESV9MmPypZS
PLYwG8/+gU2hKus8OLbf4ULXASvmluJpmmyfZ4/DVAhoHrhNdbrqF98JARxV3m3v4F1Z+WtX0xuV
7WSVNXXc3EinZmsytgHzV7y/dlpcQhh5az5EskG5/Dy5kGOTp5QC4TaPnodfh0Dhi27TMBOJSytq
5gQ2724qQvMWS0AsBXxfgHV7fuv+pB2hFVeYpEGcmqtVXJeCmVnwUg09sIrjzOQL+E80suY0u9Vk
BgGpWwddDHijgm1qNAJUMPSPeeZZxWyreJ22G70AT+T2v5uU+22ZLz+1qAShmUtlBFQWlTof1Fkw
EBiCC4C6dwUkxTiL7ImB4Oo7rwQna/caPJHHj1Zn95+o54NI3TN8Et8uRG/s+zT0g6yviYu/U1hz
WpXH8X6s5wP8ZIT+I2+5x7hNwSG5oJzX3rT/g+xkmKkUaXcHFZlPKyUOk1gMZVczU1p+Bkk16BTW
jeRnXarHn94JWr2ZbiNetSTRnkYhllKyVbfDLEp0z1b/6w/GdhI+D3zURzDSv3+cyIX3ZDp2QsHp
yk/3eo32iax5BQq5CJs0QC5f7zvDGPysC1dCN+IM8Urw4X/7U5/ohZV3mKEGDhGQ9PuDKVPgdjPT
95FsUT5odhSby5mJDfzMBy7Iab3Nje0tpo7YKkzazv7zlhCQufPvgZcobNOZ8caEYTbp2JID0mS+
v2H4aQWItXEat2N5JBHXkuqZCTQGWDqWdCsLesfGRVCXcsMmA/PB3RS/LhLJMjVmMFnTYKL24aX1
oyCOiDJVdyOcSEasoPUJI3/SIrufhVKV57BjeEdssZOV4kAIdSBl8QT+hiUjxgUl4evg6Z2N2qwm
oH8FYBvCEfGVZfCqC96jW4o8ZtkmGKyV7ICzxF3bSQCyghT6SezJQx9wMMxKPVM34BRO0lpV/LTd
Ov++zcoRcXm2NS8h9I7DbmEiYQUVrjTwqoosOC69PkI9HPPuoKqlY5lPLDYM2DdtqyTco1CCveRD
ruq9qTOh9vSfB62EZ5L9vSMMGD14VFG493NcwPrE7VxejpZcpa+gbF9iVeIGJ/K/ac+4QfbOoiQn
46DDtDpuqPnrRSSyElfSEukRBIm7/1qJMpz2q6kXPTqSkaHycA1eo7hJmNjZgcdwZqOVOKEbjd1i
4k0CR00+l2zUYmH/izqasLxi+MpyBLZbMSloeTuHMCXEf8mUVqTG4wXU+BUTiY3STYP1/xjoy2A8
mRebg618RX6z4e+eZTaENAFv/zVTjPq1qnferfWYv0gn6+XHFKWewHX4QrzM16t3H+1tYYhQEm0Z
7V2w93YurXMbtFLP57zcaG6xb/g0zquYhWWYH35fgTe6EU8DRLJD2DIkL7pb6hgs6ihVObJTdIwH
khEQ5goy1jqHXDxo4fSpKjl1sosjX7seczJnQMIC5MOXU+5NgLVRJ5ftZBm/DuD7Gc7GVAIuUtnE
mp7ktTqBa2lehzLsPZQ5oaiw9ug/1ovrlbcGK6M0PdTJ3HUwL145XbU2W0ROBQXc2//DI6XCA09U
jotEK3obgAkhYY0UMHANBz5ehB1JB7NG3sUoPIqXnTbBqBDCXGi7YAFKHmbJF7HA6+zI/GjKZ60S
Yfcb9Uz/X3alniUkCJDtWKNMdVOXR+uWhJqemPFj4NwWG3ecuShkrtqpI7EfmzsPKNADUqNPGmha
OpOVtOG9ZZ3iu2QeyVO0oNnYjP07IGd3fFB1z1erW8LwOyO5zL1vEPOYqc6egEmNrvwjw7BnP86V
25U9cgXsPJTfo4XIB35MdZR+V+gQJjmHTq+J9GiE5KoiR1gDNeiDHrZVnTlKfosQ3XzG1ttDmsOH
v9CDHjqJ52Ah0O5IIrJQr/DENpwb2gviydKGLPmGCFYYCHJUYNJTi1Uk8NHs3zhUsZPbzJ3sczBU
+DlBxkznCwD5fNaKGHYEbAvo2ArZ5t/VQb+c0L2fc+c1DfhTokV08wqR35LA/+uqb+kudCOQ618F
dU3+ljtSfoBkQFeKqAbBIKHKIOT2YmTIMujXhkHcsmkXmkGziKX4MiQKg1eqjkISIfKBDTQyLWiX
dvOae3yGXU4ta9mx3BvP8gP5+VyhDaYX32cRd7IuTlDU/CPDojJVL277QiKoWarPpKsRfW68T5kG
qbxTOuSsk5KdKAkgOnaJ72RmAh+KYXwI+pS/YDvl9gvQbxxerZG0msJ4ixB9y0CBokb4kJ/2scwd
+ZhKQfiJ+FqlpsyCBWb2jOpEbowRbYEO7CDiO2sd1RwG0LBG7+7/6j/AKz0J33KCoyMOL3qHE23f
btGQWxoDQ9XhcPwQcSFgXrk0PthXF4oeTjlv+durC5cAKFTdToN/6eUzcj1bzcO/PWiMaKKo0zli
wUO2LyA2rchqjBRxkhniCLM3BPd+jz1sCr12bgPE5JNLE3QVzq4bNO+VJ8XfrU5DN2XN0wJABt48
/LT2LzSpolkzsrzInX8/ZNveGc2sIMwSQZ9UlWfr6FL8TFGktxo5vEodQG49GUi87KTwOULJIIlN
fi/Pa999PBkTaHLfZ2oQhUUVh0Wp0i26sF50DYsRJ5OLY4amfW7Y7Zw9865L5Ks6G51Wboh0c8fi
dwhyU9ZGHZJGurWlQyz7Zs1Q4c8b79qzx88SQpXnO7hFR9c2efFQPnWnE9g6wxSXDCko0k6OCnrI
RsXR2QGblLym7sakMc9Aoh51ey7IFoddNtckJ1ohdAy/x/aEnjGD+i+57Wbx7VDD8u+GC2WiKQSh
L2A6pia43doatyGngttXpXAoLHtPktrbdxwkDWbJCsNvPP+VUhGginzdvPI9YzXaxvphOjtOB6dP
zbe+kuYfPncJtRZ1fcJfMyYy0OrglzHE0qxs/jvzN3s7Dh56coXsZcFdG2ytuV8UJYjq6xEA8DT2
VYyR9XTAXBl19qmYnG7SeajF/QFqlQPsQLrfSEhkV99MwTJWaMpH1WfFTLdMbZqVM8P7A9gYLquH
iMwrS0RntPnXch7SKrnH0l+STlS+K3CRRIdqIpb3eKpDngUN29rkXGVmt03kOtGiKBe6VEAXbTl+
U/OEwSuqYgrK06ypJBiyDkX7GMmLA0e3MqhdsPEOzU+YqZsqNcd3GVkGuIDoAYhxFWLSfH39K2wv
LGPXKUvythRQea994RX1gF88yFpTMp+HmshH5ImQk3wGJjz2t5HRjJ6Ql68ANDhisEJOMPTaeaKy
M9lhnxDqWwR57Ohs5vFevSg8Tfc/D9gkIln0E6qOGJjdSFTiJ7JeFahyDLgVngvJRg55efND4EnA
wJ6JOzrEbsIg71Bw2co6xdirFtdxPasn6GxrN25gsOCCLteRqOtnCMA1O6CT/K1tCv07ko815/ZF
lIGMa1PkyVC0here8QFaamNsEhjt8XDOaqS9nKoefrsdSaAxSpY8uRmUfofh+54xtv0xIVBOZmei
kVI7Ju1azHZLO9i2il4f6eHwU44Kq8N4fiArwrr3Uq9VYnkcL1C+Uv2rL5/BlpHBTdI0XCzcZb1e
RBODKWLDSrKUzMnxaTIAEewDHgCetLXR6Vuc/pCoO+OtqeL7eeS9wfGL+fOWjUxz4Bo/nZSsLaYY
AXQVWdeR63L3YxRz975iHmOozOnOlTAg7C0zkeyQH4a4FVDJDESP8s8ieDlO6VGSM0rwSly87pLp
durtHFHzJHC/uWq6u0w1j3Tzf1pbudhS9PNJoLc/5oQZNyEFO27LtCMV9gq2HdxP06EM6tibYIbP
ycB2MJrg0DmOaKbqhFyyfA4LOe7lAk5Fwx6cBYXaUxf9bQkPJCVouHccke056dngvlkQR+35o3X9
zdkMu8UApIGWCMJ4NSQhMjuVx08BtBUP2CxvsdVusXWzILwd38UykYGtg0U/bLlvuKXfTbzwmFqs
zczhK/giIiqGDnK+oQohFLjaiFb/stFYlL0hdadjFkhmH61zBqre9qStBIrAzfgY+t4gKr8xh7JN
umGzTmvliZy7FKQIRxATinDm2+ILfpLySd3u58SnObJvEkwebiIN/euBTSQtz+NPyNg5EJJM3xPm
AvIuci2CL9wnKkVFbmV403M+7QayDdOoHErGcUYTmQgJi0vdhC+yhHw8j8BKzloMmKpTj95XKS4r
hxjNy4sVx6/OdcvjF2SFb4Mgo3LaR7bCgxYzrBPjxUpz2B2+L7Rv6WTnPIvWzbRDWSeBuAkn2Dhz
0+TNA4C3lFUrKPYTArA4Y8SWGVKZTZupNYmD+it4FfYcwksrbk/P4R+OHz3P0XOLP8m1gKLD9uzi
/Agw6Hrw05iyTL0N59RWPsNcM2iD5firdWfGAJDhCV0eIpBJz+N1uBpcRdg5iL9P3rVBeng+BWLi
TsaCDbgyuDVoOsQMCBwrlooXvoEVkJaoVv1gp7p8ORtYtivJ9vl0WOm7bd+X4jRkIcpPSg1Zt91O
Jk7YbfXMpLTeMWEb9Vm8Hf6KGIY5OmWwb3GRooGRFfT0fM/SpM9xVOn2/sCnXNadN/SKWsmRoSi6
BRhjREbl3+UufCDheCb7QJsj3+cHGKXgdA0iUQRg1ZtgYMS5YV6guaPKosJz/PbApTKMjLewFcdP
94DOC02Dw7B6hVv7tyxMpl6Cm94Dy4wJNqV8PPNZaqRCwHLfKmoPXZdjT4rer3tXbNniNvvn2vKj
5o7w7194HBNfIMBcbqLs84lCEhlezhD6GdLgQv8VbFQdPmoY9itD33Cns2O9GGJP+77FRUbDsIrq
ZLDUNYCY/TIvSmLZyEyliTNOwPozoQK5GzOF1fgw76CWLDeRJ5U21ii6mHTh6X98iA4eZ6lEhs8u
lCO+0MgaCk94Ew2TqNomKrUT0/sbR0JnLljf0BuYT4N9K8JMIeq2wzqNKK0e4b8FSMXDtIUzRXc8
CyVU16Uq97Z25MohGW0ZfM9JXRfvqyWgdqmFw3F2ur2wTPdZ7tTHN0yJiSc+cdWuojrnXxvmzedj
2LA/gkheKQefFbWKYC4EHCE3X1kBo/9ORVC6TnSCeBqNDAfbd7GOtp5/tTgqw4uVUnlUC21bR6NP
H3FENzNAh26xzBdLT+EJF/bSvcKtJnqylOIcbRI3o+7h7SnFaB3pBV61Y0hrJAbOegmFdRu5RHh9
LsgYP+N1EJIRnBz2lEIDtiGIKs/aArAwRf+cOGm7XZMl1DmVJy+LVUdW9vVLnxmxuBu55VNLxMHv
4k1puw2TQyIMeH4KPDrrDEgc8/ceNSadNR0LL6cHq+F3uXQ4u7wi8C0y8Sf+TadV8TCCD+k5g2JS
gSIEplCB9WuddGSXpKiaFPObp7lXq7N0slOPZQwW214JhEEFul9epXw+fazyB4rQDTXu2/nnfRjz
FfU7kJyyNcNz+o4EgivBs9M581uwbTz64Tlu2aZI3Ms5RQmwP276UvzkNe27L2gjtYmsy61Ug2FF
F/KbMHR7kAW0JE32ETsmK88iRNV3NgXCD6nFU/oUBPWaq2TA9ML/OxkOAMEXhEkp11GFRnnVgHg+
Btov7XTmqlhEqfrX6kjU31iFdCjolxqvxt0E8HrZwfCXbZNvX97Pa4mctdlvLjUoSc42EuM6GMSm
qcUhdYdZLgZyT0Cgzz5na4bgRuK1VDHCzM0LbFd0anbVrYxSA8GBnrL44v8nujKG0bfifMyPKoih
mI+6sVnQzQQswqLpCpdTpWJYA6hK05We3viJ2L9+BU2roH0q7gFr5t2XDaoxfRxwx10GXTFyDIbe
OxbjUhOzpxuWLUTxpkRqr6fQGCXqkho4mpKygFS0CM2qqITI+SbOzmrl7h6Bot990v8WSP1cG8wV
eN/fu80GO+hry18a8N6Ceow0vnteWsBKieqhqJOBrOSsZ77ZPrGtmuilnIaPkme3FDagbPjgOA9q
xkLCmSTGuAkmtbcCad4pCFnXNzpFOvNgfrumPicZKWw4G5TpGw5pkIbOTYubX3F/MnFY/XwvV8cn
KV5i4G+6eMIEmsOBUfbraTvJx1O6vdG0+GwviStfnx8uWZx0WYOysEAJC22Obp+rrR2zlR2LXIUq
E0krnWWEkjTaN+YOve8Zo2R4B3jP3Kg9U9ld5qx0EmKssO7orOILSHjC3aOkoAgDr6Dyi4I36G3d
lw/uF4127/5OA1Eh6NqIR+X8MjR3zCgJM9vpTHdUcTfp/3PJ9f4/+WKoyCBuLwn2YoFALGS5EdzM
piSjIabCjFnF4zy1N7WSRaA53xp8BmsIfZ7gZxdIuDPzx6/oHTbr9tEbqMZUIfMOT+06HZa/oVF2
MlJ/fk7IoGljNY306SZ1csvfWsUl0xlloTqGMN3H8SwrXc8nP/X+K+eJy2/qyHERL452tmkcp11H
uvqJLWcYayS3yyLDqS+x3ZqxoqT/MMp2UZ/OA1hGL5BT0Lh28iMl4UbNNl9k9H40rYH5B60gjFDC
tb2lBBtNJC+QnacmpLr7kQtzSKyMcLgYktU/sI0cOq0KVfG0ZCoijiDFsAwVbQ88TwYfVBUZRL1h
j9SXjGj0mSsgFaQM/ukQwIHSJPb6DILqgogABEdlH8xpuAHUENCmE94wQbE/3fOYYMFfqV+nPfnC
MmWGSPpYXrOnlThJYiXKGzEMmx2q0s8JwoGTA76UY4G7+bhnvk0U3lY6niHs/U5CkTOyVbGC1IDu
xsMPB7r37DRyL1RgYn0fsbvnW9QnliJdWqx0vpLuuAgE7LINUNhqKz1e9kmQs/4mNBslxH6rl4Dw
OqbcHMzOgQ8WSDxkXJqvPww1yPOkEcLlfswFDsqIlKBYKWLO8Rrop4VLw17LZWc2YSL9HGYxo0E9
A8LSYFMZDM3EVH5kcPAssRQajGpeIZiKxmBFKELaNqSA/JhB8CgNL2yXT6MYEH8CGXih7rWzsBw3
0xVReDNTMd4DEhy4qWl4Y8BUWsqhSzCRufuW6GfVH4LuNtdWgJU7uNcJZAIixV3mWLS2xiLsRm+5
Er7i7u/+yxIs3qvwFveOC71XBXslKTRIQUQm/oZA1Yfv3dEuDjOmypPN8ymJWlORaRFN+qFuedIj
weNWx+zaf5jlq+LxpmcVw16Y0gEW/ru+vlNJRr5G0vOmFcL0bfiCzJKvOEtv6CJ3bZqVaPoi4sVo
AUyYKLG8My/k1+5K5wUV4VV60zHsSunimvd0OkY1juw1NXjceXAYU1dAp4cQIVdrwX3Ya8eEJUvB
fDJq19TFRbe4MIRpjAxjrEiyF+Q0QjWSQbfxV60jtHrODfQYUYKwpQW3gkad+pTwMFy+AEYsGWW3
Y71SlozLmHM9pHzVjU2FOBoceRicUw8bxwLcwTpSK5BRJwbFNQos29UfctPvAxS1lxO/SKRAyj3Z
KMWYZTlbdktD1r3y8xCDZ69KFm86xIEe2+eYKQh1XNp+Zwk6Ph/r4BydIZfgnVLqjmrvU6c2gorw
IrcubJTLWx1h4HqjuJK2Zq4dFbbR1U+o9STcLiC+Wr7uOHBiYOE1+3yjccK7/7J8V7P1pTMC0kzU
9jk0e6Bem//WATxu/GXE/y1ZcAkQrwSiScISTHP+OE5pOsAu2bG96u3Gcy6N0RhsJHFY0uMw7Ogt
Pd6SgUsZCjAQmBQMPLg+bXX5emRdM7AvAChAh6MWHCEzY/okdrLZZyJQsE7NoSoNTb/z3mYsJ7Em
CvQnHzphrBj+LSDI18/Um+bXkTqoA0o4+sjkRdrb36Rnzrju10ve1hNNU3tejK5iAWEpWr1eh4i8
Exzj1O7hULwH9oTAQhA9I70u522x3s6+VAoc9v+fwRhpTw+lGuS5QbA9S/EMpl6YXH8C5nx7rpyT
wQZbQmRATIs9Ngzk/8noL2TXKjk9imvUAus222qBFjbaKY8fNeocJMVvoSFH4OSRJckJrIjnYGKN
JYo9C6hfd59KDb4nZwwXJHRe97EW8Un73a5lawgILjup4pMRXO/7zCtpIKf+tNHuWlyLYWGIjL3/
ngQ2syXAQ1Gjb9NItdXrDQ6VAqvzvVahtMIexb9jy95qlq3aaedSXJCInrkc+i357IfgYI+/lDc2
RQvwZJDaYUxk1gz1Hxc/7YhyK1t2scuIOeiNA2+hHnMlavH3xYpx6UJ0vVhbVrF4uoqlYbjjfbGd
FWfUIs3ELfvRsv6ynBjDlZNNCUKu23+eVn5X+QLe3IgD4l9VgptC06HxSgQnOTqLCaoGmDHJhBES
5IBa8ZLAPz+FKYGa3IUbHkb8cYuCOuMRMbKk/6YoRteCIVY3aOYWXNPC9Xx11qmeqgdRMFcGfeOk
BH9duzsSFj2IkWKwOz3qjFcaXgb/OAom9T5aVO365HU+1NmDMnoeQrg1gd9REWmvv4WV6wVZ8PBk
Ohxley8K8IwbJs/GKPAyx2XAZFu+xVFVn82Bes5NxPa8XP6ViRD3thcJHsHvmUsaTumpPePKxlys
ANVcfhUXELQ6ZLWr1aba9k2GLOCRMNV1BHZ19I6vMYeA9pjWeI6RrCBnr901LjCDUddBk2k1X8OD
n3w8407KFe807D0FWpkvcrQS+PJ1uyN0DxaoL6zfqafG3NnCNVYNFL5WOVqTsw93C79eE2oW1v/S
Xxv/pSWc/bypjx9cf8ILipwOVTSTSmyxyV+mj+svssypg0dHzgCGwFFeDVRyHyDy96kVhtML+tmg
+aZY6kD4s/3MDlNgtECQ5ltISEWSBhxNz54IigxO2lQIEcI/Nwf5EFyBfCP0/fh2Hs0HfJtFvVRl
kACj3hQn0sBkBERLCZLhWrmzA6lxeXDjfdf0jqBETi5DWrlybQz1mbRoE9JUwIixTGXFDgwtslEf
Kiuu6iXDiWagWBMIqjaytm9+2VpQElMi3rD6Lo5deDQyF9Il5p7ISRbI7P6kIY0FuqQ4lS8ttoVO
VbSiaBgK2TfI5umcWsGhc+7uhE1AJGDNWe8PMHDDjq2ch46XNo5M0d9kmKkca1t/YXyUW2KVI88b
C0h6Ll1IicTy3bQAMmdYhGVE3Din2n1QmswBtPeX82SRUXab2+vdPJg4GJsmpZ/pD5S+MCDttIPK
bhefRLh0CiiMhmjnKcXrKQe891aIzXa80N1Qyhsn9nu9UOvv8dEZe6pxsqOou6ZbPmb0bWigjoYL
0957nPeRQxmlGmPDxSiskFeRZL5WnO0VWVIbz/OKGwjKzz2hHOHVrFed4OeRJR3u7ULQHKqA+A3/
PPJH0RjkJF83X0fL1hBijQgcMmxvMgTxx/keSj+DaFKC1qE6Gs3XzCel6+42KDbpKYoKIAQFdcVU
9oiwO82lfz4ceV36xk6Ulil03vYVIUGR48JE60s2rXX91/ERTafs39O3Ni2abQmizyRVLOsAbp+1
johMNzGOHFXbYeVwnd8y6JDj2fx08P0oJYg2IRfCelj2n+Wc75md9siCEdHW/6kvm63ET9jpDXqR
PVdrBk5t6fXbowRqWhDYAJnkw0KgyQeikzdAB988FxmJgLgtoVum6HYLIxPHeWQ6DYtHz3ehaLqL
T2vz0GnRhO1Ssd2PV6+NUM6bgIh58m1jwM1OEWWSq8J7uDq41JLHoJozLbenaolw33cwNc1yIH4v
+9XqrQCWNLxqJnUJKSAvIyikAAe2o7DF9klrg6C9av1EwGRgCkIMrznUAiijtvA6P4qRPMYtjWm4
ZYnWTpBGMGMCuGKq0etBfwcc2AXGPp0N1Wi7lBFF7UHBUoGC/9uYkyH5Z+OPhzNGELpEexJ7Iomd
KDJ/ZfZrIcFKyM2HgxmQgiVXvdPUtEsWLCNIm3zKj2MXVyELxWZDlh/tp3uXOWzWFT+OrgRUKPM0
uSfUCbtmXBuRn0+H6oepFrul30RFS85vL929gEz4G6zBOwhCbDWpBXfITwt9KoJmH9Zp//iP77w3
IzpNSxhvPBRGpArDOZLA7K31qfnnSvypjUY8d+W+Gmun5TMiKps7QFo+udPtV5S+2CNBLb4Bk7mf
tXPcfX/7UUhGtVq6PWSXKVyAE9cSQy2cN8vOxVcGjmJqoQnqhF4YzPepfK+7d3dYjHmYl97ozgyU
wZnpXC2Gh7tD4FToJRCBUhT4A1UMV9d015lOJfOLKRn6w5Ku8Fw8/BBAtYb7fivhg6GM7YxDDMGd
Qa01R6P60of9eadyJYPXij2ZqZjeIlpBabcuQQeVgIrAJZJC72T6C3VAG91Sy7wvmPq9GGQqzLeI
6++j9L3URyEbJJ5Kv9ZTi/U11nhqgA2VaNSZ/9YchXawswHbeADHLymZhxUrGixogyh2s0xKqZl2
69BVYjUqrKyyJiM6bs+pMmHNQjsTa/S56mkPN7VjtHYEhMN+mvv3dEJcHTcN3Hqsl95juANkNNyz
jx6rfnxyCx2gjIXhPcpRpelEq62go/gpl0KgTIz1vklBYqyWrPzP1DqUcGKXjN1ASIp4t/ysttpM
JejZK633VgdLHWEe1XSP1I8pK1EPoSk++dSjzO7s9hBahsbpltUuiTSD8DwDHX7JcP8cq3BbNyQR
JxFYQBB0kpKF2MjoR1iv0z2O28oznZ+MkzaT1r5oLZrAaNwn5zgsu4cJ9lrW8xQqaU0OhWrqZ0o0
or65u1Loii5mB5Be2ar6RQstlT+3b7w0FBnei1ibMcfvoLmnZPbgp3U0pCVkVn+y/lsplm0CFdZT
QeXVn12bShqaw0kWNlyKqGyo+4bpWyp30sheJwDy/7ZYQK+RDVvu7aE8Jkvie3/N6VMRUvbNhkLZ
9TNbTE6RU76WnRLSG/CsjcZbNONwqP0odKXWj0VttwIQh9IuAln/RTrU+dZWBZTe+yeteVUPaCm5
P37oiHd9ktwcmIqvhHs6eSl4Y7agY8ziAvk+gQcN2li91yfbHEnL1+jNnRMv5ncPTiyIY1yxmnZM
Hv/a7FOYi0SSFKDTOa3w8b7m1y2dkaS5CIqSZQiSuINHM22v9+TV5q3yDh257tfrv2zbJhzadSMc
4W4T1dkCODkzRIo7+/jBSVopAaqI1oD3wB3azNqQiRdjGB4eMuryQGgr4tRqqcQkeOZtAo005t5F
yI1bmHq3JJDpaBiBT7C/fOim5fwBSwRu2YdTfggE7TIOCeHY3hVA8u3L5D2egclIKzJabTEbtLCZ
cn2ujg41uQxnhbgjlYww9UoBpdv+Ztga5hqlzQGaJpYAMI4YY0W1+ToeUmD29Cs4k6T5RSEURLQT
jbAg0r3eGbgznrn0KKbzAYMldyDF++FUP3uyP0RWOP9NuVvbRHErYI5Vkf9VhGYSLbkhJafLSK6g
HfDhKNVAaGtbxR1iWB8WDmNh4z93N0ifAxBtSmmBOQEtUimLvnpkHLzY08xxZ4r0G+CXW3AlhwAb
b9QeZH7N3sUzqeMt3ZEsAehUdSOA7FICoQ2bicj8/hbStIrHKxsM4SrdOEiKh1g/dIzZBlGEl5/B
NTDEJBhIh8Jk+y1V1ECtKt5ST2Y/IYOKRVKgTuBeuUjpFRcofirsFjm+V5hvXgAu6IrndTAy8Q0i
P8mseKJ0kacxZRCa763vvKhFVJVrP55rYa438pPgSM/4PSeHdPX5wl3ODE9SodD18zjK0ZhaATxp
s1ZVdizxWF2zdSi23eNKQAXZYMtdC7EbqxgiM6VKuRUZX9BTW9Ht0DM/aPxws6W5AxA50u4i2erz
3rwSEyXPWV2AS9nt3J1mfK0KwdwVy9/81qE2st0lun8ofRY8fQX86A9q6Y+EdODV6HmgF3hdhh3k
fuatEzx9rE9nO14pCBnWKVuHvWeaEghktGvu8qbPOTXsRxoIU2IenvldxvNz4t2WulE/++0hobxm
La+P1MzzKg4EDqMb0iLktBQKot+8yzGmOuil/XIJawbPfkJ03ClGP3FnDNLilVlzE/Pgsgn+Ujbo
VSn4U2t0wwfw1cV8/Cj5OVDuLSSZ/qvjMKt1R1Azl/gijc8GLxWr3sklbXX2r6I+P05NjIRyJaCv
xVo1yguA3n47tYhtlPhIHRsk5+OnfrSHoDcw05cP3CTtNkTAu7Ddvm/uCJCtEqCBz5MOn2CIDBPe
BjbLnOYmCMqN7VwcrAKmJBuMivngipYXPZWjCBVbFxuNEHIcJ2h58sSY4QD/J84Xggi2Ytv7Bvqh
KPQZFVmB5bPJSFWOIfV7wdjWKSj7yt9GDSoXpiFLeLUAaOf1zmL4jlzJPNSIXVatLivZViBLj/b1
eW4oJnGxw0d6EGkgAaIdnXF3umshGxueTBe2hApMqs5f9HyDxP6lT8LOu6JxEDO1TFTUjY843H39
gTPxGyziQ7PR4gVukaFxdbx4AiXoDZRj2kwh4goYPqPXn7ASHiRvX+wadGNItsR8io4KTwh6b1+B
nR8Qyfj4gyboaabpMBVEgcAEUQRWYomheRhp/EptoKQv6WzBl+wfqjm78VbWIfAgLjwDDUJHLay/
fdt3nuiLF4C6fHk7nQ4jz39V5VMo0uaIZASB+EPRM4yGQ/SbKa0XMKt826JM/JNmsQeAlRpeMMKo
gGtz5CQ0mttHdY5VEdGN5Gaik/ThfvnfvTLpupl129i2S1Fg2RVGjKyLP7m7WEvCku480LdZ0pyW
vMPGXIcG074jh1CUOCmtJpjtv7COrjHs7gAtYpFy/YvTK2MEv5I6uNAtjtqCawXRS52cR04qFwsY
0O2gdSr9zpA5T9DOTfNg+PYgjO14xBMw6hslVskgoEZURRFSx3tDc7twRYjCPeLaUBqHgmVJgyya
JEZ27HibCE7NGUNvSAdAptcuZdrCspY0lt+xcbTKSAnCbGrT7hicbDd2jL9glMLW5mzs3n5yNwzG
KOr9J/VTCn3DPv6B90fZGlpPu6h9k8PkIT3I+el2v99imySjKMlw/SZ7H9hmq1DtP9TOTq5je+4x
8ChyQslm7iABsLY72JDF9ry+eyL24jjb0Pr0280cvIkSpmwv4+NiTa154Xh54jDsPJv30J3xT1lp
mDd2kT1WWrNcd262YjP2o+84vRz/BGJoRB5M9h4+jLz8E5S0l2nCoEIQrt6L0wSM6rzyflGXbijq
fnqvw4aALtFcRduXbcY4je60xJJfZsKtTanfhNq9SFBYi2xUYZVTsi7SHgSxbFUkUnarzEMsOodt
duG4AbrtXUvZIurYcAyAFLVNnj9g/jZIDATKC8rbl37K8M3hdUk6BlV1Bm60XJKnaMWedsdrj4bp
FJHtVeYU6siuqQYYhCgzu7afbRDdg+MzsY9beog6lbECdji57Gy9o9cW4OCDjhsK5gD+/Xk3uFam
lhdl17Tj2SbhAxJMX3TOFzb1wPvBr1cRl9SAxsNsIvZaI2CAHy+c/b/JgTHsM2SECnbKasZkNX/R
BetcAJSM+VKyTIVR0mkDsXosTiarCqpQ9xZmlZB9s5tIiThd4rLegrigeXe1lbM48FeZ2JYxtokQ
talfRT9272g3yVr+aMe/3QEz2JNXKg2/rOagOjFC7wlJb7aci7hogEaLeY7eqXxgdpvxbquKAq6+
Ns26im7Z+7AEwqX4ynAraeghVzd+hqMIdy3QIrMA6iVEcVST42cpTfYQe4zvLKPVloRc2NgYUbI4
Z9faaDq9WbTWvN4/YB0op3cljZ9ljb6g4tWbKxW17zT8b1nYe7cIU3DRsE7nV86/mMKhirPKq2ba
Wope7DEH9Vjeb8RhVQkzjasP47uGfh2wHMRfCxKB7bVl34volL+7KZE5oid5GBL3yi8PWpIwD1wv
JBTqIaccdgbKNC7pRPAWUwbeTI5RtwH2UCp6DkHmWi+f075w6h8QJAcBkGjkdtv57cc7cNYiYcd8
rRhuGxzRwwMTGzKWyT8CXKqfgxL3k7BDrrqWgOEXbwk5q98DUzeRP0ReCs2oB90tWaFfuOhdXI+v
Be35dNWp/Z/+CcelGe/AeYCio3wxvN5g9PtCD4cvXnq/VX6bIzsa+S50CEFMUnyqgzRT92sGUtpm
36XloTO6ED7NxbUkDC6v59JSjjW5M2FBv9gIi+wvAylJOxBkGkzc4y6+f4MvVI1qOkrnb4Ve7Z74
0XcQdSRzlK1R799DwmXWNAd4GmlqPFQfR77s+pt7huR889MPXCf2Me9D5QbbddoSXLy9fvAGMeTi
8qlr1OfBJuewFkuQBUwzUa/uDC7AHct2IDcLjLRen3kq0n7G2KFCu6m2lAaFh5RE62TNE/+fAnrx
ZPo90vIuny6g15gBjFRvcL2sxLG7tTLSCmmbkwcCKnW5MUWrMO4e1e3v4WFme/ZxU8yp7FazxUgO
5HwG7rfaLMyF/rv4Zic2vgbg1yUbVD38lqpEWjZAoEnrbvLs39IIY1yGHHSOi0mMPBz28pG7uzqe
W/pGRjVlvOmBQ78sE4fkXdWRkVFGpQXsiPdI/n8nd0mwVyYpycJNihgV+uLHkGZX7ZcvsVEp61LB
SiVQzkoiO3WbL5SixmG71Z0PQF+9qXQGzeUNf240e8hzaf1KVpJt/3D/co9/todEgFMzykHYrUQZ
cm0NhZvnlo7iJZMhshhcdTS9UK+l3486eDMb49Xc2/2KREGLfqdmn1SHwUNx8LeABN37UTJfdBFq
X+n6t/oGep5slem5vxqKLTyFmxuFCHw3lMEHlZGQmH8dCPe6XiJ8+jQfCHd1aoLVH3WNbfL/W7po
P9U+5ml8Jn8eCmZ7KMleKQXlxJj2RxMd6OFJp9ZDEedj7vW1dm9r6jsJ4vSrPL8dwdg2F1Wsi9H6
qHiOnBUIJoyy4zadnGegOFJ7RDSprwNdDQr7jvUMUGbq4qDQTCcTN0ohNG4+SRbOYvdRsl7OOYNu
3ZzKTSi9dN8bffFbDaXjHjAos9k5lCoOa992fw5ZiAudsxiAu56Hl2Stve8O5SHGHQQ31sE0ds+7
zNYFIFaJ2gXptBfNgtJxab86DDYiP5a+u+CBcWr7N4ue/PaiJ7UPucfhr+l7Kdzr0yE/MglPklmY
DbuHrLDHwFu2e8eT3cWSOHsrTUUAFGPgf/WhL5yoC2LL1u2kqsMTzZ7XcW51hWauXnxPZqQE7aSO
tGoW3ySlNiiUGc6oWjtdsVgGxJrSpruYzKUUDVVjxHe/Y3+OUOgl6EdHQSguc/iTqCU8QwHD3rG+
m5qrFmtUkQKT6pMcBNQcOrPpDpz0KZPVMviXaL7EHUDLMWqAM+/XxrYUMH+P71cDExrm5GTBjmyE
pCfWYY/0TvLdzcaV/t+y9XEbM/aSpY5rKwA+DV7KjNGlPoSsFc8cEwLdnsp6oAl/5Ubc6gCuCtX6
aW+VEfUp8bbV/DIf9irSCWSLUvy0U3hVSkO0I24DrHipOn2lcFkz4WWP2btr/sOlXKMLsvEeqJ7c
9biz/AvKbmVn6Q6X1VMzUt5YWVa7kpOKQy8kd1oyh8aa182le6ylp6cda0U4W9MjPF/xie+qELut
p1uJMG5fXedGbwgAhcWx5ABdebDT5a7Jkxy+OX48Ke0q70v9yw+aMvaa2aQh1V+RcBNffc5pqyKw
Zk1J8nDzi2ykT5ILS5+jXnya7v/E3A/0sgqIan9taF6jMykQNuYptyGC0sYKN6OI3ON1CD3CprIV
UQJV8UbJz4+efdtSOiMWHYWonBrzJFgNEQB7sWh+ZP7rJU0IIFsup5RxVe5fDEI95b8K/M4kKlA7
EK2G5fFabHFVKL+wfU2XuHJwD31+qDlLxFyUEhidiw92jQakxUpV4OpT/mbe8+zcUH9VX+1eiwbu
tZbcG9Ck7DLB0N5067LhRHvZRnr+0DUWWNkJdacK47DaaPAlvG3Un0j2VKYp/QCw7SQgY24YpBex
ymODYtQiEWPq/XrE5kCi8biQo2E0KkTCCyUCJavMHukYfFY5LONilulANT3HYZK71kfLNGY/4wUO
nxg5lCbZF9gv2tv7mXenag2lU2WTi5NyRnYY6IrJkAGDih7sRuv5RafJ1oobGgnIjMXHOIpNm4lp
K8CudQcRB9A9DecGDVyhZ6gsnozgvKL7kpEFka1Drhgd5aW6YUxZ03HxONUGOSWl11wxpRYco4vp
EHR/zrnKSYgjY7KITAsEm4ePOkOKRGL2EHX+gaCEIRoQRyWkZLm35TwykEEleZUQL2ixNfBn8q3P
u8HIoa6RBhT1HYEVPab0+ENbB2Z8b1GjiWp2abcpSQbUF6HLGRBloyOcmIiiboxBn6gaRt1PgMlf
CgXQlpMBJ6gQFlRMsSEDoAW7n1VqnPuonfkNYGFxzuGuxu9IpwnB9KCtSCINC8x7fGRS5y91SyNQ
p+L4Cx6iIlP6zyHS2y90i7cjV2g2ozSEflJ1o/4qxzGOXQX9ETXba5ZgDrS92Tg/7uEMkQNGqvjI
nSXh32GkfMm5gQTDB/NzSnBXaj5dszM26P7dsxPwW0njyZgRRqSY8hgxXKcRYqnEaoM/IDmfuhB8
UlUamtMz7kM5K+w5N8uaLm7lbdp/bJH9owwTHuT4wBP0460aavbLVsbTcsWq5I0CqGisgr4aJeCs
W44niWkkLsmU+MJv+wCxHMlbWlVsAU+FDo3Miu8wnGaJwjAdRobIz9eoz7TsoCO5G3iXAlrX8UgQ
1YlLMUejdWICJS7Lo4CoXumXXdLGeiwd7n53Yl6Horz09VP4TYzo9dtx+TmrxmdGDFF5qZgS6eWH
7SRTU8XDb4OSrfNj+I1HmFBVREPMvfDGfqnlhGb5Ctcl6QUl8e0KTX6lRGUEFSQ5oZ5k7jDHO6QD
kcJ18O3VaYXIqFCzPOWVSJSCOTOlPima8d12CunUcPKogovnGSpW5IGHKoaPGFtDqckQOp0nvg32
Gh46IBZXltsuYK7ElolYSgItE+QpAC22vLe+dAK25BVb6fCt9FnmNg+7J5on4lh5PvapMFWYFugJ
V+4fS+nb1LzXH7hgdUV4hf6ME4AStOf/aDk7n2+5HZvjavyGnI0pPsFqH0xZgHz2KpM+CZH0ftmj
h72qnGMX2DAvDUA152h+L+eXpDQgupiWWLawBxphakNM9//K/grU/tG1QLN7Dv6Cq8gIKY8wGE8z
GUfvx4QZkgSjJLYKuPjg84adziYYLBfdcZv8M3rUMGdUyoQ87M/NeI/653/ESyi0dT3MsKSVdakk
3jsT/ekqAnfZGK4a8j1OxYleUtDJeP4BMxPC8QArcD3zYX34LtjvTwb+2AzlPOlDy6w0xMZP7Sfu
tV1saILKhLBh8xJvsZGk0nFJ5Tm3wuMYE9Yc4pgOv8cXR4p0RiYcwz3sdKhzyYKaTEplZy7skWrb
HYpa8j6x0UdjNQLyJrA8ForyaaL+/yoLHGcCxQv/8hwWc1NbfwB4e270PSxPFDdFtJCGojru6zLj
BvplIB0s4iY2thRHR+yD/sS5oWRuYGySvH0ypxVp79Evz3lIqYQftw4V29FtOt5IZEIiPmvUWzQ/
WOO+1wfRwIkzhLKWtRovI30Hb6TG6NMqX0lqRFfUqxjHSRl/cHtiG3OizSHfxrH8iwdVfmxqeBpQ
CnCOSXLk1GEg7jc2DD5TqVzm5JSuwpfeIEvh6ROJNCnT7gYlOBH+8/quVvpsyvZrk+HZAeqpKFHa
v3WdwpP01jVdy2hZvp6Ise16uh5GBYiMqwrDXhsxSo9ThOpoCJUtDJa2A0iq1Gk/vcs8fJB/DcyH
yh3t+cmof4RMVEw5G3PyZQ0LiHOiCkFe5JEx5fcd+xBgA6SGfsK8pKSOTvQJHxOh1X/BVt/Fm/0d
wnGFq67MZlpftg/flV0478HEGrMqMm4cZ+6F+KmT8tybjsV60AH/0SsyJJfhhxOPd6JwAdfT9f0F
mWa9WtDlkO3zPP4ARTnWSKBLeOLaxGZ6jyUwXTDX7/bz50dqP+E2z+u1Vm9cmu4x9Xy3WFMbEN6+
a3QBpo1Aj1BrBNsGT8aZJ8ysfBozGGoq6X8r59ruimRKDe/fcZxCro1KjIui5J50+JLJttH9zWyg
AA6rouxxtofqtyqvkrVemTOryJeRq7P42NhKWwApYL7s/A4Iq+kAHfEgn+h5fb2p0CrjJcDMX/tp
5g49Mrhw9tX2Oi7atf9Yhku5kaHV56yGIIisjKYBvkD5Wzg6+Ok3t97W+tkNwb8EotX6i6g0A2Z1
0EwTQChYwegC9BrqN/Mjx+sFLFHBla9zyZQrvO4/BBNj1zXhbG/RZT4NYMZ2o6CZtydBqJLF9+fy
MNtfek8t7/lX9fK2eiardQtFnfw6pt3qHWhdbvWy+BrDypitFdI0ozcRfrDF8cJfO4NGamLHtOFI
5KrLDxOeUNF2sfPkG1kCSp35xcoVn2VJfRdohG2psZ4kAaXr6HYT1kWEpS6xKRXJGEbhTbIStR6x
Zq0x30hzL+nDpX+M+RIzP8uB2XSvXZmTcrlv9UR3M9lSOQDHaKwLoWksfe+nn2dzxRfIdtzlbumE
QGi+Zo4aG6SCu7WAAXnSAlpGQ+u645lvJvBCLmEgpd6t9/Vj/lez7bwLztX0ojrsSjoC4BRKdBi0
w5DrenvUR12GbjXNynvAEJLITRPkUHy3XDVByWxD2f3G1+mhGECKuqiYKyOw8UEjooR4rWS5sU8/
3BEcF1pA0huFXr40NKiMskzhLb2JYCZf8XHqMuEdWK2CPWGDVFL6sD5wx+BDsnrUlAn9G0SFU89o
+BNNNo9Zku2T16obIOGKecbGfhAOMwydz202RiylNNF4hQlGZmi42qoCk+N50SOe+/gvENIwElCi
udE11dvcS2vQLdhh6gITrKF0UZaB0+7JkA90xMOr7O3YS6uvkGUOzzKdr3EL9y2obnQ0lNJKwHiZ
ua/hKCH73u3EGb7fYuaHiOWPdN1PEdiSD8lTzgtwsKvqVmbBH97s3/I6lEa1fTK0Jii5Rx0Hwcya
+pNZA5VkT/EVbClslwYLgYQ5sqkNfRUBPUGpPdWE9qwxmS+IvWaXYRfA6Plxglxwrd17nHvwLb6u
XUyJKVyuK2irUYmiWosBXqoN/GMI32Mpp77R6K2M7dtQyKtbhH+rwiKJ7UnSI/7n7KEQzUPoeXBK
U/fW/Uz7RgeVChwTmYcoMLPHazv2gsUNn3KLDnhLEUUOw9V6dY/5u8neIUhfVfdOwLyWdeqGukQT
ym1DdhMeicLn+VPGrG2cWJpo6hkoZ8PXmEbKDV4t3HVjjgQaeB5UOPl9PWCmbT3JLmp2yNQu4eql
/apLlpJX2UVS6uBQMZJ94vpq3vTqmQsfaLzxm4P2i4tfwd2zmTZ1iKNKLmzJRqMtRid/SRYT/lgl
iMKlmyUHIVB9/XGIzVzTQRKNcPbXGP03IBE2LWAtjUpCK1SIwwUz0CkF1suAIXdE/qTMEeGmxy2H
X+UC0UhsM+Spa6mQ4QZVPDgsLOtmeVHDpnSva4scx0vDhm5r8e7jrygNNIVMwQFyfX/sF3VeOMmf
2iz1nPHfkC9F0J9p8s5T5IfBrussJ33gZLG4vNOb305oqhZ6p9OJr/2terloLCKtpCm3RrXksj7W
ha0+9Mp/GpIeck90+AOXPuraeiZrG99iawCd8Rr7xJ9FQwcPxcOPXAnwcYuGhTjFzYBgKAHWwlFC
IoqnTevTbVtO7Y1dWNitPrTbaa/cpY5jYnE3u2ji+ulx4ZYKT7OclQ9j9soGf28DOTA4L5NpZm04
KL3vvkCsOrsM3t/ssSMFD4MUrx0G7y9jooMsNbB41FuYjodaNPH4Zk8RLrKZRNH7BQrFrWOwuQ55
V29+b9Gj15F58PWgtMgG/AbmVFOWODGvP8iZ6dKwEQJaDQo93REu6tZGbpkb3WMEZciJZtuePftH
k0+ajjU70CVgt68T+ibH4U8FRNjTBz0cJeES5wVcz/PG4NlRYQ73LkQzQTpuvUHQEgTa/JRJ46N+
57elennByirgQZI38laczYfrxfimMjDSPBDt+WPrz0kYLsTKD9XKVkIRsq88Wnr9CrXgdQ57SeAY
zYgK3Rhg4v6kT0+xQYomkQGzG0gdo/rVQvUy5F+5i9VXOPZbmIglF99EWgPCaEwMiha/M4JVysW2
9ckkCULI2QQ7uc8fp02hcvV8aRVSNF/qwWk2A/2FoCHiF7HnJoSWFC7TZnTJr+dhSevFrPcmOcPK
b7ukYEbKCsWz5XKPcoYieHBv5Pb/iTOjlIc2BuFAL5PefLCr2iQhs4nchnNOaIg/2OCtCLtULcoh
EoMET9q3kQ1QQPtWtqVSjybq6z4Y2fT7KSb/isWvU8Yp4047NNRbYl+nSc1iJ4Kifk1BwxqiFVo1
USSBL0BO7sx6Gl9Wj8j7oL3w+FQxKJ0bfQcEtP7ujESURRG/mPZBDNrIK1fK8JxQ92OAhp8562fT
hBCqV6tUqG+IpBx0U2oIb4emXDST+K4cBL41vrzE+kHmqJv8KCv3WKNLPJdj2cZ87grnSoPlNb5g
CjhfjUDXRloofE4/ES7PBYh7aqBp55+dCpa80uCS4KQXWne7zpY6ISJs26G94712cnB40/lGVOHf
GSlu5OZ1zfmEOXW6tgkl0E9L1Vhxt7LmdvMIw534mn8EkBGKIsOxNUuyHWXAPJhzJOXRRnTk2M7K
hbkLrwoYjEDrR5+wSoGCrOSFQz5XC/iQxbTBbPAvLM9fQcEwUoVkZfacPXyTIUE4WP1SpT0eAk4+
ubSsgVnBmpr+OCuZ+ijTBTkdH+hym8YZDb+f9htcQAW1v66lY1c64/XwjlPwV7rtUL7p0HCzC09B
b0eLjnYjgdNidyKu1aTHMRe61DFmrw4R8itq4AWJq/nCKS9PGBczoPHxoQFXKHGCgLIDjX1FZNit
6J4Dwg7Hixt2nKFHZhboUR3G9GOirxLJjbODLsCe0IXJYa4DGTnTVBaQK88dLCOsPYax0eapA5x3
d0gDbBpqasMHMYUaihHHf4ipYsfdJ3qBD2ChIr1eSSd0sE3wEdvAaXyGlwNSfcgoSncKA38jPPV6
y2qhBx6+6fJK//7TtKy95O5q/La1VOTRizZ1OuhTtXQUaxc+UNE+4QwSu1phljrv+F7eRl9BRRoR
iRK3aw2PRG/+9Sp0IMmTB76feXXUMcMECkdMzg4UgmB2Tb6qpVU1CrKrpJM3hIDkrHa44iJ4W0GW
N6gLUPVkm1WCt3+I7lWqgSxMimXik2032AfPPAHSqRJqNG17aQTBY9kvA59WnTpgj8Da5ogYiroe
8MfaiVykwPKlz+2VkGGEX76pl3FwvFcgriAJc6zw24cQBABqdXtlBR0RzptTDZ6xDW9dEjQdBPXW
74vQks4UkcSViNh0DmQyfS1e8YKCYtCSOblEW/qMMouwXyh4HiIg3IqGXbvYIuFH/0wHHC2cQAWi
aDdfb3fn3ZbjcKK4+WAeALYTCSN4G3TmKuda/bWzt/svcu3Q2B8uFB1aheElBpIy+HccZqWLCBfq
LugVgE72pqOFi4nTKc72DJuyPIw8ZQR5k02zAU1Robi8swR4VXQfiNHS1g2eQE99IhLClZH/dBca
6hct4afnYNLIyhER0quWItldM14Of5Q8TXqvVkFp4jcllXT+anjuW39cCpaV487UGnZgGXI7RAj1
BbAHrJ8I8+1+zIKlWsHLxIxKyVuwLZB6YUpKXBeUYmn2GkDLB7wA/+2yIjG3I5GYlC8nYp7JK2xV
Dp9LlXYCYf0VBxx92tglPJGKAZ3K0+lavEljH+f4DFzLukuAw9MD7TsYx49Gjb0ko6FD038x+xby
A7PA0GSOgIeDtjZ/xEWhIv4eEJuw7GXCatL7X6xube/gQJXUVt1Qw2QiKo++xKTjPtWesIeG+zEu
Otcrdbv18EV7vP0VAh6n/CsOQ3PyBDXM11isZ5mHSzPybnS7kLhurO+G5CxxBl6ZeUQ+7xbz0+Iq
v9l1CpnQGrlaZcdbzKR7oug3HUyagp6x3+k1q534QW3TGbvhdfYMJW2zVVdJM0fFCQ5oGXBsK3Mz
LqmYbqMXPxm1s3AzjQ9M0HD73eA24L6tA4+c0z/fndvBm7Tw7zzTuZyjkZpGaWYCwP55LW0I9nCB
GyuDGJRVDgoGZcFmhUo1QHvkm+Itz2um/ENIQAsinAm54UEUK4vMQ9EE3A9Ljmedqta8W+oiy61V
//JGIySBOU9n2NiKyK5q0XQMdgtLwMMJRiisedlfODjEk7ONYNDGRcV4O7tu6tlA3h/UEtTEmTvg
tCPwO9EYMPHz7OTsDZlxkAZBkk/4MSmXN/XXY9De4H4cSAnMsBOeFy919HfDLadGH5du+y+njJ5Z
LJFBmunuJNnXJ17I4w0l1rXCwvZQUC10gvhim4ATPeZKjMO4Y5MZG30nXolWokbVHopVYQFBep1p
utPCIshesYNvCuev+mv635TelfDyXC6tRx7ICigmrEj8TQuro5LUBlFgYa9GAiveRRk7F5fq0qxy
/hd+bZS3g2Yxxt0hFcCnqPY+lKUoot6T19aG2mraBknf8zShuczXUxC8Rpw+BWNyzR3H+Sj+QQlB
1H6+L5WKXealBLtiZyW6l/5trPzbhUzI11gMLGxVnbnQcxZD2nPLH7h0Cu81Dcva+rSDXHrSVj8q
dy6qtMXy842K6bHRYq1KR+flPAxPH00HiWonE7zaPKlvcT+e4Hqx9gflAHvzQkzB3wM4Yo0WxziK
We5eRS97Tr2PGyZ+xXwnKlN5PODlPPdSpRimppbUbehJExFaPdPDdXcuK+sePp5cAUp8q6eokEgO
2b1lnv76H2/nPJGT1IYw2LE9iR8oL0vuBb5iouQ5Z/W4jT5yHi8adku201UUYIBi73gHHKhjCZrb
cOeb1/Cwt9XgfyStU4XfuY9X0VFPzQDKTRIWhGRBlRkqIUIN9wHWBuJfAYw7hto6xw2vkJx6cjUa
yh2jtTQ011L9G2lFmMxYFeoELRd5wUjmWx2EoUNm1f23wuDZuwLwijPBWw79OJ+BQvJYMa49Bn0n
APTn4BfyYUU0xvb+VqUsSRlV5AHZyvBahEU9fkrsA4QeB6kU/+OaQeLUA1Wp3owesqUCMwroAf2s
BjLbLpSsApsWyl+EreGBNzcbxmWbukWwJE1IODjbNRQdpXPjRCjAeMLvhsHau6B3js6Gd+kB7hjz
RyneqwTMI9Dco0XYMLTok0XAMX+exCCDKFOcMxfp6HagYA4OIzi9H6Ht9tJruUJpCjzpDKvKBFxv
BiFvw4F7YTFijFs91gMifmBk5Yq+8d9LQ+XvEY2o4orSqdM3h2Viu7BsN5uvdCFZrSgUnhO3mgQd
ra1NURojcdFQNV4tVSctDqmDVD4c/QNTw6B3j4zlYGKeSapqvZMi6QyjCI+9wKF8SRtOXoh5vSkf
KFvKGs73LYUcU024/4bwZ8meb6RjRrrv2d+JIlMVne1bEMYBJClMdZIAxUBxozRL5vZdJdkoRxcA
2A/mgIpFZA7F+LbgcE/VimHv6XiLi9nfQkRfiDpBbI3HfjzBnGe8xd+pHdD/ltmtawHfg+ayF6iv
79WYJDfoa2sHYeecuY2ZvJxo632TzhnTnUHzl6VlG1t7FKmyGgRV7pEFssMHu+iiH4p+wC6gQdCV
gAq4oljEa64IZYud/ogUY5ie0eLdYs7FkzGQMyj3F9QrMED7bQlmZOHQsCh72TRWR2GWfNKjiRuY
P47hS+Qqr3z2nWz3f0xtN1jiuMVL54WTcg23T2kZusD5/XGlU/SsCsoOwHvOSjPFmQjashSpicdV
jnA0ltoC7zpaehfM/HKgMGtqMR0uY0e92I7bG97PwLrrIGFbqJ/AE2RCop8woknKoBZNQP3IBAAH
Xc5J1x7Occ1W3aWkpGYI25xtNCNdh+KETNf7ywGlfHTKUtYco4/+gKN6InWwzF/Lf4Sg15eScddM
aHe30ZBkHg5lIV40mouwdBlT+pjkxvPxoZhHbuQr8Bn5nbJ7mI3/1t9igRd6+V/dY5O057NKScjR
M5ScHjODdWMVGRCGXr7RcXeM3Qfk7o6Hw8Yl9B1dpufhzNL1rTyrBPzeK519Mti4FxOm9+tTmPsc
3O7OZquUabdK1EZt2n8fmFRrsPK0zYt0Bj6c/vCgGnjDOOYmOV9r9AI298zDlCswQM3TNrHYPP8I
q9drA8abac+zC6RrAv7lm+296x9P3J/O2rdgajpoBcJMPQhz7fXfI/2ODqxZDa/FfnlyUSYLTjLn
j38x33Sr5dD/NM4NbAGCUYdk1H8qiopQsX5iGkJGDbD0r8/q+2TDoy8ovUHws31QydiysrwRh0ac
2haXU23Fx/WpDL3J8sH3+txtEc7K/GQGAIOw0PtU+l0t5NtQCOTvtGrvkxtkDMIprRkArjgL+3jg
0bDHDgwgXWb/tJi7FwTFkxCAz/m7NOf9Hqx+D7bEBQ0Nfyy6J8rhd6DxuravIty8pLniwKY3GOL+
2PwcBUmp5isWmCnRYpqwB5BaFObxr2opU1o9ILkPe5wtV0WufpgFZ8Jwc+EShrJ1UzPJWBquBqnK
reUCDwi1VQI1yleQBW9unS19eSRh35fLMz7ItP0jiLb2xuKcxsJz6/rO+uSDOs01Oyq9riIfA+7d
wybsNItK/mGYxN5COmdnSKHzmNoKT6QPX5Z/oldNq9Bvum5YLJEXfPpdq6MnIBKjsSAnylQrgq9U
z0RVyX/RzbOwh3sVC+3KiYKxmu9Vttx2vreIabVqfo+0sDCwLqshznhfI00XnabSE8v8Zx7w/Ors
grpxdspUKYqtmSG+q2UvSGio4m3calWg1odL6GsOZTM15JnGhFlN6MJSf4qjiK7PPwQ8O0eIvBYc
vLwp6ei1Gc2ipIp7tntI0FupBxRfNuaLDpb+pJgCvRZNLKGEJH+PWcw/6w8CUsSeUcPM1/tkDnBR
nXx4xetbJQc9xM6Ej+e1SeY/b9mAZ3N01uAI8UjuPbFV5tJB1wDuQ4lukMboXIs0584P2Zc8OjQk
iRD9oHEXgVeaLPTg42JzH0xT9HEh/nDfTQnW8+SqqWC9afMoqIiTOqIPNuGkYJt+lHmUDNHa56ul
vyd7i81B/qQUWxV80KI3PfBBV9AzNC6+dxfLgEcAf/mtSZY/LSKd1Mx+gY0hgU2bt02cqG3ewz5X
J7hI9dVJT0W/jOX4X9WbEc7755Q52vBxXp92edkn4AlJdyczHAA3/Zxm8P7PY+X8oCjDiJ3bVpAF
gjMsalU+Z1IMxs+RPx+cLSfGsFulptMhQXuZldcNUpixt+SJ6fuwMk5tXOM1nzr8f7ifE3VBwlKJ
ievke6Z19PEiWtmLe0k/FsrcWsNCCk7i6Uhv7PkY2REnq5BPkUcLxxRQC0XMCOuyyrHgU1shmmyW
RYzRqai7iE4WlzAAOY4tXhvtfVbM7xO7TTAr49YFXrJPmHfQrZIabDT5HEMFRrZ4KK2Ntmlo1cJV
UozdeFfnhG1NU0qlz6jlDQYGlBw25LnCuisM/F7VvlP2Xszs1UIaObZFkxfNsOVXhrveVvn6nbxx
ICN3p3zgd8Azjvx7Id1VUY57FWJmiNPIKb3/rzxFTcA0n7O3us8qXWjGpkdXJ42oQQKVGHywp2Ob
Oo5RmA5z2NNJ6ZSv60adtQVd9FdqFvhfQjhhW5f7QAJ32c/krp5gkkPrbYKzzQpVdJ5G5ex14TVd
e3/0cphn25vOdI/9PSiuoCAriyJ5Cl1KMSNHgj/NsJDKSInko/aidmgKD5kKL3Z8DrEX1ciWxHh2
AGsSLjNMkEBmyixxOcQEiuVv1GSkAhjfyb7gGbiApjmuDVBwixXGyG3GC0a8m/BZw5tTa//JafoZ
t05bPN0aOetJHAivgh1/u3vUcx8o5eg+adiq0tch9DEjj26NUvBQoJ2xAZjDDmAXx8dU0pcMDJd5
te9PmL8BI8InJmoOUlPKVKKGUQ8yxDZSF98dXLuj2Cu4E1yRKFuuGPrOCR92w9U2AmFzylokx2n1
J01GrPYGNDqcGKg121sjwfQoYutLsuWPN2if7QhbbmTRpCYOy3jI+yRrt4fwRv3KQIZVS8/AUI+r
9iPH8VgSedP/ULTmpG9HLS5wJUmB63NzimR0cbgmmeEYB/YoqUEZw30djo899yjDWdGN+y6ubjIe
f+bvYqF85ETW/moB/AN6jazIpHYgdQIylf4OnQR9AtBZrtP1LjZp3XUkfwEv1Ri5VTlk+ush1tsj
I8seGapUbehNoEYcRYpBF/YQEkkkcUaZK6neac0sOlgpnJEwQJBfxUCZfs5tH+x1xnlSjHQVMCLe
WVYXqmJciM4tLaBFqLICMe5YqQqX+djqcoHQrLZ9v/bXWoy9ugIBggXS4XfgkFVrjdt3BZBAl2g6
6QmJpyk7XjYBicLNqy/M7SwOg6ZlyJYAicE+wHuMAtq4VW2N9STHfHOi/ujxSqxbIyYC7MO60SxX
SbYTWp3pK1WkKxI9pqaJudLDGEp4UjGGIFkemunzA9wJLOiOBAfT9gmrE6HPwkz7grfOv4j2oa1L
bUhvMaTrVe1+DNCoXWRf252OZ6QwLbkayMdFgPBBMsF0KoI8A93YYTF5Ps6NGQgWtKPnhW3zciz6
66qwbJPVsQ7poslVymkeJMjWjQWu4wSo0R4a9m0SJZL6B4jtgxguVxLDts/XXF3cowEyAXR09BxH
CTl5TyAMbb4vX5fEu1olCUuEi2WIZJRerskksJBiRIyLIeuX/2HoShwm5B4Q0J5Cn8sVn91ht5K2
RSN6rxV1urUzvWOZRF6eOphuyq/qcqaTUR3pAp00Hi96qxZxRC8saejBQnDayHWHwTh8bzTS0dA7
GXl31OEz7HKjJmSwGgnmxThg9qc5jQTDk/q/C9euTRASMm+4d9yzY8JbCJlEnRGSO1EeOZgJsyEd
kfy/T6l7Zbglpe6PoAcujaFc2u/Af9fdqqfWrQ9bN/DBaybGK60cXT9xYAJMU+m01YXkBdbqRfih
238dnbXXPYtai/znvS2YPJU0jCvQu5qunMVwZ94YOa/AC+fFqbYL13iKNrpIiDz6oqn7+lv60O1p
vOKfM53dL0RO4Qb2LBs322nzmu8uhjb0+6qlL+NfVniBagdMIMqEkp2sOaNGro/bA2rjgtKw53qs
g7UKVZZ0NMJeIAwZedLeD0P6XJzx/k2KoFaTzHUF9iO691Mm1iCljVLAcJXUI/L3XtMZGZCiMIuk
5QO84I3WcNAAby6sCbz/yWBNnaQ3/V2rs04zQ9qht0mxuIAE8KW2pPMrDG7j1q7I6ZiPkcUEKz2J
NXDr/CJDofYhOieJnOWctkzB9+uTjRWbFi2natonP59d/8o3Fs3Unj4aEejzG7z3FwrW9EbZG7K9
4PYcvQqNk/SVWBvPde5Dkqj8uCD/PHkOuXkBBT0gn8T6zjGVh16+196dActhqm5/0RSIxOYrYtLb
S+W1FwNbInoDLtkeVclESvZL8EB7U4ulioBLwoAmUKiqy4x2K9MXmFNgiFTYIThYz6VDq7y99Sxb
/0PDIMxn3lUmntgah83YhF9/Gb9CJZAw0pC7QZJ34nlsNuT+4TFegnvIbHRoxY5Qduxo+epJMfr5
KdWUeLBK0iPpCqbvKzeBa5X8y5UvOQUsUu+xTRoYEdvYaK6Ckcuo3J86jYsSacs1NcJjzi6Q+ZHv
yCbFCLJP3dwpSPlx2XAlWVguIvWRgUKNTPL5sDU8Ql9xixWBW4oZk5l9Nr0Lx6pxfGmAfUKzkx0Q
CSQIXELVrbSLpnNXy1PRf9sWQcE4g1J34IlcwYNcb6xd3G+bWWLmNscS6+Iqny7gvT4ZsmdiYApA
NRCMjq6IHQmy0fMyCX/z9Aq6d7L3hw7HUi79xRgrga31suyE8df1ZJHRG9LtMqLSJHXFT/XS+aN/
cmFEZfVIsFZz/HsD1HqCLY7Ufm2dcUxkIZajXUqGm6UNtc6TMZhSL50YYmABQrqHete+neMF32TT
fYNmILkN7CZnVac8ctxn0O+hn1Yense3n4n1pXXYkRrHCeFoIFxts6Eb9pfifGhpmuGHlaqHo04k
CMN7M5CSS4rLZ8gluhLFmYPJyqk//6YXoLqsuyKZD+eBINg4K1i68nSMJNzocSU8sf8KA0E7+EYs
cBJSJX6yTykmh+xN+sVzuOsgbcFgsLVE7vs9HpY3nFyIdGpO0pfQvy+U6iykSgLVNPHoy7RqoZvg
u/HT5PmM6x3kbPceuJ6VEbll11bb4/g+amMFcAB+5nYkVqwGhtDAHSXXAueDBe2jSXeuUaNqDpwO
uqy/sz2c8v/wGUfAz1TC9wpzFRedNgz+tWZuSH+i2/7Mi0DfmT28SS4XaEq5Dv1baA2sgHr2Aq0z
ZjygZQuvfe0z/1FrgCKuJnaF4Lo4P8Gfk2QiQesTG1OvnaxTI/1Q0EU+GErAoY77jPgtgHnUo/KV
avAHMXnT9W3UaKlsE+gZqYQgS+f/p8OxZathQyjpflCvBdVHj0NPU3KezbWvPIB+jJQVZENUvjEx
rjE/NjNuNRhOQgjheJ/VXEY61R/GfUt0EOYwFL8leCh2HvUQ/beegt4UswHfUwbbIK5K2nppHe3B
to1y3GFmI+KgBXH/f1Jl2TexiPqCoA1wjWWoMF4cQLTaetR4vxtwg7x/SnpKPa+tcYKOnykQKzCj
jC+FD2fYm0yHdcbEomPb6t6jUYJX+5dRT9y2fRjbHHhLhlpRhV0Paql5v1x+yzIvXUi40kza0InD
UXxnqpVuBMwBQ/vjRA+OjSwjILWo2edPiKSRoLg+gmKt8KbIUueE5mDo660cLiuu4VlsAE7X184Z
0O2eqGqCY9PHapNfMN4d9fuiEKkJY3Te3hSH0mhaaTnlf63uFrMgDd/TtyxSf+dyNylRbCcZWPTJ
xU7qjXH3yduzsnqbdcPn3BhPBToNLj3rKc1C3WBbbJaBlu/MBLQNdhrm6uZ7Jsnu5Dgu8i1Bd/NS
2ewGwJqNrK2xDM83ZSxL9vutAQIU7t1lHpP+2BBZymhYyNeEzOTveZC+5bNmfhU8bMwyf5FfKxFG
q97Q0xAx6XciqpCmvSATvFV+L0ySOSkwJcQdeteFKZf674OlCNG+GYsfTcu3HMQma9CZlfBGBhXk
Yr7La0uWWNH9hyv3JtBHmp9JXnYGX5KTAmqHRy7rq//WUY/R3WJJUmcc02kCuDoPA+gCRyK1XzP4
2p01RI9qQw8cNaatI/hsa1H/fBMi2H4y7R9B5/h+596VI7Mpb0y78lg5invFIa+a3jzB1xd6O8aX
r7ciT6JJcVWCxLva/UgJ8oD7H0o8m+jkXHy0zw8LbAYdQinv6Un6QkvEZHjWMiXr9m/fbIk1GSVz
PRI5pDQH5fTKsYWmlUwAj70rALynPgKp9Nhpizey/IZ8CzzOYw92DrJbbr8e1FUB7hsceMJONu6+
JqPRcyrIk4jMs5+JbcTvPs4VLMpm1hJRDE0/z5T1HH5os1JhMbIW2bgbx9FFFIYtHNVBz12R6i4T
wRmcyE7lkhDVZV6P2HC/pRcIYjdqynH/wGrF2dnwUZYDZZscrmcLgvfkNfCHUX+wcor+jP6mVI0x
Deg/iEFaI7c5m+TPgPtMbKNTTWBRmEi3NKsWfsc+SWQQ4aKuwydCNfjnEApgmSItAEGMpumhEZHL
LouAFn+YNZOXLXRt+hcPkg79Lc46knoULGLpqKVqS/jK5tgtbmP2ccL61A7ii1RS9v9CDQCeFfXR
SnATrucpmwiKr2a+boFils+zCaTcEk3UlW4tW8acaXdBcaL1qBnm6+SxDMf+ir2Rnv206CRImXSM
6nf5x9/fBDd5E8LvLt9DO2jAODgI539TDcfdvj9drBBIITEsBHlg/48721E6Nt1EoUcyZwb9pYk/
uKCRZMMtDv5Yl9c/woyzl+KC1+0uzsakAGd3tOHUGFWTyBqtQorVWhAdfvUbMQONXlSqqxnArYp8
Mj4k+DY5sJbGBBPs/r/79a8ATi40jSXUZSSTVRBKX0d3m8H4QAqUSC/udek6fABAhqj0j+XiRmGn
wr/bMrmxHd/4Z61A3MZTS9QqLaAzloBVy0Tmx2D2G0Gboa6mKKfxWfvMc1LpbyiWuegC87RqXp3W
2e63A/09mvjC5KkItt44ItMSQzuIFdj0HTxjNzXGcrkMdfiwpXVFEbCUOgR7q+uoPOkXp6nilMo4
jiphhxfrqSG6XdTCSM0liANVOKyDr4kxiq5rTloh6OhtwiSD00g8rTQUjWeUL1LSx+T1W7jDYq19
FnsyDhYhif8BaB/6VivFlwPGiyYMdvY8KnInDVVz3qQ5YzPReb7C3G/R8V2HwMT5YOI04cHXLg2k
hJLphxCAY4bbrJZT9/DI5bicVw4dQHs7NBi+2QdxvkGeB6K9jCjktTMylXVdHgFXAH8sn0vozeFt
LlJtwOV15oSc+k62QOEAbIAQMdm8R1jCC4kPIImgcJ2OAL6tdv0Ov4cS/437j0M0IZKnk8iA6KLv
P9qU4S5j6Bea1HHDQ5hcXP2izG2FI/1LO/aEzyocjMAa3PJ42Qxle2azpLIkgknlWuWymD6OQNe/
+KvKBUp+09Dy3bvfBvuMWp++RQ2GR77NuWthzG5fWzNqRAvFm5Nm1UXEOm3YscwElv67d2P+jGQn
evrTArKjo2ZdCQa4Vfepjp9ys1H7a66F+K+QPf2hdx4oavgaHG2cDDdUBDwkp86OqCAfo6CT/2bX
zsSvMNiZNv/eUpUiHg8tV3Mz7SVBX/TMw34zq6KuUTXPKlIM0oGdlqdAYXZMjNXeco4+jyHtQa77
szG8APZ6hf9U6bTSVATQyNQEHFOzZ+H9AieET2HhocYLIs8iWqNDue+MFjflJj6TXBuQ0yJwof+s
4Y3LsgwnXACtC1bcu+kZfLWcZHUg5gUkYf4QZVzDaNCB6kTmvHUtnBjK+7mRCoxXpDkJj3bOCj36
s2L1v6YUAi0fV4GYXW41TgGDY3ghdVwfB3BZF1q49HYmgFqfVGIeoa17oLD3/gCoF6vrUtQuPjTE
/2TwfwqKrWk3/zcRH2C6E+Npi2oO5EZBUWepobl8NzyXtPxlCaGc5HYdxigiZIzEuCaaRu6ZJ6TS
OxFtBakmbY0Zkq8Pjzf9256Fdv9BqdIjRWjFQOuFbWxsEPtahghaDM4bA6Qn3a7n4ew8s09P08d9
5M2AJTzICl1mbB8y3mGVzjlvZNPdePDMWrjSaMRf7+4Hc/53XwFHu2fZVkgzfo0ptDrWW1TVXeeT
gG26qzywOrfMjhtILJ6fG6C48KekNMfxMUh2DijOsKDGCkfuww/a7JEYt41pZWc0gEouQnz+b0sE
iuTA52sPAMcFr5gvDq8GMwpnMXlVyNMeEK9Gyt4U1R0dC5YZCI3g9duRaM4EYTFgTU9OKiGEfyUX
bbDVYI3C2Q+iSiBEBip/akfCK9kTgvqVGP6g1inK1wVVpIEDV6XfqQ5MbQSM3UPa24pAvLnCbcMi
PB+XiOPNEO+kAYhSyWGJaqnOCk+An6mxY862eme6OpQUOPCy1KptpuCz+ygobSVP3Z9SpeLN2xwf
z53ma0ozpjuQ/B5JfrQHCFm1IChXdGj8GKpWULxQ+wA7/m1WT3Lj6V0gI9XV9nHhiZcS2ZIrEyLM
6l0cauKJCx3UMKK1KdWiPT6enfDzm5COQ1CAibydA2E+syNsZjRlgWQZ/PPtMW0DCAuc0X2XfpIj
Y7ibx/spUd8KgcB2/OeWDMKii9B5ofv2EdZq0CelBNd6PFUVBZv8w+1SF/da1FXNehCxwdpV6HlV
eE4SYxg8izu93K0OVUaCqgziguFNwgvHpuzzrf009JBHQdT+bzwlJwbi/x7xUZZphRv9M426VAdY
wi10ryg+DLN0PjrEs1JQ7NyrvqsrEYPISsMyrRQn5IjbGJN1oeh2RhCKIhhcYWixGZW13N/t1FYp
Dky8bcTxI4Jr4MyEiLa+gW/1e7sW8OK6VtQUX7bBL88uMzXPWdRD5vhMNhJTMZjaNlpAarj1cxsB
0hau0zT2YeoRY11T6kI5sNSWAy4pMX8VJ4XNmvAyg7Z6xxZVh3Hc5rsx5rKF09/vSZYowDRUM7QZ
nT2HZyfb3LBK+Fh4c3aOiq8z7d+1jQeyjZS8LIqdtSHM5Oy/aYmDM8TJZZFuPs4cM4w4qhdEsMZn
NG+l8rkQohiau9q/T999WrssumOP2EG6J8/HiqEK+7SzYYUjgpiHeIfEwXUsLpIH+7P0VJgJ8Z6+
MRxolusu8teFMitDeFKg9XNpIlWH/aVsNZAzb3OIWc9Wh0OgeWUAVI2zGHu1YSOsRpVQW+33sq6Q
jItfSf/ZFfaBvgeVO9o+JSU7A/Hv6JXJWk7SQXdeku4+YYWXbop5j9eufEpN3iNH74mt/V7L4biq
wPIjsOGfByWrptEO6X9eS41J9e31hgd83HVhvKoehE99Y4zUQglGDqC6R6lIoUXshrpy07NizmR3
PEbv3KzdN4jlbHQqxDMDbJ/Ck8iyuBEQuQAuifneOLMnyCfqoizfIH1T2HF6s+Hhf5WBDRHM/CVF
jAt+K0bjgqN9SwFMecPlErDfivrdtwfU76kUwNGVSCR66ABoVi1cS2kVF49oU9fk+K/JraUmYXgp
MkdHs+9O5aOyhVevn4FuvouI29lOln6oyxoZsI7JSwLieKhyP6EHKD2nDDnzQe9HciheVprXDNF7
IPpOEkCm8CauW/Ne8UZRkp/tVaddRLUhfQP0NdV/1vjGrH3tvXci4vmHy0vj/3lGi/NS0AS+IcX5
mbzjoCRzcExil4tonQI+Dwzw+sJBucc+CwyPUx1nHSaTNU4H44cPI0Iqo0G0C3XTaRjY00hZmlze
G/R6PjjqKmpFxK2WCPRjlix/bruB8/n6/Ybtiz9k25qVYEP8zjAyUce+mlhtVIK6+ZUukqREbD0V
UlWpdaggT16s15XE90GNE9RRQkZMMVZfveU8ALrholwx/YzgtIedGPJntdY1TiOYE3JD2R1wAZIV
hf8oZk683Dixg1afIMI6z16MmcEyAyMcatcV4kBR/cz+p9LI6No8tgC8ddqeE8kuQhyPs5geXotS
4bhoFOM44gDeyImXtvnVjcKk+0glKnu1MZUXSQj9EE4mdSJ9reTkNet5sWm1FsNG9RL6v21wE6Tf
Q0cr8ZQo3whvk62d+zPrNqOhvcBPLjzhyx9tqiHQMPuxvDFBMT7mw4atBKQz7YARk2E7ElQ5BCCu
TpnZptPUR3QzbEkOP1Dtr8PnymrRuVPcfw8yN/oGc6KcW8tPnMWkLKEr8KC+2a6Gv99Nt+T0W5JW
Of7x6qsHDThZ/CvNlQJ5uvzItF/riB3UMNRWNzA/hA9Ts4Q0ZQvJJC7vH+o0edYvCjL+piK/P1te
/aqZ/3kepIC7RrKabFvNyrFhOo237aSb0DUeKWUDbE+jw8FEINDwTvPuSVsPDixs8v3jchjrlyLl
iWpvgIr/qak9iN3CnsqWmwfLZ1vKuTyh+DqLIREIemZI9+IYhWeJPqEsbWUPzJ9N2/Seh8dSj6mK
LyoUfGOFvT8iaSiAXZEyIBS4cWXmq//hEc6BDqkcnJJvWDghJmb5+fdgUeqO6NedOLIz5bR5du4m
v8I80v4eaBDquDLRNoyTDzcm34+xttXERqIUCu1ZDFdZ7Pywnk+VJqkQ0LgNyaAgSJUeaTStvWU7
bS3rMtlVsFXmrTiL9BXU5LZ3h/lRlN9NgSFULr4JA3reRn0MC7qLbBE17rRDi16MtGLKXSxzQjTT
TmrBojEb/zS2MrYD0f6i1eWRUeHLUhmKKIvtMT+eFePIGt28N8Y8/UlOKEYJwsAiU2GLLmZn3LLW
Eo3omfNBpyVW1xR8g3Y7lw6K7kOsLSw+gdYdiADzgW2wRBoLlkdhQaA4JwdV9WA4+Cjyvt71LIQB
hQSO2H/VrTLyfisK1YxzWWc/c/FlTZXpJI1o+2U5dXnulhyrMAwOmdp/P/mWHTYuGgATp3Xd/5MU
QWXuddkJJW+huHJ14TR8NPpVsT31rc0y7PUYTcoe1g/Vse9/LvZUE+GK3hzwQZhPmm3HNdNY7dNy
+khMF9UWkIdM/FK80PEuN89nh6AdiA0fbbJ+x4kr3WUqmzGzWzQ90Nce7tKcptTL+eeKwHRDEN4R
soka1w/g1RQyKt+JjvGC5AleYeIsjgx8SeBKcD+MEr1mNl0zhH+wEWu4vj55S/aP/e8PrD87U5Sw
oxwab2RfGzEq4FoeHM5Q0k3o4DC1SZeqI4TrYkFbwL4d7QI9C5dkG5s7qk1cI2Ck9UxdezgaYRO7
CG7eSA1WeOJF7ZjcURGDMxk/hk9mxVtBneecR1O0sk+yjcJDCdfynPjzsocqbGd+TWOtPJYwXt4y
wh72OnF9LU5fmKNPQe4yL3clop33V+bHPhzropQyIV2oTr+TqWVnZLEh7I3co7deVvreeSEQIdKz
l+xrQpjtp7k2jF8r+cmoZiTTkL6+TTH0z9DPjJBmMIR7BSb7xfNqPoeVn2osBqPqFFQC2GU8p/KY
uqsZGDja1ykR5t8Pxf/ZKgBIZTapdCXTZO0Ffi7skfxgX+YCg/be94rwTkQ1WcsUAkqxaljlHD+U
f+y+O0CNeJaxQc53/DwrBCK/hUlp68GOb4Tyq+O1xAk3VL8f0VFeM66ymmN6CUvjkJkyJDDoBrGq
HJDUJCvshsQtllrBMwTUL8Fgc1nNwg/y7pzULa4iZWG4fSYMDbi6vYIZ49UMf4Hs043WTplhyku/
eTokB1daSAa4u0jscx62/wnsOuuU0kO+vzo1Oueuk39LTe5ew79qezg6y1JTAngLCWGLJQlHeMpj
Qfg10oK8c14df5nZpNQNsGhOB2alWrKcbvTz/t9jTwqTz1d1bv88RlrJbtimYIGf7ZLkX3shUSwG
GPZqiGlXtjNMASXi5sCowk7IC8SFV1uA+Y4Syrmppp3gC5sW1kzPVjgZ6kNrr1Pk7avALh/J02Rd
K4AZAeKDBnnvvO/yKv11o/5u2tTrQs+CfzK+ZRfffO8wZfnrvxHUgM0Ugtf3E6x5evShGXJ6MlJj
KWyMSTLICbNmGv/Abr7k7rDwMM7v8XAkAsHSHhwGgaR5JcqV8aL2coIAOQF/d8S4GD0n/R3j+tWy
k6qq3pxSSnNqnxAhRQBx+Qs2CcnZQmrpWzzz6lsGbnxgazkgKqUy6cPHyRdJT8Nmy26f7C9NdQE7
LX9ldd47PuboO8VHkl+UNWcLMPRhPfacgBcHn+xKaX6KT/Dkr8Lmf1IvBiO38bCXmvPw0/C7MjTG
M+cqctVY0ZaVLv0bFBVx+q8tb6VJgvKyIu1u8kp3cX7E9GR32LX/+1xoIaGDLk1dOqKmlEBuZDqq
+cqk9HOetfhbhVIUmpyNPnpxPkOfHETEXDbA2fcMwTW3l22Pl03wdaEHg+6aKeoNOoCa/rU7r1oz
lji1ACo6DmRBL9RFHxVRutY5TMhHA6zRSeV0s8zUbQX11YKuB3c+Ol0Nnvz7K+pzA9odqQEre16n
9Az73P38Z6UHTC+XteqRom/BBzW4TMlMBM1VMCRYqRq3KuVzBsEmgGZw9Y7tNDv6KtRHhrZUdLaV
IlmSOr8W1u3oqoIRFfo5Y1JaX6XRNyYqkHNNIbhKZWKd+mXNhj5CM4jVhERXRko8nl/RnVb7YwAO
1aimE0cZKeQgh12S5IXZNb2ZezLOz2VmsPj4VNUe+NItYcHLvPdyNiRMoS7JV9e3/z9tN9xR+bYc
ch5HxTtLk8ZZSUoE2qDq4jGbuxW+2kGvxjogGndvgSf0QQGh5DCAAd3OHi2VDiWuY+PVEEsSn1jm
ioZBvdBRIHAVgSoeD9Wy/eVyXCALZngSVYeFBikzyDV3PaTLQ+hMUvKVR2nnh14lUxWGrgrZMvCN
U8J6aqOLD7lxkT6Ns6Ltize4R21VESWWxDSn7qt9oImACROAhyam7ECz/4luCf5j8G9wa4Cn1U8p
I/9tEEiBdbA9rcXRHA7oAI+Yn6PAvHs0mYaZH9JG0tqCu+OfxssTHVt1Dl/ZlebaiSOPz4AgXnD/
MbPQLnkG0d5TLsjcJKVRpehORv4ZcV5Xx5EVJWL9dC4QCGp0v4nIHaNFdGZ95MxzUzaumzdQ1gMk
TvO5FAydVeEuQVdALT5RNccjX1cwkB1aqlhSKk39jbnGu6sPD7nrmnUHMrplTS6JtooEBlg+uK4B
7LLxZecV/2ecRB/v7xhF+9tzsQRbHa6XJ7z4LA+5xxn/vqOY9/ppWf2YAU6FB3PAI9OjWWxR/gmB
hocu5p/0sq4KVi0QESqb6xXABb5HdVkN5WGukmDiuJDnkBzSsHWSbswHdmnlWCpVaNRmfJccxatj
8mKZLT0lQtHUj4b12mBdmDXIHk/qoJHbb5VvOCscryQRgU5gS9earo9+ERf3pL08JaByBIdi3mHM
iuU1rhwj7jE1Rxiu6AYHw/yl+0AoFVWFK6fQRlgm7HvzNIx5LDQECevn00/i+qdsSIZ3488CfMOy
YBPPktkzYWwcGfgvuWvpP0umtpP29W5BvvOy3L7z3LK7UW6oZ9iprzmgk2mPUkPRpp/KNgjsbv+P
UayBdORFGfyQuNLOzV6imfLSjhONSLCxVeaSx7Dj2TaOmpBj08rWlkEB2Svb0GwjRulnwSUjwTNz
D/aJd+pAF0ns7HHtJkH7pr4Z3TL2P0lumH6pGzyksxbIxeiBPr1KlVachevQ3n7/F3Xcw3SLEp+n
lovvQ7DAwId+tiFL2scex0BcugKInDm8jVvD7Up/FN7uoFxxV+rt66l2pWzlBzvRTWmDZh/bLyol
eWhNaFnth6eDA/XwVTWzd6KiKcnEFYljZaFyiSzvRBNGy47u2MOmZuYje2r3gUl/os7vOs20Vr7D
6eIhb6k56OM0DTxL3O7TPiFm9FvCA3aZXZDgFDSMcwRJRfGLor49d1FE2BlBO6Z0xXNtmXtDk2tB
7ZpVRfeK6QVlriIFNCk2R1OS4jEGYCIs/S2SvJYlKnoplQewiTEI8QWmnfwkAQjcskCIZ/bKTPuz
Utj/RoMgnSF3hSZf/nvySlklJ+dQ/SMUmEXxvdV57ozwDYvfKGRrVE/k2TCZ4lmV89D7IVU6pJGY
5E4xcg9nOMSN6dbVi7sscBA12T8orrmpIw2p88rytknaUKGtGL1I0Wz9SYDb24Bu1VcpbJGtuhDj
L31K750Eyqhrr/rRbAGMsytFKn8OWm9Q7txw2rf7WYnnNDQ/h+tM1+p8HH6Udb5H0bethZQj/iQF
uGvZGm4SDSVizuulbu0EhvQxlmhDBEtln6Sn8MfPRAjOtlszouiowbBvw52KiecvWG1VvyJQ4enD
hWshYCk8Jz/dsUW+jnQgNcDZ/WBy+l/DicaPGS9Xmnx6OgmeE3U19r1qZ2lxvg1P3EKrWY3bOEXv
GM7T3gJ51VXGhzArr7NJ50aX4ocV96EqlbcFCuI6ShK0iIDc1+yyGUGv03jCHo01eI+EpAVHQnR3
0IEOI2c1+naFWGR+qEl3eThZ1uvJjnOKfv4IyjtWWC03QVuazQh3OCt/fKEtAfSCqnvLlDeFo+h+
le+gP8mPJGL+SuX0y499C9hZhvLWfTBmbFV4VTb8TyLo3kxQCM4Fig6vgSxpML2GMqIdeykvTRug
zvXbZT/Q1aduxx7fsM4sW2KNQblkKgitHEgIp2vK2Bx81PluX6O9wOqJ8Z0FTmLBIhigreUtMH0H
RccfHlwx7xbwhxdpNjNwW4LmtIJLfpTBatSk0mSNPNGLqBXthf9hk2y826hm4FGWe0awpVjhmsLk
P1fTkhP/tWt4L/R7CKIfM7txhfCY0SWdLcliStAbGPQqdFdRd5MqfYebmEGJ+YqFVI0kauI3Ln+e
nQMa0B3yZnuClpDwr+MTnqINePZjMxbjsduQAU9PNjthCRKkpbpnTAxPlgY3NsjDvZaYSEQFpJAz
KG3Lql4iwjWrPXsgGx8F7gctqWOPfE3tz2uy54wVsqmPvC5tsCRGAvGWnqpQA4mBULsdS1HQSr26
QCEIL6mErk1RYKe06cpcqKA68ms2TkxpQTl5tXY6XynSIVpBqKTIaMHUoVjP+x8EvPCfANysLOT3
S7HPH49QKYn46qpISkByTSjV/suenxNs3S6/3K0Vp21w+cJLHJX3A9i2aYrsQ833bQC2Ice90Asm
1RfmudziZbjYCPdnXutQrQk3dd9nv9KNbzBgu8tahZKLhN/16DrhB6Iqca6a1YefOfY6oUHOiAL8
yM6JejPB3GF5IF1BlkXXRD+/viaK7ibRslgKIWqqpchPeIncKxldjQB5j9mAA0B07M6xAWCnDZZv
RylprLEtSbOSbp46pfvZHqcotIIUG/2If/htnOWN7CCO+QdwOZgjzDF55bK7MWbKb77jsL8MxuJK
ME72+dDGjrEM1xZeBRKCmlx5c1sE95ODyaaHuRTUkNUBVhPtIPgdxLqVHNb7JV0qWSKbQasa32wI
EjkDHb/95fBB1xVVli+QEVYc7x6z4TKUgdWlCn+wb/GqqayWtmfaZoGE8Jn9Fh78aL08U8LPng9V
pzx5983S8IB6AFz3L+dHmMFbZCJOLgmDPz1c/vzu960PWParQzf7oIMuK+RxkAHBXGgvrgmpnjee
a6ZQ0CGkApoMqShQIUueCLUF3rCPofpVhkmDkNkFIjbLeB3SPltQ/ReYxQPJztfZK2ZtuueUOXqP
fZDTkm0zI/FmT5gGQUoNdJRUmWSpPlwQiDUATk5in6aEeuhVtCJFeNmAzERW6hBc1RfAdbyXbFAc
VlBmDy3rXYgHHoyOTtV742VC4y9mS1J5KwR+QTuwlAOMtjJU5jc941bt2YsbK2P3rJFFEFWdaWBR
AE/JwHRynAXWgwRPbhZOZnFpDv3gAat7EeA1W6jMTv+yZuBCUPQaAsmXAwcyAg674azsflK+L/PJ
nK7ZUREcac7ia379o8iBLu+hYYGNInZ/Q9e0uX1mmFF8hn1ojCCDAGNRe/eXU7XmrFurnRrzp37t
f0qL+X4//Lgwr3yuHbTzTK4BhPcKNraQF6q7B9YiUYKu9Ceds44Kh75i3GpYurIxq5arwC/wsR0V
WKj7FqR8qwTN6GXAYVtPN03gOkSG2+HAY0BCKU7khoCWYEkP8nCfWC8+gacVtNHMlJOGZRfZN8Af
3PfF/FVjNLaXn9QENYDMtUtIvCzwBcTuh7kvzFI50qxDp8y5w85DDEE8IL40J2JDxtS50O7RlJBi
i9hTi6dAt8hMlciZBKvfCG9eRLmc+A0q7xRqlwY1/P3bE1ayI8IqyCnXxNKZuk7W12Y0EMRkEHQA
Eju9JU7JkIqdfmdz1I8H4Nz9UEeb1bzYuqtn/Fxr2VxtDywZgUpYWFm1MqJv+1qoJA/Wnd3sn0zq
Ksqoi+roGMGgLYEy9k9FOv6dwdeWGBNFHUVkGtn7YncHEaP4k7XY3FqJ7XtW7XM5yl9lgpAfUd5N
yB6ZtLWJf/ufAE96MGJ/dIrboUiS0E4fUh9J2rdDGA+7B2C0jTagg0yh1c/ncsIoPMtYBG/Uf+QU
qlqThEFaJyEfcI/vdQwcD+Mc3Y30P5kNFYSA++mHpTNk+RdLhV2YSfvb5+H0wSbUcs9NJiFFLPRy
IfLP82Wquiwo0WjOnQ+ijsbMWoNWtj6GvHcE5fgyfb27HLe8rYPAd7bHThl94nFamTpBrl4zTe0g
tQDOMuruUUdKsDSd/avTRdPJU0E1TSXcchdgaz0Ov8rMPjaEAJvHg1cWaT7D/vhufr7RPfoP/q/g
wMXgOP9HUWse/SR180CGplt49ToZ1LHCLcoB1MG0JFcv5Ktht6NKHeB4LrAOfiqQ+laOWfgUAZ8U
Tp6ITbfHGvzNbDPXAiIwX8RcOO/+qPDveWMFOgd9Dwm3e/ubSZ2X6a4VUUGInDAzpkbK/5NuY+Av
lp3ybmEBg51kczZmtELcXatsfX1QhLNL4T7esGoqXEeLI+A8hw/QyHFNNHHQvL1sm9pU3F0t2v6u
azXM4NqDSdMLdpmJ85wD6qNXIsHp1wkzw3hdzMYa6CiG2APfu+OLYhkKeV/5vtB8kRPxnEweG6zt
9Z7jDcSo6TCC64hwVg7NYHZXYGDMH5uclgl2LrtX+B4H+EoW7nFvI7vvcjFbtCDRpU1Bo+3XnpMj
tetwwOBi3c7YSb65iLCcIc6STp061bSQzjmstlIMrv3AR7M8ml+vuWBEtjC9RrhhF6mFoHMhrItU
ztmv8bcIV1SgHipFKw27x5Vyv8pHFm8h4omUoaY1MXImK6+ndT+NLTPL1/LeYakWYkkF8RJX84xq
Ax4sSAXlwYgCMGCp1Jo3xzmBjlf0CPibz4iMKPqDJvZwduuMltMPYtuBwlph8bB9xXQIVrYGsENJ
8rg+nlXc1JnFhsQIxOWBo/khItMarroA20Bu9xaRccxmw2YcoZUFKfU0EIKwp/TibcwSa8NRHldR
o5GHUJ5RArIu40z+teT++X8oZUuwIa1H+qiErzhpCS7+d2YyYowrloAPgCNgIMow1ZE1SV0sEcut
0E8MsRiXgJiBUhbPaaJiZipGm3TMenvmhLsoWpqO4pe5zMN0FHBAyvyhUV7zPSU6aLvP3mwWoWgJ
xfO2sLM12HlER2Pg7VpoYXd3igok/z8UTD53OUqAIqsf3eLkGKDzwVy0jlLESItMnhGo8Q8CZY9G
3FSndQsa37L2GlencVBZ6i9sdFINQ/r9eOQzJBqmfQ04RXOvak2ZVWpN7rI3kFFhSkMa/59LtrqY
N+g69K6VSUILnOpwA2d5c3nmo5TdAGtorwBh48/1JrUaYy67SEIDihwY2SFXpwgW4EDMKm0M0uUs
mivEwxH+mbcwJGoA5NvlnSvknHVPRA5hOKKDXnfZMMoVgZOEo4nFrhHlWZK1okltomak2sJ7dZsm
d7X3MA1GH+gG7NSDn+mhMz3UYDVNuifyqMYsbZiTCGK0M24WesKYBFUTRKlXb7qQY920gT7SihYO
fFxpvEOFbRTjoxL9R+cKcEq+Mh+6/t0zjfUw7Ke2XiNF5Uud6Rpqrbnz3aHospCvA0SfSpjyxgnG
ftNEpCqtU3hEyPdcthNmF7SfwNVBwKlEiuacgdTOSUWs1FCbEKB4bXiOd4BwMqyQVsljwkPod5jU
Bzcsntb8hEgs/KwsQG1sA2WqzNIRVyBfHWRvk4yeiu+p9tF4K76lB34trmGM4jirNVwI7sdPZ7O+
fEyNA2drj60dgUTXymdZunNMA7oTsTwx4QE6fJ17bdVGBeZSFd2/sse20E/y2UYUV5BrxFPaSKj/
9RdomhxXUHkjBIjzR/85pLF24g9yREnVGdC+0sA7efEt7XupCKLtlf0P/J6eFTzx+VIxQBRS39H3
9VfcVhVjbKGzMQU7klOlath/vFKFULZma1duaPXNaG8qZly2DCTCqeug97NVHd/xZf4Ucvah1NbM
pZaS7YxtsAvy82kA4rx6KgqDNiaH83GeAj1QiGjdfSfwS/xMF/7uQlUzjit01BlLQYKD5PRJ4FS9
taLqOabsBeq4ohJDu2X8fgdeObXYZjqsX8D2KQ8rVyD+ccvMmRs8oNWa0uaSIa2j77CsCpkztyZ7
RVOntvZNobU0T1NhpRW3tEQccPFXoYso0M3t1lwhr1HXPc/Eq02qP/bUCkyhVQFCF1yVZca3hwNn
9EPuW9c7O8PNKjZsXNkaq7uFzrQSmVXhhizXsUn/mdrrEpCaAcivm7u2ojeWIUNmj639+Le2bsHj
Iv8Z/yluWN59LGwR3ig7wTv5/DoyYt/Pt4wvktHwvfiWI1dDJexRubLRSA3jItITLOnYzHWX2EeI
ChshYs30xzeooiP0vdBApo064pM5LUx2ANHhKOdSHTR54HAbltd+Y/j7ra8CdMtIMQooiI3UwCtm
LcUAOaeb2wx4iJHyy7DaY6YKzpXIJrYeCHT7CNzGZmiMtwEoMxN+c83xUMuAbKAXZPlfvnRq6e6e
1Zxv3fufsVwqKjsACvS15xFA4cyeDrK4z+invMue7upQeNk7uNMUH7Lp2pYpvoEIwGeJhOj8Ohul
8M5BcqP6NyKN5+6FQmCkbme10Gvfhtey2mth8piZvHlZxh3ANU5wnhdTmbByeqLIF+NKkmqbK2Em
U7eI2qv3DvA30G/ker8v6k7BjnMW6Ejyf7aTZBE2N8o0qK6Dn8uvBgWr8YwWTrPoakITiqkvsnSg
sdRccO8oG3DRLvxINequZ4zQ26HAjVA9huYefYiGA6cOPciejTNlTe2SGK0quUNhb5wZU9tkpKDB
xzhDoY68GGfVG/9LEB4jx9ryDqSsnnd0leo1MDVxf0LeRqAMfrIyUJIyOztvBROaw2WLBZVhxEe5
rGpxLA/kl0hio4yh3HkGFMx7ZknAYr1co1gbHgRyn4OBj9znQKc/KS27TDMKZsemYxPU8rQuY2b+
gSSiALIkmAqDab9p4d5QnD8foW/QBM1B1zUqS4HgU6aWa9lPYNkfQrRJv1ce7ojSdW+Cuj+YsS0j
kJfahkrAD6PxqBfmSCRodAo7wOX9+bfsw221XPeKw/PEEL12JF7WKIfc2xv822FIHdC/zEy8Xg++
OGahMzK402+GXLJt/+zq3Kd/nUtXsrTgjaqNC0hu+GdzltoQv3HuwMNEakdAPFJ/RMcUK4Y8Z2ta
pP6gCH/1rQA3nGG+k0PTZWIjqK9qqSRp5uYijMUxZ9YW+Yqz040mfDhzyeyM0tuW9JdNfW3JKzyD
qP/cD7jMUpZ4PC5kDqDSNgVRB8lM5xoHiKz4y+20xZRUjP5hLYK5SFEgyKuo5ehS+0HZ45WMliD3
AhXokNdPXNzerHAwmfFYL26j2Qh5i0k4GCwmy/0A5RVLITrSBr0wKZmaagxgY6PbKHnjzftCj+hi
sQviL+PBJ3TeaChpVnwYJM2rY3XgFyMwhWW8qqnssial2oRSPV5l6kJyvGHiQ8aVrfOz9RWworgR
EYD2nEEaN46T6J+6P7lqzoojM4lokPlyQCJBMv6UTISMaZle4df6IgkDgDPRoa0lSo78Ai/Udw4s
X8I89bkUJfWuOCP2Ire66d+zTmdK1+rzyEZA1JucIanH5DFEMQdL2UY5bqXUNj7Y1gT3Jy3AkJHd
ZqkHoOOfbh9911QPAjvmUN+modlpVNrGpsD//qwwXnCuIpZiwAChr+4MenYpryUo6SOciqfFQHN4
vRa43lUf31IJHHNCMYV6yY+RKl9PbkSqE9aoYdadC1R8y+jIaiYIa89g2zKbyGC+aYL22OV01SEc
6A3ICblpadaNPHhw59sc7RBPcgfTfmCrNy8tRjar7GfH1un3VTFj0OP4+4zPMitvgXvXT/PkYLKl
vC6pTOfsQOnuAl/U1hMymyt2plyyjpnD4kg2YWoTsMz7IFxdFPsgASgubcTlgznm/x9pP2QBT4P7
bGFLz3SUfUuaekESVYXWonMVqcEmAPXJov7ECf4wy3Y6TQRKr+fB8jquoVO7l3ALswmOQKi7jjiF
/U/xBLzJdtDSXGIgzJMB0Sua/9h6nCVpCnqpcZIiEVAJlQ2416tTrv8ewx7BMKMBqLL9pT8xgynw
7GSOyHTa+MelvF/V2WZXwsWxWwvQqm0n14JZg7oVxwXHcwRufQOTQq4wIhaWPfc3QEoAJ+H5zGkR
nsiy6RPRV6KCn/aVxx7ejJ2wdZ45fuN82g2dOTocoL7MPlLbSDi+cHXiN4WcTcF6AtFo+GQVNYmD
PzAsifSrNsH8ZKuMbkXYt/XqqXDgnMTwlvPB4MphspK1/GQhsLVPGyBqCYz5qR0h1thFs8NYG7bN
ysoyQaqSUAntE21Rg9L4WQxky9htuL60FLrY69FZUhNOKW5cXsR2aaUC21W5o941HH6pZAWV1vlM
XE2fNn19ykLMTf/Nn8Q1RrSJEHBlitrQ0fyVDGXH/m1nHEPzkciwE+EOJi+1KhFlkaspzMjQoKJV
0HD+pZtEzfmqCLdgTRrQwwGlHOlgD/K9JG+Ej7kV9P/Z/BHrHMGe+zPsxHLCeKwgFx7o/Cma/WTE
AHUxEl4zlAN/rXykZBBz0kC9gz1OawN+O3+rOahXlzAKso4frhiPYE1lsYdjB7boK6wDnqk6OOhe
I2PHPN1JTYf+RNjw+ilJ9/Pih30H7pOjklb3LOK6WMMuzugy1a0ZGi+qwKkClzSF7fljM1a9Vpnk
bRnxLyA66jyCW6yjcbHTtQCQ5TXT0l0QXATUYx+dJiBgjBbdzKyYHzJnlDgn6cPkODcfLVH7Im2g
DNgLovMHH1OmeHVsmAQTffGmgKqU7QBm716e8BuZoKpiHaTF6Ma+pd7OPV1CYf/zFtjRzfR0k4xh
1e3VhnFKoH4RETyMMBqGejKu/iorlhg6aL1+bQtnakOaye9+iUP/ZdDjzMH4pfx0HRdzDirle06q
nZOG96Wb9qhnX1okluBwGmFTk0LYvUpPt6LVGFzuCeBYcBgSwOkIlZ127BiC2/2bEe5GbT28QLDe
/BDrtarASHVvfdgeulXMlNCqMrD5yM3/TvGbIbbUK7ftKzszdHhHMK1q2hXTeAZioYaLYwkUEelk
ixGMKIy+BQBC8Aua1ktyQ7CjTPbdws2bqG0JPkFeDd1HnqjpCOPTwqP4/Fl5BaD6laxk9dxazG6X
0lPibBho2L8y1sNK5iJ7VABgHWT64NuCuTdKSfJwR1J2QJPhVHNWZIaWLqxaIP2C7HyDj1Nx4bS+
rHJz5VDlwTo62qe7U8K8eevPlwSBsUd0soqd2jnG1BoDIuxQMwUTKHM7V0QeBksqEThXEP0QooMA
p0flRJSyAwWpDEWwXGxV9/QGbd9jmltNIlTzJhPvQJoD01Mkop3VA1an/9KFUHW3/+H8K3sDDg3M
hY9RwMYQSK6MezupuG5z9o+lXtL/HEQyIeh/LkMJmqM6+RvK7b6ypfV8kHwIB25Eq9hqyusva/Kl
4Ce8FvteZUTbN61Khi9t2Jc4KYAD9+Qfa7hoqyZh4x+/T7lKBhC+qottZHMCODKCnLeJGShmN28O
U9qZkZDzJXVewYHIhWfLwulQfmLIzhNA38cA/z7wUamEnaieXuv6OHA1RbsJd9w9BcQ8EhvFui9d
lEuAIqaYqjs67Q5FOp8BM0oO5+nkOdEOeJMpVynjtv7ZCgiMV21fb6stKIOvmzG8j+IfNxUAa6N5
4UoWZyqQzH+9LObp90H17lne44rnSqggn0tH27YvVI+ko09sD4nMLf2VAo5cODzj5kwpghgquolr
xBVw3wYohbvtycBRgCVusBgmVOabuSEagC2L4BC0ZD/69rc4SLPrJg15Y8X24KwosFB/I07cLvhB
inVrNC38LMl2i/+4gN1FkgH6eCR3Rjqa4mbU7tOYlYEhTa19VHRdmzXltaRmZaH80XanUafsgg9g
A1+CP5eCScKfbxumPYfz1AHrck5azUKSJdTvRK3KSXw2Agszk4De5cPolLZBn8VLv0lyO6XhyRBS
S+M4sKqRr6EfVh7Yj+wGGdgIYh48/VJTj1VzjwJrpqCcA27ExlSzgUwR1c+mi9VGVWZmtExga361
GkdLxNB9PR9VlM9UUHLZrVP1b/Kc6WzkKFdSPXK7mpHFY1NFcOZJPYywErHqq/8HzpEx9t8ANvYA
YpyRDoXfJw76u++d/Rdp02mFd5eIBqE1cmzhW8aP9hTX1GaIRK3gt2Pq3UwASddpJ0+Ey2mHItXN
Btu7+sCETt7e0xWdY3wQ3B6cmIOX34Y0CvZa6AmOVessz8eh7b0s5L5Cwd1DNyxNJPr/Xy8OePdY
/qFpEZa2PS2VHAXn4Ql8WNXK5VnXCFhGdP1xEHJ1rTuSQadfeIxMOoMm8PrpGpsnpIR3SD6Cwcps
joiksVQSP9jz6mtyrOneA+dUgaZPvGNLLdqmTy13e78xeHGm6bz2RjCuxHCpqzqFrELmbWAaD4X/
kOqgcFaaI7h/TA0IrjmvE7zGjlfYVai6Mg67tvvQ2Geb0NZ4zAMF0/2n8QxPnG7b52u82HuDLQL7
5bx2eIFcqEKsFE1oMbRBmk2sOhf+tAH+/ACkJ6TK0nYJwioWfOXKtCstaK7b/xzCxt10jAoSN2nE
Qk3EaOb2Dv3rhEEW7Rz7zuidXaCFFKT3nmOQY8Pgs+owe4IR/yWDZ/r3KEn2KrPNEzSvjAErXmEn
nh9AmhqJFIWCC9NopGFkXVU5NVdHMmvXzi6Em1qI6unXdnR9KVqs9NV7nRD3OxUDw4mXkvByUIYi
zSMcAGjDIyMI4wVXkoZzhan2COPk138rvRKVty3h81N1wktqyr0Hbj1TzHL3DeAoxKWd5iB5N8uy
zWibLhyoMFsTcXiq+54agUki+f6/XjklOR0yYdWqQqBw03CuKFjgwdQAOkvGUkoGYnmwOo7AtdY8
j6z+6parknOQwGHWQVrZbI34jNHBW27cy46qPeIk/1jdhgPpQsD1tiNPTwjwN9cEqQLjXmAbkfuk
NkwrG/NLQjdafO1UiwdSObEtPZLxqOBe5bJU8+kudQ/omRy+o8lrkeYaiIJIpfX7Xx+xgNqLBJ6u
Xr8qV4LCQa83TX+oaN+frQ2TZPdjvgy2eLwRZ5hvCBz4smtHCzVvZBT62WUopOSzVEl8sITGCTru
II1tdFYNqKe0fnX2qQvlBAfQAPOEw4Oan7KsTpgBwFWS0bVQrG0RZgmWQKSwgaRPoJah2lwAWrVM
6uV0A1RH5WdYbf8usjoz0aI2W3pJqp+mk04GXWWcXmN1nsS1oh+lfBPj5Nkhrl5RgIkCnMDqMvL1
Dnd+v/rnUxNrT8UhtIC/gYnArtGc567ArPKePhDbBCUnkmJd5Dkw7sZFtADeC6frYae40PW1xaFh
+3vYGuA+y0VurcNIb4AetfMCnYPtxLQVmoYu2cOnR95rz/9zpuCEQc1z+086WnjZATaVW74XFfUr
vwh4zq4oG1uM3+hE5WdB7g6sMj/TeCbA6gz3cL4n7/JJlAOuhzarNHaIDCCBDq5obCUSYaM/d62k
MMS9qgIXyJRvXSYdefBS/PhCqdHtd5tjK0GS3YrQUuM3TK9eayy5JfF66J5hactg1O4+A7sVoA/F
WIzw/JC176lrSddHGKYibFJEWsXgQjAlTXEdTLHakg5mA2IvjjvNY9Ze7NuX7z7h5RhmnAFzDlPr
wpfUcvkRImDVHYBMhiloHktYHqONpxTLlaoGMPMk9KlqCzSvwOCxnMBA711XNs+X+RQc+nwVv8pw
wRtp2bj4afwI/ik6XzhxL5Eiq/JiQPMbLvFn40F2yKHbY9euQaaU83bNTTfK9WIT9yfkGyUTgBnt
JgmZbvP7QODCr2utZnvjreh1Fvz+tae4XAUKNDI4nVodKMzHiEJAl6gM5zlyYugZ4s4jCSviKEeV
ZADnK2hgq2eoqaGrwt5UQOfBC2eOjKMR1hcOemH2jLkTmjFJdcGvtTQhdP06nmPs7tO5KJtvRVuy
VH+fM8GnL0tSOQ09SwWm0WlhyWoC/tWbm1Yxqw2p1i7lIwjjqwEXtlRLX3+rLRNDofLVdvftlWva
hVJU61qQ8HW4w+cq1jaHwhZhEjWfqRItFjzQ8q+DuwA0QsPEjf+vgGiqIsCfeIHRF3E/OLGSB4bx
ml9qIaj1OXou6b9M1siwkJnr9SKPxT527dKJ8Pz+6Pq2yz4QPY8zBuK8dOELejb/ZAWut/YFAvtd
I2SRzfWURh4qDCkN4k5WrbkthzLuUBL5CjAfpIEoNMBkyoEsMy5DQF6oVM+37LDmvfKiUzfx+NlV
VGuirVa5D47ZTragmWlI9jfuYWbn3lmYjNrzicJgSCvh1tKxfVTcAgeKihuhW2Gr07Jno8FadJbF
Xz98v/ryO4z5wU6a4L2vmM2gMA8CT4Z61W44HfCtVdKks+M3JhdwbYbGD2g/AeUzi5COPbIGRkvL
/uDoCqbXu8dR5SlNPfNFVjtved6FZyNZJfLFFQ+K5vjoBoAJ+A4/hKQBiIRv2MWQFY9Nv4x4l69S
FxlXwnaMQQ15zbAOFTCNGp3mEH5P41Kyp4M8DIpEavs958klX0b9Yd2z1AYZETmEVMa0L/AEaelo
o/kni6/fXimp93h3gyD47d3zww6Ir6R9dG0YE3nd7lT+I2Q2ZRKrCHjnBqTfrC2j2LB54o3z3x7G
L2wq6NbkJFR8U36fDKwUWjwoRylKdzkQOqJgShhaxdRjQSI/230vvmfZcCHuxQZmSpdrRb7yf+aE
HVxS6gy0Z12c49aKSINx5LkTpaH/sh9pWBeSNT8Nj1NAEjJxaE1b2ZJFNbIPmTE/cy0Fu7Tc/Cj4
GsxPBTiuONJ9KJb9jv7G/to6j1niaoa31ZJMaX7+Xpi29GDGCMQAJotQFFFTDxZx7hobUTmLDqmC
e13JRLikM6tkGLROp4nvQ7EZXTzHz4+frDgSucQK6EDDM2fkiTDpBN5gU7ksprK1mrJqszQCRLcw
AL2iM1JryIvhiwE0EbGBZLYK16AMFuAILzemiRicZkoD77zP3Ulky2rsNg+Faf8eyAocw3oYDqxR
sisWi/jAYaIaTst5+bwu26+7huxz4vgKI1G67YA4FWtfSchfbdvYf1IVpoAAPa9G9mOLgKxwFPQ2
3zCFc8uq59Kw9vt25Vi7CvbNBwBJ5TFi8EiyamqauYUUr0ymMqeR0yPy3wZTdQl/p8Rd25JEmVzP
MbgGWqp5nJOAZWtznnyuPRnpPGf8gLJU6w9ZSCVyvx6oJlrrX3F+bMJ9Zw+c0F35XG6OKbZeV715
EiWgpEJqiUbtPN8PqMejii0jWLrQHOZGTQazdL+ZXVcyWsV+3wADcL5kmanFmpPyQ2Ty5zirJPes
0U9ne23i9cgJj1kRqgZ5Kg81oTN9sAJqHnoSapHfoF4aQcjLussK19jsbQ6j8PLwidW6kImEG9X/
WDiWiMKUo6zmvphtVveKNEpjapiozQXkTPE43shuThw245QPh0Vr9+x+Zj8LtqsPiz+iCh+epX04
oRMRaDzX6l8pSDkYBONdyl/wpq6fS+q7MWIl00CxIjF462wANkd4pMLMtYnSua4UMvHBqrO5vyHL
8ARSgoHCGRmtNkYheoNqNHyRosJNBNZ4dCSrDyoXZDxIX3S/Ems03fARA9fmaZqmS0eiXU078bHb
O5ArNZO+qz/HQUWyg4OWnYz+kClD4JBENcNqQcy6QEE2YSmvK7gShj+9LULRGPNUEbcyBvxWegB7
UP4XNhbsLFZkKfRLUssVJIvkx/Ye6wD7vVpIcMhRiIdpbuKqNFYSXAuA7frRG5+PiejHCA59InoA
UW8OdmunbUUaVO2894kGlQZ+YXhlUgRqMsoCO3M+iCnV+pZt6NJX7oDfzHGn0xi6kx+a9pTrlm/l
h2YLxYClrb/OV2fKz2/mC10FAV6GSpGnV+D4XzexuiDNPrhc8JFZOLsa9z16qWJr6d++BC6wLxfP
FrjNx8ih953qkvlAky4eKOIo8nzClySIMkMse+ohTPgNyJW8K9dk5g8F+FKJoVe2w60ywbVXgLF3
Ldc2dU/nKAIfAGUEVaRuxwcwwT//6b2WRpUEAnz62V9aS5x7lHTYdxFyswLE479BEaou+zrSjszi
dIsXXOdQ1s6O6nR3IIoE2ZdkbP0C1MRbKGIhlVzSu6ZXcG4G0SulRgFVMa4gnNbxPSZGQMSIPR+P
JAl+bqeKONwMIFgSQyGuRD8xVEYF1oBC8xtW0P3jaKCsIt0QeKYxuQ20SjtCs6NsFtZAjrqtRGvA
lCZFPztocUWj52n//POr7wPKXMMrGEn8bwjh++H+r006JA6Js8bDMmNR1ELUDWbu1HBc+TUt571v
VQ++d/v+7isAa9qwgmRn582oamWVViUX6IYy4cgNZ5F1O1VSTOYKNRFL4l070BcuXrG46zQv5wt1
BBD0nsxQPK4r95Yu4XGjcdD3URfL8H0O5cxHKlYvVUN8biG9urcnpilWpSKgq97M38aGUQWiAPau
/XTKK7AJuSVLzq7mDbrv0pTfgvf0QaYgfI7cuFw24g4sef7rbGW9Uw99nuYAgmKtKrAGwgoDVrTv
Gmdql880lOC9S/pRa9qSUWOSfeJAk/88ZLwzkK4Y4NF0mYEjmTBbor9cGGGkXHI1XyWbEJc2pTRX
1cfmJXn4+t6TkQd6kmlVZuskoaziP+8yb4S17q/KmKe6LhSLMIK62HoHuZhWwd8MPdFjUZQUbdKB
xzPzOz22i23R/3LJQSGbkNQfCK1WIUm/xk4G1dphJadOyDmK/GxeuYwXmA+ve5y6SdhYgbJ5uBxQ
lccHS4sqF3AmcBRuL7J012JBK3ou96BDBdcE21ExNnGNpVuz1ZUAx6DYOPe6k9jhKEpFZyfucpI+
4ljorKia/ZwMrzt3thNV5b8tKa2DtV+ZzQnMgSUd3h3pf21PWgFujB+b2IdihgqpH8RrOkTJrBsT
b3Pvcbhs2UO4GfnBt4416AoY9b6PchuBr6teFSdGAZE7dwV76oELuHlZPmLW+ighNDS6OclU2jVM
2rLNuUdxw8HfWF+wl19xFKj/CaUjrr2a0h1FZ2UlafOLRfxuTSao9pvJ0mAUqnJpWmje2Zi5gp85
O5vmOo2FqnR/GCD56ftU2jDP4h1zy6oj0J5+dBcGGoeaVFnUSWU8rFX6fAHZQcsUOJt+Yx9nMvZ9
cYXFOB2MCJ3SGaelZpTIfLRcOpJa3oecAVQVYBNQ/YGLdlG+6PWcsy4KwwcuJAWP52jJNsOYIPN/
9BvFe+5P33gBwfE2SaPZlQ7qKnjFq6Qf5DRmrfb0brWCB7Jf2Wl5Ht6A33s6wu9YaBK0glWH9BYV
1IiBFVwQsRRXTzzn4l1QG+vSuojWfTiP5zHry0dDAftgn//FzVOfTFqxdGflN9BkaOTn0CqnYwCE
G5d7HEOHxEs38gTReaGfSOwR8xKhOzUQusY7FrXOGkVl1K99PT9QxAvmNT1HYQ/bIRoTqiXAODb+
qSTSRqK8iwKt4DEYiH6DeaKz41YdPsUcV5PHfkaV3jfBK2o0bivtoWhgFfNC8B8K4DyJzLlb05tC
j6J18HE6BhlCxlyGHTMW3lUbumFJJjKTukwIzQia2WiPX1d1/pwr9y+RwmI4jFoyJKkl/UnEvRiY
EL6oYgPvk+tNfG7+3kOWMGps+9IhpXcZXw47LFJhmwqnsUL6XoPsKjosSCGHYpKP2sP3al4SdMMg
W8imKPqPJEzE7CFyG8bVEjEeBD3CmDIHfAidYowvf03HAtzpgffsTtV0cf3K3hRlec/Ts5xIagHj
lm0bzG2T8K8nOOWfFVQXOmDSfnc7SXxTneEWgir3stU/Iuw9Lf62agE1uy5Yl+ttO7D830By2Rsc
EHrWbJOCzLuiCgg+3VPQO/mfX7fN8OqdCIUWguxGC6RSz/WkXTWaDUUByNi6YiP4+98eyYaZdjSc
HmQEEMU3BAy0Xi9dFz7K0SFKMNTiKFzaC2B6foAKLpnpp8U24ziN8WmULVPMdEb6PnOizTwSg7l1
rL41RDiY17EqdDmQM2u4N5NpBoiNjeGrT+zRjgBBRosgtaysRhe/B8oSUG+54zcsooAblMAd3mFo
NrUrWIwhx23nhJDc1n+ek/goBbvzZqKqAWnh1UJIWs3HVkKONQghpCfzE6u/pftZwqowxQIeqUrt
T3GyYJTodU368J1sSGGAAjYDMuF7CCvBaCK+GJxPrbITCd5v2vh4+nLL98ogjKZ4h9+IZaWEeafI
jdYwdCP52EicjwewpH7jw7A7y3hXQZOdn9cxZSPuAIV7xRI2DtRq5JIHr1F/tcv8wtGYvIxT3EgP
CFY11NvNMFtiVBo3S0h35Jg1tol2EoITsH/maUyTTzgNT0+irzd0iPJxKIy0M4ao/sB9OgUbdP3I
pUp+/FzXKHTGqji/c001BEr/CHT7XXu0cmrYE+6hNmHS5RNaMFbmH6EdYKp/f9JDLFssu1aTIsE5
0xVKGb6L1KrlniH9CcY0qpTeDn4ItWrEvUsPIJ6NFxkxDAZIu8hLF1sCiw/bZ3TMUaDt63pzQQ2m
QcJ2Cj93WbBSCgLhnNhoM5NzDxhXbn2NOxgPj8MTKBR6RyORLIJ3kcicohvxnNMpqyBsje03HarT
JCNalHHoozeXJRhqvxe0FwrG+tXe/7loMS9DVHXQ2LTW6P0AYFjcqAyR2MuXGg2bq14M/53ZfX8n
9Xi9jigW+Rry+a5LksX/D2FcOL+mXm9Fjn3Q0QiNvD0oIlAaykQfTjuzm9Xj133C9MU6v9nivjKS
DMFnMHtNiF9Wl9Bt8GBWpwBzRBQr+vCMlf1QMSduAO9GhAiJk/jp8TezNh652nRQL/h5PZUk4wGN
PvjY+KYshTHGL7gMbkuf0GgYBiAGPvqRcJnaN6+hxp8XZmfo5tGsbtWuodEtiE4y5/lYfgwNKXUg
XE10b5PEeieJUV9piD3fjKwTO6a3BulqfrDZDx6JXawPBdvJ579YzO/SnmYBC2E2JtQb23G0eiB8
5p+dvUAseb3gvB4962HdmLDEssf7iCktO8fqAcupbElmBH5lD9ApCVbtlUrCwi7IGUCbduizt7lG
zws3CJr03m8jv0fIf6gjNNzjq466wPMKQOcRHs1XajDG6SYYa3ujqNUAigT4wt1U4sqQ/a14khWB
+Jm1iyfLfjTtOBtfYDfMFHPDolpF6AlJEKhksgsz0R1goTrrKTf3kUN0cV9mG9Vc0zVuI/JgaF1b
721hpdgf/UzHh+EsgqsSRQMLriqkLV/zEDEHJuaWu9dy3ZsBrcAMtzb53InJYbtIdjqcGhNmqw8W
eI8F6+4rC2ZEgEdnXMXk9dTir2vhdZufRxPGKaSBdxRAVoCEQK0fUjHj6rfC+tXmTNddyekBopKl
6nYUF9yBetutpNWZq7VKkpoJQgV8prJ3ITnKabhs9TMpdbj5vjSz5fYRue0rBIz5X3CGtszV+GcU
v7dUhhBDJo6XbqAiTVscdfx6Udk6u1L7sB7UGtFnJWhLY85WqhuKFdqX/ScBrAq+mhaJDOQUOXLC
abz7os4tBG4HbnrORJu+wfBr65bsevLD+GqnuPQ7d3UtvR0Cc0F0OhMCYIYQiS+MLvssboLIrPi6
Jk8AhsdAqztHAH/xcqVkNFXq2fq2Y6SZb6ccKrqSVFewRcFKHodi5E6T6uyxaVXHHIlJuU5TqDmi
rbozl/ZWFxp3vl5I4qpEGPF1NirnCUElp7HGLhfIE0j8wn4AuNer/81LzmKAmwlCu6H03oFgPox3
fFo0Tkqn4PQ1pytMQdSglJ0XOeEcFr4MzwduTUZkPesz1oYk3J9AJRtyWA+H18x5tlYHGcxZ5W0M
I8DrGgRd9oFbGu8B4Qg1Yv7FVRLrKf5kuCaTN05SXn8hyp0+1YzzO+yneBQwrwLtbRwj78k0PZSd
NN3A9M0nvux2bLzkE+jzczuQ8aZjR94VvJ98JCjDGH7Fn7rrdWo94UCeO7ILoE7eV38Obxst/FZj
RjP5NNypFugU8vo/r12VYCm44mCl9XqRNQLfQWdRGnoXLp30JhAtUfLg4lbKqkULsJO60HXUq8jP
vyA7riMpwuym4x8ia+Q/YxE8pf55BFkWUaT67zyH1wOgxiP5xnaXQIhCJpYe1bh63CbLGesBgxaW
ejwxb/OmLnk8Ji8i5XaJjuNdW3rbwESRwOmWmbtK0nDnhvz2ZFZCFMkPeqrXAMci8XVRaaUtEUaX
WFCGrM72AJfduuU6a0vpLc6cZ7mO2Rfd42PENDnwgZ5n7CSo95YuQoSEizDwnUen/pjzPwUnB+l7
vTfcYoZ+6o1pl/gubT83zEx+n4HOMlnMP4PKKuonsHLwI1S4xEKWThc4OEkoOses8CiPD41pph4d
R1hK6XXFEdh6ZrM8j3L+TYYqMHEujkM4AUW3hMYsOPSJfJ3KcXP4+OVFdyEyKX8CCQNaxDGIuMaw
F5g/hrNVmACaFIjLY4+Vzj9IrA66Gc0/mVwlfnMNI90aECAT/frx1D8f1MxCKtB8CL4lAd3pzWju
OFTZaDcylzxHRWWbdC8GYbV+wBGLSpKGR51P66T6z4eDlHQ2m0gfnU7zRmwkwZzLhIBl3vUDn5OJ
eYsweR0BsU9fxO755BcY1RxWQurpvHdfkxmlO66/cE1J9oem06ZXWYJKszUrWaV+ww3aOhXTpt7K
bNAInmH2+X2M23duHH3UZe0EthodVKk8A3blR/AxtqfpN9eQNc3ZcUU87Mg42rkd5NwVyXt9GroO
wvkjnxsOYxfZVGjSl7YVvz5hUn/M4q4AtAsYZbXaeWpDmulRQBACFRP6+d22WEIdONRT3Vs6PQaj
I9F2Fo3P7EQCQfH8yPPNhxHHzmLZRcEEcgD3rQgdYuj/20BtpQH9luI/4MQskkRAxTEF0dsZ9wgn
FRAPs8080zc7aJM5zd479+xwCuyXuy7espxpqD3vrxvdPletJqGXJubBXk8tGvdH8kRssTojKjb1
n8g0IzWZ4h0pbjsZKpygWFgs7d75iTkCrt+PZuKU6CFl6JzDzc2EyVyK2n8rA45Jfhi5XrUmZqj5
3tdR1qlBMTEdiHWMUqL2Gj2uJCicvhglHHPm7REbxZ7KG/syJPYUC8SbFFQtCLv4EdBD2zYrhRA2
dG4NfijKfdfICRqpQ09SVTVnK5lP0cWgFvid33rAzOre6tUtIoOzmkMc0oAI+yvQeh3NmBzS8oP5
KsDTKBjqrFF2e7k4DLZ+gcz6eh3Ze+wQrCCSYEuRfNCxFLqsdJmvvidVoCc6uubfIJkqkewnOp2L
zpKc2L3D6bwz45Zm32Ql9LbhyWSk2GQJ2Gf/CvyvIc3ZCCRYVawyiDnwhaUgUpRWPwvdREbaKgt4
fvKcRevYG2Ud/JVxxLzmf4sNo0GXjlsBp27mMIPjV02YQft2FbJK/LfpTo6DrGXBfF0+okZm0uIJ
uUQHIPNMs4WINnkHxwPeYupts+XWOlEFmOv8NF/MC2BsfxJH+nrp819orAJ8OOPT/jvtELVEevNI
vdTk+6Cvw3cCOcSZxfnPtNQ1v95X6qGdyV4I4I9VKBwIaKcn20zZT2iPtxuaQE9Jzn3gJ0zvrk23
5wVvvcYDfTs28ouK3qV/Xgp80xbZG/nT4fRLv24F3q6RPYV30jLJaiCJhFN81uP4w+0nB7pA6yDr
sjriHTOfhga30DH9mI1MibxmK7+HWRe3Hi376HMysEAzG7YwD6c7VaSBsDByMzx6/GJWv0vp2qRq
Qm3NddPk8IQHxXmweMtfCHoO7X9l0aeE+YhNG8zGpR7PGa1ScuF3J8jJbwezQe6SN7K32i9vqlAn
Vn2s5ISR42VAU3BkDxXUhtrT1VbnuWuPAXSqdw9tSKNaycnSRXoo9C+IVsPQw2iUbLqABTDZ0Mwj
dCOsnU6vW8fug3xDmSgWR/otrAliriUNAt1teQ0SMmEZ/ei7FwK7HCbv6k0kr2YBeIXz1mO+D40r
cJ7z1RYTOKDRrrynvUG56ZuuwONANbuPGnQCV8FzR4lrIl52PajHE8h0uTDMUfGDdp+6osohVjU5
gc+O1YqH5/ZD7Qy5Z96g/yOddSTTVluVXE/FNGv+bQOaxCLehrGFVQpEjkc0b16V9I2F2Rs3GP//
RXwmecJy0l9oyD+D3B5+ulsYXryaSj0QxgEJRfEmXW5s6YspuK5c77oNCZvMKZPmQi3PgnZTrvla
uUkW7r+8r1s2I+XsjSUPab5SrspmaVVAczjR02dZY/KNm5+cGgXE60QtoI6iLYijyAAaER725jYh
gTG1feahSC9Uo3Os2rEm76kHCSfr+eutvQxLc4+po/6qCWqS/AlYVnJtx4hNf3iTaoE2RI/439PX
Yt9J4bBKWxkLiyfu+DfW7MkLyxoGEMwRWzBAzN62MYwuhbGug3S1ue55zHJGsqQ8cN6pCf6w9O99
defkxlVrK5KE604yh+tZ7LfBIqeLNund0r9FD1B7xI1tvdS4cUKrOb3xFny39eFcbytr6qjyuomY
tNDe79rUUUixlBhYeluO9LBQVhI3ExYbyRqiSF1rtcuJcSUC2QZuZz7yDdnoeXXvpetzVLeT+jAW
14xTeIsFlbN3IPSOKlVHNpdLEOY/8lbtujAXpkXqHMNcDM974bwcQV8dW8Nv8D2FWgtVjBywdYuN
i1U0da1MUEyAKEIC3y15Rrzn4fqjlW9CduOWSoBTBHycMQPDYtS+ArJ7bUD9HIneQfDnMdgqOxPq
jI5phLe1vyHQAwWp9boyTC8QMe6CSLKnHmLvskoUr6Zg4pWe1ORufYs4zSsxcvs687McD2wlwiVD
HqvhbBi9ZF3Q9VXTtgF2hp5eqcm+g52ipmlP45xaEB2d89MSkcRuh+HiVVMRHXGDWeZtm+lxjNme
d6sEIPUqdZGosz5YUZ23MXcH4Z5MLRVMb3Jgt48WEwVIB9gZUWAMHi8LYHqBdhoT+7sxSIDIxVtA
l+RwUiBb86weifiRl6EH5rMRVZ9YSpVk0nFFbU0p9CpdAnBfFiZiH/Z32lqnwqUCHqaAfzB2kq2r
zkxDR8J55ZuEcaFW7MRwsdYWgSkTzk67KzeN4wE36S/L7fqJJqcCF1zKgCMymXy74JeE2yuXA/Vk
LzQEqmC/rLAG9h+so4UGUBl6wflKsKxUFicALHPtK9hK1Vn8kFHnUET71/ULbciXGAF7E+DWlbQE
zUn9bOHwRgH5szdOIqnkw1ldp8hj/b/RxrX9pvzYgEIsCAHswMD8dXTw0YNaqBxRJ2aPcT35fX0f
tBeEh+45G7VR6Cj9usPBVrjl/TOPi+UETCEkaw6P1ObB0e3+R7U0VG2OeBb2gJNbdscvtjPw/sHG
UdWflcEzV/SBO5T9mr3U0gZUO3K/DKc6QcmcmJs7R5rv2LOjheMTvv/mELghGyzWFIhfcGhEFrHe
euMlpCS7jungw+dBlrADOPEdSV3tzonAzL64e2n4J+C2LApt3SqYcbELd407FkrwlNMQf2vo0oLe
Zux3mERSqZuY1V+MUjgt/oPLp1JaMrzqCcyOYj5IiRA0q4ncGAUVHeUqC6aAE+CFwhNKy4scviIU
b7AkfN00jZcq2TKWXRzNrpJAOlNsjvWVADTocvoD0NxVxSSxXMSJxw+mCHWN8jUPMkiO9VyjMEMO
qw/hBMBV7noCfea7R93K38zxGcbmRrsuzf+mTleurspHOqmzufL3rZzRL+oRacIQoOBZ7H/oiDHI
lbViQ86upu7JyuibkU6D5R1VMkl/LeduqQDLR4lrkL+FjS/pFaa3LdGaBJP1SLKs+11ZUJU77d2T
nawfl8AqUIZC9GS9Cfp96iC/jAqBpXl78ylVcEoYxJ8W3a2QPWysS3AQiEfpy5BBUYy0u9v6T0Ik
Lbc46oSGiRxVu02pHOC5zAB8T+IFOjs36bME8jlL2LCtA/KfU3UDHR5n4kKxAOSETMuhPZWq+E+9
8J6b++jqB2EosJKUQjLQb8nE/DSJJqp7Smo5wLy0Gk0+lQS4n399E2fJ3ny8Bcb5ed0aR/w8prAm
7m2koZBO04YrJ4Zh3lqZRFpB1sutKWqY5FHIZsX+Zq4TsUKj0Tl719UOejuVS2zagh4roquBTLhr
taF8WlwhVE81/sCZOkbaGK0//ufiYDPQ1Lpx0AjrBX1890hNureC2zhSw7+tZECIpf+BekD+GVHa
fS0J5gTPShI0Ns2zxTrX6NmifKlIsuA3hqdc8RE7FsQ71zXjOTh1eDyRQJgoi5c633sOg2iaD1wE
HSDP5lduAbdhETqJgBO4KQB6EutfBUcUcF9mI1jcH6vP9YyvT+xpwgU0Ldr76z2MeLh1Eht/uatC
upQLH/NZMtwbcTgl2nvFSbjlOXWp/BrPnJTiAMKaqJXhuZAG/+sPswddeQ0uH7Lddc9qd4nvV5PV
22Bgb3TOX0dSBrl6O2sTjDMxpQoJpgO1MLU+DrVjmOhhvKaoqWX03ITuHnweF2UR1CNJCwCRoyD8
0aC+juR2mE1uR5BGUOWO7+4Mb3FTohRyNnBIP00x69cD4OPThJleftjLJcpXs9sGJBlb7Fky6U9t
elDeGiT9SeX3ZgBocBlkWgcoJ3pZRZPfNMm16FQ7OHsxnra1svEZLyqwPFm5X6AdQ/y3sPvXg/2M
gAaHosOVCR9F/47StJK7yCC3zGLx29W7WHvU3Iad5aWKHaBMnI0vIdCFKmfRSbognj8XgO08yHgn
rPG1XvAgEtBzHNM7tHiDEm7P9QBVTzvoHxg6YTilWAV6D1Ka+0D9k5SCZjd0plPvHhxlKlt9gvKn
E5/O+DrVJJaD7kJzmVoFwP11aUF0xbrD+0Lmt8ocJVnREzSeoSiIiXbCbcZY+HORvjw741cQQFdC
AojPjbTasqryCtr+cjvAF4t/6gjTq5yW9q59O0SLy+LYspUbwxN555FeEmnPw/2pQYe7SoCRwilF
GwaaW7s7Rsm/y3sGLKxHrTgX/FEnvvTSr7G84EOrf8qOJeI4emp++c4d64L+pv1Uj9cu33Zgd5iD
jaaLliiDH8l0TdkDLTq0P4nRGhBZMqssje45AJWEutoZC+tE6YoTHncecdxqtQy2gtiP29qFQ7q4
ByoxZA6UGM/SBE/ZuEmx5DhMhYSsYjmb/+I77fYI4qfCNCEpmb8biwtneDNKpYAFG+Ld7z9H9S/0
r4NPIzhGHjpcinkfsyf+KsSSr2O6mEvpchH64HfhktfZGIjpIf+Jf1YJR4L+AT7+u+4tc7nOQCgC
tH8CjktfknFznM/b4VM+q3ncYdLHt2PRPwu4WFJQKAtA4LC+2x18C7WwRGRfE/CI2LHX7d1fGNwm
Zl8+/RcXNcBdzX5GW7/ou0VKuMoHKzrBSG4smHlqe9s/299E7oAUYRqjsLw6/vCf76i8W94knr4T
36RM8QBGE1ryvm9QdABCDtM8mmIlvZV+HW3NIimBZp9xA86jrWcQmWagZWkYY/B5zXwq2C07CXvZ
1kmrE3mEVht8tpsEcqlG5kIRehYK0QDkd2VSG225ntgAhKEWP5+6R3aK8Fg9JN088+PcdTHoYgTx
xQElxZfkmxwRD4tQ37ZzbGJGetOQQxoH7VjTMZRNzdWpnl4xkopIMwV1X3vOBFCpxlvITNkL53Qm
r0zebc5fZlQ1Ad37pSutTbrnux0/IAbbu1LvRKX1lD0wsZqVTatzGqwbhMA2CQ9BTp6WLoNehzUg
VwBxZ/pSNs1UZ9DGHWEemuR7i8LjI3m7/cElCROH/pKQmVLtQThpmK8CZUQzbiPrhM25pyP/JU5c
J/nOYg4m6841noQewM1v5cIvqE5aFgSDiBl/3kHKoQ+20UfLl3XLbsc/n8u+KXtFDOa6SYWGuKHx
1YWDdt/qOun+mE/LZGbAyB8owKfmCZ5qgRARb5GXpekhGY8Xcg2nJi0g/BaWY+IVEl6DHPY+eB59
uQYscMIzRPTdpdwW2C/YBY5LAdzDliCV4JNlc2fi2hMEB/TrjIwfvXHINpHveBna+hQs55LUTPig
pEI0Qdiyl+VNlJS++Juw+Q0r/KhrukU9Z/a0Qbr+KxXsU+2q8Bo52vZv2am7fJuae1j/vvaFKZgh
+3SQa1mhevuegF60GqtJGOjLInKU8rBhOguZradeh37LJMRKoCAPE6czqDlAtgJXUruXQAE3//7N
BA7MM1zTw3pk434SB8dCo9Jlilgx0om5enHO7k3C5g23musc1ZBL1bfCgXL6vNP9xaFaxckkHOaA
SGROqJPIuOMv5M2L7PuyPM94G1HCIpxceNJVSvW9Ps+cQnuPpKBjc1ixoCYdDW3yGyjKAke1wRnI
c0UsxrcVanNuSzFY92HtqG8Z5XptSlXrQ8SzGwpJFjw+ILKrYRrkP1j13xNbz0/N9/Tq5ZrozVvi
O3aeb+DNAGeLRRREOKrKDzYMJkQbmtBi3iorRUyVJ517cSWZcvcVXi8iGoWR+44hQ8Z+GUMN+Aio
tDYK8FM7w1kSL0ZUIOiift0WVgMtnjl9iobhrfEVPh88ZvHkWvo2XQCaGRhuaDKPghFBcppJzGD8
DIWtuiA5SCp5yqoEAv0PLPB1cEfxiKdNTSZb10RUF4pM66md2Bbtvl3k/ww4H8M83zz7BUIxHSHZ
Svntr2VmOv6O7VVfbb0jPYZTJDNovlXvnoVPbBBHAC+8Mz2GIbOEjKwkU1J3xz+RDGIFo+5+rlwa
oh9NCEVEXxYmK6EdbkANvraAsvtUcL5NcfQA2XrkeWDVChK5oE57lxiv0xpkP9D3Jpo8mvAOJtYN
JBabujdbx5i56XCH5UZOYLO4UkW0bFNOmab6JxsaUeivsLpbqEnuAsfCIbuUxm17HnpwX9/dpBNS
qCJVSaA9hXII0elBlSS3YfzCsIqxY06wwICvUpijlIQUiPbGmgw5ys4fFO7zXL+rD0qW3kbmndM3
aFYg0jd2cBdhLDBD1xUq2Bg3/6fD9muJA9miw0RLqD6IR4aXagPAwfaVN710yhveVPDEf67yHdOG
GYOZd0NJLNy+3CMEnkKZy2wKngug8wXFOxcO/BmNW1Gxhdowvv9Gz1jOohToSkE+IafOE+yMYT5e
wJmCWp7uLlVp8OtCfJbmy3g18S2GsfkdwcxVMhpBPhSaasEtowD7Bn4MU8zeTeJiIJhhigt4W1cP
qAHAJ5x0NimJCJ0m/9Q7o2+ogicrlCvnAqTpTWuJiwJNLmsAP5r6MNWhmXran2PoJQmEDmtG7T0F
C2sMvhMDLY71HVsmQBZdTzvCcD/6vvZ/Yq7BwpRfwvye5jDwH8o7XQO5zhTt1+aJnHSfd5Vcxz5k
BgnhtHOz39CCUrBOLFgDUZXpBu4zms6qt/lYTPA05hk5oUAeHgItsCuVV2xU5gTnjnar7T+Urv3P
7XolniC3jquOK5TGvzlssEfqSOGHmJSu5JjLaTJpwEIMdU3aHjDYZMw34VdFIsWE07RQfHpNFMmZ
PbJTvSCnzxCzidx2SLXRwE4ogEJm1+KBlfaSS5W7Efm2+gtYLs790/PO1HrlEz7yMTlJtlLUDQ8Z
zmDmatVbjtUOhtMZ0xX/H1dKpC+JQ0bbcg9lKgZIMv4cHgsWcSuJbiNWSbp7LQgoqvUwiUJxv7qz
HaFbjzvleFW1lXfo/wk3925eK9KlU2yxoHbP21f9QuS3FT3zRMIv6wSIj0LJzPEsH7k89D+7UgeV
1+HQIifIlj+uyiXHv1V4nZEoaRUqjdQT3kH0gFxl2SCE7jLyIIUogSONeCjpJXtGGQVUJEmGbaXI
NQNqBd8XUIBQ1g7yaXIYZDopn/13uZK0VUwHXxCxjEFzDUNSLJzDHUsZjB8cJppaUt48D5Todqxd
24zbuGxyCI2E27ZaqAgnMztOEXwqY9eHtK8lvA6ZezJOGngNNLRq2/7CIZDXgK3h+DU5g4JndNLk
62SWMY8FvHAjYAd/XxLRXkWMC8PDVYRjOSIsnKpMHecnsPCsoD26VCD1/hlRqRY6fL5Ms2NTpXV5
tGkmGTbgbkE4fo4DBMwqMpi78/+dv3ngB1NRqH/GJV+iezMeJXAxjYEdklCGx2JbZIsuqn0NB031
vUuVHE40G3luYr/u4HUiQuLHGcISyz7RKqNJNPws2bZru+sCjdeQl4anxoz9NHwxuMnatI4lZwiN
pAgp0PRJ8y2nn3Ec5XWtLxcxldFn+ifBM5TszMARjq/uytv7ZWfJaFZqJxw2jTW2O8F9l0P7TQc2
S5Vr9WxdGXOerW/DWp3o2gM3AoqDljE9dQf6t/8CnWzja/wpUPrfBWej1KPr+VfSpQmd4/pPccFa
oHOhjFDieWZqJfv+tc1uZCR7wx5RCd9blvvdYaGN8Q6gRHf2IViCQi5PTv9631GaEoGY2TbO4iFG
oxDF3nRXfIDqd6ST8rltmMxbx37LYeCOnDdsflsCfBR2EsCsGtQNP/I9/qmUrfjC7KXeEuFbEzBg
MX1NxhkrUM0AHyoqsJJZxx50ffHh1r3N9o+q+T86dSKxfI3a3S0QDqm/9HPBvzfsnVIdcHJemLv8
QGbzcikbIEfJLXf9eedo2/vKKqpPsQa74BgtmOTu2faBnXkjg3VBXNOJ1Hv9K/fJO1lG1XH2HMEy
TYQiAo/SBW8IcEmc2HBuzjQV+sj5t2UaAYI+htyXhoGbRTu6+2HHChLF0uBWKtqlnqeCa3ocakRI
7rDSaVwvB4DfH7g9FsK5Z/hXcf2+wXWV/6J8kWF3uQHYpIAjfwnNRhgk6h1SjCX6JsGv6Ecp5cOg
BvIWsHdIEYnZOCor35f4bla8LJw4Hx5qBU/zD2IMBfeevPdo4ch0xL4SqQ2X+Cx3rAA6Jz+akFDS
mJO48hxuNr6K8CQKdraRtdHf3GDCBfnXC9qJYxa3gUZSEvzu0rS4ClwN/jsM79N0njdSrQpYxdML
Lt7qBAwbaxTFG77VyHL0bpIzh3OpRLFOI8b52ADRAPms7rkDY969OGzGp48z6fI8ntM/c0pYzmMd
Mq4yyKb+CasFAUlsa28JQraNoDJ2SzXhgG8N6tfAGN/cE3Iw1cDhz9kY6EdaNvcuR/Z5KHyxrNRh
YE4bHMwIVJWxvK9BcuDdgtSZEqhE5g1ZUjmjONlFZe+4wGmBqL7NqZq9A1qv1s/KuuKDBvFrEi6d
osC7Y8KbxZFWSdrQ5HcR3CU/fbjKg3Us8T0AZEtF46hEFtePZ6wgVU0iEaYh99CzRIdLjbK/BJfu
d8QbKOf4hdJs8V4t9AMfLPRLmx210UDDEMRFYV9pO000/Q8Ue3CdvyV8awDKCA+xrx7BkYfXNsvA
XrJpM1lMlKNuVSQxUp+kygO+dFCAlYI5uvWA/7tXhHA6Qi/rfzrN1l7ryaMX35SGB74ARquoK2uy
+9ssX+lkcqLK2WoGtXBybGm0owvxPh+DW5kHSG6wsw4bcT9eFGqWgo4SJjbtUMuE0nbXcKIcQY0V
4ycHsXsx2upvAsOFPLjhNT0o+I+3nU470MQ5Lygb1gNhoWxMLf1U0MpXnYVuDiX/Rf+lSufrdjdg
Vyv4TCCn/nu5EFAb514qE51DmBKaYJUulyX/LGR8XzaZ7maqAhe8McfyQgWvLEkMkDNBdHA/5BnO
1JCA4PV1SuRre7XrMz92p4QCBCO5eel1oXwna94pQQP/ySMi8GKjlhs9ZwRa8cUecaClrc0PLL01
9eWhRetbv2JjPhPT+p+QfAXYksHvMDaZxr/PKL2wotsP1EqcPeGBS9sJDYR+FVXKfIjm5p2fMkNI
I7XA9F2j4u43cGZ27CaclgrBJGF8KBHX/eGQvZjYhmcpSVEjxEUmLItkIOi6oL7YDqu7IKj66aYz
aFkskyYzAHNXXo+DplJIhGLq2foEGDtaEjwkkuhn7VKl0g9+tz9tx7R6/CcUIFJJ/mX7K0/h5Wxx
8aiSJv2FT/4FuBbEBI/YVUAK74FMiwuclB/FsVBecX8p0aMMdnSYvx3IeMb6CY3kLseWCAVx6iAQ
C5VwKHw0pfsteFh2vYTnpMQHTbepZskZha8bxWnGCmfc873/gqoX8yOV3RDCmhg3h7fnNv8sUZLF
0+Aec/NozaUc+7wKJFXO4Tde5iymxnoFlip+aEND0xgpGc9OEg2c7bRxCxiVlrKQIWZkdiMciPmX
NKFcFrtd6bQ7m/Fy3OJynrIAMfXVh1GPM+WxnNgcaWrdi2c5yFCnEk1kXJZ7zB7Dx+oIXFR5PPIh
smnV9XONvxXVNFl/PSzppBjlJEVcegFxulGcIadDjqMeaLnuZJuPiNmTNi8F7/HkOtKOqwo8Cp8d
a0LRNStAI3DtGHtfZDg4UGs5KJtdFTN9B7fMfTgCmyJArLMr5MkJJqpYuidEyEwUdMRzlb15Rv/1
jPp/3YbNgs9xzkpJrL53IfiiVxc1wuauszDHsNiaCYneSWLHtJBMK+/UtPmLXyd6edZpcnKjcrsU
P3+ulPGEXtHTS2xebjy84NMn5TgLsQ44uysOvR3Zlx7SLAu5wkGcCDJoracLq0FXWqmMsl3hB4OE
qb4/8LUyko02nuAnj47PUeVkNabERDlK+z18Ss8KFTPzYMZWXC9UwEmQrJrK+lO3VBGS8pjHs8Hg
aa1jrkXYV4pe6zlSERDRbHgdsbDbFBgCJgbmKT0OkbM2+5PJPI+4fc66aOvYYLsA+9LlPJsCzYR+
KhQUf/6Cr3eyD4V0nkSQGqDwIcsGuNSbz8nlGFKj0Ly30BPqw4wVXFD6izG9jBT1iMBHQlAXVdJs
jdDUxVpkoCGpyK41sgQr4fs6tk72qGMJCiCokLnudYR4o9/cGbsxk8QdTm4A1Q39bdk3rcxEYhOG
trKQfoX2QjNNKI1svRqWFqciEvGrXNZKqElKqq7rPIrW/7fIAEZNxSkEUWxrcKon45W1zUiHA+8b
T+I0jbJEqoq9Ft60V+oigq1lBKc5C0XQ3ZWTdX1etR+CA/mT6iGEfGKFquQJ0O7aP2R+xnQLRW3V
TBrrCYZsXiXqprl0c6sFGTxWn78txCLkmx5xpZobz6R83ZLHL4xrBAeIpJ2Z+VlkEoSs1NwWzpnr
3uuIHgrTkiVCoBGLATUaahBrWYzkYsw0z1oTb74CfVTUtZAQ6A6QAiJvqkMnBBkfi60sG7t+G05q
yc0mDoi3+KYyGEtDT9v5SeAeuxJGL5nr3VB7pweljjj3jnzLJ7Xzi6lQZjVtemumkfkgGDkczmKe
zveMjZ8DDtIqA5VZmjmFhOvuYYr4qd3TRAtzBU3jbnKWU5HJLBlNetYPui8zgcHMsO5raNqUS4Y9
NNceTB43dGsyUq1MIm6n8x+crKs+RPlhp1fKywdE6eCkhVQCv7MGSSYykjqz0EcLOJebCMEUB5Co
lF4IAOx1ucHY+UdIgZaFHr0NUdGNK+eo5QPmfBEkz5kaD3rRDbEeP0R1NUQaH9w1lHFmB0ZuDcou
2EeO+e9A8qHii6lXq1Pu14FNv4HoraUu3zRot/xvHD4x1nkXZBOrSILzdbym+DpoWYpVmdtDz+3M
+dQLji7WuxBVYptJ5mgQ31wDEpu0D1zdUlwEb3Uh+l1MLojYDbSBcdBUF+o/xJPWtnEVsuWXn/B4
T78B5h4BYgx+MRbA3GzcE8HQy8d98RvYxhxMSen8gpx+gxUaciGe4tpZGOuUw7/LAnaQdGC4wWmm
ZhzVB5cuR7nts0708EaDCQ8OBGlBZgnnnmOPuwapqdPVDGmlEEYeds6/irz3xwzTdRpAiqLMnfdl
JOuYeRxYNj4sq5C1RNuJCxAh+6qmJj0KXXcvKjceOAGORpVb+wQVdXwUSz1u4x3rvqlgsbhIwF/U
5Ey48tMJz+MFgI7t6vHG4LNRO9ko3TUPXxEv1Mi1qGf88SCfRZpo5IMlM2bvqCJY7YvI0fSkMwnV
2XM4tk6WDqSJ9AIagU51kqJ9npvXRoe7+/lmD/V/nG8mMtGAl/RQeydH9CwKpl8vUhKsOK6ohJ7B
ggU4EEEJrCC6fyfVSx0y5nBQARRO30YIegqh2nGIpCbBOdQ17X+zUBHnfvGWDejukbiwOdnB+ht6
MCBoinph/10ZPHDclYcA7gegHWRK1ruXkPsOn121zVVboOlvIqrYjUOxmS9Po/gDxrp0v+7FPqj1
EFAgQ0VxC4nMcmVFV58USsNiBW6peit+ZZYdbKWLJtpCjr1d81Iwh0lUv6Iupa7kjlReflppHF1z
5dRGI+nMIyqOu43Khm56qC7jBoX4nJ7ImL0uoFq9xGaISOrfwJZ4o3e6fMzUHrH3Xcz4RF6jJDNA
ttAwpC1XCxTbJ2M8JGvv8mWg+fOgVNzpJaGk0vxYD+4tu+V7qvWGEbQWPDPlJ7oBsZyA/mbIYBnM
8Aj4GGj8wgFFiLFzkHOXnVlnMxfdYPUBSY5IVqmENWmKdQTN1usX5fIt5qSapTKdwffYwtb70LB7
lCDgQTaEpqtBjhBAZJ7EoJxmRRCPKYRch3g/zdzJtO31s9EAhUGmTQsoYFwQ16Ksr2qOgDktFMBO
JViNnIpsZ8evp8vGRnsA1Xk+eM7iX2EFc3La1FouygqYtnmS67xFYdOs+dJAo/1Gz6RHjx+U4s1A
N/VECDxsGNY5s99QaIKFksRO4NwNSLGB9tE115ndLR/YddQWX8Mh1tFSUGv96nDW26pjBdRpBnsL
KvL2HB550nzrAZMsnmqSRVuaFVbY6/2m2sBSschLOd+LB8vTr3j5cTWKlJ2K090N952v9IfR5CQR
+H+K54Vza+za1U/8dcL9Qy0khux3lClD8t9mMKj/6H9q/og7m567X2d8Pk5VGLGOmAZKnMYBf+mp
/BC1K1lstt7//uGi8iW1ScYfL7aT24GMxN1YOA6RMiHwuPT8oIAvKM/zGxtIioVGE8Z3hlPgpT3q
inJZYdf+Z+zdQxd+NE8E7xVp+7lNvNp15MUm+ty9z+yBqD6gJqma1Q91PSsoYXO2f3i2erIbBrBF
U8ru1Y2qy8X1JKS2klOYENAYemgQZxDgRX9OjVxzSjBuF/FXZ7ov+Hg035dAVe57ctVp/mT8SFZ8
Aszf1BpET365PolijrtMlz6uPt46PWAiA8vaP1Nxq4rPhMIuk5M30bM8qhGzcObfPXM3VSCdUTLZ
/45k2blGUY8qlYKMIgEQJkdnus00pd3k/ZQ9LoiL4cPHm+ibJas2tyrW1l0ns731znylBhfmWYF1
WzEe+udYA6Ii0hOTPrd5tK8uFb9R0rm2Rvr6FTSzfmospYjRib1ORpYYCiDBnsb4YUeW80gtagny
3+xGceH5ou3LDMqw7v7HTN8OkYbNOumdt3XiXnhbWymgD/aIsPjmraWNrcgSAQ2vJemz1EmrFr/N
bSyxBLpTZbcfojX7gkFNZZ10dnJJcbn9DeiIeHOrhOONArnQyIuXd1D9ua+lVjtMcXprezYZlcv8
D2nrP/QMCyPd7qHbAj0JkY+pBX6eqzSsOWxjwqrTv0dMXA2NUYhTH1IRZweGP90aaGN1VLh3POb4
sFJfzpJKhm+clvEmIOrPpdu5fIOU8O9XIYLZ8GbiOTWi/9HypjlUDnNbm5N/VbAoblxqKqP4B2Fa
1jpP/PYypSrXhFOXb70QRdTiXLB6DngXDwvrprmL1HCas5AKUACnXt2zcRknJ0YWKWKqegVyHxaG
WxpCA5tKyVN4pStom+WZCHyFaZdE52RbrEdYzqR6wiQG0niNNrLgp33deu6JTDNlPlLs6t0jOQmg
pZbRtlz+NYvqc5TPU1tdLzUmj+GA9k+qfBP3Mq+S4nEDJuWJKnirhtdyJk03BeK+/eKoacNHTyYW
bR6urMgGDOcsqh6MWE2Q5r2ANNlJrcf9DszIaPLbC0z8W7gTbB3AGf74J13Uhy3t9M+ka3isG1e6
cryyLShe0jiQ1SEWXnpifdpGeMexZgT61e0dQMx3DNBgfIQwXp+QPOjKGx0ZYV08PKrSDvU3ZgNA
YYH3s/+azejy1SyjpL8jdyaZAJDuod83xYBPRC2cFwqtdXxRxlL05/YScfJrRtPojZGDBtccWoG1
nLB/rSo/vwsKju38uL+16kmmVn8utde/wR80zYopEr+YRt6Cp2hLOBCsV61imqRzA63PYLMa1JHT
pt1pKASuiCe2dK82dn5QjW/5WKphv27AioDXTo3rcvtS6DLYzRFsRxYQ734WsN/LzuFDbZ0ZJw7k
+EZ0pZG/OmxN3DCaU1rr0qkCYR5t6jAvvyOmrw5HopJ3WJuKFVQMSE45eINk6fcYbyu1UIMwT9jb
umYd15h432bkSbZs0cI5KXeIGHoOV5czpW8N72xOOaPPoiPJ4Y4YqAmuqyPdTOIXBMhfBsAJXClB
lR/M+2HQvS9awL39NQGam9ZKZQMN0PBE32Y9TUM5vM+/OmtIMXl8X37Fb+JuBYitwHpepcP4M/Ti
YY7AJEm/vvdCbprg9clK87utoTZS+AN18PUaCJuZN3aqxtFJRSY6/oqa9DI5v6Acs45pOs0sYV1K
3hia4gXzNm4K2V2d7Fz5GwCdcAGUvXN5n7nSXch79PDDAFeRu79dqwfOGhyv5y630cGwt6Xpb4l6
cALGO0o5Gy9Qd9jT+MsQFrNEzS34GMvSoc14aNuEIRYLF1LWBEEMtDrUgvsVRyYzkJoApNDC0RQR
o4UwoXTsUqZAi0hz9w7iTySvlhkiKT0un1j5cZYiVeQRnMmZJB62XSTk4QoJEofJi3pkvDJ4NPM/
FVKZD0wpAQhU2fJqmAGYkrCNxuieXU4IkZcc2x9rczDXkE9xdXS3cHMCQS22T8hLXgFCVCgfsTfB
84wD7+qxH2QZfP9MkW0Iq2Rccs7MxON0vMzQQ6QlshRXu2EiI4UbyPfCdpZgfOxFZHTWnScYHvNv
cRiCu/G8D+1OGk9N1Egj/bJQtiBCoQs65Oj+jP+sobJmoRN7EZB+XqPhuD+ZRxgdaGX7P23hoLWF
/K6NkeYDnWA1GNbmumZloD6Y2TIvztTcmpGq3eZ079BgDO6NNPTJhtlUXO8+MTAhMcULcQMKfBfq
IlUT7NIWtA6GYeBEURD0ut8w3lnwNSzwRyTitzQnRHvRR3O7pK0GS/ge1gyxDba/4km+SoT2CRlT
RKrhugXS7FL+wf4lNfOUmftQu9RwNjyh4asTlmYtk49uMM27vypxCDz4eq8Mi7IUjrh9xpoH2Xml
xN6TlWHjnOBpz8OIJZcY0VPHqO9ZxGqm3jzBaO/GBOrrGfh+ZFVHuAWT03ySDyKmIlnRVs5w5rb7
Odf0l5Mg7zPTb885W0nrFTsR3irLeURN1KhbUrasO2Qaj3IpXwbHy5jjxlmoffpyGFg7PXWcCN7u
p8vRa63M54JjlmSmuhI5XEfqKiCMxaicM/kGgVzMtXYh53cPi9Hjd9qIogibolyLRDE4rGA20iDk
bVicwAztRUA5yxzNstAD3vd5FFoPC57VuLJm/6fG0B45+da2t6rHOyFCfJV94Z1wqnlQ9JxldHIb
M93xAcnqyS4K1OKb0wNsKx0wy59kQOGh9gCcPkkD8GxhzgJC/wDi7aNQpPrgMORoY/gSJ+FArnzE
xXQXSpPOB1Bfat+N3vljAoe5NjhMAPwqZX/SbZCHAmOIeA7yy54WxEY9Kke6pB410bfYSBNYJbXm
uATKqYk9ZgCgAG6eBkSUROQdiadSAQunkn2VYuuMTXmfrD3T4rrxscATOpKmubfk0Tnu7oU6n3bO
+E07xf9Z1A32SSeuoGCoOZKQtkbNePKE9vJkYKcEnrMcUC6rNI8h5+f0v83THkJ0ZD8BpJdKQoh/
RYdemqTnLMFDs+jF0QUju+zKIeAiOePIsp85DVdNp9JTFfX+KRLqCQftQ4Q9zeajCsRW4KS3KuMR
A6Qve+vdAU2L84RRnOa3Sucq4NYGBnzDaRNZc3Kb9l5d0KZ0qtIeY+1F74rgYlI/tO47VMZQhx5X
L1x3N5yRfv0yUnuGOQxNbeGxyvO6tQwm1rlowxQ1TzOV9equkJVSsR8eCHpgV80UkGs0lur1ZTX0
rFKV14UaxiQ++CaZpuRvU9R77x+BPvt27TWgNIh3HENNgWpJIVbd4pxxArKmypOkQU6UxJg300MH
jdNg5jkTN7Z9gXG9buvGvdYrI6fHcnRxvA69O7Z0uATqFoGftIX5IEy5AyIGX0zMxLErVJWbfh9u
wX1xZLkrcVbgR7PRvzfmtZHmMwCF7irywG2q20unqjq2NBdiq+AGoAFbN1QvULDWCIYYkHbvY79B
Akk4NdZ2e5k8ibrwbiBMxYgwQOwd7u4Iubi8Gcno3Whb2ipWdxVi2YUDyLVl81GC64ginqcKXlTw
Tt+1a9Llv4El7tjoYz/W0ew0JekNVN54rLisleVKtYbOc1HweLIA6mMVCDQ71iItkT6M3S2a9Fp+
oDG3fM21M0fr/NDez6Yf3vMPOnSvILftzly494xDZsn3DDHsi80wrCy1+ib4SzZRjTbanYvj59Fe
8ynRyMgxEt5RyAqrrSBWxO+9pPjPP1nRmcKdYLZ7bf6LUV9E8tQ/R2T/aLZKx85QEkOaWvt2T/XP
7HJcWKkyp99Idc6KiIIxeN3lf9R7fGgiy79aHHDaDCMzmyiqnbR6K/N7+Uh1qpzrbeWX2G1e08hC
1JCDplRPqKFO87pUFkm0+LkgfZ4GGP52/g4asYTP+Q5NvGG7pWZCcWFMJsg1x5UruYfjfsnxRs/2
GxNRkGf1VO3He0offP01icVUNyBAzVb/Jive1Kh8Jd3HoPX6B+AKf0Opu52ANHAykiZzDHma/AAw
v5WD4cVCBs+lF6Yik7Kax58angvAZIm9t5yUXnSWFRxfhSEJjhtvqVIIlQPo1looxWJq1WtGrxB1
jFY/dbHiVcovzyYXUrtPmnPc2EcoQ5eAJ3LQbi5TnAs0aoHR8stfzUhKS7L6msPfRHiEQehq6tfj
oRBBXgnU/GuBEhEKknYY+fEK+NiS3XOlI+l4E8fhHUhxqVZVV8zO4BQHIjGK7uhbum8mu41ggB9r
+3hxl7WtOhoqMOoTS8gfegsVwxyNU3ATYQBN8itvl8439d88JDszhB5LRvV3O7LtYT97AEDpD7bJ
c7LWysJduV7IwcXh8R9a9kOIsenRH61PYCXhxOe3wCKDbbozaHgvMW6yIwdwZTVD+x6A3n6gtbk4
4KEwcXERURBlTjnBMhMtxZahIvdG0xJjNPpgTJyGUfc5azIzDm6kXdCkSq+HeGfy+Y0jncyE+ONe
SibOm6HyFQGjbUJdtFmpQNvuLtXN2748i2VcYaHsKt4UB396B1mIB20K/3c4BSTpv4CqmClZ8lm2
2aJ1fw913CD0m+5LoeVArXvFEqugBywnHA9oOoQwx7igjFTBZaBqJciIlJTadSPEF9HidFyjNSZ5
IzY7hhepvN7/w1ZvCvcJpTP6x47gid6sDFHy8NE8dDo2h0xL4ViB+3HANjFwlYJqncKVvJyAGBWE
oX4DC2tDo2m9TnTN6FYG74L9/CxBidNkS/m2fViXVOA28DF29Jno6aMzw2M1SRZYEFRMsvn/Ef92
KS+QZKoTQjRlI9IF/npDUrhw8EgDU+pYDxQKO1czl2mSLxn06mE9hNNg+dnoJ0tpqa9E8Zx3tRAn
8QjiSZEbg74xz3D4rYAIFvNbto12BHFMsZAn8X5KZ2/FmmSoKCwyrryXA4X2VjCN5Bwe0aU2hIkd
tgDscrv9fLeoMzRM3FL7MUG34wetU09LGEhdrWm0qmO2PaAdVirpr4yHg8RiINSQCy/t4kw1ZoUi
J+hUiNW5yltrIe36zL5v9w55ID+TZ127SV4t1qzVDARTx3Ns3kK8tUAFXP0aM4AO//TGGVNaHa3f
0xe50VAniNRoGbbzMP46trRZ9PpPbodyqBiGfaDbEQtKf5h45QlLXn11prqqYJha1k3+rklh8ptF
GpbHz9EuRAiQl61haFtK/N7TXcm6RSROflkj+JZ4uTU19FHajnW3YaoeJO0n/vvftNYXuFZPsgXg
hhjBS3HZi2Pbo8TO27meWJrMdxkygnWeBrTfqHcnAJjWH2Exqe3YYaVJ5M4wl0lFvXTw9vov8J7e
Z0TRMf2rmVsI9YN5tYIgaed/0A6bp/Wnflf7BmIwsUql0dSm9QKQLnAloqyuJjgrLOqvJNQhtlhH
y8HFNAvxkm3H3LuIHHa4c58C9QOfpb6SI1AWsPIk2ocqXD594E2dAfi4hyAyUCOsw2I2/g1U3KJ5
1HCTrwI5grd+9wh1vFX3swKaqrYbbBXOMnaPvtYZ14a+QggzUluOdvPsQIR24ITUGr3487fqMrVc
qaE09l0PxbGaf31IhkJFfbK/7+S1bdTTkwuNslzLGvLRc+JEEJRdlfIpzsSs0MGtyN+us8+uGEn9
DB8BArohLBVAiWqwjJLO7TdlVoV6VuoJl4EbJEE6Uz8V2MwAF0Dk5qpwRJVuOGG/nMM9UDLFhJBd
DBcSXzvklIH7Hdzemv5Ir1WugP3E2xfZRHuIsgNXnohl3rzjJOmrvtE+Twcmbd7A+FYEz9FwK4Mo
H+TqfngCZHg3H/2aYvBJxt8SK6zdsokymocPYcg+gMLX5ZclKIMqMs4fz2b3SzZI9whyQOAlGyvc
lZDW49CCwEolGHcjyb9K31n/YyjwDOeAmkMYwJDqnUiZ1Jr7oudoRueLpd2UBFFdcIF5u0H5yEqL
AejR3Zg7ZuCcZ6qJYIBeX0xAcvFG03zn3VQCl3SgFVwpXFZKmd1E6U3LZAiXpZafSX11LfTupDQS
PrHW3Z87xUdpWNT5jXj2kSLof1/BckMqEe3HZRgtyFKEbR0iy6QlBKsoHh9uvbLTJoHs1AuLbtR3
XJPlwX/II0nisp6+vi80QyhAsCZ0APE9DVTfIDw4eTY7LjSPxYnfBylFrbXLQ7FueFF4GK/cybhx
Y9dPt0BbDXFKERWAsiXK6un1I4jE0MiV2TxP8vUCVOBhHd1dQUI+chj4X9EV+ng5cY7YWCbGvUc8
0eD372WiktPoU22HUZAh+ZaU1MdqMYMvUfKoIAhwN4we+Vr8Mp4uiLKYsd18JdAFwRiFZevqx7dk
7LDJ096VQk9ph7zKnITrxesL0/XyX0E4GAOo7Hj34c45ThhbIaXRlNhcTmvZG3UYTygDroEJb52a
0HsmfFZeN/OdyYovpuMJzBtTr+11ivwJaUfDriRXajBRs9ihi74IvgdzQ1sZqMPs1KB6ENDx2p3q
Sk0CYw0nqBxBeRQlELQ9HxT1dxqJHwkOv0AiAHRW/nLWB+xsK1FXjquwjRIAKxzY5/zNKcCg9rJ5
XDeoDE/jAbXhsXrPEeYBcDNT+ik0fePsnX6DRhhI8BP2XZ09Kbikpas2Edg6ycml16AqtsYiLbse
yjA93Up5N6+YJC2L2eR3jT1Z1VKnbLvM6QoYv84GFQtCgnffOFCQ/WUXndyNdjsQ93O+Vfb1juKx
53R5bjq2OZxeY2XGDPJVMih9+trXZBwaaX+sSmFdIdOsT2UIF4zPp50GX7dKNhb5at5b7h/qVMAo
JycxP3fC11npFiHpsrgXH7Uws5tAa2iMYm4CNk2+urj/hEiNfG903kX/HPNrJTFdDrl9RmkbKtrc
uw2bUuQ8rw4xI7yYaixlO7ADO1ACZc2jDHK4MQ+606cxzouoPvHbpivQzDVvEgKsibuixb9X/zKp
VafTV9kr8m27ssB96LxGDYAI90PbP3CFJX1qZrGPKrxgXX5Z61BPZ5YzY1JagK2jUHGlmodlf6Ju
WK+WmiyyFeddyX1SQraXGqXAK8JdBzlzkrFlLjn9Q0JalcbzAVLqD7ulilzWoQPmbYTgw7XDV1Ft
/7Xl/wTRHnPy1aNVQ55ck9rvANor17UQvDXkNFY7KfrSJYf5OH8xuQD9dOdTotkgyhte+Kj+hXut
HFoucsLrMOsXn/eZK+x6g/TrTyY4fx41UnAIFvNPprEZYd/bXkFAHibpKcw0c56W4ZsITCYI4ent
bBUfyNdDMwwmc8JrBys4I5khtYn2D6d7GlMcMUaoT2ucEiC4ZcfEcHOvbX/TGs2dpD1udc9Y+z57
Zgyhx+zb9aT2/3ygVGJuU6eNp2297QOANMEKZypszxScDWqbhSvciCq4qvVkLIg+H9K1mKrnI7ss
2IAIjThmx81vaK3buC7MV2OILcDOACO7GdnY0+uwpyJPleVIiJXNLU4v/lIvlR4Yo3op6YZtKOL/
SSpSFZwpefLF3n0Pg+E6rYD9VZrVFee67MohTWrxEz9ksUZzNwEEZkviomhW/SAm0rDF1w/SXJ6y
8H/jnL14xJ0rivyrNNsx9UpyNdptlztyQ5yldMMHKOclhJsW3PnMGy6xWRMbFXFWMFYG4ZeznhZb
2mX6RiaOwJlJKhemHBVJDgMwUTg1WrBT0gjEGFrBPvCSgZT3MO/7lf+XyivAjXBW2DI45usUheJY
leD6aUp6WyJwMvEVLb9MnzWzZ6dupNvCm4mziq71+L3xGpdhzskU0UbSrliimDUccENzodEiV7WX
O3ZjVQO/0tE8p7aSrU7+STKxY5MTG4r6xNRhUrimEGf+A4CKXVCghlm9e+iIrShaU4MbQC38jfnw
KGmsFH9wOmIKKpQCFPi+FE45tOGFCkhgawLLRGa+btj4s01QR3VkxTp/IGtmCSViySCbAjQGOuNb
IxltMzsiGzlq8nKNKLD/fUJcboCHOK5eR11leRhFxUstWxACnAJx8vcK5S4hj9i/ekNQnePlilE3
7QBLd8dl8asanbwxqdkC2LpXsTbg5SZbKSMBnm97OO8oRiWFwW4Jc5806atNIP4jAM6eHH2nNoGQ
HgIActorSoAlNHonCXUxYnfHQmdpFb+os0lYsFK2Sbo3MAuE2GcDOiSzuAq/r7WSI847DOUm8BMd
NNVhmsp0XmUWTBxsXVz+uGUgOOFrx3u0oKhTdbCs8HQvW0DIP4jaALaA6PGQDUqNnXVQjIkDWHNc
R+ZdWf4JCjCFk1IgeDsqzgxkN+wIj2O/v0LyIzESLjUwVBNm+5pMVL2kTS67qdtyZVC5sbozCncu
nrBbH2zbGOW5fYakcpEfYlTiazefOhEvjOY6WQOfeaWLZ0X7Qu2N8dRZS78EdinZVgDO+nha6hZo
rYPMI9YbxqJqXD8o3h0hfThArzOjKwEzsZ9WnWcCuAkuWOckTG8ODP0I/9VzyIgvaw5che4oMxKh
ToGXHMwpT7jqllm8QoIWSheQTnU1I8QShCyKhSnZ6yYLIOUgKH/kATDClL05GQ0Mc2ukIhb8nQWy
/3SRjQITO1O55Ricu3bsrwU/Q3bRU6aQVH8aZfe3U+ARnwK9SHar49SAPHcYuzSoFaPVzePnVOYK
RhlQmHH83yeXbmo2ufaUZkvMzhze2UNUFDyq3v8XXyyiOeW1rMDUOidTCWvuNn4f+kIV36TnE7mq
BegGEQ+MpVzI7V+VtPzflWwqE43wrWWaQpqeE2XmFJSIJukAKrNFp3a3N5E6JQYvubytouLkYwII
DSVVuu2mXbsqZxVcaT/RXiCsG2qZ9gK7dFyoKHPNan4Ln9Xv7gyCBkDdI3eOfuyQmdskBUkmQlC6
MZzJiujyT1f9iTWbVUVwUtyRMv87TxYyYAl1YyvIRkN/ick8tbU4JbTw/Kyn6dESVIa71ia52yah
drdUlegYNeaLfgj4kmLJTUjE3dPZ0l8Yvj2BYjl5Yma55vBvkKpSFTaj1MWjxVJOb6q/ZKK3q4Zd
iQvqMSbShT5AQRGW/KJ2eWjlZHmo3bzePWSNxXkJ1TfTqYvRXFmTjEwZzyoyPczguhhC6XdfTc9k
O6Aza/dlLZNweto1I71boWZMJOIm8wiopnqFTQsKQNNRYQ2zO8yqCtmAX1/qwQ0NPknChrpRseku
twTvigWvixMMBHlaSqzoWcyiKEwuzr90p7p4Q6SDByTqQ5NJBOcuQ8faPESdL1+PATlIFaX4J3gB
upHZqP6eW3z/4QGsVXUep3jDmc1eBuFyHerT5uX9Ed7GMQWyVqdjQnWvLTwWy/NMH8Awo/tmR6PK
JbQmfA/QmOYgq9HDAQarGqkCTxdtTGj2IAnu9FKwIHvFuMxTxILK0I0l0ML+hbYz91Io6/RFzkRW
4Y+oebLkrpXt0ifS4kZwMqITmQY5jNoMjF5gS472VhxMjb+2ZsjNeWDwE88yocVz4c2M18P0P7zb
fxf786RCp37Gx/qdfTO+1EWaQY0FdJz++BUrtWf721ZTTuJ0HnO0mqdSh1OccZq3RLYSSQeq/3qm
Jeb7lW5W25a2lFLCqFFFhlDO54RUb2wTE+wTerRkQF0rSGFbqOry+cCyfbRYAVp0zVPiCOAVDJR9
SLepWK5gXaUDt/8qM88WV2x/Ml7NqEYIt/lhOw9HxZzTZr1SVoBQY4fRKjIus3xQxO0IPiNP2vww
HZg2CgtUYLOsX8T16IoE0l3rngdctygHiLD76h331b/TvI5H4medINI4c1s0b1B5yrz4igoN7KqF
pggOP+dQnk5nn+KY+0es4kseMG6x+DexjA0a3wws5NwquBOY1HHwEUv3UQVgXrg4Quco176HbD1Z
eZHZHI9rf2QrOyzY71F0oq2hbbHiFywu3cyl5gK4BjkqLRp6wyGtUww2J5wJYVqQa3Rk+8Cu+JrD
AsGyf0NOrjsP3JVPsNWoosetKGyQyF0Q6K4enZVNiWTSVjqL6s0RMzN7+S6WwDFdpISqMOS4BIYa
4SMde48NKfp4QS3tg4AjR+w0REd1wyTztoMB+8KWuuP6OdlO1QZLaqsvh0u0mwJsdSJ87WjIRF98
PUW9MBTAYBZKBveeBNDZXSb6E52QlNVjuttcUZwD/k1GVM1CKT10HrlN5KqdcWwSBrtNkjF80ttP
4i2MeZzhb91JFjl1PWZVhOaWDXcaz23yztIt6U3RV9UorNVaGPxz15zHx/A7MNZXbPnfD+z7BoRj
V6jv4yfKqa1/+Vv/WdoElGykXg80E4XpSPfU44+myaD4KlzfM4E+mN05N1OKvOGYa3dg0Pqvcz0+
+U4yBOGwrZ/2eJ5bbRyvzDJ6QhljZflYGvV42MVFsU0T88nQHhUtQWjyl+Q3QdNbaFETYovb9jPB
LaR+MyAYt+3FqZXqijp+KecuDO7ZHhNSkX/ybC94+Dhb8Cvhx1QfSQSErCB7ENu97RGLc8emVcmA
1WzNbn3T9GOARjxCNFDFxjJheJulrl02e9X3hNFtqt7g71HPF72IslrvlHG8pPozjVBUF+a7exou
1P8AcSoArHf+g3A2uJ6bPTqeiH0HnlCbgXv9nUHi7hW2SbNBkCSQO5ybAG5jFigSZEujY7rW/bQm
tuT2RsMOmjSiXKlXCSkkLwhlBN79+Nli78P8B32GlsgJCQuznOQn553S2/Mkr2rz9O64Pf2So+Xm
MCDlL59ECfDcA+XnCkD8zmG7ysDSiXPjivphLg3VHekqgaAvzZfHf89K8AsjBlVYX6S7NeaKElNK
KduB+TvL4Ki4rcbKvu/uSooQdvsA1qvhSo5tNLC3NsYq53cy8KquLF7K3yy6ZOtVXKngZzQvExrg
MGNnDONNSR++JA0hxO/sKoO5tWSj1LDJbaJZ//PPrTDs0sX01KKM/CFgBRyARRQxvOUR2YrcorBr
0NLv5o6uPjAuEE1BmNomKtxFS24tW53oleF8dZ2DCIssoYhRd8e9fHoeyfvNSbSrOoKeTp+xc268
H4FBwVbNqvxBfnnc/HTN5elCi5+cNzGtaARXUIpXx55YSEvglFQUQlmPm1mspQMYYYDLORNHTF2U
j/t6JJuFUyPqWZnDckdW1iRiblC/JbEmKEdcVCs88EpiIUtrEw2/y5kN2X27yGdkU0nqPK1Z4M0c
JdqVVB+F/NtQFImsLiV/1jV73Q1jVJXtD5Ler2hEUF5m0ZQPbZYYzm8RizI+uShYK93Gii6pWjbz
G8ZWbpZLDX3r3TFpXuCY/4lJkQxalT48ts1OXSGPbkk6NWMvdo+n57/bTJmNCtRVTDUdtFUacYVD
cUTxem2XrAcG9tW/wa3C+X+4MqeDNLBMc6f02IcVDDnRnNtrMC9VtSubzKiRVqH8XZ09Glz7Gitx
3k0GNgEgWBcIUAWVVBN+nQ8SYr90FM+S07LmGdYoqxmSqCih1WbwZLRisf6A5qGNHVSpT1G2OIeD
+yhWAK4ghruc7nDnBJH30IhbaVoMq8NkQMZdCCVCwpGawOLMZri9CIAeNlf/Of0cyi9gkqi6oMDz
SEGQzd+44C8WX2w+4MmmK4mVzTJKHYWMuebvk5WZMv09uZZv+dFbUjF8jKr/w5TGtt2d7V8xM7sc
Tgy/Jm1aemGk+7FRkavHqZdRuMt2T9ai7j66kBXHAXuiVMhjrZjCZloWzZdGDgUz58FMch7BGWrZ
tNgjL4TrOwt/b4QMALCXp5FBb2rBN4FuxPa8yZpsmfwWZUoroSOkAKBHnVp3l808LyWs/uwcNQ90
VZu7PzzeAjcd+m01rN4L/3hAFzEhaY5Pw5OPdkqo87jeGaRphXyzLoKV9Yk4eVZJy+5Ar7iRHQrH
96j6Tnod9soZtxqEa+WQjK8AVTJPOjxId2UGVMuvpOz7y/K3NmkUZdvKYoOnfaKsRGAf9O5pi5QU
DUmytPgbpVM58uXN/uLJsweV75pKxNIXpIFLnAU9x8FS9W4i5W/lL1eFBq5G7h3iilg/+SakZ5WK
rmQfFNkBm2YDjhgNcXiD1QoKCm50NC6732MUpCGpzSEd4DhaJhUg56WaJKws9sySOk9VJiAunUt+
5q9FRnXHQkVJ2i/ua2tXSynpb51Dr/QVDVHIRzEG3lTCOhcegG3cGTkSMHpY3rM8RTRDfKhfuxzg
s3J6z8wA2VZfbRNJQoSOAmspa864ITOW5jVLBdUhRm9GKtHa/gcbXaLNf+xtyBlspJS0TamxY0Ki
Gfni0cVV9qdNmr6iwmo5gxtl5L6QntRK+WQNUwS80X+PkFsXTvBcsPENi16n0lAOMaVpljIT/TTu
rvN9FoECzskHoKTaMyuk0a6PbgZtl6ChxYZmvKmwKRfLUBpt8wYZj7wd9MFKQwcpswgOeF48Adpf
oi3+jrRxo2zwfkl9i2eKdtvQQEzxC5QJ5Twbkm+/Ij/51twhPxPjqorCZ8IFhAT2nV7GuvI/PZgo
gjVGN5haxlXNlb67wVzX+xCDy3XW6qxDMUZhnQBLaBSSB8dkY6xa/0lLpn7dLmNqYzvkUFw3+H4Q
2Ryi+tlCsqORafazMTfNTi7QO6a6mGY9f6BbK9P05+JZ5Blwau+dJKrVhNi5bUmkXeLK06n3kPT4
mi+/RUVkJWGCF5HvKKw9Bcvgb9tP18hEAWxcwHEsCa0uWiUCJ/5UzsPE07MEmX+6GCR2t72mAvVd
z2HJegSxUf4yPSOO0S6A8FeejvjEON9ebOlfzaIWdO867jxXZLg9xWCjIitcshtGJnVFXpstDy23
Y3U7JredYjxhpCyuZEm2kLPLV2fsNG5TtjMfBEmh1/yFdf4JaBm9VEPF7DB0mdfG7jqPJoWCHymX
MZQ1Sq5kx2DinmmxkDDrkZhNii+iQEr6JHJZ5Z9k6wdh+0QAA5VhjhQs7F1oJAg4Zm40oqUBbPyZ
8/SXzre3K8PwWgyHmnK/YGTZ13366zOHS8+g++9AAS84sYcwD6KPFI9g3XtkUqIrpgzj3n/9+LJ5
n0x+dyYsECkwexZBV7OhMvID6UbdDlv2+q4/m0GITP6L/5ocPnqJv7l5t8Xfi22Kkx0SQRTLDSIz
+FVO2ftHP4x+CMiHrUu2LyBY2OMisAiUk0tTVKA3mvW39vC3TRxiuyEdiM7yups8aoEzYwSXj26c
7i/ZHmJxuox4/BdEajzAaajkx2UZxWvCpQkzcm/fJQz1qodP6Y9H0yrVlwEH5d4nJyz3qecfn4fb
e18Oci4Frx62Wah0ZJx2oLFrbsWfa/DA8unZKRlxdvEJ/Sdhk4wm7ohAkyiY6bba+bFRiHF3agGN
4jzpjfbojwo220ZByQeVnFf6w3gqhSJCnWU7t9me74nkR6TUzVEXhokmX89ZZASn/TAVimuRc38R
lTZCN3i3EOecDlUWp+w75KJofn1Pv4mXbPkmp1t9fXM6cdD2uH2dnAL2F2UNyTbpG8M+emcubYng
J7B/VBDsADjNWIlfULEfv3Fj6Nhg8m9pO6yufaXkGDM3UCJ6eCYpeL0pktMQfIy5i+q1aWlCu3Ck
DTUWrP6cQzUZ8+j69lKC/FjTLjDjJRTvgQ4SL8CyCkPhsQuEtmknGFdYcVnlDkTcCaPyD7ye7lsX
OgJjSR9lAPTx+fVOe2TBw5xHCfRw3ljDNC6vB07J/xvk5XcGe+uaPR9ahhV84HpSp1afgvhtdQOU
GJGGANv2OrpUerFXvR/wUL2e1KTdnNkfclXH8ke4JNxLnKvmJWRO4QYc+zXnlSoeAg60pNe0qdg2
xKxtEsixWZ/HNt2/2/x9mpsrlERytmZ8i4zdukIX7C+oOelkjKptJgIBA65jM6ERifurLd72tr/d
ya+7uoziO1Ek7lb7zxQ+8hgtws2dRbZjOFnGTGxspvFd0iCjpZijEjvs6ylVM66gHk0bXo5Zb874
LgOdqWzyuwBk985QX4XnS1sTSJ/xaXvPkIgILtxoSt4Oh6zs3hNa33Sysbh1pxt3ckEaSg1JuRps
fTCP6w84BCATXL1U+h8VKtLNYJq09dKPuTkb4bg5rrwrDaXGCK2Se4XD9HgGqrs79CakJbA2MRNu
IL/6Fn/3zP0oSKqEjCqCW+OQXgOeMEEELKDz4ZtGa3mM0uDIcUyqsXuLdR43KRfobKB641cepYAy
Tajw+T3uE9rBQZncgVys9zR7BLghAQ1x5fY3f+lkA0mTcmufuyGe4zuvzXcuXRnqq/8zcW9gPw5H
bKvw0uRYOx0tax8BJYqCyMUAAbMgOKuctidywzpGYzyOFrFYGKeNGioWMGOwTklcSHRBm9adn4HY
JN+2CXWdzNoxM/W1dj61i2wHtlsm32bwL/LdCjXSsrQsUzF2kZ06kSNOzdkaLhu3jL5cvYGMlvT+
ysatmRh6ISUTDldt8NBLFd1F2d1P2OnLIia6ZNWZygQtnpOlTX8LMycF3wvMtTg5qaziQORuM4R/
+7QrRGc65Lp2ZWCIp0PoMJ9SxUfLmGF7Pouuuu1g21x4RuFe3gv1+iI6JZwHISe1U1XMRrNuDnAJ
Nmamw3CvBuJ7QoKiNyRZEr1YbKIHuwv9unh+3vPUUG07CpjtBOyIPEtCCGK70HoVtj9HTQe9JYhG
hwmOdL7kx1ySx4CjOAxLyOJkDBVxyH4vqH8yUZD2EsYndlUWmPosmDjXFuSOPjlRBgFX7gqQE6Du
JpWhPCpaGILJPWbS60RPRQTzJbzVZXBR1egU3rIASTi6nko4kor/uGZnC+huszPkU8YzreHINC8x
Z+9yfIbIKcMCUnPLYO7E0+KBLN4bfGRt5T+Q1XL7zVggnnflUPwj0TRSMLA8jptmCIAPscD42TWc
OVYYyMWHtPznBjxnNCaQY/we3VKN1srunnsVl+c9IStT68N60csEMck/TfoxQno6g4LZzHOdpKzM
EOCgLq8FEFaNS4+MTqxwTrkAvn0AVbUl/fSkxiis5uIRAMXsBB2N3edpfr5nfbCQyNelsrZnRn/5
HxU960pN2Yw7Cbrf8vjfGUZz80cfwyFAKvRNYwPNp1dm+O/j0DSDDDOl2iuOYVOEvmLZeKEais0r
7fFGxEC7Npm6aJ6o8Z6736obrk6WpjB3v32RgY+GY52yrntWeGRFrf+ys2PElOfrkSyK1Dq2kYlD
Ul5AfCB9KsrKXAdhTtKBR/KDyHDXC208ak4uCjNRV452RNhu0GtDtgzJ+pEymCuTPwpYVQdmybNh
YwFq7CK5RsVPCJF5hbaZ70tytyLUXjoBw1C0RO8zyrFSe4k5+jTVJO1ieT2Bsx2ZZ8e/xwuWeQ/I
jCUeZUrJ7v7W40YPVIq+C/WwBAUnyp02rcm14FCnYcQOOqSoBa5sEi9z2h52C4q5OBz9pWwxrKGF
FmEbZ6qG5cAKSSH4j3UQeccn1s7P12RUF6UUomqf6/14mpmSODBhOyME3/6TBuX+6rL4uSfUCFlT
avLVAbExgISy1cLPXiKG37ZWhbyuYVL3lukdJbDr4ux6m9xoUESmHXlQOcaiVNnHhErBhCR4ppU3
xNRy93UepiFzjBxmJkpFnDzkoXTWjjuqc/vcmo4nZ8sGTBs0scFEiF3JkVy64IMWAQDg+5YajJA+
0E9it8gCBkgoHWtj71C+6Q2Z6UL2VR24MH48FYQv7n7xQct0W7rsaZdBXmgp+5gOdWNPQH4uJkxt
9/x/p7WN1UCwA7tCcE3RENqLBVwS49DjjxG8xV+a7na5VLfKATQkCAzRLUm1g4tH6oVOuRNlrzzs
57gi1HDc8bOKW+biok70cEusGlVA+rH/rsU085t719e+CNVuDGW8AjEnYxkNYOZUkwv/+9/XENNS
K7HAogvl7+6GYx66GNo/x/1osS/jN7/+AhN4nkTLpcuQGSWS2cdjbd+YxFT1rWwnDFNyoqEWJuRJ
VbrgCf+n4m5pmqHLlBagE6/zXpYFT+/GMFJHLzy+WVM0Zzl1wJjQ9w3vYPqxtZNoQ8V/0RHESnuA
nrqTom56ABzQ4bVYSyiLLzClXab0ndRsMg01dbq9lydjxgZVOMkjPo6j4ZyjH24FQGCuSDlA4dMv
I2WhJe2O5abC4yaE9/4YHhH+UHlNkGa2QpBfByH5V61YagTLRnS77yzd4ZuZoxdNoYAChE4neH9p
naI7KHixXSjveQmwfcWNqlEFJEGKPInoLNfZgC/uh+d989nUOyU0hilMaEvaGe03mXxRwQWw2IK9
y4Eg8hfC7def6wUzBhgvPrQ6TKDlN9pIxj2DM9s7hV/4olcjnBGnKKh1TUI+KE9pKWQ3z3kyp5dM
GMUhlmY5SQQw40MwXZo5mOlubr+42C86hEVgdDhclcUnBf6uMizqOui6irD2neXdu/cIAf6Bo4LL
/4/V/088MUmhO5FkEEAjPmYpAjBPI4CLNxPSdh3EdrkanFoMbhIrGwZNXm42l2IXeVSn+Sl34PKU
YfDSh446PO2vnSE6zEQi7UbPI76ORocxbUi6wvy7lXGz2tSuYIeMZhJrQ4vOpEZp75OYXdPBydbl
SWPTSUUI45Pr1ZMS3lsTl2mN3eNdScFpz4csQOZs4fhFO1Gl5PexdKF+wtzzRR4Jls3UUiJWllKe
unw3t5mGnc7Z77COxCGm9ZTjwzTkR27ydUCYXN1xuwE0fttTsTdAAI3CKE8n7+b57pkmd0/MBlr7
Uwvcwz49pGWb2Ddf38mjAfwP6raLzI7uqzyy0JYGiOFwU8qmLETGMoEG70Vp/ozH5S4VC42AJv95
sMMwCh0dfHuw8aBXdJWdindy97zYhFSo38GXG2tQs7+yfFWI8JjpX9sAVkeTK1foFzwgp8KQUSis
NGSqQMfWp+OP/Hz3qfZH/qOkkSIA/63a517dkYdzB540KM1vyafN6DYi1ML3PqYsJgZ9wv6enXK4
E7qVArXRN4beGlh6b/kGWPETHJiOoHUEkr0SHnCOdFLoo0HMxoFfw9aH4oeoQPYPQ3dMF+ZtEZ5F
OCu+vKB+439F2wL7vxVwlJRt+vw/dZs0Pr2RL30mlTVXmVAiK3hboeuEFbQqorVnLnFbIKAkKzvM
2tHDCrIFZbXA8MTLBR8MA76kgeph86CXZYOMItnta63RCHYrDBOEGffkcv7aL1Wl3EB3y+xNKqE3
QiNiEKaiahB3qSC8vRXOMw17/ZQjiCqn6FA1hdwu3zB5ewkLbfJKF910HFzPT9W/WXkov+e3pMaY
8txBIwU3QG9/n7GMhpDGDSjqTphMMaaY/MJ7hC9UbD6GsoUUON+dDlYJR1kZJcYN7pvm8nu1gBqV
MfnYa1+rClRHm65mHIhsjOOpULnQtWdcrjg38M+G4ZMqR6iiYjfSw+l8T5R0O8FTB5/TTrKxl5RF
jOF8OuW49lz2XM1pzFqi1mlcWZq76shE8pvKAOPnyXutD/Hg4T1RNzgL3WpagdN8xqH+LQVLdkvz
x6LQt0QR0jEEc68XeaTeWaPxMvtiyGWuTBH5VdItdHd3YHc9CEoddDeDaliW08OIfU79oSrsKhNH
0wMQUP2P97oCohN2gj0QVnpCFt5v82hxp3mmqZSUxxACHacFsEggPC1Cg5L+jwrw8HAPtEP7uIiK
SrdoIOTPRYdguaU1YlKi2H+GU8STEzXlmsuq5A7PCd5nhiNfOLisKhY67hzR3zdd+9ZYBPU18rxb
O/64rqPjEy4Y8TPfRg/CUE9b7HfbFeR7WolfxNHz+B8pPYdxckAHfTegcPYnttJo0dpdamuYq3jh
AT5PPEeJ023++WEFbyu6kovqxO8l8w6T7d4GpUJxVvDP5/CEtjowP8prtK/kOEioCGtBeUj/Xkde
yg4jgc8OsHVxvKp57r8M0R2gIiuwyRCcSWT5/nki7oZGyfy9VY05Rx0/2m3R9I051IrfaOnMZt0Y
XsVYbR9nAHkbtiln4AAIpwMt8SAZvKPBwPsR/r9Uqj5dmt3Hus5SWxT6OpVJ9RUZg6AUs2sODTZb
Z2tQhT+Z4GOLDlLadjwjrpl9ELMF4Ol8nFp5pAzgOS+mMbTtafQoL2zbaaqMltlUXd7eujFjjaX5
Rz3k6c8FugpIzkiYZBYmTCuu64yEZH1Bmxe/Z4mA8EjZ6FhLYgzs21OVrO1butLEHVTzUwEcceQm
qSUVFtL/cIYog1BP4eKgmHshf4O6hKDoyMY8xH8g22eTL4H1Q6L6l9hq0i98AS1ml5/NBpaT7WZx
6/DY7RDcGAfyRiVrUJ/KvSRYIc5vRymNCEeH1T5XMYzKxgJL6JAx9YJHdOelwOKPJ0/pQ3dH4Xfw
AvkXsdxMsg/G1mZlkuI2JeFi+JOcIIbT6P5IV1sk9DA9E5TFXGnoUhHpa+eWEdCrqsuNwRyerVg6
TYGo2Itl+xhr1LW/czjsLi4zNuhXtfN0WScv+sPlH/SZjaItZW4/t3xPN1jN+d0CcZtfocMFcI4e
JCs84hywvhtGfaJzH1rdPYy5CaZlSeNxeBk7iNioAmWP1JObyrJM9Ci8/r1iI2K4akXrDahFvI2z
DOzAI/Qd/ceJk77329s4OjGTtbhUd4jZz7XZBYqSu2m7Oir0iQ3Z1r3JKU0uXcLOmq2e/xAgRUYo
6jprCY6+cnCBZei0pM/mw2A/XESt2BvjaI5OQDLmEu3FekOZlFroN9Yo8uWQgyrZJGXqYUAao3Nj
Iz3qGDFUeLKW/XOJurIcJJsF6ZUbrZ9zr0MnMsZYBS5oweapxSwl+4IFX8QhRKuIhR7YHjHoTfz6
09Ewx3+7OrcUSdETDQALtTqIup+prtN82bVquK9wXomYwUwTvB+p8RnksJwaYONkzgslzlFfscrb
R5L5AoVR93S1zsSkvqZpJAZYeTPh9yJJBFE9Y3ug1gNrmd/eUx8eh/w14m31RoFlCGDL356pRf17
LR4QwMRJXVYNotmKRSWEOc9cnDJwA/91TEPD7m89FbQKRfCrBwBgNVZ9s4JIy7nnruRDC8YWDJGY
ld/UlIEau9syIfifNrnJmO0U9m+hxMB4QmueR4iy8r99a95NiGR0tJ3YAA4WJ47pJGee41tzw6Dv
enEQo6i4Y/VuSk8W01nZmU+hLv4LO9osSBs+fuq3fI6QX2Kilos2ta1D8WfijWNLPoYnZAWi22rK
uqQXDy46liJPSpNQZRpRJuckmngH4UJYVUK+6wklowGdG6ElQSIoxgi0hej4tZ86uMYzhoF3qMtY
YwieAw9J5SZkIAtksrVn8Nl442ociWJm5JDXWWiqrgYDfKEtUr8sSb6mmFR5POn9VO59cPnvLAMy
P7UMRpOL1Vsys18fZfU8NCunR6gIPodBvQXcUuwUIc+exKA5iEva8YMtHfPVHsUGP0ELpveD9kXF
PcrcB6TQyMwct/HWyOC0xr2UORkCew/usY8QChzgr9ECK1FCwv45ndvTr8gPN7EZlwDOH2ohVNyZ
0pBcVHWIuOmfD4j5QOtpcQ4KkLPFRQ4EYVkCzybf7BECnPmyV+uZOj8ihE6In1A75QKAbUGzukxE
WYVbe4dD4irntWuzgh5iDPv7N1yd4F2cG4qe1JnUFBYGhE+cYc4utVvUHLdRmxmrbVOP2kuICgvz
kzouFcUdnf2JaoD3rw8J1DG0rfYP416VX4WALPXSs8jiDg+6CMjWIjoZkqIH0dSScAjWCPUsO4sw
YEsUyOVAVuMmiFIpzaWC3AbYVaDojf75hct1gPjgd5jIb6p+fre9HmLgt4tfSBRbY0Ye0MqYmFzM
tutLNYwpOwZn3r6Lzqzoa/ExP9n6aYwT8mBq3TNvYcj38TDP2anX2iCvM6G5aVMIoD00C5CDFyqx
BtNOCwnv29XEtkAvGBibfJTUkV5adFQ3KjtojNzUQv8FNY2yIXqXjkImEPA/DpujAaVdcMQn1ZbR
9ihxpTTNYX5tha7lWpmOlFzwIBsSN9KttduCdecSadoT70v9j3JSbtueYxOUHCX6/dz6HeNZ8T8n
hrgoBQM4R0aIzn8SqYoL4beIvx7IxCRri7+OtzjbAXSd9dxAJL+8Psk4mRPFBsu2s8T3V5v51fKF
AAHkCGE1Vsd9J4MBOBb9SWx6E58G2/zduORM+S/oMUhqOQFjwGYCB0e5zGkDyqAdYN4LSEgpfXt8
CST0+NdwJv1s9jzQXzHtuDUBOr/8PT1VTrLuJQttEteYZVSs3aq1u/PDqqfkctZ8e8NBfimZ7UnJ
DT9iKz6f4DhGMmgm+KwwFuFFB7dwBwJdfjJuM9mmf7UTXRhPy6/ZSJoz1pv0iKgmiWRjFKPVB/s8
xnLwSg2qW+vxuBmXDHoKrNssd3en7MU3XkjjuPKDzY/gCvxfoxuizS1UYLM0yOgIVIqPbv3M8poD
LGr+f70J16Mk9ObaGUYx1Dl6sPptOmfJJKH3p6cotQ5xm/07AxXdxwJ4AjvBhzmb4aTMYsEhVh67
oG4yFwAHvdRT/CbLLcouIzuGTKFhRlP62BvJWLikvijft6gs1wCAJ+U0N95SXugQ7fOgdP8w473A
wQ0oer08r+xHReKwL0wsXTTaWZoKp1YmNI+bZjCN6A3WAoRG/Ro7nnFPhdulafaVdLgo/QZjtOri
5GBo3SJ6YrUT0WQkuB/757TfGVPTZYUFQsMy4EuCjdDnSXm9kwwtXOy9KxEzmxD60UeAPoMZM4MU
6Prb/xOS26FCWIRlT7m04p4b2e/Qha36F0GlDriMrnGkdwYYBINaiMCV+fCIonNKm1vGg1SsO2US
HsBGH3V7np0l+C1oir1u6tXpYHjdhCHqSpw56qBVTk3IgQSl8vvO9GBcfNUZwLixH1mWTwOXPPYt
D10leax/XyF6lXrSfM1c0BWetwbv8e9ZgjJ6yCywxoAwhhLsZDtKZZvMMWjYUBGVMDhGY7czWbop
hqFDFPnLHp3Mx21381E/w3a0A9+edRjhulB7DuizMjjq5d7hD+MDJTAhOAdJnLoQ6FtmzjsGTH/F
QXp0n1H3Xu0ab5/gsJykXkPXqZqVl8K4c8UhNNDG5f2z7N/JUogZBwOlYRXQ8wdwLbV4peQx4ldQ
IsydG2DT7eVF9aY6jkuhyE0xZfgEaU6aR9XBTuS+lUu2HMBP/rKIgKpa/5m3MKgEmNK6bCDv+sBj
q3A16a8vTmtvymbPqeJm3C2/oJtPrfyS4KxhNQM8BafmzylVE7otaTfKgVqxAJ/zsAex8LUMC0na
YiQJ3rSpohC728mZWKc3GznHwMGKKhPTdJciEABT9MswnTPSzhSnagMI0q+TQOUBBNqwils4cAQc
4zjnlE3PeMVMK75WGZToa4tbB6qepRgY4OgIa4+b9z8nDzYMUlSeClAeQrnoiknbu288tzrZFwbl
rrqYZKL9h+Joa2mOGF0+iCTHKWVDT3V6zN2wTaBMCFPJzNmBPO+zyqXtkHXrGPoCVjElzxFfexjt
hvwdgZmz19o1LZCAei+IHWrKD/Fr8ZhrJyGG9SBWVKTSYvfObKikUPK5GkhQJ8q8hz35qY03OLCG
zgzprDCKxRzDhAMG16GkMTR2nEIrSG8S9pnlcjgYG7BJyKsK0vBYSv3+EWM7qB0RnQWBrWr97nRd
XSZlvybvOszDfrK/vJx+33jDY7aoANtEfI6PQlwULGb5h6AZFWT4SzxhE1VgpSk063+omWeyhmhG
ghiearW0RKk0G9fnZGRHWwI8/C0Jb0de7XU71jvZmK3hwQwywCgSC9tt7k9wDdD2ZpBrqu3wufC9
zU8j51a4v85+9xaFEykRGppRNAcIyq4YmESLL9PSfGHDSeKL1pDxscO7ewjMRjBVP0QkzdgELtUb
DDHAVoE9a99fRDBNWthnZKv6sOPo1qRQzJ/zH3dQtVIyjk3MUC3UUUBHeC5Jac1+tnyEQ8gEQCk4
hjsExvj46hgefKXWmcC4Q4xnvt7CRwwR7HuHPr4pFM9uB0QPr29m0sfyI7/Q/8RUpELD+ZcCGuvl
x+u7+LLy9TjgNWlCqYn/C2CoGiqnqhjgzQP2PLnDK9HA8Q7GnhX4hHl6WzP1zrnyHaL/zKYXBYEr
+fkGvHZ81mN26k7+XL7fLbxU66KK40L1CMzy/W2M+fVVUpD+9Ic8piDE5t58AVEjfOffKzTVL14A
EX+4Rs9QDX2Lman1NHAvhs/MfjFj9+laolQhElhjkeTyEuQVrbmR9W7/h/6PgJDftjz7W7iapNYM
YQHMdw3X29HHrn6ZQT78eGjRq7d70ZRkMmsQfmGKg76IrPy3DSYqKpKjmJifQTyKynDHIwqjLUie
YSeb6IXOqrXjmpibWcy0+CHzForpDxIbi2oMNxE/RBWDukjWGaiz2F7bLpUsw0oj5vQQCVGrFpLt
eRYaZGXfSyfNwMI1ojQMfKkzHgUowx0Wvl1JzMV2pPCDN+brAJ4J6oem1auA1mmHjwXv+BPngLVR
HQHENrqG5yJkzLUTvMggTOrD1PXJgDZsLrNLt8toB1VFXbxlXEBdAY2O5y6M52tVyFaa5Af5YH8F
7A+o/wnPgOCGMAJBUs3rVFOfUO/y5bKP3Co7hvzL1dNJE9qgc2duGE3c+aSB4HUpYSIc6BPpbk7S
zgKR/klh/K+dj3YXqAscuichMQq8cLiFtVS1dUe7/TdtNdEkm+X1I7ofhqUapZOQTiseUlRHrglV
MPL8H9+1ZL6oPxKuh/NugRA5bBOq7KwZQtdm0BdrE01lem6UTgptldf1D8e8FAWD01ZHMqL+jAhu
OSgBbQ+dsNs85Eoh/nmCowXE6X3YEIvfLb4dZJLYdvgmhpSfIDIfqWmPMQp73deT0WgjFvp3IIGY
00sS4rpYR6zJXULPtr1P8m3Kryuup73gQdg/ktfeDUQhUWc/k3+EVndd64aLV8ba3oR+Lf3X64H5
yvxiQJYPirdiYI/kNDpiMdfl4RaAzlND9HKFSkS0Yr2nF0PFb5IRsfKjG1pM45HgbvBRHghv6kGd
Q+RLKyN3j0YWNIkxPsQNTETkxesYnDyypcLOsoQhVh/tc4IR4f1D5+NZZSWYSQEEjVRaPcOYdgzi
dJWfJvPGHSs75zNPIuDb6si9uMxj6/EVytUWV6yFF/KE4Lm5DnAti0ye9fy1lzcc0A/EA92IHFsj
aEADMWM8G5YXxnf31dvU17pDk2MkDHjy1DXIC60z9gcTgcRHb0WjK7YesPEBzTYXehQMnImLa4vT
6Mol5Fg7vP1YvbdTMKWMVCp8jRD5PUz/HyvEsIfnHgcNGkgpanPXcC1HEGbAPcSy4SNZsO2zU2KF
8S3X0+YH0jnNv4tqCnv3a5KOjWxQzepfW5EcGFjteXag9poQXCfYTSzyVI/OzlxbpSEnfcc3TycB
SvtbbA8CKXVEQTJ+1PKSC+YIBgwWbO1L1USk+qzh7q4G8sPn1m3tUveIGQ/3KBc308Zx0E2XLM55
srhNOn0JxUuzsSXUaNLA8/GTLdbcy09v10+OdqPwxwFm0abQ8IJA+c7jWIiA0Zy5loobQe3LcZLG
eEYeR07wVUZlKAE32xQ17fGgSYc6TgKJduD7r3n3foA/280ZrAUyMm5snZZAIjLjrokoukg2i+Th
LHy/I8bRol0VOj1OOw+JST9DBoi15IHIU79OFdn1QkIcp5JFuW2t11U8HSbFe+nt94iaJ8kxHgi3
jOTjWL/vYWYfJQCM39gwr2BTEbew9b6haHnOrSfhleknhPdQUqZRPS9LRXvhtUk0cEtQynwQHbYB
0Khn0K/EZvJ2vwHBxDID159F53lvCpaP7yJaGj3/hr8NJT88Z7I2kTEu2dad/qW83/MBHP+BlcmF
3BIbmg4boj2a+hnxnVQ9qir4wCThz+JHHY66UNOWZzSa84myTGKWl690jbeBgNyz406Wr65u8vvS
bKMQ0VRBRCW89uiHa45uevokCqF0b4CA3yS/P/cI+ru2EXMEWJ+fQKiE66QkYaTlvI71n88HUBTU
xkcuU42GaB93Vd1UzU2Gi+ULmUjvJUWwNZa7VKWnZZygn17Ey82HX1UTjGHk7c/DT2SnCd+rX8f7
slefSL6dVCeRno15xi0qNl2wWahoNqfYPUZF4jM4FHJdg5OzK1W8bKNYY8ppmtDpRfaeUNoSAFfj
18WwlskvWR14TtvB9oSK74pjqG5cVOBk8Znn79MLA6DZEInHu7uvxQvytDin60J5oJBo8GpBzPgk
fODR9U5Lda6/2e0USRkL8X2dbPs9BYnnKEp1y0OTdPeZ/RnTISz1VogUXYV9JWYM0hOtEi92/rjI
lzXXW57uEe5mL2yZYeeN9d6gSei6aABl0WtHrTHTCfNJz3VkHCu1FXKq8ofyOvnjLSWWrMzCRdNI
6McnP9AIpUpRNSy7VmaYjLMk9cfQxlXZYrAq0fBQURtDhSWsL2nB2wjdPNaLNFJ8bwbF2a6RP2Md
sVl9U36Y/zKrXEC9DR4BAXdRaEI/q4y9mzuFYhB1QphS0ERiV8YliyKj779T7sY0LQIBzHsSCYMS
D7gogLXRGbaMzy6awJ1tZ+0v1KAKBjKEPgoNCUGxv5uo1fX/ZAZlgy8r6UW+V6qVBo7MddmCMeGE
XhVyCSltuLIA/blYhc7mBuaw0MZO5xmjcq5DsyLh2MRaR4F3gV8MPEQ7s8zzYuljzXX9xzShpsHf
L1syjlIkdGimdhY/tyllUh7ARCv+zURAnCRKJjDr7O23DzE9lFxZvkHS5E0+jEX7cCcLKuVaYLJ/
ES4lMhJUwXqFEKiLgH2xYFg+1VLIm7dlAwyjn67fb2zz3ioHq6Diet/nFyUHrkkwoXHLc6a2M5MG
UM6Hw1FdFq1zUJtWzfTU/+JT+b8uQ50FJ71OLp69c9+Y8eUkb3h2mvlouFAYyNN64kErqWiwcOwQ
gmp9lGAd5bHpYXbLXOwZ8be+sOPANirsH+kHL2WlStTDS66wPhrwzXG8Hd7cCqcbh57ll5Um+5pA
UMC2Mj0AZmoty875MX2PYNAWEj7/pEBCMEosMwN8ZYb+XZDosWvE8K2CFAxaMLcNYog1AwK3Jska
iHs+9l+fRurg7KKGEwVZy/W0VHRTtepxvez4VnfXlZrNfN8ZJAftN3hqYfzulpNBOo12ZnbsdxqJ
zpVRC0IvqR/jqVoF7tcmC4VQx+eCJuL7iFUTC3FZwR//XVION8i50zqx9u24BXKJCQ0Oxhe1ToTE
G15zept/7tCJlJCo1WBkx020I9HkWdiNSh5fJsV4z0HRJUEMD66jkMkNTYY5QggBbfck0RHenITI
t4BUPFq0nOS/5+eUHsa0+Vx2WRrpcBVjvrn8ePHbfn7TQckPCW6dyi01ETxanPBV4Tli3OabCo9G
Z6x5EWNjIIVLyGD6fd7QEB74p2ucvcz4y6JqIs39G2e4SabOvOWMkAcDI62PCrapDL+TNfloJFoz
J0R6ga1OqAcMgQsJnQRXCRD8rss9r7l+mPC0bssezUNBB+9H8dtDk1A5iG0ZfrgS/plShYDcr7Ye
9ieyJGAytZ/iyHODHVHnyMLsffnfHWeH4YZmC72tbhZbycsXxQj1r+WuqEPcHK2eH58E2NVTRlNX
5KR7E+MNrQwT7EQRFZGmNXcjaWaWybSjMJCxxXRu2uYCkni2DlNYJRT33ouj3w4Ofd7OBPec0ZS1
7xhsrXVbhkJad9Et/TH0HQkP7WvbvCyTZr6RXJkIN2PPe7v1JfoF7qyV8oi2JXBLaCIeenuFQFQO
XPRuu+DlWVGrdp7t4R13qj3NgqZHVNwjS0rQBFbet/zdsP4izJVDTrQVFUkvkoeXaacSnHMQlC9R
Qy2DMiHDVqba3jdpEmTeDNYe/789V1yBpjTnALf8yMkNiMhvGF/xQbgWhpObjpKB/WHkFsSrDBHI
TTMqL7GWzsOL49YK6le4ahCV9G1jfePFJEyruBd/MPj17JV86xieuJtifU8DKPjifVsS69hwZ/Sk
7xyDbfo2lXIwcYn5diS8dkLM8R7Yo1/armDrbOVZiZ3rW5AacVPIL3KPPYo+Apcgzr4WwHplIOp5
7Xjak614pz76gQU2aBEuxyKVz9dByDYDTIQrusM0O5tPWdCfZe/8Z6daRGAmRnaCTEnKKMsyr+/n
trrQ/BcMKsfDRNmoXmn3ehhVC2LIXZhOWvHSOBMO9x17kdPzgvJ3BRg/doU0VOQiGGnGJfm60cF+
rH8S1dKmWoChr255zmUfEaAfB04xR2GnP+Zn/5o9wr3BoEyhf968Hy95dwGoSRNoM702b18u0qY/
XbsCXqBgMW4f7DJJ0/XwKp+8rh36Cvuw2ulnptPg5MWAgUCUtYENJ31VVy72mzhbrM9e6Ezo3TUa
lPoll85g7F5u7cqKCRaMTbk5RFeypu4bRd2THweN4/XiqtPqGrLp8sK7yf8818OYIRtvnue0jBMo
sxHVE0DVN7+gFx/YnLM6g8DZFkBiivSqV1vJaK15QHxv0rG1U6YxBszFofszmlkUZjDRhf/+q6Yg
Ti+M2DjLRraVXbiV7g6L1z8xERQvkJkTW+pZ/451JJJ1n5LXWHlYv8+soiRCMa5TIcBU9oWwjqZU
1NRzycX9LARnCDUoSJAwqC5qSLcSgsS0itUQD4yz8E4HMxzMbt8tpdWgdzX2k9ztJw8IBfGVICk6
k2FvWobBxjbpO9oAUL/qZ5kz+46/NYJpBk0+GYm0xoBzG5Zex6VrqbY/DXghPSQAGi5+7SU4bhfW
VCm7ECJehmyCYIX94a8/OI+1qlkBF2mY6SlW0GEWwJAGjY+SmGF7Trn1L1v5i55DWI5cJCYtaX3d
Hf4Kw7RPywu7+sz1+HCYkoPMZEr16pAge/mDUXdU+V+B2Aq1NYn6ulmlqUejQAZHrlHZvmx1Y1WQ
acHWNo5/1LqsvLlJpEZyOxFdE0IdkN1lX+FOoRRBak15lrFhVzIsG6nF1pQIjhoc47BQJob25DXq
25N6fVZ5yU/mpOlBYEdZNqOGfvPePkKMFpUtmoxwj7y/YGGWPOS2RbTFaRSEbycd2g2pRUnAya5M
PDCEWstHCEi3hXu6RfHBcNCOlSqus379XbMLN6Oucb/cXROuqJYhoct0aMhEP6TGPVQhWV1waqk2
PIoVoc6ko0ajwDhdgnRbLfAA/IgFcP+HZk5+mYCkTRluU4o7H8FRcHRYgTfKfcKHJbQVZBM16USC
5wWNepAkDw32V9KdrQIoBNCkJwAKXgpmIhANFClyazZsav38fy1uGCbGzBPGgapTV9/EBtLmkOp3
yuTaDxSybaHcL2HkF9VOXoQMy3snVMjPGlRS9usowTpOtaR6UP5UYJqRFr9BPdpi3LjctPHYyrc3
CJHnvNFCGXWd9s56m1HIEHq55ZA4yuM7zZVGqdrXhVwms0hVfDnnHHh5LwmIthpq76dWshxeTV7n
YBG4A8jgSzXspB1Xp75dxspYOHzkY8INg0zyNYVSvTd4fsv9To7Uehx3loRUmkl4lpysBivg79Mj
ADn10hj61nsWX53DNdZ7lb8F8hCkeU8mDqJ0UQ0AL5xCW9hfPSc2SrtezmuibNAiq+zTx6dGfgOC
bZmKkmQAQvhpsIJDOsH+mKoIRSN2E6+7gpeRWuAr5GY+f3QuHbXoKBoPJ9qUOxaopUPDfhquxNED
nYS4pO9ijh4+PQDQsFZAMHfTwJ/ZH+qVcnN+y+u/KcweAM3P6MCg+VdTQlbIJIas9bQUkQ/li84m
3mcdNO1lJR5B/8mwwXdE5T5B3ZwgOsWpADMZ7yO7qhK+hYkdRDmZih+wrWpFFgN73RTuAPTpgX38
8uWv35CzPXSpajaWrYfd0SggejxdTYLucezpfTQX3e+h6yTzxVgDt395vNYQ79oEDizNMHtWDB5d
c2KWDCcL+qHw1+QiLAZiMzOE3BZwxrA8aXVPYKK7BWw3AOEPQTY73dc8cLc46kurXM4vSVN/lEoG
aKAZujj7Q5LFMbCYKkktZ5vi9RVScZ9/6rVP9DxU8i2DUpVjCSCh5oLCE17nCfXYmgZkPFAzSA5F
YghnQvcxRFjn8Hk3+HALR9+1oWIwZUSQVLXpllTehNFIKdWeKWwHK4Z0Jzk/QZSJsROgg5ShvnKS
+SDM34mWz/7N8+6empjx9pdoVFxMw0pF4AyQN9+zpy+p76bl8UqSoEloMVEN8NT+/i7p2xSkR9s6
d29dqjkcJm+i0DXei4Ns9SzK3/7tEBfD1B69pvl0s6/mwFqzea7N/dcMHoWSCIkeOrxTc+UGqgtQ
vWYY4zRer+Gyy6NvRThRR5TzJbffZw7wGVa/cGZ5HKbt9R/9x3hiz30PybR4ZAYObyz09ippA31M
AItoaxfw6dO5dcN2zGRg9S96pnfrl5nh5XTVPXi0jEglqiymtrV7LyBT23dLcQIp6M7Av9V1iAfT
A1y++lt+0d/2lMjQQURgC+JshDkEi5HymNG0l2Pk6bV4yj8C+debAIkaSARx43p7+W3ghsqacAWk
AoiYtIsahWVJNYlBY+27nBOSqhgj4luOll9WN3idTB18T+BRzA2F+8cjwPSykuMBWZ8iPdEw893X
HAIuPhf7F2XtxiD1Nzio+Q+Z+Sh+QvvHpG/JqAdnQcAqICtdM9JpCXLXaTgE2yRdwoGVLowpSdHY
PbBpCgkhWSMD2ufoZIh81j/qmmDM+VpGRAqqEsO91VwZSERvWp8ycA1Eao4wOEGqjFXgACgmG4QM
RQv/tFtK222DTeCVs4o1foEMPRDNzXpCj7nB76UPmZ9sif0o1ufeltJLTQ8UyQdMv7gk1p3OYq0B
Fhnj9ALgVvqQVdJBVTGx+CuzGIJEwViQnGL3yhrj73xpCzk4qnayc2joJmp2fETio6swVOBaE6Ut
nwQxzcsV00In7FKoMBCsKEwcxowvw9tcXA6fD5lpXPIuKopbMD3KSlEP/yI8TjwZZqcAU4wcK6O+
3AtJCeLxQ/RsKDb4HNsnMXbT+70S+19RuzdbQITxl08UzxEu0Cj3zR9UHdVOnjy0DGYSc4YTNo50
U7iaA0m9Jc2z6+MqVNrQsBTnjL0KJJ+10UVLPnO7RbXJ7XWHRPyE/eTnIClx4JDCRnlJrafw4806
YQyP1mAT04FuS22mDIAXksKKEUMiDA+OMWHQQ2seoq2hbHmTQ0oqP0CA+vtIWy882hybrqlZNLUn
pTeotoaZ3o5Nxcq5gKPFZ99NLXQSxj6jovOpjRPcd1iwPvaFC37ABEXkylXim+rdvN+KfG7ufh3J
TV1c4P/3buFp1p3agps0oxOln7k+Y43EPLxd5/HTjvHkFP3ntqWxOI/gRGjsbVnyON8zw7DGkOjK
GNgctcC1pKVHbvtQ2zWQFO5KZLRB0Af6ZjZq5+al77KsiuNKhPVs/6wsJouJoh5RQ214ILtaA3zw
Tj/neN5RhfoQgETGxumUI14DLvaEWduSVDG7/qxLOA09ssZrX4mqryTbSVXdRbfXPjg7WIckeFLp
+uqs1uWOF2+ylZ6GHVQYhGJ8S1SwDTFdxkQtJCtRskL1F0w07wjwDxzb1fjZ/3cNRcSinflfXSf1
kIpYiV2meGBBpNM+1UyNdYNvizFscDprt/rAHZwQ+mlNbg+2zByO6YoYvbXPh4RnQ1krWosicCH4
NgDsK138lLb3h8hnWsp7w/H5KM97LM9NdTkZrDNkUE/YDjjMTofWgDGUdhRiC+wAZsrY/wpmyat4
1v9Zr40EpCCkBlAxU3V6zh1aiJpK1U/qUpV6kEjVC83WVcrm+UgllcYz075XQXsJJE7hcM8uTf+w
H5uscYlnvzFF+L3gqaYobcwPJq5SGhqi6LVaMy9HuTGZFx64FONGpt+TXWAu3w76LsEUr8E8FfFy
un3Ec6rq499i3m9JF49MVV5W6Wy1d21wqeYHoMmHDzzEthNjRQui8u2blHZm6ps3ZPy3QW03UJmC
v99/NAQLYdnJZ0sFwPZKMfP8iySBDCa/HA3vvFUsP9K6jHpkxO4zy3EhlIJUdsisGP5K+3N3NKQK
A+zkU2/gdvoQXAIGfK43BYSjN4D2iHPbycGO/MVl04QxZ8a9HkRwE58uAIvda9Y8pOaYZ5XedlIq
haf6k0IjftrK3wlTiXCr3m/jdMwXMkRIH52YbvmokMMHZ4x54zCo8y+RzDaGm5V4UCg34bCDaac1
LTlkH4MRD+szDJsVUPCgc4KciVT8lTjQobsh5mzIl6OB7dQ/4j0QIKrrR7/G5/blFF0U9f9050Ia
eoywBdwf0nJNhaV1qgcxIbDPAngR4ueRBwYjSAcf8Q2T5rjG5QpySDtBi7CcIV/UYhrwF4rf7vCH
LxbwOD1PyEUsaEP9VLupULv6HFz+m2Oyr5RkydF89E6+H9gbFlOmWHuG+6utku5m3mYKx3HQ463L
Y6upmxyNFfZnGJxRvAEXMRyNHeNDYvuz4O1/+Z1EyZsWa35pXwBdsbju120a/5W4eUopVrj2H07z
+7RCQiNs9dLkWLCLsIubcEoSkag07QPHP622kaxgoAQjWnHNsUFto6tEh4bwtTxUkg4dfuCIZj7M
vWgNqYCmS4Kh0r7nNhXpfvC9rbQGsqtoXyFMpd9T/Ej60lKL8KyPz+TPUg7V1p6ojCDDIrlV7Rn+
nxwBoXxGCsKtP+zuiu90HNNf27EkJWe1ZlYnH5cTmTO0sRLDv82v48HQ7Usjeey5CDkG9IVhT3LX
jaySMYmHzdW9dpX91urgIdljJll8/BOthEx2WKISDHb8Wlh+Q4/9LzIZ2SclI3BrCxd8LU6ZszlE
ifKN9VdUvNVv3m1PH7/irtfHYQDD5ERevV3uiiMuIJ8ERxfq8Kl7hE+Ig9m6XIHkpbFQ/z3VtoX8
LvfRM2s7D+hyN/ls11x1JhZ7ePf7Jnnva2e7b3Atl79/1HxrEzuzwZBuqdbbBjNsMGrNPnoMuWHZ
5CJhMfWT0XbVN3N2DNdBOXyMAQWdpt8A2FXG/CRYNy0gLdGVwk0Z8WzRc7zWDyNZDMc4iQ4+v6aK
49sqQqNyzaT/Xoiy893kwIGLNnULXF+MGOQmN0Y9DlcFXYXuO+jB0ToYVxc+/KF/5X5Ilr3PWjH0
92vBqMLNpM4VeWj/6LyVZjvDJCjMvjtDiLuxeEFndqSVYirMcv07n6HCtO8iQvW6q+7vZT/auvN4
H8uAyY8PZzlpzaqjLAEYd2sI+suhbLYmYyAmpTMcySgtopjqMqB9QLedjvi3Wwr50MTMngmOlL82
rnPE1dRjxSYHa9MjnDdnlAIxy78vzBpcMaV0ysIDNNM8I32Slhvsa4PGyX38ay6a2nxSGA6nB8em
CQaeyETfrPzoc2LxEVUkf4CXfKsl2FnT2nvhZrofRvFkL1nq/Wr6XLhDEK5s3Sytfo88IzcTF0dP
kTNkk1r9oO8W3j2Yhk3iA8Yv/wdeEfaqHGGFjSAjl7mCEnBuwIn0Clpm52Ue63uahZojtlzCcQJV
O1twnKZ0ycghQw/vtMUf1QdMFR0dNDUXUFy2nEOCHdoqgFlBar0kMAjBSW7ZmNHkVetRDWyB0mkT
NhmrmLr16SixB0RkFtIMEmaLPBGDINrkOT6z1xOOGimEzajP89/W67C26Sfix0ZrS25kzgzl2QT6
lQLyOhA8UzwBpGcqbcbsSfr5aW/nyhEgcqMrRuO7Q8I6JjSPOZ+WjvMk4JQTw9LCNj1E+0Bl41GA
FtQaZMlWhyMB2JB5yJTEV0lr5uk7P+yWJkj13n2yq90WOGzPowqOqEaEk+AcwR57F/TMUMLv+nig
Np+keNQyB3lnGeIEnc3pMkY2nqJVOUZxvDNYlXvXcstVYONYrF5E3/XzoUKHwRWf+x7w9VM0R6Qt
ypWZxs4cEutx/6WmKrP6bSY59DrIml2CDKmHXnDSaJ5Gc4mhwlLbXO/Iy08GuTGWRXiHPx2JW3i4
te+TRp8j2vCS9x3SmTerpFBj7amQkpwyH3ehsuSZkT4muUtp/moyVgKsFdEwcjg6i7bdtsAS3I98
gCi5wq2K/lksxeYYfIPnd0M06OSH2GkLp9Zc2DZXAJqAaxAoV3ejW5Vm7PLY0UG8pbTXI6mJtcnE
Qb8HwkY6nhg7Ww5rBST3oT7tdIDJninD10G7kPxpwId6PuOwxfbtStyB8snd56q+XxBMSDXf2XXv
LAc++PCy90UIIN3Z/+ca6xydoXuedXYmCK1iAvuVMqBGthck/vw5tw8uNXpk8qXTuXiC7p+9cJg6
69YAU8uRs+gxxHICek2bRt6w7g+SGdzi0fVYuyiBr78Z/2R0KJKBF+9uIZ0sdZ7Fos9HhCGtJhta
fEq74guYULgA6bu1NV+H6HUjKXQPstHVls4lSZOZmHmNjWGkhQ56ZUN+t5wMropM8VZfWB6JF2vA
r2ssx7Bveok3syjihsVVFvMckrIEaeTo2m4YmnoHuvqdcMuOoXsgJspAwIRY/zPdBCbVjCloEP/s
YBOMAElvAjqBIJ5B5/tuJiaSaT6pyGa6aTEPEauwPSNhMTMh8z8n7tShoB1jbsP600A6egZf+x/O
/C1jTgtFfzEFvjA38EdblLvYwS+vQHs2Lpy9DrRsu9V74dRl4BOPp7l1zb7d9c26dh3/g4A2LlGV
fqHtHiYQCLRPc312uSKsqe6xAAlCygscR/XxwiDjTa5SQia+Qjsvkan62fT1DhL6oTcv1MEJ1jYw
1pKVlkniuk15GEGu9mAR2qXGjf2F3OMiYvifHGw9/VV9xSOAuP07uqxXhtpzr8oPsNqHHdUKyKpJ
t6YBBKh2fCDWUFVEAc8JBCQpnekM+fTYl93CoFZahusqRZ9WNi6go1n0lBkDCw1lJY9D8B4UOYv8
HAnTCWA/ER3wsjPes5ZhL8s83KuTb55dTHRwpYYATrUjF6ZZ2hIwgaEKBCJ+VL9sA8maLSXkPi5k
+YsvgXNjJ4GYYMd1QC3ZT9uRKwGAIT6XUvCWHn0Au+Pn6ZadhX/SRCW4p65Fjcgqp+4b42TMcf0r
ZLJOx43xpt+DLHuEmyu6coLlzK7pFhkAXSX2rdsvAFNZuxkITj+t1pdRCv/v39gbXPyXFpdzd/y9
N3TAMb3vctksEUpPcsF0w5HhrV2/QwCzy1DPCd4xsEZfTowKuSp87sLDrBdneq/uvtflTDB5TVwQ
kEyvSPBwNXUQQtBVLNP2LbeiKFBLEIuNCQQGam/3lidwKP1ZIVa9U5xNiKLsFMqmHPqga3x/WWgC
j/A7GRlFWGvN8D02BlBqB75Ufn4E8GJgtD/h34ETn82Z/SGyk5fTv2ni5zsCrgY7+ovbRZimTmtN
nGW0d3tXWI6cW6njsKKBBySzuqk9LKQcktyTehpput4ey6+OgLWMhxsWS/iVVVaytbby8pstxTKA
nk/M/NUyllGOo9lHpl+EtFQoqJOIIfFtXs/qzR4wU/o3CtsyXFjJ8qNp5M7IMVM4t9GlK6Udz3lt
4NdwrVYUyrWvZ6p7qIPQJzfOsV3jr0go7wHTpj2p7+qaNqxo2jujH7PKyl9poqB0bH9RwdWEVQVL
yCMl6cAW6l86lgcNTIgMqOCsZF6ogohePdEmRcl+U9uKQXqaI5uRTmOblOa1U3nDr7zeizboTURy
wtvF4p5+vRNdO2fQOX6pkm7VV6d6U2DsC/LYgphxYoQt+ZFtzz+l1G9YJ2onEI9bJXbW+1gjheHZ
Y2rPRGiwS7tt4OGvSMSCq1Z7vVL04qNlFvKWPEXU8NxFAmPB2tnlTh2ofT0bmnJwancK7Ra+0YX5
H+WSTS1NkJsCa0vrnJQ9/YQZy5x25hkHVJ7RXI8c5v6Yv+tmJkVkyVyUK9Ww+VPR6mk8vVl/0w1+
Rc6KgN6yd2J5eOBgZzkPcEJtO5RpVsgW5OuJtJMXByKSZ4k55M9LpyQArl5aa6070YhXEiLdeL7K
kuPDbFPkOM7QGYTS8sLhbpiZTdKiyn8ML9PeUKUIPy747OAJUt/pbb4wKkmS/nP5Zqwms+rM3eFG
lSp5DofnRF/XcXsdkbk6zfc09gkFDKXp+RhnfOzyxXEvuBvetf+VGFtfkY2o1HAwQX1/r5oHqZC2
bq2Snrj4xvCaukfMjun0EcZSbNPJxmhm3E5nMJ4vxfR12J/L+s0E5dDzG/8Uj18brHKd569dekPZ
ckvO4fpNTt5p3om+h+EVaMgk4ICvakcKqZ8TZ7/82W2bbq0aG8xPZIKd/E81Ffsu908OXCzgZxE+
CvCESoZeoNe2CWtXtPjHTcgKw0tPiNx+CEIfEbx9dRLAosXHkivl75jTyPbpFXJzPWjkM00vPQLK
3kQBLurJcrGu93FGJOajuZIVO+ghR5W7V8sbakMPzbiEqNYuebmITBrD9HZUUgJpJ26SVvjXIaDZ
GHAvxbIF/QemHFgVdSFpMHE2XqD/ZWaDmSyWHPzYarzwPb3QghMRHn272GZ02vrUjlcN6hHvZLAQ
Sbme+0TeFJnV11B2YvEG5pAs0x/tu+/4LTV5SoYdtlHKqy93BuPlH8LTe2A8XOPKpW+pk6A+CLe0
/cDoXhiTc3QzD0KtpSxujNVzc6d6nIcmkOVl2NuunfL3KRXxsw9bKTOJGU7qiElOvSSbGgWwscp1
diqVj9Vx6JXeUdbAKOG4dSFf3/R+Jh1sdzwkmNlDm0fjV73+GXslqDYBXEsHrtlGAQQuiIF8BtO+
xSmQprESKTuxXtwEmtx0hf+5T4sSjHcN88rjADXWBYCBWZnE94sn15NOqMd4Gf8RDZmEzYPjxaZd
zWTHJt+jDNWSeQIA3VuV9czTqMlXspUXxZbnak60o/0avGlmOTztU0AwQvKsZsY8egW89YTrwljB
z64YBAMKFnAOi3UvpkjzLdzhn6denJ1hsB2cDdNqIc6U0c4vFsYfF3xI0+vqw6bNdjAHlzxjB/Vo
0rQy+7spki8UgMg2J5GFYob7C8xKe1JqxqNmqE0AviwLjQBK8vc6Kpxny+t7dlx/JJDsbgwa2cOG
D0VWvgR6u/x2ADiObpwMYIdLfS8YuaNeeC6v7vOWPR08HUBO83/KFrMNZjabFwWAc4aj8BiOKuj1
blusYFw5hTc3sresy3VhDhFxNm4q3W4WbM/2UZ3kMbH/8UNrmLerWiR2TU9odM9n4QQZrXljh6nX
nOX5v2r81NOE/qNqN0veJfREyfJgt5Of9Mujtm7fUE3P+S1XmbQK7Ry7CQIez6aiZ4fBEKy7J4Dw
rw0ugIB6+TG93DtJR/rwtIwnH63b8NfSu6/8SMPgpuke/21bhpwBnALghXgKFcndk0MMeQ0VFDgC
I3SW+h2sJFpfx9q05rRRVVlsJgWlBbng0jpokPotZQVVpa6GawIJcuIAZhszfzl0sM/NjUxj8eJr
qgel/ReNdO3xQ81PbLTf6YkdRsi5dM7TWWZHIMvCfkC8kg/bdKXbiFrTDgIB99s9+8CLy2e87K4V
AgGHTelTXJCtil5tp3zowg88gcCkI/WBa3ZpVFKE5pvpY6rWkovsViCRjADBJeN6YwtKbbN3geJG
Lxsf1SCCEagMC/VjgLI+CgYrp0rhoY5wrJGMt5X0S5wwprXxRRIeegwBPsZxLsH6NqADno6mD3WQ
LE0H8Knw7wipUd1mqhElD43M1fhlL0LLDDy4iDuPG/dJMFS+fVX4WA/5cy2pdMPkL9HDiaG5cjjQ
SbDQp5vrBXqBkQkeJvxIN6bU++Nbz7B6BiUvpf1mm9Fp5EMhu4szVYtmo9Oys9Vr25fqxA4AbAtm
Xk3GQssBH2NfcmysJrOKFtLs2NEn+hr/+7O7QTBlRqNbJvh4GTmD53sCmPj2zyBq7kMA2kC4CUsp
44eO88qgYtvLqP6g6fbd/nKp9W4Z9rD6AL/GSWYNXs9nAMO8WLaMI+nVBIEpHK05pYH/BcTwjlN5
CxitFYHlkT/hSp2TQu4bgHsXKiGyjWYsa1YjgoyscPBOHaIgpN3C+c+/ybMzOe8sPSzo+xtrpQbH
Bdl3IsljSc07vI1gnQvnnIORaghkMGmswZFFcEYGQbLpUvQZirak9kd2cA4lvr2FVe29GjCK+Ilk
EHkrsRRCbq8kEnM2bL4w+PIV66phjBJgrVBt0VwsOV3ddh6mKz36C8uCw3xMqO9UAhAWQDrEySrW
oUuH3UkhAVI9QrH9+gDtX/O/lKthgaFwTQ9T/Tmprr+LKzec9+GyPUzr1mZ3LrXvaK0iNnaucB/T
G3AyHK8CSff4hKxJkW8AQxOus79VR42RqBlDmfDBhivwHwj+ubIPCkDh/b0FCW1jSg98HQpYA/Cc
kH9zKASd42iEqB47g2DgC/lszSQHY3U2hsJvjPWsAhECyRqPJ38hZunSD0NpmAtfNW5G3SoE1rnx
MKGPVugSw70gZaOzWYCEGCVLAFIUKxrlW22NGLdsqWAAgQQg1+4KdosnCo0dG/FqlHeev8lJ8x6f
QOQmG4bNvDMJLywJ11sqXQWRWBYfyqEMVH0b2rC5rWsoNCIXDwfzZ1msfCsLexLvYBTN07CHWu0O
Nx7cE4yQFEgs8RRTAobK4xdR0vttr/NkxWPAaceNU73LB3nrCkOidei4OiiQXTf7lyPf2wkoFt6b
5IGBSsDGCMeJCrIZKTuELagJXQ/ZBNpOow1RMsy6yo49ixptHc3ezOPDwQGMoTGYeCUYCd0RIU+F
rvcroCjyH4AQZMtF9KbrxTRQPz3b0nDvUvcqL5XEDv05xBfWFjS8Xpw95bMJ12SXtvmjbtEaWooy
LHzQWFNaPuRs9GsVI4a3g+JKZ2TJ/S2A/6KnikwImH7WdAeZOJsLggwyjeDmcBknl3m27f9xSgrA
7LcumqyH2ZHygidhWstg1z1bv3z4p2wK6LxoA740OrtUWRCdOt+JrCtoP/PV2DYkGlWUvjIgWI/R
k/Or4+oSPmIEzR3lNP+F6UstzLfeH2KjwnXt+UvQYWaohMKyiscVsfTnOh91Afi6UQmtW5pdWteo
WV3rJzFqgRacyXAV7pGXeOHF+6IJj3nOCsZR7KAR0O1o0kYmqo1dtZgrjv6+pRMON77IOPbRTGXQ
UNxe5mkOzc9vq/+qnIyVR9jG0I2AKuWcV2fmdKh4ZoI9JJoiNFq7r89//nz+2Lx+KZt4dL4SVxzk
vRAWNIuiZDhyEt1ZoUpcnyXTC68EgcR4RJsfMA+MEP1L1pc0Ot5zkMJfCfjwj7JivuB0pkDE1q9p
mqYRC9YZ8qX75d3YRTSVef6S/8ROJUoadxrSnjo7CULLi9TaK9xzq4sR8F5Tl24tQt4+uuL9mGZc
um95fetUZjDVqAdbPMTMlh0ffswEymdF3icxVV+47heMaVR9DvCwgJ1bOp8r2ffiKlV1hhWJCmCw
P9fPVKtfXiosQHHpYMyypZgke8oer3MhJ6CbremYM1zCmBtEBVoc3VYs+i2K9CJ/Q82LkuUDRtUf
eZq7LVjOpRT/pAOKwlPdBH0RrL/dFgaq0Ir4SNK4fKtBlsEOIctuWnsMww9hemmS6dRSh0gpak4l
09mCQg+3INhDHhrbo28kOz/ignY8ETN/WiF1ol4/fl++1CmoaHPZ70QTjK88yOBaZeAkC6MUPmau
Nk61my4EVujAJB7w1sfwzbLsyY+1tiO9NxUeayJ8DJrH3RmLEHoTLJQi5Q4k63/612fi/Zv3zyhO
5SZWfv65FKC9jvYRGDIY7jiv1ouPor7R4tQcG+N3a/XFHJkokAqyKqbo9WkfLwdry3RMBk0deYVm
UEQNpMJ9ouA6dOzl0Mu/H3qyw+ccplNLCuJhMDZh2One3msYrUg56F/BL05s6WxNdDsk73t0ug7l
StdVzRRJLXipZJS6swZX6/VzIUlDCeUjEsu+AUOuACu1pGKj79hBnVfYhZhh4XSXSc0y6RnD5rJg
mXFmmxUQKKz/mAWtBP1geVXFXcdsccqMuaBPfL6Xr/j6cY/r+tiSD7l86YxxdSYQKQxDuWfgI59G
M2HONnNrq8YMLT8y7cuwNVYHkua876SQbJnmeuJDc91+nc0QKHv1arWy3sj30YOFfZ5kNgqxPzOY
HQ8TUDNwnRTN8VnSdo29c1GxFSLaucGvQ9m4Yu4nIrYo1wPom9v7SUY+k7FjBcjO2OC/E8ih9+3j
p0B8R+drLJ+Y4rP82y/SkOVCYRXq/qEz7mNLPPRPb9wDtz5uLj1ulWDUPdNcOlqpPBaIOLgnh7gD
xRkreZAy4u0m8zsVFycH+YLXLbH2EY1vyej1sxgRNzZg1UonUsoJNM48V98TNdkp4Mi+seFXV+38
1WPu0m3QNM1K6AW6eSnyncsX6Mn8pNBcdMWUvTZ4NuMr9YHj4VPDJvaMTMeUnvmXLpj0VXvV+XmW
3rWbQhaEzhlyykicssV1gipRts1117rtENRgrgMEjfkEOcem4xeWFJ9A0vRNPhjq9KqULVRtv854
9xx7p1V4pBSKL/X2o3uq0yGPtXDy8htVXzSj8brVhmZO0MmE8Q8MCAEO5ifixhLXWa9nEImxl+j1
hPhGatBxLwuHLf+DkizFgjptRhd+tCPWXPMCsydAGukMXd+MR4X9q1KweejXSyRfb9PQQbTMoDyi
IbIxpT+EdwWvZSloAkmyqBwckDCIyZUiK4h+BEsrGmQMe74SzrpFOasAyM5FOCX4nuZ0XVKhrPOZ
yyNRwepWlaX5UXHvLAmn/c4MRdvnxfdZPtM2CdFpkXVDWP0ybiNBXyTH8X49fVgsSetXEg4mP2Lm
cPGa+E8sim+jmycwXawGNudn1Q1Iy9SSKNSy0kLSHX2QTPQRfPShFSlNpLHllMDih8wm6HmutEOi
yX3D+KizZVo4/RU5ro8xjVjN68/1jfcbEwlMhtHJJF3AyIFxHXEEgWZDKnVpqhL4RH7Chn7N82iQ
xPnTqVdG9RaLjqDTbXAlp67+kutrwBxYH9YwFStknpWSR4cPVIcM9QtNjzzOVKUFg3rzBZEVQKnO
vYMzVW3I9ZBnKc4alOYAxX2j/8xMQAuU7Qm/xXclDE1OAAF84qOoOXKq6DJaJW9XRQXDfo77Vc8H
jNowTZj+6p3w6oUhhixKYZVDIsWHM2cy2gcVINNU/y7PqRQlb+vg1A1gC0Ab+rY8Cal2gned47KM
F3pQ9whJOaawkIAHfL0+Vx6MQpp6jOW8ur9Tj21CzEfU/d0nk3CT5btwAalgxevy90eDyV5yCv7W
ZLhCpbbZxZBWGjF5+YoLEHUkN6C+MiuoKmgUkgLjplAAetkwWWLDYfhxl1zhXFDg1UyQuqhZW2n7
nScWfIeYtblGTmfbKhLssYBt8F6YfMMIp59FiLVX9xalgXdS73aUuGi098XcQR6mS5Q76OxegQr3
Igd/42cF53ujvwXeLHvL9K4mXSOpJm6kp67EoFMiI27b1+DEgYvbwl33Ab7izVOKYESGGUl/1tyY
2o0G0Z550aEJpNnLnp6HtBUVYFneJZbyoBX3Gabqi9gVhXTIqVVJvbcyYiGEsfHZDDJT7qknDhCI
9fbupTrhuxOIrnJAupRTxa0I2abn7c/moPnvCyyOPsa8Qzocv0zOX6tTKP5HuX4sVVIok5119uSt
uY96Ld0Dmn0nXA5qxNuEY+ItIFW+G6FVKqEZKvGa21Xh3KkV8cPfQtr18buhOMmLDX6SK5TfXRQZ
wB0V0aIyTeQIN1YkcPO8H2++XtNcq0CZH6Q4sHgY2dgb1Uu2GmYMqq8Ksi9/myb6NzkfufE8tDmF
iCtuwMHieAGJwoeFn8fp0MnfoQtU+W8vIANwEIqqshGBDeVUB5mtdRszqHmbY4vBU+KODinNT0Nm
CvQH/3yHcUjYcOKQiiSlVNtKHNzaXozAdEpIDyHvdAf1p0qyCQiPmZRfDCwCaArz1npbeNE+MQ70
rHn+BjnGnLHecz9dYGmS3pDjNYqnDHyx6Orok5j8sHPr91st/rs22jdD9lyDMWGQJ0JFEAm3yL33
l9fua7RD74AqyNVXTsuUSnECVrTbo3/aUtB3hWAPCFES5R94zDdlntGiygI9tVVlZHvztbasxj5r
S99pKndAmnqQqm6fGh5PSyGUblpESxgKMDGIB0K7bZHjV9olZYLuUyKbzYGbllWt/aY+MafoPP/X
VOpluv+SRgv7icoFLofLaCBqXt35QmSOQ30ivD+Uc3YjWhLnNs0+snn6Nmhq+NLG+O2cB1FkRQyd
sg2W/y8jOjqsgovaeqtl1T/MxTVekVQ612JDXzZuPqpYwZIOUlIfC0scBKBcy1i1pNuC5eLkbMm1
4OA+2cclPzfxQNCw9mpcTJlEgAxxsYGWQ67Eek69Lpi8WwwXbd5KEbCKmAK2OPykSt3RdJpa8FWF
6dx1pqU8clCFx3bht0AJGK8pyveaTr2ZOslkBXqGRtSuVvLK6/Ti1yLPlkhSRwlWUNRA3SnZ7Abs
5taedzynCxlk8JwIEHhuCZhor8zGm1fuqoHMnTXY6yjJ4pgmbztPJQ+ezzXvm9CLf8lDsKlvw8Zf
Aw2t+C65wcp5xQU+iOtpMFG7aSuLxPJZlBDd5HlqsQzm7aGsSq7mNZvEspLXZBSXveQTPqEzUlG2
aufUN6FlSpQQL5xs73zzRyL63zj4XGpAskH1jVGEk2Jxu4G0Qeb/m8CWD71JNVCqiMYTLY9U6U4u
2StxmW3KRo3CH2cD/zNVaJqveYeNEz3URV7SO6bCBzdZ1KM8+pTq2S1Wc29u1NLdg+W7RTTSwuZ0
myKfMrcrEJ986vZeC+xoWkr3a+Y7k59WCbIlj7YEmKxlFSRBPLMsy2Gs8R1xmoVrwQcj1mMVtJDH
XSOFNikmLGEDQ+m5QWsWCMUjMrbDgi4oHHQ+gmZOJ/fOx0wbzcHiF21CnBJc/yvPB9Kj9+T2lIvf
Bho1CyhEzPUzLfHzlBcJ8KKDiTdTodL/TM5QVvh6UkUeG7iIxebPG+B1L1ZGzDXSDbJ9fGaNeTxN
ZtUe+waS8w1K3+9RGPZL990nDDIRAv10JR0A/ykg35tY9wwC06FYK4hsU9uoNAJOR8lUhYoqOnDi
NIPj6DcjW2dJ8H03AL/XRqtDp4ajEouH5ovKOst/luRtOQ/nOmT3aksVS+L55Fe7rNyvJm/4Vxuy
ej9oie5n3NbhXq6ZUfyoMZ0HO1h9BBLBtIoU2Tg0ZXwD410K51sQBoh6+SbC3iN10clCKspx6HX6
f4v+PalRs+fTyIUU1A6WLiUBN5gXnSNxVw+/76oMbdliqO02nPQXy5uki+12YtF+V3Q+AbFQ8nOX
p3ysksQcwsWTuHUscr8Exqbd+6SIaV0hdUpc2cHcyGs76DWSFAUXAxVNqzfu1rIgw0X8xtrjZr1+
CVbD/3yjAMqhMfJfwQGnJm5I9TlIcWNCfYSG14la5UDOKY92nltsB3wm4zsv5htOmm4BaZzva70b
xIEqtUMjCm/D5vVt5YWTKfA37KffBpME8a3CMcGUSMDgGS/M7M3Tgsd6FGU8EPBlrnCbCmCA1Zw5
a6ReLmHrYZfDt6VHuuUNPMSKEowanHz9RKmqrLR7zRKwMC5aox/tEvACbpXMPLT7VjhBr52p2p9K
c+XdOoUNKuiwqASNwILHX/rr/BvxR9jE5xszRZlyrx9LDRxp910cZEisRf8A4yYbx9qXIBn2eJZl
YYGTBlpyrVysGFiBCJLQMVhO5KGd61/vKcvKXjy7n1UVWj2GRFx36eb7/33BQh5154QdKeesKIw/
z8aswCk+20w6orXryK97ot3ahgsg4NNms1yv/lwcpEWdgjW+10l5jVQIM+ucvDAvnuZ5rAfY87OI
vMD+VDQ0//32roZ4mt/Q9rt0EUCexH1S5Av6+aDMEY6zceVrnb8VdkNsqcHySLAy4M/SLFO4wxGl
li7t6+hrYyIFJ7wps/BrIrdvgbRbwxeb0k0iJPCzCGd9LJFr8ayBOURSifvgpiiEhN7elw2eOZmj
4Pj2XLSnXJgX+dSOpD5ru9mdju2XwubKunu8p/HyVlvA8v1r+KCgDe9kOeP+i3i1AXvusqX3wX3p
/tt9PIknF3BSqy63mEwCa1Hpd2xFpkfO4kjFqQer0BNbNLFADjtyK0moCxrYIN9vCPnn40NfV343
aTevfnAlTIpjTpZygt4lO+4CN/bI3GQcAsL1bkc2gayGfbq3V5P0sKBJqHS+RIZq6JP5rMqk6GMl
4ML8MhE/ZeEPDgmgi+2t83sNHkVWxcfic8nahajhaavC082VHnoQWi7YnaNxwFNWvylN3Y5PeujS
TsZK/s71RPeXpdQuHYxgSPzmnmOETf9QGhXS+ZoUmhX2GYL3WGyN2ibqFpXrimyrDcKx4xus6NUS
C3VlaXhxfVs/awpXPfEUPNY8VrNRdj9QMVpolf/Gyc+uHUYVW4zt1B1/Yw5bpy8/M6mLiOhdO7gr
g5Ri5icVGJOtlDf4QCnEY4T9YK5GL3S8FVl/iMdQuQqedlOffJHNf1mNgOr8QeMVIlkR8FUEudKb
bQirsvId97vapFvyPCgPBbnZUh7tVAzIXdwnt05ksTd30KOsGkm2/2IP5btLL+SbLtZ3qixN6EeU
nj+Wl9RPKvIzhw0ECpf8o9JNfxfa0hZH7O/g131k2oOUCnUvJdmni2/9WDdehG05Jy0aRFoOVSWE
VceQ88G14Q+kos+Qi92O3SU9EIE9c7g+wLBbzXAXKnglP9XcUUPdKUpdYXhsWmhSa+g9JW0riLCt
JQi+nDSryimTokI76yIp4u67UjEX+7gfdFAZmjhMN8CtO2YHRhxEr6y0Ts0XzWPhK1JlBLDJhIlU
6x+ZCZ1Mlrpowmm+zaQhI4ROw1dPCxCfx81MWIwfkjueReCAdIZNPzEmqJtLHF7gtS2hIMsBQptc
1QzNfd6Pye/0KoeXkuOO5Zf9xTPHDz0ilp2QC0X/YG0ZtqwQZfoCWnGId4uQo0uzZU66ZZtgPO4P
KgEZe5YuOwqyQQegDIvWdksAk9GCgpnsHSN022sw4r6HqrWjmHj3e7WbL6sldEZ9lV2Jmdmzfx7K
3RKPEaIxleS2+xWPQ2Iw9tgzLHa4zACCU0tWWV1QPMXJ8ap07FYUcythUamHn9a6ur4gliYJpJDT
3w76BSoZsMO0CcXa2I9o3z4f9x0hFDNCWlZOK+1pgPuLgYIWyiq8prwGdTELDr6w/LOKrEdwk8cU
aXpI3/DmSV43mXQ61zqe3oW0jDdQp2INJDXaAG3VN5sJNyU9p04ZP6kJKp+58EFnX/x0YLB6tG2l
fOWYxeByMinNiMw+t7kuV11YvP80mo8Luj5Tj6c6P8/JS61HBXwQC1J50TH0H5KtSxuU5+wYxPcW
vM9a8WRih+J+efAZ7hvctlYxodhKVAgxWQzyG5iKDZZnsrx6MIcjK+pi6h87RZjzru5toXIxYT7/
12dbzYdJrFjn1fIWsDmMvB11QUtxf80+IqiZzFJwGJd0f8PeDb/ex8tkeYwjJ2KiUU1k0+OyXgcX
E2Ucc821rsFe4+ZQYfIjDvh55mdzQ66fDiWZfvQ89qkEICNiroIdXYFtc9Lqu2Syev3Jh+vfwPK9
W6CWlZ/dh+zWIVx0JA+SyIIiAiOw2R68/IL+pLrDFLvm32Ph/A86JMlMozHeU3tzVlhNFtY5ubwz
4wTmGjrSBvfyjuv2PwyfkTWpqVFoBNoOKXBg9Glc7Wb7WFIabCqRRvm4LpVjngO60+aZqIyKVbQI
PrZNlShebQ4WgZFDKo4VOOR6edYclNZm3p8gGx/envqvabsf2kE4MvsiltZ1BDoBLiAFSFyfhkWT
fQmhjzzGP+egc5BFbMHNev+1W3X5twOeiAGURe5ZT9msl+woLk1wHgtisiEWlmoV3nhWISb1FPej
MUCzec+YYt8zfoVmVYEW+s0os/KFRdjm/sLLNoOke1f4II4MQqFPXVH8e0Ly1ismcNlQVg5Bvoa5
y2EALfbIz8Ry/6v/38UjUUDjDW70BzG+szPq5Ls48jYDrs88Oy84/gtUkIkfXfzMHGtqG/DvUjIc
zuHn49KawwRSlgiXiYhmxEbqle5VL9lXp5mR8YrOcO3rRdqNe1KAuJRZjtrgShwCKl1ZHE1nfrKK
ytDJAFL9CFtueak1iuY46OUOYV0342cdEBuiNZish7CzGB3SfCq7S+9esuiku5fDUr2kPMFwbcXD
zq96Ztk35e5LjSTyFF6WF4rdTE7MrknWIBvWA6sQNHQC7QsDy+c7mmmyhUqM6VRGyIjBcxvNacHn
cbbOc68IiNfpRkSq6wwHqsIKAAy4Pg0bnUs2bEcdI+zm7sHCqEqIReAq7p44bp/cBVZXydUTh5s+
oGeBEmZshkJMFnhwRSnPpqvXLXDQVgafJFDiqknhUjE7PlZ9qKzcpaAgNUYHhUL6BWa49vabe0MG
K5JAuiVuODlWKjHACMtSC0lptOwiWD7z4pJD9oi/s4a1LWQqbG+QMiBnZJW8YCVwBF4xg+8OxoWy
IHDsNTsSKSbQBENWRO8WV33CPaMCA8hgxmPIH1fP8LXRnbMP0z3JD7ErhYp8Kc0vzq5XxHtT0fxJ
DqXs58AVjIL1BHxNCIHtwqCbuSTWm2Oqh12GDqB8ooKBD7u4w5lKO0lbMNIhmB8tWy59rJwRwwd+
sFZJ0dxhSgcnSo79nmb5bMlWWUQ7ZV5YhtaAXlepVyQW/S1GzBZy3GLhe8YfTHhqXmXrkyq1fviw
vmM11efc4vbFX9B/5t4pR2ztalgaySzIqMGpsMSIOdkA4qpuvYSQ4iWVD0jxbEYnHOKs/Nsx6Gld
ni78MmX4P2hSF1XiDTfW/VRrUf5tCcie9aGKsG25bzQkv+V52ChQGs6WhFv6uGBRs2Nqetn1Q4St
GptUidvJTk48w1k3dfBaKdaYWMVQkeo2DnNmMVeKm5iFjJPyfFwQZALtYVuOjp96a6pNzH+v1g8O
22W7yQhaGb43GFpc4pOfy875BYABJJAREC3eHiZ1hQQ9Tx9yw4JRGe/NpUORDuhaIjRoDUGMdAf7
F/mCqOFxNYtrirsmGsdWs02urUuKb6oVMgwySLGCnAAbaFc/uDXH6uWvW4sKLBo7NpuCOMwvLuhf
i0AMrynmUy2WA2uP40O93IxPt9+KVt+4rrtUWtJfoqhkX3r8sZ3Il8YxMs4kM/gL3nR6B3S0aoTC
V/tLG2lrJfmmYIH24vv7e4IBIKa2EulikwgPv7goKgxl+ZF89oH5ZbD0Qv5o1bfnO8uPQy/V0Lm+
o4ParwYhiAUIrjvghZ776j+azrsH4rz/KnCPhbJ+V65GnU36t3KTBjl0Rpn0Ws3NbGKAgsHXxdM3
c3u8OUNswCPt1KYQ84HAsRaq0AcV3AgDbhlcjwsP/jYFea9rFo2PAWQGLfrXIWllFhr6Z/fIMYmX
RdwVNP4nBwP81iegGsLOIPT6kRo2754S6LOsUfQmC31Ul4my80gTWoqNNHUVUmG6torcS5bDPvOa
LXgdcL8oQBMceVKsbC2E+vgwvdYxdfcTPFkN/K5iDRNvBCRFRnYp11gMJ3Jpj9v++kfFX6p0ktzc
7tKYarz6CIblFGEpsCD0QzIxecB0vrIto299fUPJrRyGo9DIQ+SxEe+Pm4CaQENBcFcnCxM9e9pt
6CviaOJt0x23Us4XTbgbNWWboemgfM2fSqkbXY55Cs+6Tq7n7tdF7DkaqT9GJxXehVFInEbSBySK
d5fpB4mFLibhE5zmsbRG0fL+IrdG5llE5TzqDD8xJlcQLCkSxgvndgrvHcrjE8dhGzpZnlSo7BD+
sxWK7Ru2v1ZgqUyV13wFvtmdnuSg+r5HlEU4UBq14vUtfdQtlc459Bt+3cS4anfC51zOIh3z/ghz
h4iKpY/JQV0gY/XW0uCednnYlhxgFAX7KrpT/WegXIxDUzl1kc5IJ1Sygyxe6tjy7uKmXeOeV4b2
qWryiUoSpvdpwAA/18p7jROXT7LQBDVf/umiBtOhHv0wrWjqANSGpkmW791+DqZKi1ko4YNpzxZ0
bu6N4L1OLciByKlfICeNFu6K9T3jikC3RMRepRtS6+in9QOr12pFzV3zib2gWpTfMVvgQMu9NZnF
W3pYDV0e5ol3ptUtYoeYrVTH4PxtE6J+fiqXufBIXHiAYiTEo1v39ulshjSrfI8gjiu77Man8XNI
+T16WwG1GPrFe2O5nQnIWwcGGSnj6jWoT3+EkmEqOtfxsbNw4F81AJPT34fYMKz6PqiQwE7QrjLt
5sIleUSWZwMneUnEMQ13XHe3Ts4PnyEGiaxuPqG70ZMs+K/kMK3lKlEqKtmxEmWZU173FI3cyXTy
6SXHGvjQCTwQQgAJEkbcJyENW0aVvF3XGqVVibMLy0DlIkanqgwhKHzXDEpLoyU7C3cJdHpS4i/Z
AuvIdpuo7D9RCEFcNzlGr062qwu8I4hF4+Qbt8m/N17haPL5Yt29l2j4tIhFaWlHhQrGbMsgQP7H
HbOUY2SmPzJX4vY5OfUneSETf+QXfOpHjtQcySO6+wqJyQOxpYgCOUrUMW165uRpxM1hhjw8gWwS
aOYlHEC6oQXg7hGZB3Pb2CHDxMQKDPjmgaCISssk4euPNIdXcJSfyhb16hWnVMsXkyFSo7AAeZQj
p4bM2W8bHTHxuNG2W6vKOdSC390CVhJqy4vCYgoI5cqehInho+2LUmTKEziSiKBrVt8Hzoia1Anm
1BTNpQobYB4+IGZtMgpLhIgF3FVQJMrYlqj6dqPfYFgIYxA4c+1j9QLBM30HHCpUMFLa6JOi3CZg
PvO5C/MynFuw8G5QVCnZTeMjpaWJ8VwunccniF/2b+txU+Qezhm8vY+va09uIpearqqSJKLgn8q7
BLM1t6uJgGvRIOuI5NOpPnSbyL/njIptAByrGgwJOWnTFJYXOjogs9Qz4QUlJ5P+HAmpmE1uP5aX
awPJt4amJiTZtrmu6hzLUmvYIebGIvhHgvm4eqq3xImViTBE9r5ExLgbzeylXdLzv2/+dXo7sdXM
9sDBgxIQp7oAtNpuutG9DrPN44XLi0tNkr4IqBWDJI0yAocLplJIZKV2wmFVmHUfTl5f1dE3jTzZ
dOJtoCHQylZs9JJ9rZYBT/G0H9QHxxgPiQoy3zOKSDW4qGoAdbbVl9rtC0DfcNPumxaaVQH+iBhW
xUnBKlQphUc7rd6LwBffORYEyPJOh5nnGsH66nJKjAcgbvA2nba0sz8UvhIy+yKT/+bQZXXv44+L
pB9Cy+Pzkg3LC4DstdIDldF53SvzvPiyRXriSBhloD+UKeQJdB7yjEXr/l8wiyIaKge4l5OFlV+p
sCa4SDDGjzb8NY0w/lmkqqllSrXoiVWddDA4KIwHX0phgMYiVZsGGOkShFfamr6qH1IPY97BGa1p
hCa7SLHKubyO18ZR3GnkKoE2yaRQ1yaJAAun1iyFNiRb79F5KhiUnNYAWJW2/qdF5S+uUP26v6gy
W32XKSA1kCaprooula9eBQfXj/WyWnn8n4qCb/JzXlgvhA4MW1qNHNizB3k7q2MWskw04ub5979i
ANKDSqKhGWmXBj+PsnZ0hk3yIRjY0khRuKE0i1D3ShPLvWFv/iAshyZzMJ05xSGuxKRXmYN8XGXI
H3r4mkoncFLOTBInc1hitFI3T9Fz+a55bFvtOYdkX6/5pH6OPTlp2o8GiBFeq13TBMd0HpmOVfZv
kVqMXP6k3EXD5vL2EMNvkpp0YI341NiHwGQy4Szgxx1ILidsoYkaCh641zT0Yth9wq/akgSdLgyC
wmkm72JKi3psMJvYiRF6PpeOaJYMRx7C8QgbNmX9klTCmZEq8ebTuj/8iHedqj5sqrS4Rm3iuQDY
NhGDrtc/+XHbgr6Lm4Stnrx9gJbue8Umv5dDVvu6XPPIXjeFl1XZQBr4BAT5gXcE3OAhETEmDcax
6vK3C8h6I5BbzKwGIUMY25iE8NHjCsDi0taWVJSLV5Fb6m+HP0YqcQ4L3p+Fa6XHE24ETPgVI3Fv
YU9d6B3gqwrKMY3W6VAFnNycb1ikVjUC1O3npDOE+G/k7FdnGAiCmEmNcRJ8K6tfLTwlp/gQpSW9
N994SEnAoIzInJo0IYZeX/uEQ6u1MctuGxnLg3x/A/5P7Qq0lqPIKdaCMnl6PFHc1Isvml5qPS22
KzLpKn0XX/yMK4GR2y7bG9k+gMkEdaBgK5ov7QGGSwA+wBVMO72suFPOQAx1ujnm3/Y9PhsfUb5U
hUkXfSJ2jupSId4MIsvVZP9FL6LY3r2FczMYuwAyfABRH4w3vljfj1redmFTa/oQQzUErT+oeGOe
hFV5+noGqy8ZXlVyt2NatQKDK7JyacsgurtrsvXykOYx7ePXlG8BJZgRuhs31dwL8eVoCKkF2cXF
dqEULmrXGWll2gqSZyMIKbRJssgR0HN3NK/YPUL72pDm7D2LmA+n4j15Z6QPPVUfTuIxCNbZ/Yfo
YEfptYhpO+SKt7IAt/0aMaIlSpmwBPRDJyl6kb8lmfUAoMwfnknh1sCkiD+l/OM19XE1yvmPurpo
y8X+iUDNMDG+e/WFPUBVq38DkXXs0nrCYHoUUnvRdgJVtW5vaScl/xNMSsk8t+KgTB6niKDTGVbK
xBB9zCNJQLn+ALzmZziRAKU1/3UJs9UFfLuhVhS1OpNdFDv8b7Gu58/G79Hwn/FXFKavPztUtxNp
w6bj5CJq5RBtEmsjU+p8f1LXq8uKmJyCAYUvhbfQKIIgKGO6L6XxovBOpWWGSVpznctWzv0RQkup
XDsYt2dBRMaLYKre/OIh9PQxuk6/UHSuSH2bZCq4d7ixUj/AeDxPk8H3iayc65wz80qwEBr/uTUX
RT0cbYrVmvwYqap3NExiww1dWEa1SX2RD8exkBQnBuBFerVOBkPAoRQUZWugmtncReqxHm64h4IU
4SSS66A/VpIW2AMKH602bnD+yw/nTtP0Q+zIbR6/hmeRrA6Qc7whSSpNfRZfv8c4vrk5RcnXz4HU
qdOGNiCE6iNdSxnK8OjQ4WM+s5GxL+mz6BPdLGddNBSvZuWmzs4aNXDKEPpLcCLIjm1+iKJkEgBI
B1Nkx8e4StzGGPkdOnCktQtqoASUhRiixbha76/fgSn26S15XQNenK8xUivA1k2T5hKy/by1I9Qr
DmpghwV+tCdQhcPNVAgd1Ln6dgx6HFP9MoUaJcXM8ecIgcn5r765rDFzNBx4FCeF4Xw/3NYEVQww
ZranUWc0rtd8JBf5zB4BHs3mYOSwNAAN+Fj7KRG00fvX73WKJi6Pmy8ccyqgpIJ7RfWDOP+gXvbN
hyFDJ6Z9dIT27tOq0XUH+r+aPYyRgcND7IM9gYqIvhLjgvQR4qn3c/XX6CP0RXx68M8eD8mBLg3s
zfkDRh0egHQOYSHRJKCYoDwqccIQnkZijFdSjpLxcUP++GCp1sDBQB9TQC9aOPeSx61GmWWDvbnS
FLr3MjvCMEXzEKnGy4Xk8LBXs3AJz6OF/ubvNMXvWRiT+MqT1o4v+Pia7yvxCAx1Xi7gQhADyC9Y
FDSXEfEWd4MYQuayhS66S1Kl78NIDRV+gvilTAVwyx51HSJoKdm1piBb6ojtAh5IECcvgziYoN0l
uX/O22TfM+pFE/HPzgh31u+rK0J+zMjl11MMSyq+b8DAgae1XjYinKoZcQ2qa0Enc9OE/V0M1TTg
fs7ivQwHVKz1pXhMHqN0IOsunJqLtE83oajqFvYKjApsb1fEg8bJL9X4F0Hftf4B59/RlPTKV8zb
2F7NUlmNuwSbCqVqqbiv28xzlda2TsIVIIDLd7+xX9uIzumUTCzsS2D6C2clIZ6/G/+fnTeY5HJh
WDsbGdRY86ag7PlNuBVa+VfVdwoWH3H9pBIb5eGEvDcPcblLUPw5HCupJ7qtFG5HlGNcmurlry1S
ym11fFuZC+JC+DWYwU5Tr3jpxVjJ4n9kbDtaGWiX0rsCWN2f4DkZOe36XM6/OcutppLwPeMxB5rR
zVrDVv9SR0kJOFEH9P20b4vD36hfZl3JtcrHoi3N5Ldy07dI2zQaUT6kT03zva2LpeJOY5XzLD53
Ni4WsxoCT9TOvfsLiVMF95T97TPflbZ43gkmqk6QqdsAD6KPlRjQnxYmK9REIipAu/8PhvkgaTQp
FpCikOnq11p2mPsXpiAhoStLuRT7jiLL9KGYUyWGDM7XqJeIoFnN675znTpDHWU2PUzmRsfaJWCZ
0Y3Gohz7eXgVEDs24E463+KgV7GI0ygyH3lqklvo15Og0G/aV0eCir/HrqvR2PkwPnoN+Rdj+xHn
hZUf/V584BLVbs8qN2b+LyaCDK+ZrjqcUPpn3DTDSqY32GO/b3KiekT9X23k0a6GuUobk8YaDoPA
p04NuH2yMlfMTwTp5H3F4Ks+xpKmqi8tgRajXhRfCiiEoH+GzgxGY1e40HwLlS3NnddAND3iVOCK
7b8MMXMzMsFJ0Qem6nFS5Yp6N0SQO9GWMRPUinJN9rCeG/1nGFubKiKE8YfWre8ZO2FKknpePsZs
YS3ivhUG9Tvd1zHckN2mWE1MKwNrmR/W2+pWrtU0sx1xzTAMoKsN1rZKNGrqB9uWRuU4yrepzpCS
+XVHtIvwsJhwoha1HXsaEQMEmrZ/si/LPjxFb3SQA6nf41p9rOf4gBhlne3JRpRd4N528fZvmqvV
CNHWe9vOsSoP6d8nkCEgE1eTN8Biutm9ZPTMdygMSncqEzLPWkuslq92nyIYVqicJz49WLbbNKGq
s8q4igNPiH1fO9DztplhIiYX6t7tXT2Wf0Qx0rvDKiVbmWxg8v0eejYsZTuO9bVLzkwqHNjD1yxx
IgfNaJJ7EYvcstWjb19rJSceqbU9uXtrU8fwRTdfpL6bC3D8zzBEnRhZGFYA0Q5GPjXDBqUACfLG
Y68PtkyfHoFjRAfUEZ3tzhmJkJoahPXzbJSwKTHGUtTxPOJ3wPU2HnNwwXhWS87lR6gNs4AEvFx/
w6qpgzhw7fOmwqpa7IQi2Zigo4yaPW0uf5D8rxVLf9B/yNJy4KOhdATLB65ZgB5qc8Kz1dy0WA7o
ZZ/4PTaSbEA7XL69vFIRurIWIUaB6+9RwQeu1YG5aix5ETfzMJMCokwOS+CQ5KRQRYktryLeNTAd
ODGHbd3HOYtMWSuwbYkxwUSR3xXYlfx++lQn7rO92VtK39++82JaWAE3UmFQEIig3CyBC8XCWQDF
FhJMTP+t78mtnHbeHhocrFQOJ9f+LFzYVxPMVKckG06VjogT7XpDrBywSrfTFB0STF9aZQSa9mE6
XaS83hYzJNvlDTTpUyyb5IoiL+O4vteRU8sSli9ncYefBwGrOVUShMR5sckF6SLeekXv9yBJiesh
iQz4Lh+hmPEDcBGEGNA9c7cbfvaW87X+Ze2/JalFkraEEiBZCVkZDoXimiz0wWINwkgRubXNRmbb
OlcnsG/ME19Jg2JIv07dv6KFFV1N1LnMFWjP1dLlnzhro3GQsjzuidsLhdLjb6d2rYdUVuugUiDP
zjOCRrmNm0tdj/A2SN4VWyylcF673PI3G5aMCXva6VY6pvmcvyeiP30sOD4gSr3aTk8YKf5rOHvu
0CXbFXOafNRDoMa+aRTMwS6smj/JlmAvnAGD+Og7Vhrgoginrjmk0nnHNJgrFPp/f/UaOAnRv/7R
6WCLEfWNBixGo6eTGT9gAWlpwi7kzqFF6j6dO8lL60VdrPOl+TAlnY7Ja778uTfIzVcUgBbxT8vI
V5JjF9Kfe1jztGhAGWD/5fQflucevonb3h4X4Cq/Rp3NptWcxh31H/bzc1zJj25TFXuQ5r1fhfGN
nKkBXpxiSEnRGyoS5WMKzZ6sxoVBxUZwYtiDGX/PLXVIUueM0E9UrZBTA9HWH1WUVGJyqfwd0r5g
Gsvj523ZwWlUErRugMUG++bS9lnIWSBxAph46Dry0stnPHAYVHKSD/Lxzz/7+Ph50iCFQVhRzJfS
3kFqZm5QtvXF/ieCniJeMnIhGIjq6aers68W7SPJcEf9MpypEuS2W65lFWCjZhnD+kCFqwqwBwe1
gge6p22tr5ESC/muCeBx3v4EKq4Vh+aOEzNLGMG8VOQxmJ6YdNOuQBwrPa408SSq/rCcqgXJNDQ+
NrwfAsG4ErD7J9jua8y+f8G2HgewT7QTYdpK8i7s3vEdqfcaKa06cSAzOh3Ycl0DDz4D3m1rxIjE
y777HN6NFbFKUNlKOnzo6ecvzQQs+Q+owTukwLbKs8zPQMFiR5mr2JVuGZ2dpEB5sKvQmaIk4V7N
0X4/gchKLek/My+5TvMKJsDSdKhSRYtcmgsOQ52P2vnkQnte1CAGZSUny7wBl8/2WenpUoca0F7J
h7l18F7+b6tIqwa6C3IX8ggInVyjNZ0MINoJRo8XWFucRnHt5bY5tvpUtKkO8TCvC0rxJLtMYqt3
Uz+ts8VVmbnmoZBpBWcjDq7OXCU/GIuCE3nvtoMxXxjiTJ5N2+x99kVcNYAdTy2qj0z+0OeAGm0f
azwPAS5/yCec99MVqwD+gKkkA/sUHZ5i37KQ/x/7QJS5/7BXu6vVkcLZ471Lu3x3eH1Uz/R9hLWw
5FTywBPDDe3eouTWu/+NGZUQ0F6RvhsBVDQzwVo9r9faoZeQfCFyuk5PaIjA7N/isHe0Y842UoSw
+Q/uncDCO9m0DwpKpeSzDJHy7/dwqGb+u6dyDP4SfXSn2fDGauPPQ0o8wqdChJ2L3l+nObqozS/X
1LMtgTSpCl2MZdm0j/FiJotVvFnjsLPHQ4DB7Vt0kpaOfLWOXn5XuwlHdOZhYeac1anOnVrQjFl0
95SRFkoT59VJNKpx9bIOv6mchaYxyrm13inxIWUM+ff8Ya2Jsu+O07urq1QmfpIDfV2T6JnUTKIw
9sVuFk9xxWiDTcoBPhg3bM0358AzpIfceESIE62yZLdLeGrrmEdVALbSeLDsqdRn+OpdT9qIa4Ew
GDsDSLQFzVpsowmwEu9D6JD+TTmR222pMIJWPCw6uf45Y2eO6tjiBAzRHCRmvYHHUav95SGXW/Fa
LE+pvKLMbyvfgZcSlWvJGoDGXD7QhrKMx6W63nTYmGB44HWkrbRa2H5uwqQdTX5KlFiF08QV2bTR
Eg7ntbSHcTq00LffeYf8mqph5766MdfM5H9FQSb7hNc1uTv3uqs8eP7Nfo1fLxjvc29tpdkvg/Vy
TW+sECAwsA/mNI26IxESJpsHYUt/sZU03WOYWmg0MdyJebHQsK6wBR56/0WX2Vu5S6KSpQJKAm34
8UlP41LyAhzFPsxvVPQrlpB3Ef/yEAhsfaz+rhJA6OXEEsW5dU2gzPEjA+VfuDPreXEUv+y6JVlq
pglJ5rZbyafkgM+PpuhF4ICvPKZDfegkSfspq5rhkrM2qodfbxarTqPlyR55jOvFZsFZg4Bmk0lM
9/qfQO1Ul7WOwhcR5yP1+PnZI+LvolGcFejA47nRPIGtPLcsERyQkr3Ru0nswTHfFoJc7SzDDg0h
2dzfxdWo86MIGcHvrt0daIlvJ5zHOlbZIziyzDNb+HF0QcPXFCV3PlXe5wg6e83ksvLfslNgyRHV
wG3ew9sjvaCBSp5GcnvLlin65MrbNoGnp+in8j7GY2GQihQ9ICbo664P8ctwsrO65C6jaPhpdiEp
UmrpnvYWzQT7CRxjaWNUvwShd8vnc830PFTv9Zh25QZKKgqmmlW91jcFjKLNk3OiYBWpDXOzgOfN
SdI8ccfRxbHNdGsLLaCfos+TD9t25BggLaZ74koOypKwcW1qPfhYPpIvIa/T3PTsbJF0LJjIsHas
v0YyKnaahCoL1bteCkQcaadeFkvsCRhDoKAy+WBx6Y9yy6LDYXsEb8NpdORvgu7ZPMLXbakN8hYa
T04Rz78O6xK65L9tmUe029bmf98xgvkpTlnJkubpaCzteatupBfDGv/nVhcFGGVPzn617uHucBVD
ZjnepAe3znA3DkQ7m2gMEqbP4rYZ7eoUZ/XU8nIV1+CnQWtzZOsq5ccOETbIyX3ePyI/vStjAklB
su6bKsevTsSjxfptW5LrRC00SBZxjpbCzwshZ3jZDJdG4Busge4PmXuYBLzlPAqqUWM8TcUVIHvV
y6Zvzr4Hnx+dImrdrC+GvvI9g5oR0a7NzbJyq2+Hv7WtYrHnwGn9Db/kZkU75eSiWGyVE8iDmbA1
ukr28mnpNyndiNOr5ojmsZV/Nn4h592srkeNQ1Hd9u1Jy2uwcvkZOaxDs0OPWD0Fvxu/tfRebGLp
pTk1YBHpkdr1HQXSOPKK9fJLe6e0k8L96oyIS0m6z0DZhuusll3IrI80DhtzdjMJOZTia39O6Ll6
wivd+DnqkZIdn+WWughG37hMY7i+KAedw83UM7OrFI+/kpRZUL82W/E8wdITzcI78RTHcQL/mAmt
8FHO+fiT3zkGPJ8uxrZW4EvCW4bxucuRMFKYWkOk9KMlK6w3ehBgSePFOHNvSXQP0c40/jh7W4Z1
1qrxDDBakJliiZVvzgE4GKuz3EggJo118eQPF8keRnoEgo4M3UXAr9yGUzqiwxJwoiABEyd4a7fJ
FY54/uu/Fa4wVsl33O9gvORCOsKT6NgwTvjTYRxvxyBfJF1AwCZcdHV4jUOE+OFBDaz4Tp9mRqgU
KeSOGSnOe3bbo0l0gyHrNirMjpY8l7uf36D1anZWITngszs45ScXJkRh5haSqJa3WuLtNnzAVWmp
C1n3i4Q3pd5Ia7Jsrq9oMDPhg649cEjAyrnkdnTT6wNY+nHIwwWBPz6+wgFSqyvheraiHQ7Vo3i/
+0uAcx57hvTL+fm95FO3kPeCUafGUwdZ9r4ETkvdaRkiwSb01vOQ/DrUdDOst+5N+WVuAFXSZB1z
2owFokD4WiiG4LLO6ayy49too7hhlsMoNYVLaTlBu9+dftUv6B8dPxPOhDCNmfysza5/MPClGZBk
c0oO6RY2mr8VIHgSmdLFfeU0c+jAL6DIjw5m4MH1m2DDspJQSNebhWVQOjzcXEih/U7k6OojZcCG
jPzAVYAM3wuihrOTTqUymjjq0roIQYgz/v+S0hq0bewPVVHEwbzbcz4dTYm83J5AZ0GInHQLefWG
q08RF8+p7rWK0Np4AcUgCidQcqHsQflzyR7drPVznhjl8lDIYMGj1jOnxKqWaa3RrlajKR5xEhz+
9PXxPv1csgAj3ReTIWlo7ute8s3+64vLdnGdJaQSbSw9FjnKpqWnaez6IIoNCsniga4fCap7cJvB
npofvb5iYfXcOCPvruILqiuguwjRFOfn35b3plzYH8fDP6n34lk4atLf/UmnBSQL4EtZnB3ZnKdY
JM2kkmD3feiBnvIkr2loloSxvaX37dGlQ9pKW0VcrbgiY5xrpKg0APKsar5CAjlQ728nrIcDMxwa
yyyyQLr91w1GvH+W9bIpU2fQFMZCgt8ORO+1ghwLNGx/CCqewuLT+3UYJ3fNuFvhbjTvT29uJGdx
qRwPllDL9CkwdTrQjnrTnUQqCBOo4JikDqElroQ1P735ohKGFKt8y8/W4qDLlP+yh/x+F6/YxM2N
Cji5C0CfpcRoHzfDlOLqz+jemy/bN0ZHrk+DWy4jsr4cmat2QxaJuDddndyJYtwT33BWvE+28kXW
RhmQYpyMh8G4u+Kdd5lrm0Q67O71pZVLWu4zSDrhaJEMfGMa1xTTGfEkvkGe18WtQAQr2oimPjzJ
ayX0AXPV9qu1qhDXJabMGUcY/m9wqZb0xCtDcGKJSH1TaDclCx/OLZta/TJlvx0Hd2lKrfHd4EJe
WS+xhZVCIBjzghr0V+nnjERWgew1Sv6G11qWt4oyktOGgPtgsN7v3NJ03sEok61Xm0K0HXcxWsYR
ghbk0TSpdBoWLceRvhuomhwyNjZojs6smvVERyzt24qlQ9Fmj3ycJ5KXNJ7n5MWp/VO3XD2+MYYl
MWRJ+V4oKln9dBMx5fBod/ETybZe9jzapMg8apq5pw4ocHUinUanA2naSLftwzZ3rxfAhIagVJIl
cIzqbCdpI4eI0aH2cp2NwYmJ/02U2zqohK+n7vElMpB8SVb+eVePmvXgxNZKkR5X3u6pJMB9p1Ev
HyQR8pfLk5Aj7YfoSgeYEP74GVJDe9xWxFcO8Ir4ZOTAQHDVexLU4IpzSBlec/EQChlozgk1p0YZ
WT3b3gG5K2dYR0QPc1PpHb9/jpbW9Ty0xuALetndifEBonM6k+XuiTphgJGh02riZoEiIhBFF5p3
scMsg3xMNRlfhKgA4+hQpDTEoBz+qr4zmb82G4Dsmo3oK298iBmbWqpJaVEkkSf/RyaLizy24St9
3PSQa4G3PS8en0xA0avQHsMp0fYAHGXHKxJIq4UM1dBR+3MABprA/+CzBovxeGtLq2+f1NEF13fs
F8uKVZXywN6TrrRcBdMXsd7bvjrvnwgYgjQZKadSLRIxgB24vsvOaKYHjnAeQ01yhCeaK+2fJW2h
lY3wuq3VhExtxdX8VG46HJLDeHApvHr2lSw2ipxaWARZcNc5TsKpo9jo3esqUJmo/cIqxSBGGUtL
hQMu4g33tWgjxyUTm3v2OekPzdxynoIDj7G+vY6+uoETvlNuSn4gPedtaCHKR3w+EO+e6FgkpcWO
QqTv12a1U/8qc/jI9T+VzcLCEghxDakEH6m46n/02bLWkI8u8PG1wYP7VsPX/CezEeWiEh6T/77Y
bG/Ec5xmjS5/sheqVfdUm0l6pku9+YhS3QgsWUxuExK8Fdv2mQ50aMHeDLwrd/X42+wgqVwG9Pbt
lI5kHwzOrPptWKrglViv/CfBn26nT/fsKUiAr5k8n4DGWETR7G0g9P8supOTxVs4WhSIZa0G+5Bc
ZypqE0j92SxLCNrwiiViKfbtY/62u1U7JVMb470eM7GWbltjIAHiRki14f6YFlJgXS5cFcve2asM
PEQiHOEvztKk9llL8OPh134XvYstB6RSsB4EQ7vkFx/ZrdFvBil+hVpbwx1SsY5nXq/WiK4/qK/a
KFzqNTsPFUdk5cOD0SpYmHPoNmjZi3ywEQ1XTkstGD/xy5+zbqi1N2/mNsHKUn4qfvq6lRAqYA2r
7jAE71o5KDvkagWjyi6UWp/xSBPzUqZsXGRrl8NQig1mAlzsr5/vOZTXv4EzPV/JrVIpODo1/Ro3
WOfaJqNNqIosHJrn2sxu1/TsnPsWQDHhSnwuiEsCCNjiJwUtaQM7bgCCtnk+SkGxmibO6uLAuga/
x72nHZB07znk9NnDBxB2B0FUJQP1b3W6W3DVeuZrhUFBgRoZMswBntENmbocZ+y/l+MVEJuFaA2n
z7Yj3vrv8U+IglYCyRxMnuDx+VhkcTBTWNxAWAAz98wi7QYaL9lQ3zNGziQeLJSru8NPg+3hZ7d6
6/8Gksv9GHp4QxCxuwAsWyQfleFoKingcYWkLI1s3wjozXqZ3Q5smOeUqCUS3EwpwCTodFaosSPh
q4amk3FcfwZKWnpf7YzuefVZoiETcQQ+t5MQ9+7We/DLuEfObYpFWtkDg+Yl/RLtTYNWuHodu7zf
fWOKiGeDZQ+5xD2i7DePAU9vyUl477rBcwroPYM5PNm3qo0nk2OnrZe2EzaFthk5hGia1wo61kYm
sgnNW80JilquOz0w5G415zm6+WwqjN3Y97/amU176R1DWkQDBhh2uWFEgHzBa+tXQ4P80F5UQ9fl
H3SpoSnBhrA91yyxdXM7rI7Qz0rIGpoFHqKzAoWzcca2A7oL0SBGgrEknzVcDHKlOxrO+1yYZZ9G
WATCRn55TrVaD8jDnZsroOVO2jAvA2XgnA1Bc2MQQ1HQcA4xoLD2A8K7ofEJ+ePbw2QIRo3gaBYI
mgLYuSSlGgASq+22h/wDc57Bp/gm3xnVlEoWJx/6xLG2JcxtemLAZzbgVTNfR9czJyRZ80DttE54
uPB8vlWYNszSu5MjXwxakwfHlzpRtNUT8jay+Lt6Z2slZ0Z+xLQO8neJhhupkeCPNVyeit4nZOcd
q/VEedrIE70O71OVqEA+AOEbSPFxEkA4+TY5QSHkE4mh1MlgbZfla6T42R/MaOhoKo+xrJ4uI5ev
RfjIOJqbpycb4db3NryBW7PPtXKMa3a9Y/I9joXbznuzTGFV1omcSaHpIO+Eykp9ai+5JPeEXTXl
4ptYV7QVH513yLH/nZwDcZc7oSp6yyQHW1CwiHUpTzmsc4oUiK3+7fbV8Gpl/Al4M52KGrHDTP9K
EBm+5pFIxzHLu3x91Jyvsxlu/rfd633NAv39s4fmT0MfsdeYFOkN59WK5F+iRbkYn6K5aFVYsvBq
ppgxxoJh39JJ9HtsyHNHPMj+TjCSmofLdJBYI35r8IV7vyVvuoOhJ2QC0yeHVjxxiPNFuTw9w0Hj
byUckOd+5mx6ZM9uJvs20MJNmp51uhtkCoBwJpDXns+mE9ruvx9VyZbPSfTwJ9FG4kermPyDZ6LN
/DYqiv8z0Jwz8gCVj7SiQcEfcDfUWOeWV/t9IGL029yH3ECwTH7BbQaFBNeXsErhZPYN5BVMeDf7
ytBxt7Zdp2K6b4K8UR1cnWtne2A4YLWFQYULzbNsoYyo5RmdYTnreHAUvZhPPDwIx8U03to/tZZO
5bcDb4nbjMsclVfPXr6voRCeT1FjYASJMCVTw5Luu2exqb+ih643VB2HOlrJ1gFBBG6pYnrX5Bny
BPPghkJEH3lO5Vw777gwWvopwfXH3d9UeImbrovtKF0urjU+ztaz4G+WVpwbjm075q63+LITgOX5
jTO39SSxUpA7p3h5bnMxbSo0N8KsOHYoDa+W2CVTiqpCQVLaV/7Sc/8H4MgnGFdzKVgJy0VExlra
wHaOJYVsL7tfZIE/0kp5W/wKvZAyiNDZxA9gZuFQm4JiMbv2k3FCe18FmpPoDGCbErhsGr1ACXmt
rT9surnjEpRV7fwD4Hv1XWdU9T4szacBZibqko1/5wbhx+7QZec622bJn9RfsAeud4ZICeSZc4L8
FvyRnl39s/7mmb5XMXdPi4/bmpAZMD8jmpjQb8YCx1fn6uzhPZJkTvt0cS7Zw5vOnTl6v+n4ZZKy
tz59wLh0Akx4dqmR9y2eLFuEriXNtNFqz1SBmc3ses7lYCwQwzDhhtmKQHougV7CAGwBhtRWkgFk
eGSvmFCPvYz+zknJo7egrdpVS63+2IWLePZG12QVAnfUjfr0m77/qwpGeOjunbzLJoZDboi0Kf5H
x3VFFkrVt6OxIMxdatXEWFndZSBrQ6bn5uZjCw0EfFbnj6qTFLK9TzV0zWdIXMerr1Bdl2vQaVcI
9nYQEhqR8zli3WAxwu/j2IeaBWCC8/a/q6TRDzyUBYDZgGTnxigHZkizBylJfgpewVqXAjFQ2E4l
SvVyUpX2UyjjTPbERf1nWYx1a/spcLCBwAO/wLnj7clvvPZAUPGxS/uN6liqsWnMPt8J3XaOZvex
RAX4HG1HayMJxwqdvuIVKgM9JftuU6dyht6Hru/o1UVLRe8kR0JIWO5/O4og5m7CDZ6SHG18uJr2
idHB46Y6KNZMKKa3b/QbMhD6rBbNB/FsqOt3h9FS8msZhb9UfFJnQu9M7wk9pcezTFz63wZTB2uc
0C6I/dCEbjHDR4R/2AvP00E1YPpy9IDMqGNWDUW2imOpG72V7LJUwpzAk31vRGaUjgkefEoAqUe/
1OIoIH7VlYQpJw1eWvxe9C5cflXtAKU1VLG8wbLLqgCwjIHzD2ZM1Wj2IDk8VvdlQpHFxHU14286
qMu38PVa+gp1PLGbzxDLrikOKB8Y32uGOdAyucDsiIyx+7Vg9zWBw2FmtlA3dkbpgG70M9GHdNC2
rF7zkXwy7fkXSefkBTrzKZywCRhvN+v4zZNiPNUouYy2o5Y0+ZyzXkIOid7ZDXX0tTJMzwE24uRO
acrRTyLzCKong3rbyivKXMZzGoeJCkUPd5PNjRpxjOV730W321N9PG1OLh+/5aPbYMBvJ7h2pUnw
xSkfeeLVtn8n7RQDp7lthoIOdwsJdSAa9zaX3E4g+zxaV5wX3BXapgNhvnFPEeyQoreanSZvaljL
DxCkYt0+xGjPj5fdK04ZHDsUmYp+po0zkFfqAhBdcITe6xKb+wbxORIfNAeiYKbusOsdO9srjuzB
MOK7N24/B0hdJ97AjgqGB9IuLp4ZcjkraHbcqGOHznCtNo1SVmpHOVY78WYNhEmIWGI/atuU5kia
n1C7BD2jfgFnGzd+hyX0+HYgQ1J+I/HMK/ShqX1Gplht0SDS9y6Aaajv+nrKtZdMuh9pfLXgeAPJ
S7z8OgBYOXdjeUB4ibEJhhTA+Qmo1vZie2q1cbh0Z6uLsBo8OFGIWmtYcBmWmfQyZSKUTvuckTA5
XcrfddFIgJcp4IJn83ev1qEFw3qwVF3otluMlxIROYZGqGDPVAFx5MKj3Aui6Ak4oOyPNxO+2jBn
SLp84Iitd7xHgSd/M8AgsC3iTNImHRyjuBgz7SG3bg23zQ04YE+lufM5ft0aUJDLGR4SxuqZ/cvn
uA4o8GI4C6nXEbSNrBR0QFooxNtuX5grFsKdbKC5NlR4xemjFcrcPZpUER2h3cnMSaqPv8SpWPPV
br0AIk34xTRC1ebpzcwHui9WmWUEib+XPp8syJf3lqO2mTd1RnYtyeAjXbhezLxySHRabosGCWfc
pGd5BbDVMVi9dIG29ckBHWI8MBT+m+PJyM2S3+wY/lD4JDIEuMIhsK7ypCq8u7lnl+eaE4gNn1Bk
SQAOEfP6IVbS4heQ2v89JSf7uSaemv08aEeUApYzi4XmwVs4euI7LdoU9XGPTASLO1td2+4UOO18
V/sHKAaSfMxNiEZ6x8rScq3JVMymaTqE3tr35Mh5vrBsEL+SEVjH76rrn4mKHPOsp+f/KmGdjWO7
WaxxE3qthwvimJIu39D+Jvf7J7y2kHDVh+LjKc04v4M2L18bZAyVUMTwpYUpMOCMpu3p0EhGoze2
2icjrQfcNetfc+fG8ZToUkhlcXpUhvUliCHKtYgYcI5+ERDjh19uNGexkFcC6t3D6x+kX63Fxi0G
A6cUOuvYqwdt7DCj0C6z5El8fhAYEJJnhWcVMZvt4GEAISPIjjwoJM+P5YReGHKFNIH6F1l9Bs7r
nsHym+4XI0U0G+/6oVJqfMKH0aJrMlN0jiZwk+yUyfjlrEaillupH8hCEl4hxP6rZj7UuLaYFUNu
c1WxYgeVJbllFTktAOCv1LtpDlCNx1SrNtyVmynHJSeoUodQfigWN0cpIU4CzI5EQuQeSRqz2vwE
ClutsDpPx/nBsNgHGZeF8ZX7MY3BvALyH5lNl3v+ouTmzUTZJoGh7odjW+k9VjHTW2s6OAivyrWe
9bd8mQDPb0wU6f+30no6gV+WlL9XO+O3Z8UPMnt+j5T7uoantQYpDqSoGrEqm1+Lyu+ZcuyfNXBB
+QwHNcSoyLPe3N/QzO9A5K5tRvylyNnthhrXpMrQbvWqPl8CodnLprgKnNLhTxfaMwPpeihRzKjA
nNTZYsqCec7gObwsWYpXA49oMvoT4ynIqDAqhkweO2INA/v1l3W2ncZF/fbeOUdHCNQ9RytyTPHi
RgJDA8PMj3GqEAoeyZnC9mYX9Y8b+3Dstyo9BBuSVOr8PR8xST3ldb/UA6XVNkZV9VJaqconlVZa
HRE3RSLHlnLOYSrh+pAJG8Ma2ZnKaqYk/gelL6oFkiMY6cVad7i8WE0gsW7kW7LbqOVmygq7yRAM
YNe94EP2J+sao0ap62kix3/lvPLt59cYi28DP+dRZxYRJKd1fLxOZugv+TnXbta3KnPvpa+c+TkD
fp4D7ax6/+FJExICCX/UHE3Lmh14JwvHPEzR/u4BBHBanA+1fJ/MAoNjBqlJY3oPubOsfzgTc8Pq
4szDNvrqT/9aUbG2N2V+cQqjnK5cCv+48rAs6ZvZm1k8z6T+HNsuhbVeqnA+P3KLTY595LB2S+bv
03J7umSEggBW+EYonnalr0ewn9FEFO9u4Oq3ZkOkQV2WvafDcQRNub8LSVICRPjpMYDbCZHjbBVl
8VGsRtiaHlxqDrwj0W4lEnlbjtMLqkaaa+hqD/HwyBQLz+WZWsc7GxAcHkYYyFndA3vjAxxIEh6C
4yxFJXGrC/KJem1t5KCI4PqTTyDTElHtFhdcpa9Bzh2fx0eth3VvlUIq1YOrnODLvOei/cxwJHcF
SiwhjhUUp7ct7AelrKGKj9GksvT+x6BYsOA7q/NwQbAATkOo6FVky+sCmwDZGJt8KyGPha3LqeYD
n83q5Oo86dS3GEudVvp+xKD8ppjlPw9xAdySX6LgI2RD7tL8NKTW8cjYn8xMOxTLb7YpvOjncRf5
mmOHHLmk4OVXDV7bONVD0OMPf97+onqzsoh3uVsFYeLhItgrTKZp2Q2TsA/sjhlWBYTF8KPXvzDT
7KIWy02LUs9oAAOdm49/B0h34YfUlRpI3haMybhvgbNsxHVWFm4nJ3OoyOz5dZRZr0iBr6/8dqOp
JvvYYtRg5yzBTDbS8OWVEisqvlvZepb76UNelMMaUnQZb3ZgKYKWoLB+z4tH/oj5qbT+xQv1lmQU
G+KeiNnmCUz9PIYmUGxyi+CbQjEG1g7r6rEq6w4jkOYLWGSN4GNf/z9K+zpWuzIeyYtk6OrhHIFs
BNer29g2vqk+KlmPjHLeOD7xU0KMIV1b8tVp+euUuv+vE2spA7RX3ztHWJ2C33LBmdyFxwxGYufx
+GKt2565OE21AWvH8wj9qW7Xo1RLwL90CFCRb8lgJVA0MLM2Z52mueWJLnVaWnSrNNJcJwTnvF/A
ZIfS4KT5zqUE6mH6YVfgavf1tbClcXQE8mCWSCiqy4rCIEbinSPMJOquX4IXcUX0abLeiCdiEIBB
BEus9++ad9uGeRJcyQeRuF8utj2lZQCCcxSIE8ML5SbbJIKiHXo3Bgc+88z2VME846MFu13tRPhL
WVdD4T2gUYg26yErJAyoeeUtrsD1q9p/96sTGSgIyrYhbgjGXZ5/4zHT0lcy6L7GdXRZvTBe1EaI
or/R+tF9aX2dRVe64gCEWebytSLD9AxXj5yHEN8qi6J0uaE2KtkA/hGdXBfuvQwQsy8WBbhsiXt4
Ds/Y4lJfeqWAFAYPHFHooHfISPD6h3L9Q6TE6B3w3fF9xEE9nNeBPqbLuhDMznCg5w+ybQxx0jtv
/O+j78BOUUOuA4Lp8skkUPsKG76N1f7w0NNN+IgwaJ6WXux1fs8c95gtehQuJhWxOtKSrUw8dWUc
Gn58TcpyC6RyJWLODH56Lx93bFFebgDR0dvGVQ1ubkuiMzgkDO5xsNOvON0SttGBxKQhlQSrYJrL
Jv3b1HqErsDYyZrncZZ8XNxiFyL6TqHiwzaXa+Nzwq1BLMj7ai3fjiZxs01cnQxH5N1kZz9KGQ+T
GVl+tS/aM0oIYDWOvxDo546LtVuiwLNAqdC5lkDA/oA5w0VZLN1gC58eo7E6L1B6nShSI9H1pJs5
5H/sb4Xny3HTWl9PeiYe3Woq1K6F6FdCv3+B83L3U9p9fb7a64AsZ+07TTDZwnDRUdZb9kL7wW0L
WFqlqybSoaZulOc0YYoXgVAj+dKgUFScRaUHYLL+hGXd0LFZHDb1KHWYpaFXou4PciF5CJn5MD8L
z4ic0XPQ0UUOlO7sJheWrI5g3z/AQ1I34u7ULDiXqe68rSmZGSS1/xCEzM6kiTpnEFCU9czCv2HG
7jvss9LEJ+668ZQxVoXOSKPiAOd3dxT3xrEfwIHkQ/ve16tQfsTwrerGYAHNPn893TJMVNEmxlzz
X4KJ7NjQ72JjMuSjnkVl1JL787NiRQQnRV7qkhwpMFnq1SN5peXNCT7oNYblxUQnkwWuXgVXjsdr
EyZBTxAGBr0hmyXc4BCLDZSnxQ+I9SIesfvc0WtuwXAVcDyXYBdEHLYrBFQ0ytHABEsHvnRBFyLA
2etTL9fnlAmf4tc+rm/J4dCchJWBv1wr1uroXbBiECkaKiWrDdDCyaM83AmViCHMDoJxX3KW0EoA
wrboqLr1+lLp3YoG23KJye5nouBEsI3ELb0votZAHOAC5kDyrWnKc2lfaXmSFgmFO8Yr9APLkBWm
q41P58XWOEnZJZ1GkBf7MjzldlWWaB6DL93qd+iBmm1T5cd0IBc4wXjfC3jrcAPe6rxcu81B1LHf
qL3svrpriSDln3quiv/ylw6OwEI0i5CDQfQ9RfRWskc4FqkR2rAt+0VPcySy5x2333lR4c5a7O0e
72pPST+9LHoUZdr/SSwA/FHPs8bgkZCH1xrFOKDzib4DhSJ1/DfUHnZ+0kzHF/PmcbRcyP9TC+bf
kzAljtP3FXpMR/Qo0vnFzBPGMAL1NBqNjK/kOwlzXsOrgy72stqxxZS4O7ffqyRSNFiNzU8AzfPL
Afqx3EaKVq6byZ/jOulCKO+VfTV231AADgE7yQAIfJo3geL5ztN4W3tbbs5b6wpFsUcN7ZGV9rPy
m/lZCky7x+UdjpCcIUL0hnFJGd9D3ZvXNiZReK0h6NlJPLmncdpgyxlmpbZ9kALJZW5OyXKeKHhA
WzravdksnpDZuaav3mA1L6SpFjsfN/XssvG1NNc+1tpAzW0AkcKX2TEQZuCOygG3G6KrMUTF0yDS
LMOKGn1rVfK9VOchnp+C4AEiuOaKYRjRBfiUFQBduOUOP6oUsP/tUVuLuwxbIM1BWkLtzXOCXQoz
aBZKM0/7KKnniHxA2/Hr4OFJx1w6c6GXPst2Lzwd4AV5VP1iR+WCkTFn+11kYcKC9UijDeVbA7p3
rjMtBnsju04qkAhDfCzJsOW5rImycngtPsNFAh6ac46Gv+6biifXk7wZm3JhW8zeTgUZFULan+cG
sEtRussKERvzSYquFL4C9p3jeUICeQO+YRM4uENKQ8YNi5v+XtnMzBmfnYKvh1Z+LvoJl2sXrvyr
JF05zL/4KELXJ1WXDoilf5zNYB+M0ofMb5P6TP/rqcO9plsj4vfJO/P2YPRmrs/laGplGrw6DLh7
Qz6STsz//vOqa97Oug+eVG0ofrWbn3RIOka2CeibILtGOKcH6b9bpVGQDkVGMBizmb8hILK+TvmK
iunxtZnqGqoSIzvTqMTTQm0WhSYRKq1yM4ussNRVIBQKEwYVS4oDxMvg8G1BX/fkcxONoWIEsL+6
/Id5uwqSIj3A817oGca0g0MFTk5tVzgfioQ3I8cFUepC+Waep7diyurwqZBVOSXN/PZnRFXaUmnI
MC7AEFoOumTdlSTmIh9z5bZK05hgCGCc1Yo7XAc4SP+6Vdv/DQhPq0X3l5C4hjwGBhnHmWYqjEue
2dKoYcvces7VYHspzKo6ELAN+oKqCOqevWj8N9CZJkXnGpD2oq3dR+tlobGu1E8QPr2zlvEBLVus
cd4E6Hcm2PCXADFGEVDQPevHh23lOUocwwb++CzksxWV3fZ4uKXeG4xs2SQxMvu4DC1110AvzA/W
wEjsfRWIP5/BO14MSBX+P8mqTGghW2J4rX+Q11nPfl0BGT8tbgVtYdZxRb8myYmndAmEqCblMu2h
sBBkXYN2N8J3hM6HHNKq5LxZtxbzKKgsuUrzzblPoODYS102oLflCFfIegev9fXjyLbiL0ky118Z
yzrZ5HPKOZMBKxFDyURI1/g6E2/pWvofkckIwOBpNZd+EX1Mm/Hfly4uZ2bOIKIeDe3hOk73c3Kd
RXw+O9bMloV7LK/Im9328nCH/mMQYBYYhYEsh7igA2DRTqW+82Vd11WP8ccJ9ALSHOcy0FTUautg
b8YoFTAsPoRQv+m2xPYp9nQr+T+Y/Z53kE+vxOfGCgXmN/KfgEkNv8Hff3f4fkpM9w4XfEd6sWes
YPuhUtmyicZuRki3YzUvVX2tRHFrlH6/3A+bE+qLesIreSTa4gb0KC041z8dfSiUJwrc8nxnifPs
JQ0miMePnX6Y4AsDHvcEsMSsBqOaVxgvi0UZHpuoG0OzCMUrjAz7Xu1ypfY2vhZOXtW3kOHb+UWr
mJKDGcGpzKidbnGOBt7LSrBfvA9h0j11er7ax5lADg3zTvV0vlviBaQZgpJy17q9gF0ky9fAdILi
cpjmeOpTwrrbDFlEXz7VoMXus1W/7AA123TT6QF6umG8Cj8mpknJYnHs8AKw7kV3dLyYzgFDSwPh
6he0F8kkvZ42x6qDb6FtnHazAN/1jlQ0SlT+ewNcR1onjh2QCIQpu4hJepyCxXZRb9UKQ3KgdHCT
ZpqW6pWPtW2kFdGquTF/WjsZ6QQj9yxOW0+89pcOXLjoH3PVOsXBhmE0BwGqljm4jF2x06K/NhLc
FBS5zgDFgEGhTFCa9kkNdL2As9Jq1tyeZpb21cSl3yLCRdWdKQsb49pYXqqgfROuppIxGhnxBo9C
vJhY/ZZR+hxHcD/eDcxq2H0wdJ0m3odnZnCaiGNSHy/167DZbKLbfVyCy1Flke0qlg35RUyokHyV
8dca92pEP4EQ39ONZmLm9fin9RvccxhkdiJHSQh8AjmxV01XebaofRS59q9YvUu1PMWERFKzDj5a
LR4aHvYUcR5srxL3ZNAlFhITZ8uzCg7S6hdQRnvx3VPy57187VKxv0SHcMuc4aLFDSY9c+2Cw7xC
U5FlCp11YpoFNzCLfxz/KIb/ZCKww+c/XaYR5joe2a+hnWrxeJhZQ7keR+SxssttO9Z+SIOX2lKW
Iksl89Vs6H0QFF/22+SX++etmfgBQ08ixGpxc5FT5vLDFiqKM9WmUY15FEAkEUyVNOgVRi3r4Zov
znqLv5T/XKvXI8bSbBPVXlZVZsjFEXrAmIXo10AlM6tMaveLU//vm2f3Socekn8nyKc41PLBOugm
bUJz7SCHp+fAfTvF3ltSc4jP4uNwGuVoVHrzRIOAy4eaVJhhBnBDP8tEi5Oi0x+8jNidtkNl7lLo
rhP5KXhdq2PQhAW2TikU5eVQ2yA1PgYmHyj2uT/FfEAr6wcEXt1flYtXXK8iU1o1x0gtzuI6rcz7
o6KH1LgE0q5uwd/HuxALbzPralf1wEkm4tAcloRsYF0T6GQaaApPbT+IxIVg/UjiTPNNLwon0xnA
tGH00uwuXkoczqi6n6sZCng6KVtPJJkCF/Rh6+jAHiNG99XexOegYBsLK3P0xqzbTw8jjY2P9J6m
/xMJ5b3nG71mYUSKOIzedv98mBBA/Fdnu08jGh9qzRf2kZ9CBA+fTHOPx2vdsKw96RStbsht+cLn
rlHXy2+oIFkYW09jmidUMO6PEzBlifU0P2MILzSO+84U+aJTCj+VdtS18SsV5gZ0V/uewyDEke+W
2DKNGK2Dazv+61e5sNVYLBS+ydZMQmPlZkjldCa6L8j8+IKbRiZeezR6ByqVGKiQbe3FftUQRXMs
vlyaMDwiWHdKYqE6vVu75eBhyAXMVFl0T/ifjt23cq292kZ+ADKHwxoNGYGvSrY5EHreutDY+D/2
rRr/x4xYXdwwe65JVO3dh1e6/qwHz6iAty7X1/ZJvuug63zc7qCyCmMdPZ1cJgTRrxAJYpc1tq9/
/BGGn8fdK3/LkWuh1Cv/70Y5ucRw1GlxpRtqcnNtDWDQfc7Eui+l07ZuPju3sHR5dArqaRoHXZAD
cYrJyY2+yTuV0q/kj+DC8ttHNLP/IPObJUCH3/1qN41IAzYSiDZs9paIl6QvsxrtfVG0MWUJaW90
nziZua6a8hpmx5l/F3XD1+lNlE5Cz2BOqJIl+TL67GZAfLQnau4eKkkE3SHBHDOafVX4VBaqDsqP
ciyAh+FW/8Jg59Blq1FDBN+OmqDrgYOcYSJVTk8VpAleMW/R+RioiwWuSNs7Zl99j4JTYWIrusuI
NYyvJMzKxc2EnqF4CKha/adGi/2Dq2SnBKZgGnrmGMBnmpbipGGOjdJ9dKU621l0C/vVwjoLaGy1
/X29gL0TczSHnob2ltHit6+PoxhBUfxN3g5iEHDK1zeJ3iG6EVlsRLXJahADauLONLJRkYMmIngn
nA7CFRTNc+c+kQFL8zxUUm4VAbiAB1pdvt4PjSYfKhZ5NGd/iXbFDtOvmSzWGRLe09qwf71/oht5
+nlcJFYmbhp7fXnFMEYfs4Iy2orOoTzwQLSGY3y2ePVMNUXTE+tMKIZGm+vGt9zYA+aF0Hk7zSTx
3nIC/oY1laongtKVrWZfz1/BBLNb9KrcNuk2lfVEz2n5XYNOZhcxDRifXnADW7bXtos2rlKzpvJB
D9VODsq92IzUzCSug3QcjI0vtd2E1yCydhBYJx99OPRNtRFEujEiLxvdrOtawtyZe5B82fl6ixY2
OXpPoHhb5geQNeRytyNNwTuviRnsXP8YWTRz3n5WSSne57GXIC2w5G6qk2Gd1QIQWeqk7GqoK4DU
e018qBbb3qpdqBdnViEmp/O7B7AaxjlmGlA6gjtZ3Q1Thd8zi9lEq1zQGAQWVgMnP/tApB3Oz1QP
YycYLzB1r21Jm06eCpU6VNkb53jHiibwnE4IL7kce5J8ACBdxPfxIuve6A6rG0T2EpRLyo+OxdPi
2mzv/YaQ/hDHVIyuzVn2dKXiaCiCxnS26B7V3CI6ClkbUL6PTrltVQug0X+uE5rX6hfB6k0aR9ib
VqP7oD018pQyafxLw+xyZPGZBJGjXTDtLbSffHg9N/CiEE8vcQtHmhqi12pKouaTimklQC0D4jh+
RYFhC8OAir9hdbyYUuV3kw5cpKRza2+bW8B30jt6TMsh6KOpLFcBer4sDtIt2kGrSlJThrWjJRcv
HiXxY5VCuRcJC0tKtnk19MOzU92npkAi59obNzquhIGcxoMaWPvcZtkjLQm37/6IOH5VQ9/KqrxS
lBJCguMtH5N7XHK6g1OUfPvZS2hO6wxP9siW4mh//rFgdYBqu/J2I+Oc45NFtAb+zEJjGcbrUrdI
F9vqxcLtfT+IpB+P6UHMZyrdHJhQXCLf9eMwzKRIAKIo78Iz93nC65l0FBPIxnh7lMa37px5DL/W
EdNWcVFO6M701HNe+STiniw3nQBUx4o5UZNMD61YDr1d2grWezYh5nug4mhZzRK9EYuitpUYwGaz
ma/1Evmx9pQiPLrEVfhFIaSiYCky1MSTUyUMH0TZghKY7vd5tZa7j4UfwYVIPbSNndo6uCJV0kWz
Xp2bAj3u6+CBHt+jMv/jl9SoDij+3SCA/PLFCEZMsJkYkBDsX5uviBYYwxY08N+ZiUxuItefUJYw
Pa2SH54HMOE8aDsyb65n5gL6HT+JKyCvvtc9v1pqatIvP4X+DAMSab8bB1sbHDMxOVra+mXrb843
WFbrJtswu9/fSzzUHz0+HwzX1OGk4oLS9rKw/2+tSCLQjOp+2TXBAsDL8MBAqlVUVVVb2jGYtJFV
35HfB1z/EqlAgnL4XEpaxfFpGLo3pFsPq30QnEZa4hdq4szewnvIxvSY/YNnV4sN8UtoFRCpg2xN
2Zl5MZYwSuflz9JlQ1G8gtec5WYII8O8gi+cPGErj8oYCEShjzaSVznRl8K36vIbqZEuZBVjHfUk
BoihpSi0oVKVC4XGOt1aUYbWz4NVV2qcjC8xeQWzuaj0T2GFFKhScNJD08S1NbvH2P1ntOb0Sdf8
dMcQ97AQdCqzyePGv6Xwt3G+FhCK7AmBOY5fOVAevloYQBrlYVgJX++ohwE+6MsnNSaTO3frrL6S
d67zTW2Czuyva2PKISLoRp6pFmoIX1dkXjQEmL47rNq/GNzegGxVsRTefRgwuD+hnVd6Xq39yG4g
tommmP89EXAyeH9QCOSKfOE+5BkcGmc1W48Xd/UVJEOcoFKUhBnxNoETl6rJdWVQFX57i+f54IUl
++R0umpUgCCeEpLG4Xe+Wb1lUpfcjom2Biz3zPU8BQMJdknGGeiM9ioTl7yR4XoIXxEd2ye6X8/c
AyHz/pRuSWjLOoEi40QMq8ba00fKteAx3InRDj6iNLPcbz3p84aGqXSsPBNuE5mWz0zVm7xb6e+o
vJnZPI583WDPYrHsYM78WXFE1fSyuF6mWaabjSTxJMOcHEoBXwRMAmg07aDaI+sBLJq+7mA2Yyi4
DYEGI8cjpfs/zxeiA29gHP7bJN3SmbxDOlAhsVv6Abunfnnyp5ouZOMkv4A2IvrobZJLwXw9MBKd
gOIKzOzIi//xjIfPb98yx0jUtw/dT3jSETt6ehO0MAPuGThyIMMEyfyu1Q8AGo85rvjmPSbbx/uX
Mn+5VVzpR4CtQpjbNG9r7d2ma9ZNcqIu4NuvKFX56nChOLUPRiz4NOAmrHaqD36cm9g3zGbk8bno
KEn9StCMnQ9HBRsgTsWDZzdXVkXALKHGyVUhYBWADQVrgMsisDZslfBlrojbED6JrJL7pL61PSS9
vpn6PMY/o94p5GGouO1Klgr7j8Zb4Sxjj31VA6EJ4seZl7k7/9j7JcAwsu0UACCDRJnVy/rC9sT5
1PXWlQeuUpLVbuTyU3UgTr76J1c+01SLDdOHDCoUNPiSzRO1AHjYsEJ9XeQgd8zhBx1pwuW8D0CZ
lZGe3mVRikctUC4o+zTXU3KvW82KOIh76RqsD46ntaLjvG8Mz73k7tGFpvGx4XDRrDcpa0XX6hq3
NZe7u8YQwdzXUWBsXPlbYHbru7FfPDLPYiBXeqfXxENoLiKoG4u8HRpOg6GgBaERyuGiTHD2524h
dljG2z4+stLgmeF98M6lzEbty6iszawF7fF1euHjDGF4r5QazNuJ0LmmNH//xxPutOxIy2RM2RXN
O3VzYpywPlvaeRFpOXenuyLfxYT5AGlXL5IOdH/qanzfHmjKUDKxHU4Eh2OEdFV7ZVDDi6LFUOxB
Xf2obsYQ6C/oy7Ahe1Tdlvds/KfjUua02UXGLf/t10KBOkDR1tgUGUzuvvCo8IA9qIHuGjDtgRlB
mmzoLXxNxC57AdbUm7Byw4SA6JRcs1RVaY8TiG8aaKlYZ12ceq749H56EhSN3c50m5LYCicMqzZD
2ltedF1lcg4CKn6K1zXSb4ywrw1REIpMpcO0ZY+b1fXm4yM29cV5GCTn69iKXW63Nq0HsvmN0zQZ
DrYF9RDWIV0mFojkTmI2GGWEUC488Ii0fNZqHVdk9DPbDJv8NKrNKvYgk+CbbfhMWa3YLPo2cJUc
yTPyooVoVbFotSbVAiM6nRgasLtvzgRCDt8wG1x2Ydd94cDAdED/Vc5gNi2Vx2/9wtnKOZpqkiLK
0W1PBJFz80ygQTIlJp9GBOybQhH+ffgI9w4l6fakZsWYpIPkp6r2rB+pgOu26/UfufpBK5aaM/lF
izORJIwlnQxt6K7Fkq7ffQIuuRY1WTE6wGu/hI7PgtlYyf+q4A/VmX44fJDtfyGl8eKpXMiOgHUT
CEZyyckgGAICphfx8rTnC0ihjylcSrGEVCoPUVQtLr7rTNFC5ruv6lqvXNH9iVksr8DAE1Xg+449
E/EYe3MwzGi6f0yLQiC3OIZW7eUx7SB8SaWZQdkU0NdtHDrso9RbSweMzAvBT50tHBetnNKkQ9B3
YE5D6x4GD9J7yd1aGAG8ZOF+F8bwUenIlTV+KVF74DOqzdZnvRdOfn7mf9kgkQzaPGUj3yEhPjwG
fbuDjFLoIqhWVVFb3YE3bZlJ6SccQGtKoriTsVCDl+0E7Sm8Xrxnujl2diMh7tA78O91N1gra0b3
0nYUPBDZwjfV6E1wALsMEna5wAnSkQ3mqCa0acP3OjBBObnyc3mp8KW0geBh5Uo0/rrRgTN+Jla0
UZM+Rkt2naViRzq+ZlONtqw4tDfxdsb6mH5YIHJwZCNB1KlKSmsJjOt+jH/HS/NPeWGFhIhn6q9l
4odORaMsUFpAr2TTGpiTzm0fMQSOZBlL+kWBot4vy+/CsbBroKL+NpQLGn1yg1sS0P/mYZHBVm61
3p+YT5cebY7oi+42o7pQVorJQ1IZtOhJQ6mWm6tpInJ1au9t9BPX6Pc/ILW4X9vZIycJcmsXe93d
aBFUj9ZTD+jqHItINjGEKOjSyjvvWDPae2lEp20ObzfAF0U6u606P3rI1zXJWfco0OfHRzunZUok
o+t/Ffsz3ZRtQdyAAwbwt4DxLRkn/J9mCftIR3KKHL453LziHkcjIxF/lj/CzgO1XoLf2cnH7X7w
GZfyPHVPujnHszqYHoCHOBTe1akP93mRsrhl7orLkNtvUg6++JGTOKIkazW+ZtdE9/nHknIieY5S
0M7EC7BwpFntf1n8aEmX+0Khux4MnmKArD+SCICULMYOjIEc57+nRBy/6b6oJnKBG5kSBIflD6R5
Xz35WGkytbGag1Estdw1eHzEH08XOEMY4HktQKnRueHTkbim3F/1ihTDjG6gN3KW1L1WT5tWmaSd
HDxpnXBAO/wr2NwZFlCp0fnBncNlgUYLN7gMx00glvSjo0YT8lbby0j0Pol3gHTGfeNmnaVxMG0Y
VbC7b3ctgue1g+jjjI6AEuoXRUMwzNiWszucTtgNPJASU7pWKUN6oaVWjXg1LwOow8EoSwT7YrZh
tx2O8niEU33gxzcOtgZVzBqZnRnv2r91S1juf7WiSr0Ne696QojyrcFFaaP6bDVG9t/WWEemrQaW
9Z0XURMJlM8Bb28tOE5ewPL49bVRSaOZaKWgsGqd80Dk0wc2nmetLPvn/xf4ArCYuEPJCLaHSgRS
C9AbT8DAqTzdjaoTKMoqAJzvmgRZ3RQyUPObgjnQEvzeLP7ZzPXwGXE7bDcuABllypmOgwP2OMik
iROgCnfHez8oIBfLyKd8nnSS1g9MJ85hC0yrsoUX/7kkqCZ3NWCZxhjfv7YvJSw+JuQtcx/P0BcC
ngbfMoU33Ze7LoGrB52P/214wmdoKJxr4ZjguxqrmK6RT1tDEyT6U2bG40Ea8s/SlAkx7rIV8EsO
ed3apVv5jaiaXnu/UMV2GiSJ9MnKm4CeLmfsN8EldAAzq0GP6adn6YWkcDtXfDxNLupeaeBDgUUw
OUgJTiesTXzmkR327jxStHyY1L2fIuBaBszfFZfM9C73TxzuiYWB8NuNNyDeYY4arItehT4CfV8J
Podz9BHf9/6BoSvInK+IKkQ8Smg6NUp51YFt30cymrW/UTrJUsETRnkDUqVZ38LoFB579NhtIbzW
21TELx0lCgvQMXCxkNin478jfKi7SQa8JTqa2rKqNnHh2hvjz3pgQWG+XXNFsG+4P0ajDdfcKCdk
q9AO6uJFvYQOLPwweU8N7HRmeU5UqlcnS/vKbjY1ZZkweErwYZpzVEHuMwLlWUnwDwrPkuTfmNsJ
PqcVjELaqymnffqLc7qaGcVdcwz9tZ1NSlHYDL7eCSDRwv7ZkKbCh6UXBri4SoZp9uxiirCW9dwm
SW4eBvyaj6JkLIGayrMOv1yWFsAeNqPuAsRPec9cN0HEaiklMt2wPGeOslhxJX4dIZ+jjdudkntg
czeGjYk5tO0KmCYRo7cOsYydaTxhhAw1+VQEmFC3DM8hjfg4NFbRmAt06Lu9rdqBJvqgTbNgNAD5
GFiF8JVmuy1fhvHaIkWDo69LFzmS9n5QP5CZ7tzUDqJ+U1HSxIUPBk/fAEZoJWGEdHOpJcEC5rJj
yAfaVwPC3NiAEs58GlQkl1edB18JdCrVV+rLmA2LVHt/Ve6QewVJAhH7gDPXqlGZ2GB5pwv/JVxZ
ayDSqBGKNAJrluS0hSspR1wwjP3rcK+VMefcRq6K2THlbzqlrNhgb0Yudt1dS8p5UX/6O8ckSiPl
n/D9YMS9CuYqxsGbuKARd3bL0eB++UZipIZ6bQ4NI/LsZmreotIjN8Jbw9q+8R7XSPt+ZkoAiLIe
MzfRr0n7Fb9UCjPvt5jZxthPukiatUdWTRSKlWfkMaHehA1vbUu9wYpcff1f7RZcRSBz9CTBxW+E
UYWypIcx7hI7fZD4jeSPgIcLuPVjs5EUF4Iym05XTCabhF66Q+GLojm1ilTWbLGz2w6KIt+DVBye
OGY+lTbAFOYyVAgPR/cDxC47Bx+Wy4+0MnZ4ell4hc4sp+ys3Nvx1sI82f/50dtJ7Y8MTk6bgaKO
Z24iUKeXyOR6MOJIYpHq16G4ODd7ZpIBT0Al5nEyJMSedyffi9TC4M3TPGTd9rroKPfZAwse8mES
MxSihVr47Bo2cr/5q4zLJeXDuQ4XTFMzxl6njCt6qmZctFJS9xM3dpklllD2k1iQDqMFJbJZ61ZY
HdOotnZSeBthL9W/CaxtAd+JO3IVfpPyHpDZSzXDDSSXmgyjFAFWXygkfbhKcRW9yJpST+FAHHKF
NLUqPEcRtzu9ia8JzBEiDzetia77rGX+Hdu03kDnJmQkjsK+HWdy1LvQzUpze7qf5eU+0IREWkGN
wWFzBFKXU8hg+irrjDsZMomqH/lw1NA+ygVUUJE4cXC0vk/5OD6mzSnpBFaWF1hReCdMpuXibrsc
bAkoJAJ6y4xGKaykIVLRfOYwumYc1QI3khWvubk+4QkBIk4B5NnSJMum79zHQYCEXtCUq8lDidZN
eWzu+IoNgnCCetxdKZwuUPF+pm5mvrgC4fUxJLBlHXTo+aoMGhO7hcj9pfNUWo/tENzaQOeSwjUv
42ywA41zuPlZzyB2KdthJC4mtgXk2oH6Kzgq52YWaGlLCBybx1z3FqsFTSazPF6gtfmDpDQohNyT
ogtGeR/aRN7FMjd/24GNrB8qR/Hm2oT43iBW8IFo+1YbLp74UK7gwzzdX628JCAaEvObddCvM/3f
xtK/tMwE7aEM53+q/MQ9o35fShsDE40KQUWxCidXXYh6YANC2+98fJYZhYMlSs8ZTvmCC6wCdFr9
4VHNNSb1D6JVjje+ex4U8ZdW72h3envjiZ8sSkbea0nkuoB8obqmLfQ5d50ZcSmk6URxFIZFmyou
hVH/c6OQTav+BzAlzWZcrTQcAyoQIMrMV3zLrORducEqPmIdQP2x4VcdjQtdxdyt8+23lG/e8hbM
BFdFGgZO9JvfJjFypPsAkplG9offUcS9dniOdgbO6ypGt/pO0bLvpi1Rfi7wM9cqAYwJKc/iBpwf
Jsermt+lQpxD2iNdzw+FJ1NBo8O+ZG8e0h9eJUvqV6OIz1mq5fd+9BkyD3yH/x3gCCg35Fvv4Ttb
vNQt9ju1in5ZBIkafikcbhnwpMSLpa5TMmp3gPqfpmEK6njpw3HMYt7cVIcdADT+YjOEVtByv0lF
uKgVDNxPRNGPAoP4VlUhBr2JlAR/pRcvi0wk98rWM0PBmG0XrDSPdvbM2aJAhEhgzg27f3GYllCE
qo6gZ1nsB/JxiLnjhB8U53ggmq6VV/1F1gNWqL+blK8i6l8gXa9I9uw7uO2u1cV6l6rtZYY2Peep
mtMtSmTCixf7Lb3UCV5Q4OaX15zpyP6jATTep9DhWkeTrqzvNbJk+lBnsj5pYSsS7JQDsr1p0czP
wVWu/R/JKqC8WZYvzs63QMQWen90XdAM2T31Xk6onTbqCIUO66g6IB9N8oyg/Q11Vh31gW9KpK4Q
oiCuIqshE21inAvhCQFpGZcRp1C3ejGfpOVrMHSre40hWG1S9qVNdXbJw2kMaxLPgJiOI2OPMA78
6AkdXtRriS6fBrdPEMQU/2HLMJx+mLMoNmFCyiJRzIvXYMwMGmtI7KSCNZvYSD3/vxXYSs56j6ef
uam0Xgbje2euqj4yBXVLISl4PK48NG0cpQBHBWUk88yd88sMQLjquIji7xTp3Ig2gPMFd8pZnnHm
bDUCnJQ/ef1zBG9cVxeEZ6rXEU/hX0zJILRkO3VvyXdznrSx0iXeAKcuy+0bpC94+1FBToRML7d7
IpzHy8mX3FZ1y8qTc1pqXlItJuUvSkDalSM+1ffo8uo0IYqicxY7hTTKeVhO8NgXL+FOjEBbBAh8
RwedFH3tbfTOTf3P/kqZxe/rxocQufCfdGRadnnYCoCv84FaI4zLhDWduEGeeCjavjSyVde2Wp5b
6VR8zvc4RYh+buTfUCw1+HG8kwvGFA1yRIPrKXIFH0ywC10bs6Iws8vvAB5ipwVzdvoGpOug1pTT
SrNOEDVnFytedmoMMolSO5N40Sfn2JS6+LoK1fqEo14op5QhgS24mzKxEVCmJSMcm5OIPptayg21
bzjR/WfNk5exTZkfTnC9vddQ2zSm5mXH7wPI/uh8pIB3VENGZ0iYV3eWCHu/Lb16Nv/vc7sTfAfr
XWz4yz3p7dfIZvZoSbssQfvBh0r0RNRPJHkzPTZ+rXlUaEj82L2faGfWkRwmHa+Re257iq41EWA0
cyIB3zMt2F7tHRw0Da5BnjmUW0MBH0V5HHxeCB9KazkWtDQWFcaCKjJTCCUuwXpaKwKnyyhnCqrT
P7TtH83K6aOELCe0ExQTWGlSvWNnkd+BNh1pXp4+l6CAT2lfD437Wg6cqYAgF375/tuJx5YDrpuP
M/GQRHru+l1kCOSi5ZBsyRkdzcBIBMHFQ8ESEveXkCYmjPzaYVUq0jqF/rlnIqEGmMzd7z+X+LEb
V4ZPqWB2MXKQ9z1mtOMfyxGjD840GgmZXtA/rVIkXKX1eJ0dyTINvGUUEklmxpfEoXxEQoZby81c
lNb0WDVCv5y9MOoCXvEDJB1Dyg9X2YQhNvYQG2oahnKEq4B+nPQBGoA5cBAVmDtgdtQTDtSuwfVM
2U6qYxS3Bjqk2cNGs8TefNhtt4Qo7TDIi5AsgooozqD/8dgo/ec+Zn+kpyuBvnmQznrASr/RysyQ
Ks2DlIHNQGogs80WgZrX5aSvWpUjqQ3yTdl2lPR6jOw1S8bp6+FvgucroMhJLpoQoLv4WNe9WCiy
unp7rqv705ncpSuhTjNSXxZzKTtKXMa1ehT9qgKpF+bnxmN3xtvWtYMt0zR1Lv7pM6RB2ZWJmyQs
2HL9ZdswMYUIgo0CEBRgyDjilVdRvFZL7qez9STeIc/SsseGKlNorKHtxYDoyhyZWU7Cmw4Ahrf+
HlfYc0bgwZOFRiiY1v7FQRKK1e3zhjgLBHd5rKaiQtHsHUc6KzwlvaGNgP8b69KCOcWpGlW3oRSW
+e8PWGCPQA0EzPpzu+dnoBYcRYq9ZK8K7e8bzAfmbEAxX3kKkKSrzwSqlPD5SiZHnAO5sUCh1A1W
7gJGkzOn1ccYijojrCBBXoCFXzXDGIBO+upv2t2SIkl5IEoX/jTSwl5SbREhT4ZNJ9Hf0vVeC0O9
vYAlDQVrbBL7JSz/DVVGslxbUtkwbzPhsPNxJFZxS235yFQ6MIu8LnQilUVr2PEYKvpirxQ5IO+x
j2ORTR+oyi/7HuewmoTguv3iYMGpwEssuBtoKUcHU5/HRd6fZdKeOEoxR9zk5gn+7nNPaDhrtcZG
dIaK5uSaZXWeY2JLCNd7Z5xOjvqDFUD7af70baJO0tD+6FuJYxpYvCWOD9zgULh0LRMMHJEX3W+B
QXWN7sf8LJnkEu3YG/E6IqJyQ70oYt15CCT5jZhHCJne3S4skVnW8UzYSRl4R4QUjf2LscpG9FXD
6hF3Nvm70mOV31pLiEisCEbJ1jEWuj23Av5Alz3ou9Be1aaPma6y4cSfUacO2DLaRXZ6HY+bOSd8
VjWL1y7cZZZKmdS3tvGcRmnYCSdKywxPbmeuoc81loVSOGAdzXh3DpsWhaSSYBYvk3hQfZrxDHHr
gQLT5EECVQEmioKvjGhQnfdmhP2Ei/w5++VmhIesha0bbFB52cYklgoIyaMBR/FVnurFsHbd/FL7
RVxxNmxzB/xKdfm0pbf9187dEAZln7us5kByOtdPzk55J0MjY6VDGnlfi7ViWx/s2ljlP3stB/RI
t6UxduIaU80heHbIFUX5gbEGMUCCtYlfzqCo7niLG2V727hULvMk/dJDWlo/NP/BqG8PEVHaB65Y
pEQrSzoQu8PBaN0MkIQo8pQHYyKC/PU2ZC+2byYsk3y1WL/EL+vcEjdhmhXbCvBpcnq3uZhpNxmS
gH72fmvh3VQr773LpZ1/ECi5hprF2LZt6eWqXtKrwWVJl8cpT0rw/IrSfneAsz0d0EVF9vbklzlx
iMdmdAWURICM8DN2UGyikEagNa+jCNbDoLucxQU9IuMSEQo/csxJf4hq65q+l+sevtGjpkHf38UL
/MVWp4Fp25YNazOhVp5i+YVG3MzCfFBZXbWj1WFRzdGCKZols+w7ggJ96DYBTx6tAM5tyoHhxVPF
If9e4tAL90zxvmwTqbW6KX/GDU4ob8mPHSgmeQ0CC3ddYX0bMBls5y0nTumL7/+m8gqy3etcSUqe
iu3NK1MOntZY3Eg1nZJ7mV6TH5DEtg6hMhmldZ3PkwsXpxL8BUgpe3Yvy9DAKCKtJG9+roqjSCIm
t9kQ6WYhWKyACue+g/BuioW0ZE0b5zvFRRYQnLxW43vccIqjo37xi3DJz67l5QBHXRJyNia/qxf9
CoSiqWSqkOMC55dZQuiSr/u0s2ftOCdPtwXKtTwYW3bwvqQajNxY+/x3VIW889gYtfIHyVOUedpw
veBWWBhZPSCAqtYJdINtHpRAgqIEvOdQUuAzHizgXzzT4NHPEcBzrumovSbrARvbDSSqm/aD9ksd
7WeMvGZUZHAF3c/RVkGKGC820CMvwHXXwqAStFP7oKePimrJmSnY5tBBDr1GtC4RWXLmESmAM4WH
EV+jOr6lcdy8ocbuiczf8/a+mkO61OW8SMfyjOyYr1U1qZMvlffyAFYWcDYdHSpDRXZuXBkGpDnU
jSkHS0l5wEu+Xuj5oq14O5jCvZPDQK6LSHoX4eZcvfwodCRAi9JD1QlMECY0fuu58TrUkYuWPCUN
UDPUFHO+quKuexqaz3eg0rbmOl6C2uZNFVwvEzYEsVqU0nUD6KEJ7H7PQibtLYsimFAWOrPlDB0a
8ATHo80GY+QsIcJTakdwrRHMQ5tOMhu4rfE+FMfxxGLGz0iAL2p7sJafZ7Pj5HCkjh0tf65NGLRW
6uYXsd/IkNyAYg7WfWZ0qD3ed5umwCICmmCqhwF6RX0nNk0EpHalodbKEP6BPUcH3Hc8N6MYVBpY
9bqyeU/mVKEX+FmmUMq4gpCnn7noGk2gBbMX/XuE3qVglNJbK5h/jONPiC/VD5J8fJvxThy3W+es
h5SwExxalcTw7BdQc22V0rpBuY+486EvQA75OynHIOhxJnr/pJv0ke3utWH/WwX13FmyF0RgsetV
/VYKifNqk1U/zhSezYQbcBt6xt2kcucEBuTx1sGPoHhPeW5KDUUjk5O8r1BSH0qRzyPKyzaqzm6+
dEi/TpStsG4qqp71+0oRtmbyexFYLp6IlqiCxrMA6WaUNyNFZk9yfeNF/Jy2kKMMFConJ9FJfHLy
YQ6ooF09diTWVaOWhC+mUVUQOjwvuPy5mnAPCYACfowfIn+1xSRnUPXo1+IF5qVd1vQ86xoQhR2E
oKJugbMqAC1oA2YW01YOtqDtuUyCVnzVe2qfGk1SMud1DRH1rZN9m2PBGa8iDNsUdwp+18WXlS1K
rGiV/YL9hyVJ59iVUDEnthFm6cw80baZs5YurbXIRfC254VoITcilaekAuKNNTXnIfvcXC5CjY7L
TW+hcMm2R3lgJaO0d6j8YzcpSBvzDLQWtDbnTUP1kw2Rzbl0haHnG2812Dnamxr36pVf9vBkUgCr
nd3zbd1cUu9G6dVJkHKLVUjFViLBbD7t3SnWxjyi6T9rAAZU+Qp+O0AbC0aD5fziQMwQgkn1NVsH
9m4XC6pu+VvJun8ti3A79ooAazH8N0haTHS+1c4R1VGTYFZdOGL7ncRrITw5Srv7FGMe8HTjMw5A
lBlulkpUPUGFh/cx67rSADgTXuoW8jdl4DHxsxHwfWXS9sOR0SmH0C7M6y029c4TVXVDAr3Zcxqq
pxdu1VvrB9vOSM6sKJBlbOoRZgNRm2C+Xtq9OFQ9u+aPhV9wzBGeC87eBn7v3LHrg4jpuF19FrM2
WRCmyEOnIBAC4m5F8WXktftRldy1ihGC4BJ86J05UQGKwt47leruVeBv2uGJsMwFecw7gjTBz2x0
/KOYuptoS8iBPS5uTYYkdFjHKlh+5RJcR9hTEJJyF9NhGtCCbfu1mVBJ+QfySYy0ZP8yRVPcqhep
pr4KX4A3CmfcpT4Pm96MYW8VOAX2ON2VDBHBeItSf/r7RDomSv/PrTluyBC6gUDoC+ZuREgvLNFm
MsgsF8622Z2hOfwOqXMd52IpsE438mSXWzhrSs/UdlhY40vJsmULFn3LUujegBHd/vz+OgoFwfKw
W5G7EDyxlpI/narAckv/aCM2MdpHNUFQyWANtRn9T4TJ8Y6mEkuiGMDOHIwtHZ1ywByWIHKZC0zq
r4FROvnlGkbvhFeI5iRPYxR6cb3IwcVwgr68einKgdo8VH/vNVj5Q3YG4h5ZemdMNsKwxg9Vx/oo
XsDJjfW2z4ToWCba4RqwLOIY5baZ3N8S/c+02rkbHtEfpQDJLm2kXRs1BlTZAg1e7ErLYqw8PVtc
rxFl0B9voIbtLrO7iTLLK4hGpXFQ0OFcClARppAyT7QeQLzVam9PMeLWyCi4R3E0VhuU3/hZ51Ke
QsHICHVTMkY93D9ai0EF9KjZ6X6dDxCMT5iU7sBgQ4sJ/nsLT03V8zTmcA/DkmewuEBIBvXS6kdI
gL+nRBIqQoBuef4GWd24LOwGulAah8YV4Y5JRR3bb5UdhT5kumxYa382JPRxVjOTNwRX+SfaJvx+
L4yOdyv2e1T+7NpxEa4hxEHRQzV/CxiBtRwwTfMsDhMrG1e2v8MudXDKiNAKl5h2WavQopJowCfw
3a24Qk0hPuPIde5+7zqjVo7iNY6J3Wn6FtUwrXfFw0KNrqsxWpcTFCjyXDv5Sb5kVzFuZpF4Qlxy
5QTs23eaG6VhHG5dIVzDpL6FML4a+0+LDxUQJAWTme6DYaklu6r2eKIzT3p475PkOMIwZHoqKtjT
eMTPor2d/eqMKOFpFXWShQjBK7kiP40bnhi0vhZQnareX9eds9hqFClrQ+EFvyxa2mk+UrhJqYfi
/1isWhHPOLXCq99WvQseFjpA8b2QtNUWxuOcJIhhiC8RTd5WN7PBcIELlgUEvn9YUJWhqLDeJ8GV
hzEhSV8pa/8OAZ/Tmtmeigh5AqYkCl4yG46EOdd8YqfwJcYSRZUcPZz9wBWnAGqdESnSf+SwcNLU
66y8JI0ZbBPZ3uksbpIL/9YkJ+Hx14iLTG0VIposIzahV0EF5wM5ofbZd0FUKz4zVaLvm9d/eOwy
S5BMD76SK6zUeJ+fIiamzv3CUCtCPohKoxd/j2AxHCOl2inw9fpagpG3fTmBnF5er1v+v7+ikHJ3
gqPpasLzkZ4XSb2GZP9+IJGI1cZxc4S6Iz5qzYPrxiCd6aNWymyCPXBS1EaEta4YylFC8P2zKe9Q
WTcbq3OMmLI7M1az1mbjPZM52ZeRKJjawcgabxgQNgoKSZaxrSfVeBH14GPrW/+hMVTkISZlmANv
O3sdLb+mX5pdhYTdPX2v8GQoGqIhcJoY50bNVt2SfFC+6ZUivrsBcAMqpXM+idGfBfyXqV/GEspA
t/dCkVT6CmCrV8jPwCLAdgcj8JHnqB7btcI7cmP1hSFZdd2dSY6IkUlXtnKNO1vD7fr7BylscPL2
s2MZXAcUOh1zBG7efKYhUE5uqWb3kTnD8WPomZRNGAGannkijZi3E2Ak9u+f+JT06dZdp4kY+KrQ
XKZny1bci33OhVrSWLbIspzUnPKohc93IthCihgxiSpDSP6EQ4gWxgo25oYb6ruComxcpSLbmnwQ
0m7PVnR9tX2cJ6mbk2bnN0bA5LNEh2L9eWK2Ls+4TAoq6LkX5r6jSirRvul/p5PYKG6VwaDiZEOg
QFgAu7+Do9N6iL1Y1W4fhC3Xfo1vJqljSNcVjVLsnSewOkg2Tw/uBSgZH93kUVk0Lqqy0bDG3yEJ
oQbuljLaFF+g2mkA2gbXi+cRKnSaSQx3LiRVR41TiA4Jr+GHVTo3ypHeEUfyQ7CER3hZIHji8dKh
7VMyNZjPxPgKzEhj69tL/LIvfoLhmwZK1uMzMZgJ9bQz12Ueq2vd2GmupyJ+Tz9pBkKRS5pgE/QD
QTu93/5lke76wn/r6rVpD4gLLMejpErFKrWX58l+8jwcIQgDWez7rFT4XjjTgF733MWXtjaAmJWg
EsZkKFw0NZnab0iKXGnEXTmz0+WiH2Q7yp2+pjpxlv6cxteGFoBcvVbORS8PxhSu9Aik/aoDNVj0
cG4RF3R97oY1vsJL2bFzfCvizA41qGPsVuSd4qdul0jfKs7QNhoeCnQXP7CfX1OSlgSxfc7Lv/47
+4Htg1L4O0O+iLf15knb+uMK+lWCiXTS6BKbuuJ+GMtVPDEyBUcgya66VT/9jjCJi0IotmjDJNTE
w0tXBb8XeTru8dlRT7161rfu9TCsB0MlgTfHK77Gesu8TKObvm0SW64oIwHx6j5rBR0jy1GdFyIQ
K/DjIx7Idxz3jUILcr3QEoUpW6vEzEQtAO6kIFhuNfqS96NTx+GsySNEmDA439AMxSeQiZSi9igZ
0fDY11wviOPZY0k2LsEtxoKqhJHZ6wjs+wAiunA/lXRtLF6J693+6Kq56eVQF9Pjml1macivktx5
MBdRAY9Zl7o/gWpuWVZlKFea/d7zuAsb9JdPUmk6F9qUsyeIo1RF61ene6fd0RaBZIIVGkaUiuJs
rdaqT7j9qHUe4hw0C2SK7/bnQAs4v+tKY9O6HGBxS27I2UAlf9C3d8Zduvg1AbDMnQja5ovNZiID
o8RyNHa8+SfTheh4sn+ZLlkWMRz8m4h4p/Uc4djoO34UAA//5AaVKLG+1NmfseM7/+nfP2sgWBCI
YCBSM06sIh8XpDsjJ2wxecWMonffGLyhiWbfpTyPcgQn02OAnHhjBm723FIpX7sVt+Wm0AkMmnZk
94Su4Mep5NlCSQuouMtufUmN1fvU2LknBYYbma8q8A4fw5keJOZydf8o0kKaxrKDcFuxUu+vwD4I
hNaDaebpzwapFLWxBwgsUGoOZmDuIBWVzMayxPHiOwSoI/b/j7C/lCR4ULh4+0zwx1tcvy6EWdW0
+Atr81n5ARn3S5K+xqmjLnnUI6uF6vJ49cFS7ySyemFrpu29AESqoYeEgNZ1tBgNmi02wrZIZDTt
UxdGsaIlh1AdlUwgnxQVkR3cirULdk1UHw7Nx5lClHjE/Cfr9WPLuW9rhl2Iw6l3xmqu3l0HuhtZ
MaYZdL2MGyFCKB55Q4Pbmzyf+suj9l3EdsoOUC+vRYyOEC+zHlS3jQlmpmfpQzTCni5qSm64KX/k
hsX3WD6ahUhoc/9pCpASJzbv4KpJVCJp24arb17azWGghTh6njRdto3EWip5jfrP+qQWAZg5kYZD
NN38eGm5kmM/1yn3gY84E/H3fDfkZLonXa3bPcWIMHainngs5O4b9KusnlWNX5XoWbuN2yIgOG0/
UYlr8TJWRu/dmM7a1n2nHwiQjaz9I5PjDupTjN5qv7/6A/QqrSlAYFbeKdUXujJKSnhLLvEAz2EC
gulrsRcSU1AIsIMdvqiJ/jCSjz4KQ9THTI6L/JN/KlRRCRDW+AwQpWeTWUAQBJ8n7xyahrVdmTPV
mYHANOSmvXavUWgQ1KDqljCO2wo/DASXd4THtsQuv/ZLX2ClWS1otIlHVeBrtB9IMTyEhhSQmSkT
QJkauiOdDaxNwH08/MFEF4RMNZZYjYvYtjv6OsF3I6TTiBIrHsiySROebhdBVEUXy3uj87vpm6rM
qUXRWXWrKqIQeSg8KrI+it3s9xUbNWOtMLLnfW2jcjLtTgos/Xr3aDYHw2n2gpTxiWpBAaXS+Ufl
Afn08xUIoRlSLNS36y02U95PRUyCLRX5Oke6YuHBwK6ugL63V/QTBrev9TbKC5BMRzXmrCo4pn73
KVatBhO/2uadBfulzXoFAeSO72ZbK7D2N2lGJNF05Bi4a7+Zma7lb1j2/9COUEZgr+6MORKucV+z
FVv7w2CJVNpdU5CsZKsCl1YM6lmHPjOKP2RN06q2/HaNG771BEAxliJHci+sPO3bmXm/Dx6XtTBn
YNZ7pTgZsPp+M5uMpB2j00TKV89ODM+CgnwRTDWCsm4ZqjFTX5y4/m/nGZ5DbHYiZCer7wPsJPiO
TWRDGhZ5ZAH7x3/MVk0Iw51X45zvvUFIF78Dcrr9SH21oFXhYP+wTXX4jbDO6GTgLVYeEO3PKmiV
x1MuqVSouMsycuHHnSz5iXhMvZfIYUqmDZ2gPgJPqeehIJtZmQDdZvptE7bQVY8i4e3gztZ/b/sB
MUyavxxDOdkH9QXEdC6vB9hY2lYYyzzecx1viBta1nU+5AoOSy/rGi5mii+SoExarThx5KR3xrCO
YGlMJBWVSZT+t0Qcnr3iazL/L4BtXdHz5TrPayf3/dY+r1qeaasPYekQfzkd/7JrX9W1zcvDsfLu
/CZB/0dImiKgPS5VOU1fI2rR+Ve2qa4cZBSxw93X3u8rZi+SUDTBMqI5NPGrNjo7gwFWUvs3+kLW
WdLZiwjvTH/LHfcbdIHolBiTL4onu0iWUIN9xJF3p79dDFEJ6tQ08/uv3DqNgr/o9BTPz4mrh3A9
0WbHZwmpGLg5vlWcSb4Q9YjtcFYa1pms9yFlJwl7qQRlSfbOpUYpTXyQsapVKkwyUiQn24Ihd4Wh
65LMVydXRDtz6n/XK0ebGZQgq4Y4NTk5Au740wXIS83jzNN5TvTnWSCZ+2WVUdwjzX1/rts4+ueu
+2YVsqSgqxpTvzvVOIXFY8aD+N6bX02/y/V/wNl4Ux+nsFtzD9dr+SwyIDPdMRiadIRbkXQeJcZC
iBDWYRCHbNi0vWzbzAJyDcYWsV/Z2LIW3BO2ZXKmiq5gRNILaDfthVo6GlzedPAdetbSRaVXk+lH
XW8OPD4CVrCwy/165HSSAzyjRdE7IS0o82lfEa5mG5WY8KTyMa/aj+3rS49s2SMh5+VFNXYvjm7S
egUhlL0n4pK2xpC2WGsRjsZHYfrFi438SITsq1ke/cUmZQDlUXKMXEvo1UzjDt82JShjM7n3V4QR
NmUPUWa66PkouD76Xq8NVVAf+R5sqqMfsK1PuaNtZge3f6PTb9/YJecckc27WLibFqrdBV9DMduW
2tU6uRw8hGtZ9Y/M7BtTC52tuN3+PxNq5HE6+EgW/INLvWYq5g9GiPPWpptW0ZFahK1CdVCJBo4f
GN9hc1ozCjkjAqFeNvl45K5NCfd3lHrhUIfBNU5UPy6+QuzyPgAzfCHQaktZfJUri5OyVFg463Pk
X2WmKdDHkCmTMdjArz0WdcwZrGLPUsjoctFnD9s/NToCd/RSN1k5aTwZuzv4aHCnepueJ8QulkYm
+FbK5M+2XCL7MB4vxbZ4DX0yTnBNuuaP7PtamRPWus9gaYnDEuBU+fbmdNkGOgLSiyn9gc2arrbG
jydRl3UZKFbz3+GZm/1HnhcEeKtNyqQFL5VycTWdSeeJAA3aUgb8sJ0EcE7n9T+sDRF69xbAlOxi
R35YLQrLc2flEy7+tIhwhpKD6FdOuoVhK9ApiC38KJqn1dsk0PkuBzEH+0SHMpgAHCBeY2BWhRd6
YHTXEQZ58ZIAZiX0TiEi+dCVhvRNBB8LtWmInsDLdPOa5QbvzEoHM/lGiEAN9ZoCDZCEGH7O6YsZ
FyVDtJ71uuOxqojPDafcRbiCPOWsjAsgzJftQHiEBF1TR4RwOl2HrTAABlJDd/czvQP9wEEZvKsN
5evacd1MoWNxq4CUoKeRcV6d+XZjpJ6Jb56dMdb3H2dYg+V8cMG/o0lBwqamLgBNinvog8HWve0w
rRPav/8592sJlegkRBbqpxYXYibJqsc3wW67KG+xhbqwaYZGMW7jHF4gxhS5JRyXgZ178OKMnsn/
e0hQYfisGqK3liv01KZ3gKo0C2jQ5CrJ1YpTHc2DgCgZiwvupNDltWeQIp+uZU08jhIQXXZOc292
CoGjSCaiLbUDPhseNqV37AX3C7zsDM+UbgPeTdXlt/acRvuCMoUSd5zWogXcmIvH5017zKb3XdrF
40YMf/Nzps6pJYKf83CdGEyS0iifDLfhcg0/mA3Q6w1vnvG14Grm2ueRcIhKMAM3pCRi4kPtAS/x
go3IPhY1ufwzODNEo992Vc5Tu9g9GE3jOKBt35mCo/g6A9r55kVBknwsYHqvhARO2OzDsC2RyzMw
/Ck36BDzqoK4oCBuP7kE6d8FLVyOANtgUZvSiov3hMkCIUgumnQ5nLBlW6qg4mxkFe69ox+mseXp
EjhnEfsnSPZcOUsY4OpKJTOnr7EoCFpZ+b82jssoswtD3hmLDMXSXNXOoMomO7MhqQdNwBvAYIsY
u6kVRvI+XWGP0PT9Oi+ZzxX4/6qAejD0LfisdGd9jPobwo8ObwHXxFqnkZf6bmTBC5GjlKOy6PQl
KGZUUB505/cXAIJQclouopl+k5AwQmrpP3GtBdvtpXUJYOfS5dnOrURz/PmGw4zU/rTtyawPMjMq
sBdEUj1ENEhhImmf/xIwDxjY24/lDye0Un5EzVX2+iPCjKsTWe6EYHGwVuoRxKGY1zQddlzlzckj
Qtd+v2o4+Aw9iRLEaYggd6iZv6krdF6vSTKWHDFc1Dz8A3jvtoNXAtSiAze8EscCY4mTiyVgnn7G
UuLbgVqwPGT6XsYWjG0LAUj4W2tJX6bz5j6mH8LDh37cLtKkus4r1qYk27D+eFzwOXn1gE7+FHUk
yijajdHmwcX1kKUhEsb7Xty0o27DgquLyMdbbSfDdZi5ltV0BNrVNXlfdye9JL0uzX2y4fGtLCeQ
uLaZCyQJgqEtIgq3JRVwnzWzXIMnA1lXIPLE/86V2rSFeGk3Zh4hegtOh5dPmhM2El7S7PEUAAok
zKeB0bwjYMrzgjZ7kOLzj3/+JRCDXCdq8TEsPP8hrMsOWcDVr//MESW83dSkywwgirK/sBfZ7aWm
+H/ha379yXzOt/As6mzENiGSHhFxMOXd3xAWDoLaZwH7709wnSO317gSLWXrUNvDlv4j1xq+xCB+
w79Pu7IWCXq7JqaJeWP5gh0G2x+9gM24Yd03rj498HaNO0PsLpzsnBsdgk30n8uJ1dfPzWj0xuT9
KvE4t3b1/UH1070nwt55s+alu330V4kKba2EZNrmINAqbpMwaJI3b4TmyUfv6DWqDFUczGRoJVRI
ynSDhRzdEV4IBKVEfo1MFczqWcu73RmjR314yTZSoK/MM9ET+tuB6VjBQZPay0mIkG5pSxy5F2m6
XbKfKQ2S+ZGYT4AuOEN63X/WS99Ow1jE1M/lDbi9MLToRYbyfD8C7u7lpifvdAmYpqWKXkD5QmUd
88I04br9IJ5eZx9mZ/ycOH5rqNjREbfHj4uaRXtFWSBloII/DvXwbdUdpbZpsn1MfGnOgeBE+jNo
HSehIspT8ceAc+zm3dYjjSSjW4jVW3MUAPkrtnWK/oGo1ABN8XBtU4wg0gm+9A4WQPtB+Ln3jmPM
dfI15iOS32b1eywIsbGPyT4C3sM9GBbN2gWQ+uAKcb/4DFbn7EzKo0EFhDYkpAHJNQIw6yrz/+cr
Gs8/Zvkk34PS0KQA6xGgvMl2I5WSrEtkHBVWv5vEobehXNb59gn1SpKJiQX41cHSM4VTSq5fkYZp
ytJLAprISUZ3Yo5fyhSmpfj0Br2L8wRVyaI4xwCSMUXLXNW0ceXx0tsa8TFOTJyX89RMoGyb21Xa
O6e2b2i4hW1HFDIEjIOpYP0OvvcJLcdoibQ91eOnkwWYoe9Sq0Ru0qug2oK3n+57Mc62wVajzIla
0j9zWgecB05lEBKNJwERDzmf4y82m++Npzb2YfKshmCR+8/0EPHiwZUtJETw0krafBJZOjG+igO/
NY6A8bjxKwRntlaG/zDb0JndZmOn6RvNbuw5m3G1msYd70ZfMgeQyQsyR+p42uGBc8D2rD1YUFF3
NSCbfGe6V6PYvhARZNaC6PuQBNZAcNtJuQr5aPs0Sx9FUM1WfHkJojlCvXQo0d/6hTYsFZCaxK5R
+GgB/Jh6heKbO1c+L7T+WcAJpkiKo7Ziafc68M9zhxdO8os1MNwWdo7KpSa/4uS0n3SkCCZnkcpj
OKH0QTh/Q1icU2gDyfqDsqMl1U+8ysiJ1+Jgcw42tE18kQzdzM8z3KfLLJlqshafFjn+756hu6C3
ta4pnR9m3zkcOIsuIExYem+I99ft3J5ajyeGnwpR1Nieu7yTMOF973R1uqlidSI71L0GvmPm+000
iwbyhM5Hs1dv+9XIQ3ANCynBeF8OT4eYZT5xHefqXfhnk/863CFh+Of5CtDX+sfRkC15cqfkkUmy
/H2Cq+L3X2h7Tw1F2JhGhmkXGJ3dCXcqPJn/nLbYXbdKHMZnzfOIY7cLI5iAktHbXg2icy6+We5i
Dx4f/E8X5stz64ADmoAZ8wz28LOk8HUzxj1sPP1FfI7XJ30OxcHU1IaUAPetLkI5ESQHmRVE0tRe
l/ntjabez5KpiPaBVpETuS+oD8lFJSjYoZQNcPV3VTeLXVRLNNKDG+/PSNXvCvZ+4dxhNxaplDcW
AwNlIJKrcXuzC7lScqPqWPAaJ1a1Gz9r4WttJCj7DeVZyjeUmFcEKoN0nz5lkcZvulcuLVW7W4Rl
utH6mgqN7wrL5B0ATO8UIthmIe7LzPlQBttj3gbc/xeIO9J9gJcW8xnX1O3knvbWKUqHMPV/4xST
1d/pkCLKFDoBUeXK3PieT+oXc4Hs8WS1O/Cku0B7RByMcKSVChpC6T5gkX/LhJpFcD6Y7Uy2XiTz
0GUII/qXP0u452d4LIO6ighhSSAZss3PgxjQ7MeUnJpizWDPMwm9iIi76dAV/r8f5kbOG5KJcB3D
nQ8iRi+P7DnGj4mwfVg9zzQHzZa0TbKNpGeAA25JXH3A9g1Eu3wuBQoBRfM66gh1uAq28jv08tJQ
WWpWQB7Zrehy5cw5L4LAaj5IC9qnI/y4rT90UA+SXeVVrXAQf0ZHUPbeuT6cStm1Eg8e/sUCZ5Z5
w2MgNOP2NWM0jmoqxlg/3eaes1djucazPOq/1ZsAxzdbD1MrFTO45sRSbMQpuYYcHsJujr4htk2d
yXyxsdj2gvRWFuFwC72me18wzGCkdQDqx2W9KmI4tW1LLM1LNkvNzSYkX9/zBEP1ij/3pctG6wrV
9n0H7AM417ik3XPf0GNfs/5F8VP9zixz4pdLWonpzQnnlmim/1VFE1zK7d9O5/DPVZyHAn/XIi5n
16DGFVuLTjrO+/KWTEogeY6HYw4VPjGDlkLAaQjzeTBh+4c6oygqaRhPQnjOWj6A+gl87YCeoT9p
tHOuyrh+peSluGChuI5fW5+GMF7DbqXLxP1xtWLAC7h6eSVIkbX5w8tkWNQp3n0ILXY+wOONVowT
oH4soYHQ5AaW08WfoC3RoUgwXEdQmEHY4RF2vdn3fdRXdCYwjOqCkYNwbEzn80Byu9d67/HK1+l1
4+IjAwZ76T3z8s6oB4MO0wfFlWVmLKu0d067C9VSazMMAndNho2M0bNvOrj2Wa8MfRhdooRwSD2s
hEbTJYvgFHTqjxaqKT2jC2NsOpXh02kd/z5ThlbYu5GAOrKQhO4YOn4VSHYi3hvQpPUHVpJlAiW4
AyjPqbk5XM9Apu9dSo501MKX1XQPuQW5+IAn0v+nMDtLdR6AIwPBu/bW3EuY2BYQk7HmkWNjzfdU
ZrPBIGTOcEJRBM/50RXiB42VeUduWAaAf8xsvNKF7W9cg9sX33VlSyaHA5dmFkZzAit3pi3h4gnC
zP0020UT67/TxEAlzSeI7Vc6e7ZZtADotQR+VZ9/Vm82CRrEx9GtZfhFfagD7U9PLtNxjfxbCP8+
XIxFhKdpt2wTpTax4p23GEOZOv10e0peOj117qYurNdWpeK8sJVWUt8uMV9e/mrJGl4gsMSlvUER
Ph+2/6yjwPz+lCgFzHYH4sqBDarEjoxIwI5eJ29ADXp/1/ZVlS/6XadoR22Izt02FGslVZ1LDozU
vAmOZjpCryj7zxOUFWC+n98t8iRgEHNfzF8AXKgaLMUXgoRH2k+x2jIyINM19qbBe0q55wXhvvo+
/ECM3cLHbRucQoI6ByR6fYceVWHaWeRfSt3I60hk4nWr8c+0Cl25wluT8W3l0BGEZJAr1mb8q/Lb
+VvfHq5GqIwHulxqihObaOwiLlDsZ8B+K9HN6QT5E0vR1BF9HyNXom9cyU97GD0vlhhX/ksFLQZb
deF6WzLVqIAtj5W9BzDQdj4H6wNMO/6aWZypoOcYMd/CbD+Rqq4SqMQ25j3WHtlqOxxIGVnIYrdN
fkoIPDnJ2/a3ULjVOoS2Hm3L4IyE5EOvjZqI1AQrL/Ef2HVVGPMNFVQGtcm3pGiFvRx7N9nF+E7I
lrfpdRzzvhZmMW64aMxRWRUgMC6wZJ4WiAP+Po3tr7AgoKspjMHIZZVVJGR6d/tj1A3YYwmuK1lH
1QPpaXQFzQf2kE9njAIdCuMtJctlMBMft5uC1pMRhryjSUIH4YlxPHJjhc6T1B0Ghto+lJBmcQ9p
y7Yk4kK8wXlXoL1H86YztYHPc81mOVYCd8c3+sWNI4ouGnk0A+v+yIqVI/jhrpgSQBECzC/URAuX
RGIVMz2Cb3iavSRnVjxoWECOoEIn/ooWg4xLiaTZOpjVGG5trJoyhHbR9sG5vEpNxMPcS4fby21J
/+gX4LznSzthjBREzNYkPGD4yf3JGGZwV2AgEmzRsPEyfmrB7M1Z4inGEmvftTKN2evh5WSVnETu
gA5RaYNsiN2kJQ+LVD5A+oYO05Wqxc1YjJro6nXIBp44zQQlpFY2mPkalRtCm52pDMgT1O4+q7Qk
VJhn3qZ1B5AoNzJmN/w8P29AJG7+yJ5Ghtq5EWMaqfQ3h0MEPYRw4IoLVkVa2ilUNpZtJlOwa9/Y
GvAdqxJeE8qb9k1Rx2mEfTU3WkwAkzJbptK3ewrhij5Re/MnVN8uJZLYx2IQYH92PPhMYlloN0yJ
fIFr7UC+DAOjYZdS4NSHl/71CLrmEnj/2cac0zVPJhRj1bpdJa9Jbd2sUauX+6WF1bicwg5JeMJ9
35K0pHHkvCxw2Xz4UwoxsQwOgGUD6+Ujt+Us7EMlpRQxzlX4DhcYW2hGQ+a99FzssCIT4FmiGmXy
RjWmVEdpESvTA/1MTPVsmzjQZwsHSVYvcKZWpgfkQ7VoAAu4wRfOVMRJKTm4QTK4akeb7F9wa8UL
w4OiHWlaeUe5DVTxFxamVbWbopVKUOKn88EA1N2OGkB4Mqjzr84WPtXonXi3BK0gtpQDp7N0NOvH
CfRJIMsceQuuigcLXkRjM+B215B9jPhBo77xj+9qS8a+LY2yFsHcAyNVqnve8RwkdqOvGqt+LbQc
TKDgh1qdyhvXLk/r+Xb+JGJalDAX7HHr3WYAFtzwl0BY7S0AnY/Lqax/yCr39nI/qnoA/D8cT1ff
1+DWA7qcuDk/1jwO75yNMalhPIPNnQMOHB6LDAi0Nsnu+MaaTSxqnCMfetPFesVQ9TXa3PupwU10
kEIN5s/CygCzSL/E+gFh9HYOM7pNBo8yhmmoKBAc4eC8yg35QONySbDXzMzG8TWGOhmrOmMeKyLe
qFiBWElsDtvNa+BQjK6JhOznELvH69ppyx+EyKHmGXIYGZPSDmEsj90ETgg3MidEa0/pMWpScAa9
Tls9q47q1rUy2jdznEEYn4OS8XGl8Gbzi9ZcdHg9aOkbMpJNFh6L5dbjHyQsGLNewWPmDDHAB6RY
qGZN8DjhDaipcLHUTz2NXa4Itg96tNwVZ0tBbzvWTD1hOn1nxUUO1p2W/LvKSdAOmLW1e+phj73r
JwiSSyv/PppahJgLeEec9Z9Yv/WNyzBZirAbVKakFWYaJ48OcHhRsHZPdE7y7PlslwN+sQnxwCnV
vS8fOW0sc5F8CGWtrQvVOrTcQBbI5RBlLOBysG3p5siJoXhBuzciiGEldF6ee2sjM4vaFfnQWwND
3A6T4Ue9MQbfjuEj3v0J0LIAdDyZuYon8oKrU11qze3KFR9PD96euWSz4FtYzXLuFlydskyKiom3
sMpV8O1b00R1CdH7ot6JvHOPE2WM6cX7q4ujgc4IPzPpBFTDA0MFPtIa3VdeZAQa6T0OxjeHAj+Q
+NwHBCG4+LFys7TNGaXZeYyAPkReyZScZp+Aa47MBRzXzf5EQGqPQiMmMaA4xGX30XPX1LwB/fqT
Z94w7TQWRy9c+08hR6lVtUQRQTuQIdEVVVakIKnuyxU/f7QZ+lqjwhkuRu4ebssAzWw6RXHpptV9
nNEdeitfJrT7w5M8axuS4uRJkaNZJQGlcXI5efF9tlXgFqJ6ow+WRD/2RNJ+V/6IJ1W2vmUT0SO8
tYCbt89UNMmmffh52uzCslCjq82OqhRa+Mv6U8gTwMg858S894mXh6oV58ukRp+C/yk7p82OuIgn
tbkVFzcL8PpdW3Zj86lecYm5NGVmTJXOqu9Tc+2b2p5IClJANWmtLdydSkPcOIX2rpgPnTs7zO0m
j8/f4UFnElJ7RHf83w6huaNRq6EljzIEpnV+c8bOoEbT6WJhci4T8efNR3ajL11MhvFzLt8mn0IN
DQDpxAOaclmhpr3amGkTGDXT7ykfjHMtgsSSLfYBZ1SP+CLYT3R1QViuKy6fRoo1Ncm0Q06vUmFJ
g+r+KHzkGwrjuaDTqjlMKTtx/Ov4q+CiXSob2fSSQPjmH38EeYVQwPOa4qdsrd0eolIUja0N7AFm
FJi+XBgGUPeswMMGFQ/UDpmSwMJBBV0nJMuIPcInRSSDZIg63lT1ze+m498cHw7c5oRHcu5v7CZ5
QDovmnH7p9g22R80sR9vgdTGf/4P0RTHXXALIeMI48CXSkGoN/ZZ7YH7/hcvSyAUD7zB+xOEkuR/
HZ6T+ZSCd+JuoH57kp2ykcYZWKJe5iQDjQki4RqkBV3ij9vNPpR76FYFhpoCE86kfqTvR7luQH00
nGuBZiBYgG5YTkxEMz3HGVwrG/ev4VluR/V7undkc0OU+ojm9fKca6tu+1h6DvbUf5vUC7+NI/B3
N/KpTldRfk2cM/tZp0cfDiaw1SuP1HDNXSJUUWXMAB8Ahs6IIzXrnHWm0GbwSe93O4w+iSRg1FKw
C1HBYppHPJHeS9JpsRBEXEAbmF9jeXsirSoYI+HVe7Jn1NdPTcG+US/n4VvmVthBAliewWZkE+b0
RYw6Ou+9WOCmZAYOphK8v+YSG97yOwfyBw8e8P6bi6+Wq9b9iV/W5vI+wzgtd3H4IkApuVx+JVmR
QcpXnWjmFt59xeOvG7pmORjVaUv4SoOTgZVn39hB7id0mTffToHjno2o5bbKzJyt72cbel4eZlwu
4oefg8xjv19FreYDY+0HHa59RGz7U1izCp87c1Q9Q3DwaLutekQEx7abDyD5zTmYBrExCc/3WcsV
nRQzFryLOPeNLyUlnCrnzaKjyle7f+QZTk10bKbV/ERKheWUGxO3uMHQbSkrNvXAGNesQBT7V8Qw
eEyKQcLUpn7GMUWmvO5YNDrOYKYx8mFgjCqoG/EjhB+onVsOqAsJecoByQ/Ro7jXKELEPyWwwJuL
zs4tNf5mnvTy4aowBmuFRMzKfaykNTthzmAPuo0dQsEY6tqojfd2/eOs9NvtdXbRufTl8nmGZ0lG
G5m+g5AwjL+vDVhe6QL2NVNGWBJl/FY7dv1wlchVUSqg1BkhsJROkLac5GbZGvCp/mnFWnDo9yzz
OAuU/sqyZWbAP4/qS6xxIOAGKJxzO9SglWC50IarVI31FKH2uBCaADEMgJ2fswwJRGjRxThndlvn
PeWBbSdvc55JzC96qrW8ET88GvQ5a5WVIgibOu8VQGP2TqHOMtndiRalWoNzVaRDRuumrOeVVejT
YSpFL/RSPpij4xXkmr2UtUobsDWar7uTqgGuJ8lGWf5U6GbVoM9PLQC3j/AQVva1/vOAvnwu3d+W
bOTz77bDq6KMTI6Fq0zdP2IgaQRQ6VWkLZYs3R8RmDu4ZI5XV2s8wWO9L5isdoqnSC31EsDJhshh
KPmQj3L8uBKQzDdNVc4m6/ZYAcgbbmpflamPy9iHtEB6NBPuLGZrWLkeMxrUZCxSeO2jMmhqkZe8
OH8rZkS59aJrKKF/+toYLT+DVBo936o94XVQFIDSjZ1U5/somsns6FPqD3UZV1xhJ+9wW83l/hQ9
01Fta8L5hHkZhSDyLgyCnw4V4iBGBDlKZOx4TjGzWgSNBzhQeD8kMSl1G2N6h71Idh8cn/p+H3Ts
Xv725A2nM9WARp0v+dYprSpgyWXt4Bv9q7/gQYUtj/W5TFE2Bm6g2A1CJ4/JvO88YqDKL7jaZ9p+
0dXnNavTNPNe/U1qvZeqj3UuSMsoFfsSgv2Cmm8QasFt9fiS3EpE+RpZGyV4KhwSOZVXdlL6HpZI
JbjhdVqrMnKKUkv4R1k6bBQa54DfTu3sP4VR0jLeQLltgmHt+qTB8BhbE34yoSuDfWR2HFMFOhVT
9KlEkLg7m3vzgKJA6/DN7hqmhWMwxW9mUI5iyXtoP/FtufDmPE1LRaxqBofTL8p7oYvITa0wKS9E
68OQm2SPwO1ej3uziw2V9JIrmip7Y0OS6Sgd3rBwWNzk07yzsRjEs9X+g50Py3OvBkZl928g4BP3
yhTQiXmRV86izhiV7rW9yC6t/1MVgMaw+ZzGFOLC9gSmacSGWDVny7qUPfyelG5jsyrTwpfdm0+X
iKRwUW/B1nwd7m3twmjBleS+gffW23aajelWCIfhvol+yVDvcBHbHHtcIgCanRu/kALFBK470pI1
J5Bs+SFcop7N2GOjWB2JL+luPpU0i7En8KnUAAgW/hGMPkLjO2W5AgA4Qw6c5y6MRnPKW9GSZl4u
J9ppSq79pLnRuq4//qOMw6Xs0Zh54F0dlxjlrugIeYEt7qLQkOzjnaePZHeeOLw+t++8JKZogbQl
fa3067Njv0qgQmuXHlz0uyNLLjMtBL6SttEtfyJkGEVVDYeu+J5mPJkScLExoeslPOQh1eW6FInj
1m/gQnVZd2pZrvKzk/45m0LEDtoUKoWRGtcxXP5VZKLUOfvTAW/8af4sxTRfR7Ua+VVYDaE0FRLI
wL8EMDRmuH6EN8l/pwKkw3jz/0DCh5OqQuJhgbZqejM1dg0leIjJHoRQs805ezDfMnQmlTJVWRD6
FAs1JqiuD4VHa+Uz8z0syfQpLG6dCo3RtkbgJGtuLhd/N5ajdBIke/Qu3tQK6EYLKmZEipwq2o03
Ovckizv+w4X6HT+3XcfYscYDt4YYXfqLXm/1mv8X7ywSBzlXjvcNCJKGoNFAl0iLJ4JPkfguz0OY
CHMYBrWNzkQq/XX7zURG5XG4boDzq2lXZmETe3CDxpUR9z8wbuiRe/w5TUmbm9gKT23a21xlqDMo
9f+9NMW9J/LkIZbc6a1nQlkLGSDJgl3lD5qlRT3E48VGAWJ+fyYg4J44A3aqM+G2c+LY2H3TuLaG
ZZR2b2zeNITbHetN5ZtoNSTvu18yP6D0LsSQqslWwanaMIb2pPidq2xXDhjBUrqaiS7D1lifqRtD
WCVcUs1nROwXmRP/nJpb1/ZW4ZNF06v+gaAcwaZjqXm4oKJNjJgl22mEp9CfLjxwK3X/hFUEuvF2
Re3s/6Y7fAXgxN1YRpjABr+zpSKHJl8LtMCOLfxWgRx/iv0t0MsuSDo9iKa5RinujDM4Pi8HI3Va
p1oji5gVwhpf/hAl3eil0ON4SACeNhLR/juAa3VIDN9lB0s/51YMN7xpy9jTVmXvihFVeZj3NaSS
njTlbd6T3f555nN8+K/Dm1ywAjf49AxHaVEg+DhY9UgTidrNWf+MybrW5ND80ZgaIRqTeOV6DgQE
S+eik7E1GunXi6W/ERi03v3LP10a93n9Gsm8OhkI3WNDI11T2SxpJ17s4wQAVi/QXqZjQT4rbp/o
OFiJ/avEvbK7j3O6ibF5+QLYRG2poNpFGrhlM8cBzpOHChIAQK+/TKk2cU7SWJhlehkgBoT8yVp0
5Ef+6xbErikT46QV91lqTLHgnozOhTfaJadG4ShhLcAx1V2agoCH1VxLk1wEbL51OqCxXj9zGWir
sbTtO2n0h9ucmaBGal32Xr/dEe+kNdgH2eZyw5PwqXVAODT+EHldA25DMr+sGg6cmbtkZI8Uk4uA
GatmUyadcdYDr2yBQkKmaIk1tb5k32tH3xw2RqKJOhgupVjdipDKy7JL7zIAWHjeEyt7CSHfZHvM
VJ71hc5Dga3ZmtYQzHul/lG5RafXhplizs7WN04roVXgBgfEjS4wYyZPnIARfRJdg/Yrt3gBmHhG
ycC67khZe9Zy1zuTFSu4MNNY/Lz7rOmPznUchHps21Ey8ydEE5uAZhQZcxA25O0XX/0muFKQekVn
6CulZrBNX5YQMLkAQULB4f7F5fnvlMn9f7Ip9AA15aENeGAr2gFahME9UkVn3LF9bFMbN8PUIyXp
TStN3xaVY3zsa2OQcnnvGNUXZvVCkGu01AmUbnRTuQa7w9Y5aI7PiS1Qquzz8oB1mkYOQgIhmMpJ
AzGjwXQdD5Iu4g4USIjMkorH75FMFnNvltBP2e83YOeQSRxo/ueVFGolz1k/QR4AsaaoambKbb5Y
yXAxJbV1ByKAvM8X9ONeqx1kObFS7BpXAxm/CGFxfABXCGH4CacU6v4kYpSuM58Ok0aJK7nSa8lL
BnpzYV0aNHA+0XUiIvh7R4abEW3QpCntriUxHNXlbesHj3GloUgo5DB0wMs9MU+IMAfIIDRI0RIb
iBu1+2p3IEe4Xb7aE+rOnEnnRp+fwZg29YPWlWfMJfhmvxQXt7ZdFDH/ZjVfRjVlWHPsj5Qb5ev3
ghLW8Sjh91odI0RIuguoJMGlvIFn2sFWgwDYe8HHlZ6QaiRpD6r7WfRKgP2OzRotdzDMbDIeIzVZ
z8Hl+cZDLfl0HwQJraGG9glERARd1d/Xs/JU9kbhewAvvOltL+zjgh3lcNwmg0nEvyP1N4EvfIp/
3ILUEMbj0ikSBKc/Tq4+bZXRBd7ktclLheeTiWMlOiqCu3z99VPZRo+IaJD+4t6BZg2A1pXWJ5L0
TbiXdFsybiN3NVKXRO00Ohrslxx7MzaWFDul1thS6yOGoYJmbC8buwSC6nxhbD66PanghCcvAOIm
9RroWT7/Kcerb25SIuphihN+p2UfZRMWQvgMc6X8kFHN1zW6no6k1nZRYViHsREUiLe6Ib+UA2kj
PNzJXYK4zBFJK0UKpDscOTeGuPqsoiuO9oK5YE1FVIj18K/Nm4FxgJ1XFuSw6fk7o4rzbF38Zu1y
6dwIbNGGizjeCRpJTBTmHa6PDzDusMlbwLt76HcdN1LShemh6HV6Zr83FjrjnRX7mZAeORWad0Cg
93CT7oYN1bhRxOMK/NUk3zzVnxeBORdqvIqrCuksNPKc5MgNXaN7VskemnH482VD1MgtOiUeEosE
FTAje9nRrAndEybtsXo7m9Ttgwcdv7LgCf9r+zuGcC77DrLRwYveoPWX7C4hpeNu6h157YqauZjm
cWUzjmLlSyUv225yRitjPPet6N84021Vy3s7h/wCun98+NwaSzMTXpGpb/HG33NOlwHkfJDOprvn
Myx58xnlF1KTjf+AMTYqTE1jKvod39Ht9F0yeqac+DU97zZv7B4YpCGJ+nuBUM4/EAHQjPD4IDj2
mbqu/HrrZQflZXJum8qIVFGldyzF5lCQ/lOKVzGdZUBHB3f/YeUEFLSdo7pBwXGX6GulrE6OILkV
+bpPrPUn6fZUk3cspQ0bhjNn25jBVk3aj1JCwcQ3nY8AvpFwUv1dN77NwPZafZiunf7nSmRzsVA9
Y/qdG8HRa3WswbHZcB6+i+Rb3i4cVpGLIT+wjzMbyx4poTl0DzOoVuYJil9wllr3569a1mEqsrTf
8Jo7Sd0cW7W//IGGcnvICMJfCMnSyIPJa+mrIxzJO4QpD8dlyVA16Bw7PaTL4FzgSDslYF1wJd1w
B7KWIkGSNavf8EtpFciwP4g4uhLUk+w+7OfBoBk0pdItj3ec9ptn3L+Y3CQF3x80f3jBjZ+kyT/g
IYbOA5mY5q4zvUJO+NZos13p0TMwdg1qroF06L0SI5OKdomWIKa4ieSpuPWEovSBrlrKgYW8aiUs
8t+ApsD88ok3dZWd1wIRKWRpN+dvNPFvB7zicxsJEewMYN3TYr8GmphGEGVuLOwbMEk8Af71PjxR
WHvXk+7aEqQ592Hf34ISSFR1iTTRGE2OvrJXzNxUhfMtxn/CHwihccd/Q5m/by97ukEqWZ8QEsO6
gFqa1Jf0BGy3bDD3qrAokWzIMYfZ7F8WLnG8Cjq6GBJucjcDP0TRLNlxtpMKYod7WMeVmTs9RFkP
PaJoAXwlBL8rQMuyWlDDyw8V/KmxpK7Wgr2OUODDf1Dmh66x9B1grj0D9oQRHKEduqxSqKyvaU35
goijqyHdPltTH/7Hrr5KuzP0uGDkT5yM3HMWtRv5fPHSLj8n/2J2XOl0Zo+wx+H+VH9bgVXYSmV6
qVk38mpzekIJpFn/LH5SJhmnVIsTJXrtwD4Xto6b3e/xUa4gOhY4CWle4VVZglDPBz6/3iU+1/Nq
lwaWejbO3BMz/nNsc0arPBXq8VSx87hnWqZyd3Nqnj5VA6jimhBQzr4Yi9+z1fX6lRAmlfK4zAPY
MT3BsWyZfGP7OE+/C/1PZvT5HzbQ5qOg9LrSo+voD+DNEnLZFBJZ8CjiJrZhWnSj5a1wpUGhY+Ei
bIpiff4bPqN6W7gs/ku/2zPvUoxMSBhYf24sX0hKpkq/UnDSo8WdyDY2typdV7lqYqqsam4zM97e
yCtmfGG39nns/WjqjvUDqxJk5b390zNv2XWgJrndISrjbX6Xhk1tmeWpEW7mo5trYSLMPZCasu57
DRGd3GXkx+WgbaOmLzkdQ7cSD98GxAFGMj2cRH2JaeWpMqNGnoOwdB33CK66Ysbz1Bv0NtpE/Ive
PNFdD4MxhecMXnNkY9jiovw/yK8E8El4nAbyt+VRZ1h9pP5zaxbcO3KyQHD0KWKE7NAOyPKa6U24
CaUGCrOQ98Kuj6b+zAIexvTg8u6BooE7GzVPL1jMlSNa2pdpHjsiJ/1b6zs0gSHgQ4wbHXUH4nHx
DiKAl0Hp98WR10FXE23wIxqIG5HuRbHzZqxb0/pzn/PSul+rzjIF3KCPIrOwOuZVMw/T/sU99X5W
Sod34YfPIGBg0zX3FG7xmjkprDLFwPweQcnqKVFHlgoqJ+kjfr+6MaDsE8Fu69/vvuUToS0tQq8L
vkEAuo3cJz2o6GRkUJ3IvP/azU3Ta8m/S4pnq7rvF6vakDf//0a8ANUZEHtLV40Oxmql/5eutsAR
qHI6o/aMIkqfWx6FVpGRXmGusHVTYbc+0GQAb2E+VTIQH5ROTOTH64xihTTLBbHq6TVdiVSQ3Foe
VIy6uPa0u41UxpXuQV/qy3gvn0eHGYbVon7PLtZ+BI6LCQwCW8DPm8igudazdpFjdZ+i+GiEzFa6
LMFgyvgbDtpId/eScUpPwjS2xhNbupaBumasyDRxO9sv4pObgtX8zwWfBdMFfb8Y32UOEPbNZ9HE
yJWb0Z0929hzXZHEU/sAXUv6LCHxqnu5HIKB/kBB/Dpi1tu9FASV0tu4mraHWPi9YgDw4Re0IMRh
heJ4U2DhCLHO3DUpWHokf2maGjmAT53bcLHgyJHV8S8+M40LpKHumN+cvS7U7RIuSs46hE1Po2QE
HVqdS7QafbRJkCJr4LGJTvrytCBbxxo8n0lHs9cpbmi6zYzJO9VMKq0W4ni1L4rCcjakrefx6wRB
cBLO47Pu3FVYyckuKHnW7CIMIbmn7dLRRPsTeIAY+7e1L39Xb3x8STy7gXTmsgFSjHZKGn4RM8LF
h+DaW8l0Ix7vFGIOvmjpINWzOnsXxrBlMZO/KN4CH3fTVBmjIvrwToj8eqRW7s5KjKTT11L+HROD
zdbQgkCzD+nTvCh5bYFCrdBWGud9sleljfVEKRD+bX/Qv9L+fvPzCPQlnlcXbXMYYruavvc6w6qC
Y8VtQ7/Gqox9PtMBzsnK2oAsnHZnj4s48VMkaTs1kv8hpszg2G+IQZL2MjSRszfjH2e74f6xjLow
8isT10Fx+SIsiVTArSGC1fwGNbPY+EqTHnfQ9DIrq0IoN2kClWpLbe3GxTpa+EqeWlgkrrafz7Ur
Ml/cjX0USLBCNs5VwQGmhFOyWh9LogTcpIurcrRIFCYXtYdFSwkfabnYlsBalxaondlbQRVO05WS
56lpnosAmaN2a1KPcrplnzlkricvsA/udFJDAL1IvwGZf/7NWlCaHhCfssGdZQ0Hzx0tzNG89cIC
YMo7UFhECVOMB+Rp7atSySNZuWqOH/241gDGAguIKKrdPjQIBcZ7/EyStFuKnW/h2U7lFcrB3bAQ
CGgY6Ya3DYZ4qWJLHFrsPILBCdya9wUj4BbtlXpabJC2JSYjI6Uf3UDFuaqurG9YLiXJfJ49YGcS
xtsASFV33UHtCIRaB5hoX0cFDZ9g31BZUr74O1vSrBMTR1s795/xR8yCGg5LeHram4gw2vceV/yM
/wCJtjiLf39fXo38eOghHjpUvRHm+8G9HwhTJqNHGdu2nCJyujvAmrDAqaRToS1eto67o04jcJix
2kf6qjNoYBlQer358SoloOUtIdSOyWrHhQA/se77PPwU6h1g4Jny30bQ4LlEU/eNBrNMlV2xGLx7
4O80yWtdr7ghCUqjSNR201+O0CA0IxZNy79LOpiTl2d3SvFF/pwEAoRuj6TYxk/dHa3rNavMcdBC
2GK07RxJiup4zycnddsgMB6la85cKtU3JgTP56QZRTCebxlf7S0COffv67OG5p5mn/0gAjEQtL8R
G9u1GgAR1NjqDw+grR3h/GyMoTAziVoKczO1hzwDRW9p9bQXs+1TnUD4Tf+dzQJO5vYDdOZWIm51
lsQ0rTOK4eQ1SRijv2l43SHBr9lOFNNgYNk5hOAPPpoCq2EVmjtlp17XsDa3rmTjwh/5MPNHbIRT
U/KCjecjOdqa00H04VoQzo1RTWSKkHJNIYGKRW3akhNK2Ki8VOe25kMw0naqn2fsSzO+FGahuL2M
0YEZtRd5R+tLuvkJBT09rvEM0uYkSSWPpbs01YIB2iuHiy9fEf7wmT9OiHyxiGwd8cerxlpQMUDw
MkPyrslGt7F4MOWc9RTZXIPqjHdI3GETYX57qj1sDg7rPZQ9//2KMJnfOuydODLOKRGEh9apbCzT
IPQaB7JGS7HpZzea7jzVlngc1sh34eauVniVvI9L796fL6HO6XAachOv3uQl0hLnw/ue7Kkw1Zst
OG18IF1CJ5B105Rs4++UuagnL99aU69gXhH/sTx5XMxHol/Qbv7B0j47G0i/v7Obci7RYO4HqJxD
wB8ayUbWVOiKKuyu9ipWQHTCkaaGaF3Pgw75Ze4apZei/e8W2j0s1c1RoKLjltNc6Y8GVlLzcYbv
Jj2ipl7z8IlEeJezed53ks5mLRGy9M0O9iqWxYYl2VGblbIzfGrgy1Y6RCnLst2iuw2mw2LIqWIY
nPCCktrU1rTMPWptfdoKfu96tZxI2XdEivsc0uaZAZ/O05mgpRy7gSQi0FQt81Bl6BKBs/SaSMxl
bFFQR7qe6MVbNlWnRYCiCT+HFZ1KE64xAldo6C5Ptks4n70ChrUYA5mpqpPBTjRQfMwbYXOOdSAT
BtAlEOEuGkZOaisQ8r6jL/ZgCuEMt74hw1hzVWXHY9JnJu9H/ozHC0e8GCFx4zCVAlUN1Xt/lFxz
/nC+xZZn+OS/6mJTcPbOSIOs/jUVFd/z10K/AZRNrhgwsiaNkFvXxxhSwGA9wr5Im+ScMQbiq3AK
Wxd5lLb+ss+fHN5UJQm20GnY3RdHm7lPaAhRXCwmDrEq7up1j4z9lw/8XiLkj1NvCNOK7xtY02Gc
meO3wypoxee80zQKMu5nJ2EAfg74BRXn6/SaqzvtSVX8pkKhKXrn6AO5rAPOjIVBdnclQHD0ICoJ
3CJcsXqH3Lz2WeBRIBE1Vq6B5ZIhh59CnvI6gnVRWRuQrX4aQWCf0HL6aBRzz6kH+DRdhBq0HGbC
zPAp8RsI70StG2VcmzpT9f6gbL/1f2NK/QSzgEBezd7cO5+CCH2b96EKuOXk1+AaXjpeSF712Phm
ytyWQFdNYV+jw828xsdyE5aRcj3Zq4XLBp+Pg8thc+Wv6VQ0N5F0a6eHWEjxIpvsYVZcpoFCSmk9
legqmIKSGPu0mBx6aYu9jydu5A5PgfStqDssK8e4v5/nniikFCnRa/VSfqtl+Gb2Nk2WzwQaz7xh
qjwCZYlwPvrkTAxg57LfvCnuTR2KBC0qyszvyNfJzRrpIsiXIM3tRjxtYruk82JSf4TFqnR5qTst
p5Rd6wwZE5DYGLuEoEhnjAt2hfz7vqvLWLKbafwskiXsOOvuY56pEjnL+UiBacvIKDFx+hsIf/BO
v9tnh0e5SID37ozlTtdtgCewnqPmkMXm0SbrpWNC4Zx+9ntp1nz5Htzp49H9xtNhIdb5aUFZ4CPd
1yoGYmUNwRH+N8gMb+PAF11QDAZXbQ6ZTPM/5Rp2+XoNNnNmjc3fJeKWTPSsNk113j5sXT+uCj+r
8tT9zK4ie4NySOBiUCejhT4pzM2E474Pb6JWl1G/mEnB6VCU30tRTPMMAJTv25gK0t3P88zpqrmA
UiAzLSIFdHr9mvWtMP4VgOPHQZsvkLvDOx2fggiaOD4dkNeJnhneULZbTCBeROqZBXoa14RNU4XQ
dd8AQqXT3eOCDQX8WlGYqKnD34k1z/dht6Fgk2GbG9rkZhGtTI5V9ThZIIY4FTAr9q/sdDOViHNt
2exYdgN2YV1fKBE8ukcYz1AfriQGHlBFswo780mLYsS15w14ZXyfRk4Do9Kj95sl1HPShXalQBwx
xfAJDLX9Bb9wpMyOfjiWaRe3pzl1O3CEV6f2EE83uF4s8R/kX5j+4pPZoHsNzDP9oIzkPMFT5oVh
RSXTngX9Yrk6RLK2Q5gN3tFOfD6C4Oxbd2BJAXL8OOtSzPqYIkDE1fQYbA+hkgCwZ/kt9pyyRVRn
aUqSeBrHK5xe2aDJUOw+PgHo0HujPqHq34zrXQLasGdU2JH0FcXV6r84W+k9T87chqCtz2WbD9qE
peAC8dOXYsKDfNSEwHrAElq/oUsx57W0HZ2zr1hT8EHaeYPUiNdJcl8xvoXw1FlrgPHUnjZVmcxd
kOuebnc0PDfrjFq6kCTRBNUfwGnYtr94P7bFr3xvIS1pvnroIlUMAJgHsSzJBsBM7A8Bf7yx1ZmX
eISNMaFcgif5uEOj+N265CmE3/w2kLAFe5HnufWEgLDZv1LP0m57UB2UG8iXvIJVRE73kivpHuRo
J+VHSQhplC3FkaizLpJZiOPwBBTOy3zFG9D59aUY5dldYR6nMjd32EU978gGNOZ5vJy3lKa+rtwf
Fs3LUnaB+3Di7+NWet/3K8vQO6mFrxbKjeSpc3RTelRjse5idfrR1c+y1QELTJoGdfmti5oMEgib
bLz+YjqtGMhTqFoRjnPeSxEkSodK00hvAnY72R96HpZ4xMyI1ZtU36ZUnXqNKvJx/IdO/z9vcchU
9LguolbDF9TbyuspX4DLWJ+DUBCn0ZMhHnc9zMJM2rvKP7lN580KwSVACEObegFg9LPQeqYAljpR
Qoj/s1fHhSbyR6X3OKQqGpTVpmbQwaMWgM1TbOQRmCoph0XwN+3xpGi5Pe5ukkMZTY0G4i4q73Ws
Ev+9llRvo8J2C5Q/0K1AcCN+elTD6ENZ2O/EkWH1VK7VTuJ4U+H33H0qRJ2hhztq+m1Cr7DIWt3f
qJHKLxPijQGx/u3eRD6MSOHh1P8KcjDQPbRFJwMGHtvQyeUXgqlv0GIqQxMLwk82gRaWJ2VUqESp
d5G5xKEiLY72q9DprZwz46Y26Y8QiwKjsA1WZFJMo8TUmHCYB+n71ArlKF8Xbc04sfgXOuM6qtI1
Ct0DSSH2u5CqQZhsQlW9Gv4h5bhUUZSw04WS6lLUooNMh/BNOZX+DfUksZvi7CXSQ925OWtgQAJR
rKx2braNtT7HhG/YIHuJbB3Jf+wyv4YrebFZOw6KGOKH07X/or4Aw5USObusjf+TbD/wif9nQINT
L3564I3X6Q4Aag6mAJ7MQwkDjfhn36oR2mQ/VdVTjbJDAXMrfz1WU4/64V1uGWyVAp2XhIoLkNZ9
nT/mQhy2Id33M3XqVOhzOi1VtslzNuLNGGGliuDYNez5ztqhzcl5NywPP4RTEgxJ6oxe8xzixLjS
vj7JhNX+H2f2zsxXMqvVKaWQ9zLymNAlW1RZaJWmiRVHWx3/QV9c5uvl8y9Hx8hdP1JcQewskPlM
iyzQ4eP45l1ZaCOcBxkjjddVcMRiASLICBSSMcV6Tv6TvHQnrcZ8ft4uF0/QdDibh2hjda3Bd0W+
1ICbJIXsRtKpvsVIs8+DC11AkTFFGYveSFXnHLOSh0GysfXv/JT3L1UR82kWGGoeThz226sgkR7J
xrNC+uB7OYdNvpKa0W11ioqQ655MCHWmEpNqVse2es4dlYIME5iXRgDx79SHhk1p2LoyymmA2aOP
6MHiyD0IC30e5lj5SPGPpyF3cF8FSZgBn0hn3LW1ddGMMUMvfRiSzFXVIMWeH7EVLT/2PSgNl/lo
JrAP0y7O6N3dQHjcFTo/DKpiQlmUnv+tht4bMYIXtCCwsSNyWh8kiNJYXRn2R8Ic8O8UxGmoI7kn
k6wUNiIUMvZlNd8HNne5510z4Xqm9ouywYxlODwbJqizEKkVr+xcd49aqDKgmikSQ+nWOYx/nFNU
w3PPNiAnCd6IfG7jCUEfMwAnHTEgZSODZ6myjTX1qKgWQrIQM7lVQJR3BfJpzFr0XvX4SfXzCyhK
g4IqOWlZCstsFSGtZfk2QOySYlW47jiTeQxPialk1KkjiRUXBrQ0EIeCG7a8x3zpbPXUor4OUpxc
wRPPA0SpnydXJDUVUcbySHrULqd4AcqCmHJENqxtcDLVL777sT/oDv3r/gg6VlYdvh3GkCTMf0Dy
HcC/wayZ4fbR3FwfyeRi9A5xdDNwy39d5gSZb0Ahj/soZNasvecMjXCoGVXHI1JOCaHOOOuo7hGE
rXv3QnfLPN+u6PpLwmAW67QWw+dBl2iX333i2lyrHtsbBobXVN8/Uot4ZSlGj6NChFEMQ8GmPpwF
EhkCMSXeuGeJP95IZSXGC9tzGofhh0mBFXS/z6csaLO45B9HOEDdoVE1WOdgDeQzD7HXmpblwmsj
UyfRinmIWcXrUAbK41ym0UJDxk+CDJjUgrkOIpfvTert8taRdxbsBBy+RifHMTak3mNlipo64fTJ
BYVMG6E7+4QH0+Vecv5VWu30UH+3TExQv2ZnC5UeZg2j8IM/d6rQvaufm8DklFch9K6jtOOXjJzL
+ZYo2EWiI+OkDvNdFG3MR795dsZZRdE7zUZKD7SR0g9x06XERLXUqm3wSr9hto7lQk0Eol0+1VDl
QeRWoeyV59i4H+SYylk2BF07lp2odYWp+Ai0P6wtmYAn/7ErmbmKebc3ntj44yGY6ZtjnfeSd53D
2pWfz38oQM23X4GM4Eo8FJCE4amGP1DGju7txmhLFW9C7vcsBhInhs4xjLF5fHFCNhWUqoxJrDlv
szTVSszldIbhlvkN0HYdYak32N4/WZnDcYVF1N0pXpeqe3KuDuvjxb/RVEfXFnhWWOzoGBizA8jH
mcwxuyZR6oIfsjdLizKnXVK/faihxQt5FFtJgfhGsief/F9HLU7+HBuNq8UHRiChfV3RaVoxojXr
GdIKfz3FCwMMpNXTN88QpvgJZ8VQcN99EyFHSKUxm2GIw8rGPkn+xN7UZoEzgqJ/F0pGR0FDg30X
3SDPlA3LYYHnx/FQSHccHBBLWswDjHSDVXe/v1n3iBdyzFs7OZpTRJ4iZ4lsPUr+ovAgEGQ3tVyd
kQn/3cYb9VEoKdCG9liNoPYztc598byuecxDuihBQ8kdtU4YXQciFD/7kyrWbDeD1h7KvOH/NvTI
D568cTLmKbsRJk2BwIsQGDNNxEG7PCvzdA0fOW2e7Jf+oEia8TyLzVs31I5Sm3bek1D627OiY7VZ
8n8CFuX+naYWcPyJiJQOVUMIiKZ5zpzeW4PfvJ2cAhtAsmMPuOZstfQcdRJNLD9eVyU/S49w6J34
BRvIMkjld0mbFFJHQUEGler676/5RNZeyUUr+BpNEZhwfnda8hR7BFaI3CFfA+lO8d3qzmyWyUDG
MQcp2Imm3MZkWyb46qg3qsRR0iFeQ/MR4Rnj40i3JyGY7an+RxlBP6za6qyXgybYXWE1MmzMg++z
c4qTTUUqphl2IdcCuRM6ZuWGfLvCwU6UOJmPxPh6xkRbXS8qZ9a16dDGt/12PiwwX1iMACqJ81bx
mbqvzn1ClPw5qYSc+czRzWULh4dKnkPeg/2OEs14ZAmtO3AC9GqUGziDAQLN1X919W0MygInwh28
tRLZ7YXyem3p3UrAnWHsm5Y33uIy8nbvXQU3WNBhFXcDc/kK+kvzcdZ/wxMUHXsugwi8eiF4Pa/l
nvh6xeTCq49qV+hcOisTYdbcrRbZuFwgDJpyv53O35UrFqwhQ4H+c1V7pY8dmt/P8b9xFhzoX7u7
2ZfDMqAd4PsKc3tVkVdh1QZ8oe3Jh5cSm/aWGc8u10vq+xS457QTNeG6nlq+VRX20x9piXIzB+jT
Ho4ZTExzI9UZN1tmHIwbGuQcf7VKHTGImxUP8uNPGlONZa8ev7sajh2zAomjC+uRhpkiiX1olV2m
UJGT1l5UrQ1SiQLXJbfiQl7NejXhkDBxfLi4wi+d82RVHuJgZb3KkYwyAuyyN2Kma/27pTMjSvVm
Q1zQS/o05Evb8ZDAMWs98GvJ2t3XE3tKpF9eEKU62R3ww+cDlNn/f25katDJDTZWLhej2ajim7Tr
PebF+D+b8b2p/9/w+od8RQee8gLFtadUagSyzWYohFFjJugLZ0KIRjwuXjCfh7uniKu6MSBVU9rF
muLk3KAnwcUoI7usAhLb9AKybrCsWMnXc0mCMqycg5ZYCPAiXAXlSbkMT7ARTW7mn8HQcwKK4fQb
IdMlOHvdwJZEp21CCZTWjo7vE5mPjoDjSicVM01jKiDWCq8D8gQu9yx+ZDgHRDnPGnKCG0fEPwin
6lRTow9MuPFZIhbnkIS5IqMC+xrEFZpuHRkBqjJapMjlWkHY63RBF3uTR74kcqXScquh2CRyCRu3
WNHqzZB29E9NKi5HVBFR7xI6+boKx2Wva5JiiV3h9NFbbBjkDVIy0VDELawyxDnEHxMD5S2hctgY
IwkRLkOw/MLjPU5VW53eE0M3pJL3kE94lfiOayGPHAg17tPtoSsIuKcL0X8RKS2q16TVhhvJm+m+
rto69BwUuCXXA0qxfS7bDhoeI7n6b4XILafhBHDKjly6qHod2ctRJu6P5ToUAkY8ueFVepb8VmHq
c07wD1ZmNGQS4TmGqGs82NI6uITy04WBW0sNDz1du6kaft3kLz6sTVzLitez5kFcjin7xrspEmxG
YApPjuPzQa9nlWMryAutvSCensCmJYqG1z8tpzQqIl6NZRIMoonrOeU3QAgoO6FK1mQ39/pHYFQP
twcpMuDLCoYEUAXLfCHMtz2BxMj70GjR1KnBSaNzG98/MSXmdk5+xc7jhPKCwbnRCofRXlWe6acq
lLSvZKwHMT/n7CZ/+iG+GE78/vSQe/zqR2TXlW/TrPceT0F3WhU4yMxIpspqSOXkPYimiEsGoI/Z
GimotjV/BekT1XxtQpKtifSX6FocdifM5WQJt0onTKXNzcdO54ub5Y1l0wEDx7X73/e+mT7Pb0R0
1Ihl3r01DZF+NWUE0fC8OgQTSNiH4BfqIpt/CCSBCpaFG7d66C6iE2l5jvEIvlbOx3e1ZKmIKwUY
oIYtKmIzggBMJt1QkK5L1ifNZDFztno/pZ/msCSyjhAomPKF+8VqsXkDlIux93IYc0z6B+CMtSBh
Vj5aaK+PNWOe16kTt7KdOIE5uXup3ekdf5kUIORWMZUTwqF2F8hbedQt5lFKxGb36FDQA0R8/B1s
6Qj+F0nYyZ+2FznwzMaMWrwCkAsqAia9sEQlVegJAnsJn81LWpLrAE0uU/n6WcPYl17b9+3a6c2E
pr4pCO0bzte/gNSN87DJM1KFp7sFMzkTrDUMr2m2c/EvB41B9m3Oj4da+Cp8tmM42hUaZOTq2gz7
qyWwXYIUvymkYDeuH4OfT+8plCdjC9udNP/PmJ+Sq1XlDXIXCKtiO5ed85Hwaxvq9SSXuX7pzo1i
vvnK4/CX+3SCk8w2+GaBNgQj8R4qbaNbEdW0P1UJOGROfFf7IuyQYCSjMg/+3m9TXaxxfWuk1gWd
uOH2NP2HJ9FrIH473Db1hhtw1nGVLuNJeBFZivCxLkS/1+PPrD5XTfp0VreN9k4+EbIYkcAAydYc
R8COGbxjPZ/5iYOfa+Y1pqiFlnCaEbntp1asxwlvfrA6vyQLQNCLykXfnnBeeOzVb9CJSFwgxUej
FZQebdl5BLB9qIf8Ahl2MNjwf/3sgbAosaoMh8x/9sNAxuWcInkTTDsnK0bk3dpevIOPpMgQ0lNG
a8pzqogHvqDhGTUaJOOsipwE2fdNMLMVqbdiak1R5unEfOtVeTqltTv0JBQMwkKId7lp5gfHLLOP
m1VrVPJLaABvon+aDSymoMJdSTxHHiKsqTk4BMpaxlOX/ErSu2JBJHLuhbihI2HQQ49IP1usCgdI
Vr+1lTnOxEGtcZM7MDtLyTWN94ESDzaro9FPEB6HiYz0kkEizd2E5KgA+Ly8r+WMfxCXV1u9yTCW
DKx6D+7V+Tw08Xn9ZBtVlojCpn2ua31B7G7dJVDH5iZUKk3pTweAU9R9g4IxPcA0j/JCX29A8Rq9
vgDeRYHnTxQluJNRBdD6igUcGrZK/Fd03RD+pkZ4u1BT+OSWvnuA5MYLq6s54q4lqP06zOQJjq1t
shUj4wMrYPEZPr34nEHE6drmJ3bEsM6OWJBF+xU7GFLkr+A3CT9ybMmuiSEx5sWe1PAIzllQRuWV
jGzosvYcEMq2dDS6Am7Lat0NbuKGMT4c7nAqpjLd6Av2jZ74wTgwV8wrlt5lH3AiVfxhdLetIPqp
tEwmcuj4K2CsRxNDUUP12tJXllVzoVuhxNgL1oS24tCl0T5Ovqrc1nLau9C7aNd9pm6leethrk0V
RMiDZjHfGU1wuhl5VcKqbacS9yVbIpDkBBc200W19+Fmd5bWglKy/S4uYG68GInbgQyAPrsZ9pYR
SsQEmqEM3YvWXboeadQnnuKwruP6QM2xrnHXY+07Pla4VRq4T0QsXsjMfJaaFVEBkmlzmMcRaQBk
BH0AG3v1hn5sIWIEiCFHr2BJM00mj6J7Blg0WY/75r7wtQ+qwRGIwoNGwnAbLMkqPxrhe9jwFR3+
dVYmgSz93TgDeVvnpnh1qrplYvWJWMsm+wEs+utPBObwsKMcX9vNrLAfVtJEY0nmw5kCIMR219hm
IeOWorevL5iHctMZG7LFpJtpdOzqtlO2QD8AMvAhks8ZolWcODhi2qAbQqEQi0RcOX145CovqOrP
uDO6yxKescKg/BDyKQo+87xk2bOgjWp2BM6ZpB6dW/7OEVoLMwtRJLxf2VHYP4CxWDP8d2CUQM+w
mDrhtpKtQ3PyRyiZ+ev4EaZnKZYl0TPkiD9r1HxM6QTVXMFI5mTq7fkqV50IhGty1if0LRukkf2G
gUAP7B/7YUV7upS/yPFlU8odqjeOEO9ekh4Vvjv4vmxNnyIuOgAOAE7iO8AgbfkAP7gV8jrlwJrb
U2bm5+kwmwU51K8GKLjwVowsSBHNJGNoOtboiP2jhvq6usEz8FO8REdfSbgsYG5YKBq625G+0cNB
bHxX6R6SG832bjLieFXPITW/j3ls+reu151azVL+Vx6og/HyHCxqFg+uQgNmPHuu1rTHC1N79xfF
mUbQgWLHrjHkZCa/i7sVe3FDw9NHRymzpyl/r3BLfVrw8nWaG7QPgVnKDuLYm5k0so8bwCAEwAmF
42cjrbR580cIpYf9gPxJMElHYhoxp3kxKal/wdZ24escbSDJv1F+czy01oGUsfuzNeZJUFJl38BV
ei6wNXhiBlo2+U7VMlC9x8zGohMJff14zZGx1wJ0qBUQ1OmLN3wh4EZkwbA1On8/E12iGV8MTO30
XIFUu/oivvbqYbK6qiaMprQ2xa7TMmkOh6spw9OI5v9PcJIneKiRVD/7qwULvqXLtfIFkshN4JN0
CUFgoKMF8HbtX8IGhJUu0i1+p8g1swHNDBMu0vdtUEKrQfbMkcdKyDuZ/o3q57ar5SDDZgPI3Uiu
gljyQcOELLozRHLQDffeseSDJKUBrfeP3AZY6bT1QgGnFYCtrXAd5BCMmQR/hmSNkeolGCMlPDHj
L9Bo8fuCbPubzK1VYgUIXBJXD2ewW4hoQqhKhyohJb79OaAH5qy1KfA2eIf48/HxptGurayGjPv+
vkA220IDe2T31CMwAADRtDAYJJHcFXG9VckRqCAkRjibkSMAd3Ki0EFRSZbu/u2q6EeHi94CUtfR
s56eI8I2/Ext7DMr31Cv8GzttOMKlFpd1zd46++jz3RB1Rqlk/TY2sG/vEBVf2VN3Fx282qfCwlD
1ayFrkukFTIe0VFy6uPqKWhI4mouUkT8zn8DdEgPSPUHxzqtIibdxXux3Xns/hrsE4Vpv7s4DAln
naje42N0pvvPrRb+pczVXSOpL9SgmeStY+cDHu13GuYvzka5rTkqqoIizQx1mdY6W6WCh+ece32g
+iLyLauqbG7gtPXvxDIAo7oq7QSYER3pI9c1BSDoMnxzGEkLwqWsTeR9WnC2EP0sFAOyHE7OExGR
V9ymVJQt50s7WTpffw1TKyIuJFF0P8A49AJi8ojfoJg4wudQACPowpKGWET2oW/SwwqS2yIMKZiZ
QWdCH0pN3BYsqp69Mh9rWqBLTcP2bhr8Db/Nf3Q932cm1m5d1sT+6RU7f3oibsslPAC6/MBAHEdQ
7n23ulnLck2FKtKD5YM/WM6hrOG973dt4MawRsjoWq6UubKGEQBVom0bIQn48iMHm74Jy3EEH4lx
wHATRi/8/zNKFtAb7N4omsKNT6OSgKqm9njv7H0jFEQm+BjImxANt1gMmdtxxLCCdylQ4n/pQN4O
4DvdgGtrz477kM0o6Mk1C6gDzwGNnL7G+Rsmgju6pt3hZZobD4RBS1ygWX6EgJCK0+zJojsQmkB5
Mnxo5clgaQy9KyBfDqqnAj/PRUzGOV8W3qbV6t08JzK+jLVa+X2zp332x+XITeO25rrcnZ9Whc1w
Tg1HR6WJtJK9qBvmKM40ZLoxvJoc101zfU0rEtW/X56Id+zhCGBfAgLZ1G4ryRkZAQLMHOgbBZCT
JDrlzj/GjGxm6eHejI3Fq8WCliMDujfN0qcavHlfxf7BliTbOJHUVuE2aIlC/PSqvl0i/Rei4ysB
7iX8JILFvVo80V+HBSH5+nmOV5Hn+tq66xXvT5cxMICS7xow7OOhqvTIK4ATG0Kj5QEDQCxg/2Vj
4Yf73K+kTgomu6Sde0CYauxmPntjLgGtkurec32uhSn4FdqaSaAfVWFAWw9NY21nYr+YZKmqjFqp
g7R/ybcNeCVPcg8wQg+YbM/vX+62duyn9jJqZ4JrFR2C82rZNIGdslnqaUzfTOTwharN02lCR9V0
u+o3TbzT5Vhy6HSnBcJlP6uPxeay6PN1O4bocrUVnkYP0sM2atxyPJ4WnCkLpom32DnRUSpxgQYF
A/cx1omdscURoQG4ZaOOq8SFko5vU7UKEf8iUnblTaq+xyMxB4ZkAbz+3meb7E4bX0adZqAL/7hw
LqyCQX1ANkRJmb6OA4320rxhavv8Qa0peNV6CjeyfNzSPoKpnrxX9J4/trEWz5ojEikEJpKod9q4
nXS07g6d4Gm3bs7OOYWT94FBOTvAt908JOKsI+m5G6P5vd4GyM3JJebDdXa+UlW74U45sD0tSO87
Z34zatYJRVO5MiG9gHH2b+CI9jKddm1CZ2gEwprYxrftQH+wakVSMlq/SnzhbyPpGJUWi8cWUEtw
9zznJTnbcGdAgpuSzT0AcfnJyoOoB3JMW5BqITS2EboMAQqgXAoVxNETppUJ50l+grZ3u7EVqHou
/mc8urO91bipWlsOBTdbcrdyEgbKBZFa9T5AXZ7HoJqNxQR3KHxrzsQoCQ/dg+CHoyOg7FfD6BU+
pZ3S7nH6gUv0PM/zav2+/mLlQ3hH9jvqYe4XiUCxrrblv1qDzFQTl5EDkB7GBIhpTj5MKca3rB5w
LmiyuMsCF8ztoynFZdAxGbFOP+D9wuo49aMjdJCh41vr4rnhBk+6RGAwi119VsFs8A/GklH6eocf
5/UAEZLouVPswz+RSI8e8QOXIWTczYxW9746DitAnZxrvNduLsLDQ25FQHADCstk/BgjMb98Pf6h
HEd/8tImNuDt3u/X2QSeaBMu7T26WXRZ+LVU4ccgifq0CbptQx6tkPrKjl9pkZzA3Gv4CKeu+98G
oycBWGhxZx+6X3UxOuKoSd4vMsRQd5fyR9KFWgms4KedyfSxulftOwKyr5gfu5E9W+jL98tG04B2
Aqjs2vqeN9rhi3UAk/EsKAl0dh3abCzRE7UJcnf5MsNppK9UXrzDMzkGZCOUCbvkPSX0y7yonJMd
rRi+caaETvIFQ1spxeuFhAs9ac5EVzUOpgQKi5hkoNtD1KBKtsGwX8mv1rvDoAhWZnixkRLzJrAL
AxvcNUd7XcD9kGOqmnSHtgDd3jXuV3ipOAfQE01KSAWGf44k64IZ+QgjmnVEJELJkAI67wSNmria
hJFldQH6IkYhrzhGQCHbjGO3s0utneKnXLT7YYOoOfZgwMNlM+XDiSVIO0x3B8/9EL3HesagHZ0w
BK/8x7ZEFWeCTHOnXIb9aO+wXS3HH9Eiz209ot5+maOCNT6+rGoE+rOwS1ksaJwnNlDHwxEHFf1h
Hr5pFrOdt+K48yXU3EM6PCDWDvB3kAqG7k3Uq5cQcNrJbRKNFE5hWwwCAG/eTzhYQ8h/VZKcCDWU
1XKKT36TF7ccVt+9wzEw4FQGzavOgWTutTwiE27b3Ulyi8lw5CQ+0PpNOTxFJYDs3+h0DIAZwprl
2AZaACcwoqX6JZIY8lm8OXi8fzYI7AU+HF3w2Kz+k6joELStBpsDa5/mopkRyrgoB9lxVTUxL4JT
pA2EO+zTIB+BCqX8Wce7TbeLFGQkWZRY4rnw9Fs8Pr5MdLrlD3uQ7MRvpbLD9marZ7Tfr79GIr2U
/c/8NeeN+ohweIstjy9Olmxx3EiM+zVEs3LFBV4vDxN6uhIcXg1LM0ZMX7jWVPhyLkfpb+9hEr1R
7K3wbqNRAvkH9fYT5OQyMPqcHccuZ8m9hQbHaU2ZRJnhK7z3onTol2q7801o0vQZ0OrRr5iFgcns
qGnMpnvCrB3Lhvcy9SACmdSJ5kKAU+9KiuZpaavkChtrenq0atT67Q1rsCu4KKYPGTRBJ9a0KpQP
Jlw9EKuW5aD89IWG6pMQnlsck+5Foda+89A4N+Jt5p1i5avZvc28IGFAunKmangSU0+ttxX91G3V
o9PZY6iKRUyhsF9pr4odZE/cr4grGFilloTregoYx0UiWPTHwSy7qtQFqvosgbSRZiDG/HCSzaKj
2Et0Uj6PwztKtRZXmfFMI1kb8kGHknFL/lzrVdOBvu79GQ4S70cvqDRSU7CHRZVrml+h2eLa9Ovs
AX7DDTi0KGiSF+U+BTMqYm6eKNHAcm4UPntbJaV/z2pRcao2T9TfGfc+scwZIl1gBrKOfbfUbMVI
QmCXlnLAnY8z8s2rs3oYi964XRjV46GSN/2iD8a6PWbBnRtGV1kqGHU+yAk+lhVQCkGZM/xwsxIK
YwHdQul/jvG7nkWnTm/zTYbFwAsbSP2qt1q3r+J9KqLtA6YejP4rlOqyRDbA4HzDDNeO1ZQLd4A8
koZppTAI3qwdUh3TSgOKynyEAFGZQLtBbL+qIcO8ncbzzBR67sT5XIIUBMB1OSJKNaSTLK0Muwat
Poi4ZUQKjJXIF59kGn7pM6Zh2nZbLj7JXpOXPeNd8isVHe4+ZV2YUATwQ5InctB0weJ13tBpV9aZ
YcdaYSj4f0qL91+wyUtoQR7Kxc3LEtTh0NVk7bFj4f8Jabd8/RT6cFmynZjXsGpBHeMFoysDjctt
RNN+VoDhTF3K4xJlNBV5FI0/B9RgG3XahBL/u6QIv5g6hZD2Ysg3Hi1NrIqnXVpS2TvNo8EBGB3H
k3CG53/VzNyD6lPbbGOOP0gd3NnxJUej5fUoTXLCYxLa9FQ3cq1m0Q6I/zqZtCSJxTRpU5Vv7111
VUjfrdvBUjkLCt8f7XCiHZk2B1NymZ1Ui0VTeiyONhSubd5b930kvkdPnzDr/CuHoTxljtRiw++w
eAArDtyLXT22xRTsCBhbKfJFi/14mkl+Bnr+BB12xNmOVTQ7hzSD1KKoBGLQB2acfQCv/uzW/SqJ
epwIByJefxKqYHNEFM3b3d3m+C4kIRhj1viibX1oquaf0iobzoUz0bZcTHqqcQ0kzPiGu6RVNwO3
zqTzs/G38/zfsPwhxoqDTuWAEuIIioK/DMbSS53/wPhG3QSaltFtguRxlqusX1uuJ9jVX2Caolcp
a5f4ABbe2ahkO+A3vOeYykeU7nj51nprKtsC0d94jjyOfZBc+vcXgSlsr0Vr5PgQ/cCw2s2MLN0E
TlyPrk6K+GSiYml/GOrUDLA6h3ijy6/zO0qjZVTxo7wn9yjTX4rlMJwGUWFJugffQwM0mgjfNnNI
CzATWBGdDj1/Q7sE3uP1wYvsLUvxPpLqEvJmJGXCJ355KaXZ4NaW60jbOYBwadLYquC4kAkFDwU+
Pa9GKyPO8X2C5aefbQE68cNLB4LoxAgsZnX4t9kn6KD1+S4TGjIkGdXjPXF8Pa/QjMnZxFxxRi1R
HQAgY+n6kO2NXiIl/5iMYoQqxlprxls4g7OYSsm7rev/PCdc2jOaxrc1Y2XxP+cHPH8GO8xWBEQK
g60LWpXUJa9mvJNb44/ZWs0TcfEOhTYzmf5ud3852N9va0f7SKNn6QrKDdLJJQfEwkkK4bbAe19W
5JOh9xAxqDxHZj1XmK1szuv7DisgHUTH5raRcINV44TGs0rLnMVctk++ZJTiqBHI0QYTTzjzzZC2
2LcAmq7mrShFFbhb1t7FTStVQf00F0majXfamepl6vznh/BtlEK+JBF0k//CdMtsH1X1ETA5XWXR
wBbiq0TyhCc7LeZ6KO52Ddhu7h+MdRimj25onQul4FtX8gWfa5Y0QX0SYb4nZfrc3b5aK5w28VDJ
qZVjAbq2llx9cCZ4JodfYYc0MTueWbff/Te+tvInrVAoX5pb1yodDGOd+9GbetjiuGEuDgQYGxhW
W75Jbz8W2ty93SwZo7o8I8vQr+6yKhjxe9BMwkZWFTru4MiXlO9Fc6qCAoGRpFbZVltm2GyY/W7C
OedzsmYJE/mUk4ejis3BLlMbo1w8agHinh09unLh6QpCetD4Dvo/KCsBQcm2z0di2sPtqafotIDm
bvnz/K9dx9PyQg04SRklN8lT9s3iJLyQGfhaXdjWslaXqSWVfQWj5olV3Cwy5cOXmlkzm5jascBl
PGOZyS/GwoLAX4E6G60fSlABz+DV+tAAa7089U0nazuB8D1zJJ+1+Qzf9L6otScudo8KQyWpFlGC
holRVgjBib5HcN+yns9hX/r3graMI3nusgDUZjqi+1OvvGMlLqqg0jHmpS0cu7+sl+JX6ASBgOtX
Jqqwqy+Vv9PbewmeCNWmrOa2orgFio09o1k8PApv/oMGCUJGRN9jbIzZJt7WHrZjrUHVtNhmAazd
sTxKHJ9L7cAbfqXvs33griaYkT8npXg7+JIbGKuStSKNfd+uUtBbpP/6L0NFCgBSUlRxdayWGWOg
+78jYQH5T1BtaDbTnEf+nbNb7xGZhdBQ035bmPd1Mi3FwVkWKwu5khz/nK/uYFFhtppcHI/2GaeQ
3AmCVrRCUmvau5ecqT49USsYWgCnsWUsGaMw/uxOSKP11H4V92tJbdWTEPCq9PeAbsRmJEydc8DS
i4FuihN8e3meuUE77nWOWwvXJhEKNuG9Aevwn3KL7vj0hVcKo3Sb7b23fDeDUs0+DZ6OH4tIYtlc
uJGn/7ye4DJTRc3r+UJ8Da/L9HeelXVsRykaJghrzV+dXD9sdAD39ZgEUohYNE1eSeC2NIhxXrJn
o8EYMwNf/8frPk8UYMzIu9mR0lrJhwz0eToQpuiTVIXx3Tq1gY3O+nBxyKVDgBMamw+ygWmrH0/G
QpBiA5ClJSF/ogFy8HGNeK9hVb0kfBWRHkScswBigJg8cLca5kIvOuVHnZL0b6koDb0t77i1Yj7v
IiWACb31YB1lZg/4AM1O1VmA6/IOKXQ61+upS0EMu8M5T+5h2Ar/1t7NUHkPBaPDiQ/+T05E//pJ
yAxrBI83lmoqILzw6RWPp92MFbnvPMpeEwXZUG4q7eE2sshGtS61vGCp3OTdV+gIFPud1mwcP4aj
3IAktAXBgGxrd3vTu/Re+sEGs/RZkJs8x7iWmElyKWwpncv3bMi5Teg0rUYVb9r6E/A1g/JcZx4s
ujHjBIT2Bz/CNU83IfvUNzBtltNFjXC2XBuhUxTOyhuyP++dkZdY9Z95QhU5HWRA5jx4/LHRykdB
iYrAPck3jJTjs4+duOAe+vHONNKlD3WFHOMzDpODZ3lAvIcTiuKtUW0sWoPsnv+q8Ae/3wc6NRh2
6K8D0EkbyqYhodVonK6FIqNwA4GW7No0BUIMFa8c087f1fRlnNSByffsJqSuHVw5WSR6cyxCJvAG
lTDUmEY8uiWM74JdQwz1M3vbmzTCglzkXQ0SFKBw8IsnBlMT6Zm/2MkZ9rMC7dn8Ikj3PkB0i7HF
9w0qxitMnP9/0M70INz+AqDX5+6yOE66xzpf6jNZst4n44dS4fLsBQHk1OmVsJeZnULXkWLkGPyz
Qo/o65zKIwfPDPI33w8wOfdZ51nihXb2PCkhVBtY5sW8qaPIEZQ5haNzaJrYgimUAY6jCT6ClP0D
bVkv7BFxX+ZjeylWKT8ZM2T8ysOV0pjQwAexECDv817LzYx+oq5Errb91/MEoOB/TO8bkY7XVtO4
KQbmkjexExJn16nU+EWaYJSD614QqSc9PhLAMr3aemKw+8ucQs3aIP3DWOajdiFQWMNstIAkQlde
ewDJIQkk9WXFNGkHM0OIf8pz/cCwUz7Ra7jGRRaEtp9u7qBxabkLaX36sX8GQFn0ZqgWyCL/F/qE
0sDsxMebrTSUh0Ja/7/qZjEfqwDRllaHHtIIF2ZJw9Ek1ui7dal7e65pH6vjfd0e8Y2Iuc/HbkTb
O7MC+usxByGzlpoa+IOpmI22aQBw5+lx/5JsPHhniBk50Lb70OoqH7T99pZQPpjRU5ngK6ifo2oj
ErJ4xUfEpojPg7wOfDSS0qZoz4OeisGTGdqm+34hkp/aOrtPBP5wy4NAYFYQ90yK8uWn0x3odOzT
w3fwrT5/MUFcSAjIeq1oVIePpK6YdI589dhDFTbCp9Vc7S6vKYB9KwjjZeuF2wtltAKIm4HhSa/t
s2LQkYUO1piNY20GrNxORht8m1C1oSRDOunaQv1HOwzx7lUgr+xqmy7jDG0qYk4nV50Hn/uWPj2K
QMYQ4wRWJR3fe71OK2KVo2SBzF7CBtIKGpPSlC6u9TCet5dXwM5bRAHuJUYUCXLLXNR7FtmnHbM/
D3j2/2Ac+pkeHo+tEkQ8Apha/eMXRy2m8LpLketiNWTb8GL+twSrfP6hbDvtuRsrDDrnMWByOFYq
doW0QGfCdkkpD8IxP41wTmKmqKIIIuTRlWTEpsI6g91stYzPIGumImNWLgO+EhDmvt62ik3JQpN7
dXvrCMU2nW3L2V6JYMvw/CWXEsMBEc/xum9pd7M7a+FgtBohhLA2RgElSnADKXWwcbf3YUA6Np76
qYdS5nDa6b/TNZUlitN+DZqOnPbYvPTOVzWEgbhlBnziVRu0zCWP0lJm1CxFz5B3rPWdwJvavhxc
wEVi4FF4LzuMIVsSKElJqS+KnPQAuFJx+KrqmZBcSvToSVEkna14RCuJu5HNn/hhyYlgZxAuxFEi
6vVBccef1lbgjnVqPldJN1adrdMqov/rWbJfXtNtYKmeCDafky9ZQHUXlHscClPLD2DBT5z62U44
royftsQWvq6HimRH62+D55lUo4G7kH7IDv7RlEKbQpCafNn8i6MWExS/t/juXti5HDxV4g5TGe5R
YW5B3t9I22BU4044Vhaft1Zmohby0oPZuG+plBtb338aUZqAxjpuJ+/Awf5ZYaZE/8VSNT+2H5V3
HUqL+Pi9FJalJBunkb/9IUBAaRJRpvdIwrtBQlJvcIZknA339JHuA89VnUedzYzQwajBaH2n/45M
7JjAodV3PZhpYbj6tzHiC+pQrDfJg0sj1vedaOpXrjGRAkibz/LGCEmKjbgNpZc+rQATOPuZwrsx
P5CdN4t39QzmGnEnjUkPd7tq24xlC7/p07UdW8pPqm/CQ86MCZhNKdwEz3CqDPTJZhZI1Ct5/Nc8
ExVN8L7CBiVFgLSDHRw//qJhVkxhoj+52agCbjYOZwhAMjHjdl211KoJ52Ha9PKSw1EmTRVuXCBk
oP4F13mT/sm1fGJxOGJLZbZFTlBL3O7PPjCRrqSbPwO7Bcznk8hdPxMS5/yjoVkuZOxRsWbs0Lse
FxDZm5Ezvoepbp7JiUlobyoY/tACyrteEWuCCHFKQE3FMEwRNF672m6HsljQmM1J+BpSk6nSvIwX
b1LsEnPBj2teY/x1dj01ZLDDVmA5pLU2hiZ1TVZ/ykCKS1KU3FajUIeqlkofwo5E9IXfaZRZh8qF
mqCF90YfaVsxrGJxTVJfbGN8dHQOF/haulJc98AK0edPmjVgWue4BAHk4JDZkbWZ2IQFWSA/aThi
0lO6J+XmcUxV4K3Mc3bIzFrfPpRcv2L4vOQRe8TpZ42vOLFqE/8LxWvMsPx83hqnAl0tnbRsdgne
vvKcv+3gni2RZH4OankP3SS7FqLFOy3Q+H0JCvaCoFEsi1A6FnPf5kX7c9LbFS/1hcPaZkOdFGCo
JOItYrJstEEd2O+oI31A7A8YjLisu6T8Z3wk72XpkieQALVswIhzI427LBu9dT9FWA0q4OlJXEkO
CHn7pDLYU7oXmJ+M1FQk1YDGotZ9aXInIW9Qq386IPVWWkHUd8UGb8nhfSIJig4mG+Ggc5AY7F+w
RG0Tymnt4XCKsVzHOReeR2z8lEPi9TQt3rVios0ezmhRGbHKIRDvNYkVOYpsRBl2i4RCUzZTCfFw
1YtwFFkbqKBi1mhKwxbMuISN8SgSNT8swfg9I8ESu70CqsBdeC1iboVM90sibpxfNYBaMklpYyBc
S5o8BJQKkgaZGTLJ5WXkVhHg5mYuBveQMuHEQFZnQ10g6xtf4TnBEDOlJR2gU+RDH6hgEeD4KKmQ
U0XWMG9BjCerTI8SrsNFgoZ3D3TMggve/5dSevwsC0+9QIjMhi2f/XF2qwSf8sdSa7yU2Y+h/U6h
N9AWO2aKRUbF5H9Dta6zk/9s1++N2mA85xRcCcDYkGK4GVbm36FgBslRzlmXnbok3cK8Z6EExSZ9
5vpzia2PUDpqm6RvEzy4nFWCP643t6guG7VUq6c73qnz2OtPnLK5CrxJ+Q6pF1ssBZ3hdrBFZ0w6
i/4T7KTWELkT21TRf7nUSd5rrRzauiN2GUKCzedjh07bdIFZ3bx7dJe/yMWnVPmZGRlq3+iMrkBD
MN+VO6C3LIjiUTDiU0IRpeM/19k9RTwtzgkEMxWfMryTGOA7ezDGQ87BxtRW0VoTyXNgJXoLbuXH
/n6Ebt2aZojkedUM09Km/fKwogjnE2spjHIP4ZclFJrsSiNcH4OAeJpdkCnJX/BjI1z6oYqxt5L+
BZk2GT3ieoHOdSrN1O2R9O6vtRIApu9zqFxmNqEJcVZajT8jIOPguC8zfU/fOuoFXBbQ6VbOet1X
13PiI/31fHI2sbKRzWeNMCytXYACwyJoDsGA9rNJswhj5noCmjE5f/dpO24tQZH8OLV0Ss7nDqdX
8T+1UVmvFdU5H4PszaATbfCXS2WYwWQX+ni/lwb65mqE7JYvrKGUHSRdRtnMFXqG8NHuI18xMKTG
6026dGWQReGK477uIPpN4iVjHV+amsOKck/tbh2LDGBLDbznU57X2wmwwtP4ZRXUvn9T4szPfS63
7/1Z2tF5sofvHhjxyWBjX+HgEoUf2b9r5L8cBR9Mkyaw0SJbuWaDp6WZFX4CvVIjWEO2zCc+iHcQ
XSgs5Ra1fd/hTJQ7pdF+fTl53fkrsB7M9anS8IuF7bAtRPrD5kHznMySru50uAeWF2E05rSqqYQ9
n84UUohrwTa70xSIojjcWKFLsVJvrSyivHDmUx201VbMbj5ay3AT00yKRQ0FLZgP5elhtWaudrc7
5KnAhlVc483x7ARJNgKzS+ouWgN+QuLpM8+hD0zvnqIFwG48m1JlkLlHnJuiRDR612bH4KYAuzmy
zmktZXbwhb5E2FeuhNQ2ZjXaz2qa4J4YpnbwPU50li+Ejrap/KjSoQkULVeG4frM0COKmZw3dwtT
Y0o+lif7yPf5/nSbC4GLyOqcHgR42t+lFpz0twvBaqSW/QTHsFqpdYGCbhadeX+X7GHyq4cabq2S
7nIhtd48Rv/nvLHXmoulZTMfeUJYy8xQ57zDgIV7PBzJgNXOBY6eh8a6fK8CdwUsp2DS5a1qGHQ+
qia+aP7TXvPmpyT9ff7sS7vJ9OReUMXFs1eb1wGhlX7lHIS09ZqxK7JNzU5pY7MbZrY/vTLtxK11
gNjr5UZLds1riwUVEZ2FFLu3UD8jy67ToPMfwE1wCgv0vNKgYBYZXjoDC3GFVZ/5NikdlHs/WXuE
A4RfH98U4lWwyDzQ2Ssv2dADZDhP3sh8J1wZMK+TdgGx/0/oWOIc2QLMMrZUfimQVRw+EJECb6FX
VDPuvlJnV8mB7ITTz57KnOOi+KqFSRD/trlRwnF01f0pRph5jAKroL3OFFVLjP6RT61dXJ1TRhEQ
px9yq+sUjAahDJogmLVqDM7rxX9n/90o3UkMyxOF91RGe257gvChBU5ttvD1HZ10r+yUIxWEib1B
OTPxgDxHBjKHzsFuDVIdyCh3M3MgpKKsdAIP6skRQzps7+d8rfQwI5buM6dTuwr4IxoNa34lmAgR
XNv2Ec4G8Cl6dUdA1g7h7QQJpkCxhZbrwKMizpBZl0svYsrx1CZGF2Iz/QiKV+aV+m4LN5/jYcvM
fidLavHqJwi8oPWvL5GyRd1WqPbb/+sV0seo65h9fKXddAXJhyISZI/HIz4t29EVifY452IhCIYw
kYdc6eAumYKNPqGuHYJw0YmTTumJG7JWfSFUNJEAet1J6YW5JNtMtGZpk0EUgD4CjdthrOI0h9q5
ogkmzfj4pV21tOJZnS9S7iUNsjen9Re4nsPp8VmzuhNIphSzL7sE8mr78U4vTHFFoGbIPtgJAzZd
njpHrtdzfAhrNHhk7+kDUBZuyvjrHqgC9NQNX7KrXTsYl9vffkvsaWMDhLiW9bE9mNZkBbVP1uzl
PNiSaOqQNnpNccMZ8Dv0yC5OJLSl886lzNGLuNzeelmHyUQdtu33v/7LqyFOqcA5Du7H+pUhfYRS
FFMbVsIOt7e6b/kXs+P63crvqOOBX3v0s7trbil31xHx85c4WXtxV8rhFjcUd1iYRaKdLww9YHcK
qYLXaOPY5MNKwOgnBUI1EX3pH1F8JrJtg8lvI4j81K+y9OxyEWWEw+X9Wu38xDcYRjgAhIvJs31j
z14AQMN/R0HJLsO5BZ4zsmfNF28HlJHud37/8f4o0xahsLKxtZDNP3hAPgm/6NbEPjj7eF+5VJSF
g33dQ32w2lKTCKwgm70SjLQ28p4a/Sd6/OCJ+WmAA4tpyeSnHgj73Qa5a1lAP46njF+QPuAiL5GD
brg9PriCmfn6vBiqD7A2wyjInsOzmjWXfUEQRzl1hubv8edszYPY7EfF6jOnQbDc6yp1Z4iJkxUX
Lx6v07axzsTBa/AdmGMx/374mTTASgLRz8+5LH2RcWRf0NJhb+BvS1JogdC5iLrSR4pzxvD1VAcX
j+e6v4hkAXKoGbYKTQTYe2HbOP8/R0LrqExooTp0Qid084tmZz49aX8i5u8bzDrzbs01xOwFa8zz
G+MwismQhlpjLkju2EfRmyVVhxPQ9cdXHb3afTvt8bPCHS6i8mE8y8ynTAeIHcJHNVBzMtXogk3x
7wkYgmyzR6+6q4OQZpkTPsSkIXYXu+Qb9E9j9W0ysZt9AT8KmvyXKoxDEZH4wuhceSRkqXj0e0qt
xy9gCMKTQgf0Zym+dJOBR9ZuCRLKqRrOjzMvGDMLgna8R8zIM0J9JNdb+8K/WPcQF4Zy9f8+bspw
bbMJB13DEHTSFrfGlNY6kyRFZ8TS7VC8C8p5LBMrgxmwCqOV6oN9MniVtsaWSNzMbmX7cy36gToD
Cadc2y8Dbj3vdyn2V6i574+8xdxxR/PRFSIy5f7EmG4zxEU4zB7hgRPcq9krF2qz0shG8mbw8qb+
sKMagjsVj1poMYgeoI20VxXMOTjg3vK8sKRJm4pRzYM8JkN3Z1jqZeCTtE4nzW5IaJlVpHyG6X1b
IWPpwH6Bh1m+WSdtZghjQe7ez+NhLNbUhpPkx7nMPLyD62vMq3icoRvwZwJ9UMKGUnx4rxGgy2U8
S6V2aJnFnXrUIrf0PuA1htR7A4xTHmp1w/UnvLiYliO6uZsROpQCXFqQL7IAl0R0BReSviIzRbl1
OJMHYDWg3s0VSLO/QQ+/viKQVRn/3b5ilIhJF6IkkH2WioOMbvzycNZB/4wXBNGfOd0bb73jr+xC
mS7RfdrFe1Q4b743A9IPqruuHCtZOIvm2lOFBbnAHfRiE8j5QVSMSmUkxvLrgCtiSrwRpnGVHGNZ
83x5pimY2gB5BlfW4dFoFt6UZaN67a/QtBpjzf9Q66TW5+8QRfhMgUKbt963fSdOlENn8JFvfk2q
Isx9oOejqmqTYBqlxav4bdMW/2MkUtpSX8HHRtyQOKo9miksQkFBS9j7TxwoJQfJ4+K93KOP8dQ/
Jrrl+Y4J4a/LVzof6b7ePtiUChZ48fn/kq+A1b+upH31EegTBiDqvL60B3WPA8rkQJWP4WxdMqzx
9FIhbEmWxVY8dgz8js1SsqgBU3ksLZjeVDN6EazaCcXFq1hUABblVvPxMFbgbxUnXTV5INQmHEip
pzDqIZ3blnLgE9v/YLOCCwKuE5IZ10izntvYGiVHvPCCTPG+1z+XkzfLN3hb0ouhNqeWnRTPmH5D
+HVYTzJyxDYWK0oB4kiubzD9mHHP298t+V8ENDaVshL6ENtQQ94bLjXu3Zs8grXAJhbhsFOhZ1Po
sGKy8Oswj3Eqh0ZiMPRJT0HKwzgqDhA1dCG7sYlZAy9ygcX65AaoA6EJ2BYuIBK92cyk+spIQ2nF
Cd5WTmAMWMCpL5VmUz6RTaKpn0lPSHl5U6IeA3UFrVYnox0N8lBtx3gV5iUIrGQhkzxovA1V3uVq
yq5Rzt7E+Nd/TECrbI5cyYHQeEjvYMsyLXmedIFDfk8E4TafGrYdCgZ8413LPrseMbjXYlZI089E
RV7tPlVu8kh3ra+bvkh4hHFCegdHhUJpkd/tdmdDD0qRdmZ32M3GYrDqYwG2DXtyiDNK+bbDiKf4
hklqlcKnrwAHgoLsXYylVD8j1nP61zgXSm5a0QvbsNOm7C25BdD2zf8NKQ3fbuY+25YobrLebpjC
0kUA2HktiKxv8GjAqTYzY4CJn0mZiuPDkqAbBnHsrLqc9pzgj6ie7pqJTSkB9PcZIt1GFsbZRT6K
H3+5mbAi4IbjjHXJJS+1mik0dVBWZtrhmisC6yNGT8rJbiCrPxr+ZQt86eIv2LIVFfSpDIWrZtAs
hdliF2U5Ox9APzoIJkpsgepspav+Q2DcBvhrTV+rVU+oUH2FEerNB8ia1DJ6uPud3dwk4tMJSDZn
osFSf2K5pR6rEAdHGJZgNAZm+hhgLm05OA7zkC3UR/ZT+QuVfXEJTt6stGwo/O4YzUzXKUISyLCW
r1vQYZZYzWiLpCz1Y+L0UR8SkOY69jVzwzJFgmE1rsLDr13Tzq5iCVma5NyaZ4sbv59KkYZmX4Us
A7faGaIp417wQoSqw86i4kRMqzPi4EoblDo09E6pq9rFgLYrVlYXv1nqoMaeXFw3moufQGx2xVUB
jIgxoHrdASJoAxW9G8PjmAhUFXaOGxxdTPJPXSB3tzYm7+IkDL/K5EYHSJ+uWLwmLrn0/uvBABAU
/o66htL9s3N5aYROmM8iKen0H263bpwpvAHr+6X0hCotHmZ0tCWi0XYTxjgCrhvQj3KdEZKYViyI
FcDUj+HvE9HvFTeEpW08wePVa2FaC+VA2/F2TYIxzzSBFr+dhsvf1rD8TD4DnhAWMZg4H0+SLPPM
sq0LHWCryOhxD556vRXNh6iXgp7f8tWEZzqW4ClVg+gD9CDMG0zgRTV4qyOv0FRPKfRFQVqic5m4
2JeTInc2TffADv5HZGlYTPWlXbdXgp7RcjqJOYM4OTu/4kEg52w1ZBOfxbBuT71KcXcJjeCaSEWb
TjYFxHvOPf/YoJMMwn0EXb1aR1x6hce36K9ngLoSZvyy7dppVy0u/WcvlMv4UXDdYOpsX3zVjj8W
LW5kDamraRM6gRFiK391HB9wAuBXm5aH8l73nmszzjAadKAFdvZhpJMUQpzS+thV7SdPu+/eVlbY
ywVI5vmJl6a50LZWpf/JVmC+DD6KULK6dfNF1fO7bo+e9/ytbngwX5q6/iYZ80xN37q/7kQw2Lev
HphlgFn/SEKGL+6JNRaJiUTImb+evAdv8rD602VIzw8CAXHuxHi7RD3zO/LgR5yNzKZRn6oYrdxZ
TkTYh4eBnJiFrhmNDg5/xvcH/5AYd7fkWO3g9kmLZe1kXJfxkeMgunwb6JeugfpQ4LjLQyElbkHj
yz5qHplqHdW/SAkawuZZwv55FdE0dTUQwSsFBz6uQ0ab54Aml2HttBjliCtMABtZLJ6IdWQQ1UyB
u3Ms3a0JR2MkGrZcrg+A3sEVa+mOvEAXboALCdWfgrJAfLcW1OjV7dBCNWmH6kG5cAbsz9/3LQ3L
oxIwksbJhlc80vDj9cSwQr1Bfp7uM7twjlmq56L61ta80X/9k3edwbV/y1Au13MYr5c3HaP0G9yP
zgR1+Fvrxuhis8NSfvbYXP1JDsJ1G7LyMGFZCyPr9uFAVsq30TRGIK2WYndF/hosA2ZaWOly5b65
jjLgq+hvuO7Sd6a47vhd6qH/6J3RSeyXI99NYlwzJUgdLsxhKS0zIqAdblMneQ1NSxqwWFourJyC
5EJpQyKvimT/i+baNZJ6d0Foj7u79zPt7vNhpQg9pRc8CVQ/M/FD/y5PYtQsMrjRC7bVjm5qY5ky
whUMsqs/GMpRo/WNaU2nU32N7i8SXPAa450iALyituRn1BiV7SgoQToz17DxMVuDgpiBdRfxdkE+
QE4Fk2hExE6o179iAkaRaDlTB9VxpYj2Xf/5lwFBC5bNI2BmJCTXYAEocSt8Q4OmV57TZmmU/G8P
JG8WBkFde4Mw/4AXGM9w7fbbwFDkIi0LZ/7MacVQUxz6zaQZCue0Z5L+htRVgv6rVzypNtpAh/jA
s6N8IERKkdlr3LEBK8rDWZRBmIND4nTvIj4A3otqPmxKbqP6GuOs00hkon0XxTrdjMvndHRg/12D
039GJTlwkpxAd6755sSz2qwkUDV95EzxWpG4mTe0Amt7Khg2t3QHw86PWv98mGfMOfCP5sXCue+v
1mhJIE6n4roVHf8E3HMVhW8h2zt9cq56W4MPRqJ+fjDD/xiRCRUr+UEkwW5ukPg2cvhgsDFJIdXW
+Y0ZjNOaRy+019G8ZOKXJ3ptpLYGaOlGaf5Ln1Ock5NLshunYlGKiiVFdpXrLcnSTiFph/g1MSaI
De+ReG1tVJtHnTWGoTqjnSiflt5nNlbcyhvVBlkepdJF/D84K1VK9/9scgRh+pmVQwKWMrKVxID2
DMbGjcXV7q3frNOp+L2ERpX/8FuP1w5+lqjGExIrppbVfphwvbkaEfU0CJayy/YWKMiLO15bktlw
aGM6oUTE5Ac75RSUYCF7SKS8Wt1D8uEnDIvCfrQHTLatsk+FgSmDy9WNo3cYRBnZRKYa4Cw6NJoc
/kvdTlLXTXkn76dqUPGBxok7bKGLoEIg5BjjZYEv362LFlrqMz+V5wVPALGyi6S/aOxXSFvZOnaY
k/iptWLFXrrffnd8UhzHJDTaNSsW6BMccUCqZp8aMvbysIEPZFNU07lFUbnkRNo4v/4F7QneeaKW
QPTmeJCktHod4hrGhPSya2XKHJAt8AeOy1nkUGoVC3wDTaG49Duo7p6OMy4lGddeDbp+eLepoFV5
9/EuyRGzO8J3gUIFZBEBAPMPSjIBJfS/gSNy4OiZ/sP6qAWV9DfIlRWkCiGCmmQl2vswVnBnZwq+
isdxqYoF6PTSj3ZvLftEsJ+8cynQb8KpFGvxJWhbRtH/piE6iGCmWnKAjM/sZ9GCC+cVJLrvrzOP
btOGoGYGCEu32rjkN3jVvqPSFnQdvyyPsLd+fBmQaVqdWr1/NZzA0LNPm3QHDUwBuyqXytUmP/Ws
yehdHl3WfuVv8Nx97X9rVGP6XSu3StPmJ+lI6cQSEzW9k+7AK8wtm3MDlfbGG0TW5TgEyZ5XQuRx
Z8WNcSccWOul8B/FGtr22AfCpztmpH10yaWNVW84V1SlZWVQgKAVRxzHnis7o+8x5ggWfohVONhb
ePkUGIwPokmhyIhMBRfQXWaU1XSenxZdObciV0PcqZwIVEjFhexh32OxM69OIlO2CnDpSD+rPQck
rNBnPRTCq0fwy8b196PbPZvd4fX++c/lKf1xcLR52PVOXyb6XSs/c45zoFbZotO/Q9LCD9uK1pll
QjgnvWQ4H5cAiJs2PP0l2mDb6BNJtGbkNE91y6Z+odHu3rXv4PxrPNUs2XLw9on+GQnK8ZPfDPhy
D9rmNui5Nuk+7YR+ngPTKKB6fB2CsgoljuHfHE6RY5WIGM8lreuRE+WzLbfsU7yploZEt9TV0m7G
M4eUyNC/36gYgDblQn/rvBnA8HYreh1Hokmjyj184LYTFct6xa5+Rrt874cdhViDyCuoF1joXHsM
uOlKi88mhXEIryAtxiP0LW3oFRZiNyWU10hAvUz8Vim1q3vQEzFUaOIVTTMEmDYLzYoDVET6iPY3
WMZWdCk8IU6YnqePoveAGYclhaMJ+Eeslkyob4trx3pPrH3wwxajkj2AGqM1WBzj4HYHxi7tbdcu
w+LdO/6H0RXN7Evw2O3cpLBK6rOI02VslN1n+GPqHPOt6uDVuoTB5KbU2d2o3KWCuMq+cUIQwLaQ
UIBoXcjTuTI9cOyZIdJGPqWoEpyt2umt7H/ABV/5QM9Z3EjkfEZyhN74mFHOFpOpXux5ly133CDr
Nm3NHTDW2CCtPE9EcI135JjL7DSCzgGkPD2Oc1xy1iUP321zAObHX0TFuFJnzbFV/fX/RkMBcSrt
MDQips4+f71fAARjwWfNNFNui15opnLTWwkJh98wFcsvPVyD8LRRoBcnG88cANYfSdIf++CAcnSB
6hq0Bh/0UfKfLYJlmPZ/SB2XgZILqcZw+62WEpuCQBKecmim74OQOxywQuIMQpgiNlyW8R0IAU9M
g6WR4uVSFxzsWa5INfD3R9Zcs1EwUwGhe0IFX2ufzBwHCmFS3K4cjnvnN8dtYIImhBUQaACl3561
8lSomAgfR6bbuLSmpHE1e/Hj5u8kJTNy/rC68cFyvtiApVkFRDDk84du8sjFOeLjHi0DAhiORy+J
JZpx8+8/prtdBVESX6qRlmlSevwn8mUNxfHPZSzHdEn6TErvKe5zMpIAd7KhPGPlRQwytChrooA5
FUJBTXJK8y6QgevW057tLqrNRpbjKBo8oAekQ0dGtmur72iVLSBe2O9kVeTFiAleMDqSPjcN56m6
qyA46d01NS1eJOsgusbNjKzvA0X+rgTN61zkyQZ9SA25e5suR5dqqDQSCQ9x3vZuTsDGOMWLYgh/
U1knnneWG8UEMfa7Qgq18FX2Yx3fFx1uNW2+BpShC0+Z/NnKxIzChcpU7wVeyWRKDo79+SInByYb
XaVioLkBnaASJRclQlcyb9AeyHIAwWhuhCwYrosFuo6VpTH6ePmx4dXFOFaN1pZYVy4QrWt2tcnj
xugxIbrjFSnYM9BKYpkT+tMawi1UJpGTvZAagvrvFCBKg53N0LVRXZLzvKRrq59WGuBUSl2McZ+i
MfAzCurge6ANGbt+pNy1OPHBy4RczauVGbNH9//GDoTzs0uziZ4ZOsVWNGnvw7abGFFAST4E03C7
t4A+IBD+WGhOgCs6Hjrnn37OJofb6vWeHZLJ0oUnsefxCwDrnzlBuRB6my2n5Go8Fa4i+e4Hd9m0
7barkyosqzwKaUd3rF3Pgs4EvubJlvhxF/rOVQDudeyCQTeVuoqcn60xrNDIH8ucOHp/7ZMv7L62
A7C85wpjU/D9nDHdZVFGUo+SFlIuyKQkTjn/kx7QUGaVjF2857spBN0NTWmtFZbwX0f9y7qFeSCU
zOJsfz9rulKy3CucwzqGoE0Qf+wfQJqOZ2g6VLCQ+ZZLTXGGS1ECedrYgdutpKdJLBYizWGHXfHJ
VJakYYfckj9YU3anYyycCv2sMayIeAlKbeJHf8+eKOO1TmTdJ3m7Wv+Tu+83T3bti/MKoUyWKnuD
x+dKmrcUgXbLL0rCoxquAOj081I+1o31EDxO/+q6/g9mQgAVkOibLOMvoM0GjB4OX1RrHeQ1q2Li
m6D8HUIqQSohQkBeTcvgkmCkhewPQqUpZvCrJ2N/ou9IuvSMdMIsIaAAo4ksgTdCUroMc3lHzvD1
VAkkDuqB/cA95SsVbpxDUNk9doupdsJe4BeDvWaOjhetMej/DKT4PNtATeM51nmrA5+TuITNmEan
sKQz0uThF0IBIEJCzHwOCZjnd1KJFyJWCFSG2J9LHdGkTHMrkSZS9N/h8MfCZ7k1cjYix073H+B5
oAG1eENu/K7xt3E59VEVT4jC2097i8eyZ5r6GZRMgnCOPmRfp29cbkFVblvAqKkCUsdIAZeDNvAv
gOidHlhH+Ms026m5O3Ar2IRyoxyOO22pkK4rihz6T3rWX2Dyuw++dS4wd0RppCMYdM3I9fcfluFr
KFje1NBsbDzFD64xw5q0flHwt5G3ZZ5gaNzV3ZWvRVJVru9/69BlLnxhLJlI6Vb3jXw/omxlKT1U
ZPdi3EToGdEBb0UDIxScwsQxOuluUzAYnWSYpdcT3zeUKXzepcX3zoJqhLuYijqC1OFy9IW2yvMM
X4n9vGafjrTLogsfm3xUWGHIynuSqkUzbEb/+8Np17ogxEHRjavbF4qwlq1Ma6jPESw3eRBDODWg
2RVVgQ8904X773SfTYvqHom1xAJiDhb5zuL4FhpEFiWGIPKyRHpvCK/Zc2EOa1klom5J2n4vbo+B
ufUBeZQHVz1iMWeSTIfPUhvpMv1+6IHl7guwh0fbI26m8Svq01rllonEVWJ9wjns7FTir9wq8Jmn
3kNljOeFr9quzpx1stA7SUv7u+5Ac4UIUsbQVmnD5/INaNJdJIo7gweXpSyA2fwi/9DXMkJAL8oi
WF3tKLeu0RYSkIabXdkirC2OLirEU46Dn2K99SzG8bKMVWARh/YXbj5sqkkC8TDzwksRic/cC1sR
Ao0SjE5rnSSGJX2DPLmKUf0jNKhzFC6E7Pa5f065wfR1JAmEJKb5p//4Wk43GyY5kxIBGnfS3jcM
HwE9df80F8TUUTO8boBA7F64y+F75JuYIIaymxPA1Ylr8I/wshl/ey2CLfTHEyyBJrOoq0WDJsgv
kLDCMtUNkeZfMaoJ0krcQHFXipK8n5DEdEXpVDAgRmgOSwrwyYUwWZRFYpEG6faZ0pTqWy5lIrJQ
X7N92w9gkCb22FZ0tpuQ5kCb2OphaNLVVvD4uztujx3mN6Fy5dpPnCsA3vCbNuzSWJ2V8W2wfLql
FY67DTYUyCUvjWt+SZnFrutmSe61/H3rLWyukUUQWBj4dJlHokt1vOfGiHTetCOUtE0xUz5khzni
cxBbdrgDwB9kivgxePj3X91z1TQpgI8uzHgVtFYjUfTc2EvV2tleZodmgAlD9HCtF8xHBBuMJPwY
CVbk01PHegqujQaygWZgm7Z3n1agLfIkh8A0LDN3vCcpx5rY0b5BaVLnKeI3n6KEQ4oy6wNlr/eh
1diFIlhN3wk9+WDPW1Hq8msdzQPRj+lcwejWhiRQMlb3BVieV+GiKd//ElKJze/DmuJjPRx3rldp
BDY0Glft/9X++eOAHAmbe99r1dJLe7+vqbzCwouPCQmK3eqnNZSe3sYDM4nIT97SFB/1rOjyAa16
5X67GpsvOYaoaLWnfXnCKCb6iZ0emveo9NvOMPS/s+444jFgqiN1DISg2abWmeFuPErnrq8p78K3
V1lbp6ynCmkYYHRCSoiJ5bt0vFKAiErN8HMpIRFslvpTpF5OT3UopryibrXAqu9CfnMGTGz3Np58
NYKK4+scEzPR0T+sXsJM0bv5CWgD1/FxbjTZeppvVMyJK25UPbKdzK8fRKGQ6DzbCoHRL2eq6Usc
Xx10fkp92S8G1J0pqph9T6qWItPl7r6HQVF7RhcLhGkhky8ZzdfVtMKmAzgExEsQWHhc7QMdnk7j
7F/EXLssmRGcvTCUYDShnCsO+zHggSEBaIDI8JWsAjTqbi3Re3PMw6ewzpspc4t41mocp43UhUai
a/aQN1YbkL4jrbMUBXQs1wBIXQPdXL9XDZHMZGuD2WITxxo/JkCTyCMcGKNA7MFpN2SmvFPY0y/t
fLxXwNLIScvFjkju+XIN9KdapnW2kq6MBhngcjAnB1Z+e2wCw0fwIIfay/xS8asL0boR4laL6VMN
Wpk98ei92WhtpTZFarbS5+TmyqDg6ju77tFlSMRy6AQOvoJOgR7+BGCZZGnCspvjQSQD5dRcneo/
oatDSORT2gV6OcbAeVfxV6W/XvHrYOPGx5Ap4LooNPtNmpUHOtf4tEA8VzztuBfz20URVwaptNQY
NZV/L6D341X6ncRZmZAFCueuKXNYK/aF3+l76WYRxwYFT5PsZnwTzN33kZoLdhQoqvmTlkFQOC2y
7HjsI7hloDgdhhreqE6y/D46GQJ8FeTw1XCWWPhuQAgbQk3WmjHDMwsnNddd0DgkV7LY/aftOADg
aIRfW/zTr/rwSa+6H2aS+emnLcWAub9QSfBdt8CgIy2WQZiciSJKR9WhkCsM+O6s8Um4GFnhV0X0
DbAVLXCbp1H2ASRBmoqCq+on8T3KIqCqihQCpxEQ/lTfBsTwTFSSbr+TLoprDNUSrwXho5GaKx3m
17R6joAHsUT3fJcHPHK8j3fg3dc5CZkdtf1vMWMhoHVWfKmmyQaLZsWgzb1NslUcW6WYIUFxp+Ib
XmMmKgbC4SM84mwRmzbG60SIsKlnY6P6sLgki2Fl1HzX1BiC1xTh2kHpuy5JWAYFoZVMpHaq1qJP
rqK1mrvweFNp+KuaSR2JNTlnjg3znHS5wZAoojqj9wtPCPjBMQjQgIQ49ZSZfDPPfsuPIhkHTJOv
nc9TIlEJy62PbuzrTPyCuLJN6AiDuCW7qVzDFQR6sY32LqF88awQNgG8vmvTmgwqYKi39WGbMFwB
kIihbn3PtcOx0+8L4MYd8jvhiyerFC0U0AsaKzKe168unHabvb8HGVHaUnnRzjqlYedOsf9WF4TP
1jtre0Tn9S5iOmRBLmyK/HI1p1MQPeFo3Mme5xPOqgQggtrnWs3h7fovdm11Vp9ext6jVDHgGhNH
c5dbRtEIlrmwQNHIisVcfvcYiWieJSJ5t5pUL6MipYWyZUl7pCc0ZsDk1BkwCM7CKRDW4bWHivxg
Cd3C3tTLRKFmJNdYxdlm5jrYFwa8IPjRkscuAe8kPF3xrfxkTqtKk+kR4BlMuUGrkeJmc2l64YDC
D3XcvVWAupHsAZx2tkTO10VXZkh60oAoPYg8s5yZviWcm2ah+cz5FhltecIY56A27Q09L1W77T9L
xnNUSpAv+F7VBj0ZbSmiZtFIKsT9rzJBAY7AqiGxqC+qMN1UJjFoJihlVf38Aj6NWQ8ZbNUSbdjy
wGT4NOubx3Iu+1EueHe0B+OK8/reekOU6h1ZEeqiG6ZyH590dQHOTNIyhEL+oSLhEi//17cRJagu
bnG+349ab2BLjxUdfqTqhC5+y1DONmHS7aflEwPIegf+UQd+Nw8HIdsF+K4I1euoiJyEl3LO66Fr
vG1lFxIT4xjP5CnV9ItYZXHXfJAGaZuORgo7lp/2yVouRZztD4UxEvHIDCIdznk8er7LNIFrluFI
laqK+QyG1mXxYtyErMmDvlTMrg8igMCixqdIf9RZ5M0CGKdTeSq8TsGvIBMbymJpPzYfD3AijFDg
fbv5N+o1LsPRBJQG4vNv5TQcfy4xCaUSG2gKPishTbPDQwrEuTUWGoWpngqU1LqszykwpBW2cOrR
L9mKjMeMvtD0d5QqikcbndPSwWYeQTZ5SJETCfmW6y6pB7hplFuV7WyE4M3ONSgH3waPHE+XjJJR
WYL6ZCU5YJo+0dwK7/KgvHIREc6jlNxnxJWNJBWrCXoYwsP2yzNlyfKvhKlSVP7eeUH2itohTsnd
APKY7J8eVEHK4XLP0Zf0fqTPA8lcl44jQ2k9pp95DBKFY6UdbPdqLvxopLgrKp5rSOFYpzlm5p1i
5ZDx3qPEw9OJFpoP4plN9mB8h+NvDOeuaopE8YjqfABrXihA5PxmOw8pzlZo+weRSw3DzafeDbN2
zkixgtXRspyPau8UY9Vd1Qf+iEM7eZPaKv9VKryBYFaPnTCpz48xnJptwaBqH5ZPzmEjAaV9brjl
qcqg39i4x5x0KuSndRnw2OsLDY1xJNoNx55AtdkDZYY8DyaFaF31Bbt1zUK7raG6RQreCFYjNJMD
f+aDy2HxGGLgti0dGmJYMgGFumJ7GTphxo+ojqB8VYM/KYzOqk1kLgX3FvQjWt03/5qTqD95c4xO
t8cpjJCUeCiaN0zb8pYp/xmPTtZubBxoTK3J7t5OYw0+y3GPj7H6+m5yJ6Tn0Ctjs3+TVv+YV3fH
9BncCdoo/MDwRxfB2KDzdi1sNfJQHgGKZEJ2c13JpQBTmfjFhGZTx+paySd3peJbTE3Bf5o4q1U6
1f7Gh9f/TVev6aiJMAfB1e2awvQjsP+A7ycECNUm+8m94eHMF8/QW3UHmUI/uEUB3jDU7rAwY0k8
aKNRz9bFps0biqOfY7ZjSq8UZzzKpAfuvPEyLIbiH8cUX/ErhRiM6G+lsL1jcrDjuQASwmkkjJpU
rZSurqIUSDsa6E1vU/3n1Nh26T8OtrA3F2ETZ2k4Z/RXPPculY1E1ZvszhiOZtB1aevGts21NaYY
6xhZt3HC8DAM/MfYb5B+LDvVwc6BSRTXPSa43fpf4OCO4puFba8mAFzD3ftLXxyhVXe3SHOFulXD
tZ0Gv2/KWP405aBE03Bt4JePKK1D16Hww+KMPZP+sVyZ4r8W5mPh/TZZZe8wkxdTGPopab7j+18K
5DQ6kTAnW9CUAxiMY3o3NHKTH4L7NOeMYWlTH2AEYYM6urkNWyAu0dOSgXq3AYy9PXfMxOJZSUEU
DgWUazXy/z4G2q7RhsjH4lJZ9f9JZH4FLCa7Ki0v5pIEGYimt9F/wG33P5UiXdQsghjHS27TeDuy
IAWdInvY+oiUx3gnDzCCcKj4KOy6Hx9Udd7uIQ+WsISqEk7hjI8wgvWnaM1e3ZXNLfVvEU+xlvNV
+5gOWtsNRIfNeSd3uSkEgGvNi2cKrMCF6xRmxoLRSxNs3RdhnV9mLOOYnXEQeW7keKlu0my8rrMp
kf2IIa4xRx4LFW/FZZF0VH0Wr76VEUeAJThrnwiZBitgl+h75dsFCiT7cD/1u2jW32cVH5D8jF0d
gJgRDGL8aWUKCWaaosbOkeyDgj2WuyrzJDTtjFJ2GzCtGfySKBMZDaHHhJpcXKwYPqXe8ptVr3yS
iq7fmCsZOysvtCtuKVopIJoRSTr6j3+opEE/lCoh1017zIZHSIu3lv8pFlxaCsAndYWiKTDZvIoe
o0VEm7cqvm6mQa2E8c6C4gWNcHct/5SxO0TxrsgqAk1rOEdKYxe++yXkbjlk8BJqtt+rj1bx5/tk
aV8BD4m/Z01yFQg2iRMIz3q9LN+mFXPLgT11mGAJo8xrMgvcynLFKbKAyKQRk1F4UI2fLuU6vjkW
p8/vvUjPro1bt7J06Wy9Ubso/A2k3g+BTnCtnrpWRiI5Pf4OJ2jpc9C1SdwXTLiFqAAb516EYTnP
BkjvndmChRowSw6FpunoI+alBu2QRb0oLAPtHuFINpD9Qe1tSxe8xdS339Wtr7F7Aya/y+KqBixG
fL5qI3Sk9/f21PCXWJpJRWZJnPDBLIxmszM4BeNC8pCEktBoENsAZxUfb4WpGrBb9Zo/COJCcOyH
bHVekiG2KcLyJMDMEq+/UsoDKY96JJk/izhscPwdhg2Rio3by7nANxccMuVVpHj0HKwqHtwmByYm
VYV8/LvsYxXpZy3KBfV+ek7+KQfgF41OcimA9roVqIRAvinknzeJsSL5zqaOv4/enxA+do3MW6xJ
Jt4Kop/LEptnr6gitVCqBjy0AdwlvUcFXspiGdzYfFmpaVp6kGCt5P8AKdixc/XwkkpSkOHKsN8S
jPHcJ3x4Cd3NwJ3hrSj2lnWSdPgDFVc+oz/2Th4t6TktIiGoiMi0tE/R66hEx+aOS7TPypMjFIID
BfCzsetG9GQNiN2PpUSfo4fa/3xWn8wxXQB4jr+onOSx3f2hdH7EgshGSby9pBcOYnavmPqczanU
y3N7HCr5PKmFVOhopJEIDNcx0HFg2ZxcsOHfMdzAW2RbSEw6nkAsSYXzUFTt3n6XtW0VYmVFqmcM
Kel43uzV/qDYsyJO2PGfoHio0xc8RHohvAKb58XMm+3GOGcQRBdmJk6/Ls7MuYwHLimpYQVjgD9y
YmADOEnWqLcsSBh2qjxQHlkvaWCJJEizoUvOKqKwhTFAAV2VGxI3SkXR5EAv4+GauoAgLK+reqDa
5GfeaerBzI22jIquZM++syeHxcbBPpv07zaDfBrdd0XsdKuZHoDRU5z/mQbl2kQ96o35EpYNev3L
YGR2cUeryCV41dLEeBFxSZWuJJY9zHHU7BM/j0udG0za6Pd5FTELWq2V4DHtpgOWmccsOrocrOIY
vLJyBJkMbF+Rf6vnjMa7k4kJBWohnL78ZpvUHxZj0wf3h8luqSAdXEfFD67p5mvSSJ3r4NQt2Udw
Nu9LncwFMUiwp8rqNtXZ8eKLiZECy6dhT6FAm05LEbZsBNPgtSqhx8xASNbuMYSs92BiCbAk1/3j
O146srHz8J1I/FAX4psTGJcwi6UUIjxXseDv+4/OfKr8IuNCLhPXiS00CPOAvJcbtWttTJ7IqWhJ
A2c3wFAOjaU6ZdYT9b9HMfFYESiC9cpLZG8iqvs2xcxbYl5v/iXQLpz1eUJ3x6l7SmIrpg8t07Wk
YjeWm+65hL8EUpScfQwOYVVtsTj2NA4jg1xnkTTbg5w4Fi0XXjmoogHvwmYZMBU407+i3CGiENVT
LCuKVOGzx1RdWTyFrxkadoKnjjXVM64XH1EFn3U9Vd74Tux3eiMAv2SRh/s81pe3ygAc4Q6z5LI3
cRRoT9lR4FvaU0OP5Ip9JA21m1PUodRFWnh7vCBfdd9JnIbSFFCnaeRvH95oxTHiIyecLC0HzcDp
6Rf4TMOO/JjP877vCgr5pYmbEzKpBAzNhaiA/BhnokA77h6Xp86Y9P7802PgTqibI2VFMbFGx/B/
Reo24ozS3C1pJvcP84uiHMqdc4GmHmrE81FW6onln5I7Lxglh8DuY4HGD32cf0sTxA8SAutGowJ5
Z8sipveuk+5sysjUJ7JE6qJT1N7Zllgui5gsLQEIsugcY9ruFiIenyN6FPB/T9bN66dZyzSJCzzN
CC4wL18qvjM+QXN1IOk6H4ZtZOPeus23Nm2SjymohQt8VwfCY3LlSeje1Mvt+yc8Vu05rsmav7ka
lIHBkugDBp/FVWsdXEOoVR9Fhx8nfsIUPrtX1TAgHEaksnOlkqYbV1ny/AsbN4lMg1DugUP0Ffl+
Hh8TjO8gDgsb8hCDwZERCKN74jPPi0CHtvdad69TkqGid40DS7rNe99qXXD20y1Fqcp3IwmzSYLe
uggEM1srlPhB3w049WCD03x9MjlH3owbfJ8a91+Oz64pzVbLcDAGAkhGj2LbzdqYFOcGw/GssnaE
rKZa1WRiet34mBY9ersIkcWt/uA4gYCo9hZrn3VnFKDjfm+PC4IvzkbBYxU5GHH6zuApM9v7oFNP
In0WPHT2gxpQcTiI57/mOZRW9ccwD0TC6sSd5zUhdjJId/jsW9sqQ4WQ+BERq4F6EljHfb6Mk6HC
Ih9058AtTXkWOBouj57Eox4f95tqwJj9Bc5vNC4ObJ9429TXbZErZLQZXL0ZM2YuVP1pNKpkjlVL
92aNj2oMvvcPpF//BmeW++/T1DUziD5cwHmpLJwb/kQt2DlcZV69he1Qf7bIKYBIJoSReBGQTsfx
7/mvCQkFxZzWA+RH9sQ8COKcuxtV1zGUoGm0tTzg+qEVzpYufTNIVs6cb8agy8l/10r3ZoOMSJt+
J9OG1DFZIJTIE094HUjcxg9f3AGj4QBhB79wA+yC0gGcq8o4GcRjcoExxzIHa89xVVHlnVaE5L/3
l2T+VwTs1FVdjuC4IKEbYxDOr1fEbWr8JYOMC10u6YTISUHoIssULp+6km6V9NHRr2v5Po6VfpeW
UMJ03OMkDRi35pXuvfC4jUAVBYlR+JE9/Qnu/LAxZAH/Oy6C2k6hDH5ukiSEyxhwWrg4sDNBtvDk
f51nU4QGrWK/MwWi3MWJRk7425J702ZYfIFAG7NRk2k6UC1eMc35aBzE/czeY9fWyLPUcipaI1VC
fdg+E1KJsfV3dQyLyu1ikgmxPVAdlAUtJq3yFT5ubjGJkUoWgA6/6v8GPnDaGmlZfg580TLErbJh
Q2dddH8RLoEHMJo7+nRON1eP1PSmPa/XB+lziwyuJ17oEhEmZAo6mnVZxQTk6xjmvOJ344YeV0t1
+32/cDwyXNbqH6T8uN9D95U2jufkSus78A2w8iaZtUao2msVodNEyt/RxyP4K1RlwMhOGYQ4vXDT
O91FwAbkiDBRJYQphsM3hQ0oS+Zlq2nGN9zRnFnPLDZsFN7bsN8DRt6QHBl5bePEhOO42C6KleFR
I+VwlbnRiIHOSdbYMll8GKnv6yD/C65V6zu6VcYDokH+XCsfv/HnpNbxGaOHGmYKWNf6vT2Oilm0
CPDRrpmlzEGKDtJIdPJ3Zy2eRlYH4zv9SQv9JfD8aGX7PK3qnVoMi7Z8EIhpYWQGWer3+1Fp0Ysq
VHfmjwzooNI9wlyqNrhp2lAhYJoKl27EDXdpzC2l4knWPXnVdJnBBlgYO0jtO25+wjtsSTqx5Lq2
k4LtolqEaS2/C522rO40fZJaBgHMLkp5y15rEacgc7TH0JPMH8oi2NjMEzaCpavx+m41phi5o291
M0L9yHy05i04glG7DujK6pGI3ZDh6listPlVHXqBIsTq83/Uq+cmEUN4zsL9YGLbpwchwcT07I51
0OAIFOpsHUzEKSIfUHaedpDv+3amjl1WabUE42/RxyQtcq6pHPWXflWjHW1/XnwSDdtc7piMUFCv
WKOIiAFRWwabn3MXxjT6whSw2BpL3cXmaplJiiNcpR4zgz/crdZhioR/7K1FfV2LWfiuvW+xZy+z
9NzmJb7t/MEa0TfPmRMxAQS5/sKmBMYeI3cV5gFRAeZeYaT8KMde38rqHOcL7ZpFXbGdcMmkwG8U
bTkJiTZ4gzqkELoQ0/KpSeQxNjDTcLWH25L+v6fNapnoU8kxD24ktqCJMMABub7tggPy0vj6u/tA
Ns/vaKL+QOm7/RE6TuKrPQZq5LeXc7Q0O8JKliqc8HWTcrx0RSf3W2drlDzjdaiwFTORUATmOwt/
dzb4o460HXAIOOCbY46Aykzo5Km3i7GGFtzV1F6f6ZmaHUN/iJUkRbmFX4pZ6ycl+m8TN54CkHl1
pX2+0dwluetYfkUIpq79+JEXjYGi++1s1JorAhcntI1rY/1sqbZST9TnNWU+msIMwMGqVdFMzgoJ
GnlEEKhbYXrBaap2GUz3wXK27buZCvcRoIdF6sOvbtpBA3g1qmmFErAa09LYKyNQioCY/AjWABGa
eyVUEDqT32/w49LMTLqCM7VDxcm7ODI3KhqDREAdmdsOFsVzWsGvIaJhShq/HDwEbC1KzCKoyhBY
OrZWFm4D/I6fuLds7PAOlYOyoe9bqCEYIhbnihBtzWRgpxzw0Q7Hh8U0T6cuPHINXgkA0782Qz38
MDZkwPQgEIu51A0Sgl983n90bD7lhFGwMFw752jrM4d0mHxzMA49jrEeFQbwJs2zZf9Yp3a++gIL
RTd6yHCenVJElZy/G4K+ArOCA5Rwv0xzRVg1Xgd95z3pcUF01TCVYvPxzQm5nivVvVkjushCCgeY
YMjmK+OC5f4d7Q6ls70mBCRcGUhLvk671HP3AuwAzGZUfyFr6vZVhFXmpTu5v3z4qm5L/uI8PQZN
RAkMuorHbzYojWV+bP5jo+xBqXD7Ih3arfXoGQvCpKXnR0PINZOAh1P878QjmNWefk79092d4dDu
hHNHj2kIu/O1vlXlUm/XuKEr8NQ4EjAKvgygaNHa8/ULll8gaTQsn4HRyi/L/QLQdWaLc4dUUJLk
S6zgBWt8SeAmDddnpmScUw41Ok7NpFmWRsCLadjLmCd+I9/5UaDLjwvuiJTmcVavhG8PrERIQkW1
Zd9JvJ+GlNYNHyY3HIzkqU3riSjDm2n5vnECPMGG5eqSC1xciSTBlkEeo6r6zBbFm0ZaAxuDXTww
9hTX59Nrqp/iBGByi08cY5fbQiA60kP6z756AczBg6/agdwyMaFeMrg0q/fQK5jNj/mnP10b+bzq
rqQv6Ts+18mgdKWzIsBp7R9mG8/lVu17QR+wz94oIMN2hPsnvhU1od5SvIL47WfddvwzDh9qLZuT
xTGXqRmH2S6rUOFJ26U4ugLTcsg8hft+JcVb62gRmqzgGk4GFvdzp3h5lO3fEov1avNTVQIBIoYw
zJ2kj6Q+Kon1EAiOpX/5x0SoKXOkot0vcT92bnPZ9CRZ3RtHrBgsuTHtFJlAptyMJ48AaG9NSkg4
ljR5WlyEydSwVjGR2LUA0YAfj/VB7hyw19kxTLF0zydmMkxaigQgsVT/U1OLDDVQP8RwuEUhZBRM
q8JyNcEe0d0gSHC8Rd9P/Tobi+rTnf/2QR2vt5krB1BHfiJWC77aZAF8r1HEuSrjHP0GABA7e9ZU
7wmtg9PD7W3lBwruqhbFrDXC8/dBgg5UI+XWObOWQpQVzImSjbtK7FtFVaxjvjFIjf9Y66iotUxS
Xqr5ZVm9fZqifcECKtxYC70RS6Yv6hPDo6tNrynubzL674L6gW0eSwN3DYtyHCPQjMxlYNJkiQhx
8vqJqqgWh/LLEO9fL+Q72LU9stJtvY0hmSBHpNBEM700lFvN9gqbU+o4Z1mBe8niGLkhbms5WdO5
lweqcfAJEebEfWho2Mc+I+GR3dLtsU+Oh2x9Ax38f/ovLJiaHRiU0tvubD47eKvLU9NyNWSfetAp
4+K+6JxQODiBsZJK1YlVnImLzpDsi5AauG9JiCbZ065UKycgq9b+9+bS2K6kq34RdvMQT9YmxT6A
vD7ik07C6IUq5j8fJmio7ABvAq6qPDnbz6+Q8NPhTpwqh2lPIo4jl+8CBlYC6vJA1cXsFzWJMQmb
LFwWgngzSWytdpQP9INkZYfoy9Okb0aUEwyiSZep/w/OksurBpPCy4vwbI3MsuQnpJ2gin4/5IqE
cdlQRS+4RebOD6ysIfYckyU9l782U+50rEQcGWpOKhfVDjaZeBlofPEmWAm6MBfsTSviBE9suJN7
rPusANvlKkv8k/9wzXOnonaWQ9ViYojzn7l8TEpoaeEwy2WXtZvW5xZ8oA1D+XwiH0aSINjkDB8L
/O9vkSeHsD5v7KKs5m7gNSepDaoxQPT1tt98nPbBKReV+n+9DMO+Dq7+xzbjLmuzUXRXQTa9byiM
CBBKyTiRFKlGJVJYXsdUGL81kwhjJV2vGykrZ+tqUN4CAcOCumc/y4LvgTyYe+msHqK1klV2eypN
B9zsIqapvbhSW2ViOws2aTJbJZlmcFs5c4mHKFGK6eIlWlTjRckZojSogiabOPfhDB0CcQzXSa6l
Wguac3CIlmWJKbdDnyq8+y33WutmiPgJoLAB75oWbP6cO2cBR4e7m83FsvMTvZJe7LL2lMhF+weW
uklIcpJ8TC3hcRo/yGGnAR69sA35wqhYEfvjfT5H+xSrHIFvqTXEwESTfwi5TaT/YpeSw8pUMmzW
hhr7u4oV6gGnmY0A1F4e78hTqveuBKul2tL1/8bxaDaEmfhlWDNvVSAeJpKnXD8PzWyQ2Wi3Hlt/
s5eY8zSRSq+F/pdg1tPpVtTP6Vct9ncrwapldFMYffdvWJo4iURUMciIDos7pM1YuVq93TF3RAe6
hOReKSpSq13H2600d4DzvWGh2WrbNeRNMmwk/82RImYbPfJLc5egHMZOG83cH1kpjvP7tJqKXQ6b
xQt2aspvCBchW/uBI5KSMsFdrDgpGFoPfckJjThXH61s4LgGB8yAvHjEgdojY3pO0sy4OQoue6ss
q0lFwlb9ksX1xwcfdApkIaXUB/XaWI8lErwHITZQdLFoWZNuXs2pCeXmYKLb8bNdXEhkphScfWqb
9K5SZ4IVKyXBsptoherVnZRe9kOH9N/1UiEN5gpl2jqTz/TtdGbF2vdOEzo3V0fOW3FH1NBVlIwZ
/SAOSi9WvVsWkb7jBsVCFT7EI/+B/INvL+y5Jgg6iE3hKX8O/mHtWdL5W6uheqC4ebNHx6keTTgI
a0VHEjXvyzpp4NUhFnGOByawDy0cZmpgU/RtrFakY8eTK1xLM2xgxhfdNA7sTq1PZYHN3ijL1/c6
5Kdw8ly33Ki7+A0zfMa1SV4k6R6HgjQaN4tyjvDeuF5Df5O6BDzWgIAGDtR+dVjdCa1eI5MIAUHg
yaXHDYuyZQsCPO9iSSAUAiPlHyxmQyF/1SmcuVS2L45b7k+i3MUMcHS8A10Hv7LaMSn4xRgrTh8h
bdTelsgWwAN8ZzcU4cUuX1xbFnPJFbdcyDuLhw1pE/QrzNnXDcmYkLrH0nlduP9LuQo24oCL6eDc
k+9Xdj1kn6ohES8uiCUJ05EPAoEZAzj44yzzkQG3v8oSd+WO54R45lVfNVjN/GpiI4RbH13setxL
kdkiJuK8zR2ElNEDdbgImCFVqW87KGVMRMLbLWwPScfpH5ZHBH341kvleF6IUUXcK2i99gnFyKra
o6FDgPiUc7DFKSeUgwB6PGpnjZWuFkTiFT2+1QBzJbMSLKCGfCTfK0QW4fjzyxkCs1tYCMz7LNoh
7cphyaqcSAPNbOKFlU1pBxc+qhW1xegKklEsN42u2qOaEBIvb4RjYJLB6TIXu5YL8/fDG29m8+aj
Ajc2IYcO0ZrFLSw/JveuSZ4WVsJt9eQtWd1EGG2ybrMliplbIGedo06pa6zwqhOki1tJ2E7KLyU/
TN1g2s4Q2QTX57OwyRGGI008fWd4WbipOiq1D+XVfpTr9O72MQ1FtTSoFtrFW+eQWO4RxeoUdsRz
a76F2OX0vQZJ5V0Kis0mlvCt6CGVxe0szVGLUNd7zzY9JIJvIZuIs1cR78plzVoaFkS52BQ2DMTB
6fNQg05Bx5123LVJ2Q47yA1CgVuc3ZH6yqSmvPCG/rEXsBsK9PF25v0dYnS8uDETTxpv4WihAe6J
qA3NTWlSefxa2u8t8zP7dUbhj0R1rWi0e9fq2yzzxNWDHTBuTalfh8N/HEehCRZ8+XwK1hDtivjm
+DyuObD569XskVAEISt0hLLmFZJCswRN4dg=
`protect end_protected
