-------------------------------------------------------------------------------
-- Title      : 
-------------------------------------------------------------------------------
-- File       : 
-- Author     : Benjamin Reese  <bareese@slac.stanford.edu>
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2012-11-06
-- Last update: 2013-06-13
-- Platform   : Xilinx 7 Series
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description:
-- Used in conjunction for a Xilinx 7 Series GTX.
-- Given raw 8b10b encoded data presented 2 bytes at a time (20 bits),
-- attempts to align any observed comma to the lower byte.
-- Assumes GTX comma align is enabled and in PMA mode.
-- Comma is configurable through the COMMA_G generic.
-- If an odd number of rxSlides is required for alignment, resets the GTX RX
-- so that a new CDR lock can be obtained. The GTX in PMA Slide Mode shifts
-- the phase of the output clock only every other slide. This module's
-- purpose is to obtain an output clock that exactly matches the phase of the
-- commas. 
-------------------------------------------------------------------------------
-- Copyright (c) 2012 SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--use work.Pgp2CoreTypesPkg.all;
use work.StdRtlPkg.all;
--use work.SynchronizePkg.all;


entity Gtx7RxFixedLatPhaseAligner is
   
   generic (
      TPD_G       : time    := 1 ns;
      WORD_SIZE_G : integer := 20;
      COMMA_0_G   : slv     := "----------0101111100";
      COMMA_1_G   : slv     := "----------1010000011";
      COMMA_2_G   : slv     := "XXXXXXXXXXXXXXXXXXXX";
      COMMA_3_G   : slv     := "XXXXXXXXXXXXXXXXXXXX");
   port (
      rxUsrClk             : in  sl;
      rxRunPhAlignment     : in  sl;    -- From RxRst, active low reset, not clocked by rxUsrClk
      rxData               : in  slv(WORD_SIZE_G-1 downto 0);  -- Encoded raw rx data
      rxReset              : out sl;
      rxSlide              : out sl;    -- RXSLIDE input to GTX
      rxPhaseAlignmentDone : out sl);   -- Alignment has been achieved.

end entity Gtx7RxFixedLatPhaseAligner;

architecture rtl of Gtx7RxFixedLatPhaseAligner is

   constant SLIDE_WAIT_C : integer := 32;  -- Dictated by UG476 GTX Tranceiver Guide

   type StateType is (SEARCH_S, RESET_S, SLIDE_S, SLIDE_WAIT_S, ALIGNED_S);

   type RegType is record
      state                : StateType;
      last                 : slv(WORD_SIZE_G*2-1 downto 0);
      slideCount           : unsigned(bitSize(WORD_SIZE_G)-1 downto 0);
      slideWaitCounter     : unsigned(bitSize(SLIDE_WAIT_C)-1 downto 0);
      rxReset              : sl;
      rxSlide              : sl;        -- Output
      rxPhaseAlignmentDone : sl;        --Output
   end record RegType;

   constant REG_RESET_C : RegType :=
      (state                => SEARCH_S,
       last                 => (others => '0'),
       slideCount           => (others => '0'),
       slideWaitCounter     => (others => '0'),
       rxReset              => '0',
       rxSlide              => '0',
       rxPhaseAlignmentDone => '0');

   signal r, rin : RegType := REG_RESET_C;

   signal rxRunPhAlignmentSync : sl;
   
begin

   -- Must use async resets since rxUsrClk can drop out
   RstSync_1 : entity work.RstSync
      generic map (
         TPD_G          => TPD_G,
         IN_POLARITY_G  => '0',
         OUT_POLARITY_G => '0')
      port map (
         clk      => rxUsrClk,
         asyncRst => rxRunPhAlignment,
         syncRst  => rxRunPhAlignmentSync);


   comb : process (r, rxData) is
      variable v : RegType;
   begin
      v := r;

      v.rxSlide              := '0';
      v.rxPhaseAlignmentDone := '0';

      v.last := rxData & r.last(WORD_SIZE_G*2-1 downto WORD_SIZE_G);  -- Save last word

      case r.state is
         when SEARCH_S =>
            for i in 0 to WORD_SIZE_G - 1 loop
               -- Look for pos or neg comma
               if (std_match(r.last((i+WORD_SIZE_G-1) downto i), COMMA_0_G) or
                   std_match(r.last((i+WORD_SIZE_G-1) downto i), COMMA_1_G) or
                   std_match(r.last((i+WORD_SIZE_G-1) downto i), COMMA_2_G) or
                   std_match(r.last((i+WORD_SIZE_G-1) downto i), COMMA_3_G)) then
                  if (i = 0) then
                     v.state := ALIGNED_S;
                  elsif (i mod 2 = 0) then
                     -- Even number of slides needed
                     -- slideCount set to number of slides needed - 1
                     v.slideCount := to_unsigned(i-1, bitSize(WORD_SIZE_G));
                     v.state      := SLIDE_S;
                  else
                     -- Reset the rx and hope for a new lock requiring an even number of slides
                     v.state := RESET_S;
                  end if;
               end if;
            end loop;

         when RESET_S =>
            -- Async reset will eventually get everything back to SEARCH_S state
            v.rxReset := '1';
            
         when SLIDE_S =>
            v.rxSlide := '1';
            v.state   := SLIDE_WAIT_S;

         when SLIDE_WAIT_S =>
            -- Wait SLIDE_WAIT_C clocks between each slide
            v.slideWaitCounter := r.slideWaitCounter + 1;
            if (uAnd(slv(r.slideWaitCounter)) = '1') then
               if (r.slideCount = 0) then
                  v.state := SEARCH_S;  -- Double check that the slides worked
               else
                  v.slideCount := r.slideCount - 1;
                  v.state      := SLIDE_S;
               end if;
            end if;

         when ALIGNED_S =>
            v.rxPhaseAlignmentDone := '1';
            -- Gtx7RxRst module will reset this module back to SEARCH_S if alignment is lost
            
      end case;

      rin <= v;

      -- Outputs
      rxReset              <= r.rxReset;
      rxSlide              <= r.rxSlide;
      rxPhaseAlignmentDone <= r.rxPhaseAlignmentDone;
   end process comb;

   seq : process (rxUsrClk, rxRunPhAlignmentSync) is
   begin
      if (rising_edge(rxUsrClk)) then
         r <= rin after TPD_G;
      end if;
      if (rxRunPhAlignmentSync = '0') then
         r <= REG_RESET_C after TPD_G;
      end if;
   end process;
   
end architecture rtl;
