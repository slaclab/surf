-------------------------------------------------------------------------------
-- Title      : 
-------------------------------------------------------------------------------
-- File       : i2cRegMaster.vhd
-- Author     : Benjamin Reese  <bareese@slac.stanford.edu>
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2013-01-22
-- Last update: 2013-02-04
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description:
--   PRESCALE_G = (clk_freq / (5 * i2c_freq)) - 1
--   FILTER_G = (min_pulse_time / clk_period) + 1
-------------------------------------------------------------------------------
-- Copyright (c) 2013 SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.StdRtlPkg.all;
use work.i2cPkg.all;

entity i2cRegMaster is
  
  generic (
    TPD_G                : time                      := 1 ns;
    OUTPUT_EN_POLARITY_G : integer range 0 to 1      := 0;
    FILTER_G             : integer range 2 to 512    := 8;
    PRESCALE_G           : integer range 0 to 655535 := 62);
  port (
    clk    : in  sl;
    rst    : in  sl;
    regIn  : in  i2cRegMasterInType;
    regOut : out i2cRegMasterOutType;
    i2ci   : in  i2c_in_type;
    i2co   : out i2c_out_type);

end entity i2cRegMaster;

architecture rtl of i2cRegMaster is

  type StateType is (WAIT_REQ_S, ADDR_S, WRITE_S, READ_TXN_S, READ_S, REG_ACK_S);

  type RegType is record
    state       : StateType;
    byteCount   : unsigned(1 downto 0);
    regOut      : i2cRegMasterOutType;
    i2cMasterIn : i2cMasterInType;
  end record RegType;

  signal r, rin       : RegType;
  signal i2cMasterIn  : i2cMasterInType;
  signal i2cMasterOut : i2cMasterOutType;

  function getIndex (
    endianness : sl;
    byteCount  : unsigned;
    totalBytes : unsigned)
    return integer is
  begin
    if (endianness = '0') then
      -- little endian
      return to_integer(byteCount)*8;
    else
      -- big endian
      return (to_integer(totalBytes)-to_integer(byteCount))*8;
    end if;
  end function getIndex;

begin

  i2cMaster_1 : entity work.i2cMaster
    generic map (
      TPD_G                => TPD_G,
      OUTPUT_EN_POLARITY_G => OUTPUT_EN_POLARITY_G,
      FILTER_G             => FILTER_G,
      DYNAMIC_FILTER_G     => 0)
    port map (
      clk          => clk,
      rst          => rst,
      i2cMasterIn  => i2cMasterIn,
      i2cMasterOut => i2cMasterOut,
      i2ci         => i2ci,
      i2co         => i2co);

  comb : process (regIn, i2cMasterOut, r, rst) is
    variable v            : RegType;
    variable addrIndexVar : integer;
    variable dataIndexVar : integer;
  begin
    v := r;

    addrIndexVar := getIndex(regIn.endianness, r.byteCount, unsigned(regIn.regAddrSize));
    dataIndexVar := getIndex(regIn.endianness, r.byteCount, unsigned(regIn.regDataSize));

    v.regOut.regAck  := '0';
    v.regOut.regFail := '0';

    v.i2cMasterIn.rdAck := '0';

    case r.state is
      when WAIT_REQ_S =>
        v.byteCount := (others => '0');
        if (regIn.regReq = '1') then
          v.i2cMasterIn.txnReq := '1';
          v.i2cMasterIn.op     := '1';          -- Write address bytes       
          v.i2cMasterIn.stop   := regIn.regOp;  -- no i2c stop after addr when reg read
          v.state              := ADDR_S;
        end if;
        
      when ADDR_S =>
        -- When a new register access request is seen,
        -- Write the register address out on the bus first
        -- One byte at a time, order determined by endianness input
        v.i2cMasterIn.wrData  := regIn.regAddr(addrIndexVar+7 downto addrIndexVar);
        v.i2cMasterIn.wrValid := '1';
        -- Must drop txnReq as last byte is sent if reading
        v.i2cMasterIn.txnReq  := not toSl(slv(r.byteCount) = regIn.regAddrSize and regIn.regOp = '0');

        if (i2cMasterOut.wrAck = '1') then
          v.byteCount           := r.byteCount + 1;
          v.i2cMasterIn.wrValid := '0';
          if (slv(r.byteCount) = regIn.regAddrSize) then
            -- Done sending addr
            v.byteCount := (others => '0');
            if (regIn.regOp = '1') then
              v.state := WRITE_S;
            else
              v.state := READ_TXN_S;
            end if;
          end if;
        end if;

      when WRITE_S =>
        -- Txn started in WAIT_REQ_S still active
        -- Put wrData on the bus one byte at a time
        v.i2cMasterIn.wrData  := regIn.regWrData(dataIndexVar+7 downto dataIndexVar);
        v.i2cMasterIn.wrValid := '1';
        v.i2cMasterIn.txnReq  := not toSl(slv(r.byteCount) = regIn.regDataSize);
        v.i2cMasterIn.stop    := '1';                     -- Send stop when done writing all bytes
        if (i2cMasterOut.wrAck = '1') then
          v.byteCount           := r.byteCount + 1;
          v.i2cMasterIn.wrValid := '0';
          if (slv(r.byteCount) = regIn.regDataSize) then  -- could use rxnReq = 0
            v.state := REG_ACK_S;
          end if;
        end if;
        

      when READ_TXN_S =>
        -- Start new txn to read data bytes
        v.i2cMasterIn.txnReq := '1';
        v.i2cMasterIn.op     := '0';
        v.i2cMasterIn.stop   := '1';    -- i2c stop after all bytes are read
        v.state              := READ_S;

      when READ_S =>
        -- Drop txnReq on last byte
        v.i2cMasterIn.txnReq := not toSl(slv(r.byteCount) = regIn.regDataSize);
        -- Read data bytes as they arrive
        if (i2cMasterOut.rdValid = '1' and r.i2cMasterIn.rdAck = '0') then
          v.byteCount                                            := r.byteCount + 1;
          v.regOut.regRdData(dataIndexVar+7 downto dataIndexVar) := i2cMasterOut.rdData;
          v.i2cMasterIn.rdAck                                    := '1';
          if (slv(r.byteCount) = regIn.regDataSize) then
            -- Done
            v.state := REG_ACK_S;
          end if;
        end if;

      when REG_ACK_S =>
        -- Req done. Ack the req.
        -- Might have failed so hold regFail (would be set to 0 otherwise).
        v.regOut.regAck  := '1';
        v.regOut.regFail := r.regOut.regFail;
        if (regIn.regReq = '0') then
--          v.regOut.regAck := '0'; Might want this back. 
          v.state := WAIT_REQ_S;
        end if;

    end case;

    -- Always check for errors an cancel the txn if they happen
    if (i2cMasterOut.txnError = '1' and i2cMasterOut.rdValid = '1') then
      v.regOut.regFail     := '1';
      v.regOut.regFailCode := i2cMasterOut.rdData;
      v.i2cMasterIn.txnReq := '0';
      v.i2cMasterIn.rdAck  := '1';
      v.state              := REG_ACK_S;
    end if;

    ------------------------------------------------------------------------------------------------
    -- Synchronous Reset
    ------------------------------------------------------------------------------------------------
    if (rst = '1') then
      v.state     := WAIT_REQ_S;
      v.byteCount := (others => '0');

      v.regOut.regAck      := '0';
      v.regOut.regFail     := '0';
      v.regOut.regFailCode := (others => '0');
      v.regOut.regRdData   := (others => '0');

      v.i2cMasterIn.txnReq  := '0';
      v.i2cMasterIn.stop    := '0';
      v.i2cMasterIn.op      := '0';
      v.i2cMasterIn.wrValid := '0';
      v.i2cMasterIn.wrData  := (others => '0');
      v.i2cMasterIn.rdAck   := '0';
    end if;

    ------------------------------------------------------------------------------------------------
    -- Signal Assignments
    ------------------------------------------------------------------------------------------------
    -- Update registers
    rin <= v;

    -- Internal signals
    i2cMasterIn.enable   <= '1';
    i2cMasterIn.prescale <= slv(to_unsigned(PRESCALE_G, 16));
    i2cMasterIn.filter   <= (others => '0');  -- Not using dynamic filtering
    i2cMasterIn.addr     <= regIn.i2cAddr;
    i2cMasterIn.tenbit   <= regIn.tenbit;
    i2cMasterIn.txnReq   <= r.i2cMasterIn.txnReq;
    i2cMasterIn.stop     <= r.i2cMasterIn.stop;
    i2cMasterIn.op       <= r.i2cMasterIn.op;
    i2cMasterIn.wrValid  <= r.i2cMasterIn.wrValid;
    i2cMasterIn.wrData   <= r.i2cMasterIn.wrData;
    i2cMasterIn.rdAck    <= r.i2cMasterIn.rdAck;

    -- Outputs
    regOut <= r.regOut;
    
  end process comb;

  seq : process (clk) is
  begin
    if (rising_edge(clk)) then
      r <= rin after TPD_G;
    end if;
  end process seq;



end architecture rtl;
