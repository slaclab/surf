`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BsLKlGOMdeY5RBZ/8SZP7TZdMKY2GAjeE9r9yQWrtub8CY//d3+2El7z6jFM5yUZL1yGBgJmq8iX
IVH2qn9akg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dWLTiJgtPay8aGdTWGCZ4wBl/hZZBypc7MHe+FGG94Lv06D3dXjlWROxt+QTzZJqZkMAnskTwsMb
N3pU1JlMqlZDQS36Ox6uoB32VLDNtxE2CkaGIa0sFUpH+Lm6kCDBibYqC4QhLcfK4SOFjPOXfrU+
AAHgt77b+zoaGcqTEPw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OecO57YEu8tguvMHHYbBeQ68S9/ek3Y7gGcapIzzStiDMztG0bWCdKeaWalentqVLbUu73tzJmfe
751MxmwZb1rwf9lc4fKkhXV+Gm+HFuMITtJjJcoB8pKjdvA+HEMcufPjPXJDIaoqcuiAnm4Y9Ev3
0SczOozgAXlrm0afUddTt3rE5S/ue/WE4iymSfCCcsw4r8JJTd4f9rLV+swW27rCacWJt8q5YV7V
Vu9U607PsYnOMJLn1h52izf2OII7Yrs8/qY20glNNOmUzspqOLLSpTfjhMwzCUhxr4Xzyok9AmGK
2HodxXwvDM8a5LYjzxVo6YAAat36hnESEtVn5g==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t0cDrXZR5NuTKopWPL1o2DxK71KtsmYiCkpGYbnqBd0K0qa9tL37gfDEmKvrT5rAsqzPk7ozsR1z
Ytc4X+TipbKlpStJwkPQVXHJmORdcef2nxPUwhcUhixG0EMWb0tX8CyXvBFVJfEoylhTsj5qqIJe
bKtHnTNp0aXMNzFZmuPctg9PhQlTMJlS6Pk53XEqohyeOex+Gw2CPjW8C4Is9LBz5Tjiu8trFfLn
+8/rnMCxZ9Y4xmOi0JS+cUM2s1apHT8ezIi99NeQMpD9SgwRE0pZulRYDnJteXfmH3FQKsHrSCgR
IkV1ymUBGLjeNIf2V1rTYjTDs7sPm69rwrOIqQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u35MNEl1hY6Ryf3hxrvZPOEd/zo6q9y7p976xJsrcdiq7Tz54PZQsqbcJYkBSfiV3DtZu42g46p2
23eIrPhoh+qSBRtHie9eIlZEE8JPYeBCFHxFYGOmQ6L8dJoZ1JFakQgzV1qQR91M5X0WkfncTuC/
t1qCdMr6/osCLNxViIYuULwrnC7urOK3OslystNsnn3tmurINqnlHCisVzBdx8X7RYN56qG5DGBn
ohZLdtJpxYUMqfsqCH3pUlYQp2sCgyniMLRV9y+Ypw/f+/fLDxwN8KiksMcNQWpZPS08j1Qf7kTI
BJn+4ha4PNDhnFoG1AiFsCdfQUmgCqxyaAQvow==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KxSzBCWckkn+5nlj+daDkPkET/ouwdClQArAGA2Q551Bc3q9RO5rg7UtGyqdXCMoOgEfbjD42+Dd
IpiFo34SqLxPuPDtxW3YZmjaJVuhVq5O0AR3tyNqvEyaelNU46ct6nCvSzWwQo+O/LMzAgAsC5+y
0hAQuNeYzHUVoiqkjXc=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XTnHsfp8ieKcuCeXmN7ZP4tmNRxmuGMFl+7jFgaumtMmikSewqrvtKtmi6t7irPx+Sk40+Yr+u8G
l/iH2+7PmTp6wuIMb3GEZMirZWzkjlkC8nBEi1zFAdT/bq494xfoT5XzagYfkXH04OTfjdUa39Nu
iZcQZBfzGlwKk/oyxN8yjr5pj39843/F+vKU3mpaCrWOIGBphTUCF/LISYWix9VYfJB0LD40kK7Z
/DyJCg19VyXaSp3SLGN77dcKAX/sy+kirxFn6fJ1BYz4byJW8BjKwK86fWXFRlhnidQMErq2xfmD
H3nSlYP7ng//oGWNN5kFD2qT8JpNf3R+yCkrjA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 792016)
`protect data_block
XR5qC+/4bNXsAfLHtx9fWCsaGLwmMJyWUPFYPFoluK8Yuy2quoXG4mBVOgAltsn43BjnyXAJTpLn
ml7TJ830cPohoaVidc+r2iQz+FQCIvZTKtknrfWhZ+BLbjtJUl9Jh36ZpHfjKbNIB2sijKoRu5KF
eVDbuGPcp8P0qx5bP6V+jTfq90p2et0gqZ5UYe4BOHfoTr0lPyyVRs2HY4gGuAaa5zdkBVpJNqmY
vxEcsepHoAKYtbQnvlKvbqDkpQWJfOp2h7qjYVflJJsHuS1XIRneiwBNq8Jm4HX2PSaJPM3+t1v7
xHY5iQ9X9HH/FIWpIqKjO1NNVGHVJErgKueRBGPU9+ja02TCGOr5WcRdiCil9Uwd1E6H8lN7T8kU
m7AURdycldOl+1gFMcQ+gMwb0OrRVSmWwCpA+xWKlDYieVxhEbDmGaKeQnOg00BdjiIdLkREnlt3
bUVnCkzUicuURbUQ6uoaRrsu0hhNk67heVHxIdBZ/HrpcqUBK5XR/Yng5XWd8ZG+b64OqAHZzAIj
LXuu2mYJ5kMpspXzid095BV35+x0Q9R0KjMHKvVueZ63vOsQesKhTyKbZxnz+995bUbH8ELnApK0
ChnpG6LNuYoeHyoSxpg3R1j4x4tM6hZ7POkJR8kCJuzaHgg1ykPOwiNTemZLmM+nF49P3UOW5jIF
65WhW6EqkoChxuafqynPwAauYA4qrnY4F41O6gi5cexvflH/TW7TOn7yul4eZE1qa/P4I5hAqaOu
p7SXAonS93Lr1EYAXIjFbFR9mXMgM3y2R55qiTtyJASqVpkNZJKuOkRk2GLjtzioz6Mhj8q6Phi1
CCvUHI8YdaFtf4aeGO0/W9VgOAVmrnFtblRoT6/j72OAkWbJEyNAYGpzhco9Bs9PfDjzTWkr3T6p
4LdCl0/j4H6umPru+y8rdoTlqh8m1NuIVuel2RONRz4lWAN484bl6Hg9+i0W+mhmid1u4cddWt46
NwcTXYew2zV1bDZjiVZG2d7W61oj3lvw0l5L7K+4I84n3vzmOGcA0pDMmdQAawWhxaIOJuTNhBR+
U2J1jejmUX3Oe+bezc71NLVMiBr8Q9pu2huqLqQKZEGrmH/O2ZunZZJv6fsEg/JejYUlnaNEjPSn
/J4hzG1FiKh1UxSdENEKXGryfKv0ktUcaaqtsEq2V2F4wzV2aR7svWVQTOsai7LPLScmRwqtDK6X
JURefSPlcdj1CuaYTa9L5YUv4MHS3cWYT1t3Vv4+fHqOo4md9SK++pX8OAVOglSfgQVrYInCUtw+
UEdAp2sAIP0ShNWCLm+FJOOzA9gC/RdbuxJ13hZysajBs3TNuvZdZJxQVWjgSK283gzWEKSTtbGI
OgflK4LuAzVDhJcUmFbY2vHBWwbUpLN0c5/Tyk63BXiqHQnND4fN1re4lkdlmdMv95UHzTOF3hjO
lB1BpIL7HddQsyZQxc4a6WTvFVH49JRBdgaEET1/AJZtwJaaVJ9UkVGUiC5W98rNTkKlHGkY1Cev
Y0yFNB+dmCNP/+coAnX/Nw4fFSQkvlktTXa9VWa5oDse7u9ryOxiAyIti5556t3ZgsFR/N2WVzu7
qT30mZhg+FEXIgUGkfWW5UclZwbPdXqN2/LM/f8vKVqQPIwb2R9if/3hEKAHTN/PUL0CHfM4r6HQ
CueQvf2v71dVqe6rfmEHP1M4vNn1uzJSLYp9AmIArJvyfuyevdMz3BQKZ6IVJKJ5f/tuknBUIIO9
nrsufhrO1y0BKPs2g4A5LUR9GKc41M8f6lWJvFQTWL9oPe1bu+v3/lRDAc2l4/aAZ3u9KJg223D2
xcraGeIAlWehsEPGiAMGIKOqyXlc3D/PdFaCHMNesz+SWhftEZAmxf0Yrerc4auJvvVCcXCKomUS
OHtTyEkVZw9nxWnxVLvUtkkK+KmK9v+wfo36kNw8lZgPteN9fH60zpfgEQMnhjwayFbZFS5Sp3Ec
K+eCuPNYWlEC9zdH8ChhqFv3oTWuFExSwOs9jHUXBO1lR/GrnvQ8pV5QoLdOZ1veWl+HykrwU8Ce
uhHogP4ir8fVrerdg9N419Gj7ik6q78Xz/JSTVqMmjModC4L5Byxt/ekKWei/5fmzNR2mFBpweUm
WSqwIpfh86A0vYnM+HAopbxbtjmSLGIzwF4vXK7S7kN/FfX2HqS5FwCXv/YPdijZYMAnKjYnkkt7
hOkoILSluqrxpd+OlHjL3Ozy41CqcOoX2Ms2VIELqT227ol4jlO+GpAI2GRLfJ0tbURFo5ikxWTg
UMot9binJEpxsuxneGumql02FODLGjRijlpkGH0CUYJ+yzWwaH4sXWkQzEO5kP5Lhp9oF2oQTG/2
wSPtMCzs0/LwEZthz093SxJoCjCobjUAPQZyGZoZPlsHh8icDlUUWFZ4cFW85wvgLfx88Vmdli+M
pl2kzd1uMWKuvLE5WNt9/GbTeNJ98cWkJcc1+OBX3azgJZMN8mGjO6F/0qozMp5c9v+VMzSXsVfo
BhRnLr51i9T+LqRylqmmOuMjR0FNnMGPyA5ly4vL3PqUcfORDNvLwWsF7TaoFg1r7WA/y2z2gABp
0LjnkptgrI9ArGx8JkriH5zHZnY47HIVcSgyMET3y9MAI1ThYvYFZ7t/uHALR5J3JKtM7/wIfhJm
I1aEr/Fhe6L5DvF8dg3U9RAqewNlViXmzy9M0yD0mP7lbJWN0IZhY9dV6SDKdMlxdEHtbDKevXVn
Mc2xZelZ+jLBrDYsqMHMtsk/kjFFU9W+jTgAtPpHXO1C4RcoD5ws8Fxai7XNaprvGs8CVhWR4RWC
mvFoUJzipEZirLlOdTdO9djyKWzn+8o5lbqvEfaiVuydV0BOcourrXjqFzMOgjdCp0Uf9QQgbRJ2
9qnD79XMAplkTK/I2xkJoTmBKYhxzcx+hhqBwV9+AD7EYwWzX68kdcVHTbCwe8TXJQ5SBP47cbVU
gv5YALHXmZH5/OX4rSMbOtd0v3eLawctscrGcNeKuI9Evv2KzChZFtmL/EQICT6EpLFxK6mPvtaF
4ibaOFyuuC4LS6RyJYvGz+GR1OqU2eizx6cnvPO56jsNFx54/YZcEX60d5vboj+pFiDNNqIAzN0y
ER3ollMeHZYH5kyxoxlw30Dn2j/o+rfMAmC+CBUWzkA6ufG7Mllvr1cra8MHFAWmPcL8+blS9PbG
of94zkfTGhmZHCfBs42VMnS1b3ZOEfaLqTAoOofj9Bjj+729tKjMw3DNTDUlUAZoZlhslgiCq9eU
i6DSBE2F4Rp6NuJFKkFJr+rW73LeAfYKg2ysLS21Z682gy5Oasy6kGn1hG/Nb8TKvCEtVnAQB/nl
oOUfbB+iY5mlZ0btHWGto/fQZJlCSXfLtv44KJMKJbxccWeVVaOQnGwamoY/nPARfBl1WfsIpwK+
BJKRqYYBk0xx1zUOPtxB8a3Wt/B36yw1yDwryC+YzguPHTIFZbC9unPJd6hTFZHzzr/C+Vd1y01N
s0Cbi0fAA+xHT1QZvczj3iphigZ/iHlKID82n4s2JOPS6+envA0IOo+BjBlzaBwDmMux0vVEIe5A
QBsWqi3Je+VzniNbCfYDKXulpWHEzj8D2TrQy+QHsfVSdGl0xRUt2yF4nj9KrE75MdqfQ5cRUt7I
TpuwlqP9HkfinjTKXIwrfwyD11yZfL2VByUGxJG/hwakazZ9Z9NwB5GVmkZ3jdtPx2jOXcA7dAH+
2k5AtLVFsSd1B0dd1UOiYNa2V9st1BMsIFhLPC+Csd8Urn2nXaTgNT/pMrC+E+lN7xQTVjrumuSI
fFT1ERoy8lmLsFii64cyEJGq/tafs2CWlJ52gw2d5josCd8zKzdZb1azJw97TcczL+mh6LowKF+D
QRtKJKVWbR52h7chqOMzq1VdwLJ+2fDg+HZFLsiK615xMlU/Jejp5VVTBPfTSr8mkGr/0CQ+RvWv
8UPvHCF/A62l50u31y1Q+GOcKpkKXJDUixfIQO7AOwaB9t3WA4EjAga+PQMETF6VPrXQJeqBZieL
f/bfGSXLjwGq/umJLEpBYUeKWTFAIfSv/zJiA/vEFF96DvQf150Ip300oFLAHFtSJFOS24KqdP1f
tAFCO1Crrr2z3l6N5Yljtgg9+axsy9G6i9oWPjId9HparpHEcFPEFELWu+y5eBZQWXRjbZ6TtfX0
7BH2Gc8x8KRro1W7Df//5eMlYw51Yz5879Kk6im2QwSga+qJ5ucW9ncKzRxxG5VF90J71GJo4mXN
zZwlXEcvQxzQKYE4katInVCWpZXH+y9HWDrVlZy88hUlfzZvaJsvD7IfjJbANWDClEAlgbVGmPu1
ieIUxcTdP30zuQFI4+9LjcKJGS1Dwd2f194GEH0ciQhLW0PDhXaAyngf4daypL5J3YRhiu8Ohbvz
X1/+l7epPz+g2YaxFCVyobLncyEmo7NAad2M/brIi1R3XucmDo15DE/9v8fEGg+IJkYaXH9QNPGU
LD47feZiQNnbyCUgXaK1Y526CrNfDAhEUj0AhsLA8z+RsDfEQrflVljFQjE9PpKJmq0vC/7NHAvm
v7DZVyM8I6KuyG+Svj622LULgfP1DPSjX8xPptVmW+qYO5yX2rK7hvtgH48CPusieD1M8ATGbQpK
DqKGtf1hF3wmnS4oVxeIkD72MKdgZd5oU3KDdzeWRc/KWwtoN2lYP290clphu2HumF/qnNoFNkhZ
SueDFkl3NWz3gOadfIcb3D6aMYIVf4uAUqmVtAGfdXeiFoDN2VdfCRCNYJU/xoJrQM20xNlXRTay
S1Ah5PniqzLXORicpiTLT5itJQcI1w5BMKPj1cxPfRCiY7VvguXD9DaNzTpMum2elgD0vHNRMzau
8789Eh4dJoe+pN9BCWmv9yF5q+S9JZHJb2Edni2KkhY39ETkEHl9I6eu48oNUGqTCJe2xPfFan0s
3d7cAUxF9PNZUqmcFEC1UBOIVUPRBdhDISBw5GEbU16/qZHG5BPGOIIwcKT7eIj7XwapiN4p0YdY
ivSKwojHQMMixEJA6QUaD9XKyutisYswdWVktXWjXWRmoMqwdjRWrWRUXltMqBuJL8h484Ce6QOf
j114GcChF3WySVfU/Z5vln50YAc3AkdBlWA+PjyoDOoJU+27CBciH5kpgNg58egO/UeGHbDEEIDb
y5UtBEUczAWgQT3j3X0DiwNKHVETtUGq/FrgCWa3FUZwio3TWrD35Wz0kBhbD27rSLqGh2Xc1e2u
seZVIl/H46hxW0u5uvpuvvQqLDK41e84yb4b1kBiLciC/34MKYvkTIO29asJMN4kaiGwXB/H/Rbe
rzxkQC+bWrz0AugLIuyhXQGIstr/9B7DoJD99AdVjUuotPW8l1z/6eP9Aywkct6a+33h2KgAQUlW
Qth+8LvaBco546N8Nchj9sH//PyhRaN6uNjbnFpqJ5qUgSmr2wbd0shEOsg8ujikzB6+kI1iLHuJ
pEzzKaEqAI9705YN7PqZ06Ol2nYakW/XXkMF4ZGxRgcCVeO6WMH7q+Qoxm7ViPczKlpldexWrwR5
jeDLBReSz+qhotkPWb6eWWHNsrIFFFEEkumkjbfhAH/VrZzTwGetpT453lgxwidj2iPJKqFx7Dun
v55j3KJ0//mpPszCrCIyipRpJt4wvntZB5euaE9TLXpVx4n4/4I8EguPwN5Tv+nMeeuqPOM2JbYv
FOAJ8jf8NqjOCsT2gz3AzqTOJ0vJbwhPmqQy4zjd0Tlo4+tAcD1SzqcdVcVk7ANEaicmgqrUguzY
PigHvIKTTgkJJZNo1G/TdPNCiwBFdG1jFDiQ6Jz3aLW90ANNz94YPQcukKyAadL1p0GVa10YMZkl
O4O/NVI1MokzAIZwwB+zMKtkemGZCiGYph4FcvBpzR4FxhR9I3W1RCzG13qh5l4KB/MQsxf8pbN1
XlaUWNvm+Hdar4zWNOmckkPyMr8KhzgawoUbWUFbottkGznb4N34edCJ1LUADuUtBQgogjKLkuLo
jweiHBHc9XesxE9hGyvCygsvX7yB7X+mceF1ZhXhOkko6I9A+xQeByPQ9/LQa8/VdPXEJzg2NBvL
4fQPf7WsHSNpv+1dC91r7as4tSzqOPWihcvUymAK2RFeT9Uuyo4n/zzybygIXpwyMg5bvWhkjiWf
YtF4KOC+Ivt4uivcC7XmE077QzyV506RsHsC/DsderXGhVE6zmTG9hgOJkF8Yz3xXCLzdqtlw3NV
8U7yWAH1qCLhi97Bms64Jk2drYHJ2eUEOdMY7FJD6t95UQdKqBu9HUeM8Kh15hNIJmeaDTVTfz94
G3q0il2LdcNAWKig7Q5H81donkcm6SSme/xxsxZQINqSBuje1ApUdtWapvzAq877ozz6kOQTNT19
8sBJWwEnvetW9xLDDJ23ZF/C2u6MspKGtFkmOWPeCjwhum4F1gaqFsvsoXVLaq76HyKMSyPBUT2I
0Y/VMQTU2bFFjoIziHD3bjtVORlFtte2ENwBdOxXXSP9UNCiXVxzpDFLJnI5iqsiBiDPAMndJ75C
rTWyi34FPqrpYmxKTp6hyBAuz+NCqm0auqDMEpE6gVRIMhRH6sKzhJDYuPyGL7drgNIIIgpyI0Nt
pYxmscnugocQlDHNGgKd+4rTSMrBcQyDbrFdsTCP/3NedDLun619nb3ehCn00joTrp1vIBcRV7qn
EEGawbozqQYeAJud3Su4hYyRt4md23M47/1VN9ADKxqsQ9+/nB/qcVbTL6LcvnRkdOpHBNK4gt7+
V1O/zy5aUw0M2BMx/xOeXso5GqQCCrszOiRiKJSZYXaEo/vjz9Y2WzMjTCfNx9OAMEG9VPCOpA6K
0gvlutQXYOD98dZrtIzRnwFyfTyxOUuvxKQUCkP9yfZH4ARMDlvIjvNM0Mwz+Xiw6E1HvOiTD6Tx
qk/jNaMkdQ15suJ9uqTmi43f7eqv4ugqVJSiTMJHiyby5MXFn/u7x6pHQoX/igFrWTGD73sDhNlM
8sc77QlaLiWy6tK01XFUWucCoLzdenrX1xYnHYG1MGBTWwgzKDIafaHiy+nmSQ8+Y/EH9zr+CmPA
E4N9BNfdu8mz39eoAy3JPcyeZlY+NddGrKNixLvBreQT0yXTXrXYjOADXDMBBBaQHQ8xgoXPeeMb
O6O7YHcrmpSb5YJfI37Mf5+3iiJpqA9z/ZRwx3z2+eXIEKz5JBFLD+e3t3vmg+8ynCjWR8AFY/ic
Y+lJ/9uY9Z1yd3vUrklH/36Kd7QwEq8y0kxQm3lNd0V3QdNGAHq7kZ6wRE0rqR0yDQl7Z11pFdtE
u55HJjUKWvS7E95PRunRrk94CAr+NzoeACjpYHObCVgfj519mneOpHJiR/RXVbvK5EpYahkvLqOh
yMzPF/Zpa3Xtmn476gSoH/VkWlj8YauPl8F3m0GaleHv7IeG+psr4zCYQq8sTpJD8RRsDK1F3Xdg
t9fBad0IjNmHNapup1kgtnR3WK5gNKbRT3hdIMNCkpgnq2HQy1jujCyqIdKm5Czho/QCrliBHP8X
5dXGeu/Bmqwl5Ltg5XjjgQYvgz5o4gy/1UejHGDE/p6xx0vKJr/HhIjsRDtLhWpLiWsu+b80MKZB
Lf4tsbJfwAk/8TSL8RH0qHTNU2lB1F+vLTj2zsoZAZstis0bfLa9NEhmjkA7gsdC8ylLuueJypkH
YNrPpddwfp1EwKyIsvMYvPewGTYhDpPOF4BfEm7xiWMJ+Uqz0JxK+FowYoOoW29HIt2NdISArQ13
AVuzwnrgg50Okt/g967o2lTFGeWMNS6i6V4vYQdNfQzg6RbHTeOasvv3WCJ4dY+2277ckZFp7120
pprG2BbzoiRO9tsA3Evr11qVR+4PuyS0wrXm0UJwdLspaHdnCIxavwB88kPa6bGv9g9o3etiyttb
sHRQwqx6zv/+6aYqcRyV3JPIY40o9N+8dpBF+O85+VXvrtBs6ZRpJ8mtki9fxwrBfnyNmn1OgktH
SRWXIkPJkENkmOIwMuxwf/wAToeb9KBm9Uuuy4CldMrIQ0lGzGkdd3CkQkRQ/P7MI2bijhF+L83s
KeQcfM3jgnxCL1Ebc4D4Y1XP4lxReRw/o41vQamCqY19mUzlSnvjSUE/u288DKrbEDweFl90ojr3
wA6VBcWB51AMbieUPFCeWgzhnQtBKbVv7F0D6WaSELXaZxEQ42HioBgSiQ/qWGbXSJdIRA3EGdPF
4ZIAe1SaPUyd/mvT4NIw6YoRcsPX9dPJUF7ZH3hCPIXOvNHVWewSvo8Y9myFeO7rdakicd1E5kth
2mfshqq3ZTwHhpn4te8PF/SujCnD/SYlnslzDTHL2R3V3/MbuW5LwpawA/a5Je8Q0MYFwNcpo7pU
SXHx9SuGyh+7GdUooVXi+LjjlT+4IpF/AqOxZfqdz+5hdvSURx2wktS+Nj7wbKGGaszhpNIuAoYo
nEwU8EM34+YtDl8B2gJBe28L0I3U845MvCm/eNgQgTQjnwkSjBcKWXR/hs+c3LynADe/vyx2kv0i
LXdEXO2s7b1DYyHE2iehzJ3go0F/mJ5CzPyo2CxpXOoyXbHzwQ+eqv+Gijjf6uixGfPWQZmXSi1Q
+lc9J4WbPXIFaXjP7ThgJBB5r0038OO+/w2+ZtLpFA0ATHrWIp/rAeGAeZuDQWwKqXU7j+YMxDEB
xw7hR9a60/Y9+4zkNmeNBT4Ht0XMH2sz1Wets0w9/huWRk8LKmIzCJQAvfQDlnUwz8J29zkvaefZ
su76HonMB46IKWG45h38zoDIBcEL70I+zEGEZK+ajY7P82m/gADTy+DjJbOjzZHUlX5DJ7l6nLnM
TULpnCMuw/OYzNAmtYyIwNGmxxnEWi9BVt+JcoNqc/BThAKrdUoQxN0fgZhq/9zjEam3JgrGZE8k
pks3y/YEJ/YSqntWGkPqTS1ingqNKvsme5mTDFxuPn/0yAnjQxb1roCs3AcfTAY+7FZtcIBpwBKm
orzyrmQz7TW9OXfj3504r0jTzNYtVjX5xKWyak5tHw4IrHKV+7fMkQf09NF0/NCUdRtGwkxRxMTN
QYYEJoaQpJmo3CYzvDYcqgXhpJ4fwDej5vXV5KM6EP5c54h0fSMcSxWXk0c4LCTrrAbbGsT08r6L
G4kwAOPKPvsOROmFfAyLNvWduLZcShWFXJhXv4alZ8M/8yy4cYzUtvR2pfaWgfzAl5MQpe5graAQ
PBsOIEQaSifDkU2WDh3kbi47pu+PndlK3BkaOG0WwCPQWUHlbkzgI34DxJY2/UZK8nlnaQlsRc+I
EZYdQB6/BK7cFXCf9e57048ZzfIPBlch+aeDy0mgXPLl69QrTXyiPF41IFP3RyO420EPBf1JJSX0
VX7wPhaUvB9hkDQd3JS7WSYiuu3dx/YWOO+Nqof2MURu8CZt+n/GVNrTg6icrBHwPO3r2xLl5tN7
Py9GhOSAMwPdhBx/UsjaaP72yNV5Dm40x/eAhRgtrMM0tB0ymCdo0JbQ5AzuoUr8sIGrptk8ypzc
qCNMQQYEsQgAAFbDQqHWymJcRYzHFOxrbRMsfBSzsVLY7qzMJNQv+CBX+eUuR+mtMxGoKOm3YPEu
1H2T/A3FuwCcR1Gwl/6LfFfHPrWax5lMBaoAApY/BP2hy9pZAuiUHcEuD1yDm9fzpDVrjXt/saxE
dB62VUjMW6xjGgzDixao5JX1j2lR9D8Iy46jgARdpyP/3qsZO/OMyExQd9sJBl55AxiPjoR5e8mV
P+ect0yNSZOc5rzOt6JGx1RETlWQrCParB3P6m5EYHclzLkVX4KLnSet4xKxwDYzWvtW77EeefHj
AlvLE5VJHLeSNRzzXwGh6dvPvQJiX6y9/hV6TJHGMmHNl5wwJxJQIiU23iRhHrjTNJy00GKeMt/u
R3gpbEuUpvWJ/emT89eW0ov35z9EPzU9VW494GcNKpN1qrYKpBnr88vG/XF++lfZWOHYLkfojNOw
VWbT98p3vzg0clj67zqEseOJEsxSxjMFXX0EVxO0ybBumWNWC8vZu+LegUU8yabml+9S6w2T3/Ga
B7yTA9unLEEh42/GlyW7/m5YzJMAUQl3WHWreFmfZQQBQBLUKn0/GaHnPthpjmsslCJhakGFKynS
XwvCiDOl3eSY2p7J798XjAwp2kOHkRvJm7iCByLpKzAWXwUKjFFlfc2A9AEnGa3SZfC/JW0LVqPJ
SG8bGjqNo2m7/fH6Kl9BB0XwmzSAy3qLyDoav41ThNeXEtbTM+ZqsHD6fKrmzOZRZOAc+HKNfCx2
aTztIjQySfmTrKRHz60CKCe5gT3bz7wFydSPhOfpDmtidJwWTZMgo6Ev6YzqvzAEESH4VaJsvzKj
+hrD2jtV7AbaTdP05yR4cVMyj2BuP8F9Dad2aoGgMS8yXSa9ReSNPSQBYMPOV5QK8fzqzjn27iJV
BpcTQ5i6GC6C7b2hXXyqfc3BMvZ2Zq6BG4fN6xYzzAyRZ0WlWQ0zgCKkK3J0j3BkUQXzQeGWLRcA
JLnkjPgHfO3rNnx1NH/LbyDX/0PJdgOv1n4QKnHNdL3kUYgLlWa4Cr7jVtutLUiJL+7i4aHscYP1
GQ0jWTWf95k8pL4kJrLFoVRKSHF+9LFo+9RY8W2v2L3O20TWZI7grmRTmvF3B+arSw9Jum03s+Dp
vJwoj3YXqGZAYvEa2vNwzvlhiN8bgoEG47k4xiHpC/PiQ5UGK0hFn1fGOIaxHgIqDM47zfCgcyON
Y42HD9zwfXT0flDTzxBs72Zbat+INOo/G/vRM61YVA/ZnAGZstJ9B7XCBpoksH1GBeQBr6mvdDeC
dd7ZbLwoayz+fOEwg3G3X04tuDIfEbYfnxPmKPlPmLUZp6Kg1nAjOU4GJEHyu3Ko1+cdGi3uJDY4
KVWbEJVpqA48SG3LRnA6wJlv5eCHd4ZxlUoa+bsi+FyBbo7XW8IKRsSmZjX2Z/hg6drJVLynjPBl
KF94YNr35bzy/qKzkwKdns2Mr2vM6pkUH0mPaaquQ+GPFXGmqGL6dwRu+x3Gg0/gr/yqeEUmvqqt
CYYYCz5flQloct6lOoawoxfAA/mdQvokCezE/XxjH10T8WSQEtEU5s9ZB0P7Omgy7J0EqvWyQQoh
xtNkg+Mt5V9UKFEXDWpvs0RFLkgHj7D7KoMKoUedf4zlGYvB+pUlr0PJi6R05+7KZsX5UbimNWya
KqzdDbhNM7JiTfEhW0p9Cu/uK2j0DnzHQNr2GNrxoF8oUGkSczzqRlgGdxjJVcHULK4fJDIdDpUN
vw/9dhb4uuWnKMA8xpXz5DliutEazVIBIrmZEzCHWn2Q4UqiNSetAZIRDSPcJxI9+Ne8zd3C6Wk0
ytdeMr9Yo3JmKYyg8BverHPlmBiS7/LsR+yYXzZP2AOtmdZ4KsqVgDRJL9tRunrBiB8su9VzEn0y
ybq1SErzK4eoRps8GCxuNxM63A/dwkl/nGmoqlfWepexiuGqa/OcfqXV+rOSMe43oOu3ZFUMR6GA
nB9XpqN0cBaW/Y/jGsPmXAjmyChEMghb0qbUiiLeXd9Tu7COHd4mhAB+3hnEGBBk6c+BEEjuRqY5
rf639lg2VF5C9Z0Imjaefa5bY1RjL9DfAXaKtadn3mhov0ZaW70R/ioxW8UrOvnOx2D52agmnzbm
ntMMhsXkc383iaiZwZUEqlJVsYGZbZCAtW62bqXAd58eVEk1xwAKJau+XdLdDIepz38q+rrsX1PV
1i8riidThMNpNdj9MQENnVCpwqyk1EE4SWsxTySA822SRJeMbh21caRGsSk9UUHvpy5V0Ea/ED/t
VhQBGT5+qTqUrcn0N5qpFs7yck7sdxT4hWglEXWEMrQSNmVfcA8qasvv9UbWBbopWlSsE2uj1AwY
S1yLBqT11CZqxPqcuelrNdM7S5WZMbzWp3AdZZQeKA4qneHxEhoA26F+iOE4yUenGl7oqUf/EP6K
yGEg8USO1vU2irymb/likXf0+/FJY6Y/NB9Mr4SFAJGtnlq19G8R+A1/m60bnsJjUaPvAiDTYS0P
ejfRKwCsoh98gx8hHJqj/kwtOB0wMVwuGj8barViWkRF9n696wgoHH+WS0rEQgWcFPs/UfJrn42E
cBLZlRTdAJhXre5CrO50+kUBQzyu+zfUcOnkOauRshgOyJJLlIg9etKJi7kKpPnL9kdMd5q3Gaxl
QdOjVQuQcQiwDuerhq8E4EAMmZEhxKD9cJjbtPQ/b+7D9dTEnEWxgYRm1msGbctnl5L7SOITcLg1
aJ/84KIQsx/83ud+fLtjQTMHndooshjYiZC2Ep5Bnae5sOro9refFaAC3YNJ5mOGyR0AlS/Nhvyx
gGAdSQYG6l4Jz3tCSRx0LLHrqMQBTaTig8ze3E66CwSHV5dND+5OXFOqpMc4Mp9fgRWYYeu3mj+W
YJaIudJc013nbYVxswWuIqjnf4xlAaNmnaPcZPBKjQIqN+tqAGYbYrGKVInmFpcX4IaoKS0SN88n
XMvVSrC8L3a1Mb+wIb1v/BnSFO7GP8D6hcbrHOPX9RUQpZdKme/3ADqkWDDZCYHqYImwBsDfDhJL
8S4sOtYWE57TEr6lxMAn/caxti2VDZOspSrHHXmExG4sEu/mS/+Kz61K9zKafTTkKO5Lx15kNqzM
+QU1C+GR6sH9ITR9AJ+VgRjfNhwrJoZXTW8IJlmwVhkEzlyQJE0h4Y4n2+8D/XusgSfaak7XI3dS
DMgird2EsJ6g3DC3b8v/qUhugPWdAUYFSmmK5YGlDY3ZWUfsoHefxfDsoR5kIntPEEpQehSPtpsv
9zL5KdQdYdCsiv0E8ssROBydkeRb8dX4XasiCYseNpTPqBT/qc4Wq8gFyONLMWZLvDMTSlG7wd6L
iCQHyILwZZ3yNm9cIIHA34CuvgnhDCjcVszqdJvkRu3xbt8DiYNB0rOO/1d9z1buff5JHJfOrSFx
a2+Ba8ULhKDjY2nTuNPUrsLmAOzVqAHTcBcxmRaIfYGJMNi0JfV82+fGURpXwOABWPDGCkKhZRlD
hTipkkbzAsxOxFDbL05AUqiEDMsEziOKTuUSYREaOtKyGOqFjEYFPIG4ZJDYIclTXeCztzZ/bX6T
gaaMU6bwLgksoQY9VJAy1ltEvfvIovABGekgDWiWOu6Ztmab0IjRb6/gnhbxXL1g3F1dHoZeMWiv
nsMd0aYvCVsKjTwQM2MF/X3nM8RhJBVYOMnQ1LD1OGTTbufKLQpSDRDlNkGXk28TMMDY8NaWtSNl
nmFHaQfaCwClS62mDXTwpVl63ey1uEmrSuoFWg0XJMg9ymg+GN5FYjWC9ffTJOQe/vUfidiVLgrQ
ftJD/Oom/ncgV/BXHXkHBP6duWIi9kPG9/77pfTCHE+7PmzWpijmKUiHP2IvCeg4UD42SClbTp2b
K+fBcSGjkSd5Gv84poTgAV3Qys4u2w1oooP51wB5Uri40GtYmeWYoDpvMHZsTf9UrCH529DYoFvg
0aTVvpVQ3xY3IMJBXwm/IACdiWoTubMLTBvsSjAnfWniC4x+Knc5PP3CCSdt4QPT4D/CJ9f/O3XB
gRCedH669dcOYT2GuAIlQ142A+5nTXo2bmQaU3C6AuS8mlyu4QlSNMemyLdAv4uVApXkAFUNy/d9
jJKo1E1BKsTAQXkJZzIF3LylDrLWpiRaHxtJcixbsVXMoP+BuLfIw9FneLO1+tBkPU+F/imqRK6r
Kwu8gV6pj0IXvbePebgwl4z7/kpTgIdmidxkU6g02WsLD7a36JWsNe+a5NgRjJzkYeJ/lbunL0cE
ZOYyPV55V4xLg2GtaxJLa/KAnFfHGqQOGpe3sHbBDcpdyzhwaV9JEvw6vggdzK/eKVJmoYBf9CcR
B3khuiih2fcQEQ3eY6oViVn7MA0WcfSC+mhuvuPsln/UIDyvYUYUFeRqL1fiSHfvtVQihkOrhDhy
YvSeSxOo9+TKR3DQu0n+NI+WJe+s+igITQm+aH8OvpXCBzXh2WPxxnwW8CIuZTVxMZlI+qUjeMMS
OOXDZvDzFWpviYOWfIiL8Q0zL8m9uom9r9rR4UpGzn+ghu/NPP0LvjSvjAqWdhard6mBSGaMeT/Y
v5PnvL1J/HPxaapoEc4kwRMWUZ3y2eYvK8x8Tbc8a4QHL4uKTiJUExnrBuWwFxfopuvO9N8VjOim
Qzdw28SSxgbhUAAkALs2O60Ilb+3tP5sfE2HlG7JaFPibPwHO8v/A1xoj9hVc4SdkcB6iaR/8VHR
iGF7Q9xBjHCKzVsERdvE1QXBHNQlpwkrwyKiG/qg7rW8yw5k3dhE6AZ+LlGX6in/Dpr9+25rtDYE
c/eZAl+wj4TdNDnjuKmyWd2sc3H0fMNXt+bCDFSd3sR0BWjMrNNg+n4PoOvEfFE37loZBkqoXQk9
1FSQFIhU1RsUHbRss7uappQgbhi3Vt/Do9nHobTkCTa/au1WZBeqNwN93UH5Kvy0fGKVzmJNNKmT
YhcSel7oWPFx/OSFz9NbnkHbEHpLRahMXDQBn+x0nq3D1MCvlyRTPQFcmMOkQh35mFaj6q4/MkXK
CC1e8m4Qxh58II70C7kAaOPsmpFsIHiOwQT6PmZtDCCQ2Z4yIcC4Ww3PwToVPD+5U5S1iP1+BZcd
W+ug1jadyNK+3CBr/9Sgt5xYNesvrdaj1M0bSXdztIUmH4YfrjBJV+jcxRfg185gH0grt7JRuxBy
ACo+x2XNSmXNbvigf5JXM5vDZL38VYvS0HOMVNKXOdJ0U7hNNg5mkxIOTGHFXdmuaNHrdOAgOTus
uGDI57I/aeQh9E9fEEzzHC8Oj0j8QiGzKNEX9rHCiSesk6kdyCe/qAuNkiZu48cTgqzARbaNDDh2
APQeyLz0gBJcnLA1qXhp15/Zri34qSDYet8IA0We28vyBKvaHlp4f/F18s6f0XHpB0ssvLkXRwhN
Cxda0HwYGtKP0ru6d1byKtWrc9TpSQsJn0OxIS1I+UuAuGXuz3N9ozpHdqF95CXAIWrJx8hZs9W9
eefDu17ePvs0uOxEgKO7lVJNA1UcMoRFBGo2tkFBoOyMJHDRdrGHDJkNf8WKdEmZ32X68myx3i/H
YGJHmw5bLtBfcgyHpic+m5I0K4eU7krRmEv7qsz0qC5qH9v5lhuwTuAZ3ByAdxvm2rJ8D3XqR+Ou
y37ewrnDjhKP4z4fMoBxWwGgUGoReVa9KCvsaGaO/jSi5TwISlzBd1tDdQE/u63jMBD62bKOBQKA
GaY9d22UEoJtxX40jFlCl18uXPd2ZAsh1wiFLm9kZ90bB2zZomL0nI80rLbDASIOEPshvdsA8zXZ
6rJvm/Indst6H898egTDN3URg3O1mPMwO/mP3nrcyB0aT73sRGpnKKQpGwQi09sADiuHF0RxT/Ah
gk+EWgnUO93SK6SjdKt3ImwKxEqkjA+i1cZWs1W6m0aMQBAk3C75rwMIjHgyHJI3qplTYgDdunpK
jS1y0OExtKwcb0D4BdH0+VqZKti8mgJ4afUIUk9GL+yT8dCLOkKerOXkJDymATJx4XmJKfILr+B+
FT8pX7/9izYSp0nu1fMyoLj2p575eOwoWc/geyTOjhzUxLrr7UW0Oht6edtw7/kdNdD4Iprx6L8g
MpDE01MsX/7MPcNFl7we9eRaNfUaLKg9WfMREcnjOyXzripyQCjFYXyZgAk7xNRgHVgpEwIl+d1U
Dhjz6AsJoCT83fFDxSvMALPM4GhDl0a+7hJwMlBTG+UJp5XHR2ZvgTC+4MU2HQYKfcgEexctje1C
N1fOHf4NeQ/2i1+F6sO+DzT2ukq/A8j2HlL7BqR+h1NWTwjsVmd0BUIQp3cvuCQEYxe2Ges90lrJ
4g7Xu5Yiir9zJnQuEvqt2V7w12DMmHHZudJldkm73XfNNG7ty8IpLoKOUt36x9W/RHar6Tim3QkP
BSORwHgnzQ0b/7RTUaHz2N4n1ARxsp8biHZYBc9Xq0cedcn7l9qwf65SytWtefaDD6h3ARaZ9H+x
oNnjx/BEjBACH0kREX+fUu2CxsAZ7jvOHexDgwUuWSuMNvFAq/1uqEBs/cCNGRidZezzIN8hFg+U
Wrc7oJV+nNwAXyXI+F7Xe2zT7ZCxAjxH/B2RK9WGVjme2dK6ViNQl9xXgoU457YDDt0PgPPUg2H4
uxtGRYdjtxM1EpTTIaGCC3ghHC0Va1rEZ8XW3KJLzEVMiI45lHz7LqUvrUA14HGLi1WgFdiatzlJ
Lo617U4OGUGkNOTlOSpmaPZqCzkgZf8PC+8BFpfnjh3qU6qZ/DnLi+vJ1rL27IyxN6u+aHhmisIf
ZzmkMdnIrYGD7kZAuQB0b0za68pEgvzq16UE1xr6udIuBSODeEYtGUL1nn6rknilSKUGGoAUEEx9
/T1IkVsg+W3EK0XQO7KYg+Ruvo5b7FVrIIL0/K4RqfvuwzTIMq6NSzyS0DVVv9txo0NtCkszVYO1
HD1PTzQs/wMgdu7GOdfawVuEDJBmRj56155mBJQI997R9rYIHrMqIjiIPn/J4hs+XFCaoLCq1Ozl
iwMQh/95k35zTvnCsuffigMWth8soJZx01gVp4KAKDNV+FyJFCNi6pH5su7duh0kjKS0h2q3QO8T
GYRxO+eT1heVJqMp35M94p4A7EAJRKRXylb9CwrU8o2Xfj08fmS/vX+akfgYQwJFtNs6CD5zBn4+
YqvJbNMB0flNosB4rhBXNzMT9rDmBHB3v0RUv5g5bcVdsj2j3UnzC2G5rXYlC75ANJQAhqh/Jh5K
iDpQSHlQIZzP9/Hrp6xPbgFefZLWQtfFJY6C4fztfzFXOte5vtz7KuoYEaXGuZF3ZeHF+Uu0kQ1T
82uXVeYyyeyChagAQrAUsr4xdnrgDB1Ok0VnnIonzZ4kmKYJBWWhNA3TEaU/ekJ9JbncYujBhGKm
a7EBtZrV8jbhDpnMNJuwgCtH9eu2Zgsz2Cn3oWFGHFUiXWtcLDt1Bo/c7n8h5VLUkXm6Ckx8qcTN
tzGaKafjFivWiXUpQbbcUITMPmq9hblV932rwdte2UFm8bp1mYnKJ+9H2S53siV72VxfrAewwH8r
JPVFMm4BYdjoA1UjAoDpwsEWHHbXBtwnGyIrNlwQzShcB6Pe8g4ZEvVhZRfDLNnStJKcn3ZrgM15
mXI7OThKWU/8DL+mP9onjxDMaMekLVUpah+i4mGBkGZP/RiytLZeN0rgdgP5V1qgJ0uUSM4o/Uiu
xdCMUYNjMiLKQEBTvlfyxlrQ/dzHzQXKXW/lD4ZSgX0NwEeKmePj1KnOn8as3jOhw7W/x2NILzZ6
mzOCa1CKxwLrw2Ee7cVpCsQTpaecZyEXNjJmyyYm5HyVHDqt0ydMyDPgbNe65Wsn3hYmUc4fCLve
vzdZFYkPka5mqL7r8394ei3MGrIkCkgnOWwRHPLWVivMbsisZO6zCcBHkJpbMM6XdFitebCzRvDb
K+bWDPQGdUV+By2E5ayGmCBWgPHHjSWZYlQ+YNk3CwWFBuRS6PxLtct4bkZr/l4llNlBiCgQDCTY
bbJoG3ILj4V6kXNNfJxjstB5XtSe4CjycFcHyZwydaDPS/gh6BlxmsdQ2SUxJWbb28CxMYx9QkTi
+tWPwEVBZbM0l8hqNi9LsqAXNqpPOxVEIGXucTmE/R6rcXmzlAvNJ/L3wYhSUAu1YmVvGoT02Mwa
J5hSCbokdtXcJp8PVSsmFHYrMPXWAWmYV0ANvEDoQSlpyCZzlZYnlKQk97uGQ/jNj0EbENDfi8ua
I9Mv9kTgMzGIP/EFRRmHyS+5G3PNMJEgg6+uLJBp5FGUYw5H4HmtW0/6sQvEGovX/5ydMMo7Wln+
cLs6JEm/tx6MUJRHnzUeEune3o73Yfkdp1m7KXIf0qVAjpVu9FF7zicNXFUUwvSbmeBWCPEEGbj1
SolH5NhUsojgy0/wxt8qK6E6XzF58lv+SxBiJegbRgdlZsWzVkCcHokARDAsTZGlAFhVUeAHCxNV
byJZsfNBxGjWLOjf+u0jdrH3D503NylmidvBAcJgGs8rcOlqm49WYSeg/lzW8jdfx1YyHfuf3qwC
4j2tI163h6GoYwvnZH4zbXw5j/0jh1TwvGKezumpRbU65t8emvV4yHVLT6etxxHm2foqMjJ0eGHr
3iSVGRe0NDCJynkiJmF8qyU2vJNkul3OIBj1X/4rugtusi3h5ZcgzeU04k351Lsow4wQ8fDtzBD6
q+jG30+04NCYIxi6UhL0QvgwnFo7T1H8MqX7PG2i5XToCMW+42pgbYFFgsE2xlzzbOgG4uIQKwgf
8SJO6gD/mRvknfvEgNoaHaQu9Tr1jNlmLaQU3rJ1C4Hgp4yXxOidwQvDUPi4MdCN0kiAF5gT41eh
2cSdWgEdDO73jqI0bIrZMu/LZQIKSSIU73dmsH11rt2q1Rj/ZFIRH8rvs7m6mQekZB1hP2I3mpmu
wybAYqLix+U3+R4luDU6E5G6mwCj+I9fm0PALeb/Kxuh5FQTylZssx4Bcpu9BWI46Caep6K+ZC28
HPKfpznMZ1RCzrD52Lnk8PXEsqZUucRbkSAQfQCCHgEkeObRkCmZw+h4g1Em97g1n3r255vlGoGm
uBbKyVkyOWvVE39pqNuFCJl96ACJcfc/wzIIBykS0c1EIKevumuH9lqxybxxA9lfriP8D2Ov5U4r
K9nsB8ES3nlEf9SW8giaa78+SC/EKaiBcULcsZMIs4cu+SuG7lIpBBaMLfUs1GqNpHUaI7mCFhpR
C50Gdn94WKijb6UHzibPIWdd6+V3vWopaJUoX8CTtHyB+S/AO4n7CdKyCBLF8DCtB30RA4+vPmiS
H7nOr+o4PHUizf63GP2/3op/DmEz7q+51b2dEszUpcNAqgoboRVrSPduen4M3QucPmhwR3if2KZX
fDtofWmWQM92kIQqBqn63uyTqtPM+JFAqkoeeZWGC32Sf1BYqAgGFwVR4TQh/cDFnPPF9bCU/NoN
uFOwg+8zAG5aBWLkEKkWZTQWOS5I1YD32SPJDfEsmP2sPZM8xoUqhooH0e/4KNgcnSYG2LYv0OT4
eLiPSEB3GZK6JIXibfqJBklCn8CcTonQGGJ1PQ0e7VIogkmjF89g7OoW8O14AJtv+MEHWGQIbjKx
RFuZ6tbxCC8Ea8XyoTnz2mBA3jImtzmFM4V1aAkeQbA6R3th0XrQmgPZztu3gNA4fNNJ3aBMQfUT
Eo/eh1xerLKXGE9JyC2zi6YuM7VXejB5N1wUOZCzhs/CTQj2NVfksJbkUZbK2s/82+RCgprKmgg5
NBMTOzFagqwZML5weA5SYM2acxtJR+zdBld10PzNGoXGEHYCy/conJRMWe5f5WznJ57qSHevmwOX
s/WHud6mrCfF7z4p+swnqME20o1+lLM1VoZ3BMKGIecIW+ufwmPdVqSaHRyRFK8bPtmeQb3fUhki
rYFKtlEhMBdN96MieomfHt2dCV6Od5SxcH6I3y3V2QdRPPslfDg4aNDp5cxpAT1O4c97Bgvb3WGc
11sYOOS6K1ZnMZl9d6eecbJ+cW+vADCCWLn3PvrKCBLW3LULu9CN9V6lojQNHECnl/JlqgCO2X2H
A/rsOQ0rnUhPzv7vJTF5nPFiMkoaMbSjBBpdBSi8JP42IcHbJD01HF6bHLCNDKLNcgdWM9xFi4zq
U9H4/Z60M31qnhi/eeF12H2Ye0me1CGMySyVrZ6fA++gDX88HtREwkbCGQKtk+iDynfrCa6WcDwN
atxCP2RKYpr7lzbQU5SKq8QrT/QGRpq9Vom5L9u498APgCJpjeU/aNTMhq00yJ1RfZ1v4E7ExLlO
bZ7o1UV6D5Jnf2prsg+TDDd8h/Xui4Ieq9OLCNMT54+EeToxW93hkbUm9XQg+Khm+vuUPPSylQgn
cOSoBo2RDjm0TbqogqlkmNyhfmIjhPn0IgPgryzSswEa8c25BSq8Sw6vThlbzCidOOrGX2Jjf17r
KMms6MzFrX4RKhYQnEwwy+cBxOAEPj5jH3f0AXpMaPOvZEG/+Wb0XQkYmg9qf3XvSqQV0dD7Qjo9
c/ogquTD90SETZiapXksL9DCHsyeK2C4kBOqu+EgmR/bbB1fP0H8XwV9XBX2qw+w8z+QwJEX86XM
ziW0jGffjoibDGu4dMAVwHsAi6Yt8Av89fwt0V7k6sMXazgmLy5FS6c2Q4JkzFdjvi8COXWWE4Nz
9E47y/DuRs/CdoCSPIqfbw+PT8NBY97QPzahDvoYxlynjIfjs7TkiI/wEedl72tXOKwfdu9Y/8eE
Y35Na4NSQWguGl/vOEqXw0CPdZ2gbbAxhM2UWnhCcRAMGpWNUy0lnDjGJboyQOL6AbvmJQbddQfs
ir4COFXevX3cvNPX0cLnvHCFmC7qA9Pk98EJvucGbjZghDzS409pC7JpHXFOY8CqbDVmjm4cWlS0
Tow6tYiKLj7G3phNfqX/XOu5wHCKUnaDtAE+NWJeUpjsir+ajUTTjBl2jMU5cVzAs1mlx6hgZENJ
pcIwUVRARsKWhdI0lNbUDGPCNfr/Y8Ae9iOZUITJEb6yRZAn11DbD14QLyol5RQyxLIx7K5X3+tr
MXckNCDuZPcpVAekn8cZpVAfoaVTGwjC36QDnbpamkrr0iFVDE2eezKGBlHroufH9Och5JtJ6Y7Y
dtQH3HGzCWoIB/Srws52i7eRfW64nG8mhTliK5F4HB3cTaRoqN2yUKPDJd69KRfh/c3Qa4vuLkNq
mEdhF3Qc4OpIT2xjMXbTYOe3C8lTDzjgN+inJiH08y8Ep6zxy86jV/pufXrB4zHdCDzCv+Y9wFY2
qenpXD8MNVkoOgHzvURUrHs5SHh0dYamfMOKU9zXc2+qlIB1pkwxHsbJRe8bifHQu7upIWAvr/sz
GY6A8U6JQq62EkN05Ot9V97uAvcHgAqiuTEwroV16YpAaj85avgFgRe9zsewsbK92bQ5tDv3Pho0
Vhha/l6SPz+iM6SU4Fg0+GOJY4HaulJZEZ27CdxQSxulzX4aPBoqxlSZpYZCf1tzOJpvL93M6KBk
d8US254yLG2YgjhPxViq7pEUbTnNtPsE+0xM2MTS2dchunpbVZf8/CV6QtB7LDSNwpAhccGyVRQX
RU9ZWBqO24qOGaPNEOa6fLIDJSEe7/ohB/m0MndLu6n3siUeSb231yxFjHijq0OlebfCdybiIHy4
o62UqjT7PInSyTh1Hf39qSKJ+WhCr//66u6qEZS1TwAICv6WPBGbl5HuDMTBeOynE7AoZ8aj8Son
IAcQCPf1EwKKDakwwW0qbJovE3FsuKm9A0B9ubpfFdxBFRZ03BLuQujuHgKr+ue2iMfUuqZIhkJK
F7we+9r6tCHNUCVaxPrtkhSaPYKIKSIQcSj8TkMzUs7ZggQPMQVlBqiMg/6TYfcO9UnVFkgXQe9e
UUxDnWLKyNVx03jhhbkZw+YTnkmA9VDOABPkHWlYq9nErBr2nHCKUf2XQvH1evHL6G6tUNFkSbL8
3ELEJNMriNPgA+UehseZPKXq5xA0gxw7TjYDcMSIo/bH2DY7xLiRzwBNSsSuQQSDKNK1tnM5zs7w
LVHUBXxLUeJQnq+CAT/aE2PL8Aay/5rA3sti7vH8KWqKSS/c7HITDA7nWrL1TIrlHwjBItoKHD1p
if9iCSORQjnxGw6xcjbUzgWG2TtdbHHJCPIk+H8akKXExYNlmIszXMGwtGAKYAv8iU4OlDFTWCbJ
1CLnylJ/9y3KVDzY4F6D+Q7KP9dKX9TMyTH4atk+Ywex0XYoX52uPp2iO24aDhdhMGng7AYoQ5g+
lYJfCSwWQ5edHr1QJ/t78+WNMj62jN4UvgPuS5/9/0qm0r1G91ZU5sTYYLB3MEWVBkHM0llo+rf4
X2AmXXRgbj1BZNXUqJhTS7Hz57YF3dQXokD9+GOsatSjgXj+4gSd7ukSlFbLvC5PQV5TfXzLVU4o
QLC3F3mV01ZkX7AHvjLsHNbLDKA3IxTQEjTakt4UD6FCE5tCzF+hJz/0ET5R4EccBoix5fW7KIl8
Qz4YYMSifgpDKyXsvS77dHa9WqvMDdStTzqHWJaw9sNYFamNAaTc0Xrm7hHcgyi5wj+GzVOj2Dct
D/gQUyUk5+8OEUk04VgTNkyUWPkYL0MXIJYXHbSRMcE3y7pzs1SEiNPgyoyULbj8G0G9RPzdPWjN
R7GbrJRz+zg+kCz5SdE0RUWJAAX1tlm+fgl7rPNzuGdwrZYDcWK2kkCgXLvbvVM7NQFWSviJmukG
/YKXLF2R++bhwmqgOINhef1Q/1yV3PHvOMG8an5TvN2G7/5nRlIRbTjc5IVnNjMinRLOkb71dosX
lDPBJHR827CIYsMANwgupirWONk+lYNzdLS36HM+eSM/o5YPuK2+Hk+8aoJRCGmU3cZrP50gdOwJ
VA8WeikwcpfMVVLZhVNOxLRdZ60GQ6TLMKA/548KY0w04rTBbSYNC9EzFVvJAv6j+p6kexhF/530
4Bee2w4YMNiR2ULw6MmzAK3MBvpvLdi0vQG3YZUw4l+siC3Y2ZRJkR8UeIGZf5ulzudosrtVYwds
papBFBwB1qsLFjH9ka4lC2q6ay6nAq2ZfmysmvP2JqzIskcYVJOshUwJ27NOOLmpzsqXFAxTpDrI
VIpukJw7ZGiujxlYubkxSPLfKb+fn5fVpM5E2NepJ+uyUHCg4KYpdZVE6xJFB9gNrBLHa0BrLGGN
nwD4/i5g4LiPEy9t9Ig7LDMafA1BXPZmYD1AE26gr6z9684UE/XoDyU6x7euoqsMjElAew5U6PHh
/vpRb2Cp9u/zLIAIjzYR6F7IbuNXXongvgItA4kLu9G5EIeFsKtyXlEVLEnn/k6/atavTck35hpS
c/alOPQY/wshZ1RQ+4om02hmSNF6FfxV4CFtwi1ZgIPXUK6d9/ZvZEWAoL+qHNQcA9I+A3I8H4Qt
xOl2siSSV4Xici+Cr8l80y+4PECpnvnFSN/a+FmKhKeetYJlFqTkS0ShvoiwYWqM5Yc4tRC4SEXO
qAPV8E+GWkTwidQGebtRnaFA2qqjdWQAN3iumsl9S/v6irrtE2AkkUU0XVenlgR9xcqE1tDHskMr
mxPRhDnb7DCs6JjASSlUsXybZ4HAvhY2WYsFFwUw5Onl2cMzuD+gxDgY0UGuYJAWZ2f0BAL6MJNF
SCT3OjFeCRFYjMaH3IBz87dlFU+txsvG30bV5ffksIS9kTL9nD1RdyaUDJjUQdzhmf204WQWpQFU
J2Bw9ZSNzNovs2n5CuRajI9YQn7stH5t80f2cbhBEmIQWQENQ+yCc1bMdZX6I5PE/yZSbgxtxUAA
sy4k+FR/RaQ2poWwGeskvDuvN+PowNRhHxbmsXv78dWASJEDNTNP0+uRdte9jxraXG3/IBizhr4H
FCGSV3d2WhKWj1OPJlaExGZzGwA76qGmOK2a/2N2+79eLNNbT34y03c9W5P3DDgm/28zHq0ubqZl
V2aQz9+tXUi17OpFRThpm900re3/ltk727fQdrGQvZH68ggVGGPbliFDtDdCUnya/9wojH1RWg21
YDXrKHNOgbEkYwLoJ3zHaCqFgkW5oKywhYYUnocUREfqxUglBPRd3NyZiw1SXJYem0fTyQk0zIs2
QbOxhSMVsx4x/sSPxINkZvq7Bctq14rH+ObcZUejVfFproywY98ThjYS5cLaJ9j/tU+0DC3Cm+8f
gC89W1SgERJ889ONvF4cLd+9BQ/g6+KOUVm8X4AiWbsosTpbXjYOEBDydiOlkuXoAZs57FoxHwKm
np4wcQMjihf8HVl7J/61l3jyXr0T6nkVU/ky0cnzS1NE6PT46TP/oXsFeInDmq/la+CqzkK1RKK4
PE/O/rtezqJouQag9vvunNYKlVeCIccJ7FAEZjP+aLzIEDaD2AUNCq5p9VFdAtlH/uxP0NoVM1Wm
hDQjzhyxTwTUG1QJSp6rrtZX9ujAgS7rhBmZ41iu02sg2VbarkOBPO7xFxE+05SOfCOjxMDBSUlA
bW2iLA5ntw+KxF+rGJicoBL2U+EuZaHeT+LJrZCFYGn2H+ZdQoCBixY4/eOMsdSYxUyV5NwBOCTX
/dpNwjeRXxhW6kxQh9ipFPfuHxQOCLZm6siWWDi6dC4JJP0nyNs/QUDXLaPstn69TNehMouJ8+tH
HsphYVZUKp2PUaau/tskXtaQZBpu/n3JcvOA108BauhPceqEeqAbXw4dqr8Zzx/XCu+QK9BwOPrW
hdrNViNwDcMgy2CDv5km41lrpgQrucDTnbeggsdb6mmEwvyXVqN4Fe0hGL8IsA1KEU7DEq8lcdsv
uOLCCLjNiaONmrBApS/7x79J6ZBUSqS9ylwEJeluC91pMcqQCSLayEOKphiOQihnZRG90ye2jn/9
yzguceBLuEs03Hnp3TAouyOUUacWaBq4vGUE+TxA7OFj94I+CacepdgJZKVQ34EFgUUjzC8JiVuH
Qkw3AVlEeubUDvXZea5KpACWaohfY2vXPn2fqdwQhHN2z7bS6b6a+bqdNCfmOYuFd2xO+98LTse0
9Pcos9XqxYSjBtksYMwTXEYvgWB8nVABlAnIzSaiwLuosL65N8fYFh+lrAyiRrJQaS/hRhcQt7Dh
gxaqAyEKtZ16qDw+HdRYm1Miswt4ecQH2Olji4H9yojfQpgKY9bFYuLGMU5JWkRnhrHaW4/rjBtL
nOlBxIrJ7vCD7mEUiU5fiv8/ioQfj8LxyCipqUsGQE66vifJyPE/VIcJCDkqFsmLnZGgU09f6lTY
fmAbiiO/iyelWxUoExm5YtxiKGA0gXT/C2d8MACzAHcsZLjMBzbVJy6aXX6V/ZJtNsajYmM23p69
T5/CJmoPYPp0MDYbfTYZl2vvN0U6Jvl63ypRlaM9nMFrbP6tNBDpMj0XN8zCNEZRNCPvB75onp16
fXqFbOLS6y1K0oEgaTTFACQdzaToAa4WOW5bk+TFVy9ZSM0pB20lOcD0fX0zRpHKwz382qUwLVha
JkJ40Wqa48FBZhC4W2ZwOgtoD/J/FkJhqC5LeX3z9QG4mETRSJxB6EW3k+eKyFpJ5hTMZH0gHu0E
3epoPICgynbu9Xk7v9U0zPTS8RPufROC4dKf7763kZMh2pcK/aO9uZPZGPGyhdJCH58j4NcHR4kS
w7SjpSgYmKxICl4Qe7sQN7im1fh3q34FlGWDBpRz32gRLXDrPgwCADwMFM//CSlqjWYCumnxhXEw
cbowoTJ9Zo0s4ToW81vIrN2IVS0GGT5qoIiGvpmYfqahMxrMvw9zdSO9GDfOu0a/vXqpJPMS0kXx
IQH/QhYmvkUOvgXVjw4AZrVcYB8zSK62ocoCxratp9x802QdbFs1pajhVE8D11AEkc3WoDQUh/zF
nNHvJZBwgs1sAPCuWUyCiiWwxzof1BE684ZMAzJRqYmcZ0LHvzCU/GrZ7HE66HPvIsiGznu+FZtf
xVranyIoGmzS4/qi1nCgD2zjJ5iFIJoRzuJWAvzreUYSG9JX3sbu/2amI53iWXwvcXT3+h+UmSZ4
BxGlEqsVPwJBP8wsjNQwBIOUfUxEIUlR+4dbdtgNkZ3UgqX2oAlhxwC9qT/IbPPH31RWTyhwZOGJ
qi5WUuLASdb+YodBQbnXpfz5mf5fDbKR5DYXb962NLJwGXv1dDnu0M0iZOqfoMzAdYUCQsDL6HbK
d3+cbufB5+LDcogLesntGp0yoNGIfx3gImmh3MAVlwQ1xvBH+iTFRxMytUHb/tpxtvIBt7pZSJAb
JEsT+XgupvM7enqudtRVDJurDtB+7Q7ZEY84543jP7O+yeeXlWylsLUgxuiddIdQ6bVHC+scyPVH
XgStedS/NkSwi6wctEILxn3RI6PAv3qahEL2El+yteojdxC8N1mTiD5ABhgBKaa6g1rdBMwYbSD7
PHi7lRLmzZleSATHlEZ5fmMsoIhWK0hq3mUI8zIjLLoEMmUKsJnNNBYQHfgWcgVVnMwxzrUE/7iO
xAO//mE4V68MMb232+UHbnylePgC4WsHBetPTq8VJQtv6D+2PJLiD8xl/2RZ5Dc37c16IRrgx8PW
4f9vkNdZSd2DyB1/LNaEObuHLL2uP4kvujAZ6kHf1Rkxp1U+Q6zNQb5hxPC2RcMD7WJgpAmnb+bC
eh3pO9UMKG8T3iqHNFRuakvf+yQae7RXVGHiqUAvUOYlA+UhOl9tYCh+H/u2NQAbbLqDlHJb6o4s
UHjlh12l/xY90D79bAHSB3IEIjyzG2BCw98t1d1zXF3bbiocx0iaodbTLaQmI+xG/vc4ooCDScmh
bgcVl/j70RKN4PWa9dSWCd3afuMF/Ng0RTj/x+QK88HT2RbhrSal9Lldrv+Wg8qtgXhIv3G1shH2
GJXtxaj9H5IMIXmnG0mYyDBvoEMBeFQSpPXWEg1KW1AeQrLtHr4rDBgyLPE7O1feZJi70ZsNmMnK
KcpCj2FEPNigg0sMdUppciPe2QPYp0tC2dJlILlGURIqFqPZTig+as9+WkPDCuapO42nRUM4v+vf
et2opscVHVUI6oqzlcDEBThnWWwOcj4wcdCfHKiJfaJfPsadHUEJ+WTaG8Gm/0xHA7QsqzpB8P4G
42mX4xZKykOEIOj/3LZb7mDs0vUjrxWZ/FwfJ9ybKTdFVMq4NwsazfJlA73iGx2qwZZ8cx3nvUZm
JrnqeEGH5f7/ziXG2VuQdaMTQdVBfIS6efR8znPoElXru69zHhQO8sLg/Wk8IaH3pktKetRpcPxn
ZjM6dJQPL1DUUhZ68mgSd5S+vpNKz7VpFHZ6RjWLLdBIfiyFJy1UV9DdRDsGKwDPx47bD+Y62mEE
sQiY4S03N4vWGFFU8jVdi9LhLWS4ucfruG8G6QAi5iIZC9WzseZhf69Qd+oy+p4FeLr0swXeuV5Y
0qFscxss05HZ8Y6Fvi2bhwkROda0kHP2IiXBlB34Ir1TF/p040qgS4TbkRGZDc0iObNhxq1EPrun
w9MkB6ADSsDug6YqMSgBLpvaEVZWrnwWKjWpe8GKRNBC0UvHEqzRm9wOeu3okJObdQRJClqvDDtR
TH6qNCoKKcsildKf/HnOefcuJ43JJihlYnr5sz2//kR9PMOs6f7yckIBprBojUUzd6aWXoMHJa2a
zPnv0IxH9nd8xHQ/3u4ETHCf1mJQiIa8YkQUp1Su209oFM4RxmaHFzaV9FmWjn+9REUYx1Ms7SHP
ExJ4ELtvs1Mw02qrb+1DmNwQmRAgAnSGTG5TBoIaQA36xA4lYusXQt+QXsS43jwtFxjo4nPYLgPi
oqe/jWRGWuALHB7F9QOi1mUvx655y7G2rT0O2Y1F2kQVlDu0r4Ag33paANoZZCRR+mwvjq5PGU22
HXipa/M4vm0Zdfa1avdmqLM4PpLOoyjsQWTnMH5042bzjOZaF5ff2jf0oJlM2Lz7C9LVIdgj3IFG
LfRzQuvYrGAPuuI7eFiryBOFhBHDxi/JeZ69qUWbAteOPRvGvA5z0UMdbzeqlnYwPRZLcijUp5tj
G2+zOHyCmlaZG3cDg2tXQE7vFBtmizDT0irP+XBNTMbHFUp/z/iXeFM52lYLE7U3CX+Do7ijYQ7a
pkS2oSw6kN6Pc3/UVKsaAk0trbQJIO3EY8TKN1JZZuF474glIMEjdwpMwEZW67meUcUBtS1KU9NB
OoTPiN4+awMQpfMq7eGjuRt4OItQFrEJFHrpe09dpUIhrgr0Ys8VEyNG48DcZ1tVJMNFOrSikE8X
Nbsg1y0+OYhxT+frevCu/dERrzMMTaiZ2ubRikBnx9bb0zMVi0oSiwgIRi40J6haEYWM0xgxIfih
b1IFPX6mR+dm/jG8c8bDvlloZGi2Wc2P2zJ6ld93CMp8sl9o9OIfa4hwBeFjaue8YpeVKhrs7wze
RqVjRBjOkldhCdRyQCoOsl0EnBV2YVRdt6DXaW6eK/vYLtpoLdmjRafx5TIfYZbnhcO0kKReRDf5
zWNgruMPGoqVahUI+B0AsaUggvHGrwquWBW+krvnsfgLOeFa9Y+nwYK5nIgW6bYbG85P7Ob3f/P6
1qRf04ZncC/JvkpBWTBiyfRiPMCIjgtC5Nzq3pNin7fzwRhhnZeZKoC6FtUled1lGTdwwdy7BiWV
7rVip1BsgGdPoS1UsSzAB/tdx9yx/lDszLdYvK2A+i4/Kaihi/xtycPu6OuX3qHSLN+LsaAzf5FB
isFoXw64hBG/ilSdcyJ2JTHLKODIZgKTS454dZgKWsk1OTgtJ2NSQJD9VMbBZcvyXm5Va9XQsM+Q
6wB3GTxxnmrFeVsUtfZjDmq4VnREEaMKStavhOqCoagwKwmo1CV28EXLN4btCk12djPELRGlWhXP
ZixlSKDmDyXFZgS7D+a9DSxIncMtgBsj7hdTKqZSkPPOsNthHoZiL9kgpjgzpdV47rx4chirQVAK
uM6PfosJ7GglsNILPqg79el/BRClASXqeLK9tuXx7HarsonYE0hYS3mQCQLBktmv/YzGklzBH/aL
ZWjBh1NQ31MFYCS5wsvNdjsbafuuiPspWeynBltvHr5HI9q90t5GYtUPEryUyQmpHSL+SlDCM/ip
lUI53QmgaCeJC/qStGN7hPzAq6tEA21BCUoWU3KsCgazsoL55awqUUeKbTKaxzX5ZdfnZhpN96Y1
U9Gl2wgb6qc4LpL+Gri3raF9SrRIbXQKo1waKMbmXyXkVew+MeLMWmL3s4OUxKc5OpY5p0OGUMKh
vbY/I+1zrYny9CJsFKfM4grulvcHYudGfzsCmQz6x2geH+erEnRf/AdtlPlIHSbHDH/pjNCEUXn1
jX6sWMVJn659LX12amrNvZ0QqFvzrdZFFSBn9p+/O2wMQVQKymXS0s2itBD5OHWjl8OCwypsxb87
GX20hlde5MMPR93G7tIf0uvr9we5ON5RFqLRpkf+scR7ZwTC9gouyGOo7bIQ3sWRoV2YXNt+4qTt
6YKyk5whbWBG6TsYEZpxfRtzcZbGhVrKPW8MIWy7LApqeFDpIHnH91RKhI+TwLhVWP5kY3WvK8/S
b67GsfdKRsIraAo0G3FoUuKNkgPTUAgluAmu4qy9W5KM91DqXUITIkTJZ5pqtkwcIJmuDl5+/0fm
uDn2vKQRSmuJlWR9sbfNywrAiLH+oO8ABauDBYtw/5IJZg9pLFsXVYhNmhHCcu4oDEVpv5yqcWaY
+LlyDKM0l9LZvtJgL6m7gB5z6ZjRjB8BvFIf8qqPkExI3GCTWrSr6GMikzHK+3vEuNUrbzSTLB/7
YiADIrPFDkCQjgWHU9pZpkcEQTmQGWoYbocqgC0apJRKfpLJVZrNy+LOWFk50Iht8mE3T+eippAW
OrnRPPnHOjA3mVcxq8SSW/mK1R1lkTRP3XdaCVMu15pAdZk8BN1akNqah8R+gvQGuU8euAsdxWsc
G+n70txCxAsSX+Tzpo6M11VRNKF5HtL5UICitcu5FBXMIA3QoCCxtO25EJlanVnqTy794kC2aown
wbdxXSlTQ457CCUSDMbDU/y9RAT30buPdIwgks+MMrz2Di2G+VC3MziW14dv/gNm1VjrkWoNiUOE
SnR+1dOO8U6N+uj84zEGKq2qveXG6WXufWyeH0OxXlQLPG35dLPqd1TqwMPM9m45rmc+3x0GYguz
XpravENoqOrauEpURZpjBtLoq8RwvUlApVqbOQBZ9Q73S5Dbxd6N5O22W+/XQiKWW05klFMcQ9cG
XpkaTnh/Er36OqKIYLIhbTgIfuiOeqXIs2kCU5kJS5/sfaxW/G5eeQi6X9pD1iy6y7Ebt5MqIaUj
X9Eg5bQhibHtv22xZu1Qequ/tat2Ct7H0T1yOxDcrkg7xPQrRDy45fW74kD/D44+vB4gDanCkZMG
S/MAVbbv2pXNuTsWJOI501YDlNNcnhErkzUJhSeJqakptQci79xIo96kV+xMMldcFrES3tHGsHyT
5A8mx93hjLvC7MIM4gbu7Lyk9D48W4/nd4rn9iAMf8JzLkpLTzYdY1Ot8K11MzHMLCCVI6ZHfz5J
v9oqQKMujIW4MRkeTasrDRsKEkUOzUBLce8jmmae/2pS5WXoTauSO/AeDEKnLjH6+kLJXnMBjTks
oMEsQQttHYcvMf5rlvVm1n8ER4hvzCUL6sDc3VkhMqhM+Uuc0Iiv5Ervw1M9G+spc1gPKtjmbwDS
HEZhcwHaD7NemJMa3+J0/IufL5XCAwqypAzD+ISawoI0gYy0STt+hhmeEmv/QK7W1Ie9vJfFc+x+
IpF2d5iShdbuok5j8Q6Eo2oP/PG0dscdHTfaW3vJ+sdNAWEKlsJ/beupYeOOdVIUSjO+opyb1iLh
WYd9WWAVHJWpB93WW+as8EYI6Ir1TbrxJLfMJtpKiJJhbq6XHwb+drqo57winR8pEABMkch/un3q
rFMtNHZOaeVvckp6UvzcYYBJ10fKPuL+kq79kVJu9Ufv54waC3M0VlQkPBYq4IQhb3ruQ0xj5Fu2
Sr+TONhyP59MCVrcPwPVuNzLOWWm9GYEJSjurJGU7Js8RecqDwogSrBHYtGCNdMZeYxAQwXBiEaI
gRttKV6UCji9l7tbJHwYKfzjjj4ZPLDdksan6dcukcQZ4C5ccLXyiCfitqHnBj+sn9o2R29GOLWZ
/Qgcu3rHDDGDPRhlUqNtGcRzFWWD0svawkyMtEF4mcPrZuy///FTMmFzl6aGkmfFGovm8jaebvnd
iCpcfiDIuPpUrIoI6pkog2PZdWt3Cf36jL3qr0vdzP2GsF5zfQHYEWGGFz4dyOuGu9w4Q9Rlohm2
vN3DayS5YZvTHOmRXFR0XoO2P398rRcMtKcEj251U/BGQ93S7UalTSFIlsvrx8eiJ/sh3XTpL+g8
p2Pmju2mBsof0lF7NIvID6m+uIU7M1ncq1dhst3eQjiSB4f2qdooH22XPL7KgIgv/ysQhLD105mt
HTzHaS5nSI+y3xnnEJ8IJWTm3QswUPQ9g1G7RxB3f9NH28nvjg86tyiFBgCus+4R8eVF0gvG2GSm
O86J46hUT5+/5dnqZOWWW637CooliVU+kXYLXP+9PfyzYR2gotjI+0AGoQN9aiR1Pn9P3rOtAyo8
xuSP6FcnFcywwdCzVkvfaVFSD0EERkW80LHkdiVlG/P1lXv/RuCcHOh8W1TkYL58qdpUw+IK3gdr
LyabZok5EisATz1OSvz0LGO3658OLQB3afp40IK4LV0AK7psF416zk4VP8xZtGCvL3LixLlMIHv4
xbGfXinsbxetbuceShstf3HziLLODHorR0Yvy08p4Zpyc1kTb9K4H8XktzDp5IjZ5mmgYXArlCdO
QA29rVzKzogGrdp9aI3jtom2si8KCOODunWppFfMsXJ+T1nnnOVIFUj3QfNeKdwqHcrTeIpVdfvA
p8dJpiRN1kWrdB5oHOrnHtLcQTM7SctDQQndcEipeasIVeXwHdDbq9nbGj/AV6GQV2zJe0uF/l2W
6EVLnU69iQQi/zwnQG33Ov6dAPhp6WiQQ4KMwN0sipZoH2pn/3oTGLlZzMJ90OliKR0v9EAQ6loz
SrfST9oMWJGzsUwWFspU3PtvOzoSI50yZfb5zIc4FwZy1N+sORKWg8UYivd6BNfutJRBObKADA3f
mclDlPRY+IP3aMPdMBS+uIhfADGx8ArIVFQjibW/0ka5qE681vcwCzN0bXihbVEp559iXgPnTcFq
NqUIVgzABJjAE6ECuigZQXI0+tVD779NsA+psjhm4/j2f8Rdp61EFrx6LYbz28COixmYTjDaLAUN
p2690VimDSdd2Ou8XNnHb/q9uO1yoFDmyI2qVkqvyYl9hteA2GTw0X9lWBwlUAXnomL+yZma7Igw
cLhJ0VYjHIfS0MsDQikYFCPZ0FHd/7z8/crsSzGxcF3JQ+bZEfTB5rdQ2AoYzs5GDqdLKL3vpiAv
3mS+c0wOurBkuJyuFL0B8aynTxM5ttXZRptp6o2QCMuh/w3X/HPxGS4jlTx40ZFKprLwotMhSi/d
NyGu/wUmugJlxRap+ISsneQwBP+hi/0FYihmCpNJd1KtAdgrFVAZM5sUONLGgejDWSUdOhBI/UNE
efOm4jfwkpJ0pP+nXwh0dvkiEuR77mVd7bYYencOVXoPjRZHMNu2jXOA+jbTvahRR1K+HNhfwNfj
Et4IvxVOtpsL8EmDltIHwiq+JNEoiUa1WG0wIFjnRciV61qeoHYbVZ3rrvu8CsC0DxKRl0C8j+gs
kDg9YfhNPNBQcxyiOxduD2fZp9rmaxC+GAAJZ6iHQvQbYfbaDO3RateA8hYtcvfKa211ekToP/70
Sjl63RLeYQyKT74NCATtmFXXOx1w2SnopV7e9DjMecc8/8legF4oA16uk1VbTfKj5ZdqMR2ApN4q
9pq2Ja3FlK8skwjcGtoWO+vu2elcsb2JNTnqwNs6HXSzGa7TqizruB2ltJM8kTUFiOd5zDeyxP3y
EA0jBM4QKoBldXtNlGD7K84igU97d3qn7/yZMu9xuJPdXW01QtmO8fhWDWrNpN2D1a1K6+PVx7If
eWKiqGBKpAdyg87+zMlc4g6msUyOV8GzTVFomNOI+GSE1WO55ZRplccfQrirVxjwv2V9QGiUoEwW
JEQQWrFvaTXPjZQaM8cAdBrHS0U0sNx7SpAELqngoPg2hecMls3++Ka47nviB8/PkCbtkAbbyip0
HgZNu26y990HJBE0oOQFD7G1H+F+JpOsLlIwFrPf2deDoUN2LYOQUWc7dW8AsvxJNSIpRYitnXQW
ZNb/oesZSbYqS+wV5J5EQlzemydD2XwcsxwrTpEb9FWT/dx0Ph4DKSsOqX20+LH8IPvh6FZkc+vF
IBs/rORVeSRhn5yTdpoIXXW6Wt/w1YjwITopisoe3It4fbgUbOa1CjiTH40q7k0j3PUousOjbxkf
RjFYIQd1kbKQao/dKs7nvuXWkWkmApkTNnhvExJu/znkQG3q3s1zPSL5NHd7bJGp1RBXbA0v1Fjz
EIuuyCyRJv41m4YnCS1mluH2tEvSb224kr0TR0LdGo9EI8ER17zWTF/lPn/jsSCazMKeGfoIn4Nj
Zjr7y+VhZRHlCy/bvnQvf+GChbjZB44bRLwckkDsvuyninG1B+c/yNMxx9ZdDNn1EvsVhIbFnBj2
3SCfJKohtvvcx9SJA4Iy9xPjoDrIGudV1VI7wRU0yqNcUxi7UCtOjFHW//M9bP5MKC/0IQmFdQ97
EagIJGjg1XWD7H0HOF/kyE+C/rrt+Yhox91cYSFKLdVU6LysJ+ul5Ifa3xbzYSv4vCnb3rcC7/EU
ZE+0+GyNxh5jPUkoGkbd1Joz+pnucPe7qmKOovA7NNcCQc5N56edxGMQsvF81xD9XyZo1FSal2Km
px9BNFZcpybz+zlKbfkcbVYqlLrvGv2rcxaAR0++XIfHf+2keUXP+/M8VbgW7MPTWnnoy+5z1tLp
V++ng/JCsdoYThytugI2BEyAgsfPBR2hfcZtpknjw/zLqOCYdrItU5kqhZEHFvzyfKGmWmQfmoap
w6NDEHmRbQ70ryuFPdA+LVkgxv5lO6DcfAiEsEFDcC5tN5jYn2gyTR8VUcT6rArOTqBLAeqRpA0R
/1WdPUpK/oTyJO9+chIs1jqgXMIRSVtMgT6hJ4TqPY3+PvS0MJpjqNoms0b9N6G9TV0eC5HPnhgf
7w6iZqBfYdBs8h+1Sskl5M8RA+328zTcTSInk3ubbnnOPWQoxboy0bxB1R4CkX1m4r21WzMC7lxM
dEVB0A/JY3x11PMjRVcUmBB0Qgz41iizfRJ/XEyqp0GFk6XvgQ7Rgj+DRm0Z0yuRk+hGVhEjEhQY
TEMKURaj1ZOPfEmRdOrFx52FR6qqGwyvtcHDqf31p1EXS//ri11wCvutVNT4deIRSjv0KiBv84DV
zl85HZTi7LyiaqD4Gf9GxF7tUfrAmj8I56wSm4DnYOX+T5+QO69uWIeSh2YinAuBPF9Us6urmERe
RQet2CPgXc2gNRA0pQE23VqstIhmta4AgUngJEyRiyPgYhmOPERIengwxop6iT3CboGwXZTW/FtK
UovoGxj3zI1lG/dZoSzHXMBPnFFOQLKeDBA3Sidmq58sHn3E//rpm23+3Cp1nh/JqRcxS83+n6lp
zz+aVOPlvM7dDbwqvWafqKeASuC1eFMwnpE7E0X2DOyBYweLORcTa2k7AHO4xgAPbRcJCeGk3jGh
12p/gKhDW/f776jAavmXbpsYN4wjXow81mBPvy8bFsbI0jcKLEh4wgBC7jw65OAUQZNV/Bhoo1Fq
KDykEIXouLFp+deiG4IvofWt/FN8WivDzeXasTARHCft5mENj5KhDhXeLmg8V6tE0/wSLiZw+GGt
+GkyxpDgK/vu2zbRtd+lVauKuHRGzjuYJHaeKKke4SQ0Ht7G118hBLnUcsrp18K7b46W3LH6HeX2
kEUTk90CK0x9jxDhyAo29BS4ivvcrwd3OGSZ//P7w3Ywd7DomzRG7eDyOsWu8HOM8O2sEIb7ab+N
oZ+29g9JF6VCG4gXkXoJTu76QBpRPsMJqmo4wIbid6FnMNzBiAWvXvEIuOuxMODyM9pQFTiEbeSD
JKcNNnGP8TUOu91jRX2qv40LMvhL5Fz9EsJbPA1SS7WzBBdZ8HcjQw+zDMLipp1w7V6uNgOKx/vA
KBE8/BlJ6x8rCtqP0yAAHVZKYEXUKYDxBx58pnQOskpqut8sTIx1OrW3QF7lsXiT3AC4mZp7xxuO
l+rMai3yGLSJbqc1LsmbBGmlXRqL1sx95CVDNbgqzlP1hAjV4dYwYyTY3nJ6UfUK2VuTs0iT2DFu
v/fdaYl4v5vfYTM4KVy9BlQ7Ez+KoBWZWzm73rkf2cYuej3SMDN92kg3jFvDbwZ2ocwHoFuSHEdV
Lm1pWflr+Rrrm/t4W/EI57CaVAA+7f2Wbmg4Co7kdGfkfM2wT2hXJGSqfhEWUhy6xp4veqIkwJIO
N2OFbKi6ONITIyVg9b3fDyz/REJDTb5M1zesAn83DWQ3UfMo8TqBOstdsHafWU0oYsRH0oAoBliw
UaJ553Lpj7v5Yi6R3G8T1kveziAmzIKjT7VYFO9YTmR1BFQSq3K2h62YD4dA2BS52T3K7jsnjSUg
BqBAaKkak/k0+hk8RKrFTA3tEI9szU7ipGIHpNgSebSh+qqg6CEuIOuzwSZHTy3Rp5T/pl5vGolG
kHmz+CsCLwPkc1tL05qkZ/EV84po829G6fDsEDGH6vGHI95u8NdMDwPSoFpgw5aJdKucHk11Mh0g
7CZpxd2OzKu/ZXswNJP8YsZPf3O8vOlmhaqdi5Zpf/dkiIeT7iiSxDR7D7TbTcYh5VoZhPiGUMLM
4u1xZvD4mgKLpkTetUiOAUBCcliy4m5wJ23U2Pvj9W7yRymqfSW13uoI0w8UUiipzy8G+v7XGQbb
F/oCumlu57sNcLJpXrtGJxn9M15egX5RSAF+hYMMw83J9Xq7DBwJ2m+iBtWXVstTHW8wUQCtHnOH
6a0tk+I/9BV3FfE/rBqSQxMuLZpJZYTZxNg8Hfv7DLOyy9A4eLgbTRxPlvBc0oq/D2xlCQcBRYz2
EuIs5FEz5P6A2dK7K+3X/WeeZ1WoioC+/L6pWkEpSEiATdOAnD1kq7v1oEkl/K58/CbuRL8FMR/N
M5o3j2zMLudvfMu2hKIOY2h+wtNwpolE9ub5w2q3iDWqoBFXUTG9kvphCfJv1PAjVqiJwWjEPgwN
s83440iF4DNwZBnrOHVTDdeXe37VyKNJSGFR9ALN8HDoZ2sk8WFfPDROe3Cm5tpsApMB4duibhf7
3PbvFC8VNUpRVWrmU0YBp+duIjSgovS128l0Y3Y0w3x87jQnx5uWij7pdfwoxPtpEd379eP60sSH
S6MAdIbVrSqtyUVUIhUjbg7o15Xlx18xyXtloc5P0eAr3+LKA+kswuRq0R+KVNvbgwVtxYyQk9ZQ
u5/N3T/UGmAFWdJOomw9yjuKLdh5HZl/DhnUI+wuxHsIXyRWWAJmwiCTkvlATmEHHzsglUTDP3p1
C8fS/DS2qbfwKgeImbg/+o9cV2L3Web57FMs3gb19fL3vnmDWwxzrHFs4ZLhMMKu+nxyx8WyNhNc
qO1iyCw7GBeYq2qwy2IjW8oRnlYGtb14MU3IOroIZYa89Uj3bTTQVQcIemV9sV/xWGttiJKDApex
uQLnc2pJWGVTVxZ3vEgrx+vFXBD8eB4QyN0kCsdm8ueNGnvRKaO91/KdkOJm6xmh+lrLNgWhTCFf
xULuZqQpJAOztE6d3VhdXCWZ3fJ9Qx4we7k97P1i1OcNaxP4OhU2ICLA5WXpzmfcs/FXD5xSQ48J
A/PGudk44BP3H32Otnn+1jo2x2zNpT2DhMSoLfHeHpC+RXTW50av3qunY1jjJ8O6sTce3LDLRGRc
2ICKG70uhsk1Ubbch8FEs2FOyatqg36Yw540tEEgz96hoG0vQ4zeFJs0qx32w4BABeygp9hYuH2N
Mw/N2loB7DG0yLN0+6RJaOZuKX2HjPbIbMVUdsn3G7kMBJyxaXFSkavQCaHE7uLSW4hFGRrx/5ZK
SnHRf6G5perBh/gZqO3/0SuU8IUAIbYOflXQiCO6G6ZkM3iV7WzrD/6mlyGiQi7D+NG5O95XlaU8
YQal4ZtGDNde1yUuAragmlUtvHSRtMBvRPgFr3jH87vziVnIlGaQNInC5sBw1K4OQ2NJvYy4XYQS
nMvCpJyF6/a6AY4D0MzBBqm+3mZ35jr442VIanXZwG3AARYM3sfn3yBlT+/gGWadbMU9BJUllMlY
Hd8DieTNnqc1fArbW0Mf0n/s1/95BT75jehtRbtN8di9VlSN5DbqkjqcQUOOmSKmn5fk20Q/7dN7
lSLDTYTi5znH2r2C8ZslWEbjatmblMbDfLd6b8m3Z9xETd1t1QZkW/vUUK6hx9Ic0TxNtsaamQO7
Xml4fB4TEbVlbR6qy2j3gVHeYABmfw9fuWTdYZTGktdOF+WE7MIKgC0mcXCyx7Y8Rj4szvs0sPzr
M4Fg/H08hoq1rezgpz6sSEKYxrnnA2aqHP3ntNVMQ8CWfsCoDVND//wJm229yBkwbc72SG3NFHSa
w37r+5M6F6XstVr2gFEA5uyb9qCae1w1SuVlVV/4TQ+rll8Fo5g9s676F8V2uc7SELdITwjwMSeH
3lG1TWzFLmK+Fie9DHN6YPXgHKFuNJPshyh+tX1kqByXOJPuwWZb8KPfvACDs6Utudg/PZKdf+FU
YB2Pp5zwVIqGWkenoCXNUJx59f7kPKoES6jmiCaDKKmOfth9kqEoHid8bWAZ7D/KSHPlcclNmbPX
T3VOPmuZq5V97PIghmRVXEX5u8r6DFNLeUOTVbKdeGvjBxkVwE9kn3G8NeG0f4gwkj5zk7LeZLJA
s8Jc8EzBMP4FifWoGu20tm9CF8CiaNA5IpEkRMSgFThQXD7E3rCTKls1nL1/42PCMh9FonfQr8ij
a8ggQoSHemtAbj+JJ3wjfc/19vXcGVKBacCFes1PLTrg4Rg7x/wsDnGTNXC0LPk8ZCt2xIpNdcrr
JJCUhoZj6BEs+s3DDKmBtkQS/3It++0/f24F5OzbREY04QkeId/BDzHCbfLvc9lHFI8aHiurEcZm
xidn80pqky4uiFbMVCZ8liwksoZZXSihcbVZ2fWaWswoEmjGIKs8Bl6VMdPTMfwdPIsIx4IY1N1z
Bdb3yKfzDFywxIOloHNNzfy7h3YNoeu1/xRReCmV6MyXOpYZQ6aAl/GFjRQTNOm5vcOVv7sq9cCQ
lGbYiUhbzuthYh8uaOUxRzenuyr40TyEMTlygCJZ/fp/5J0KLNGrlBbNJCVVY/fTSo+j5SRIWbB+
5iNjTM1b5u/P0u4Kd2M3NCW1YslZ1mdOPPFPRrcQ2I1/Us8RkTAi6rJ0shJCJ71lqVM2MxOqte9b
2Uxm3J/XzVh+9v67p/P6HRONs72wgJ6Xo6PXrzhPS+BUhqhMF9ROP3adkNGbjFq7+hyLTe/cJ+AM
iBONFW3osUsUzlPLht7ALLoS42cZL73wrB67HgrFR6wBIq8YdsCEOkQ0J8P115GwfQwIZi54Jfn8
BmH37AVe8r8nsas5LDD1BeFikVbWUMw72+0u4AT4LllmwqbtMgr9veM+rI3A6w5+8Z8IbvyMwfQw
2aWmcKRTS5BkksnBK3PP0TTkHmQ7HW6GJvf6HYJy5sUZ3uMYy7aKnNzJ1YiUWbt+yabGDJHb8VoT
SLfETnLHUtJEt298fX6Xipw4tZb2Xj8oDksNhegPjabSUPTnnbicNDxNGQ/FlcaEmi4QwqzvQLkV
IJpFxEMWxV0F9NI9jT5Ud2zhK+tlGuMJUolOwmAW10hxP5x/jiSswexiMY0BLYQBrQPRanPxR0/X
Fc5WJ3Q3ViszM+ymGM45zBxKOjz84rhRH4NRsoy5APCbomSsVBc4nMuGRHU0fuSe8tLmCMAtAwUd
ogl6kf2vZtwZ94klM324OQRxYHkYQq+aEhRgGGzponUQhLg3wFt2D8RiVkvpcGRdZ14joQuLFLtd
9APhVaNSmzZU0srpV2SwdiRMnDBV7HFLxsX6d0r8oEd9YSYhFBzQ28oYTBRO9zraO3hJ1kbzctEz
Q8gNc+MyIUfcWQe0WmXzOn0Hc/NDhrefk9qPeqzI6PF6KnXXct4rBZS6W0MMBvs0jgrH+/mkx13j
iQqCCJln+8UBvYbpQfN2+wIxv8F2ReBM14fiVFeWu0fKaYxrHr/7IqKGpsmOa7BjuG50F3aFbv0b
ILEKJwU8lHcmuNHF6e/8kIjUgPSA6mL/GoNF58Gbus9SVX4eha10kXtKcpOXEtvK3oE2774yXOuc
4qPHBtKqZwFYgKGQMyIJvh+es6eyuRRC9IXcZtQ4F+oGFg/pp6Uw/jcAq7eDwW0EAlUr1XQUGZza
iY9oZj4iRCmQ7dUNy9Qkl6OnugBHk0g9qAFkKMWQlXBOt80DqdqR6nICXqG4BtSfzX+xakKGsa3N
8PHGH1nznikspslb6Q+yx10y9ZViCWDqCF4qiXgtk/TNHqwP+MWFq85yOcpqZzA03YhyLe9z221G
1RcgvgYml/rIScWK+oNBtsXnhTJAYPOTsgB/y9AuUookYP0bOYWQZpEzzrsP/0R3QVaRKazf51H1
gmsPitVI1axVNuV+IKtNImpEBIngaEqAGZudofUBGbRvPlm1k+E0OxRxw3aiC3bOVWQC6uvJyq2d
UyhlMWs1D1nSi13YoqZAiBC8oIPe914hXl4Jxg2wKsU0r7o/0EHd0nmP+/9jAu3yUtVy+IWx0Ixh
p5EN+DE8xVA5bDOX5IbzOpjZd4eFn18PPV+/arUzAm6tAMpICiIDGohqGVitT8k++zNXiSArzmKR
oboHX2fHmzspFeLgR8rJW0L4kkPDpaOygnvxCqeJ/TREW2J+2/CAG6i3y+7rXi0zTIgpSThd4+pv
KzR1GJ5ThRKnXmmuni0GJrjOOPQ/RvZyycksCdk4t2o7e14nBg3fHGAf+UpOCfZpFB2KC6iixQEw
7viF1RYpeyQ/bkKyy8SdxfaQspH0VHC5W2MI/k4WdbCXzL8UFtSrOuqA1FE7yptGC0jTIUlqYCpc
LJc/sDUNvRIRChh+2xEjA4jX/IsuV0ibuWbQ0yvji83Kf22GEmVbTPIqXONzp9T07gu19KI7r8s4
u6JjLtV/55iD/YNwAR/0qM9MgxPt2iYfU2WXARIOu3tWI3bQgzbeNrRMka+TDOfMxKBjvK1iPSVA
OXGVax2dEqS64z/1CsGagyC77rXq1jxP1gJIlXcBAUezE8y8ZZOgQtGI9NWSi2l5L62oXNjov3pm
Cqek1hiwNTtRgazWPfametofTC7/ZskkKfJZeT+Y3wWkTyPNL91qHOycfIWyEzzVPHIHFDMnTU6E
x7taDugqkecXfA/mJOneFjxBMap6GQXbAGiP89KEb/500yzYFF7P4FDTPdDmJ1edaxHNhkdJOgr2
tIvwF3F9LpX7MTNRA7n88hjJPTNoG24MH2y90fbD89Sp+gq3XBG4av+SZivEDyzri329gFFlIPID
mEnUBCLbFgYrnG+jFbQ8cfsP1opr+H1uyvAUAQE8qL+RR0Cum1ExLAt27qdD1xrc693ithb2WJ2F
umhb51Tflvdav9qJ74q33MpTGeXR25GBCSIIZRhwSmD1gJK+lwzLPuTTZlNNsILUaCyb27W0amJw
TaDhQxbzM5uQunxiPJCwxJr1FBmtM6BMQwTsKN58isdQ7JF8V3H2cyJL5xHcJiE7tqLNWncKxWbL
6BLd7Llyfs3phoQGkjPXoN44vkxZvdcm8WZhhLMIWxoVM5Mzac2cFqb3R7EOrACojmf8FTZ7v+Rl
RTv0Z4Ctd1gY/fd6+w+RSsfGryFdfyoNbwPsL8Hg5/UPGUDr5J28qagWudKVrqWZgpCAysqdnjCI
IbHCoG0V0ykTPZXnkjhxHHDMrfxJxr9aSD5g4UFvwbUdw6AMvmEAsiYmslMm9ywj2IfD1QLty9Po
qRkfFRRP+zgESvmJe3KvsUtA1MP0h6e/HPDKEUeiU1Uk06hIB+Vvkw3i5ysuA+pmmHyYLQPilVM8
i1unOe5D6w3JXAbrwaadTdymr9NcG5bnojv64Py8Y+9gUamf/NmMi4pAAgnjPoBIw0fmRAvn2qLT
o8JqEXUuptUtiL8iYJW9nWMhI9LK+xAiGyQYS/M8AlWb6P35A2RjoKtjIIZmGxiWtLBVNUpDABQI
GTaD9r2gE16RoeYGZvf7YyH14l7IWAvXKHOaxlELqt40ofQtnplN6UqqQPJYSDrfJ+01uN6vvb5t
kz33fajDALNWWQO8iKYbvdW4OQAb0ayTpnXy98IIjpBlqtAV2GrsZAcEYak/lcTSlBM/1bXwglFE
QUy5uT4ojrWVbmK4judL80SKG9pZ3VZEw8Z0j3KMYc2vtA4DcupzDDR7NzlebRbwj+AJqS5Jmku4
zdv+36/xJI14MpJ/GFpmi7wAPQPd2EpZtGBg7s8VQbIsKboA/bBtQo+tV6HarX+MFDrfN+hRPfor
uQVCkdrBREEOkRpoR/X7k21G3nSpLLDYJD+l09JEokfM8iEM04HgY2Lhb8RE45fSMQfUUFAiQtzA
xqWSNpFga5GmR1dmfCyPJJA2m+nmC3b9kh2pUPPLr0yRwe4J0FAqTZlbh/eAz1PYol860H7JRfav
XPuH9tu9XFF6c2ZZVK71OFvtKeqCYTigW3R1l+yEswIXIX1zE7PVISelunQ0nCw0Rtr/P57VMSR4
eSJeeDvGiOzfVvmaGmNEjZq+fqy1OEh57P/OgLaAMwhGCMbWYiiUo0DgzsMZomzIrd22gnbwmx4+
6MSzzg5Qh43h6+wsSIv82ZxGfJ+fHqRFMKjk/fCoDhzWgQ1cBxlf5sU4iMRUcH1ncUYZRqUSzmCU
s5VgmDdw7pLU6/CrTrPCcZUEqXOjESSfVPl3+r+0Y7Fpe8CatBiVEPGwK4qUNvpHXOJ4OmlfhYrc
UYrNlgh/U2DWFo5nk/rig5hNniW8dYEkrFR4B9IDp2qE5YubTrZYMV7LmizlRMXfxsQVnpnR8fzY
tf6j15Mep0sxIX2Snjcb/yH+k5aDi1tWEv4FaT1JDwYYB4DEqQVdqftBoi4kZ/OZpFwwVmUBVG74
sZszgqAwbp1ttj04q2XyvrDJHxFPcz97dxeDW7agnJI7GRT5wdutIUhPkAHB4uyukcR3T9MPHJ/7
n6qLR2TD4STr8ti+AzlG64WShbwLXS/qvZFc6xNRxkbVhbst/ygiql/LVTF/Hv6BRgqPGKGVF/pi
NTk6EGON/c15cfbERZOEyIPmI4BSov/jUiyi4qfJyTMFX9zAkWUshIBof4u0xKGF6jrAamKupgoU
rweMPm6Vnjd1V7B7Z+mMx7TkvXp1pggC5idBwsCaoWT2LjjRYqfUyslxQTOcT0+PSdCRivOY4STB
0+tQOHeLORwbZoY1rxgLBAJ51VRdE49TaDdfZaU0/N7IDRjbrUhWjn1fX7cdljpzt3JwFtKFPPPe
uJ666KJrR/IcAnK8jVpu3pttJQIqJrhov1Qc6wIeq83IYpfYimI99PBNO43YOYGEYrNOf5VYGpbe
r3IQZWID1JKg4XkmomdXHUrfFLpEIa8IufValk19BYGwTA12O6DNestplu5cmaTBCR588BCWh27t
6W6MbE8JwI2zxmT5rLrpmPeAu/uDv9Z5J1YoQxz8pGie2klTp+eMVifS6jzBv5TTljQLPL9hUEHK
PMzdY//vyfoJ+4XFDt63zKaBNI+fOLO8pJwBTRL/hMFJoTxIFSxVcu+ikcXJbGZ2pCq7/DalCW/u
DFd4ZdEq9lS5FaCkjOWZ8Ob7bYeLUL1pLMs0VbsWB2JaJK8DUvodSs2V51LXkkWHNqiRUufzGd+F
BE/xjZ9Bc3UvRuxSuL/HgBlX1X09Ky/i8On5iJhbJBdyQKYHQ0wrAJeBa/16qi67JOa9IOjJXRuk
7x5tykM8SwdjScG5pq9NWE7B8vseKgfjTkBsh8Sz1VTHDWbSzlIbe7ppSIrRWr4d8x1cximijIzU
iJuKKnvgMTJs8Bpr8S8/rm/x/4CPyKgijicTFMi1kBNToRo06zJ0ve+hpl8s+zIwL7iJ48/U1C5y
eqZ3ddgz2nEQ4I0VmEgdRVN3LXMgj2RHnbyXm1yO8aRQKajMVGNkqMB7fZxf+GI3Q85NPWfVniLG
dW97u3MLxifayS3Qae/oyYo6UFVxILXcFZ5F+JsexBJXDFeV1YbJF7+27W5HNU3NDzkIm267cAh4
aDeaL4JTXOPYZrR8AadWFPFt45R0IMbgT11meewN/obXUCHrbbpLrXB7qIl/GPQp5FjEJlE0lhHp
xS8BmAl6SYlCwllehuv4IrBIz4qvx2xeoUqFL++hzNXipVBrvi8dlQ1JXN5/kMpohgf5dxu79M4A
Hckfv1OSReBGaFPIu9Jng7yb9/JvJwuk9zU3icQWffioKOOcDv8ela8x2NBGa/w9gKsNUUOyhSSE
sd4JMUUOKXlBxyKGZ7+5kl6HfZKAtidpXPkkRQsAyeT3K37/1N6L8WeZxaMLJh5Hyji4VHj2g47Z
r+dLlEjHoL6tFZvXTk7hXq7R+X4BRqEcekIPzMWOK4ARrjDa6qWJp8By5w4ogT1FrdwE+TCKpzsP
bTkcpgzOv6ZVZ/YgHE3XfzS6Awj1chmi5TYmHftXd/6Muzr6inOnCzXWPTrCtAKnRU5kJb2S5Vwg
ye+5ndTkgLyx881tLivgcg0tdMc/00LfeP6uHPzdzjUY09XenyNK1WgoQT/3Ttdcq+dDLhtDFnFO
qc+BkBbyKHSxDsTtHIipFKuJO56xdB857AU72zlYRnEPCLaIZ950wOZ8OXZSus1ZPDCNmil1YVKK
zsoWTUOyvmfnTyLipJJDxHmwIS3HSlp3/0aapT6b/ZUJp7ZCRsxxq1m10QevFWaMMB493Bef7bs5
BEhvYZI9JfOznjFPlIJOtLMG3NfjZFWJOQVbcZas62RAi50uLm4pdRuSm+tsj/dghooXayAyWJSc
GMTRKjrZ0OJKMPJrFSQT/6ZjXArXVYgtvqeVN+4fHGEhkVZBbf37aZd3uaac/7bXw3zpBygUI3kb
ho2mCr6y2t+C7VZrsH7/6IV4ZobELFu+y4OWKIVrkuAtHZCg06VKzSP16UTxbNM7GxUMjyXFWp5U
qxKotEnS5hZCzqXTEuilXneoUNxMtI96uSwPv8lX1ctFT1NPckRrCa3/gF44/THrvdlKy7K5nq7K
dnK7HUhLyGhh0M0nI9KLT3wiRLkEdaqFsZulXrWayq1MenTuM2xe/GA4JKd4bZ+9pwAz2CKOanzJ
2DOoJJ6RNyFGkXDa7vJxVqaPOqd1IQ4WP3DxhxvnaJ2RtH+mUUQp/8sGRemsI98PpVEd/+VcyZb9
bYLfXoTfdlTr3H9DSvIwKjPoobo4WZvSLZ84c3vzjAcqnRndsM2RGjSDFwINpYnzPv6mJnQIpvYA
8HJPpdiM4DnY/r+DTz8BXbCGQ5bmfMolW+DIuS72t6dfox9MXzOv71ct91G4Iox7bw9wSqxQKRHo
4Ie02ifGfHABxdp8e4GCQmX8PceJ7+rXhLf6xfzFmXolKvuVPWwQrT9FCzLCSiMzL4b/2Hyo3IgN
8E7kRVYgv2W3ZmSJLvwhgx8bgF8kYVgZffEZdpIL5T4dED/rvBmsguA//6dNj7JHdmpT5xS+8XFg
tD6giTJiu2ez44oDKYwKXOH4z2XAlhPPrTsTm2w7/ADM6VoARpRZ6Lh7MuKJQFjhsJ03+jOnW9Io
oobCtFdM4hIaajsGofUf6zEKAtD6dwYIisXjBpF2qR9LRTl8GdJTvIGEIWmuVCW386xYX1hnPfmG
cducBsD64VaFomca/i7WzCgJRdAHT9yWAg9DZwld+iTV1AIYDMn/GEVqV1wt1IhiMRTyOSnTZNwk
BKfEuPMluce9IP/4s7PqNzPkQws0zKorWtS2hb/j6aOlhYdKVDtF3Wn+kjojBKG8IF2ZorVg5SVi
h2HA2x6FG2aXm4lasTJBt80rDA200oiTlXSpCFBCzatgdVT93UT7JznhR3XgMYZ5cF/NUz/0GFOp
ulYm7pYI5P2n6b3e1johjctcXRiAg+blSArgkyc720I8msNIsvgGHKd2SDZDLucYfWXznsf9LjBm
TcWzD8lR3mK6SDeMSWgrUOBuFclt+fK5nRRJ9trQvF4WS4YViSmPRP0wbKc6dkH09fKR1bN4WMq0
casJ39VCdjTAJJJztc/dCDnaaH6UQv0lnYhuHgTVx97oxu3xdUplxlpBpCrTFE37S9LV+4m2cy2a
3372IdheEnagglvOHuj9YUxGXnEjm7sV55Oj7aRjjaKLGR5toIx5JBW2p4fwt77UVYellfFb3vGp
lZqaWFH4IH/ciALDAmlGOUs/sUTxrCxWS/TGofiwKAanIQdw5wTOCJoqVT0x7Nju3Ksald1CtAGS
9QNZOhmbyMnmzVgl6vMeDcpxJ9eRdXfGuf+rZSdo6wS7vAT9JDnGRedMDfxU34R3cVv5vmEkgVRl
H7YYmzZagCg7GXqvNfZXMg09nL72D/hYvqwSKoRFlGIa4BpuLmBZ9+dEFTkRYrlruR/LFiDDD4GT
aZ6AfHDmC9S7LF2eXQSjrH/P/8FXtQPn/9eAUswX5s33Kh6LqPRHHVrrsP3u76LDOdZB6pvoEsDW
kl3VamL8sC5Q1DMsSCcWJxwCUkxutMpjUrldRLgBTIKg3+ZTjgboazfUGCcbJM3XMHGj4kJO1AQ8
3Q8wPbxrkC0LB0fm/CtX1iq3wocFlh0YhW9tR+oPcRe8n4TQNdu2cYKBQRvBX/5b8aLdxMbgvnsq
YKwdoVqB8uQKKzQgDixFw7UGOedfMwtMieLMwmN77FznYOOM4QxgMmpIluxFq06BQ1Kz7MhR1Fs7
UFyuYeaJ6ryviQpvL2O0nRHK1s7Ig7X3lLlIdS2xzgqBEdaMfrmBxC1tHiUgDxTV1JBO65Yz9TnJ
L/RHhS7h9ZKrIzuXlqQ5l4upFjF3GmcUCft5r9l5G1SKK0ObMFX9MNSlTk2znZcumsC7Sk10sc6q
Z1lL6l1nPUBjtKo9NOdztwld/0R5XZSxfd80uKO2JBdzWLmUv67QldPz4vDObbknXCNbKKsljHWk
b7dY2WhfnmgF1flT/IL/E6UoykC1PMt+XHlQ7hWQiNyXys7YyQniuPsUcIzXo1YC7he45nUknaOS
DpV2bFMprcKHxQtaiXhSkkaYY61y/VEqVpQiUSHKHDcAmRev72jgfzbZYcKxQAuINSlAdZH4E5r1
lTpr/slrl8gdjadVQZggt+S3bDME7M2iRV9orn08K8fjuzML/+Ee8wmKhJ4iTy5vLBAHwN5BVW2V
bKyF/JpN76KnQIyN+6asazZEOfx7nA6s3f0gGah7wi7MDe2lD08BEp6L9cfEhbcvqE7mym4QWCG1
30a5JNXaSMiouDpP76xp5pFgzgzwA+U57f2FkgUe2BLK6ftQ7V829oo7Dk1Qt07hgC6Bq9F8/SVB
2UK79mwWTqTYqM6qVB5XZFv9lhw4BzWw42PJtfZngNMM7l3iQOosCprlBP7D6AmTrAGKwSqUUS5m
oqnEaBI1muSVM+StFHPYzg6QE/do76EbZY5yVFxxVIJ71gsk8P/f6g10Ojrbzqi6xNb/MRP83ZkL
YC7pbsn+uZyW0tG/cMk2mCQpnmX9SiF/mauhVcnYRYC86LAJ+7jsmmacXrzcBnF3mSUmVKTrcGDQ
s7McEB7dDGUpE3w724nI27v8VQ0hU0R88jU2CY4fkRrzLReiOqjBss/aJ7cED+Ed6t7FyIjHE3pW
ASUp7gm7Beul4Hrge2TAUlG8ts/tlCfRmPb7MkwoMLmttVAZHo+4B7VVC/Ha3d0hyW1HeFkwtrDO
eqEQQloP9mhSIptb0jfEj2n1t/RRQTJIIvMmto+ojrEG4rOTfUA+d2rmfi4pT/lAigvqdnh4d8xa
xdzPMgWbtUQS5uP1A48CAVcrWUj4zT6Nb4yiqduhJ4cjZ6EjJjTxYjOiJRsgXIYwCwiYAMrm1WFF
UwKOCqQx17F/PAiqKHhOyhqXlyczzVFmV1Z5DI9A4M3PYECML6mjqaGuK5M2OqAdcsI6ptr6znkP
S88PFnV/7Cajba/oJK0HxpONyZ3uc1odG81GW0sD9jbun+wvgmqcjSrXIwpjfe2R2Bcg1XsASLuH
JgV24SccYe7SwngCBfBwaFKFCYmjVjp8RtXmVOfnpx+R4+jxqyFKg6QD7LXmEfKVzlDDgxtI7Y9/
uXQxYRaVxSuk8sDU7qTJR3+co+EGg8IPU0WzwcVwMcaJuDlV4EBQgE6a7CHKa4n6leYrKKKKlsRJ
PxQnCUBXFYtAk51nfvafWTWIak/S0GSpv9yW8tDxsi+cQv7aRiYg2vRgrSIuBSbcARbasFSXvTJI
pwrs2yIkVZ2bJc3Fk6esQd/av1FzWqtPSI8vhxfy320bLupEa5OrDYaFy93eoRGqhKWJ6RWhQi74
GAXEJNsfGC79tZUvAohRSF0tM1umym6PqtycvO/3ZYCPEvYqcUV9afuW+4uKWNU37t6Ixj4X39X6
A2zr0p4vNlLChDZo00ad4j5HfaT61Ew4DU5KshTGFZfthsUyl8DDuMiLJIu78CXehEWkhgRMmCzU
Dn8gAx41ObHdLo2OXefbT7HLbIgabw8e1IZ32XOFxfhiGODHxECkQSmjNg8NqkOzjjTxzQYCyl+l
Q6WUOwtB4PwiLKe2/RdQD4LGNM1XHVXG88rzZqq3NI5tUE10ZIzzasYHlaUGY/kVZgXx5TvBuT4S
xrNni1FMtzcGuufHilyTndIZY4WsIhOYZwP6EPZd+9ypkObVIGBzViW5zZEW9HYyw0lvBdyR5FZh
lOxTeiVZJN2UobJKwamJSMoJwywTSjnn0MJ9XIOdoNkT5K9IMYCup5JKNhIqcGvYCf73zPhrxfRZ
WGcdAKuJ2Fjqb5I0hj5NyEdYe5sQJS5WVaOEpaAtrmmZcc9j+FWS0vVNS1eozEf9YAMOIV+HyAmS
h6yQT9g80ciD82q03wyPYFvJiUe4btpbWpUXOvGPnee2/rs8teXIoMyZwtM4rXL+VvhkSt0jRw/6
1SiNteGk2IZQzO1MUlwEC2ULIZ9jNYplAsBF2PDs/VVdu+yhgThq4v1zsfhwxUaNtxclN4rM50c+
MrBWN9QdOazMBy33Rv6V/veVMYFoSPawGnkHsFO0ibagZJdUzXhzF8nSEHTJajXad1S0efXiSOk0
lYLjlvJ1rvHGyyBhFjh6uyUchdqguNqz6WHvJbDJofuxsL/Hqg3+OS5TeO5CWMk5j5RpsiWVD/Qn
ODfulJMAqhP6ZRAaoBcv82LcWTiMfrSEpS9JByHYeRFVh0+8fsCXEluWGX7MlgGMSixpBBYj/O/S
dTTdClBobpMuJIumUXZpSbW+J+lWItgWtnaPP0BMmywGcbFaspSKB3H6Ol7m2Pr0oilUQVECkDuF
xKOoJNjoAdgzPS3vKmVdq2xybrrDUuoLU1cnYn2Hla4RO9hNwnX63AfwGirKjVRtMvMTISxff5Ik
GfD6Xa9JRJnMLJ/m7atoyDOmsp4iE4VcI307iRTxIk0kCmF8PCBbPYxC+y+EonLfu8TG3UWHjmcw
aWSzfmzVW6ZCYBTyiKbauv0mSkk9CrwtQScnKsk6TgXi1qKQPwuhhv897zmvqRvBk6m4vXKp5xdC
jS8cCTEF5dSR7n1MOdTounHBE9B99xA2ZkW1wCnodXefZ6WLHbCpUqdbfb6j9HiBOG7XJhrfslj7
tUx5V559IEEnkrAOv09oYOlj6bbItseDw02eqkxGJXqgnFBGS1u1C8OSmEfpxvO2jJ/k6q9eoMJT
aF1Bu9KCJRS7crbTp2Unkd9bII8+CwlEEzylizJyqDyaFxUY0S69oJZ0ihl6s15TzT+59Wj5TVdL
a94eB9Qo7TrfzTmq6mm+mowg2Zm6Mt0/THmoNIcQ86OH/AYOwPeElywVukiJxTyt0KFGT4DNLqjo
oUDLrdH2v2rw8KdIPoqg6wgg84IoSf09ZFrK6MXwFidO7dk+jzadgljBEaO0303pyzbVD4OR7d3w
dJ9IgcS0mGvlGP0Nbi3P3rZ1UkFq0SEQnNWQ0kML2gRxU0cE84a95qORik3GwJq6ycPCwk3rtJ1U
TAwJX3XEBRryrtccNkqVIcpI/Rq7jDoI/VmMOCC0BnA6XjhQVIQwp9blPHcNjtpI9akZLF5uxgiP
LkXZWmUn2OyvstmbfN1zwC8I+QXre1qC1X1Tw3Azk5jXuRF8eyaNrCz6Pk41iHO5v5ez5CvHPQ5f
yZDQmpZjc84TrE/gsvez15fIvI3LuOl60aUluOh36XskmgQnT+TGfI0cJtPNfOGicPxXNoxHCf0L
H1VxZ5YB4Sr3U0hoLZ4mqOyXX39IINFufy5Y9A6/9p2hs0R/QB3GcSO+slwP/8E2tcX2vrk2l3BA
HnxSnY4EWkd5ouxFOv/cZLzrmXefvAP6esSaD+Q5NtenzIZzZbTbQRd8tw32Vt/C8TKchlO/FsvP
mD03i3TCAtwB/rShMxmzbRanp3/BMXAQ8HGIH+8cSIo6PSt65s/3gBRsi+3ciTjV1btoq1UpoYhD
IdRFg4reioyQD5q6c+PiT8YllNEKNJ5Pb8im3L8gGZKaCHCDeILjWRO8NabQdfJta98pg7qlCeA8
hYKmh10CDd7yxjOyS24r9l1/EWDhDccm3M6HUOJLfXsW0xH9ay3nuoSb2gOLO9h3sIlKmHfKkyet
bRp5leo7vgT3TFwL6fuh7Ha9twhoSKqCXSCHEDASdMIsAKjaOJ106lIlqzopImOmNPPlykM9IL9e
tkSEQZuGKvbE6Il2I7x3J13Z8imCFOBWADKGsyCbTg2pS7rroCAzqaVjv1rvaBA05XKdw/Y5paOo
5nJe6yVYLROrG0G0NKWG7CtCh6YR+GcGjEb6j+iMKyuwJRF2iGX8v3UUp1Tk0LRw/3zREIljajDr
KYE3Un6nTQkgyzG3C61gSEHfAz2QGX8q875PkNCl5dj3HZtOlrWi9wbRs/uuKa1sbLjKcXGXr1SI
V4mCoqZ/ZvluPvpP2/08Eij5jjdUVK+I5GLNNL/MYXuKbb73Uw5kh2g5Tbvf295TsCOKfaNgZXFu
SRUiYpTwoGuP+HnbY5CtXLixYrV8AYmj7PEtUm71mY/hxDaHBvm7DkH8TRxdncRCRU4jvg0GTnG2
SZuefkwFCvyHaC3uRvF10swwAbx11i9x0ZeaoDbCcFq+bMPyiUHaQmvZiyk/fbmcG5CEZJJhC5a/
Ojenx9MDPh4rmQxlvBvhLIpy5HfDhRd8YPMxeqRaitmm9KAntYM84bpYh28jAIIVcA3C/Hlr083u
qShzq+iOmUYymdLPQzzLzYhDf5xlQrekTji9TSAe2BrDjeXvhb42DoXHGr/DfQB0SrZ2gArojypf
40Xv0UNcuojZefd7+BWB1v1lVPqxnPDzdTO0og0XJPr6rUCCrtKMi0uWme3QxirZ854mJ3RNQTAZ
KK1Mwn6KaJtJ2ozXyT+so0bVLYqVMTgj+F6oU3OhqeUPDMnjTEBw5Ve/iRz1+TlU6+n6xtYgy6NT
a0Eds74YxAeW7hdxS39ItytDVTGD2xGFLPQSUdF2t8WzcY0+wC7h9QuhIrHTP9SsMk5e5okdIhe4
jXgDA3KECVtIoNyzIl2RT/Yy6BdjUOjvQUV7LcaYZELkVyAYGdJ+c3JtIvBZkyM1NmIOyNgBiKtm
xyRcytImmJtJTuu2iM1HxEHBte9MbGrMBqxCbufkcwkx4JBYSahwpYC+QRDLyK2uATLRSwOvcshf
sYqH8PYKGuQ2uMtaJrKqF/wvww+E0JwQaig85t6e9XMUyjtZF5e0J8E+K3trUB2cclatjsmT5LZE
lyrTpMOjKomgooocHeWT3TCgehG020u/R/rN5qPkhv71CWspi8st+4xP/SiwdqyZpK4Y4sM4KNCM
zy0jExoLqE78ZzmjoyCnAVMwPvnH+EnOTu50+fSzeCKOo1igdrytcvA0l9tqjxm2scMfQrFP+d0l
Qhsf4iE/hAsDFyOjrHBp3UCvc6LdUjyXf20p6TA6iXo2LcBso7uW6O23a7EanMI0p3OZetbRM2/I
8Bum51iM/A7sFMRieoOTMocekbZG+sMa4mR1X2Tjz1H7KhdbGTmJzusCn4NNYa0d/R10bPv1gr2o
GgFgPp9XnnEvBpTLHkEjz2cXpFCff9Rey4371XrV/CqUmqh5T5+yNSAd+rEQjD2ubOfoVhHME9az
ZyII8Amzk/ZQJBiePJ6+Si4Hl5PHOkAN24gUG2QLm+n7WQBFZwed3zC0qzHJBGiD2HO9iVMjpKYO
XQ4QxPDGLCS6hla0H+twjxWY+VTRplA93yxvaHba7ILdYASRg3MZNUCcWZ3wmYZRaK7txeW//KJ5
zTVDidGxppnswmCe6zvY8jV2cORmi0WsME/o0GzSAyALL9vpwmGIatDQf/lMVJmUa+qTkVk6l+Cg
Y2UkorGyh8BaxA7SochaY1xBKWbQCsC7aLTlvkCZMhhOoDFmJBCOZj/7hrXs9KXBTbw8inYtPGNE
WgGfGF1lwVIBwySh3b1ddSxa7421XtCKlRbYRLxJ/tOB8T8fvP3BSmKyY01ws1E1YPzAnIKbpVK6
wqHroTcSX5j8Pw3eatg6cb9+U89IrhiEkcWA8Uirp/pTXZaM2T4uqm6A9kV0/grx+X+t+B0Ht7oe
TfMe9ZHb6Wp6SA+gVgIQUOsrkpj75GPJawqgbLDQ2RHy3vx4/kbCbbhYc8Kux9Nl9gIN4PrImAKH
rQudtkUnOxi3dBOwXmCCpVSqXQjKa04whpGO9NhzVOxYDeOFxR0iNmoIFOJO8c418BYnmZfQvqZU
nJ35XC8u1s9mPu6YByBYNscAGGvqlOGafMLFnlXsqpAX2laEH+bZ4QHMUzyV8HAv8z4tS64+4yC1
sNdzjSoIxihzjwSDRMj1nVIZAdPmR/PpqjjnoD5TKoESbi9cbz5u06go3tvjj0qf8K4Zk1NE2rrC
u1rtkh3HHO+X0v4pVqiwnMjkbz2LPySqQYEoOa9gr9/uXAgXBfBKhRVmYfWOwx941V/aZvE+BWGc
7CWmHYULJSuZyT81ERpoyzTpN8bgec+E/n5vU+dXXQWvvBdnoIdpenfN3DN1gEKMN3686WoLonp8
DIhQXwyR8chShdX0iF7tqhqXWxRQ1h2bz+vjg37OJMS1rK7t3aFsH9htzYG6P1e8bg44BmOmTShj
4jkFQLmasAbqR+kMFSeLihgEf5jgRcCRGxSDoeDYuVSO1bjH65aMxQb0nCSnbnXQNd5ffat5qYNn
He4zezGAag9v71+TOmAtTmJC0emvVMHwAn2hEBWTgpmaPimDZHECjWD6lfS2XnC1y+fekXUWK7w8
H1sA87x9lb1edfTZxs0YmBjm7W7wVRcJqmaEO8ekHEFNc8lC02oL1nRXPQUJcTSgijx8gTsrqSNs
V+lMO6c8coLMY41SN4WIkgMesjoET7k3dUILKD8scsSyvkEvdrO18qfL0uyu53mpR/RGz29WbARA
IT8NXKRN6giLJUPeiW4SI0OcIik1fQcvS2ZRfRp38VFJwz2e/i1pREQSjn/yVIhTEp0KEsyGNoYp
btBGdQHeezAeCDLHtwO0plen6S+bWUtgNp0hFG1UOcQrBNHQDR+9VPv6kPODY+5XVUV/CxEncElV
40PsN4cIc28ceX3YoYzLogztTlnhqRAHnUBGaJhr4IsxDfg+ph8rxvnWAIXkEipzcCqiCbmbQABe
AMkt90bImfJVO2iTNIAizC0S17pP6DKpKw7idp+thSKk8l2CVp3t72ewD7HsJwlzLnV1dXZaAwnK
9SkoiQjQfQ4kOdtqZ3bfw7dKjp+ndlbXmaUM9/rIDZe/QQvlksmHSFnUbAjbiywpk9o3DUF2KkBs
thxVW/Zc2WzOBQYU2gxfHAlMuZuxRebUzEImclzcRGwQfLKoE1z5QkQMPUbP+0UeQ6NyrSkLr12b
EFVf1HYn9xrxV2HB24GkDPi2elRWUiOjE4kuzgTJY3xFFAabbuVq3F8oOjnHVmeUTjvWHoIqHRN8
hVq5p9LJYc+ME0nn4ztGaCgiII8TVvhCUOBmH0hrL4LtGiwQOSSoEMx9XPtdYnQQmbPLIwyvw06+
rT80E4Z/mlkV7C3gVn0hjLuUKf8HXLy6OBD3JBU9e0gh6yipnP3BUqXKOstlA/P4Rs8FJglEIW2w
1YsJ5hSIetU1k1HiagYLHtz3EStcU+HOP3nAykJjq785cidCrUeExGnoOwaoUQlxiChPNJ5wk/oF
jTkCZHe90GiR7gfz17dsPYUItRCHyq7c1RO7rAvRTVkyatxktdWMoMZmnTuJIwjfFimNFQ4evpDs
MSv+9s4zH3+vKN7P0Sj4aGhKTjJiLyD3kg1d+vGv8KgBmZGPvWiE2PHZqhXcsuBFA16gJY8U5cK3
TBAtfUfaGQnkkeyicQc2ayz3CjnwnGDclXr9GbaEa4DsUWOZpuPI+qap90VULV6GssLqh/wN25iW
M+qQ3SNt5JXO9dEe0/CEkDusP+4eYraZGELew7xEpSg7QZh+TSndjpDMFGOEXXebYRjFzFff2iHo
mGahCW1NjO5jEVytescgr3tiszw/2JGHrO5K+8H+44+rUBG/kShNVSXsCgQxb7p1zmSY+yOoOiQN
hxrJtU1iiiH8/r2SKsLJ013TDcmCE9ryoRyh2+6eDZIOvbpSd0ubvxx6x+ZpxWmPBjMc9xqObvDN
AlUcgjFEJHkopt3p92ncUtX3ygFhLRVx1mODriNvtF/BHGzCCUuyEzYwbsVrQ4Ek0LkypE/f4wkM
d24Q7+BNWcOHQcYXmb9BCgpBfQc8YoGYgBfP4Tl6PIxxKHUsPoL72A6XWu74ML7oZ03LuGj4xKev
5/U67iZG1wwLgvTjv9JASOxchUGYP9jY2s1lJR9iN8g8AWszlwMKBjEOkCxcleLG/CGjHoJ6aFjn
6mDRLjLYIqpI7GmDmSGRmSVMweX1p/0Xq9xfK0cINa/WCUIEEJclQCGZ3m6Dn7EL1mSXsqSUpYKS
FQ3PgKqdIs9i3m9ICKxGC+HZZdX//dyUyKdS3ByQ6DNwNbU/cr2581F9DabXowLIlwXG/W6EJMdE
ubAq6JedjdxvLuSPgpj8bF3vLStjH27GC5dCi2WHSQx/T6t4J4tuBKjSJfVmGv3kkQ5ZsSITjkbD
BqGiK2l9UCa7tkz11GrSyG7o/D/nDAvi4SHPexj2Tzdk7SwjwxgeaULcSnHo4oi7ZtZxAKTmiUSL
13OGW9Wlo5rWlajNraJdB7Za+0rzFdfSh4Rubpx9t4wBZnh7PlA7mNvJjma6RBJWkkjen1S+0Lxm
mwDHIikKEMDYkUJpeSWi8F9GhDWmIt6uUYWnW3ET/9ytzKzyAS1QsPfWcxqLn+n+0ciL0Sed5cv5
ydkcf63StBo7dw6GjLtjmN0h4jozQ91m3W1sSQAKx/B8Jf8rYAf9OBjsEv1eG8BzcPlSokfSgUgR
eMjhX/zVQbSeB1L4/DwjyOXEcbJdfy1XhJ2z0aZ+DwwFYyuT0uXJlLmoYLTUf0aMS95WuaFdwYn7
/qjZH7bl0ndyKNJiiyYlNMYmhf07aMYQFqSuFsjzcobmkviQ4HFeR55W5pB5oVqUvuIjUfdXyuKc
1rozZ2SMuALVWouj6VcThToma8aJDE8lPcIefnj2LM1oauNxCKoTGfjr2Ev8xgOHMVsiaE6PyJbW
OuLaKgcyEyOf/6LNVpZoCnjs5hO+7zslo5+QIlPN+yQISkSf48nZyAa8fZA5TWAzm8Of64/Sr2y6
hpPuPbR8rcwoxmPdVTXbmErRgZKN448ksnWpgp7VZXN66U6d4yA00Hl9/spJkKsmn/YvGdFCRuj0
nAQqoQ6Bdt7dcDHmU+dFCqxesXJEy0k78xKVh2C+cWrBTmS9yxzi6mgbzTnY0UV7xQrPaW+I2K9k
j8g08ns+H6ThmlWCYDigoJmSQJuOOJ7p6nksLaKSSzBSk3a8OMGWboxOtfv7Fl/2cjNCG18+7gkT
8+Pg/RZc++okJAzoocWKM+xpatwNFeV4dMNZW6hnHM9hpgHAyzXq+E2m+0Q407inpgWi9/L2I6jV
EFkN6GNDBY1OG6yx31+Pc16T/VEjVyyVi7BSyXZodILrvED38Tht5L/+Torhn+Uwne6EdyaVTilP
mFS8ADjnMa9LwJvxvSvZPTfdXMu1Svsya11HBmQK4oHJ+6dKBa6ZOWYlUbl3iowj+vpRtZ2jnA5b
A4mwu730cfS2GEErDmA9drb3knmXXYdJ1azi1KWlWXOy7Axb5UiLV4iCOOFXXv4IHzJsr/MUIcye
AuTahVki+ZwzpjVNXWsIpAddST8hu1cqJV8UKYRg7o+jQ82tR1ekukqLMFtl73Pk/ByDZ61OAK4Y
75tzii/hN9xPeY6Acezta1iDqZeVLbPA5v07oZtuWusA/3PTbiYcVEvsUwVF+hMVxlCf3cV0vfkL
agQNDA577JGNVf2kmM67ACJ+iWkm3icrAUhisyk5REOcEFuMWCNFnMUdpC43qXp1dJB1L+p8YMVW
TuD+w/IihvWq/dr+uZOqaqGMBsSCbLf00UHfFbfrb/g4mmAt1sLdzC/tsFoycJGnNCwxlpSwvQmQ
UMOEIdZMKuVWBdl5L2iZyw41FyIHVP26PPT8d2kCk+jPTNAfDeN6T09Wi64qV8o/pUhucsCmT1k5
bcjY4KzlHa4cyLvHTwI8H72Hs3HntDz6zzoj94jF0cx6hfMudfDVffiAfjC3emEZDbWI2ffGXW2N
gMM+qOfnGYGz30BDbxGvjjh7Es4lngWhmri4qbHM0zL5k/XxUtS3PT0SDu05zApYFblLY9iypy6B
rwFL6bP1IPekzxLnmwINxHJWyAlE9mGrkQj7V5YCvunr94roQXQ03asbvWesWkgsnihmkYz7xnIK
Bx2UMgAtKrPqWBhhehnU9fDa/oVfxehm89VjLNXrOJcTgpuOxNBBW+5MP1pVOLFlil9mEZg7tx7r
m1hVgEVKPKt6M3qKHGCgzZGC6qta0El1h104mnS6uJiRVLGo3MxZ/rODmoyxlHefjgqNuFiZvVuq
wcmRmMhR9e3pV7IkDGFGQQj/prWd32vLp4cGBp3Oyd813xtLDk/SRKphm+Y/g2gNtPU4ORQ/OVXd
vO+jdRrM9EV9W0MpzxsbKAPSj9T2CcVBmrbNDlizsuWu3YIY7Rrh9tCPh7XCk4BQUDnetvx8LAY0
Ala1O0i04Ovwc64jKq9tadt5wNm3EnNdcfoKZGRea2Twl/yrWVy9DQZbRWHZJoLy8c/jrDmr0L2F
A6WILHi6XCJOkfYXLqGjxxzmjuIPWBSSAI7RukrycGbZIYg6XFjiNlGCNxh6aDt4je1rOhZev11U
GyTpW+P4cQ0CC7JRjQYd42UlRZCQC6w3Fd5oTQOI8bW+BDRLl3b+NiQz5Fw5QaZK9THsXfghuevs
Hw3pAVu5d9rfp9a/xDyWso7gMsJZs6OZPV7dZxljrc7EstE/vJ2os/BI+2jNjyxv71wvclUWz4Mz
bLpiDy3kbrEWA6xAFPNTmiD4XX425eogwAE86lxzpjBWhv0Mk7hthWnXmCPO+i77RFYaoQd3VMBi
RK9ahBkVALEdOVPYsqH+oWkuTH9UmKNtMvmgh6JITw0b32E5SEN+wb2sl48wz9Quu0fwb9noXGXf
Qr6NltdQ+D0KQ/f6Lj1kk14cCj3JXuXV0t2UWsKKIGPUdGAE5tCizU55KEOAyQ5YTTg6KEwKcGQB
8tLACNy0BxlP2vFUlKB55fo6vyiLJY8g/wk29Ylixld2iBWDnwNt87q0nOUxnsjT75EC9Rwns1m0
0zemC4tcAfVsIlHvcuGrJUp0jPHluEN3X2MsdCm30l4GJ+K7ZS2KzIGrY+Z9UXaxnx3Cy7f5oh6g
vy1IhNCuxugMnjUIhB1CGyv1ABVz5ZQxalK3jG26L5cazTgEdraodhu5P3ZtmCvoMMExNvJX/ULg
QyLtdLT94YyZgtIX8v7uHDv4RMo7zPzulWK1jXjzEWCDcnjbN7OZPJlq/pABz/LIQh1zhhO99lCT
X2aqkwW1ZHl8ApfvVvYPMCnjp+Ji3czJThK2Q1LBrDNfa2SsN6bWXPq1C5xkIrOBpfVLE+9VYy2M
n/V3cuhiHoHdt/uKY/gRR5mgzl8dzvvYqpnqsCfThpDVa0uBuRlHnHq9SOBvD2Ziox3QJ2imjmOI
f5OFhR+vuv4lSr+Xdf1x5DpkTOYkwV4gwiMv2d2SRr27/RFgzrsmt+GddVjyQ9kMHIOqXeuh3QWS
e5GhYB7Nf0P6wy/6ZKTA4mDTLvR6OdN1vy3XtQOzHAbMEmLajbjoJTlNzY7uQ1K44hZCHoix5gtj
zo5EFJPhKjzVif7zDWmHdz47haRCEldhLARrjgab925FCqsypccY8ZnQLLm1OgBS22JUT4j8fynS
NALUBiruOrDGfWy1iEMSQ+PsuUf2+rPDboXF4lUgscHEWkunIqvk9YlayA7fMV9xdMu4XsPRqyUB
5DucqS97TX1MsPQNX2MtUij4NkmwbbsWG83P6UxXzs7/KiQPtiKoTk2QcP3lZuoXzGZnwW5Vr1Ni
N1uDVEUfdiRr28tpj+PJo8wPOdnBJesIJuZbqC8Z0kJFZTe7k2EjXyypEoIQojfMciTd209s9D1p
HhySt3D0iYI56I5YxEFXucm/IXnZzxptlBaI/CmgRoJIxXYsTVcwogRkMR9OCJu9P/UgXR0HqxIO
Rfk+VmgUAyb7eU30huvAmGSLHOX/2QyCZ932rcgpYvzIG8W7qE98fNwaNwUA1DfTGYEkZqbe0VZy
hKMupkMOgbiyPPGBd+MTlCKKZlimyPdlYtCl9fWXnGZFMd+15PczOXMTqB787IL3vqnwuYew1U70
k49jRshejnGJcB6rvgRhJHWHoxZo7tZZwhmRGM+I2t71o6+/o8k4rOoucK4m6zWHl+VbpZDwgg0C
blj2wsHcWvQvm/acoq9MhQykyw3XTiuhituRNnWQHwJfmp2ewyTWZeYgkKOMtS1KhaBeWarc0y7W
FtJyR2j81kFhxrADhK/JdW08AHTN7Q+0yUFYYnOIhpDYFL5VDa+7KnKmtRBrv7bueqEsrpI8CPEB
nUrUiq+D5t79bNtdmoqYGz0Mho0BrUKIJkQxOvmYPG5N2sSCxGUgZksSG/HJgaCt/Nukgcf7oZBR
OP7Xjfa+GHvS7oFpGmqWUyUAYu2hsmGUL+4ZJiqNKNjvoQYvGIs60Mm4oloOriF2adlJDuGqkHtL
Flr+QFa1LCPRFXZ/eBDCg0m+ClgVzDU9X+3zD6N+BAPWGe3jqpCEuwJT1k5tyqd1UGcuh4/ut0Op
/4vXzMpiiEGCeqrgIbCi+S1ctdksDFAAJASlhgCIdkWzrFOh/I04A2QbLLsNo0tVkuXsZ5LbNnPd
OhtuTRW4uNk0Id6LXNJvSDF7eYzYBXJb7Gn2eKqZQjDEPonfyj2L9dacHDTHBAXG8vyqsDAat9Rp
MfUEvZmUUP6NqGXJEFVhr4GAqzYVeH4OBvkgq8UI/ECEfx+hJU/5Da1fLvrsY6F0E9JqcaChuLX+
F5yK+pH1WGBuiZfaREUdOlwhiXWjVc6L3COoX9ngrQX2Q7rtHZNdRHb/HTGr1qist0oFu6H1DXge
STJwfiuz1XldNIN5YKQharuAQqbUQex8ALgv0y3ilHKuAX4c+jh2sAjYRakOTl2GZ5fkAW7VqXoW
Ex59uq99uVHq0GJFDSPr+8h05qLKLJ1jwOzu7oq353EG91H2Ri+lM3CUoSs4z1SGVLdI/ZT++vgq
hJSaKJjf03jkT5sRh8xQqsPioJPLOsrMk57IWDu5/Mn7ATz3A6elFQ0IRj7u6GJ7XayNnppcJVXE
s6/KXTPuhurpQzkiC3o14sM+zczKjLBrF2P+X4+fvwQW0FO97XbrWyIYetaKfrGnaN0BU1NxxQUX
rGAyJJW8wdq1Tp6gATVgRGNjoY/BkFQ/nUhSJJEBlVnb0os4EdoPj7C+0Vz6+H7TUrLvlxpTllJX
GLCheI6DK6lPf8yWkv159alJh+KYOvJKcsE3Iq+melLR6SlppNLDqDHKiHoG1aTAUiENAHtTE1Wd
VOSNUOjHz0IrXglePA5KSMbEnWoPK9JTuYannhmur6W6xQciLPEGC5y2kxpEueMvmdnHAXwEQ2Vr
a4WFy3lPVsqO7bYfznv1FwC8qhIRXgxwtjODDY/a2pP16n/tRf62u79VzPMfm0azxRw0r167XacI
M1QdOr1vTIrOChH5nm1KppmVSS8vuKhdZOL12lTLDOKLXAyx+Iy2o2s4Mk5WEXDHwyiOu2xKbYQi
TVyVlkz03UF4rhdLbl22YjOJbm75hMhL7vXyNdj0zXqSz7DO/83AZU38dSSfnSYqBucvVAflMXcd
DIpvqkpsLWBQ37HlQ0pTMKSwRV7gaSA8nPdABr83gASSSoWN6i3rAPo0rz95zvDC8THqIEgMS+KZ
JbAxmqFZsmUhoKuy5TBSrwPCZefWAPrE4ZWYFCALGOXh7piuD3S/M64GeLxnSH71TjEqcLwy5Hti
WN3kYI2X6LBkYUubBuKnp9UeUcHayxYhNPGB2esC+fycSbVmtrK23pHoQPx5mtNajHn64DwIqTFB
+KYFYc5tAsJV5IWLyHo32vcwqjRkkv+NqdZqRvR9pCSSofl09aT0pHUN6/rUc3wMqetxg6CID518
qcCEdinhFU2NQmp8T1UN9vgrOQx53Dl1bNFa1JfwnUFAExl//Tn1txsDOUaRJ+pdjmfIisyaZu/f
lRwYeuOx2fc+zEgGsDng+c/USmhVstEXKR8l6RNFLhPhj9SMydqAtiN6ngEr0VB5qgtmVgn/dcF3
+nYH8h82OtfmaEyp+Gml2MwjBX5QGGMCjgENza1f+TMQqC4UeGvUqkTKBAajenocd1/j250da0Tc
9Dhs7b3gaBsoOQKfpfSPNjW7TpXGMll5A1Y8oBGer1QaPg3rraxrnkm4ubguWFHj/NKlVWkuG2Pk
JninTJbARsnpBG+Cp4lr1o8CL4YlAt0s5WvsIGy4SiOX9fypxKWQdv2jerkwKDzjmwVDvG2FYnMv
grWsbcBrNaeAFGaB2wT9U6AZLVhDwNkoeq+4Mrw4jT6scg1Ea790DEVzgtcCR6wFlOurprAHeheX
UVgTZNOBNSW1kTz5ewOGT5wQPAJ9xeQCjhABLZTAE04e5iicSBji5nWAt48EzzP7Cq8Q7FG1S3uA
/LJ+fGYFXOYovpzYlKh/Nnb47FK0PVd+G0rPOrohMRwD+BGRgUV5JV/p7mlS4vUPe17tMdHKef2Q
zR5SAyMD6QghLvEBAsTRNiKavWYMFvG8/fdU6b/+2OAILLoYDWXMCF9ie5wD+5Oog/eyDJLE6nVC
/N+28D+LErWeH7e7ZquFwCuqWFLWAZQfsmwKiumoyUAqwU0O5yBfD5JlPNOFna0qfXEWXaoyAXKW
h3QJT2YHlHcvllZmlzTYdjJ+pDNmhvjtD0d0wNmhNPsre/YOyqnXBpndq1xZdzjhIYbw32YHmLLQ
UrSMAp1pGnKJHgnbkOpHUgWmV/xBVk8JqFiWtiQOILOQULJRMT0uTDxFrfAh6+IPCzgqrxOkPh1r
Zp8OMEvtOHm2YGPnD8mX150qwUbecxo8mFSoSR6Me+mW6HohbHLnx8+G4vl4jZXVkEz3SBdTTb1u
XALBb3feA7RuOWpUXAfs77QeegFmPhHUkxwVwEoWJRyjCixllcjy6HgOYoJqleNHPJDDxYO9+sx8
uaV/X5tgLPHqaUxRKEebIlaJKSt4T7H1ppVKBdkeGe7R3vZX6jL5WoPlmfUBg9e8o9Lnwq86kXHp
t10qSxMfQ6I2Iallt8+rviYesBvxbdRfcGsHufoMQ4s+HmNPFUU9a2M4um8yEfW5umVaKSsrsmSh
OuDYOR97L8rdKJtedF5gZqOgIyorIszv1J1RFIL+RB4iZufpKjyE/59uCcO8XBPGUR+ZzibGck0A
wv8h/8GJI7yMsmFL6Of0yJmh9J6atXhW14CwUUHyekH4iUueEiedSqLcx1kaiQUC61BF7GgfHEws
wJ7lA2YJSm3b7mUESmisWF7Cw1hIWH+LM/D+wbrFrH0nmge5IsJLezqCH6uovTaf9NT/UtcYsvNJ
/wx6EzuXjkc52egwSl0WOLoDOBss2cafG0g1D1zjyepvgitoyYUgZ6/s2hiIV1tJiT6I1cMAWue8
9K6+KNfLV2WKkpqgOnOVgx0HuRg2s4m4eRfEtAcse6LM/B/3Ihm11iNTE5up0BFC6enXxWWN+Ixy
xiSI2svgG/GGA4qpvAtZ0BrfCZvGsvyB/Bky9OABfDPkqovumv97r2g3+nOkz4JmRv1PxFHYnIKc
YYa75wbM+ql/BPpGIpYP/xFGrEDXti3hxfxvujf6+dnjwsb2ewzLefRK8Y8gxDeQsZU2N+mSEe7v
5hGqvuwEAqJ8UCZHqNwsOL+xC3FQE+/y0AAHnh7FHvV/Fx2ebudQ/beQXDj96AFwLGSDfN1uyVhX
J1+vkKK0mttKtmDBhiGPsEz1aHD1QcB0+1G7yHY52GDSayJYwXOQovnHnDMU/8boVQcT7gWXxg3h
YGQkGkk5v1k+cLV2S7fIMKc6PPV/BZJ+yYp1ftjcdj7SztcyX781Q1+hrlVgZ8NxMMPX2Mc2+EEB
F1yttoH4aOA9hHGthSmx9PnUMx7KEKCT+CKKbJSlB6kz7AHaIR0g/JFKX8iKYqDzXQEVARllD5bZ
4irrMz3ETBv2qsmqpd4sSwHd4E2vI4LRnwNCPQ42mHTd77LyN+VOtMqGYMUrfDVJRbuSGoL3PiJC
PddyOkDvBbgk/w5TdfijHzWre+a+tt5d/pbG9pHN8SoCnuK38dkDNA3sfZ7MYIMe9WAuTYxVf9AP
Dvk6lR19fVOuapg7NYHnFA8RBE4uhJmLAEsr5/zLLMhmFCGAqRY8zCBIc9sCR4U6ww/ZbTy7V864
RIPETpZosR83mZL6SkuQxUAu9d5H50DjREPTb/0Dt6bCqN/He/+NRxKLjbZnw0tAkEGcC0NB5sjV
JwOoYyBkShfF1BAYLoPagCh4nRtpmzdnjQiIoNRTP0dMTGLaWfa2BgB5qfUnfNeYL59Cd6OwCNGf
R9U/f4q/+6J9RUhQ9I/R8r/SRBSqBe2Z7/2q/gHuiznvlvA2pBjOA0LvItXYyBo5rKE2s4qvB4Fr
N1pCZAq1kW8N+RR8fNLf+JBYP105TjBRGDDax1pdQdYC55frGqmiWyfl+rJzYHuSG6NZ8nsxhIlX
tLW4rFsQlqJ+GaCWRUYHGsmAjUKXo698oSxJs+1rmdeRYkItqRrASGJNQrZ7SGgKoPS5wNFbLcn3
NMZqP1FJ1xLIolOzFDRK9MfRWTxtRkFZAufuXK/tBMb4vPeZEYuUKB5qSyrASf9/sx2zZaGMO5O9
s3GIvFIdWjrudxLB9Ogk100TBpOlzlp7k8b+Ja9OxEwnlCxUgjmTmdTJ7AWJ2haKIoES5+/cIpcX
skVt0N2nJX7mGdcrfPEOIS5X2gQZdSQUwur+VHLyuyaW/3dhQeX8vI09t9wwmFRtlUMg7Wr9X7dR
hmQ6S1L/kLPwUqpub2J20AYI28dzNm2pPOxDmAbM1AmaNx3x+1H2+8EyDuCmpfczv46AJdeA7iwI
K9Xk76qKP+SXQbDAfgjgxWnCIyR+aXcK6myJ6BSoXXkaFtNwnnmWII6X7FBN1jUON7aoOMU9JewY
0utfSYGkdtm0Re55vADqWXDqKRAAIifCWJqMX50TSkwh0t3il6/8E/9ngCHNRk35nNrkEz9rAMiM
ReFAx99uux4fHarqAVmWgbnPsr7UiygTXYmI7M22/RLtBp6fgZWdtgf+1En5/SdBu8M9T0MoYTBv
Pk7+kfpdfvgWH0mMy3S+DPvv0AHHLJKDOSDXBU/+5LToLWbcqIyn5YWdt4r6VM1q01wVrxxouRXA
i31yU7LaKSTq9L7PU8C+9Ol60U/jm6GMb38n4ukm2UKd7CvuAwrn2VirtfjygGwMVjg3UtJq1kIk
bQi3sGf2fDAEZiWS26FfN5Ad75i2sMyYzV9lZFpn74dNhiKb7s4wlI0o9UwdBbrfLWQOQ+3oLLTO
S3GPdIY/2l4bgJhX5qIx+n1/tYEzWZnBp/GaTbtxWuirdULQ/Qglosfh/uQGkKeVvGu/kmDSUcRV
ttnRhx0c5oPzOHzYyVKN4R7KaUE6GWUDP1M3MNttKix+ZovKA8wzd9DELeUbeNzCu0kgSUc8qE4Z
lTO74Of+p4KHxSEQ05VB7g9CHJvuLGMXtd33lzwLk6bSjNVPDDcIhwVH+HPG8uk50BXu04N756GX
6mcEYJuAYBAuwakcsT9036Bbdx3fMaBnnph/ES5QUMBPaOC5Ps/OgwEYWhZRE1d4MqgQ229nqsyy
bm1y36QZghBHprVQ/9hW7wXlb5Fb/52qUpXK1T1cdB5dlZ6EKLvOT9K7Q2lYXUY6y5uXbfqQYpKU
sY7jZDFVmTkqXMVew3O5Ty9DISNmvkkS1c+ObHjYNZaLve9fbARsyiI309fM6coD3KuwOKW8COjQ
nNHdvzSL9ZL/IzVh33IAYg95oalbTFDJVdHEizNXqUamzQK8jCKOCoM5Je4T5uWarHNRV8YEZ57X
Nb5OW0HhFxtGoPCMTWuro8TdJH1TR3bEaPiAwCDTffSTTsz0BNYglqZfJdJc6q88O7ZAZguYqSh4
AjWA9l/lhdqMqYvLKnQtuh92MQQy3zQHugjygE7/lK5vY888/l8C2ZntFvEi/Cy9y2qWk0Ct3pth
Taj4VysBDRCtS2gopMpFXPSBULOo7X0dXJ40KEtifOo5/AkyXfTz+QPQo++T0Qksd95JxGUvMw1X
n28J+qMHGQFw8xx9K7PhSgE8QBJcoKBZfEmZfoio7a3LAL9mDpFxocexe3zBi4fMRLcSMAZ2e7Iz
tD7dev9XV90LZ+9w5F/QCf3bX/DpjSJNpFIQDOM22ebrwEphKUHjsR7TxyqhNP8ShR5C/eo8dyEh
Xz3BXLU8U3nXgVsoqw2ypmbkYiFjbdUFcJ+mb5pR4bvD5GKQ9k38rvTAm1jg4FPGKbGjmK0HbN7D
F8dMJYG1XU5V2prlAcmxgCVMU5OSRET6wPHUsAOt1uCTelUZHOLsGaTRm8uzTUYqmMAjn6j025+N
gfJK58p87m5hx4kcRGKgIwmocyyLnkwcTnfkuRzqv8IXZniuuEKBVOJ6e7G/53j6Z9vv6G1tyXBd
Vamo6X28+pJniPDQrycTGLZmpMaHAq0n7n5HxeT8diob2jTKfFgpNGPzap2wp2dKjyerQtKhy097
sE6d/yaaL5qtvRE7x2eSDEq8VIddviAT5TSv3n9NjnO0+OoMaN1/cwEZ+UZz5QrUdbNe+Jye654C
mNvNCgBUxM0FlBjAAfnJFq4/hZYKbZsCxSJunePPwZkACVgvaM2A6dX8oo7mN2LzquGXswWFT25X
c1tFVj+tf+yOJhwYlkH/XuGmMTwqx7p1hZ/DI72s6eqjFv88SUT4Th7A/fhRSEbvHbiwf5+Ug7xv
qqRC0mR6xbkLCYynnIS/eaEG9r7sRsoTZbR/2GHgoYpTBST6hEAZ/9awFwkGrX1bi3AEl2gz+NuA
GnM5qI+dfkXgN9c9Iy+D/WU11S6qYXx5R0u/MgmprTM+ENcI0RjzjExtshJJVQDqcxG9D0UDeD+r
z/MRuFm7wUPI1UVZL46HiBbvg83j0fCoyE8/I/+ehbxst/wg+J0IABNarnvsPnjl9B+ZIVFmwcXS
H3gbolRS/e21QMKMT4sBxIP8tYw0UKH+8B7Wt4u1x0fCX2xtC1EYWvfXJjXPUaFLX6J8xRZdsfu3
8QZIm/mNO3hG2FHvZeFxxZWQY2LWbi7opyMDYIjqxjuLeBToCa7ZSIn5G8auP6vqppylSJx2np+a
8s2JjcxNZVdnp+q7VWcHRM/yZ0lgrn1+8eFy0CgL0n0d2fokaqRIBnDywC3+E7NJaGQnCvGcOfVw
5AEcEHK41UF3mvDzkAncADvg+2vGKSwJKwzZvo06+UrIpaoLEE0pVgx+xT3pVzQwTNSMbLITyjeo
lOtQTcwFonXQhHv2/lwenD7qJQfGxLO85gq0fDYWc4jD6ACV3sp+pRRint1NbZplA4GgXxv8logP
EoSt1u6vcnP6WIvhMntNxt4gmOb1+Cyz2Zv7GkI7ILFaJFqt41m0BAU1b1Oxw1HtL6Fs6jcpr3Oy
rUObFtvoixE4koeFhTXA5riz3k3i9iQ9uDyaElI0S2EJBGXnUxC+OSd7jrvjIQiGyJShykUZrZMI
5N22U+YfY04EPOv0CfHsPdywOYo7t+JJNg3y6dlHcg490RU7lw4O1JHWAkn8a1izX9T0CYPR7Ork
pyn0DiZgnlqyQ6bYLln8UQ6wGzwpTR8oBYfrAt2ngnXYb6BTZnhY4bF4A792hQSvK5HT0cnbmpwI
9dVjQAGRHpDcsJgvN4ZeHSQZ8pdMKW2uPLakfAPbJ+JKe+VQsb0LuWVlQLysVv4i8yY2OetfwZ+v
3MPD8XohcHHxLSNKH8TCldj3b4Z/EmGbo4O66C274rODNvEkISztu0ooukEzvCn+oecjHozQNmgG
ayAffkfRpKZAD0aHSzSnnSf5a2Dk7WkcpO0Kh36++KozIxfcgVG+SiW/bzK2DIAQZhv/8K0JrFW5
f0LJjIlA6Sr6Gnwjhqw7LxuuVXqpUk0ClOrEhYRDx5+Ok3FJL+aUYXBv6eObPnD4iIn2unYRZ4mb
jvFFh4oqZp5UCPryE1/AwvH6gtB9N4ZWXiURcxTrAJTixwN8diMC3yjIbfwrQLns8xQwho5XOsWj
7ydOz7QS1cUqBRyNUsIV+ULjziQF2KbSVVX+zYYsaR7NS+FKwQ/PgmL6Hvzw6l+FWNz7OGHTqkXy
Y6PSazs4mfL3gRVu272Z6v/CLHWK7RXkNEAvG+10rn5wbsAMeTiJWWkczYeRPygByLe8C3btHNK5
75fD+adUnXBG/U2EJN3zVKZ1q9Isoqz9VOicLKEigAMv4leGyWbl0TLucfTz4v4lZJL0NV7UR5Cs
uo5NbVRBpQxmksoVQqGT7oPehYCeoTUE7XzOQNILMBHYvv4kAGt3Z1Wl64VdRyeYZD1Dov8BxH/6
xlQWFR0ICgFJdoJ0CoFKGE9kQTaU0MzX9FJkqhSxG3f/WVTb1McxBq59IcyZfjGGukXoXYKwwTJp
DfPK8EIMzYNmdcaSUTj+9krr/p3H9LyIjRQc2p0vdYRX/s4SGT/Q7iYrqoTxbEeb7RcEPHagvsxC
DPR7iuwrkMpx8pCb/jHdA0H4fD0PaU1VOmIBQNpGWB3gBYOiEoDR38JTxmyXk24+JNAc+qttLKZZ
fXwdwNU7rsxLvcZvyliw9qyhRI8acWY5Z2crvPn3GTC9oKawnZQbLMuLqNDpCv4v2/4Mwizdb2L1
pT0yAe1SRydFVkSmKNyPWHrZV6bpzyMMxlgLA2Q/QxZfzfleimjYjUnwhx7ZOdNTYuWvl5uKTY76
5U4WsbBj7E1ytDItkx74M7zaOwXQgzvbprhRy50sAPO9w7p2P93PlUItRnp//HmmApgl1o+Xm/zW
gfi/aNlRnY7CPq/LIYcocyoeIYASHT/6hvizt3miLueh/2LlETzUX/1An+LHbwzPbTop22DpcpbN
MFV90El2viqTFA8ULPEGyQ5EllU6dX3pR/U5sq8DZf2SITDu6t6bbQU33A5KvE4XY1cTfoXFUMJF
a8gNVMtKQp3Vfmorxk2h4ToGJQVxHyPhQ7wDF1NwX+LzbEpMoH/j4lf/aAYsXoX1dAle7iE/ClWR
hYv6OsXcaBgw5GgARdiTg4lMI8cz8H/7Cp/oloOC5VZI673t+ymrmTUpvy8GGW4Mim3cd+0Yvpui
eFd12NR4ZuSAUFlcu4eEZUpNo5dQsGRnXzrSVcZoRpGBMzywqg9kYtnQrHVCG4BJZsqtQF/Wc7aH
aSqES3w8knz+wZ0gjgtWbS2z2POJtRX2yxiunHYLAAGSjHC7Ed2hlnx9hGy1OyxCCIrnJI7gtgdl
A33FXHWSkHyE3/2IwvdJrsnSwgmslZE/I59hFIFO7WnkD8+qSkLaNGU968lpq3QzJeD+yDPKMkUY
x7EEGzP06uARnx0d+E0rHqpAhclsSyQ3mwBy4ogKwDmXZAmNT2hF4B/v/aUK2yY7QFD6OEaK2ZVA
NsqS2Ha98D8rR9bt8Y8Ka95QvHN8b0ysHvOFnjMrkRuq4gxoWL2bOUr0fqIf5+Yi66a3JZkvdMqZ
P1hrMXGuG26G8PrG0drixF2KqC0HnRTXKPF0o1wL6JyQh6hJ4sdymG5v+KIRQ9NiLlbAeujkAiL2
GZU+5ivDPJFSbMQyhJZ5Vm4SQ5rwtPUpCC5uQZHfqu2lWEPyAoWkEy3I3BJxIEmGV6Po7tdnYgGz
IRMagDAw37I6yUbNHtxPSP27GbXReh/IDkjM2Mtkkq9tl6I8eS3QOMbXlvE2terEtkB2a9btDf0m
VbOEvcMlGhgO8Q4IiOdhbBC6e76Lf4U/Ci7E5YUOLDhsLZS4Nv0kCp5KRGjOV0Cq3hJApzcv14rr
nMQl0ejKoCZXIISnx8sAc4KnPX2FBg7vaLF1djmv7+95P1Ojob8WSNEXxRn8Cq/4umsVSCKSVqHx
8TygmetoKdPYZrNbwWsnfKtP0a5b4lNBdQLasYwUmLOwKxKGKy9W2HkMvQHygpFE11jXs5TqozFQ
2oxwx/M14Xdu3N+HFrYfBUmuFm7CzEvQKT0GgE7+f4myQ4O4Va1D2VnJY9fvD7K954qb3A9Kv0lK
0seIZPyZ3yWSn/mqjLVq7m0bF2qbQu8q10UYsJA0xWBsBXrUU/Me39/vM30kAbTYeJ2bK3849pCr
Gq+A5YzY0npHqmsSkfsmfHDmP9CI+CyufhN3dYsp+5D+vrzfHn+mSgdmuWf7K6s3OXmALHO6H80I
xrXTIDh48jtIt3Rw/9aMxCi5QXzxrAn821ypzfTaFZN7snTwAK3onWbcYiJP1DPmturiukXB69L8
lUFy1ezMtOxhfHI9JKD3E78+RiFaYdSuxjigJMJIJhLdvqtCG1bagwv6nqQlUAwBMJDKsTjDId8X
o/mIhGpL8kRasm0sHikL6VS2N3sd5HIgoYPwqyD3rStmGC89TGI+FJKBqLaTmcGx3QqN9PkW7PLb
5sY2EoekNyXkgGh3pncE0qPp/5sD/Y9b7nYUtlaHuw5NPY03lQ5JPY8Fz3eEGJyAD52SH9TBvmnC
elGBe4lZIBiIrsbyhstfOQU3nCtNabMDFcScm1rkbufxtoFfPh0eAGKo7fhum8NP8pG5KsoeNMjr
m2IhdhVrteo5K5z+6hw1Aq8jLtMZydWdx+yqG+FsopAkcrc2q5s69tp3+ZoiTg2uZIrW31GQtBEO
3ds+8kfoQqmmcIbbe472dHlEegdRMfu1W6aCy44XGhCs/KsCNGsaIh2taPZDN654E2fb5fPnbCeu
hCAS3Y2tLksCeRQUwk5hYu057x/V9QSipNSYl9oz9GenthUfH9LKTH309CcqOZ7Kd9E/J+pYmCzK
lts8h2rlvBPoibhE+YxDLDJX0ziNr5S203DjtGfiHIQTTgU1x0yqP7zBzy/FFP0j1vcjz0smO7/5
HoS6IaUjC+T5dC1eoeS2vho0M+XcTS7XVQVWGuT60LK06ky6Qi4QYczVo9Os2AJI49z4JPWiEZeX
tfLhAoS7Xfx2EfN13TTG/XJQ11UEAPdugG+vLRc3WWLIC28anfeADHKhlxMgGqUy6ubs3DdJj3Nd
B5nSpZlsEl3Kf8dmOc53Y045cRWM18FJfZ9p8Sqmifp4++YQEeerH5LCeUJPqj9mn59yYBbsgdQ8
TP+/Tr28aLhb8cU+RJ94gOoxyx0zpHwx4LwSbkVD++bY6kQ7y/TBjpLsG74t2DgEdY/h3LLA9lJL
oXIggUSMLyt+Dn42nMXTHPvwQnzqr/t2H+66WSEow1bCLMpovkVbqhAbmJOilX1lVI+ZR4IeY/Nn
1qpriJ0A6TBwAL0yJ8dbtKHzZB1KSCUD3C9hn+U35a0PLqBm/mT8CMZADpqoJWTRw2brPNGhA4z5
SJHa/kRkSOXNwuxzjGzPMe0AWJ+eXjpRxMOEl7iHgUGPzJW6qVbnqTTUFe+x09Ys60jsv8ItTyvx
DGBQLT/1PYBpELf1LXsvSNHR/HrH3HihUHBLFZJYEIfK9MBNxRUrDJW5HsonO63Xg/Af24e4/X5q
QYbi/b4o72NdfcnseXUG18JZVqdufmb4t5uhKj60gyY7Ia1UQUpqQwake0lbKduf4fviFxXcmgyA
srnd5h7r2fLl31per/UG3Ad/iFjdj4Xhro81khTENEMNGdk29xTIvZgWQ4bcRzf/eLtmmSOzYSwY
30IRJ5+J+qzZvPmhxxy0bq3guGnDS7laz8mpGD34M0mCP2YfBGiTDySutiPRyVyEdePj2TnvtyiR
yV5KsI0tcfSHIBehWtwOf3n+mmaE+HKpOYnt51iX2eBk9oAxDXPKp3hesRhI8iwP1jnIZJ2uzK9J
ghDnFLGKvrwwDCGsf6nwr0vUs/IRu68ivYddkEDScjNRjCiK+/ErQ5bMvh0dcrIeLkNM5Dl5Jr6U
1jcyIT4s8fWKr3OSTsOAoHlQGvvaWjwP/jvg1rdP7KLciVan8UW+NVOyPv01SOrAUFb3lt72ijVx
paC6iF+0umEZ/kl1AXZ6Xm3Nitfpu4mAhAeQ2NXKbe01Tq60BBjdgcZ67p82e15bbuZ2Bx7ZjWdH
hTrwDMd36VVNGH7lQ/X1QiPz+p0ws3Si4cRg4sVWkDd82PeqIiOs5EjtKE1mCtpiR5tbRCpSF6zq
MikZZx0Y2Ona2z7Ev1CUXwEgyvcL2j8XnymMoQ4zCU4khq7DUArdOvW6nX5zGjn005xXS9nd4NBX
RBL0Pgf6X9xE5/0oKLYRYMfryZIexYf4hX2fN9Ju6nG4FL1h659EdXL1jIJyZrtXzIOQ0YBzSmvM
754+b7qX+qbXCDGR5bQFjMJpkv4baJE2MwZtMbL2qA4BEEWvcEzttaeG2UA3UMqprftJv3D0M5vJ
FN77O1maLJiofsSVUCIelcIS6KDxXgtZ5nsEPRzBDS+u4qB21KUxhHRvYUgm2McKUki/vivlN70e
SJT03aFHNJW6Hs1wI4OdayhYQAyQfwjCpNCNkTWuHxIHPUZuW5QFaTvvXPZQ4YgmpUUgbSqSYlk1
azwQkLz9PnI2SC3J2iDV6JwkQheDUMJJblFrZXLo+JKjeUc8OSJJvp9HmYTo8ms2wAnQjwoMBZha
6+w35z+uz/mm4qO4lCwEM8FJwVSFQBBDxxN0x1m5RDpQPLkZ0VyS0X8jnI+hsM3hdCaJlQ3iNnDb
cExZylnUEuuto6BIFV5g/3ZEQpV4VyvS9iCbdrJesC2I8d61prKebaUsynMA9PsJe88PyauePi1A
1xSfZ+1RbPeTlaIIvmS9gIx77tkF6pJF0U38tMGBX5A6lekL8wuNeyCt/2fJZSaOgjsgaZVRsd+h
KF27zWacnMuUzbjm2YR6s4Gm7zXjRCB4JTUqc5hOqMvwGz7fK3SfzE+banS3axnfI/u0s3uI0m33
T2zevGG2LtK20AmG1WFkbLqN7woTvFx/7saPS7CrBKPHjgjx3R5xQ4UqBSX51UDockKPUS29qRPv
8W/3NCSkxgI+xMKK45bkXBvzQnVXBZuhCmDmbx/DQ3OasfUjfrzvet+DyJMFhVJtwifVhjrJEuj+
7HHU2ibDskzrIYBMg7cTz+Js+Wg520g9LysYocZJO/bQvQ+LbXKB2T8QcAGpcRMsR49Uubiz6Y10
jdtufScJ+RydeeEQKI02g+b/0H23DD3B92JNVPr0aAoIYDohF9lBlpqxTZDKCxs9ynrh3jEz5hme
59vwJLpvuyy3Jntya/xUxoKRwhC2L9QukKEG4PU65GlF9cncdzWxlt6CTIPp3e5b70ItJPPRf7JN
1pRSdhkocavYOafNAvKKoixoBhfzQTsR3XsDAIbhXuS+9uEkwugFiln2TlHWDLMjp6nZ7EQVUiu/
gCjiiOZcboVWxehCOzUr7Hdbj3zlx3qBlnbu3BDJSP7bidwS2TrF5WGJIq5mm0QAgznCxYOnOnZx
wF+VzyQqT6sP1MGeGkhxn1Bjdv1ngkpKN+F9wVPFw0jioq4Phnqh5Wf0RD97rWE66Y69rUfWATny
CqQ2U3fbOdeoY2uYkEYe29XEv9uCwEqkpMZ3fluGN3s4KM0yhKUO9P68VyefcKTLvlKOMdOgyXWf
GlVkNREcbqbejhRH4mc1oVTJ0mmkulTKJyIYuxTTONSN6VIN6dBqy+JsTBj0cjMNpSfYpxYmUdys
AP0Z36MRjF/bWPXg5TPCahVwHL0buzJpOj2Gj9ZPNnlXQNHvJsLRL5ZY6/xEfVtqHizpJ90ZrZfR
6QxJK9DuqSvBvdW5TFmsDxgDnBxddDnrjeGz5eHcj/YYV9sfr3ZxiYLHHBq6JlyNnrnCGENt3YXU
EtXCzMXErD9wB61Q8YdilMSRRq7154lIktiuJNETknR0j2te2Vu8YbUlDVQG0ty8Prfywx878b7M
2R5w0TpFZrWWrIQrOS3dR+Dxq4eUs5YteuDl1NnP7D4kG+sw+eOF8XfEy3c0ExDPvwXWMfmpxT/g
z8NxXVEE8hKVaQpJbukc006QQEC/ri3RjX6YLq+TEYcbcpXME41Gxc2A+JU8PGMFrgCdXUZdzEkG
2gVRJmJWb5HQfi1Bor7oPddbZcGHBilekg35tFnGDulGBu1r+gK9fGu+7tj+aL7W3xfC5T3VNErO
5CpfuCjiUDCDYrAPlNHmjQNzMeWPTJIndugH87o7YX2xoLmUzQozfv4ZIO021SUksgzjzznrejAq
o6I1TL7rQgIaAhJZDI9eAJSKHGJtm0jvmV9kqHoTX2EzhrS7S7YlK4yRbWsIbxcQNvv0SP/21UJv
yjeeFvGKiTVG3tayE4v808uEjidNpkpFwkzQ7spbvCGQbRXt3a9ZLpQzHsiZSu+2vahFOs+M5SCK
/nBr1JOduXPUkckLZab90XqIdv0Ulhszb10vIMyKBqOR4b02cIZUexBseT96lTfMOIKdh0iXDrnG
XnwBl3CWUNAvWQEvM0zJ+gtHhKSkkkzyFS4XI8HbdaYuEB+vBq/5Vsxo3AoLhoyD3GIcMfDpWYOW
KkfKezH/JhtopNsXofn5YeADiSVw7AKUrZbY3Vs6jtGsE0kaJl7ygbO1QZxD1DuQhH6WQAw9gxhV
WzYgjmLKbyl7e3FjL13qFYC7ZLm3/8lLy+9x5fvV5P8E9iYh3WnZEeC3zKE7oIKF2mhYPyzAP+g9
vgZj532oZiU5r1El4Q2ezy1yqv1CRamr/z1+ZQCYkpLFVmAPEC6ErWNcdTNjZPnXfyyaCSzgNJ/5
RssOvQEzlNmTUOLSwc2Hj3M9VITE7Ihq+VOG8A8B/dIiM6AObgJjZpww1AoTbae60+53vlEI1B6L
R4IbyCPt4Q7zNjM06mK8cqCtughoEQWQmQDJmCcCV26hUojX3xIYqHi23fSsjXKVaA0F9Zm7H9Os
WkdJIXfrDiqqBebOSEcOZtgUpNxwXC8JkUqvHL1vRycvEkStQLgsz41IHB0YWmV7n5llL0JFjmP+
+Z2zGEVOjKVq23tFVpRdJIcTEUDUrKMidYyu8oL3Pno9D8J/vUBC4tFkIxB2OwU79H9MpIYnyKd+
E0Z4mKXEfyXJBYzT20I3VZAdf7DwgnQO1bMvoAO01RKhqATgrwYf9/o1a/oZboNusrWhKnUm5aCt
4KZAPNsc5Cd1r571dkoTieA+hiPeKjb6AavhdVOu44u//RGk7Gq1P9AldHnmcqEIFgqxTlxCCOkL
feiPEvcw7/F7EWWViRgsQShhSnM1CBLRwMFBtf+ZuMkRsXcpOw/z3NDIYHXrrvuk7p3HG+oXGZd0
zBPGJSIKO/yLpXmcJ0Otl7bRTnNxPngb9C47tPhSAAEnpsldJIt/yyNTjT5B7b6knSGmnVsouLoC
nL4Zjrku38qItoZO9mzmtdpG8etDRzoCPAS2Yqcvh56K1CqN9qHIFO7sXSwIhtRckGHL10vWuWxh
D6fp5fPk/SL6pxVBfr4Kg4j7GWgnaCOLSKIc9nJvHe42oU+ltvwIBoiTvmINH4Rox+agbEIk+3p5
x3Rmv5JD3p43NpBBVfbz+oBOlnbTY+FIVaXkjpLo0WeCGIqz7g8A8+NOd36hVcWD8zfPNebszRwe
mHBFugsdq3nKbWDnWsvXUITQBWHNrFblnW/kRaVLFgsztnRUWl720Okpn1hDrRvHtLw5DTycoHj1
FO00xcFlHb47xoIHRPXwJv2nDRwHp9mGfatvNLkX9K8S6bXBiHldpR/8EmlP7QLIsvQmQpZdV1fu
hGjTKXkqcTQQFZ6s0R+iH7Q15x/CLwxynlgrJ5vi94iBx5kxZI2oDb+zgUy3mUfe2hm8EmhC8AKD
3C8Z+SPKFHUDkjnB853VK1ziWaPyANKIBXRZTpfYKrAAPu+JCPFnw9ysUJgBssW4i6d1OSlErUSB
ZmY69+/hXD3XGEdoMDc6l5dJXkhJIZvLtSIsrYkC4Kr3K41t2eDa5usPj6qzqJsn7XKOOKsOBfoP
kevu2YlO5U5J8Qb/9HMu4FRNNaJE/aORpNS+JBQ5Tx8WQ1WAIuLellW2wvQlVS6iFKXDNoB/fmOR
kRj8lILACoBUcJRdPBXpZV1CoHP6x2qcUlE+2nQTXMedq7pr93WI+Xf8UED/eRylXpXpct63rKuQ
9kshGS4TtHLSYQAcmUEbeKRBFaJqnRsy/Qr02bu+ltVr5+PtmhIxGmrqajPHrayAHkMO7F48D4Hl
Cma9WQhO4REP6C52bhF/4uqqaQ0QfyCL/AklzUD3gUcOHPfHUfGioGvecG2fEfELBFc0auxaO+TH
2g3QakvVkEcMRmuuxbaiEEbYrMag4ddpVxSE8LrRubPnTdBFPK+nL3gQQl2GTnG1yOhi4fA2HOyy
vSsiAiLHkipvZsWPOPmIVDdQGv5jiKKsmqS9mvdmqBOElT1KUsDcK2CMMSa4QeEA5PEgCA7YgKNc
ADnzfKRUsjKZHFVgVTTFP/dk/RoBT2qVl6CuV20wLyC9mvxLjgYjJXUrsLV1660pKbQ+WJqgc7j6
M0zY+URbYSMpnTrffwkdBvJXs/bxXL0K+3V/NMbEtsr0H9+KvCq1YbSX0Y7wdoO6oYHnbT3t6DWP
/YV2//T8yNFx/5UY98ibHAPTNOkpGGWfJXDpP1tsSBqnVtKVLDjNhwVND6n6wqCgfWVj42BlKcLd
W6nWIESGl5fMUrJW2EomIoaEOVtG5J+OtgYojyLh01URAKRyyvs59w1ZHF7AoNEpf2RrP8KzUPLd
oQKiUaWZLm8eWasTJiOidZAxHOE9fZr3rCZFTeh5ZoWZnu4KDyOrOJvTpr2bg8bFN8TG3UKx2xqu
p+BQqksw4LoX6bVNRlh79jMxWpBdp/7cRsmwP0zdbykpq0+SEdE8IGo2or/6BEb7eJ5AVQS4AYf1
ZejqNtheZf1H8SiScKgCIx6Y38tTiB1OnHzUgIqGsoOGHk1hnA1pyJgTGoY0/4ebMEN/Lo5tqXLB
ybMT+mw5e30/zKYjuwQwye0k/ZVrWrHImdZkDkRHDksChVaAtMY1r7hzOSHG4c131WmmCg3+pnHR
KBn4wby3xX57LgZIke9GYslp/Q5nd24iB43ctwS2Fb38Ks+xN/s0kMlGVzJacLC9R7KI4A7wQHSw
KON62nuRjklgnPyNktFfEwyMW+8OrVWTR+zlsDwqphqjtJAo53y2Z6zsz/4WXSRfwqOeFLo7OsoN
bb0RyZ/vCMBjSf6p6le3szZY4VjEa0rGpFMMCX5BcsNjBn7TApo9c7lmsq22IEPxaB5cdt/Kk9pE
A8Unu+uOyzNouywD71xyGIAqCY4ZywGtRdNV2KzIY8YFFp2ipdbXqWXfwCRtcg3yMdCurMa9ZkOO
UvzYFhWC60HfBpcLBqqvavoDJmxbOD98dgABe2/c7pPvDLUPS6yeBqqYaxI+1p/Z4NgQ4qQla2a7
Uo0VVnfnTxfdtKCEd9XTBjYYJCER4XBwN/gGEK7nSJjPrMNThOD9dY9yu8941dfs/FoBh4L20Jur
H0/3mGNMhuxcKKvkfOlZI3YFNId+9qsXy3vnSh7Fl3Dr/AaXZ1pH62PPv3zoayCU9fLFVcVR0/B5
1m2my2RTQV9RkKdZg5VeDUZ+WSHMJ+U3v5RRi13HiGSlhJdMbnUHnwOZiOHER8rSsayuroPVNHDr
0DF3oPdK/jszrRIUcBPQNuorL0KCLc8seb5uCgGYHCYpZI+GJNSFLR5LbNe7YQ350uenEMLv7h01
j0jx4bfD2WasB8M3s8oFNUcTr9jB8H4SUaJKhccK/3I4dUhC1dIxwxbQ3UvNqnAHKhCg7iFsrE/J
7K/Uj+DuCy7DKehpJ2zoRC6Pxzy5aiGd5QT6sRaLZ3uI6PTj9+o14h+d4REPLFERSUmSUlDZZQsK
IBYxJb7QezPAUgbK+mbqKTnQxz1FlkGK/POr950UqCtfVdk4BbMOfvtFrhqvfqPqxXB/B3d/9iuk
xOQ32NDkxzmh8QLfikebtY1vO9XzVf+9+iQ0kM5z4jwIxtd+es9Lj58mJpzydF2lhi7vofse9Vc+
FSQXnWov4oGAs7etkcqxBIXeYcVVfqwYoA6v+kvkOb9uxXxKuF3jZTIADFou1GpPEZWDPWdZMtxi
SVb3oabtAmvn5zUM48r298/hgeYY1W7gfPqdbBD/vvESCMuiJno9rdzO9U0SWW73HYQT2TvnP0co
wBFZMcpvx4WPYks/lIVzQZCrupIyR2va7xsWQyBZcPLgquJg/2a+WWqZr6IuCmhnWUdUFJcrB5oT
NH6aSN7ez6hSAmhogu0hik3atPozGKjV+eyMkhA86VyyeklleRiONkSKYDK4L5Xowg82xJNtUpJv
MqV5oMAYhJJqcrS9ZZOTuYRLuxdAxvaYvpLfUh79jcMeRRV2hx+W0kPvBu1qV0HGq7li0MHv7Lxx
5nBuD75lEQ3c7NFGDgwkb8kMLC7USouA8tuTtXTYXyvn2BNzGYxdQ+s+YIvch4VWx6NMRZxXVMfd
z4lZdmV8/skcuTEPcBhNuwopOuMWM4k7NeIFaRpshlkIdpbfryAABKnzp8VcGTnbkNOzZaSsodQ4
Wg4WLvUKB4ua8SJ/25dmhmf/U2e/Ji88aYNRB5p5Ng5uD21uZDtK94s4eoJpQzI9zqO43h8K0zqY
ceNdXIbqMboGFjWdYJR+5OBlV2jrpO5QEeQ/krvU1gEIkreYsL4w2/noq2gtxevbx/uPYSAcEOaT
V7fbV4VmwkAE9uw089NfsL3364CxutUqAKYBUSZUpao6CdvstBIqhlamhz5Z40ZdKIo5XK8eMZaj
qmJFAzCUuseRHD+lpnaL55QHcVO2MIa7dyKCOmfXamYTiNvukDVCof4GMUKbVFse20xqx7Dd2wck
Kr9eqbkPtWBmHZAqONQMCSOSGUuxi+InnCXorOGLGwPgLFGR1AmINugFvtwxLKBxYnooAboXD1zr
3tIAhkpUncgfTphPnzq71opY9fouIGUFoT6pKPwwaxjt/YfCEF5+X29Qvtw8DQm3bFWn+sjTvvRH
EWA+pVRy7NBzUXmO6APTS1nruCdUHdcD2L8HGERkFx8GxbsApdo7fA8aVwQu2fSMacRC2F2c5lLM
RYP6P8ZRLeSWLxMVOuJK7cBg/VC4pvu9qJBB3LtlXm1N2JMp4P2HcOxmix9aEa4mb7CUKBjsP2AF
q5dWVEK2rMTVuXypExOEACnENnNedYPaA9p8Mb0JozqCHM0xSVE/gJguMJ4AFDb9hEved0Bon2pf
askIw63pN3rZkO2QTsCLGfrnGjv4+gZIk54OPouT0z1VI+IOH6JbOELGKnlH0pde0wPLoZx8YWod
WbsPhY3/vYR274Too5sxdt0K7502l48apAWo6GnMcKnhQFwhh1LLxRGCuc2VQwM0ZBSNZkWKKFZe
+YNHmhHgwC/sN7izaTVikxlUr+3EdZJrPRdMjMw0NUxdD7DPscsu+UzQ4kgnf2ktKzcOokyXCrGL
Op1NbpDfyhkjUIs5nthGpnecXWY+Re2iGWw5DSRO5Fh57XQToPFzda+nIFrN2pWAP6/xbv/KwPFj
KIDdEcLaj04sdtwGF8Mns2hJT2KHjZp65Qj4Nb4nd+4ZaYT3xWpX7t0E4G6UfqumUHZafBpvTgUE
V2Aiz8pBviKhBqVGykt295e/z2R0vLp8uPRC5RoHuxWR9D0rlgU8jYuONN0BNHvB/IhQ94X/PBOQ
xCehyPfw9JPRsQeU+Hw8xcgEYFxSxFnw/QGKsYZyYTy0EL7q8+2LB6w5Ka+IdkooJsrYa/MKwHoA
q3IPuw43TwgLLDSn18FqYptZKgKMHFVjz0SWXEC7krXDG8A2piXmEhE2LFj3ujXbnxBZMB6xwQsR
+gyP3Mh3iiR7AUowsMazmA1bHTukl/S26mr0rhu3bKFRWgo6SfeNOE8gDn/+JyPd17yW8Gr6TzAy
uif7LQqN0ilFq+0KlIPYasllTRRLIG+llCfxiM3gRluwvmToA1QduJC1AP6cjQIm2ZUaDRVVh1XT
XBcHvHeZ/wyMmciKWWsrGcTpQX3N406heQwBPStwSw607L4fz6BQbxeMZE8hzCZi4Mept4LNy7VS
NWD7seuPpZ9TS0ozZpnv7JlBH3muHkEk64XSjViYrmUusnbwvHlb19QNd+sBgerIE0yeIabk6XII
qVpdzPIDjPMh13yQHKQkd9WQUIJpmOUDs+ujHBwQALt4ZbMgzrJUlFtrQA29+XQ4VKAlewBlzou/
DF8gwo4qhyHYxEhmMsC+n30oKBTDmzZJsDboh8/o4fsnXv/G0T5XWY/Pn8yJsO+vS6UJTd10nk5b
oCUTPc7QxiANuEWCSUpel+eVZ0YtrjDlGYIaWavUUtJi1etpEclrnkdqcHLqzKzZeT/FsPLBiULJ
JD5ORMVkFuBMtg6TVH8cnjSTLS/1ixmYKAiPcnUwySi1DAd147qZGsyIsJET6iW7NpPL+ZAW8Ym6
7kCEoh3Fe8IhN+cd4EbfYZj3GaJgdJf5sCCuDjgi2wfZ1yHl9mZxc9Luf61sOwuLJrMa41xM/SZO
pnz7eJ3sTA4fUXlvG5TaQPFY9XSROnqWonXl0gXYayWtz/OzJsTth+H5A8lA9g5QASJbovJqlNE8
fwNQtlgsNyzi/lzgLFLqq/O941LzhE1ol8SBvgZu5zpXFvTNCszjouhXcyVHqoYFLkM/aixRExz2
NxXKvnnf9AKDtajaBSp5h5v0QQZ5amEEjj/XsahVA3O/Rg7AQpPV8KH8xZBwvCD/Z7m4hNdDcDVP
K3rBUVdXdw4KIp+snwJfTStzB6UTPa4o7dYxSx6ffLORlgO3M49SzDrdOkPXBrzJZRWPWl9Q+hgs
5l1QnVMHndjWPCQ+WtEbsFFxRFKb0mYpZSWkQ2adtfB5XKKcWBniaF4otPGorybhFdlV5uDlzRbi
e7ywrqNWpZJrxH1Flo3V8awYxHiY5mH+8mdn6wI3P0eHw9T10Tu8b9K4h+zP/DeZ+wXAwZFRSel1
PqlnzS4XNgJ4pufNaf+OFhBcQjDPUCFn4ff7w3vcLNn0Sq5vbpWH4ZNc7pau+Emn4Shdd4JKC00F
sIlV9kgIcjFXmKC1Ba+Cw4THMtffq0gdeNy9ksZeCKF+B3acA3SdjNRaaNob7KTXVl7v5sfNZYK3
3t3ywXZCqWMxKIQP1qGDeZXky30MN4BCLbKcYi01i1gH5ORtQsQYkHi8FRMjlDLYG/vZHkumZIwX
PUjI19HVW7KO5eEX3XPkvlgdJXfUSree0n/3nITDHZNrEYYTbORWHLpvQPsGFXu9mosLIMr95EnK
XKRgtlyXW5FAeZVZz43mQ0ga3gV7IRZCpF1/JZ7TctneUnUjshxehxzUwGr4FZ2XX7q5R+oHU53I
iHTi4o8yR40FhEFkR8LnvMJZ8MXhLn7NES3cX+KGlIBKgJCIFGzzVqEGUm+m1kKtLZEDFV7QCA0u
071icFZk58rkLXr5rnIIaiiQcUPWZFDpmXMz3s5DQX7iSVl3BemMccQHzrVezgdgmtDA0jUSFNya
h/lrDFLMV5IQ0Mv8pAFcZG2XMQPULxg5si5QB7gUkKeGa+6yrDLYv6pR5fyX1E0rFA05K39tZiRl
XO9tlUdIkubxxlZ/aNizQxAkfjt8MrLhUihDhVbdnR1XkIouZwdmUZ6xZHW2KsLGHcc0xJqkTMgm
XmsnvUH3ROef4ObA2SYk4uJ5rwhgBBH+d1dc6VxfY31ahS86LJwuA0NiohtPGJN1+l33w3VMniMU
fE62tmK0O0HIhCmhpnQXKCXPfnwzzhKrMeFkwyHC72S4BINy3A3aOKJvv4JPYH3NeItL2Zo+GYaS
2+TF42Axk1fszSOaTXRO/mQzK+6gQGCk8m/vxf/hNCG7KtzPbbRjgmPQ6EqYbS5e8B+j0ffZ0QBR
y3BoBhBCHsSkyVbN2IXnyNb7zzz+Rrl5sUM0sxeRTY4Vs2C7ChUH02zwpgDa5T6IEHtFKIYr3UnT
giiVtyD54X/0AAf6VG6D07mTEr3PW3MiUk2lYQ2qZ1oc0hbsKaQq2q31SKuLLrXROl4SMM4ppVQ7
7xaoQTtAhes8e10S/qeXvSP9q8pWasS9Pjo2Uw5KdqtGNAG7tHiaq9SfX1bnXgIoSEKhcVpYgWPy
AQMnHmKzkmG1CqpF3FEH4FjAVYMjSCuWFWW0EsYUOpgL/UFrTQ/NzgJ+EhLi6CfUijn4t0RlFGHJ
OO5w9jXTl0vIzCrQWlVhc6K48AVlZtMqe44jVnUKZRcvJZFU8WWSL9g3fi5qRaM/p21P9qtfILQE
eyPBgHAB+SRNqv2Jn4yKdP1U/RUSmHx9c91dT7L5KzFqvSJM/lNi4vCqp92vTURHCN9nxNC7tqr+
T6vnLuyYeVAkNXeOCLhj0Xq3knHRAYU8duUDqW30yFweBduITyBBvthnLnjhyhQBZVgI5XkgZgVJ
1eFdSlhy2FCwk3hpULAWflnRwxPPJSZGult5fGuibt+/iX8FCVw9aRqND1ShjHtlSwUtrc7Eg9hs
zMidnL5N4qulGbatrLyzV9qrU+yB29kl/vqJTmyaklsehtKsFxOlpIKiLBNs5hqyJeA5nA5FA6JV
k3cP7SFfOP56MFFp9Nf7diBX67X/pLhHi8BdIVW0Ab5gAztmoGFqk7EMSDwyVU3eSgSzaSbiqy3m
CUkIo/1DL33Z3OSZ57J8NYo0vguf7hO/vlb5PMmxzsS6w5AWSys5QrpvwOdqceu4qOpRVKFHbvRd
C8ZUF22jryRKpEFiUdQh7C94EzCsJ0CaKqvQDeMHaQ6i8tTg0VVJcq9St3P8gZdIHfrJ3GEIv2OJ
XN8lIr5p1w1h/N8+t27SmAXB+nbTq1tDEYe/D7EJhg7c7Pl+db/Hhg+Y1ClmR+M2I33as5BagxNA
5KPK9xR7yK5PTXeuIUnVU2xXoDRz1wcLmrDLahg7ST+CPNsrTjGTQFEutp9PAUlENw8QlYZKhp/U
RYbKCtUhEtscz/QhPIkmHjuuFSQNTkBFRfabO9ZphwfT2k5ZKdTw/lN0weG7OXvYjPUqjh+0ZI23
suAZwlOGdqHioHuYRKWIqrGV+ynOFVRyOKuAkn9LQFIxGfvwouu1prWZhYxtVEuvrwE0v8K9AL2F
v4QGaW24zw5UJyExNxF45J2YR9gYrAoiQBX+AB+Xm4RWRQ1fKcyZw9A765R+DoAZLH1ftLh1Eruh
sbl+a7BIvLqeW938M0NYuWdAXAoac9w3NbdZDlqIT5vzNU8g0DhDvmShnGA4LL8tvB/DjO5JDhhl
RXbbnvL7x3AUnBpEYjlTk72Lm9Sn7LboaftxQsqM1vti77K/FS1du3AfS5qzvjhpTscEZicRZTBg
8Aev0JzMl1o/iANKp6+IzzDB0XAlqLxV8XGlQ5u2LA4jR5zrzWXKYlLkd6xV0j8j4YXKIAnBZsAI
r6poA1oCUam6thUcZftCgUE/shuwph4gU9q+AhgLEfuNvYO/yD053hSok1GRxiVI2hu97dguM1mg
fP9cJ4n4HSWlGFUrW+vPnxqKmDAr7384cuXamQzn19OkDvydeX7ez5tweco4S7RigqYlOkkuWtgQ
ZJkUj0k43MbPJClNplTmCPAIWxVm1+Tn6pU+d7erRJWvspQcnSaBrOoINXwPWOxKy4CNTfWBOAS/
Jf98GA0sqUJkPs1RI4DdYfocwwjKAg+RXC+63boMw/KrZF0yQ2xBMoUE//Ic8lL77VF3L63Mvw+q
aL0FTebY9ZQRbUhqANfMk+LRQ7GzJWwWtbtpdC9V7nkVSB21MZOrumIE/VHmrOzsjUVzs2q01doy
hSFFb+wVDEvZa0IjZPftjdHVlOtwQMe6hTvdZtQJ05gmGW3Om+M6k5e0e5XHpjP0oDeKoSlv6ICU
voaSEt56R6Sng1rOxT+9i9esr98eI0eObfQYv8b3mtTvQ7iee0L7SHf0IZ1Hvo4uBmzJQETy4oNl
OoYIizKeCOlf/oc0TAGUrJberAYdsgg+YOrkf4xNGHsz6z37eVl/ehRucO5z5hf5Hti/zORgpkvP
hgGCJK3FUHgnXcPVGwtDrdEuylT7yGP6o2sXKSBBiukhGUU3SY4+DzmTWDG5odbujfST9jfBZje4
l4JG2r8opFmcd+tx8xe4cxu4F3OsnBNa8/lbidV5vrt1tibszYNYAlO0pgd3ux0WsMVFY2nqSVpV
5lOfkGk95C2LyBCXorP71eBuvU+eHLZ8JuTfICX9YhhOHumfq4wlCNLjBn3QR0F+80jXzRlw9bBl
WHRWowomthe5t3Ht51bSux00plpIpMVvt/BDTl6eOwb054LthtfooqvfE3mug6Gpct1+DDwnaEFq
Ed8w6imTWGYq+0Eg0ITncvWVBaKhGMaai1YcL8i4IjJoXRaOXPVDszzcxRqroQFHxXAlaJBRh77J
YTTSU89aYBAYMxrFPqoVyGJtwV4Nj4BpWY5m2zVOAUy04hMobLOxW5szbO3g836VOPkIGrZUqANB
b2nq2MRzzETzjuexO8GLLmhUQm/lpQDk22fpmSUJnJ3KEurvn9GEjccPeeqL1i9F86m8aca5CFUO
nmwbl0qxUy5xEyhtWIMeOtrVQqw0gPh+SyY1nyHizTUKcVOmsSEdB5mnKfFNSsdpMJBfsf4Mya8b
dcsUlb8/1e4T8j7v4y9BV3+6B7WxToNCvlFGlhz1xaM+5ktZm5YNWztbc64qeTB4leMzahmBjBVf
WUFZeG2MOijNTVDiPwnwYLSNJqlX7RxK1c+CF/lzT9piUMT6HD11Zw7h7vFgjmHOT/H5CavpfKE5
xRJdHvImvAS48PCsx/SZCUMK5cBkmp6BKwJAkhgzyn5KN+unpZnPDC+JWaqJYbyO3LDK6ujcPiYR
4PoTotfiI3UFgkUqBF+gw6cBaa18La1QsgE1qM4yPcbGqyUX9WY6Dp7L6IeIIDwwXDJnZ8gKh7dI
2Z14XaUBTY6KxbFdBQRdi86u/9SA2Hy0E/08mgZXI2h/VWGu+kHsqkRWWPpDj4cD9tXOqQPtCQOt
oKR3L7uKTPSd3TTW5bxtgiTbbIYQMU3UcEFT6MsVqUF2tOzTXgj9qLtOobhO7pg7pri4V5i4v0w1
w98eGaZAsW80fVCem/ZQBHA+bCkEDPEQwYjOysjSVmYR3D5d1sOd6KDN1aeB8omaEcQs/PBrrkxP
guV/ARxvLMJGdXkBjTtkY4lcfKCjUp3QYD2JYkBwNgFJePURnmsfmX1MqXZNx8STtb4ObmRmQ6jH
UIk2NpLXBRQkfEDqSd1+3icEXiz4LrYdbKPPIIohuOjVrPQ1qSTCZUrbMYMczMoShMaW4ETyREJ4
EHElyOFstdLTS72OU15aSZhxxeRo0hkGJCsDtVlyGgG9gEwwwOWzLgMnTGiURetM1kw288Ikmgxs
78+JjiEoWhnI5+uxLaaIBEhh1Y8X2tFpip/8Sr6mFLN3f1sNEUUNMITvJLq2GIq3rHDylgdeNtpn
JBjewu50083qcWSP60XPw2+4BLNLkhN3VWK4w/IWkcJ3mumQYQeSpDCCGT7y85le2iE6oq5lIpRW
mqQc6pxHBR+bRavbcbS0j1BKSt03WbFk32K1VCoMu1GMv02KE586gazaiMJYfwPfr+XRaUASzA0k
5O6nHucwZ9mUCYy4EfwdY5QhGONHiKBhH+cfmCA6R/+8TCrpajJ6F6K/60rZtGkffXqnNmlQNOBK
MG7iUZbUehp8F4ZLCyN+cPmvA6Qsa5GTtL0dKsHz4ia4K3FLuLR9NWicMWZ8z3MX7wba8Bu71h2x
EGknCnDW+Ymj6lR11qTjqIMF22h3YFX5QLiFlpb65rm3rcNSBL70sUQfH+QEKEOEw/+t1cDcv5I/
NLD00pgPdkUWMNCup/9GmNBC2sVrAEfqVsFrJmRqWNrUbumMbEZ/n08FpChAzh1nTQHlpM9ggwZf
Pz5Q+UcIpfCwwlyI7pFIYEI7GsYBasaLFCIpuMcPQU2uR6p4JfL8VgibBF8jlbXO9h/HgkLlQ8kr
/RB0vW39kCAzAh7tw2yvPQv+xYP47TrlJliZgGy72CFYPUzPqm/mWfA8LIQWOZMeILTdfxVDSdZ9
Y6SLnDtBkdzTDbNNG0SbS5XR7RDqXGTBQha8H5bSFmhz9IjDN55Xs5tT5Clr2IkTOPUAUMzsh3qf
cvhtwPw14ptR9Q1i9r6pbKcUoy6HSQ6664fLHdPaxGkgQC4Lz6sGd0cf9+b6OyO10Wm4dCMO9DdS
v3VAYIpyw9zDZr6Ibz6R3uj3hP4uRGop5v44zwMRwHMro7C9+en6NfD7O0ZEKaNjtpyCsY0tMSWg
mO1zU4CuRcMtdT4YRTTDZ3KMwCmDMP+8wvq+AXuXDChWMNgBPOFetzutSG4c/p37n36JABzSX9P+
gNpKa4YgxW2DBvDPljvXvGhGRmlMtMDz5+LGknCB3YYFA1LaPqFvZPt7WBib7FGRjJlY4fg7La9T
w3RBMYW8pi5RVNaJV/pJrGMDKHPk8mxJmf4u8j9vLRUTqoIA08jZoD6fUpyrbfLdZ50y00sIrJh/
Bwfhwppxtv0U/jIpok/oRwla27Q6Ddj+/GYS9ps6wcrrEePHfCizOzE539NU0Nm1BzSRisMKkupK
cNDI/EnZGyW4eJ5W+zp8AxbvdiKulgyy4lkeVE3ydQ553JOx7shpYjfgZx7eBZIRUgOIzFF7OmGZ
LGMN7mrsFnkY+3rFWDkOVyjSmoaxX8dzYmo8Te7SjLDzNIVaLOH4y8NNyUb9ZouVnnjQONIlAXau
/ZTfBAu7pL+1/Cz2VGInWl8iPk/Vi3nhbaDLm8awtopmEqvK9Ae0HqIJ8ZCFxO6Z/scpPQiLLMqN
2I4gCA5GHt8VnSHClloJIBmNQpKHkUv3Cci/Q2UAO4D48LedC+CL2aqCQkrScGrRPM0SgnaInSkB
iQL0X5C5/MOZO2IqvF/HqxmUMZN4lXw6e5J1Oo7C0uB9Ppqx90/O3mFft0ufEiN1f+fTdEHNWZ5y
sF5Bkgx45fvRafzyMvsXAPl0U+qxRaURkgNv08ist5hpVhrymWLFbHAy+VxVoWVhghEk4PDMiOQV
/2C78obFSv7+CdvBJ9VEjI3i4NaVUGX/ckEUljylfvVm1Q3BkLNCVwJaLbXb5RP58WCir5ouezFJ
ZUrg8SiHssTzTFoebz4H9B9r5bEq3rrhj7GbbFmENg2PG0wj4yi3eQxSVoF7hK9U8L1bpf5uHSg7
kES9gby82ypdEkH3JXIg7yz5A5jXY4pys7pfDHLJua+j2vP2c4oJOZLS3haS/JLijCsiAYWnvAXP
ygckkJiGay6MkD5ITzoNUMISwjiLjzJhQU2KbBt/12ArPCrlQaXPAXcI3BGmNWv31MT+9ElS0FVE
hAi7ndiUe3HqG+8LByrV3tYpUqu61tzrPlP38OuQwXg9gQ+q+A3A4d6UM4pikr35h9LBmj1D4ots
NQvznUcXt6ddffPTWR5EKUhAoy4QRjlyc08Ex9WPH/k8259xa+C7neA2AtS5X/NhfmEZT+i39l1r
Z+kilIbfqmUIvasBFnkGG6wNUiCeY1fNXUlhN3C4tP0I9xMmLMo21s/WPP/utOCqaHDZDrDDKEGR
D6tFlSke/DAyAEz7qVTcWHidnCEWUpnkacJUI6jm0bwHsIoQl5mU/vPgV8TBtX9cfvMVqYWxXlFv
pNBOWc/dZQ97MBkjplLoQRXmE7TJ4wpGTrbGGbU1NpKQTjvts2By4Pw1S+SQ1tNLjt4X4W6Fd61t
7afeSg+Boa1G5iwst1cV2V4qR1hy+8iqRYLtesW3d38eivf2SpgtKtKJg593CAQKp5/KR/wf60RV
q1S2Ux9WuzWprTSZHCJugY5mQJNn9I3TltUY1wFUpVeDRLZoZM5vDo24hc3AxfG6opSGMUghxvpe
1viFhE07n00YD5i70hXsKRkvrBOqMRSJ9t9wkl3CPmZmNVqu1l1Ukr+LTK3cOUVlmxnG6lA6CAQX
wetcozzVXhloKwK3ccseW4EypIzXn0hYaOcIIN5RwfrUJ/za4UBqPBNehHtMANa4fIwoGU+OIxL5
rmChc1V0kt0JNGNbRIr592n/W/1N8mKq2s2VgZcUE6dsi0rhHofO0qOjB0+GdwcnH3dzBNT1c7h8
TRBjmI7gcEnjywfOV5Y/+uxK53GePYACKug75NlH+7v7Fd99B01uQKaQXUh0G76W+ozf0Mm8tLZx
d6LGDMSm+gDe8dz/Rm6xoafBpk3sgHhN6uYZtYakOWgqBlIdrmFt0crzgovy+yJiBdy96ZPTvrjU
sg0CAzbBDJmfp2fsTu/nyeHqq+AlwRgstx6EwVZTUIO6YFuUg6Cq6ngnAWY8d2rWIPF8BXblqUnj
/MabuzyZk+hFe5AB1/CEcpuB9OFHK8AnJLMzPLuBNTupsRoiiqgJrj6EQAoeOK6fHr+7TE/xoWon
wH0pk4eTBrXmbvLeXOePUMxDE57I9KN5CrSQwVhgVOd8II8321oNa7pD+KkZXTc1ie1H2JnYyeMG
sztf11eWnIUEH2pYscs+2luJWxvyVu+MyexQatd4rZF13WjwqD9Dfvog2slfECPIW5sbunayvbvy
eVC3QS4zTy9woXnD1HGkrQLCXULwsjgVyBnBR+rqDbjZyyRyZSacCHAiNgKsQ72wHXqB+Uxk6Vf9
fjZX94RJJ5wiIPg/vtl6t9N+Ua4cbJOqf/zv/ODxxmDLF90H/vDy87+GMFCvC5fpeUSBu9PoeWcw
MREctZKigKVnVtmQAXXXnUG05H37CvgXcjKKwI4lmt5USwT3VXXYqUHB4JyBP26D8dutvLVeMCdY
W3tADv9Grpn/RHipkjgiYbA3IjA8S2Z1cRH+yJhsg0Bd4ODD6xR+eBdTR992q5tXxLnaGQSFSgNs
H2FhKzWFAVj4/i46BwkGtBgjJH1112sfHvAwDhuOXcjE+FFuawO5hiLRMap6qTLx7V6nvn35ULBL
i60dbUMhzG6TRKg9Hqb+xtdBP2NYGJOjFZJOJ8XzBI4F6AqJ1QZ1P0R5YRrqKiOvY19QFIkeuD8L
NV7y+VqKSHNB0HAoxZjDEZIA4nqxxJKzSektYB+QMjnmhp7uY9YnlWlFfrUysgUwaVvtIhwLiobI
nNQMjFKlyNgkckzfCwqHFAttWPEx0eogXCFCJ9PZ40q6QbcXrVJneLRUS2yPJOdL9S7kns9r9R98
Qf41NcKu2GuSh0N2QSpIQUbu8e+mzFidHqdM1LnnvJNNmHo5w3ky9i6m5+V3DyN98rGSkcGpPMYS
olSmsJe4DRIYuGNzJfaYUVMpoPQHGZ+HcewqQLnx6nMr0B9IqJkpFaVLzT2EagVMzMUKxVuVbfNF
e3QnxH/s8kkQLyd0ckereFeBAxFqgTVfUHtbCTTMe+6KCbp8kIiEWN4yMv6hlkMaaIC5KwSrB+J5
1jm31tPbV8zwbZOsmx/3mZMTikjfwt1yfyOKaliQdTVjB70IXnCaPT+x7/p5qxOdB3DYADcKmv0l
xEHSZqV5F8gJpJEhO8IKU4Eau8rSBQvoyhLFJxtXFPtWCzhBKWv8gltoNgcwsw+EQMpGjHPvowXz
o+FP7lwr9C5wAZ9h9HyLMmVP6FTofkz2IUw7KAJZpA7ZbuJ7UZbMhBdjfHunX/VDaXBN8HqFxKPW
hf0z7TqbPIg1C6dCZQtdmbi5cz611JWfnuapCTvzyT0oe3zY8cndKQX1mIeiKog15zCJ/X3Wxscb
yVZC0fDnRHUudhQSSColVVcHcVIHxYDSvb4O92noDjEvxgbB1TPH/+3A42RZL+lQ95ofhN18Kl/y
ZFIhkaNbFnn1WeqY/v61+a/qapBVKHbFeQTQB6bb9zAGyW4AHVsBx1RYCABAAO5YxUnidmVvae9w
NL6p9P5CzZUEV7lAf2dASMzv3qWVgcSWYoS+dyhFZGF/2/BhqK5sAqjdkFUtZIF7TfAhQMdHmlQ/
9/D7vSzTg3sDqWBNgAlzZyxK5miCDdRYS6o5SSkKvdY4IlCauScZRz6QcO+hzuneK69x8vFfATC6
WOL73M4IKwOhw4oG/x6kzUtqDwGTuk6mHxJ2zVHfhDc47pv/TlUlePi9wnYTlUQxAlIwgqnMQWhM
eBRpSyUf02+dOVZ3uyCI1ucjQsfObeSqZi1q39cy6T9CFG0bcuwIXiTArJy26jTjTM3JzCtc/VKM
p2h8pJrejT16yxqCrglxYGt5/Q++H4jADx6uUtWYOEkIuEFzrkMn5exyv2KaAr3loVAIUELKOyeM
yTALq4w5gGIfFkbM3ANHRSX7G463TdfPrim9IxM/M/Y7nhNo0sJlVX5plTUqGcbZR+QlDqZ6Bc9z
oyZO5C6XxBZ0DnPhGK5Zgh4AuIzi3N2ufxz5Obno9GTnSAlB8Oaj2sTd1JEoN/86T7yQ/vl/vB3r
RJmNoUmQ4wL/4fYjpZjqj7Ip7q1zV+/hooOg6gc9bybzMlxF9OEZ/SLxe3Fx2ZYK2dAkNgzY3Pni
cmF3jQYajIxw5zTv6AZWK7wbLVvFcBJnJiuq8piwtbgTnHnBenY8SfK9U6Atqw4bKjzohI+N2PCq
aJ9K4bV+HT+s1fFChYdSMS5rtAc57iir6LB5+4omYh2QJltHhaIJQ55uJhmYbAeM/p6NZZfVjZC0
UUdpatLtwoavt512uGF1w+DqR0wwQUSLKMkL7bk/CJjsF9hWHENH5wrRLrdquhICpYilZbCOFZnL
HBqKob2Aars3XkkIPNXxsbYiMwLjMuh/nOS9CGJCbOrtQ7twjT0w/lA5VN3LIfmpqy2N+MpzFjLv
eEqomy5y+ITV16WvWduaRwgtTTVIEWd0S1hUHjOvDKZBAA71OSWFnbrXfOjQZMBbnax9I93VBNG+
PaV507hqmU6aw2dKXNxhu1Q5SY3zwznfkabhfSfednpvIObXulxGPhpfL9X4fd4G3NXurB4Tr2vL
Z46M+meA3gj7oazzyb0OAMK8sZXhr/rYLEsrAKF0i59wcwncmfVDug80xQywF8lB7XumkP0iUTDe
PE2ROs7xqx8sKIs2zn4x1D1Z9VCYU4xP06VIHVIjGXqL9/h4wyEo2yvDVpQ7ngyoXAr9YyYe0DKS
/Cll9s6yPYCfZgZpU0aRfxum9LGxWmrEx6VgfmtpvfpuoVOPZZ0IF1yR0IanE1z92K7j9T4AgOA5
BXcXU81Wzlue19n8d1bBKFsCqz6y39lvemjA8Ih3RpLEr+yaKBT4RjFLjaJ3rIzTZkAJyFLZ5PYC
QI9Yugq33TQMQV7MJUwpGvZo/HyZfIy1Gw5aLAgI4sDTkyQQ+GZS5uXv1JLUKOfO4d/vfCHyLabX
bUU/bAEI/hV9ZpuLgvxxprayomzraLlp9EJiOqVpOvB62EsiV5SoCzsp25dOv2aCdBeEEakqqdeJ
eacHqtoKZNCTg2A6WzgVAcw0IX1eddEzx+x3Ej/3LC3KMGtD/fnTmh1u6z08AGT58uqx3JcsOY5W
yjgi1VxcFIMb+x0bnbscf4PbO18Z06rC+1rk/2ZB/UJ93UHcZLuGmb2a/f2OwT3Ujzhw9y5mzQ2i
uK8BAGjGvHifQZrr3RUWjEvfHZm+DD3dPPKKtaXuKYFtFA5/1vVttnseBeKRdn/OlT1EE7M0/jhS
Hog6TN1/Mh7yvqQwzXFcsiE4iHgwZrxwR6PVsmwUU55AZG1yZGFJFsoXe3mZlsOCKiiIRstJL4Hu
2K4VyUddXf6tl3SL8elMQ4v3b9b4x0nm8zn8KmBIT8Iw4gtXzNAy1CwmzkU7lbcq8qP/4Wm72fXO
s55z6paJWtm79StHGHggazgALurPtVRGskMPOt36n6F03MO+MIB1wEgCNTPfglT/XU5u03R7fwl/
9pkyQOnqRU9hxgXzHCTTGMk1jBgbEkCaL1cb6waQ8N7Jaae0KesbrbzzY+o15BvNtsiqH0QgbXcV
1MtP4CDwopJmE9yEpfIXsi3S+0kRPYCiISPjUGCFDXrD8BSqO0Ld4tKGBr4ISJUDjtVfKpZZDVD4
sVdimlISgzS1PKZc6OaHw7tSggJuZBD2TTjvU5XjFil0TaFy/+/ySW3cKJHUx0fpWVbWOfPcIM3M
0ZBIcG8Mdi+HuhXEpCx6mBQIAyL4eiTFYOm3bOsGyF6w6Ya10prhl5SmXl42nAswxShCXSVpCrsw
98EGQdAjgc9/Tnsfmy+vM90ImzE2Fo+g0Y40GvvBt+aDrPHj9W8sK8UZmFsRFN68YyMOBCZUBPjZ
zxrjiQZ7ZWIbaE+/y62MSomtKb0KmFSIzk5iFAcXoDcRH1CpEOynlWAKDmZeJqs77YD/ASb28uKe
DYGFDCMEvCTIe98FsShY7zNYfat2Jf4GlZbmV+TwevU0jMGQF5RWSC0/OixGrJ2EqUtQWxZKIiXK
k+X/su1wWxfCc6FsS0zVuNxy7k7koPda1opjVtvGnqQTK3Xz7yjjHx0AEgA8HyS0cZGIpYbHHsou
1EnqAmWBsYRk3vYdxRPTf9e+DmjXN3NxjD5uR9B71zOIH7L8bMuqI44Gw1M5i/ia7Z/dfic8+cW9
VHsCcr86oNs9lBqsftze+QfULkW9yzONpqLz2F+7y0cbW/uUIb63vzt32VNIXk+KREIrboS71hZB
3z9lTexqVDw5nGTUy9l7d9SsQXeQw8zXSJdMi9cOxXxqVgw8TLUAp7Zc090Lmk6RTGCG/oUyR/MC
SdeinZqJmQDdeLjztxXjgobebKqSe0mxjiiyuHpVhqXeKSievrvoGg/q6ExMAX0zC5XjASvT4Cbr
mLs4LOxozG7W10m+G2eBqTwn1qfR//AdEx9q6Qk098iITzcVwbv+oV/1NQOG7idZ4beBU23Ua+0B
s4fgO/HD5hHQnl6xKcA66hUiL9MbaKqqzYFDeDCsgTOEI9REnxbsr4KZWZI6cOt+BnJeF9eIcWhF
iedK4l5cuJHGHjk8K0lahKZkYmCRdVESdgOSDph2YFVCJRByi/g2c+YmqGUZbIvEfAX8WrC7hNCS
HpDC3j+dHfeTAUxOcNfwgzLSb4OIEsKJjeBQs9QjzTEWer3mLEXYDF+vylNupvx7/fD5WptEFBT1
TYcAW8g6YVXgL+ve/VjEereGODp0M0sDv2Wosl78sTt7dPyGZ3SlX0UNCmqhYSaaqS6omdU2T0zR
ygDQ1LG5WrpjtQJTj7aAxWIBm1Htko1OU0PQhdo6lFacqD3wDrS6t0/H5yh79waHA0bbFsZtsQor
VM1a9u/bYmWsldTNs5ytnGkdwcs6iNWMDF0oidZxPrLppvu2ncxtTZGA419JPXHKh0OKj9NXQ9Dy
N0sFgLpzp+STDoGxjO6Seqg1z6wEw5HO1XLQ04MPiqz0SqD5QVZnp+/sBy+cuwYYoL8svNcM5zmB
n/oE4hkIpu+5TBAocEv5XtLv3mSJG1YPNZ37eb/Vryhla4tySIxlDxMXxyHaCfjT7Y2CTW26RrjW
iago6woDvtApce0AjN5HY9Em8dw2e9L6oT414ZThqGMQJIyRUo2GVClnLvjlaRxlVuvuNWS48rFy
RXYcqwW4ncLzW6AtgHNQJOErgfaZX5DgTOVuyK2ffG2bhcB40Ta6qlR+UhMEdIPu5NAbIHVacVGd
YUm/tEE2IuqUh6fhF18M2cSzbtOTtHb5uTK3SupAXDYi8C6scAMFLj5q6a1bOVH5rDtv6nKOEmOl
7ZISN/lgH79YBAutfllqgMxUp3DrIBLGV+Xvt8rympEYw55lydXhRAuh7pTtfl2BncrZW6c1K6Nw
BUUconRzPm94fam98bd/SpOLZ/fyOBdDG+fmvbODL6XsAwY9Aai+dg/JQIcxttq5jELu0ZyENwio
7MOpALbR8Noo4P/ZnPVw+g5V4H09JeNxzq07QCibQ52/LR7BCC5JhuwUWDKQHNymyttrKBY74e86
ZD1rrlGKAL2oBvSoF/7WbNpNS6Al3o5inpa3xfiYoemkdmDBf5FYpFY8OtAv6T/G+X+SFXRFk2r4
saz5R0ujTzEeBiaSvXtNmiP2UOZqssmSZjUkUHA3iC64gQF6izIf9rzshhLnE+qJ2eacNZBksnTh
tfG6NKYMYNiyCi9vF0WZp1Yqi/h/ivLs5YnjQOpynaQ+AA6ZzuLIhUT3yv3g88FAira2trHiDZ80
0/TifkHl5bQ+3oBRSHkyaqryOwaZutIyRk1iHkRy+s6PdwFRKqn2VRuULlZsvyOzwdSX3eT+syGR
K4Zs6ryeFZ9kOMNsmuhVwG2i6aLpW3arXCrxGkpgKuMy8XhmwGjCnI5frwqC4bPVnSmvn4kVGiod
hfxWTBMKfQAJzKLaFnEMx25DHsxMWyqB7aceT2NytGJXwAaAPlcu0Zdzrk8eUmfnrORsda/A3iUq
8rQbEdxAQ8UNFxCPEl7LsNMXCVddYpLgCFiDnCrVPdfq9PxOxWntvN4yYuGS3LqWr0rjC7Urlcj/
bbhZaPmfEVgOrHM10We2HKnSE6VcGOKP82DqLUh6mqtDNJNch/OS9M5WrhH5f5IYqm507tnkfIiI
9BFp46PqlxlrqsKkTeFgKusqwyVLkojzxlPeS75Jm8wQqVHPgkWtatR16hHcxxX7ZRGgQowCxOc/
g/ai4CFt3SUCOieYy1Kc/KhT9ZN32VTjFM5q5DT88Xcv9jCwFxArMNpy19zaXhdN7SYwktm4fNTE
IdrKZDHG1ky9g2WtPJxCMhm7+kRZ7eB7T0cyT6xRSWhbvnq+HlHcTpYDDademAYzTyLiR67Wm+tP
qJWODIte/A6K3REJP6e871dFYbnU+Bxfnv2zYUJFfxlIlFeMHyy5vkMKDLSjrjZknrJ6K57ECXsg
aVOHBUW7NfYfrkESKISQRlmNtf53/lIu1v4vcLtIkxOtrCpGSTrW91/rDL2deQW61tdTxQSVWSSK
vSeHznv0N8pCQElRmbLwXrBoXZ3ZUN0Er0HtFhNjXRLVYoP1Zqx3RVYxahk7nIeF5i2XdEKFRKJ3
VCWboDt85JjW8aGvdFzhllwVWJtZtnRHrfEJ2/Tkaencgw1471wyOqW9QFwGMdZ/N+xrmqihDDgT
4ar0jSpTq9JoUBFUHqgW+GRhuFqQTDZzHs56482tv8dgN4ORhFbalA3kgFk40yR6FxqCQlXp1aZa
8BdLrHpl80h3mVyNKkyfO25JdXt3taff9iS1mdr6rYilzoTO4UxbfHbk6jbvEPuVFT8Hud75pKxM
p2D81BrUlwZ36ghOZvJp8tx/unPUTDhVwhgLqZOPhgXyBe9m0gE0XAz7etH0dPce18NbGkQ1wO5l
aHv/IPhA2rzjaCxNg0FeZ4pRo0LN1ove+0ZxsuAy4Oh/T3gDo5bl95kKVbbbJnYlidj2D/SoGhnb
9Qhwfo35e5mKe3Kg8w1j/YGy3Pe/raAJUgbCHhnHcu8Wo+h6Schj3mMV3Exakk1/yJSP7/0U/iPL
7R/TmcpCJ1xTpCRuF88TNHT81oLXCfge224RXNe2JV/rYYuHwBZac4/LlKcPfSDuqB0tPaeHwA9N
k6EWoEE8aIzMybUjD+GUQZwFY8IS6kL1ToDpzzBB6zCyoE92ahWfr0aapAYGMhZzaGTGRQ2kkJVK
PkcZH6vqzDi/ObgCScTRwpGzxyLy0SPKovUKeMq0sQO/PRCUFvoIpVSx0F+miIaQZaFNzLM1lBwZ
rFAKbAAuMaIrPRxd1Gcy4OcvyNA6v9b9odVfzNEMwhhLMYC9jx4Z7ygkoXLjahG7Y7uLiDss89ZK
Qv6lG/me78uJxWr7Ocvbbia7WPGIrw2Qs5xhLGFvwSdPATdzdtz6dPbb/Rssi6Hu2j7UblDNR32T
M/KccOUhYel5WP0vlGzudqfEk8RpBK6LtnLR+EpjKq69lYTRObr2EjOs4LPyzOSbU0G4J2MvIo3I
D2U0YkSfO76aySPizBZykim+Nbb4B3RXPKYmZ5kfiNo+6+vqJHePzak4h78msAUBG2gVC+6y4+si
+v/EcYqx6iCyxo/AJdW/SzfEzTx7x5lmEYAQ4U5t/DFJKFWBuXK9upWfXIV+l1qtKOr5506f0Puq
5fTV3hZ2/hXX7cgTSy42jCTlgqeBa0cc2pBEhyZtlglY3EKoWFVLjCE4E4qey5RRpBMViozRiv4p
RUUHkCtsxLXjVLekLz+IB9wQylC/a8U+14dzYlSFHfl/4x2AWxFSZqu05otvMFAe+OwJUZuPyKgB
EtLJR2bB5miVXbW5koMfIjUp2lVdVMdulSMT8bGlfUfYh7Jz4Hh4QLXtC8tAhvsCtDQlIU4HZ8CW
4iNZ7N0rYgAfqcFzGdbWackj0W9kZgSVjka3nwHfKJYAbDR/xveq5X4XH1Zynjse9YdCvYqMgK5A
0abwqilVa+Ux5s22OUvXKHG0sKudy7hw8kKjitIRQ6pNpR40it1XNCe9yTm9vES5o37CmGSJHxy/
symoBIwG6JN6YrkIYbezvx4D+ORIeodvNTsT2DByhkPsqKVtfBe741Daw57jNyayabhNWiAPfp76
n37gHoMFzX3tXV3qOaM/LhqiIeAzV5WzxCkanfrqVxwoXpSigWWljLuEtcoauf05fvXoLiTYTyRT
UN7fc6wqtGoj8DFSKc0Y8HmUVgRejdy9xXNEWL8fhIRanahj1gAPDF0U21pnpX49wSpRAvtPN+14
ER9kFo6xrRrIUyT/HMvLEmUvmR0f4NKpLzl/R0nhy8qg5Ogzv3c5HxGU3PZa/PLsckTkuQYzRYL6
AT9tnb1u8b1mhpV3b1P7v8xfh/0bMrDzl0EmWiNDuvUpzliQRQtuj3btiFKt9cy7Q7O8/M/ZXKRP
NQOK+Ag35k+c0uO4/K7GEbjsSwsj++EKDlDXvA7vosXUXsmOjrnnVo8XPD8k+54BbskcbABqNflP
2G8I0Jqx/efByQKTGhzwVcoYEb1/Fu/gyrzLWeTXcT3qUSJglTAS/g+CHBPUfIOsKjs4g6I5nPjX
wkTTkp+U6chnr1Ahjf3V79E9XzwB5EvN8EIsd434loKv2I/rvhZUuwYy6q/AzPZeGQE6EWnMexCM
Svjva/BsWCGZR+e9iZAXXNM0Y3mLn6v7MTFJpDoglkW9KUq1vk7Ga8MHOZ2d9XQ7Qs73nzx+qrSQ
CL60JiGMUoceKRI36VAq6uJxeBNJnWhmDkd50dljHLbMEBhvwc5n4xvpvNNz0M1BXdJSKvMK1Toz
CU78Z8W9w2CFE+CdsmDAW12jVagHwWJtr6LVJXEDN8lCffO1CdFXlNc7kerQvFY2mlwFHjqSPAvt
MJltJXUryovVIS+e+trw5eJ250YU4H3Zmt5VsppRgklLPC42qebbCn7To4mkyu04CzNZeOvKn00k
3jZQMtE7JyUGug7+/EtR9Gb+1GaHJ2zNpRNN9LMXPjsOuV8d5Zz0m2d/CKaPs3uPqzvbNWqoj3Au
9D8reW3GD2D/bWDyboCOKypqvzBE/Yp7PxIPO1N1EaFBN4ISytVmcyrL4oDallghxfNTCrTCj0rd
QbFk2DozyLw9AsdBwTaD0nwzMPfIGWIi/AcOU9Veug0oaO7Ap5+hGG7LXB0cWOhmk9AO7IvxQP++
4xgKJ9LtSAW4VOAa/OVgz3RhtjJixjcNAs/OEAVd7n8Dr6WxAMNkW2hOeAv4UCmO5oTZuaXHlBoO
DKSiDRKT51GMBc8jGogv7aotGtNV1iMU4JZW/QCmvDsBldPDI8eYmy+7GB7HV5RWLGItomlpY7s4
s63W38SppO81kIvY0F33q+6yhE0ttpStPoi60K4jIJ04O3LH0Ln7mO9tSW58SiTwYUmv2/R3fCyB
1LzHelwaznTjH43lu3BTcgairSPhmUVC7JJOtUKxfeWbYwgFf6PSEHiVL3S+3ZYducem6uwUXP70
jnMKB319yklCcwDRJt7NnX8EXcGJg13yzpHrNAiigPbIX8CQmSsW4XxSHcQBaIRAIgzwgJ1ZW4cq
4h33PEmZJ9U8XlqrxhF3ygAcQYtdArNDHaTVuyt9PDIig1ppiUBaKmTLCEwLQDBGdc/LdPWUng4r
5HowNkMYXBZTaj5MXRpVDIVdxIUj2WbtvV0lo6o1uB6wE5GVk2cbW1/mp8ajFtl5xjHDe3+KDkWg
gaxKTb0X55t6gIozFtMm/WRDZJNclzQgW//RBmurK764EjLFBbR5Q8iNGOXlcguv5PsAWKw4Ma+f
MOHliY2MPTSy6Ies0QkYxsHyBXapmAnRf1//BM8Wg2fBCo7ztrObnEgQya34pPhacwthNsYHBHNs
31rgv9QtI/Ler7Ttm0FarXqFQvkHKDr+EsYeM8zVC7qiykBWmDlWoI1gNh9zP/RHbr8kJKGBDKCv
ddfNN3uio0wKfXTqdvl5DVsFS9JATjWFIz+cB4zEitNHSZQAM2knmCAY0IFg/Xh6uq0hPHNgz89n
uyntcKEqhZmU+rD3MuXgTUDMzXTwetE/uz7uz015RNTFN29/6nQXAaBRZKBsmvUptYxjpRvdsYYd
Reb7BkBX7oOIvgMpLxDQSBVH+z2o48InFwFgLeU161O3C5nJhNALZKdAlS1xfukUf/11ZVxmE2NB
9BmzmhYqAE6p5flYG5f22kiaVxZy6+EilgW6VQEqUPpXD8O5GqSidMQLQElzXB6cKdFLQktEysIt
ySABRQGpVlceZ/Bm5Qtj+MEC4TRQJ3lvDLU7Vs3CJzUPyhht/I2Kyh+fY9BqSc/A19F39Gr2mp5O
zHtgzJCxgtSVFEpfOxUnXBibxqXxb55ki0RhQaCPYMSxiOSmJWHSdSCoap8Lzms4kRP9SZHqwZ/c
nqcPNLpRN4JSLFSsd9C9pp43D7GGLaXgupL67EiYxHwqbya04yjYJXHbKidZc0J0HeQSG1mVhGXC
gXnjQGeFqHnqgrcA4ygwTMdd5gMDAWqWsgaoTm4C2zAjjBY0EFaft4FQ/L6QGYoNIPbiogQcO+WC
x43bUwfhgH6PGxVKQyTuSxx2R2FIpaC8tEPG8GV2WV7w1JhlsGlFT+lZJgEM6UOw6ltLoBzLRnWF
8eRurHPO0vsrWTGtt7LEB+wzQStqYI+DuULgt+B7H0nQx175Qu9N71TX/sTmRiHd1zE4BdfpniNm
ohBprUYw9CSsWgh9+T+cZbWc3zOx5Vu3anKGX70m22cuK82+R4mSdy27DG68Dv7f++Wj93nhli+f
SbTCC1rTt7a950LuBCoIPqR3bQt2J5MwcL8O3pQpHAlf3j8WRYvagb9aQlNH1f8oKcTKk268HqXn
9f7zi+++hOzsMER8+EQChe+hKYrDB67N0NuwqTPQT/NMpiRSRJ9uzbTEKy7XVpNbMqNXxOfXDN80
KKBdZTtGrkB9SQbHmOuGrR0PrXvhL0gMR7VOewfmp5Giik0meLuW0PQsx/RvZldtA2Qg+qvO1/E1
3EsdGzvl6qPZAjyAB7da3tRGswD8Qrb6sxqTDZLCr6mLQ1Y+NuEIgaXbybe9zM/xni/uVuJSTEZO
nNwogVth6Hfh6oulltqYIwZJIF63Xznm3NBQtH5pL+t+j3daJnGawf+RkwBBDZzfZCT7iLql/pdo
DyFnVC2eyQYdCcGbBg29POOeXCXU6LzMge/6VVf+gg91xVGXf8NDWHq60dNzbcR520tMfFi5EH+B
ccEbPQa/IrjXQL5q2TbpHyrFeyDPJS7LJ06ZJoCWif3jnD23S87Iu3/LwAO85QNnl0+H5dpUTEF0
BT60Dy5m0VMRUP8H+zll+rA8/nqFEPtuN2Tt7AvmyxqzKrLQLQQrQozKz3vLmtivGGe3mPHYGCME
3h8iRzSzsxv9/961kNq1BPhpJVgWmVFkX+mvrSD6wi3pOfop5Ztx4a33IpNtkvRz9KGK1xGqw4cO
7ISjVgUsi4nUQxgKMkksf2LYGadda82TqA9MLIfBsuXbLBQPn+hr8ovxt3xwkwa2bwjBzQqPnJXS
rz8NfQTrXgzKrghrxIe12TpnLCqpVb5gCdh/yi1pHOmIF7rwhvT6AKUMwemgkc7fAYf15Cyu6UOS
q5314ECqs3vQB1zMGUZvnd822yoYdMwTlHbYzJ5CqQoxY9asrQ1kf+/Sq8NaKsLNOb8RV+nwpMWC
JbKPwYTdGqOO0zyXNaTYL/tSrsFCsTLvqIXEOYpoMRn32UrDf2qrj46tASWfjRj9Yi8j91YrsZ3d
FU4sqye03do3qcHhr+Gyy+F7Pr5NpMHVcO/YFrgwDr+4IgInuqOcxwgdeK5vjhPIrKTVpv+CVIn3
fbz7aGUUMGB4W2ADUaYPFvSNuSVPR6GA+lBHHw0hKVggpmyG90eypSl5bo0uuToL0svB/m3T101R
xLYZCOYaaTDFjdhERLpLkDuo7xvwBhDlCYrWaGOGxzphKUzscjK/EXSUTu6mRr+9OhPV3Qouhimu
XLyXq8zpQq+IBZfFL/4nqUOk1fPGmoFZyQDrAxv3LMUtYQ42A54DWpxq7DNndnaElwb63OY8LQqS
Ll3VKu2YvYCTDxTr29FDoW4t4zZEh8kSNGHXAAShjWd6ViUyKsASuBUnrmE5loKDtt2UGsjQ3azp
q8HmcgrucIvfARkldDfdvttWa9DuDnwR/CebjqMD5xk1iZTYHVJnTgd0D/RQSHWJwQ76Nj04Qhz/
I+ZOusLRAG/qsW+vHvrUIY9ppLNLGVJtPTINIhnKUQabt1ZwfexNk6khYaKfx0rNVUxoZea3HzkB
0tR4oLP2RtgvJfqb7XBxlWKLx5nlWx2v0VYDaNgPrG/B15zkxbNz8rTqJLffCwYlZzywuuRD2tuC
YUI8Wlpy632NCDG2P/rMF2w4rylOvrqXEtWGwVpVuUhBu8+3fii8VxrRIylVIsYRzmuaN1jKb37E
SxTODWPkr9BleqsObspLUdGPROrSXNKQR60P0KpCqfuACAdBmAmL4ocRQkvqs6/erZ3GbMSZxabM
Aa4XpMbOSutFDDYabsBRWk+z9LSRho3LOpWFmusDx2k6LPQn93kgmVN8go/QNVD7usWy/qx5lT53
o1TXb2p0EstcnkNGLdVkqoQTqTLo99h8E4+qS9asTPnnDpDR8T0uCqPBMuWygA3McJLeNvrmV3PV
kqjSGhJLI/913/MVYV6gAqqQs5QxvO5+BAPL02BeDwMHJSi1HNvxPmPK/qdokEwvKmvxGt/IYb7v
dd/Mi0GFwkznVRQd1UXvJ/xBIl+HC7vLkf9LDLNox+nKX09YGmgafAYgx6jR0sQf0yCwSQtjkmN2
D/m+xvE9DS1d2SdYa9NnA8956cfwfCbcs6s/4ZhhN4EHRbHWQqt9djHGWavoAdq41vvYC1ELVDAI
9F6f8K+zduRXUowE+22RIHrL/e/gKPFgLVcMZzVhxhhcEDTKzgunG07smbmgfprTST4NVSV+UZq4
D03zPF6mzVzpaa4xkCz2xXsseZOVex1uqTpjw2ohdNjLQoBCusNf1lgACYlb7MlANZMA1FmjMiZl
Innl4LcER8k1pmP67I91dYBiRZeuRNF8XOgmJZzx2J+0B/tBClVFHzQ3N1QiVUvFvaSzl9J24mRS
h5VGqZCQ6ahg8EqjWJZkWjSMgKERdaUJpESF1ZpB1eG4UTN64O5IXxsW/51xEG9O0rnItZucwYtt
uZyDaoKdym5ZD+ftxBeDm3i0TYmwACQLNuilGvniscipynSzoxUuufE5/1dGuqFionGGpbFvqbU1
tzlLFlYDexDqKEhAKlrQSxf1BbooiRZK25fu9srpw+6JXLH7iRzHQjGNBpOW2dbiXJQ84biZ9Hpl
sBKlWox69DJG1vSv2h/TJQL5JqbcZcC14cTFZv3pUPQEhyVM3QqUJ5A+sld0u8tjC9DIHtnn7knE
icn/3fDekcfInUHJquv71VFsXsbvEnul1lE384SCYspBOB45HXJj3wuJRv5nrLwRvEXUvIXzNgE8
S08xAUSadSQLz4RvJoHUCR3bZjiyJkTVzLa+jTxOjThiresghSe237v6sIH00Csw8A2ZQqRGvs1U
Vb60rfJEntKPl58gbk0GAFoctaXw5thBM6Bgse4+UXOm+qqm4jDY8JdzKACz0lKTuvWAq2X8vK1p
Dyzo1gCmqnCF7Ky3H3AWLij+bRZLnz+BidJraN4xd6T8T6ZhBHmJ3+JICDbZiI94x6olG38uziCa
lk2vmd4bYunJrXb5sjo+vnhEk0vNxwq1iYEhnYd6Kanx+Z5qCs3hHaM2vmKynkbugxW6JFq65YIt
Do9tpDpfm1EdR3mpDCY3PRj1wVBhXpc2b+ULmpExvR6m57wOVE8XttRtqF8IBvLT3YXGpcNz8ekN
cDwUlrFWpn2VlJUNqCjyVeGxvvnNx2SIyL1pDtL7biu/4V8MMJZ/uB02N+Yjv32RZOLkLnyHfjXP
fV/CkfQ78POTMSJFVzQWUJb3469+s8HwHNKnkpqA26cV7jSbB+ufzghew115jR1KN0URn7CWp+/q
jiF9o6jFNGIudeHZ52AwawzRhqEehNqB7lyD1cm2pd00UxL+l0UzLCzVURlQbUrjNggQSAKEDFXD
OQRwJAPNd/ZPAeJx+GZSvik9WO6b5UXhqc/wUgO6lr/oCAaiyw8J7WBU/W4q/ka2QCZjjef1CMkn
M0uJ17Maql0TfZZfOd5CgAEet5hFqY9Gl0B5URzaJ8csP4iUB7XP1v+TpZJiprPa0Z1cOuTuGqYK
LwgNTdbJaqm/xry8gXHvCLiQk05GaoWaSVm/Flc/PUIvUjGUJKpZmFG7+l7V20LtSSJSYzMVNwEq
87YLws3fgr/aQVPzQzoVOtYpFFiBeZlFeSXuYCG1JUGgma9jz8tMvIl/UmPQ9NOygTLRp2fGF0dM
YEkx1YJiWzwNVTLWzw2R/1I6jbNyTOX5EHGCKQ63w89P5ionqeFfth58qe05xc4DTyHNZ2LspGLf
4s9a7dYOOGuCxjfUbA+jkmMUmHiVuTDQKZnmwzPGRkg7H7u3Q7w9dNYZ+NJf2opF2rYw3/GOexOl
x6hz8PmUt6C/7ejVK58LeYQP40FXMNapzV5ndD5zMbCBBTfOBHt+iqgLdlU5ISYVskWBTEqkZE/3
k74GGNSu9fLDZY7lSK8mYFD3gVtoqiDg708H2PXBGi2Wm8Qc9sCTDM1X7+pTGqZdyxL9UeZUNvr4
em6kU+vPUWLUclqdLctUFSUSisPq8Y6h3SQN51nMhjHNUF+CXPbi7KGweCyNwlEC1sKEeeShVLUf
snwlYQG5FW/s222se+igMQJtg78H4V2kyOnDcCylnfINZeAiKGCz1luiTmBE9dTWr++1tiR3oyuB
54zeZRuHtlZ3vDPLqDtp7d40fG8Y3898EHh604eUgturzwr+a/mn5FC5bhCiZuTFrQHlXIAiKXnq
kiwcznW4MMEGDXfLE4tHFi9NGPcbgnJN7D4Xd/k8Bbmg+wtKWGcT7ZWImB+8+//+4tQNz6MsYDa9
HiEFb4TiWnZo29gYF3bAT+ZTygscvKzK11ArVFv/woLfxlT0L3Rf/ebjRpqtv4OS6p7H2fm9nolB
uGnKEEKdk4n5OmKRYxMPTJgAg+pFBhef05iDF3S4n3YFgG2GkyXhnk+9llWTSdfjyc9aykucajKR
lQlLs/GrHa6rQMZepxCY2sfMWPx5Y5EgiQ50/+fGUlvcq4jsQ4z33XMq7Wr0D47iyY6IDra0i5nM
Dq9jMgE3Qob8foxkPQe+dtNNiBxhNN2/Bi9rrEO5Wl3i1e0qNAfDA/cfbKOSSUFqKC+/uT/cTpW6
zPBcF+dIFIa9GYcYVzot4yrw6OgoXZC6ixEQC0PQpsfpp5+2RabP6RkoZpwZVFVMOYffY0vNWo3O
1MKHoMjgiexNcLgwAUuMMAa4Oyi4EhAUKpsm5ypUfeSpiwslaWlJoagM3sqFmop5/SrHBsNQ8uC4
parjP5/qrAUHv3HYeIMTk+vMtNP+iVLvJRZ8DjN/R2utS5HLuX/MCxxO6pUMySkmneUMMvjQj91T
6G9/A5/HmokzyD9BOtdyzWbvvBFgpaqXERmpReak/WfX8wy22TAPw6izBpIkwyH9F0UnWcO+xGiJ
r1nIhB/SCzlfWu6jybbxhx6OFcRl4Ixrfp8oEz+VhMmu6OXzNOFPsPcRNkCq95iViinpMitH/x9G
Ys+UNf+1NoCYyGrr3LjVnIfY8DRa1XZhw87G+Xqg+7aeRnn8WebMcIk24tPCiOPozgMEvZUUhMqs
NpnuzDa2wP3QgXwouC25WdxO2uOUhLfDkJN8CHnU1xuyxiHt1VhYqIHJ25HU+MSqi1H655XxxwBF
Nb80CI6EN866E8vSnM1/yn40R9nOWhw2V/JBZ9KzalrWENtgAgVf/YdN9YysvdO1CDSRF3hsLRqD
EN5cmEc98J60tCy7uLK95oX3JLPhHGYwlgXI3+Tn5YcdzsKPM9rPQPm4s5aUtAyvCL/AIV4/THbC
n40C/puAQLKaD8bQ/xjSzQWBguEJM2uD3rURM+ZHvvieCrx++2LOQi7Abd8u2GdPhEn9Df/2PIQH
WL0wWj7RBaw7Y5SSQO2m8B7IA+g/Rf/GxccCIQyByN9j3Ca+td3ZN4svdsILiDcf+p6wPkQh7v6K
xW86dLrJhDcjdg5+FcoPnYKwD9Sbb/OutSKzKxCTzW28phfIESPoW4iZeO+SIGefeDPAGTAVXf5I
cVd44V6oQpFJRu2wDxgt/2EBJ9Ps3LbJ2/CdI4f1fu+LIhUKqx/jGmqm6VDyHkNMp+/0mBkydcLp
3yP6fJmX8d5Cm5AYOK20y8QI4bqMJC3BdhI4YrNUXb9l+B/1rgbdw69Gq1f4SHuuNwJw7b9Rd/Yh
6oZNAUlE84xAvzxGUHdIx97m9hA0cwTOobLGoraP2mM8SnlxPtfT4Ze2Ac8AZNb6gNN/vDXdLFVv
YACOELhDI8BsKF5CgRaqhufM2vBBPJq9UVBddE6ZGgPra/TXJvFvV6B+OWnGJreDTDatrSet8zbu
QXIHFw/1fw8GngFfL5GbQPgP7pSFHglMFrUVFv26LNwZz0sujG6h1SxS4l3BFYyqgYMVE4uTHFQ8
7CO8nhrRPuPWKQ/KWAi6KPxb2VeIVqJWt9gn1G5tfWR1CIcqqMSMfZmHuAjVY493hrtq0qW8KtQ9
VE7jlw3MxGkEA2lFZ+BO9F8LMzV9UgxiMhdee7XNNmeWpN6zxwvt4FnfF26lZuh0FNuAZSodh0H6
Ji5BBtk3415Nw3X4CGNZ7yJRDBiPS9QPHwJubQj8Je4bZgkJSG/8mwMuwC+NeHz8HYrO56rvWD+E
Uks9pP/n+OUTJ9y1rbHfXkt84g63nnA9LTBOT/tJt8sQ5OHuRy4df/yvGP3qrwlDGm9+5qWNaUaD
oKZvv/DQtZg+D1k23BdYLvYomSrdXGR9bWhn3gKXf3+F0PsDiZCfetmVvpI3MWWPyL3HNGBPptcd
QArn6EdSCZwZXc8G7Jru0zMrHqt6qd8k2xFsMPvKJDOKoXsWEr2uwL9THsHlFY+mBw7ekPqDZpc4
LEPmHcZ+VR6xB0YZ4nj5eeDKJvlf5JxJRqIj6dkXCjlO14Ijdan8oURsCXcM62bfzuBZ+KLM9FzN
A6iICYyXDG1O2Kcad3lXY1RLYPLWcB6bc8KQjMbHiIXoWmX7jEnMGmvIetEJgk1IdNSCfb9qAkbA
2DgfyjbzFHdnb0aYiFMRcOi41DCP8vWAjheYmsSqBiKANlH8odkcxmNxyxxMgc2PMeGyGNDcPWx2
CHxYXZ5Gy5wGT2dksUz8cQJZRucGqoGP6cjuovvHlBTwmuUL/jGzg9e9RAKxKzaepgavGp9CdvwE
HZhyQpsVKceqpGpfKhbEsX6YbewXE92pbPx2RXEgtbxeHAwXj0gub7t+i50NO/nYh+MBZsYVKiWx
Rd+NCRjIHO7f5ba4ne+lJ2ItMnKXbdulHF4MdN0o9Au1H647VcRrTcn/K7yR2tFHsf89hj/TLfoq
jtOCBcM+NZ/QRbytOvKNpTgw5XjSG86Cu2JhyH8vdMVmljv6MVdbmtp4k44nZMI1rB5f9Pnib+jj
KAUowkfKh1lmPkB+qFWsEslSF2dG3j3N6quUFQam9nrntGBYaol9nzIG4BBspGxpAvmIOR44t9UY
BuarySCVQOF6eXVI79BaH4GoJOMnC/YdTcIISLEe07qw+41rQoYeGQ8A9S+yx+3sM0EYMsbQ/roe
ZQQ/+7J7WovcX7MGanCtAJ8X0SiEjKH1yflEVDSV79YW9ukztV9YbWIOEX4NwT2zjJYD1sPwgP7+
FkJG502NVjP+hDaaPm8RwGeA20umpW33Wp1rhjy7cAPJW0b+tl0+yMqO9CAdIjxFeMzRlBJlsuD1
2AZibz3YIk3GF6dW5CDj3RaYcm2Xza/fb32M4/tpK8GMRTwsQ88AROiHdOzem3k5pgAzHIfFx1FM
7WikgW4ZDBZpjbPRe0wXHhKymG3dbiqFrrf5FDglfC9TVFoO8zitGcc3V7hvKpUbs70Xs0oN+XXK
hbALC5MuBieRCGCh0ghsHcrryeauHwit1ykkqUy0TO+07IRs4I69+dRZ9u/8SAY2byl9ftcq13Nw
VmB4lbHyZ0qUf+X/8kWT/YRWM/Irt1xz68G35yieRP4KcN/5Siib2P4MiNpR+kHSFHf2PS7hgvCj
fKipsMXklgDZTxLaSHtlp5qKRpkkShY1IxWRcCjo++rsTgcRuFc4Wv3sibnQQiKjKl3l7bk3WCui
+Thisw7wi2Xj97MA5jerI47wXJBaNIb3epkMYDepNwWOZ0FKh9dYr2L6dJ2/A/mvESEWSuij7wnx
h0wbxhaE61zB85yI1efgX6wWrKwGeznAi9gKoZB4vIOkjZScSzvqahsDJLYD9ejKlQo5/rVl5Fbk
thJTyeCIVz7kyIDrFcQLyg2sxQH3sx9Edl6InMaR59odtikv6lUYItG7aSm8DMQxS0u8zdornH5Z
76wEISDtdIC4KXo6tl0zY9pF845Kwqmhs069qc24oO+buZk/nJQvzfiVZLMpD4YTv7GRksi/nTpx
pGSzXLVpgW+oKnGJtEnx02CHMUdeF8DwKqiXtZOMegtnIsUfBnmjFfzihOtJJsBV+KLjJIKZlkGO
5cvAcbTDPadif0SaukXbGmy9t8kHFC6C87CsYyGdHTOEoW7XNPP/Hry138WlRrCmjMG2eUABbSYB
dV2qGhzBF2+svwH4Wq9RkIFKrCglvy2ocu7O+OHnKpriHOBuhTfqs9GnsCX1gjR0X34uQvYZD1JQ
EmC3oco5Vp7fUtwMlXwzCew3voEBBpKOXY5m6lrjeZAyMTGKeIv6YpC7cTXl0uFTfPk3OCJFOiTK
2deHUCxvmZ4z72DjptJZ7HAXNiEbn4+4x8xhTC+TjoE9uoRU0frANkBPJXCd6+BX0kJzZvY1aX+a
CIJF+87I2nVGbx+uYmS0vKqGD5GKxTHNy2jp3aeib4YlHu0tdvsJsmvEpMAbr7nyn9P6G3hR7WrT
HY1GjtUHBpAlpDRPbrb+Cv8eb8G9pmgrXst3Vx9IHwee1gsNb8AMKoxEbjnc0DmmWU9pys1HX/7K
FTObh5eivohwElIAh4rf/xTAAXJTZYa1L5NXe3PgSxTRtrrokdlf9iCMB1ddrC3cRjJXGCMILPC+
RRmYfbYXuZWGgs4TUJQUAd5SNYvTDkEmfjIHu6m+UzqvRD5iVsHtWl68P85j6P6TUPEZcFDF6o8N
IYqkovWmBAnSPs4t7LqtLKF5orlbLnXMFg9PogCs+uFjTMYzQpgBlPwDxYOJkIDOZ4duywXKNRdD
6IbJ/5ET57apCZzmXiHo9OoMx26CAp6MBUvdOZ4O3Vx2+4mA6tKzaWhCZLNeR3XisHSJs5W5l1v6
IH908zMUNSH41BydF+wrLQ3j6UgGrLlZKCpK788RRDoYXlXhEzTtoZRHdCRB+9eOD6OlWJXfsn2g
Mi5HCzZH9Unru+oO303yj2qoc5sY2siSN30jE7PO5HZudlDwUVmMCRjFBQRT2yG+wqUxHqzqfyW+
iiB79g7Lj322q8QZ+LqqVs6ZGpMsMuBNejvFq7aPRu6IDXErGUwwE84kVsplVfk622j7CEpGwye6
yGMDtnskk+W3/DhZUeDPASgaJVWCrhUMWEMXyEsDrGa9x7izVAukHWwDaP79D5UUoxEhA2Z0ZFoB
ry3ODqgyXVNhDc+1y6nD4fNQ6Z21RUfVLO501ThQU9q4XX9ONm8UZpDYhC6/kzsVpk8/+3q5oN7n
7lLIZ5gtnDgtPkeyE3hsh2ATxgmBOXpLPwN68yIHRvl3a6Yqj0lnNEY9Q70CIgYpXNC47W3QUOd0
hmyd8TPZzGI1qjCfpRax+YL4SPK3od3c0Cd3jUAfQNnjyab4Yol5kLkL+ehPw7knjZPs8Knd0QPc
rNEcyoRD/Bk0IQtrvIC4s2qnbLopJ9dLH3uH/jjUmh9yKiUrvk4q5vhMWoztAiIJ1XsdPWvHx2Wk
ovQi74PncAMpsfF5UMNUXNvexJaruy4KQRwC0d2g0fZpKQvW2/QlIx2t/39Bmio1jyLRPD1WiZTn
xbOFCswEHrV5wc+BLuy6skyZqe3K7Mq1Oo0FJ0s805aWbbf8qNs5oqo35TyMmJM3DUONGqxEe580
SVmHN5aMQ/gniPmQJ4sUdGrpKTxJVjhgBNcketjVV76HrgpX4wSZI3SqiP9HSXnwB9KyD9bmvn95
Bj2OEtS4Vag3oRTmMm/6srY8b80NTD4H5eKES62+2jPMZYQzd809Puy6CaA2yyheFGQwdnvgEdTi
QXUFb0ia3GpuCTHQ+3li53GpeMcJ0oko1dJKkPBtXyraL+J5ueLP4qkFoQNbeTeH3dAowcv6UZKG
oOfsEVdNYVLyFIR6IR+Ifckdn0T7PeIq3EAp0xruGDZ2jzI9uxOOrPLnOa17yGvm5LC8eAitHV6f
haPPHCc4ut5I8qepGxH8p9h5bkHPm57F1M2kWFVYa3OpBntOE+9tI7OJkNgXqAc2ip8RcVDkm0j0
X8hsXC/oA0qwENoRlNI3y5A1lQCr0ewGZvr1HJT94gstm1DJrwyE8HmxZRKrKR9Y+qH900OF0QAM
1dxrUimBzkHe4RvxwtZ78MBStxKb4aYw5cxg5tiHz0rKkpEiT0WlzeL7n5WN5jlKxJR4zaybNRZA
dI3pc+/ZDPwe6i8T0oGBG6MenxcsWhRa4VJupixro7A1rJyK74slEaOwjMZpjv8IyhJh74A/xphz
gFL5irgDRqnAxpEIF1IIq5ne9J0RU+gzPBDsR/xFE+X8eA90p0dHSGJQ7NNXW/4tOoUr4qOMGTXu
KKiqXBCCVKyPas9uElImQABrIlHvBbZssFChxi2gJDKCAhq78TapCku/6dgPyqWiJdtkLK+36ga7
M8oYZmE7bvjdlqVlUicyFAgqHAcGNiI+WxJdc8tNo3qy/gCwfvcFkuRuspOc0JXJpwgqnrh8y8cx
3QRtWZjHb+iDYAOt0V0qDwdo6gYVxpAPxR50WWuPCnpl5PWwH4NtbnCfQ8BCE4JkZvczWzcTxs0X
rz07h0UnYnS/qTZNxOWiYzaqnMkw4IWh+qlapHES1UTaKVv6oP485JLa5JfVrj8fBeBpvN/JRGQq
L0iWmugaglRJXwsKsfObxC4JytTyfW1VVwFN70fHEAHTp5kC7efVGwOobHgMgEdEA9uWRzkeNOXV
KQMlFG6HHuu2Xujc3oTyIu5lu+Oy9cNz57Zv2LEjmbfpVjjt8dDFNv8lC4jLmeO5u5BYtpk0NFer
2vhSa4+ypZs048h4WPSgKtIGy1SxYiNIcAlL78pDAI6G9rP6XBw+TxA+Kr4LykTvT+7spks3+bS+
Kny2nZMM5a4/A3YZ+30ZvlRV9gvrb/4Jr7J4kQ1N6t3BAN56WhbStxZ3fyEJNQZEXbVUDtxilvZR
rwcQX7biJS5IjHRUMz4wl12GBFGmz499g69vVxeJmLvLeYb8MQFK40AJAr0O+ojArrcMkImAs/hw
I6aDDJ5pHcB5NI1lHZiooij/Owq7F+EUjAXwUk9XKe1bt1ICZXVBF/0dUNxKu/dhSne/nDOjjaOa
etmw0NkjvixOfdwLYJmGXAaMRCIJkJ5CEcwCRTUIC1ofPH1jFt2lpwXCQU0y+X/ZnUH16G8LJ5qX
p/z+k6617PM+twj9X6WGSguLufiYbfU14KcyEocJ9GkUFxwPVMQH/6u3wbwlJff4jgGIm0spHAyk
C0sdCuXMBlTx5Cv8ZLtFO5fDXcuXfQA2wSO9pqZ7ROjFIhCYAVbrhT2xT0KJxlgffojnxvJWyw1w
IW1I8u9qeILd7+MnUGZge17G8lIQIWCZgoaBb+i1A6HNUA+D3RdAZX9f2GeLZ6s2SBU+ZS4PBjgI
yQUx36TVtGVgzOVaYmAMWpQnQn0ioWDbEkiwiIyeA3k32kXmhnjLhgd22LP5KmH+AFQrBPTRtONf
TrAmMkthJdpyukEhAzvhqEBKHfP2eP1APeHzcaHtZVE4LxSgKlToOn84SdX88yihIbuhBLFns6a4
BYENYFDK2leixZWaAC81vEZeKI9N09gUkaMW/kwqTCQJxCxzGS/yEaDWjl7qHBPHrW1hkBJa3Ksw
CBjK27gX1bf8KrY4F7/UmOn65WSywCkUwT8pxYhploQ1/6LduHoGJVxmtpnpMqik5UdOBYVCQvI8
gx8RbhmtePqVSp6crA53RC+xmAD58rNpHFO78oGGA2EBSR66pl/l8OgN5+gAVI8xFlxidI7efEa3
me+TLNZH3nQRx2tLmil7kCmHf/5+8mw39qs0WeIRGrhqZ4Tr5sa+gC7NlgWpihrOrWucLF45mhYG
oRvHKwq0qt+mXtdx80II/PW4vhbQo0MgcRaXsGdAnaujBg7JC4hgL4VBToAAxwfgoTSQhH5rnNQk
7MoxQ6jgLc9/jqwhWdxaHWjjOeGljecvqbRyhfkTZGk4HTfqyh9YUVU6i3T7Qsxw7CpVJW20GXEQ
5P52qscauvOeSlG1Rnqxla/Eb751x8nKf12nvJTHL7rawIaL1QkNqZi4YnIlpZELaMrMXGLCY6do
E6862r92gAr6rzj572xFZ8xiB6C5JsAzKhdQQSRM/gZV3z4XVO/d3bZcs5gLDLlXtfnzAofHIuFe
6uvNL+JOoDMmXpt1yDNIGJBKrMEYAerexp8UplBkXUv1ODain0syWGibQ9cbfwX09ePIWzDg2lef
ge81sBt5T+xz+sxzC4bNU0kyVVbAJRYlLyZwWDX722wlXE6xhxqhixFDMpeXvkfybhX4MQbQj0OP
ljrMr36RkV1sQb+C+5aSDn+WeSMQ3PVS7bS92HGTgl5n4IejLXrF5QITu61sQiDCILzkpP79QE1w
TZ4ruVCYm3DCAdbHSlxVYEgF7wUgroH9OO3aFR2ZN16dujy4I1zBIyg2LckVKSLIIeq7mV1MA3hW
GQadhPnjvOAeXyb0OeZTfr3spwMFt7fmEqixGGL0Aj3W1OILRJJ4VgELIIsOcdp/yZ8E75YGQIgx
x0nYmjoVzF9ln7Y5aQm+WC6RSZaQlaqMWgy2ZNzptJ6i7YgTjuQBxTi7M0RV+o9qLq+HnnGTeVI2
Nf4pI7q29QdlFdtNMZrxT+XleGaxd6nflKwb3oE74WK7szNEryNkgkJzFZpqnAHFALAtvBeIHJMi
0fnhIeO9qYOq+zQZpE4JfZwQUij0fcCULqwCN1ZG77uzvf1Qmso5jPBOOhd08yY8Qsmyz9JMC+eR
ulfU2athcYb8Oe8o34SBV1+0nuhTc1W3PyFlFGykuLfqAJTOpGGn5w7ExOsSCaNnex0K6hrDFdZu
m4ZbY0KdGmvZdX24DsmKbmu57qkoUN0GWSFP99Bb+ChVXdea0G8JfkjB2RIsI+GgfOkPzvH/ylU1
psEm1K8b89fkAcWdvriqhEX4b0G6KL/DjQk7ir7C7FKTr8GL8+AcWbu2YdRLQ79VKbeag4VpWiug
TIH9qx2OLfKVAaf9Ev5mUe4P5d/CnXMlM9duOm3yd6KAszKPSI2DRlBVPL8K7TEb/lx6OhXDn3ch
3L/ulGmIEJjJKx85q8wHPtVowQDn0f10U7FVDaK4PrTtoKhAQjyh54nGZriAf2fckGXUx+2OWrwT
/zQ9kzjY9eXAyFOcgpZ6+gSYrNDbLaXaBKW8mCQJBOdNoCw48PmjyZ72u1BjpDnmcpyYssC4RAaJ
WA4tTIv7ItoWBpvIPVzlCwpivpnU7anuFe0QEvpEhd6eE9pIqQyJsNo+V3+gg3rMAeZz340jH/Wy
5peZcXBDrY3CCWE6lBPTHRiprhnA34QMBLXMo3akwAsaz/0lUAbGLCfIreRmr+eSLFTdl1rN+yvt
f62/crXf0EKqfQ2o+pwvEvU8zo6QT/EsKprOF6HyI6iir1KNxr4kFsb3+BEk9CdHn7/kWMvr+HGK
41efxr0+sHz5iKSI2i5rggMBmmQd8xQxpGWTa9atU0ttN0llq2PO/4gQ3FItQS5DkGQ68gVEXj7m
9tGOo3I7+JkuenDakLQSvxo3QymjZo52+x9gEsm/yNw/tz68C5SSOxTMP/5WgDhxOciV1HFbFXal
Ds0EVZah09FIVqiXAsIgJRZ+yeNMGcZKsaKsUA/mmQ1uidddNtfx3r+1aSNzRRIBOklUX5dvQLi3
DaH3gNOCS8tGnttPGy2o5cLnxl7LccCj1m9koJCMoJ8SppAVi2CE9fFb0zp3fAOg2LywvIrNSTJ9
jHwn1HTyzMmIaGrYMmAwnZ4jxqySoBOAAb8Arhj62KTADz41S9i7V7p4IZlh3qRi8ujdwXb3TOhr
/yzscJzaURvryhptAMRzX5h0vMygprJBEI+ED2fUucXyuJOkv2hp8mkxOaL5fOhRedahrw4gDqJo
FIts1Jv6nijkr5TQh0h2SgamaJZ40qPoF3JbLdU1ZqpcGmxwq0cEp8vlDT0KEzxRRtLFWDA4Jzx1
Y1LjCo2TLfMSJGybmU6gJuaoTkNhHyob9gAqZMVe4p+fTVBiATnquqDehadoWI1eZZFIzOBtIm2N
mv4mJjgxJYhARDwliZ2Fu2njeFESaRRGg/becvnZlyWGWiFL2V83X6tH1BgrA90byvluhnKvaopj
iLPFi/rkAJCqBTD2FIoM/A0J87+GJrL2rvBHPlhGDwJ6Bue9S8wMLPz1YZP1YMp3I/5m+GiBOBJt
HIEDcDAPkbSA7GlgdB4DjNLa5COo1cKo91NbrDbgvm1QlEq9CCH9XP6+UGS6voETDPWj/F0j9ZvF
zJgcrlZ4e4DrBdueexha7/wN0VLFF9l9MCzAHBs/dXI/5CU7ewiZeryrLPSelKJ3CJhp0r9m20Qy
Sf2CbRYJbUQmJAXTtdc3ZBy7op8eV1SgfwMLh3blfW+JPoJcgjJEE4jW7QE4kUAvnbrW2RXHLjXs
sFrHoVwSvWZcX7AXo34d9rGJ6dbpOs73QgH9n6p673puOAUYLTyy9TNeaxEwMTJw4IGogk2kYWQd
atX2maZRrKTbunJGr+1QLKvebtcujMxeowh8F/KimYt7Fxh44WoprbgXMlchsYMA1CDHHE+s5On7
oE7UqXVZeUBjh2R4k3v4Ohc9PIaySa6x2jzltK3Dq+ZC7dxt4t9zuDF03O6dD2DQI2fFRWSLQFep
hcChsilOqZHyMwaqew8L/OH+h9ES9YxzNGBbU4HRSg0gEXbaY+I/SgnqY90ZlXMQ7r4tRu8o1F9o
08jK9/EpKJBlQjWIJZWZiftvS/zIHcQJIn4DrbqpZr/o64wHty/3ldcvAPZFWq9z1gRDMPSubBj3
GYXh1oerHHx39l0x/0RvhTUC3FvfEPmFau7B9Zq+st4tCvH/1cFs2+BHS+cAgzs0CKG626N2o70w
kEYkzVgjCt59DtELEnsYyVY6lY6/GTbkozz25wOhOGe7KOcfZmMDws0ImQ9r27IcZvpqqf5BnP1z
NIYsFOMihByw/z+jMB/SG4TAztmaxjKAZfUuSfoGQtOa9ZXVXlXoP87EDptDxYr1y38zyKkBgcHk
Nkx5jiCWcXLlj35osDJGOAJnK0/c+qTjStEqVlCwCKMz1Zk7glUzKUxKC0dOVfwHB6DtX8AYM7H+
kYLdvFfw+b2XpY1o5NnHbiNPGXLJDNwxhtwFbdzkXqo6ztiF7lFY4cwR8dQEUMFifg7MquUqk9VC
Vc7QAu8kQbL2VIZRV4i++t9dBE9G1bcM0ngGJIvLkyTfq2AWCJovEyhu3wPMaHeuIKH7dc1TrUIe
q/zPV7GYu4G10w0G6C6ds4VB5khHP7FMPiJGZ1J40FxcPtWj9Mt2la7vbm5IgnRAcQ9Z48kb/bJ2
pUc6DFAxsAO33jwTici80XGxOeyYswUEy0VCk6Tp+kmGTB0ZbYAYBXmG7plvmrQ1pON+oWQozlLf
ZZapuly7amBgncfW2gLwijQSuJHhHuzeK1Dg1hD1XC8sAOflnSGjRV85XGYtRBLF6mIzKXt/baXm
KTtkHORJOR3T134d3lI34gTCD1JRriLA74SlY4TF3zV3R8VKT+vm2GnSdVhAMCYzkNMnjSM0Ch9a
QmfzDpnlzCrXv32om1X0P9Pc37s6MxLZg3mWsyNyN+sf3tUgoyuFn6b3CISyCeqItWg0/eyeSiTZ
hY3+mtOMgonbsS5UEXJNvNMO772PSJk1B9mzuPiuKuwpobH6Fi9PSfcNJnZHEUK37jS4ib2ezecp
tQHz2jkhJ9wmjw1v0Rh0csComY7S8aRD/h5W1GygTVMcIIC6E8turSLUVAtC8wR5F1eYiUxeXNTd
66FT/CPpgvjZgsMEqDF5Fu6EOwBJ/RthVaJtyD658En7oYd9HiZrOhodIX4QQ4s9nXDwfpk5x3dX
HwW3YILgeP1Tvx3rJmfJstjlFKimze7vGYpvGJwZyAXHgFRcWMiaANKSp8ar5K2zTQX0jl14GRkA
LzI03gQNueYWHYJc5UaF8/FMvTz6Ro+hoVBNxKDLjxgMXhum5YEK0+kj8JGtXaOlLteCjCezLdLu
2DLXja8cdMLdKKsnLxoDT2+lTQyEwWFjhe7twzcVVrcaJEQgZtkEuGky95lTV0dzaTX+dnBLwt6L
CnvKCKAjAuHRSWOqrK9Xh8lFYXsUEU56GotpqDMsClqzLrnuozNIeex4CidEeOEF2U5udziED+PG
zRVumwEHUZqgqQjwHOoG91UggIdzv13KH3SP0ZgN7/NxbXdrUNkvJOQpHIUuqKLcJamkpMEu3FeR
4I7HKGJ/6j6X8hRDPyRxDAABPKvqOxN3tbxQRq24r1UmAhq+InDl1+8tuwrTPx+ryFPxgZTu1kJL
KdFGJOFUueqg7O/m55i3Auvd/kzPNQoRjS9eMALtFl5PfyEn2cMAwyJxyLaL+MgoeUTQdpmfayc2
ABYqARraXoK9bDZcS0UfYs7NX/S/OxRVermwtQ1bQygOx2ArgH61Us6jGDAYoj3QgZmet11mHbwS
VXFRb64hbLlaSTmvns14fAWsIfh7KwbrZWNamGT+5HtkzPSlBCh6maREeKPd0fTEMLNVqi6wamp/
AE8SJvEkQS6wtYGvHxGpLrfM61dIRUKQFKiFFQFBpisOCh3t35sIEoF1TYbPT7Mb58P8rOZdDFCY
gUCFqssGJvFcAWf+Ur/Ij8HYfkt0jliM+tvpbwfTBqkzIb3Nk+aVcvdidT/n4hAUFWNqH709utPC
jWRA4IUrdQa6GapsUKF7myF/rS2EhN8WMt6H1j1q5Lv5QEl4cUk4cX664z/4jjSfQ2mXdhSFvviK
m3wmh6HHatNJ+Aal1zIoqQfLLZCG5DsBZR8S8R1PQLNpEKlpKwYyCoPRinwgLPxi1ELmRPv9Xa1o
wM2iZbQebYFKmjuCxGgRqykqhoacVNSFcuIIKfX8M94l6xi1UJAKfT7fNcUuLVISu2gZ6dA54D41
GBkvVTd8zIb4KGbTlpjZRDzMgKTABdlVHcyjIQc7fnB0aqrOPxWiG8wG7JbjxinWeDKbSyhsVAdc
xpU/NDbP+uz9piv+KNIfBLnZmX0fshOok0mnoyL0ogt0HRoKtc0W0aVF2qb4/n8nmtJ+pcEzmhk6
kfaii7Qct+2SaZUwNIyBBAXMaVy09Kz9v/UwzD4Ui+ou6b1+MXq+7odHaJQ5GnGeieZkSljvPwgt
BRHQhSGM78cKhK5fSSfNk7Iu3rFdxcnxMlzSwNbs2VPX/gh9N4F1ujEk5IBT9XALeapn5qrQLHrD
j9Fd+4KDx8fvPtg4JyBBroYs/tyA5F7LCDifJqDbJr//RKnqSciW1jTliN4u4RfAFLV22POxFQvh
lR/3udaOvHw+YovEMPjEkwoM2T5GlJ0l9Y/0fO780HUuWsEHf2DIKA7tQXcSx+I2i7qtz2MBNF4y
UdF/Ek0bwpB9AD2z/yLFJKrgLINqGjV131RuFCuQ8zqBb0ApF1RrYbgg+TE8E0+krSHG8n2dVlOl
vKrdP/Hv6do6ZbW08yfL8nQbHrSUaVzs6yxEOPmRYiJ2EvC7kEeVy3BNRlnuSaiu4FTUJok/Oqat
v23GS5buJml8n4KeS8LolWDi3tziKyS2wE6o5OMoM41VsyHwKgR73o0r3nzWx0qsjbp8aZXLaCFf
AGFTxWTr4xZmqhEQOjXTLGgU0oCoqmmI3SlEld3cXptMiWL3jMSqcXIm8f6F26UnOxQESzs4SptS
LViDIQbVhDXzl8cfWPGGKXQdZv4/jS12GaIDr854ZfW9tQPHoUffF6hgS7V6iKxgfv6sUvT7sI73
1xMJuvWy/+aT3iKQ0xWcrFMxMo1JwSFqqaBpG8RGGd5rXBfqN/ddVfgBpaA8mDVEfM/nDEFNDzSQ
iQNSBXpzQTapQoJJKGNJJeeiCJ6rjSf0kMpTruWIt+388zS2Ckd+NCzVoDS/TpuqvwqG1MdRrR80
ug9LGzGrrbqGPXD2jnBrFqTG8LAGCcj036wTqVBK5gmtN8Z9tRHrA8r3Iag+FFW0WbTHCH+sNyQ3
wVN8zLNyT0Go6WOPDOgPrtQqmskjIKMxR6BN1liHri2rNkMpcBqlJZIgo+irWcq/lZZKqQMKYeYg
N7ggkoB5BYqOcSoE8CiVgrXoTISol/NDHIClpBrZVmMt2C6vESje8nVmyFhuLEDRt7hVd+hbWH7h
g+bAxhfXKFbIkCsUkoy+QO5/uHpsZ+M3JAe568sd234LRm9oEoFjdTBMBPZuG7++kvFRBBpQG5/y
KLyTbh6A6gQb4JQPADeyiFcDpJBelLNBbOdUzN0V6keoiMb7CfiUXbaR57qoyRb0EuwC//lu3Gmw
u/xHrotNed8m/lfhv/sI4D6h713V96hO8jVY5A9bYDo+X661E3L8rwZljPhBWYCun0rbhX0QvbDO
WFPmX7iU4hPuBXOzs2fTO8bC62PapmsvqaO9Kpl6xYfYqmT21lWC2E4DJK5o9tVCFW2QDZvJNfGw
W/q95owgFjLMMrrY1r9d61x4FaS4QHqk0X+hAiqU13BVXVb0Y0xX0CkIw3KOrsDdkBq4j3JqGUcP
7gdVJFQwWyF0RmCaWGKO1HEWCJ+dh1vjjoeMVbGmlpVNdCJBwY/JZd8feY73RWEYZD0bKqOzZtDH
iEGl8/0UvjEQr/Nrp2AdQHrwGoIRbps1nuTlRqQWrbYtVw6tjes0kEJ3nduVFTlq+xVT0wzHUl7Z
7vab6Qc/5pfhV2YMLQW8ZJ9+PoElJl9T1+hgfpt7LeEaVfzD29J0xab+7F6mgNqW+39wGqMCu/Gy
bZ2CbD13QjCI2mouFXJsteBbGQcRZ+xPpvWewLKvOwMjTRDGwXBzRIPxrkmQMoqzWqU8F8rdNCUV
hUA7BmRLamKrwKEifqupFofxF05HybCq9K6CUENJxHF7jXj3YihS1ktCtKM6iiZBZjZZSMctjyWw
+nhaFLGXR2m+Ec3XGKhgTPIqum6OdYjVXA2SpaQZjI25s1VvjNfrp1ckmg9Vk0zz+4mBdjGE7TXo
sIaLQiCUYre4pe2Dz3C0OBLctpF7n4OniZXBXC/fJYdGO6ZYCPj3+AjvuFzE5jUGlCRiAX1m5Rqd
7k0sddl1sOYtyo+owJTcadcnjD8T3UCZfRCYufECvsNoq9yhid232z8rQSWQL2cIuof/7abPQ05a
05V86q7MPDHtH+X+jFBondUMVZxsS83hbmJ+Od+3Z61S+yhsw6XSFTBHUpqRRMx0TiNHyRN9dJh/
79Vk4poFPXbe/div/x4wq+J2/Oy9AgaXB2m2BGimlfuFRh3S4Hbg7KX6tnM4rYkdgPSvRAV2xgFC
GzwQCbNMhrHniFQhavjH5DJLVTxw7TfHYOfXu+0HSZSmrihs9eKGF/o6od7rLLswXGPGwrdn/1Qi
JO6ylojUxwCjgra3mGp5NEK4yq1PxrA62+4psitDzxZcfqHlEvkvG6d2Ira8lea03nEJ93275BW6
hjiX9chuE4YAyI1Pr2JOQ+UgR2XVaD2P9Cun3tJz20fDVPYBerVhN4f3M++KJi4Yg9o73Xdfjy9f
yxca2ixqedMu3YZ31uegeU5EDgjd/gqQkhdmjGET4HVsrqRkezPUJhe76BTQH7hQ3UhA3BWy7L8L
lbD8tP4Qnxr6zV5ZwLzqgcjO4F95apJioSrbKHDl1sw/T1Hv/Y85+fxqGm6aasIcV8O6OwMd+B+5
MWWmdl2QIwhd8gTu6yN5AL3JOkYDllCQJSOAVc9tvq8DgZSQ7Wd7wmsXF6DaJ720f797jjzq8gGg
Fyz7FLS23Dnu7lX75JE9SBMTEO6KsCKpIjAgDL0sRVRDU5o+GNpvutqtDF06BuIAZZyrmm3d1vQ4
sfIwrch2w+RAJATMC+7idqfu8EungXZei9PuazzWKaZPCC6lZLcvNtxtRlV0QfeC9U+1xf6lTBX1
rTfJrRG1Rn71ntVbApzvFAJ0pONUR9BCuXVfGuqJl1orQNdbzwy99LF+rSY3aSwvxYrIC4xdz5bu
zHmDqv4k9KOb25D7qZ1WdIsxjWJaAnx02QEdkVdhK0pTy1BucgJM3eQVCH81bBXhGotrhQ5Hd+8V
u5Tj6sFScFnRd7VlC/lQ9YbPG21YC+FVparWasXEajV71B1x+rjh/ChM83E5D56EBDdOivpkZ/Lw
4mE8V70gbi9dfEgQhnfyW4z6UIiZ9gMKpWtAePoXoJybaUP0/b4um/p8U/w3Mhgfa9AcsT2cFbn3
LzMNt9Lxw57e69N0qS4i+n99ZF4F0NZg1simhZ+KWWZ8EmIWtB+hO85ltYo1RXNwFJaYXEvvwgKC
QVxee+hlRbleRKS4Azm3Lp0Ni/VyipReb98IF6bRk2DDdPNTN5WNrF0AdBQdddawfJFZvaXeKy+B
njiLotyJ6nbv46xZpQgjpFROaQwOeCiIVJ4hlCcM0aSptxn6WtjUQSTgyR4dgSHmBBJpx/LceCdk
DLHl8OUQtfntv93yEKEmQcc/Xwl3Xd4f1igQGbyOUV8glaIV9ic9GZf/xrCfvBaziCBuCtIq36HR
77khANijlVrMIXJHY6jYwuHYP8+iRKPjB8K+w7MViwTxXT7/v0TkRKJuMafWtCLQs25wtrgCZI4Z
4pj9aE5gX3U0Dqa3E2Gge6ZHBPjn9wRzx69GMHqkeUsuSwj9PTGmf56VJF0l8bA8q5/QCmkERnA7
jM9C4Di7P0Ug4HAJL12wYhw4fDgURF3DdkmHu0AB0hiNGW8VQ6/V/BGVqBajlUhKsHdsGZyelOx2
GvgMvZoIYf0ka7x7MPHCtRLTIAiBjhINz3pkz7yxy78J7nXwYv5xHiS1mHGcJs8RgonFxZQarTxn
zq0tGmZSYVaxrsJZmQPHlAmFs7Gkc9q0tY46Ne/VybUR4cHzyBToVYUYWW2E1Zg+Gs6hhy5kBaW5
uY2XmJvdLhTfe7rsCy5Ot47ntpGRb3wmr/kmmWDV/6lvN2i6vBZmvWpqS7c3mF0oKM1RipvC1Gnu
VV7xnFTD8hYjWzRrYy7n0ZChqGIlioHBHxmd6R18EMPYSJgBnMaOzSSzN2D4RNP8AoXk+Mjd71yB
KJW2bRcauXRzJN9f56Y+V/m384/akPOWcxcWgxXuzMBJU9FHDqOkWjkgoyIwBExVMkIZv9/W6+5f
ia9KgTgdT+Gvcfm7nN3SvlO8AJNtEtriL2YE0d3jaiHoMqz0XUo9RHnE/R0vtShUA03s6soTkpyB
y4XlE6ZKVKjhcYNtggksdt5hpJvv/miH4C6jALa0gq4Y58TBL7EDIS5mkHLN7eYIBDjb9WR1IE5s
G13X3LId/GoKqKSBdrkQv/M4NBdomNQP3K5eX0Zj7bM0gg02wVim8M/cXfcGtC0CG7eoChQ+ll2h
Kg/vRecbH/esz4sfk29AvJQLUAXOXLgwdPL5DSGV/t6BX12WpJpWbf5/jcTegkUQXHWhBNfjKKJe
PohvzbAwsCZacT5l+AQV6IRejushs+h65Rbjwv2YLbHwll4zWkcyuWHR4La4JUXCdvQdoYd2FVxB
kpPzc/6RMDXx6iUoaY4rOlGOn0dqb19Qf3hnvu2QyVwJ5U++CVzHWD+VrEtSOR9NlDmoqipClUW2
d5wcS2a/RLoV9Ze9XvKL3IKsZA3OFDZWSwTRSsGmXDmuilFfyGTkR4FKAjWmKAoT8FzrPdMofs8E
wbyTpy33ZEB4Cxe/mkWbCbIJFadpnNlTaXna93LbFgsMm72+lz5XHy8buQ5H3qSRZBxlEpFFnAZW
LIk1nTbWA5CqaYMJP4z7RZpYU/T0Ne9LJBa3Vn/mbJRG9gVIJMhzd+mSRhjBgEtoeHwxZ9VoYZk6
eBKc41NMZ2rJD1RM0IXSES/YTSjmSDrU9jurxekTM6TblaFk69Sg4/A2mJiSYpw0XgWakAAfsr7Y
bD5v13Ip1aNVQ59uV44FLXPysfN4RHOm/7VEm0K9sMSb5CFLSDQjwR4IMsUHV8z/HJpej9j95YOR
ZiLKhrMwXUPl0oqznCpSILc1ZoFq6LvGQW8wk7clNcT0GONdfV8yCFnfe4vxqmTXRUEMWA7P7oFP
3n5ooeaey3m3vY0s1AcjDbs5ETrYGR8hzQVRZ39dRDDrq/ud/rnlQnRXWITmlTZOyww9cptwm5BA
Vn4mkyG7us3jPJ9HaZ9zTsRibGef+wVkY8vPF+IeOWDmCHG81V823S7cRLhVSig41uXwMzdX7w9J
4d1pNkogsXDtoS8vbg4y8iJamcIqLZ28qVOHr2fR04n1ccNSu7tlUvDAxFsVNhaP7d2qShEcYlaP
SaxsY6JbZSS49YVBY5yVzKtzH1G5QsLE/pwhi4RzR8hIkO5gQ0aW9XXF8sjkWkJShr85xO4OIkoB
KvLHN/FfbHoFNFcjjT3ZPDjWYNkMIXUaVvcyLjzpLoGmqbbdFSC2rveAMavMfpBhFfyCM7F9aD8m
4kJ6yiJTQO3CrI3RW0h/ijRzo5ca6aodz6shDZH9EOdtOwB7LvGVNGZs0Zu3JF/odm7PPWmWxghi
f6Rnzb9yLn0bB+10NUXamQ42oI1GuTuIRaSik/nuFlUsYaWGH3px5vuYc9V5txk7zIwLmwGtbpdD
fmPNgJK2SZROkPep3jN/7QePTJC0btwW51SCFCDf88k8+uQOtQANhz2Vp1Fcln+0pZ+MQhkGp6gc
QEedLkaY9rfEyvGzkkqvZ4pDDYwP8QBWaBDP0secJH1HCBHMqoPnwmDDP23Vz6IQ0vKIjslBZ5m/
A1+TIAfbvX2lqdGpKxrdhq5YZxNa9YUMqPlWEo0KThYutWb1OBuJfQN6J68Nwpt1hlLYBrG82yDu
Ivkn2DUUq3SIk2AVEZ4CmAbCA7QhMELpWKA2pGXweUuKAcVc8YOM4siFYiVId+xpBymoIepii4Ut
nRMgclC3G9we9N+00cy6cme8a6mQDK4bIb6nAAyuf9gIUvB/DXak+T8gK5YRDqusmRr/0a8KsP5x
vV/QINZR1ng5sgn+P46ORICv87m8OmwBNCSMSQ4FhlJdX0EdcdmwXTLZwOfnJNuA3QpzKw7c26bb
ecjGgmOIhoRkrD4ajKkFHX0JmzbI/Xu+kvHYcESxO+6uR7VxG4x+YIwScQuIeT76NEdmz0kOpYn+
Ph9Z4RWsIqCOmQ/ZXSy+td7a31NBO//zjgQ5HoCEXAaxeheXLja7n7OtWyh/Mzemdn5z0BqytY+K
5JsdhK9NLQTGUp/mAer7qj3ana+XxXTXjsC+zKWLAP3uoY1OU4KKG2CMq+HaD9p0Kcx/OL0qLK9t
CdfP4fc2CXgq8OvlVzAn60/guEKtcOHCBDz6st1UThgLwBepywdys/oWPZUZokIyK2G/RA6ExoFC
gDBXxAJlYkkzwHNTo18r3HbsAxD/kgt5Ox+mKrYrEDiuWdI1iD4inS/Qu5CMMN12sM8raaivMnDJ
SqISddOaEeyKDXzskLDlHv3ex0yPFhAy2eKBgfZfuL59qXtKO6HkQFQ1Szl91NOG1t5GTi8x3Lq2
RPhSsnii68Scn7/159wwyaXhqSkpjR321pzxgRBej2WqP8W5BBa4gm3hoUDsWUo4mmUeBBZ2Vob5
XoUup0AVzcYHItMvkQx6PluSgoijfhlcME74C0thxOzrL0cBIFDjLppJMWTnKtyjzyktEJV/n/Ze
WbW8+blWwz8+AvjT3yNK8MYk7mxmk6rKqOhtzgwUXzPou673H8sg2AfdPLOpM9PuIijEirIe7JE2
MNaTod6K2QjrBBKgAqDcYLUtKx3trfSapploNSiPgmOTLyAHMQoPadZ9uIEa5jP0MI0mTDGOK39k
DYJndKaSYytcoAPYEUNbqIpbnVg5DzRdo91iJIzDMFb/o4hcMmU59P9T7NeoD7yM0KsLc8HGwm7D
x29dCyXr4LOsC7/L72/JMAyZbAJazVZciBnvjQU8LTDiaiuUzxqQ4M791T5e73WviooacUFiuCfy
Gx6IPf7No/1JuBegWn/v6sYm/fmmNS3u7N6o894oa/R8ID9lISFILVpCmLqh6v3Cl5oiieiZcR7C
mydOHHcNip2GhpJ5/Kz9XgkDqfG2jdJAnZTcc2YeepI5G4mkeheh9HNTlxjwdTCTcFtOObqZIaxE
lbNAVEay2JFWgNEVAwhYxE94bTZxwsPR4cpMQX3Epn2t4aDzAmN9taxPbAGzOsQtZRamC4/kI50S
TK50DO/9TrLKpXYHLlJcGU3u9iSEzVHNJdZtkltEawphOhWk8I7klR7aHOm8NybFYhq1kUIo7zzO
fcv4tviqolgi/UW6hECRqLBZVt+LjBjSR41bDeElFyikoX1bu3SVOxUDQE1XbYBMfp3aatxngOZv
9QnYFY7waXnfnfbHlUyw4MJRCjE9rsT64xBWHVHfUyRBIr7B6yW6S5uH5l+mDJoRQZv4Jv8obaBr
ephU/sFx2SvHwMRYbQALqYepGQuNFmsrk8cTzmRdUKaYHe89txeEnF1Zerl5sth7Z5CEXWRJgiVe
xtDMQbDev0+iRWh/xdQdlNp7YYmba4Q2oRqOvHXUkqJY7hLa/xVs83QuULy9Xu6OvJHjRqkYiDjV
Pm0w2gHpUA9EScPcxHByY5Yf4eBQSO+TirGAKTXiEDRNBcORcChSOjM0Kx3RLn7sLqVAHTaO1DMI
bmFrbV23n8j0ge3TvOLWO9mRmboZ/lKoZO8Z/AhDbQJKKo4v1Vky5VzQJ8hmZE29M1qmuyxhiZ3o
NMW+A1EbGLGzKZyxofHRkHAbX1AMreIOUEODdT5nzvUJ2K9VLYQGBD5/lWEOtBoss8+P8jGU4nL+
T0JH8YUpT/5Urss59MJeYOIV8iYuI0kksGhPuOGBpRf1b1B/nAS5BdgGVOeMfT1/tnYSLVAEnHOB
f/QpzUdUAJiKyBTWPxHNpp+cEeiENjlKOj+2bjI+v4uc8ZnUPXWW6YBqxknTnmjXAFdy+gq9MHom
yK9cJC+oh0LS21pf4LLiwRqlsLLidZc6y5riSNrqWa9CLstMwQSwL9Zcxb0Aw8HpH/Pzw5FrHAFo
BYMtwl0jbZDZLB6eN5DmgCMNQH11vfBWKE/w6wEwmBBcrBB2tka8bySQ5bXNFaDIsTKRmjocwvY/
JGF119QtYV1vlX1YxACI1MKOvoImgPPDQxSfCK+GdRSb1FfxtlSKZtClxUnJm+TPVwQEd4p58CCR
yonySrOe3K4paiyu7GYmqIglLaxTj6oKCS94UZJ/8/4DxRNJDAN/ztF4psbtPL0L8Go6z+KsWy+Y
t6WFDwAI0mC6sIU3H6k45YfrADxHdx5XFsPX11k11qs03QO2OKqPqYTJNNOProU1sjyygNcQKrMT
5fkvfwgaXaiO5iFR7F5g4ioiVtO9xB613FY9cK4++RfF15nSIY72zBfGvmjiles1MxoKTU07mEyl
S/dIHR7QGPhClpyiadNDPtjNULu3Zdl507N+pSofYAohppzTZu4YbBxmim/QEYISF+NI5ly8rEt3
ubge6x88vNQpeD1sKinXLfiHVNOw+d5CAYj51tqyp6YCpqKwHM1z4+QvvY2uDIzunHO8UxxlkdBa
242fG9t7fdueNyKhCbkKffTjXtaTIm2D0kgcpVOil4npB3ELwdTOp9iRzcSLC7xOGuPRwQ5EQlTg
xyEAPvq81Ck5rXsTrrsJrS6wZwLRth/Fr0HFrAb9DDg1Hqz/nXEEyGdiqkyUeQG8toLdsLcXbDu4
yr1mpHiQIwpECcScy+BkGTqnXZUTXNmjwxv4Q24BwUS9ULlpsb7xPlCdHhvfWHqWYHvwyFpVJpVE
l2w29rVKLFdHopoHHiAxhBpQuSQy512SmDmuBJQmaLIQdEKR2fHCtLDERxqxHUfKAX7tZf7SUGdZ
oEFx7iCxDwxxuNmQvcU18jmHxF6BmKH6uuwtza5tGnWCPeMsQsLqVvfx8FLkjlu4A3lfDHK0wLXJ
F+5xAWJlvkiC8cIQf6dpleyYB38clX3Q4gaMqHCCoAuLuZVueVuur3J2T7xCNHqj95kkz0J6tbJ2
zKicdifa4aKLn2Pepqq5ZOwKvjVLTphoc8n+/X1vt2HYpn6f5pvYQ+hS3YE8zSn0wVWTAN2qxu3D
IgEK5jGXS0jXPkXPAWdGE+YDj0B2IBDEDa1dtIsrvG4A3zWu/ZfXowbAdJtV3qk85MYQvpkvg2Pt
PmTDjIvirAFKWcDMSUtAlfoF1JCpTgQV5358j75Q941Uz4dupjX5W9goUmlnhvIsm7jRe42iXpek
bJsvUw0bNzXCk2vht8nXjeTKxT8kj5rFhJZf3Ks6BW4vBVL5e5ZPw50OY/J0AaSyKxovJ5ynPzMl
Hv8fnolWmjGYD7VSn5FAp6BmRasrcixHb/WAQWPbTcJ50vtIdF41SZN62eGGUXKeSxpEfRi4RgjL
7ZnzG0OzzsNit93MMXCQNhYt3yWcckhcfgIKbEBq9Twy7q35FhRXsrSrKT+QbjpFPBxgZ5LgOMVK
WdZ35vHchC4vMViyQ922JjlT7PueVIqzEacOMKObyTdTdulr6o9sL4TLn173dTgiQZx+vQBrNJgX
o7SiA3APbRJ7EYpGhsdYtVl2Bf55cbAoAQooIw4PtwpMKkaYMihkCUzAcFEtBxh15MFSuU6bwqUF
dpofGcq4j+oBwDqqgYdUKNgsF7p5mUHsmMNsWOZMSSeifQ4Iwry5uLUM2f5LtUa5vkTpOwYRnX5s
i8BtNEBxu5gwhLSl6VedhQlt9HEVRoMs5ClujNPJAMilnoLcJrHDUw1wjM1kRulLU2aV0JqvowYs
jMH1hXGVy9HycHtI1LDXnuQH99/AuG5hY+GYtd8j5Os4F38Hi9VgRgKkuKklDGX75dKfFxtsKI4Z
r4NFk+7DXE4ey9gWMIXodAQW/EecE79HkUyZlUR6q7pJHJSUbXEWP3jOxxsM27LfYgpTiB58KQu+
YyPkHHFGCusMej0S9l1wAVeEglCE2vh31g48AO1Lkc44Q6IGmRPM+xEIkoZ0UnRgOj1HDi8t6EfM
BYlzADj2HeuPTBxucRC5Zs01m07QhwAspEuuSXGb8Hr0N10a82DZHBFS1Rn3aFLxfsde4h3w0FH0
gFyqfeVztCBnYoMHGZBwdRSSj9MGjGuIsZxIl+GzR9mJM0l2olT72qiP44xLWHFuxMDPBVmVRzR2
qQBaqJKhm6ygXz2145exK7qaZUgopYcbAK87mGoCXI9+3/aqKmEA/yLX004dygrOrU6kTkQsoeVG
YgIhms7sWMF38I6WO0kwmWq/C+5vP00PM94nSU/UdJLg/D+X80dAqxBqA8/QKydefDRtxRUQvGOD
OglIs8W22/PNor3FOmwJXYsFxsT4sgkfmS1qclVtOKtPnNmXEOKERULJzREQZ67UPvkLL2DTpX8O
ERBLNfIw6U/P0GUVExyRvmsVqJ8i0/YjSIJ5wq4wxjF9u+zVxM/al0JjiyDj/xFQXI+XA4wQZJZs
WwZPviDUb/tQM6Up6aKhIMWIom/og/gkSVH1PuoktLqE8KV5DDR2ieshUef69cJdzSjVzQCCcWVM
Wl02EJBad6msohGKgpZ6AkaIoUlG8vQme725/36+Zrg1QyQcsgpe/1YPfh0U0H9ZbF4ZJAJeMHOO
S96U3y6ofVD0H5iHmpha7nbF0WHLrt5CXJFyGJQx5yyKdglH08QFViOpPfcpuZesV4ZRx0rvfhn/
9N9dNlqy2GT2Bvtpz54KBYzYGNfEF/F5gL+if2YHuemcszeODtNPYq6NH61gJABTBMoRh1GSEJ1r
Q1peU1ofeZny6a8NGULMYGV1KbyakUSJV+YTPJCsCPGzA1SD7ucMm4RteEXxmZDYte7OxyXlmhbJ
+aFKOpeV9VzYfXoK1sljvgHtvUVgnR3gKOftLsX/x5yDjfatKxzmmGr8HdEpH4CxDl2VxvHp9kFk
zBfGKoaV08bzMFbpa10/L/xqJEEKZuBgmCR/3Mk1gbd/RT54Vpw+pJXZUizURZz8YviNenK3f1/H
diHyKWk7i+8Mmd7yUUDDoKrvbrnrxVfDxkAJi6scozogspCwlF6TwSaeZYyVyIu2HaUQ9XEJ7VXZ
QkhrvRF4q0pQvXjltk/jdSCDBZ3D7jVzHJO3iMXijIDe9Bunp7WxZygnaYKiBCE9MJP8tUHszpy/
T/mOBvV/bl11bvSO8cx/i7OVaoW/z3l42ohecaLhKW0ajLtydIWUjx8Xk+yayc1vu2nIqSwAM8wu
hbPrtzkpdLnQOUkedCzdxLgYpsfSTKZRlaYu7TRpacdKYR45SwWDn8x0wBD40ebv1qZEBtCzjlhU
XjNvHaPKBwQ6xkbat+pqFRRqda+yoLVD4KGEcVw/QUtqY3w2ozYR+q6+hfX5n0vuy+xASKRVdV8V
YmX8RsNv02a1tgs2UzdRS82sPL0rG1Kv6PiTJAM2EQsFGjJDCDFrmQJPqgP3yB6fSsN7rlYxMnuT
zD8AkndCDsCR+jp+oT5A95Y8z8VdZ1kEBvlz/svqM0mxgmxdkUHmpSQDTGyUl5TK7clI9L6jrR6v
vx7kpaSQdj6DNxMGOqWxc/DM8/CBZuxjSOTMMzTk9eK5aT1lSoWb5KBQYPB51DVsb/4zt5/SpUDz
G+7E05QZktNhwAMr3pvP3gKbGXCJfP33trhEchROH9KRVZrANAzb5XhVB/zjRNtZR5FgPQ5ujSdP
1ybKB4nWk9QcbPYI78wSsTZeviiuO3cjIN/d1ZLdJ5LC3yOdiHTADOr1HqOYHDdEPRVJ7cYdgWxV
d7SM6jeG9rYLtk4E4v3Kjrt68DiCj4R5btPhtqzKeansj9hHQevl/x8z3TYNnJfsJVJywIlsTvdy
RbiGfogoHSEaDf9HfFFIOJwH0n4SJptW+0p/JxtuU/PkTIpF3IedWA+DLRasIAYSZ2VhZDeXrRIY
4Sc72EnCNhDyx7+2W2nBsl0E36OAWRd5N2cvbN921HYGz72+zXuNf4mjZ1JiN4+0zNwi1HTXbf7H
+PljSQVWBJ/40JDpt34ew5SZ++5LltfZxbqTQ09GosPtCOa5E1fVeqXNy2stmMxwmBJ61Qi1SZH+
IVod6+ggT7esPMMTmvnNvNuBrLSjFPWQ77Rd49jgy3Oacfx8KALE6q0y24kitOvTbIkIZkbZZeho
LjWwu8eIO+sperpWc1QRAUEac3LAudwgaLQbCKwgDR9tVXtoTEWe54691NTTXWMJTfuAVs1EJmNr
qXd3IcemCVEWxLoy8tLXR6wHKiRo4TsRVHwvxHOPjlpEUs0WjkiBQirFYlzno6kTrNrkNn4SPs9g
kM6PNHeV14y/JqviuMF8cDc3/HI/bY+mgBoghgrmYFa3Z4NNhRJWBn7cbhuEidIGLSFs0ZoxusDv
CQhTWNWgSzb8KP9KlUYOyjafEgRRQJWhxc+JxxYVAuNuG5+amAc+oZdQLksNOzCe1hENIo2w6PRm
IMUrEysDHCDTFVOUR5WdIZvaX1ctFwE8GdR1Qkt5Zcol9dtDEUumNs5/ex8qVxagp2MMOtWPl2+R
h6e0uXc9tWCJcrKbo2y4CN+BC2GsXoPjD97FJ934KvT/bB3iJBQzWtG+KGZgYE3XngV88SlmRI6A
fZjFgTaT2Ux6EbNOAsK15fN9vDKEt4BQRQ0pUvoMzzJcSmR59ZaS4NJwR5xKfIUdsWGFH4CkQkSo
hfwUiAzLyRnMUltg0qolJiifHwcXmEYRTI1C4Bjoa2nNXckmfFzGufuQLKJ9gX57YMIyxGbUvVGX
XK80GL5Fjnf+T09jvDycrnURVud2Wb7SHpMZoWxCaHGynbZgk/1a6s5N3jTAf+snKue/gp+ZXnaN
i+dwePKPwZnhibkxQC91jzP8Czi0Tb8DYDyuh5T/jTD7hjOICYXjVdrNrx/o/zytbWqpaNXd4Xjc
JRQAHTRGw8c9JRl5LNW23NV1K3a0B89XfEaeGSvI28bvXZSSyUtFEBG1HCgH/SgQPHoGrdqj7vJh
UcMRqnOdNKahYED0U7/FISDICiBnZe3DnRBb65m9cYqB97uvOcgnATZQgAnmAkgsgWmfY7H2inGd
SrYmxOcVLb+CYnmoA+F27xWNohm96ThPdXguIWBZp/KpBpuMsLqEMyfUuhyfZCWsAFcfH44mxD6H
ng6YC2GBukWj/CDcTp2pttyRy8FeSUi8qCDa+ScYu87sQISgNWYgiNFG2h+8tbaPCxMqfbDZzES8
krWMEHK7CXfBqYUIcMgjBznxsiU77qVyq/eG0i0wI3UzYIBaJYG61WckwfycFBcjHiTEUmbpFpb2
UrMnpdEhITqqEwVCMhHnR17yZ4xOJJSv5750I8xI6OXPIqUVzL/VXIFyGrU41e8ZfqeCRpeqoafT
jcsre/9Vdhe5stNMgHXdNUJ6ph4KH58axKSeLzH6i663T+LoqTvac+bfu9xW2wPvy0uiy3C6eDHX
gQAzLBtioKFZu/ZAQ3zjJeY7QhdveZKRtPnZ91q13cdiaEJbsUHsfVGzZ/LICECZ3BK4CYwmgkwd
8YTOtJAedb2d3byDS62OOCYaeFkVNFMuLnuUlyJWnby89wNnchPh/jPZmXl8RXFRRXIZNDZ3dtCj
5tDj2+fkWLH8SXKvyNULvJjrtpK48YI9071HCQwPSKYuerhnuCGoxmLiZPmUZ5b4l1oOScmrn6/w
2ZhCVeYRZBxItOms8C54k3AmGdI4CcEPCf18dtGZWkaS9F4f9lTrSPi4lLxTS08OAQHYYLzYx7q4
yKzUzUBfScPwS/X5+DdkLz/E01tt7S/GCgGDwO194QZaXdW1V3LnUQcrXrfF9peISJR3vNYu97Pt
41LXucz9opFpUD5YE+WH7cszSkdB4rTvqWccJD/MEqxcDDu3VoYzZWv+XwNsChE+e6y+JX8TBKmk
rZlJpsKHXDtpwMpu/2vKPjFOGiFSO3nH6uB+JVQDycvXc1yUu0yYzvnmajWJEQ7gEfHJVrQbRcvF
Apwk4/fszClFPXJCr9mDUCWMH+tuBJmIZitJzvSX5YhdMTnpRQ6sqzoXY9ZBXObHgTn+tez9Cg0i
4afS3Tuv8cS/LM60xCN8+cx8Aibwfb4ax0FyTjxzOoXH9c1ELhgFO6CYl3lkI5kP/xtIV+wqUpI6
W3tAkFZ6zBoIyG2SwNyI+DmUHvOmAm+x7Fek0Bl5d68eyDTEQgN1jigufUgUNbx7jq/kXNkPN1Kq
q6rxUBxSIANOW/oYkJTNQaHD8MyRVuPcc/fwNVT8fe1YCpPPSmxnG5r9v277JfZYzui0C0rTZUix
xMU4pfFywSuGqT3Qib2MIYG5foemAGVNndWGEk/5oD8PQ+taO5RfVGnF3IOtS0yHX9f5ASK1NG8r
DJhnCQfSAuMXuzWZRWL5ZeFSaxB+c64s0ciI9+z0REQtw0BKqh/tBEEXde/s+gYGTTnEWSIMP2dr
1UF9+F3vEOPBrTEIWgWXTfiuDZ3FBnWyviBSdFm9UHRk2YeIlwz5troey7+c+saKsp9d4niGj+/Q
sVOdPQdQSO6AfdnHtq/psD+nKazrlwfpMm0cmZTdqhXGd3bcyjSn9hVwjHDWUf3AADAfG6DPAtY5
P36lzLsfCDel9YRfxg6wz3xTjeVWb/daHlO1WfAmRZ/QWsC6lG958fqLCJ1QA1PS55RrjR4FFiwN
L6LA2+iP9ZsQY3phcAhTp7J/D+3zFsYBKzGvbNZoQsStkp44xSaZnJ6qsEwCWzgzaH0SPVwmCWeH
J6gAts3ReDSu/10C/A+YoAFFD2IrKEJ/nGmxSuqaL6xLI08RTCc3X9DJNOHprKEldQ/8cKnwygcV
HJ8dfrsn/KKIwisRVI3XpnSvl0nXgoXcecksZSAUnOnfMU4Fr7mSJeFPUTWVCVYLmrpY2DCTguGm
89aNG3tx9Ssp7sFr6TLBhtYql9ZjP/L7VfmPBGs1mKjMRiQs7u8qTzNZyuWAvLCYjQM+btyexCku
1YsuFQinj3iBNGxPFS32zwFh2deJEhUUKRC0xi7mqjJoiho8WEq5r1lBdqsief9Ym4CX4sGZXs8s
++XPPPrK7rbUrFf1ZGLAS3fQES/gQPlO5TpkzjMTP3z4niv2xfXdsKh4A7+q7mMbz9KypdO2EbRz
BEgXmEGQIq6JxTlBuSkMeZ7dFCA7EqYN/UTcDOfr2NP2OrlD2rDmPXBZ8tax2Wv1TzXSDxSAP2Ml
2d8WGAEiGLUXV45GYp8cMC1FfCgfnFqMkJkjgs+ABOqdAanF8uWaEoWMjAg2SDSDPf1r3A8/l4Ag
anbpvwiRH3QnxMV8rujAgrTu3YzZICSC4fXbXL1Oit6mOgUza4+TRhgZ1hUpWUdDTVTyU7JlDW3N
8R9y+aei/TCsEMxSgEcRfrKEG/uu6CprfsyZXZO5wNPbxw6gRBhPiNcRSMuB/bPXJnX0dCxsEhep
ekVuI+WnakcK7Mxnkd96t4kPrdKmM+GrNaI4RFed9Ku1K32H3EdJ8SA9xnJsqvL+hchCyBWiUVg2
VZc/5dYLwnKd3+u+/iovGLz1Ubtmv520d6ApgSHvS9xjVivFi2VDfJ5bDGnObEBOrJgCAYPVUgWK
3oBlVhX91cBSwwlBPujCUs/Di0mX1B66Zh1QokjM23Ehv1S8y2mgDlamJG4U6nZWbXX7hEvIq3cL
ovadmR1jPPOtdlFpYP1xVkGCkuku99wxYz9KVS++mKhy8eM37jlmV2/zMl2DtDr3NqP5Pgy6eJwT
0UstoS5HAtJWA2hF37zl+0qJV4DuVEqzpsQ2RJ3PbMhMmy1QAgauMZOWoPpn8+tX7OSU57WaBsVy
N183QcbMIAeWm8r8C4FsunLbtb+y8Ujyq2rsYIiPNItUwdqmh2V1FBrAh2PlYcGBLiBqY6mngaVG
U2ZJa7RGrJybKHKURUot69Fxj1Qjwl75d6PBsQuwSy2GvOfPaMFuhdXEgnil2Qf5oGrwkYYr4Mqt
bgAOWpUryNC3pjZs8APh7ifGFb3ZcBu0pWc3Lh46/Rf4s1GfV9+eMTu9AP1Td+hCUNlbLdmTtnRz
VHx7SNhZMbzenUFuYVW3ZJQ9uwVUDjIt93J2lEPKWJyijQ9za8Q7kKhDLZRC8SiE54yHG4e6dKuY
LfEzizll0KxZgHQEz2pvc/Vs3VEj965m7IRpSSydIOgbLRxObZ3HBOhY3s95cdXfGskgGz5mPfDE
tdkRkP0cnQBhan1lWZa3TE1jLcmfGEr+Pmz0o4A9M7Pfn1i5/Ih8vBeN6mCFJvu7bUrWlRY8s0WM
epXkEiKcl/R4PlV/M8fispIC6QGb3KnUEC4y74qbixgsdtgEF2dcfycIMQgdqglj56GBKgOCY/U/
u0AkAbxfX8dXvAE69SwVoNzVClAAxM52FZrlvIcyyUM6a8O6JAvMbnZzKb8RIUCMwjMOSvSXqbKH
/yU2FBgH9Lj7baVgml1AuhiNA2KhMsGlOWfH9c/NSYpqLcjfJJt280xJIEv00Js6CrGlmG0I6bpB
/d8Hz9iDVVRJMHK/rjPKTBSk6duUU+3PUvPh6CaDgcc7uS2GGNQKnfH47ypRApCX/Npqjtt7gm8R
Cg9Sxc0lNtNIo46IidSjWCZfVNOHFERWigYyHIAAbWsq4aBAEUmgSjQhBZ7ynqAcYiah76rxIcfL
jLP+eVnf++ugkEX85eVaHqyw1I/QbC1njFQof6MFCSb00+AsopGT2ho8YMlGq47tQyqSVvO8jDmE
LEGKliXc9RTFpc2YXgNEgqjPzAJbK2E+gDWk4teoyveq47JEgTvJglP/Oa6P/OqlJyAQJefM6RIO
iOU8ns9d0GlnRAqosHWUIJH4Cg+41DttBkC+I60zNePqUoIQK0b+1cWdzea/sVZfOpnMJdwPSARx
XbPhW1gGodiwshNciz7JyEBRfL3v8g+zaJRSxAePce7FB1/DF1ADzhI4TtF7BbNMIQm59kgAeA+l
eW5IZGGF6b/InoHj3Uyd3PoLNd7xUENDKVpnAg/lJCke2/m/dcQ9CXHbR6XohgGEQrZSuCCc+pnj
YpaLGWObSHA8lIpgl9XmNRuE9yaPOmO6LbtDk+mgDH1ScZ3EhwgKZ79gBV/A9Ja57LMswj+4Rv8v
mqPlNjLHnbDfMqCMRLEhb1qOxnAWXsYzvMYfR4+3J/zWmirbac+vLWD4OsMFNdY84g35ugC6rDzO
Y6NQ9tCF7Me+d2BdQt/Bxbui+jW6cosA9jPEEz6j3Ej11cU1B7trZcwcVpOoAyzcnfZ0mp6mapYQ
AtsncqYFIrLBnbMGAbsLYPy1m5j3RYg/qwuiuNnee+PJOnhEF1Yyn2cWoDWnFEaa+5pylHzSe/Uy
6e1fvwmu3Wq19hnCZKFsyzyuo/QFwLO1wVGU3ktRj9eE2flcVb5GToC4mPpqlyiDs1hvYEU2SKe8
Rlgtgj6IP1ct1Kn1JYFr4BNZRoKnsPajCS4+aTTw/+RpSHsn5mm5ipNr/0MONgyKWpL+nrNj1Vjf
kEZH2s8tXhJvGrSKtekhl7f4v3UIrHwwaPAfmFFk6E5jZoE4CbGsI2IP0ZaWWBSUPtWBxf3au3EG
U5zFL2L3/vTHJRNanKge1p0X7ygFFKLU5aa8wirGaSTbcpUMWuSbD0lI18p5c5nmtguWOjmassvP
A2toKY1+cn9zoCtZ3yAr33lbE43ZX2wKqIPPxkKdBTOeJCqCBcAIWbgPHlT8tEEJ7OBANZZ9vJS+
Zi4TnsShW9zPxjwvqlfJUMSIQygPtro+HVu0cdlAtJqqlpDwHmxwQqetMbeE7QuQENFazItYjgH7
B9puTLrMLbMPcYubECv9rWKyN0cSXUyGlVaR6+6IPVbOt1gRgGWorLsflAt5UjGeyHLFIFESYWRq
uSQL/7poMYCEfo7MoAD7gCy7Nuz0nXQ1+s2MxyfbX4KwsHE9b7UmwUjF9qwrzOC11H5Lbcn3eDbu
dDsLNOIhNmcXtMAYS3HV0ubJzkywgX841aVv+rfM53WWxfsKQc9cDkKOwW0jHrUX8asM1vp/YXh7
dwHXqM+03JLsuyL5sfbLf37Gdyabgg+GD7z+JpqdfnTECsv4d6Aw1D1OfD+f3MehzD5d8CxzClLA
rZJKM9yucYYgWU3sTEU3uyLG/QuXphFgHAq5grA49qveItxT2TcJwvn0ivIC8WvY7LHJm9ni7NGB
XLWl/wTvW1bnoO96xwdne+xONtiXkq6mFbJ/b15lPfisLuWkighp5fHr6WcUL/Z9o6Do2QZ3zwtq
Yj6bJcHcJ+uc80AcrZQ7wFKqHXbzSqFtm7OGq/dWE5hF1pNwB479R7T4d0Q34m/OQSFUYzznkyAB
zooyRoZaBzzGs5mDPD5bJ/naOiL4cCh94XzC+5jOSVvAE8sRadEgzycwadYhJki2b6hAzKEPDGTY
4jjeA8PZ2WBgQhSBMU1WywAj4FKf5El40ibaPzislXjAfBatgrYsiqvNoAhM2Ev1014SYLusAh7j
vHr7rqdrUjKYG45xtjnomVPOVfhB8Pj67+ZXuNbB05WBipzGvIFe4I+425H2Mw0D+mCtcSQjIWuB
R9wo1pYbuKqtVKXKd4qXMeLGGS6Od6tkySf7m2jRo1vjF2htV9JjPmJETgDDneC2vc5JEAuOhghr
uFp8vDs0dR7My+qODR+LzErJ9RygYIn2zx83yCSTqnxfcHAchOGoepLrA7NEO4PbJ248ynX+KfAt
dopzOBUq2lMc4F6gt61zTiRukgYYjbNzuiOSg5MvuRMBPC+VMMBWueAgV4erXf4WVWT7+8PDzuZj
ylDtaUtbIbDYJAfBreDU/8iIEOPsCrYcEyGJ8QfGhT6L8SdZC/5spHj0HGye6zDw1rqrsOul/pq+
Iu3/oLb2IudgoMH9N0IAobf2NGoBjDT3xy/rnF/DJvwrSpmcOzCqIKdEQDrgiY5r5vr3hCloX70f
+zOs3SGe2hQtv++MDAagPnZQ6HBBYLDtG6IdGuSBl9iFZIkXl8JsReCJiOe0m2hyeHomF0B0VlyI
bHUiEmug7ykSrMZVpHzpqd0mVRcjj7w7gdAzPyM4MrnkW8R7DaV3egsT+Cd1+AMirGKge18tXqLR
ggNRfOGW0rdvknmF1RwaLnRIdkZCWEKvl2nDBSw7ywLSSyt/4AFucqSulOAvPTdjNbzGgOgLEAVj
Kn3gLwOJ7xq4jAX/zCOtmOAtrwXa1J/hBgs1Ru11IF5fattaSEiMy5PxLFcWZrO7NpMmBPqZlx31
kIQl7Z83so9PvQul6xJ7fME6HjT+Ed0hxhXyGb5RSw8iJOl7SVf+sl36V6iUVIbyZdeLeSmximSv
QyeDvLhkJoKaECQk0bUWqCtj2vmPdF2qQi2fyWvh0r9o87OJh3ud22ip4udhL5LUKwQ/SUJzmJdL
knKqlbxpqUiutYDKxpn77vDYyqsoPFW9gWHPvKdqliKtiM7jZb8cpkcZA7ANphf8X1aMTDYABv6M
m43KuZnCgjV/XhUlJgzW3nMUQVO4pxyqbN3uE9FmZ8I8j1fJwfabztoqzrR1k8qX3bBXMYNEtIdo
Ae7CFrmvmnx01da1NhLQBnjRKpFeqTgQH15ZQh8ncyTi+g7crM+Bq2a/hIeZLRgxqHZyVoiE7FU/
cFFOlM7BCiefDaeSG+H++3o5weXYELF0ZuZtngXYe1se+5TvbBhGO0lwWNfb6J7q0uCiru3SPPM3
kKlV69YY3ue1s49DNLnAu5EZ6CgT6jSEwDLt3f3oDUuny2+MD56xhnwsSjyYTUp04fPwqRErFNuK
GdaH3WcceRXkaOXtsAdD/U9FCDlzKUUYPsoymGrePe0TbMPB5yfpqpSx0L2BkCLWYKTCQcOFJlZL
Vp+rv545/zFrMjJgEVgvJsI8GLKuKgDLn20UqK2P+LHvwA8/rG5UV2fMFa5sUszQBu731jFggsod
V5NnZLS576Mgav4c30KnSbiXtmYAKu4YL7Cgw+2FcHpM5aIlUj7NBVoFixfKCX4YC/1SKB5EIXWp
2gBc8DJ7b9ZW5s2Qdkrsn8S1k1vhtl6IYyEZIEf1M86pby6wKVFVUc+BSRtMOedS7TmFoXMOXpEX
lhuslafrPtFLKXpMshYEbtV8V7cY+ZtbRD7haLtCWFJDlehCdmrFz9eaTtiHMGMoBRqC4a5rHdJj
AqcgI+bz0Mmkl8GD4ieWA0rNInsRVpVjaMrX0D0hwqHVSnKcYk3SSZOWLfDtKljJnhB9XZ7dx/hx
pfrN3rz9iZfBNJrtletKLECN8m+pzD5AilKf6EX2rUIblvuqWXHG8LPJXH+f7wsY8ika6/rZgnqF
4nQpP/D9V2CNXsn7GU1HHdwb7/PyceZRnfzsFJmpmaudvpJV3vWvR0Cfq/6VqjsHLnBQJdGIhYIi
SPsIWlnOAGjWHgxRmt1I26o1WrCIf042I+k5wTooqH10jBYyYUklZRgQPa+3yE0dOh3jMQRNwXwY
vUyfTBj5uS+rJ5sjmi5xNqSm5Kk5Vqw5q5mkM5gGU6cLLTeZosJ7YpUMgPcg47oV91Z/ZzKOLHNo
4doWiw+VCBPkU0kftM+kbsQOxrJ34LLkYmrE+xtBsoNMBjlgedj39GxwAw2v7ioT/FlccORc3I5c
3BiDQFbiFIIWpCDnlBhSOGAyv+VI6YBQloVmmE4EU49igdorndyVUUJmj0T9ffZzPpTNXNNxwBaE
eQwsdXlq83r/DdK/Ws5kU9aQdyW/NI+jMpRnBh4QZQojk2gWiAgXUzY5SHhDI2m8TZv5y8olZG/n
y+4MJaiRzSC7WdxZevIE3GgkY7gfowo8KKJ9BSpuMq1VhM4WE+caQ4sJ7kZ5U2BXxgWlo/rhCt93
hdlEYOGldCu491DwP1FcDpNVdA5ic7lXw2HklBSDBuc87A7YzJGt5DavtMRAwzWE51M3wCkf1pll
CFJBQBuqSvJuTvrEoYSZMttrNOv9F7v1LBLPw4Pve5FaV9pm2e+3yFXT070lI+l5kLaWCgNxTkE1
12TGqQ8Hw7qcCCfuQX1iUD9huE1mop7Osnj26ch+IzuoDtC5MN6CCsI4WgeG19QmJmceZLS53iNC
RlR+U1SpfTVC26yIxZB/eCfGIUG8/qEKNLLyKXIUM1S5yVIq3+4C4g7BNBzReQTxQ7gGKTs/zerg
yMhG+M1WgCbP+alWZQu5Nti1jkG8+mXWj9mmlveHkgHX2L17X2Gr0NlTew3hruPwtFz/Ue2Xpxww
oVKLvKzLik6XQaGLa8ph5WWeCPwvOZtCYydC0vOHAUBIJEDQzqb0AGknw+x5xAsv60QXM9SSvx4+
48MQA0TvdA9uJIh+03ym/L/jZioTq4jrTErIazmagwh2ytrU2YqRyCMkOKPJba82R/PfgCF/Dkgg
3UHHzvDquhyuK7p575Nle6FcQ3RW9U/gcc2LtJ6bBn0tZzhHBGFZjkDiT54sBxkOVdXBfKpHXbT+
OVWhbfX2ZZznjatN1viAHyLbX2DmIc00Yu8rqKPOtYQsKvYoC5vURjkw1SAb/unvZZaKQ7uK3/aw
AXqgtja7yFo0osxEgQh3lXwnZGHQITz1rNBpihqdUqF67kr0UwdnVu440xWXtb4s0ufWxzQgBzVd
dqjGo7KmUe+/p7fUV9TwIYq4QqkyAFCJ+4of5SCeukK6Swuixb7YYs0I1SbtTd8MHAZCZJ1TGZDo
nNYNaKnB7YAmxABNsuBVb6XY5iCvA6PKFrPz5Cj/I0tCugpHow/d7C2B5lVmatUt/RJnKoMEXl3j
hFLExSBzJql8VmvqkTID58vgi5CsQOBnu8oWnuUwI4bBHFCT0PfFxiXEvXINZyA6PKWVrPqbJhQF
QpVAGQJ7/DWuNwevpLJMLORc2GQfTFWXppIVTP+DEl5MYzjB/MlewiS2UBGXCkstKkW91S3F7ReN
R5EelRTSIqs/Eo6ihYu4isjrYFAYhCetODhSW1HHA7LCl5mDsYNpzIac2PZWS7s61DjA8GbJjST6
zP2weDuzxqv0y+Cd7Q9vvrSmdOzS4mkaKrIwse6gxnbVLSZvbk1/vXUFs9t36nySxhxaINfcP6mU
npkGRr+z6tSHQI/mwJpRYQO0eneIgqfACUruFFpOoP0/U2Lcoh15W01+MIDakNu3cLmEtn67KjU7
txL7fp5KCCdKLRNxZF/mh4B66UHNKXKngmHo+SA8xlREZfvI93+ANwh5FNPpMM1A1sfvQV+aVcNj
wyDd+81p5HOtQfaN6mGas3NUG+Xb1QV4Bbul5e6blR7cWhrT+HuRtbCopy0brqhN0cD5p8Vfw8Ya
trRnd/vRVLq8LqBeLnV4hVMYiSXp2dYmX8lyWSHY++y58pBx5pyAEgj92oUsR55tlRrBA/dXEWto
rzJbm8Su5+TyTJ8aBwZmI96+l8SrWtPuUuIMJ8MdC1oCE6+4556BVrEIRxlEpnrTWEDhR/zIv+Pi
3MQsEV8/HXhheea8mdQiiUgxjRxDrJQC+JgcRGVKpseqdp1xEFxxdZVSD0GqK8iXVUsPG0YH2fXu
XvPx57i9QA5n+XwUVG2wuj0zljjtL4ZFu37pxpAl1SjibzyOfIhLfP5MOYddEgfFZ3kWqZZdfi51
owlfebF9mXNYTp1JARso2TDIECroGYV5OrJl/eallSHJRAlGRb5LoU3+gh2EJkmrAwHPUbx0pj83
dmaLfMRtsQGw5e1spV124gdYgRMcopGfhp/wYZVYHi0YncohDkJry2PnKkOfqQcHjUQRhP5Ical+
qhy2znuj6F2F1/p8X/cEvvHasJSQyceIBXrWhbGX1cGfbOmJAHHNT5/hcr12wOpruIdKCdQdL7f1
Vha2qSNclXrE9XslwHywAic4COUKR6JTfonMSPUh3HYYo5SvZZDfrSo+15DA2AhXP+fZUz7NnO6G
VyKvtgnF5llcvCZlU/kH343l8G1OK6MbTpHLwrmYjOgR60b658UdrvDNWRy42a3yXvG8zAqWiGHg
5ZAbJI/LdXbcSYdKKZq9eK3AdC+ZBNJz3Ey53TXBbsLri8Q0U4Lk2wnVsWiqzGGI7eBfFiBcxeG1
Aacvy2Hpyz3KnnDNL6nacIJdK/DxdB/+2FsN2VhYMzFedqnuf+subomWT7BTRNdKQzQrS6+hiUJn
y6yCxLfdGtuEnSAhwGhHv0WpdrBzVQKPfChlt6fWltd0JvF3QlfaGzG62IRkPP+SXoOcAAo1Ok2U
fdEM6Y9Rvjz4qAeN/EISJZtFr+CkP2FcVQByjqKoodre9H3N49Ii0WriV052zxGKjyDsJG4sjH/w
uzdPTJ5DsC24SJ/uJbqzsDp5NqhF7EaKb7BoLg4ybz/F7DgBS/2uJIOkCMqm2+ajj65vto2G9iZK
ccruyjuwu+4QPKSYO7QyvYvek0DIvSsY4zL3GdWMorNQafCTSH3P+9wwsLzqoEaO5fijqTgNKsvi
ARf0yJ1lSx0nJnvBTQUahdNdnPjsp07vZYf+xgHthUBkdH8LzBwyp/ziKbLsphZL5yAcAhM0IAhM
9TLRA43CP8cZ9mlt9ZH3i7JiJY5yXjY8d72l0OAKV9Z6sJhVa1TSRfuUXSzWbqow6JSILw44O/d+
NJcMIdYhJui9S1f2+G/7+PunU7Jv/PqlA5LVtDS3+GweZwtq/odn7QdCQUw8RDe2dpY7FE5N0ZQt
QuHGb+KpN5DhFxx0PKGrvwfBtfJ/BwLRdBs8xNC5VxPNZOfwMBhIcgIHsjQBY2ZBc6BTTIuZ44iK
myULf4jNHrpHT0czvFvc5Bu3Vxy+nvcMOd51CZLRpULf2EZMdBZkbmG/GDzb7Ga1G+s9FuxzCsvw
HDdRmx2dfq7mY3ODp7oMGNrorZpWcuN/VcfNl0KTV7enTx5yAo2NEfJkEH5A/y5hFoC7aD60NyUa
w1G//e7C8LvZmZlPmj1CgokS+HvLemB0/ndzBd8KUTl3UEo4wR15ArxTiVUAzujRQAEuc/0bWhKr
c+lZdTVu97AZvNdDxF+ZfMvu/1CXmlznp1Zxi991xsH+cvqOBslroVHX0mbugLl5SM63EZUD+zhY
FUG+IMdElQrTVc7bNXonWbHcw4OCAjRoyD+vSqnKlgcDYFV02iOcjAyyOrBQyI4vFxox/3P3XxTe
wQDs6H0uM0ujs/x4J93QpktStafTWe5KRbEsRfkvX9qkAH9JjNuNqjJTTIPO8oUNyYWbNaWIeMy7
PdmUNfIBTUahqigU7IN70nWOhbihvLjghCi3jIBJrev5sAbn4l8Pccr6x+4flKm7rkdbc8gswNJP
SNt50x78+qs1XnP3WmYnYe9Q9wzxQswCbA3pABEUjdNBhwz/BY+dNwVFnaK/ScZKCbukr9lIPZS5
jBKAlIw5kXnLAAEi8aAdiFedMHEWotW8IQURED6B/VbkDime5O76ce0qtMDiJM8UUgvf/K2OAbQx
4Vw+jaCsMOS2CamPVROT+SbWs3AHzVeobfau2GnojeULd5NBuRPdLbPOs94CxC/GsuJCaSCzupXe
n5AkqxNAcdk+ecupGR7TITBKdiLJBpt9oU9hN6cb6xcvwQONgqUrZALwX5X+vZXSS8+3Pxw4lufP
CGLtrFQTfO47Iv9JHAQK/Ac4hx1yw0PmrZpoJw9nSIqJ2SXa+Sip8ROVwqI5PQLxmvpIWH5k0/SL
86qJIPox6S3yD/gT8+YXjQFoJqUISfn+RyhIABNNWJEEtN0Ygtv2bv+eYAoGcoJsTOE6S2XyXu4c
iOHi1V/UYHvRan2+4GYm0+PT2I181stknKfKqg09p9/l4CVbFcd4x7yReHm9Ex06KKalk23lZvfF
VMESWIDuLPkMNZ9Jrs79O8qF5EvZid1OEz/Xa2lnHPviUWZrPoY5ut+VuQwLBi2X218+v29vLr6+
snwD6afJpDr2UWpN7Me4UtnNeKPmGoTrPHR/YD6OompFKYLYFXJO8VyXs0CslQEud7v8i3RZ2WI9
WfL+qdtByL5Oz91FXDQ4zfiFooUR9UAslFi3j612N2QApUTtzeI1fghRIrjpn5Kn0ypJr1htrYcd
KrjPdY1rPdjzIPddOfhnBrcog6xZrwsfzwkqV7Wgg2+tEn0HB0Q8nHqXdBPKQOYFAsgwNbDY/cnr
Tisb28A8UFKCxQ+zAl1vt6EqMsr6M1HPLMbFI3bj86A2WufVyVMf4WuI1uUbM/JmS0g1zNen2S5b
QKeTuPBeaWsdyR5rew8ittRWrl35q4gECbr+eE0SfjhRdoAnwxEgsvi263wOEjETwwMSdCIlIwgG
2KhE5/1A3f9bjY2CbL00xHjHt4L66vuyLUHeQrNy0gcjkstpRnn486/Dz4ctqp1TsQZlSAKncigI
aLetCJ9aS5w9Ggd9ZLLeeS78GDopu93eLeodA7qeLf+Szyyri+bjFYms2ty4ZljbUN3Tv6Fj9bef
xGJqmvZJ4+L9ThHpeT4UQ1rwnOwUYb91koM4350H7pR8dFfCWgjugPS5+frGx6HP+NP+Z6SuER6u
qWJgfkvkSMqKBkGr85nUkqJF+qceQnUhccOpK5duZdw0EuRxtIAPpj5q95c+hvZpwYnYwGQhknH3
CpjGjJa041WDyOPPX2B32WgILStVvEgN3B+9zexLJAge7yDyZPxywoGecv6nd6ZEhMDWuAqDg7Ie
i9dShyrzlhwh9Z1Casm5mI5LTOr+ItW2wwmucKU00kk47z60DOgqIo8CkjlXUWiUFfHe3drm/LpI
mYowawfNpzCqUhLzykXt5zNkZNKEeuHWlHHZfAlsm60hVmXr6Poc0PB05aIklaEikzxSyNScBQul
DjxasqJhQAxfsa8pV7YdccVc+uVMF6tv/7iu+SsUdAT1PlI3FSWtRgefNKAVLT3kVeAoL9CwJzXq
pZbIYSsQpYFmhJIkFmRLyY7mQJVownLPlqy8j2f1B/hHuvKNmOTNegrR/hEIzj0bzgS1VSmfZLmy
pX83UiwAHiAwk2av02NhBC87Na2nF8Hmf8hhL8fca2lWAOXXRSqGyoh+jnrMiat3szSEhmvGuYch
7Do2fhkBbdvDRB+q47lTUHVhAbPosWEjRbm6TDP5g1sACbxYWXDPyqRSN3/m+vXOyMlwlSyGL6jz
2lFu1Fyhidv6kQvTw8qT3y8IqpDN7SaVXm5Bi39Nuc4bC1C3tzu03GMftRCe3A2PhuSUdFh22t89
8y2NxTffa4+FtXgUXPs+I3RcU1XMLGrh9LFb+PDTO7GTmRGgfhTqnGgBJfDg8znd66Bq6D4vFxkr
Zu4UGnZi/KNd2TB/swKo7iC7GXexcGBATplXuAtMh93/MHKdXQt07f1ysKgO8eJRblGdWS9/xZnR
GXU2U2UUEA3v3TG/j52wGHhFGHnI2akrFj+uavIBfzYijIAlU1hdYF/ZtnHuh/DFW7bxKPDzSK3C
mP3lJqRAFXN49RG4OSAgwIW0xhRy0x3sWfPOz0xqXF1KPzrJWFyTMghbwQWCmP2HFuclaaQeVzrp
9UA81XOsuRnrWCEZik3xkeWHt2rI5OrBk6XyXSDNqpdQvh1Z92yONQh9F7oTd7K2cHZlNtj4IwD5
w0oxgi8dcks5t5AN4EvuOIjfumN5Vo2LqcBfZstsTVVA2H1Bmxaz03oHfyiKLGZsUyl+N92GTotT
3xPvNVvWuynFKeBuk/x0yt8BV6G5jah6zressOkwnVKVq2pwdvGgi559pYt6kab0Pt6NucSZoV99
k+I6iXsPEjGobXrp1CaiPiaxKHrEowM9ONk4w4p4e59x84bHFTHmVaPsT7dVjE954cgJCt7Rv1rH
WdXyVnyvkRwUEMNQUGamDujoIUVtXk5dR7I35JeJAqDZz4Min5CpKYsZC88cdtKwKafa9T+5XEXF
emApKv6QRpajthrvKuxY3FBW+uxSZjpFaEgE9295QRBKXVN2/yWmvIyAM6qaEphDUqqrOnwetQaM
SrB9UF3cL1vm49P1FnQCgrDypINRjz0JET52G42Vyc3FPhEC5PGCFogSjqP6/4liIe8b4YzsYM31
EFkur+Cd0k+uA9qhUc5P3zTbPngz4djFQu1NqTQ5clVRXi4h5L7/8ivcHMtiOqBFKux6SQ3gcae9
bauP2Ll/3PbMVOg4O2hLxRUBezmXB6nMfXM/FzsjOFzFm/bhwy9cbps1tUHZOxoL7Bi5hUtvu3Xo
FzvrdKuAwz1yy1O0RqU/bxwJbMtCDppFYj7GLSdLx6RWYTWjifG4N2sRujB7z5ywF3tbqxewgfkR
V/KwxoSq+nb13i5GPIPrJEntcrJq7USprRldHu78mT1gNZzZq2FAp95tauMQpZx5K5V6yORwLMc7
4fk+aHX/8Ga2GxxuWRh35Iq+EN2YqdJVuw/ywLXVUqhunw9xLH1169p7A5QQt5F1c/MQZBL/XUMF
Vru+U61+C9UeRFUqzaAqMJqTi9LHcFuN1j9ljI6R5RHzBI7DE/T1qBosHUKRqoz15s7cwM4XnvXP
oN6OskNEH1AZMlD8u8ubVPyvoTByvUub78CFdB+Wx1gU0OON2d2N1jgzlCHTtIysC/aSXQGrASQ7
kiqWgjOhH2MaLOI0Q59itHZiSAZifHs25XKJRRjn+YVhCc45Eo0BShb1RsMeZeyQ1Q+dSqz4xrOK
I8IUYsviPfHOG63hjqUC07iaVdc9k1QMqHJl8zTdiHAhFlJqCCGtEdj9qz1V8M89z4zVgNTXjoXV
JS4CqLEGoWDGsQzw0dXwA4yWge5bFDpQo7frUcGditiBcVdAkeyO1dBQ7rXP2vW0iI5CK1C9PCP2
JV7Zuh3g9dutLiNDPMFY3WwNavYfYoWMc3Psb/zgtV0w48sLf1qvTorMTjwXmaIeu1BNX0wedWwu
UsJcW11UUvD79e7xNWKKd9mtaadCCv40Rp5/5DaOlp6cZZ2iKEGaWd7Kyat2P8oqNKs7wIQztGSp
n3rz5GopBKouy1THRJejmn0lbZ03fpEKRl1IEGSuOypIBtOHqmG9pfFwPm/Mkx7ebuB2YzrBRiVa
f6v8FNIpT9bElwe38ON8SsOuoRNSHBulpDCU5KwSQcASUa4uXIi3CY2Uh9qP5eqAEKGzvcJLcLO2
ng+aDNDGypmgskvgFnlkq6o0noX9d+4pUBQAzMp4PzQk/9UbSHSjEYJwCdxdjm01CsTx0m1aQ61V
bgCcjIbktIQkkAXunXXKFQBiFyVHqUv+vC/SrrXVdEvMeUNTaviwMSLYAOdeAAX+xS2n5q/lxEgQ
DptazUObl35BUMjMF4FnXPRiNDF50nTvQfufPG2VDbjdntSER4OkQgyujg37mwmxvpRWPRUHxq6+
mgAQ8DI8iwQaIiAlMHqV/GffarklLQtOuP1zYy8F1rnoYumW5uHZ5/pnjOwQuRmxzn+/CHgWXzo4
q4OKZWlWnKYkkxdyc2Og3gFxJjN/go6EA8lkVQRiyNgP0UA4jrmwyDU200lKS+D/qQnMzIqCMoEH
1S/VahpBTSAZDrvBcuBh3IpfsQysFhH9zX9cZUfXxu98ZkiwYDcBRmSyNUODRXI7UZAFg15wYZeN
sgGJTTwlPN8u5g5tnyEyZ+DMLaXenbS90h52xEEe2JfGhfLoaKPgQJtZx8/5KWM2abCTlelVzaA+
AV+5LsVFFQM51lbtFD4HObwet737xbskGrVKPOp6HjAxaM/kJzfQQjoCdNNV1aclNz70gbIyCnVR
N+emr2MVaNVGuWXbFV3vaK3YVFGK2sLXnCa2ygUiO50gT8tKE/suyciP2upklj2dkFpf2hFN6ZqX
UhYW/pdHqPHZICVlVKiMl9GUZr9BxXzfFLllir9G5VEYprbFPXroouAL5dZBUVvV1NGtFbyUlUzC
u6SColh/jjTwy0aKyGuj13rrdITfZg97TZqxGzZgB5YacLqnXSo6N3Rks0+3chQlpJDO+qD6tn5I
MSalzQRvV02D+SuB3K6rkGy60WvRsPc0eC7JF+517ZzgzYSipAdYNXXQnxCHmk+VwBvpsxIvxygB
yav4U5AMcq//aBfvtDTcXH3AH0KcOIAeXIa9Wa+177TP/27vDlk8lLyt6Y3iA9TpO59CVlG0YpBH
FZVtsnUhvsp1O1EPVMWvSl5NLp7vaPTDvMkhosDWDwh79sl7jz67KZi44BAYqNf9q8IlC7kOJWRP
Lh3L+7CBzfqNdAlzCg0UdsWTaxsv/a6bvsfkRhVTGDdVBInzLgMJPRPHpI0sop2ltRD/2pWqZTCo
F70S8Za6OpT1iipwa6G6UGGURQhleRLrfSLeJakUZ7y1BWr4oFjmjye0dWtQWKDc/7jp8+G5oZc+
JzTdKvPcVmmpNhlxe/3+ksH3JiBUkd3rySiSt2McbK+S5ZA7VZj2/gXpO91GXXx/eqQmkGB5i4e7
hI7joJ3ti4Q6Pszii8i73VhlMqiPRpyDQHprwAaKtayOTN2eiGnzKpROO5oySAyjmzLJha1Y2IQl
2O+X+OuGH9BUbSZ8xOlKGBGBU2IeCTBMLYuUkGj/J6gZr24331toS8jEU2mja2NEUO90f8HONO1J
ai/ScTqrpxQAVlgPPJp8QUMoNaGazGez/sKXf3j7/rryss+fXLARvQQf0CmjNElMT4iV8TtB3dMX
AM1IG6bZLmeGf8CReEsuPZwWJck0nSLw1ATmmYG3xEerXRzQGlt+PCp8zNBRqUZKOQiU2Tt1NIkb
gCIxAvj/RLVVZdpkXbFndpRtLL16/7NZ3x0l0SWHd0z+g2Q332tAbVfN8leQUWslNVlys0Yz0WiO
1m9lhum5Rn/ah7rpq8zXTlbMeUhirzO4CGwRClkoe9CYU/eUy6VaSwvqqLM3NfuwPyBuZljae/3e
u4XD+qdnsMKQ5VWHst6t6LrEE5yUG6jUiB47fTKlbhz61NNIrzn73ARxSRdaN5R45cNVGzABsSq6
HgcNsS1JExSsp7BR3PBpBwSTCOVLmQmr1Rfq2IIrASHsyKXojEY8XVNxUFPJN5M0rg55W2YoITiT
AW01Iw29BXiknIqOH81n5vPQXFJ5aMrrma8SFODNKTxS8KJ5n3dWA+i/yHSMxgW++KqymK6Mdauo
XbbyQNBir2c6ud2WGRPS9HA8AJq5zASCERLwPbmUV/ooSD9yn8/4SsHpvBVwwTiZq+3rmLSIzkX6
UK/Zf4GDaJYvuXyW6uuoMWy/oH+Ces+bOEyFQiso6ewBiAystkHy4b7njIK99DzizzL5n8kIwr8V
HTxI56q+QaQxhbE2B5H8qqYCyyywFZXYQUpQRBqhY1p08HfylxyZ1WxufrQZnZtKHw+4pARdrNrY
pi22BuNf+Or/brO0n+cR6lypHANx3KktuUWwj6t6ZqNwZN5ewAtSHA3/C6U6iVCzd93LZSC5WUZ0
kaffv7e6ebyQOhe80o3+T7UkZVEAWuBGAmMWDz9LMNZ2qNwqBUpRxCDrkpobogvRg7KJy+tK9G37
i9iGi0QfNFw6NhlZs5OXOZ3gDEHgafCkv5x2l8F0jaoaA0oUBFksDH2G5HbDLtKfQlaLrhtvpaLB
PCU8fz3ZPNYzoG1bQFsUC2k2gkG6FiJQZqKRJEogc6oOaWQbGcRo0xeMF8FQ0aGCGa+vfWLkq1nN
kfyHmyN5wkcvxlUq+E4CwTedEXqGWodEnNePcm+T0xxj0POcoQOl6ttg8fq5dUBQaBYwptUx5eHa
wzW+nvEEwmcKNFMJyfm80W8LqVS4zf5/61TDE4Q8vSdxi728l/sCJBM6v5PQzJJaehhhOml0LyzI
oXvunSWZfwygV1dM/9lgoX+hqq7lIphtFu0SyBZMGh2htcfKKzmkX9Wc7+ifYz2IHLjAEOdrVrYc
qL5RpuvIFHwS3zLDk16zpP4jCh7kvrHKljyAL2642l9I9LYcS02akq+OwyD1ITrmT1KROkdW/qTH
DSlEzMAZTVL2z3+6RBDY0KwLt2aHvrXENL9H3oHKvZjT64+2RgJBheuCMTQbJ8nilHkLa7pcYQ69
kY70N35lYc0uX/3CThN49BdROSo9QJAHhVDvyPLPozPA5unWdHSIkipcy4eoaKZBQvaI2MgtM6Aj
3bTVYWW7i2nZqoTmiIQpavg7mcuXK5BSKgxUOuE5SaFadb4BjW8pki7K6iLToaCqgnvb2anTKLnV
oXzkCJLGGeFEorQUe0EsBVhPcrdFkJNVOuEvd7OAwXJUSi1VVMXtNHAnBznFyvQfeddq5tURi7lQ
br8QOygRr0N6tetIWAH8LrKqEQslUhFxj+sia/9PNSOilWEVIYdAy157MbfGeo8qwVyo9yrL3m28
y8HjgI3FTvpq7Wi61nufvmj/+tuJwBSLGGBGNJZA1DJMoO5GD7W7WX4QwSm/X6iiMB/lRU4+UFVX
+4E50a8/45OpLa8OpjWDclj0n1C9A8AxQCLkQMOidEOByAvMJ9V7YY4wd2EBTpmFbPCbJ/jS9+Kg
dhGMthLO8ZeSq/j8kEILkk0QaxzFee6l0yYBiFzimE6anCyL0oiqosYbE/u7FLJL33GSVdhnH1Hg
31+KE2u12KT6sYhD9LinZ38McvTalFxLZyBADTpVMn8L/gPWkz0aO2OICY3cmlmBvINhRQ66SX+d
1f/N7ckJXaSh05WQKI/sZnDJNW8R6+074zU4bfGbGy2BNT27HpU06/urQ2dB4rqJEthpsk82s36E
sJiU/wxdUK7D0HdcZWFvfg0x9bnAf5TyJQ98sy/LZktcgSatFMjaNfVnMuC349xdwBS8l1+5eWIK
oJ/RZboW/Sg5AZzf9znF4TD5DGvEuU+tDhu8b7XyHF+9LDtiE2bGGt8cuYhPFHr7zlJsAKYpCjGx
qfUOfZ6FqQh1owe4QkpZ0V1TBEFdSJI4YGeF7UJbw+eOUUa/fWDGEKBfGZhX/1p65RD7QjA3i35Z
5rj5IPJvPZXbHiSxBOVmoMPdaGW1K9W/qWFQ7hkWxzimlcglNtsYSr6uPw19LqX4nbtsaTquoGy3
Rkul3k9Y1T729zlESfX5ITntAKGZ9YQ1LJsbregAJehvdZnk4GJiGlaSQsS53B2SjNnqeTBFqgVd
hLdKh8roiRgNzudO/OjtjFyroDufNRno9J21ZXKJFYjg9fPZg4rKSsWq0vuyl96UPLsQ0uMHjrlg
lh9errPStz8ucu0z/0p6sgBXtYe2ot6N49h+vkiTKlsXP+jm0eD8rF0x48//d7vkewGXnqr+6c9y
4jZjV0C/xumVSWV+NLq5Li26bqLOvXWoP0FXvCzEMamTcfll/DajQE4OyoznWSV9Y8CGJTIaEs7D
80exbedJgPdZS/bbx4Noqk44AnylRk5YxuWNj0NgG7KSNhRUoQm+Bznw+bR7Afd9gcMf3e7V9Kca
D2ZFjS3/7znU51OOvqs0mdjCxenXoSxqAu6726Ze3kUGGu7DuC3EXky78NCNA1mYCz7Bk2K7S2zV
cd4vC+hNSkTg8W5pWwLuq6vePV8H6AE3atS4zsJf8qn1G0y9s5OLyxmT48uk0wGnj+Rdh1gfsrD2
5gSWlrD1B4dV0xvzkOviKMd+PNo6tto0dTkGgApUV+7uSn+6wpKpfqNCHCBaUkx2RQU8/GPHndQA
Wvhwt+kJSH4elOJ3RjycIBQRsnyrnjVn2+uS4xr/kE87BdJ2PSE8LN+q9QNb0ZDc+NVe1f+SWoGv
hGnYBYjCospDtATCAWoI798wI19CkxIqPGVIVsK4m8HV7Cg8yyi4EpAL7CZZSAIrCMhTYBR8mz6N
FXafQ3/eEtd8lzLVXROagQnY9HtHVzQQkuW7OwihKkaoFvTehC9uEkvL47VKQuEIeViiOiY9m7Mg
A3m2bkeVJIedZKQoXyWagju4OAMyNzW3MyC4yZ42rUuUP6bhgK+LNvPWcf76NRqlzoZo1TLYa5XP
o8vRVT9QlSnx+f9xKAclv00nUTsiofLEJm5fm0ReSZJS/AahE1Oc/ZtE2WYjEbm0KeuPcZZYSKiM
AuKORLdU0iOkxnXCjRSpQAVbTiJY0c/wEncLuNBC/WjCfTjmBxd2rnwyZVthKGKcGs1IM9KMpTyn
BtXBy61gx9I7FiBiDOk9oeQVp0r8Xnan01bI20nh2UvlspxXKpjMTQQ3hijaX3q2iNTg+018DGHc
7bEM0rIjRynbPwLwxJ3/EXaf7TKPqdXBhjIZuaDhD7VXEgkVcdrzz0w31UeFZKmNVf+I7XgpAzhh
q3qkAmRHaCFOZQD1YcJaI1h4wVUfIlMZXS7Z9Aa7Tsj8s2wv02Kxh+O5q7UeRPcPgB+1ZvqCtIjg
bvx0U5T3DCXfH+CvSIFQ86Ql+ug0HU3gJhOKLcfBKFC4/f6kyT8D2WIl4UU+cn3Jj60VyT50gi5r
64eDgbjvXqsttRVkJVnegGXWUcpQB1AMSQ/Kh7R7IIgepc4xzBuy9tbeHTz0kdqNDJI6N5DJ0zJQ
0q5VqwLFei5QHP3B4JxYQNR9TkknG8ftET1kXMI/9isyAt1AfgNLVUrgVbjJ/mHGnXH55UH6fqxO
+hduZ+kFBTiv3tpzoYT066cYnhZxpdr7c26Qk6ZuaGObOSZwOmFx8GDT4vlu43uTHPdyC/i+XOer
4B7FgfWvQCH4De4u3ybKcRoTY8Eb4Ks3WE8mDuxbX2D5vxfbHUhYeyfhJN6HYblbmsIsMUAGKT5u
fYAvU8IJY5zwyWReLOTckn587KrhV6IXAm7orv8DbN7kJFKfIwYX+ll7WhIdnu+O+J+dxPslQXtf
6oozEAuxzCm6iFQmTOzeEcSLiwzIm1LEN5LLXHhZNsAuOGx9z4jZaFZxv1rWkJCak7myE1GcZntc
+7IKy6d9bEmSpOjh4pOGUu6z+xJNpoGMP0RWRd9K2VJWbLmHrfZLOrmFvGUYLXCPvy+Fv/UDge6/
CtL/kyeqFOzkTvZL3mKmbuFoDvQgAaC072Q/2aSmC4Aiz0r4NKzutXYfe0CGaSFK9jJ99026bQWi
N+tHgEdkCJAJ/q+Ou94jcW/bSlyQy15xWtMbL1xsM+UbXMHCpeFZE77mzr5bI9Tq/i8fODGXghu1
OrSt2jf4tasVFs8qzlbgsAZiu0SB0c1cjL18Z8II7S1IJJQwwNoDg1eRTlbg4W+3TvvW667Xw3HU
dyl0wZ7Ym2TFv19fneuNZG77kE+ggIUSCJl3+whK6zwYXgRHqM561cqqvmRGgstPKGYKj1DW6KuV
WzvoHnOqDo6wN6+ywY7EVGaOI57MRZpmkT2nA8Mr6tbVpN/p4Tjk7VKQX74J2fQxGy2Ip3C0ZPBR
gj6e0WLP9qC9nw/bjje3Y+b/62BvnJDDT4gf8Imm0PdaHU+OmKQiLZANg4JE5/uLVivHxRoE7k05
WLqzNbi8rs7NZZLmvM4exAaDVMVFQp2x7NoBCzxE9QCHmTsOViuefCA6Zr+sXzPr9ylPok8oNvIl
PEv7Gc6F+O6psU9KxI56R0HLCpMCYlbef7l218gmfPl3EkaiXhxq+EbKFkIqg+9aCt6OJYlme/NX
D3N1XE/OpWi8KiDQni/2bB38UB0NIzrkdRF0APj/TrJL/12tNUzHPqaiW5BDhsmV2fNIxoouB9Pw
7h//dN5leaVTaaaKnbnZ+ddorw0TSeb2mle9bKRa9ef6AgGNtKY3pJtDjtJ4iMBxy+TU1so/shes
gse2Pg3/Jen/cRFRDfBut0kxvqqN5MBjmfeXvTUx6FxpQN8xq/B73B9+uBUVwIRXUNuP9mzT5rHA
EahrevYEuwvCEtXxPyjyV4ehahetLF/yGrqaVO54XyUTL0MyCuf4mtIeRbT7rljgYTbrSHFRieGQ
GJzKltyAyxtWKxiATs4zOlFPF2b2tajuL8hMn5laIlrbDNZJUIAHquMMUN+q2mGSoHFneliq35Qe
SqTfpIWFNfNAa3CVGQU2JZhblSinRL3eSJ+wg+11s5QhYRpNzoi3HrJN8H1SEKbHEdwQZ2oMMuZ7
msy+Cut0VnCcBZ3t1fOvRkCmCkpm+riu7mceQXSOM18Rn+NhauvK7/nKymw5U7bBYPvQ/ki5IT4e
a+tFKX+M1g93kiRrRO3mtSWU1WL/b7BqnSFY9sSh/8OCe+ZjBCHxmZ8g/IAJIPuC3RkWuKDKrrPz
AxNCjiNwv8vz21GP35GgUYmhZo9Q4UK6NPhK7j850ZyxNtYXGTcmiUywrqPwH9wSChMtqO3kdRPy
cKiPT9BkwMXX1nb2LjpjvPSGvw+Eouiw+U6UTom2d3lnvIaIN7KfAcOy9p1hNiwrYq29cxv9TNeZ
Q27PCSeAU/RPhZFiPFPiYzeGSyb7E4GLYzFeZFqEFFkp3I9ZHdqlx0BxSt4zB8IPGL/qS4rV61XP
wS1tk0pZi94SFnbO19GqPYeQH8aoayMCzt32MXgkioAnBZTC099DMFH23b97T69n1QNRXNiG1k6I
sviP4Z9Jhy9S+4B5o1fhJKZcsH58HLPJsW5C16aD2/uN6Ufwn94XXcEBPo10/yaATWUnxUdWxZZC
CzsMiFlDjyveEU/iV88tHxVk969jd3w0OSIGt0NZR1gKorsHiIQCdLFqwHh7VSdk0jfq0JWczESs
Y7GYNcFz+MNDNdJBv3Lounaj68iy5zHe3nUwTzYsuaAzVpO4+i/wMh7YP8OIkG7yXLPjdh6pI65I
Jj3AR3600TKrwwM0isn24rNHR3WhyQY5stYwE6cm/HQLAXDrO1SwRjMJgkC1cQ6onilsBEeTEeZu
c0ABUZ3DrSP/3vbH7HZJyETAXnEa9mnBIo5cSuOsMHE2NH3xUtBAkLW3gL+9oJ8HzbM6yCGEFdNU
yZyYA+4Xv9SYbzgb2Hm0YXBDwexoPajW0FNkXVD3no1c5QwHYvfrh6gfOakoxNoKz4c7y/JeehDm
f6NLNVBIJoxAiVI5aRtrEWSinXL6yXyYxxkok5mRUCPFi3uh8pJERrs5GD61Sw5JRYkDnmS/iyfm
1qLyFOitzgmdlhwuW3m0BKaTWKxee8irDuFtHd44giHKnzSAJGONTW566CZwP4QABWBpRGYVr3w9
p3ywSiHpzS8Xp3jrkBnLfb8c/Ld8YhlyH75x5fGeonueSL4VMUPqBKTFl7VuuTI/jhpvLoDO2Yb4
6DRAnx4EFHRsWFKNBkxgQNm3VEzwhKISA1+/6rDDLgXXqZQIWuTEhv4Q3eYAjZmMwTERClYffzqa
13yDg47jzN6WJeFujE9CAoCJ258WoVwsxfdz5fldCvcy2eUTd/O648nelL7QTho2aNRA4Y6ae+/T
air2HXUGiQ26BqZssRPIuOM+yyCUTAnJromTvnralu2GLZHiRLzoAHVYfFwB/7iCS49hRQK1aDx5
xAr2ZHGFfxGP6EqPw5ZFk/rqi9U4uhscbSSlvr6Q9KbFE7+BtUfd71lHpxKWyzlwcxkGBHug5fcI
0/GRyfiM/XN5AOO101wSFEu65XBInpktNMWQrnt9VOyiCsoizWCFfNiY5yMrcGeleAtRKafsOJN9
cGMNRVBC4KTjs1FDilVwJz+CZKF9cAc7Covo0xmEMGEhVruCgp9lgv8Ff2G5KdPgB7tIwnsYOvtK
oXgEatvJkDVApZaYqpS5+WumwvUOF6bV8fwEW56Xcz1W0O//JeU/owO2a6Fykim4lK9So5wFgu/G
HyE4p/uxz8wyUYz+PHZNM72LPuM3VSwpF6hXWDxCTnYW0vpRj7NZ7oWjL3CD7ycbXWXSKCaK5dlf
5tMREsdjikef29G9JGnlSTeXUb+lJ6x2+2nlTWcZP6ypBLrIEs2cJ1o0B1AZ2h5oqf/HxXKi1sX/
1hJm6C3X0Iqpf7urtaUFGUL0qMBYmIdhdEZtoqycqk+8qDWFx+IrbeDHd9k+jQZHdkENenGBNgvL
cS98fdoVM8lWqAzhcNfavWpl8DSLOjuANU50tR0eeA29rEdTdjRmiYTDvEqq4Ik9AcR53dSioVBb
bt5zxfSBjq2whfxRwWdNPJ5vBmitRKf7CuRT8UTiAkYiY4VY+KK3xKqf4llTEaIdsRygHC4Zn8XU
lQPexAR+iwVvt+4/QwxNtKtsWpx0nyQWqFnvTc1Q9myyZew+xo1x3U8f+xhY8r96aYTO75gt0u5f
/NmZSrLb92Z/eP6KJ9vqkCzqCTRLWM1dtwYZaK9qFELmkGhDnH1BA13ZjPK9/W0Mbm2erK0shWS8
0seluB6t5nKrSufnV7wzrsWtjRxsN2dE5aR4cPWwS06B6xcqkY/G+ej0cJjVs4Ra6nMobbtu8FCo
5JRGizHv1Gd7OHzSoVFjTCjH02Z6upLpca8Pb0kAFzzgtuPKGQf/NWZuQqakFTQyIgLfp88dxGu9
Zlf5NcIcIYhpJBEbiAZhHXYSZOGnAbRDqtIkM4w5PeY7bs8gxGRBwoj0SRYQP+OJ7tz3exETU8R1
+YMHd7ocMgk1DFuJdK+9IWKpiz4M/t6liwsAyfC27PeEkGbnE0H1/yyAKwj43b0zqXhUFzmYMjjX
XNPMx5ga/47dQqNQSl/ePNP21t3eNXPfc3I/gytofJ7B0mBBNE3YYDvJN8xlZrQXt9U2qTNANYu/
I1/EyKthOj+G12dArPkAt4kIiiOlnA/TrJ8aNDtg5atonNwQUw6RBmEx4pGP3n/S1SuwvqZYh7p/
qhcW6sbA3Wb0PkMX5vhVcjVtp8uNezlY3zfXivhFdYzzn2fsZ/BBuYLdURhUVlntuckyTjynqNmq
n4eglgzJV7nYl3sBQnFVEJ1oY1geLBshK4BW1WoRpwyk0o1vq+GFRgaL9zCTrLkiAWffKAu5a57M
0NxWuLeG6WDS2LWXffq3On68E/IYN6onabZ18tp5RzbUw2k7668k7NZhx2M6Qol4HBFmvbc6pXzR
c7+XItp7OvJTz8rw/OUMf8HHE5G7OxQb1JzdVBBdzr3S1lSoiiWXCgnaOzlqZJVdxEl+tPspGVcJ
7l4jI5EIdpSlDdurYVifXteA0XDwcWA5rbh9hqZ9t6diUz2KNaBVvTj41KRfSlpwrCN0RfRE7B00
UQpD3bmzqm7iOLTT4kIyeGWpbR5GO8ynlMINeD+RzSM+IXOzBisIoeqwb3ELOnzEOR4fT+KGkBW7
DWgt5UWBa+ECBVi1RL+dmGn6Bv9qxm/1kxI82bpipjBIAZgQYDUubDEH+F6WH8wQzVyTZlphiR9S
c4/7Vs5m2tuFRtb9lGjPe+cw8llhVTPxMdM5XLFWhJrK8Uun8SPgkjzm9L9vmVVBBp25EswfWd6h
WBHdojZ5WyqCXF01LnrA488eBBXdeaUed2FBo4jSZkDm9oh8vkYLeEFZhrHI2kqDecjDLf+9r20m
HD3QbfRW4HKQmQrpqOZ/9tx9Q9got5AQbY3ILRhahGfiD92iax7a+H/UXgE7KX+/cqaAtKIf+e4+
/4bGZwD0vXh04z9mEhb4Gy1WJZIOfzJL9WaS9Ti6Xel8+WkTVl6Y3yQmlWU9V1MQpf27ThDptxPa
srXVwpFakvzsMyxgUiCtSLxDNoM2yvj0e6RZafdl+iV/R4TikVdEyFC8GoeWgvRdgni9VQx+SGX0
BubCfGhg0gV9Lk1HXuaaW2lDZtq60QV3rMfkXisgJhmwU9ADoi7BWLdtvrNmTX19fhKIBCTLB26x
/w8ajPx+HoxRdtriscoEdEqwmAnNB6I/A+iv57GbhRNN5ykVarZuTDH2PRNrJDt+yuPxL4SxiSaK
A3IuHDYsGpMJNoJARK5egNVQb/laux5UE+yU0HP/ro2jQi32XUAsYOdXFMGwjPzgSJxqvV/ZhE3N
4MmJpDKuBA7sBqx8pCovv5RlR8MJEq0BjUc7ALnbk9yadGG11bA92nXMeh5SyjBtZyigSGSqK4Nf
g5ZiyHb89lSK6C4lpTGUUqomkr6E/OycR7xZeJFrCqkEEnqm/C+B6OsOvJK5FpRUgrCL8rORlCdd
9bRp02/8mdQEb7/Nd0CHNTkcFTec5eYkSy+qZzoN/XaL6TNo9ZjMHgozNZY+b8r3CN/UAzfADztN
9ROnFZ1RiC+b0BHhRNioOMG38WpNq02Kv6iUF+vKlCd6yULMUDPzMYsObL0uIANDX/zqCV/yJtLf
idVzYKT9xy0Xo3+uJTWBOy9d8XU/bX/k/rRJovRChTxPe3YuVHAA3aesphiIOONGiSJKghMsg4f/
mDHQoFpr4UYjY+D6/JhHNkkk567NbA1iUaLJZtt1zfKXUyYMuvo6XDEb6TdCSaO7qyRj4iBwWdhL
WUAWsDBT+rTSlzFOhAxEfN5L9Qd8hgAxPj99MYUxRl0dCJGeEJnNxQ1iGsLwc3jYOCEbwenEdL22
DRQVCEjHIM8qAKx50mJzG5zi3sJ1+iS0YPGnb19zKPBhtuBA1sp8pdQK0RwrjfTON+rUquJFozf+
HabLuwCOCVCLtUIzgsCn6QDEUCn/J8BjQDfqZLvIc3kWZwaHCeuN9pI22ofxzPiOI1/37W4JAqGf
6PmhADr6Vpq0BtUcYjKUfPYetghs6EzLEDmYSSCh1sK4l9yOnuBHFkTCKqG3EOxq1Z6wHSb5scnn
JboV2vByswIKUbkDblwphS6DoxFXL+pzp0KE0QmUHM2w/Pbye353q26EdARuDZS2h5/p0YveG6sn
rxvIOf/tfrT7yGo+MmP4V7ux0axGh9nGLWlNB3S+3nhlESx7aT+tFMwj4gdDRUfCsYtoHtntJPXL
4qjov+NJahdvzNgIpqGkbbSiutAuHGrymsB5sQjHxhG0NifACf8KVZ4RqirS18bU6nkcYB7W+vsx
jnS9b2ImVXctOr/S5c7HaPldrwRcsw+Q/Ifs+mGEHKndeUKWrLYIwIY/Gkmb/VFEaI15lccpXy+0
ptj2NUL4VJ8wUX4FLNFc+W2nn1VFKjhp5AN5V84Hr7T20nbNK1hqUQul215vVh3mHZBr0zc5bcQp
CA4tuW3rUXy3qO+ZNYalvf4eJ+dr4pN0/15oSBHM6OoJyupNdn/Z+cve4WmQ4igulFz41zvCP25t
gI+wKJWUjyAscHj27eNmkh4Ew2HT7zP/0OYMp3WUbLOWSDHhoVde23zi1cFVweZ4QZUMliqbUOGt
ph6VxsDV/d+a0XLO1Qqqap++XcVB9Hun0PJvWbSpbj/RvGOF3cwkxPzZDabg98DNQ1B2ND/MT1nX
0xZqnx0E6HipLzHD7vAQt7Ij755ZSGx2zM5A9pc3C/jWxFNPXdyJcB+7ZxCCEfx33OGAO4DYl2xc
QJe3fgHJP8NgV4+0hfa2oK/0SCZMtdmRaynh9M7FUWdDVVOaMaJVzxewJ4imTENIFvu7fdNwW7uk
WQuX6h2mvayeBoZs2RVJ1+L5dOU9tSJVPb+hKRxR2AnEcg1zd6rjals3AHtxgZQhO8TnvRkzClT1
+HFM/jItw1/687t02V78DfEaZVcliEXnsVRVkOy2GwvFPY+Tcyw22TQruIAstsXmtJFHTVuQa+pJ
FvcK39YaXWbANYquU+8eg/WZ11DQMyCTO9Pl6vOaLVLsF3ji9gkcgP8uWwC/5Ti0TSg5XhpY4k6S
T7Oww3sKoFOCs5A2Zkd+4lzBoQRUDQ6N7TR5Z7NUQtxhisC+bQNl06e86mhHUuDj3RPw9Sr+WAK8
SAHtHK2n21ez7S8UUuI1TXiyb/JSShwYrwjnMaiW/Ge36Ueg2P49d6PnuPdd36mL/a2XuGK4Hbs2
m5yxMYqP7KmDvgnh4RrQyl2WY7e07DtHnIUTRvRCix/TJ9rGafkurlKhC2pltIrWa+39t1sqVDSD
Tr6BbzvF7BY2Gko38rwpAqrdEOqdV3HhNlESD4vq+1d9mFheLvudR0RaUwCzLxg3a0TXXyX5OJLy
6HeEYVBZLG7MB9kLcqUKuW3CnfnxAGDVhhOM1Wr8+QBoMIKMC/VaVO+8mHhYvetPCEwWYzQ6n9lK
eRHpEn97avdmW2h31eQYF51qR+veG9gPz01Ka7RkGeGQXoDzlO28zV8hDo3Pl0mH5quKfn/T+5i2
U5tLLf++spxThq91qF8nHQOQcfaQEkExev1NR7AdOk+0x34JlA83Z9IwYG9Om73Y4mtpnJZWw1ke
UZkhsWrr/fhP2y0Zfcn70ftpyK1hotxeviRYwnGhezMIIe4uqd5pwh0BVE7PTdf35payX/JK3IZZ
cxgDNG9Q0lmBxP3c80Sq7rZ66XviqJgEeVwqGtc2TBWpJdVvtJ7H3W1oSeZHgEl37G6/LVl64sKw
af7EBdAdEmizlmeCBDKh/A2gWILE4c+Kwpbjk6roIdPZ8DVoEizS6v8EHNHZyj4QF3Lr/biIuz0q
KE7+pGWJwqLdecqPOBoyuMXH51W1zp2rajj+xRcpGG2VkBFVOubFX+kMbUsIOpwubQRgw22oTC93
mVDgsJLSRNp0MQJ2agSFL6D7C06N9cOOoJVDRf+Atto1kKEt2Y9ekNE+1PSb9id2y0zWXK4fmKYk
NMZV+8OEa7fXnuEMOAuzQfwpkk1hZVKMpv+5w4vGvYxhBZk3VuHvoLI0S8/wRzgp/pQcDS/ikU95
HBizMFETHzqcdkuYb0JGVbCXJKfjXfVaA9rkPbaMbsB2sIFPB93yqCFJTx99HfwbPQMkYA/StVEr
KgMebbmsKYDZUar/+DZUic/lCDU3AM/MnD3qzWaMKz3fdEKNaAjh3g60Ks0tV777qCZKzeJ9d81f
GI2EmbXjO4RcwuI63hTJBjc2zCfgG3gQORkor6gkikPOd09UgtCeSBzF7wvvecUmnHdfu2Co1O66
fNysgfstLSMc2RWZG+28TcOqNsChdtoPO+F38xvgkaZBeqCkrF11WoB6FncH508jr0dmG902n7fo
i9UXJtTtApd69Pam7rkRwz33lTgZ+Z8cIXcur1NzQ6aeretHnIYmn3rH6zHkjhLN1KNJp+WdChDw
9UHiDVLmEiE0BR8F9Mal0GR5VJzh9GLS63uvQDhO188ldGUu3l5N6zrybhLMMQD82PowCXkJg1hK
YScvCL5GBFAI49emXLfBfhi79qNSWrejPjYnod7ExZnPJ9q9AUZvuDHnRugz3NY4i2AZQAOYv3xe
d0OdtWcyVuMUtMUoixJvdv6NnvB2buTwNIgrDinINpHzNZiYGs7Ec5k+5hW4s08Bh+DLh7AwdoyH
czqEBSQhrVsoEgYI6xDbHqyEZYctDCVdUJz2rnz2zict57pzixG3Op9Ztif2rPc/SFpvsxQRluiG
Wg39xggqfePjTJy3wC7U8MwzlmPuNkwNzGUo8Qh3nr3GPjUVim6wgx8mPRPF7zvuJg8MNYbA+Hns
yz+cIBuEiMsLWKOkUsgDPUSnKJRYel3A4DHxWtywjM44wjI8SkdXBFnSAMiSkKMrtEGEaYWR4H3t
CiCLNGGkfbxtPgLDEqZ5ukp8hNpSBRZHE9l6BFI0kZOUs0lB2oo4RK4v7Vurt5RfgpaMNBP8CCgK
ABvoLYg28aon6FeDeSc2OWksk+FSFoFubZUp8+iLinUbR5YnPfktbXGJvLNonf6TVVcFVzkgwD0R
+VVdsnUtIXNQ6afOe2RpvNGFmMS0tnldhxE0qLfhPPHR1Ep2szeDGXTgvkSxX4+FxPhET2zsKw3b
IC2Sda/U6JPHCrxp3qOct/pHvr40cJSFjaeIm5jOBj7k8xs8PEYpzO3bMdyQDPZoLiyngP9wWdhK
ZtMli+6nRyiMea3j320/D7S2RDuX7aGvn4B/uCq3UaEkUZwMzcoJvyQ4dv9kXnjFidlFdtenVb00
ffU7k7J3hOFMtV17ooefeVp1HZ/8STrBEZPCuTI/arMP5tIuopJafMVxxHspqwexpWxu2g6lUfv3
LdWbxclE0tbAIXUNyt8PLcK8la2aqPykfE7elg1FQF88/THZbiX2Mgk+edO8FHh0ZzODlidq446M
pAgTjmkbR+WaiEGeodQM+BGnS92YOQsdamolv60bvE3ZDt5lA9l4aAj2cEawf/qYbmeZj12QRbrO
G6XEKaiRnGWycOdOiI9egiR5AFEAPJY1RVZ570gwiBrnQlDMwBGH4jYYpdJImn5Om2/qTlv5R0ms
diDysi8y3wX34L0Jzc++zdJ/jWYh9Mze1ZEZQQvDzUs+guvcNRksFeUjh+J4ogXxTpdul1ejmHQg
sVEuWlmQ/jfGtCfTcNFtcieyupRnR45+BVA5+c56Gs5RcoxI5CFDGgTUxy9dBvuDv9xYQhkg5KPT
CDvQhNuiSyh89t1CHp/09MMchhaZjIVKAvvpxXkgrkz5JgpkYfBE05nvijNatFIwY+YxDqBazz+2
a/d8V9QqK/Sd8Kv0sjpXNKtuCfaNhUcbKS/qqdCbgXxnmMh3OZ7zkr+PEP0JOW6NYISwZUr9sHbl
Ofz0Ecdlek5t/GRD7+Ny5llv8AKIDRAZ5n6harMfyQb+KTE16nNbikjhTVj8m0UMrIcPPkxsw/Lm
yBIYX/iY6ipJtZ31qrRS8YBlmSs2Ma3L1s83cqEXO9A0T0c9ECrApQVT8pqkmViVVoINuSFQd4Qk
A+g75fFKBnmQHmPutXeq2Wzpfjt7fQhDGqlVCtkDjJVa3XOLk8EdE9QgRdvYzLIPHm7jfMPGsQX8
UWnaknM8d5h3d3kPsK7q4cld3WMh767dahS7WBX7ywMeZSi+yeI11PMuMyW0dYfuVnHK5xbXZbyS
DjvqHaK4wQ4xgYCY52qqKMrZXJ6VF6y5eoYH/Q+mXvuv8yQsA/1GrXzOaq6YUpkr2CMOj/2CZXkF
lz6RtAX8d8FENbzEzZdh0ojoKWLlwpnbiOaRc+/W+1y+Q1zXXTvDsGHt8CImQ7hliqFWGmmSfnOb
9C9raT3LyZqphEoH9ualkWPAuTuKdTQEuLxF62iasTmXQTqSg7lUrlmNeSdt+lj/9x7X/imcogBd
LTON37AkzV/zIkNvJm3xhlyHwmb6WOab04eP66V9x6W+RZtPoH8xnrOWPNRQ2Mz8qfSKqsenKhPi
rDUxN/mTu0BV73pV0zRxaokFNUviD0afz/FMZfWLIN+1XL930qlZsAN84VydUCHl6jP6C5ztwy1K
JbQ4BSAT+OLhL+Z6SAeAK0kaNwq9McyTx6iCT9NfpiYKvqZdQS5s2f2jcJSYdP0EhGItfCUOVyi0
+sEIiCKGMsnkbADyWC/TocF/fw0iAnDqN1nJWWV3OgMB2tYzDDI6AJdFnXDR9NewtW9eBzMGmV+q
KMswRVKfiFeiNuwmy3c25X8EUpnRqe7uGgTo6vXNiFQz/mEAcxF4FJnsRB6jqoBPNgj6H/S+vN6+
MoV5xgK1j1lRh+5YQ6FPeCur+8K7qGRGDtOgjrctWeeCEOqTG0o7PF6bzEUE98bzA2Uth18XSXwx
t6wAhFcQcmskSTJ2saHZc33ZZ7guOXzrkfpklr/u1SWqK1Zi692G4YQMzL3nFpNlGASRfwD3ooqY
SzAe1JUCr/pe3ul4B0x4CNezxvS4ld+hZMcHdatZdRi/VDnHFHd0lnA7d7AjBOE/AvYb44KvTFe1
5/FdrPyLBVvznQ47Bfl9x7EpuCEcbmQUcdb9cGSWCXGxHVE0U81+a0ZfrdEhCVEUjB9S5XvHW7wn
qyvmoNlj8YeNWaGyiNsRVea3srtguiVc34p0z/BXaYfnv7rpCHuF+PZmm8AJluDMHF9ClRs1vlxP
0FpBkKZ92gaHDeuMGL3gYXOXQu7UgpC/Yrc4DxAa1BgWLOgUMbgZm3YgJTwNcSqVg3hftI0JmaYU
ZPmv/aODdY2t9JtiQhUYhSiZex74+agYjJtUVGt5CeOK6j5FtsFCBMcCkMV2LneNi9kB17xVYS1o
g5jvVoJd6L02Jou8LhcJsgGnUDVefWYwuIqDSZmvHVX37NGi/D1hDJQ9D714PAql4JpVqwzBT6DC
9TYYfleNiBmQL3/3loqkJsrKqs+KtyYHI7hijaKf12B3MdN18gKFBeN0Gv/0fGQouzx3khq/Batl
RnVpa6hoE1Ek6SP79bLw7PAmiumyEnrfm9/6mlq9IhzV9NghMFlH3d8QR0I12HFsE9Aea87XC4B9
PaSKNYQa0aNj/uyw7v9GfLO0zwPmtM4pJL/70KAeaZT2PyP27HztJS3Ru9pLp07yfLr7A2n+tZCi
R4bjFD2zqrj3QQPJ0o5H/ZjfQs69po2bJZawqtaDcwCAAmRN01N5jJrX73kM/T/Cx/ZcSuJzef+Z
xjjXvAJ1ozuapJAXKAP0Td6msbt5dgfd0Le9Mfu43Rz5N7ik41nx66BujkaCxrnLI1G9dpps2da9
SMXf9VtVOkMUG7RimlqXKeeGXHJb8UpvkW1OOLrTma5stI6abncev0qIWLrqmDahdk4Zsju32RiI
W92Ze2zZQAj2nlI3XRYjHRH//63VK63LSjf+Av5kH2VMMi3QH3xrFbZV4++I2y7PyYHqGWHKmFkL
lrxfYtMxN/LI+3Xo8PSu+rwICyKA/UjJLYOeW5kRwKv/yyBfkn4Ke9DRoOdzlhFb8nR1wN3ddDaP
Fw96N1yGRR3g8BtexbMDbWHmM8t96aAJYxLL27ndMRVR2A7od5WabtIx5Y+xkeCIFzZ7Ej5NONDv
5w91jrjuAJTxuZvXzGzC+jvcAoDc6O9uoTDVEcbcTebW8PeU19q6t4e2pnSFpFEgi4FoCIvrqKYd
M6vjmaqLY2weeMcgXe4bJ1i+M+MRFW0xbvqdLeb2kNn+AaO1/kH7WHrUu1hnWyYlds+XcVo/7CjA
EAEnpIsthBqxiI3AANSpMZJapnXJlMW63MeJ4yvLUOtfHiz/pL4FhhROWZIQ8DjfPmzTj0MxgeZD
RfdLsJnoF5Futu09TL/CSvbupkYJhFCGcTc5ujdNBL3rlZmlz7nhqZPgoFfr+IDSsvJ+hPjEKty1
UdkeVnKs/XzoQhthI7BuGtGOdGtTdwo6tckjKCnDM1envOnpBIR+f/cCrBM/2XWddSUQAkS3kpe8
5tyXLdRiBeaP20fbaNvQr2GLhCry4AJ8ARpVIEGjUgBqZxW9HpQTf8Zv8MuSiBA1gOD4zqJQNXJ9
ttTzPnnYqmyNTXlTeme/xtJhUiSI4u5wtzhxkzQt5UuVxiIw+falOtpSq4JkEf6gQsk7iK1BKz4a
7BKAGhRSubToPCBvI4p3UiMPexiYuRGBiQG4KteWoYGEMTxOjJ5Tm79miBY+Ejp5RDIt1dEirogG
u6pVD9VZ8JFS0VmCJkPFWZV7PkYmK+odaOSrcYNzK/eGkMyhuRsAwrL7565p/FpWq5weQWF58v3o
CjmLg4VuIHAckDRWSQx+OxPVknLDosjHAyGE1w/ZEruCfKx5LzlTUaWNT0llXcm7T8b9VDj03C/C
Pqfqirb9pHmaShX5QtQGGb70yjX+ssWyfH8tGtgAatFYqx5+K24kqcfJJpU0wNRV7fn0P/EIRYEJ
TV7ApNIbyl0Z2KTTdeoFXhosU4VWNkh6+7ULoo7NA0fXgB01cweArA1xWzq2SC7jvbmhxbY6taV7
yrf7AJ+UaftX9aADW0DPrQM+isNJFP5Ft2NXCDXGtSyd0jUMumGZQtY60fLmb4Iet8UHYH6D2nOQ
i/pLcf9JnN8Xc31wlgCNLxilXhhlVlHUaW2xUsuIVCphr5dvI5FyY2PwOvg/68f71hZzboFvGadn
e4J/YwBAuj4+jvFKc9r19pvcaoIdbqbU93HFQm13WCA2KA4FocILFTVngT0oRfZURD7jGyvVkGKo
tAU5HzxsLTT5o6P2rEwln7q9tx7yz4q0AeiDXhydbS1t99niJ5SaysaXZx0GMw1VDznw+S/8z9Px
WAK6JrP50/uPjYhuZpvbUP6j4M2huQhs/W/Cb622HD/EUIvew5jh+xLsEZOlt8EmptLXX31Ho60s
5YVJ0n/GaUj1bUcpXeeV0TIPy8bGHa2q+WxO9tXTi6RLEXlBtpwpO7rCSC/KRstggYKRoNo8HoYn
i09fctviBB9OhirV2h5B8hw1kycvxcFwHblyh5epC82eAGuSvTy2t/0HweZXrEKkeFLnnInaKsx4
xlSoVE/58yEp5i/r9gAF82lXMlEaohXnGVl0V95i4F6gWvgKKy9AiAON7OMUNng2vPwiBYrTfSYE
y8kaTH1z/8/1Exov7Tb8TJGrz4sAbngD+HMm4kPlZTOsOEBoAcqy4Xhtl/5jVbGq4088MoCP/3rk
zj+Bu0PNTid1wPTmVS67nAlMqZFQoV5D3zG1meT6EqBXHrOcQLiJV1dAeSF1SE2oQBUaeLzFBYTN
ojVLDQG2HH+5Fh7r2e/X5ky2+0BPxhGCCJm+uElJwBZgm8toFbkcBvpvmvVsDYrjuEQn4/yXfAzc
5nQSrVt2z5+fP79WID8CcpaIH3NYm49KDTYN/KiRztpGh8DoqtreW+SvR30bJdcA1qjqW8sKAg0G
RnOSJQv3SzDLL17ESUrWxGxVduBirlUDLTmjt0MettSu07Kg5S47A0m0prLCBMi6QPLwl7+8laEU
OB99a1ioEttfmqeqeACo4uMU7+ifILjWt4nIJiflo211Ss7zjmVAe8WwkJhhLTFqFhzQV460Baus
Ws4mPyS3VOdvxWtVtXTJykuYreFoEZ8lFKmlb4AFrwEKl8T9ljfqq80J2T3jz4Pw7cayRNr2Nv8i
VbMf57wlrNtWBvx4QA+8KHpUA9d6mHOJM2YCYKi7/gwPYiWTlv2KB7ulib8LfYOosmJn96m3aIcG
oWoOloBdzTdPJ+5N4cZ8IzP3N/+gPugVhzWj3NS/C925doNfSvMeEobv1Eix4pOuuAsCcLLnFzXK
UpcsEZiHktiwMwNbla4quVW4BlHp5nDgFK9h7A6PpA1VMIBzz27ksNWTbdSNh6Ps0Ev6f1YPHbDW
lvyPHILDXzRmWtI+exbPC0hoHGM07n5sL3tbN00xM14GxW6qFxloYynCzKh2dMdJc8m/ma8qOVnW
BuTqfrHrLix2qlK70Mn2ouaTijKA+quCBi9RnRAJD+GnO+d6AGc0sDWVq/WS0SW+qiuOWyuqXtKM
SO6xydsbsvbAaydbDxky7C9ISV3GPI8NxwsdfAF5nA3VA7LlzsHELi1y87MEuA1r0X/yners8zyY
bJ9Ofq291J+fahh3pL8dHecfXwYzAcUWxXvwUvV8lQb1R2HPzNYQ2vvU+7N4+BroNbvSvJHBIzDa
042DW9aAi7+fHDrE+tZSJML/eZepHmRXWn0A/C/G/gBtGW825AH9E+XIq3CSFn01cHo55/z/Qman
SuNXCFsSOYUpnzLNnG47pEw9do7rNd+wgC9HUyj3spBUy+sXhHZ0uV6reIzruoATi9SL5HBkHqtr
92xNKSyboLqWfHqDgHWgllPKdXj7L1o4nNxSeuCHysP+CYi2aYOatDT6qDr9+xHsBmko9DdfTAd7
KyMKn97LDT3dWHwNxcU77RvLrYly+H17DKvX67dAMofsLZHV/aj2R6/9Ow1a6Mz/RbC0GMz+g7iJ
1RA06wNdgxh7OzGs5SCIPCQyrQRTIQre9GWPAY1WUtlga0LIQQeDDXrUQncaeeU81ZtfH+hsshxV
rw/4Xef8cmbfKNtdCslTvJLngSJXSv4BL9PKWcTAtpVPncGOCCdkgeCvl7UnWhI7PB3F2p+2HaFL
/j8ynnO5wLKi5uJHhjYVXD3gN4tnN080Zrd/Jvz+C1iWIqbNHNJIguOvJtmEJ21jewsCvm/llUHH
qSTKgjgjMw5Z7YOvrSzEbn92GdXiVoCMj+FL4JLxZh7Z+ZQ1lrS/HnVKhsDrdq6BuwKak7RS9hBQ
X9wWe45XCcunf1iY/eJq9yBMczxGERGosOtwX0DZHTUTssWlrePNVngPCQ8HFjIHYkt7ZhBtoJCw
688MvHtaejNEhPRuaFBPIsvrdb/XysXYIEs4qGM9osiCEydXRSilLGgFpdSU396VFg4LwEWr9u6j
zlI6vgoRka+5Tguikiig0RsX2LTV0FhPraAKhGZbimkNwPsLmnDVKZVeeXWVtYr2pODl1pgV7wya
Gvj9OWAmVezUotzjE2PSppaWqvN5Hxq9KoQe1N6vlcCBNxu4x5gamgQEt2qy0bG5CcTRF2mBV4Ck
S6oUToKqmcxfIj6ahhPF6m51OM/yaJCejhosJGVkEV3+hivpUl5llcp0Z7MZ6dYJtMLGT3p1a8jo
k1qw6ro29bcxNrGYz+hQfhWYgRC/e2LlimAPJvep5PGGlhn3vxCj/X5sZEww15C+X7c6Tj+DyoOX
fvd2uODylNvxiAS9QkN4HNQLACwOhgYaHlkIgvdyZd9BNnnlLBvfdhQiZ2UdzMVkwS9OiepH+/Jq
bc1+f6h7JlctVtqRVmCFYdHTy7fcvzWo3mxVUdogHCM6JSxe1BwCZzW25GYi0YFPxmBtzhByLtF/
jkQZ07b6Y0RVQhl8rKbjnN9zC0hT3IMYrEm4CE0V/ni6huUO+VVr+h2+usjQ6mnvX8b0RNjZ/vqD
N7mV3Gn+ZtESMOYNIRhgSdeZZo0ngdajjzrW+hvO3pzNE5xhs7x7o+6uVukwgUBNLe1RtVF5qIyX
JVpnnOCykw/NrREaQaNH0fj8AhGGFTxNYl8NfRCZ5X2hnWu/UsgQKwygv7AT3PP/VdB8gdsiTY4F
Bb+ICJYuRkwzgNLfiUf3nXOpFWjp9C2zlK2kGnKgc32BVrPj3Y1g5HApvhqGIfqfMDbLaQukSF0a
QeS3XJAy9xnJDAa+3vvfR6wv1TYBoUaHNMZpFCmn53smX5gmI5Ms8eqysUzegzJ463S4bgUnRjNw
OZCrH5dJRxFGaGh1m48uT+i15YC+5BRUlDo+o2kbFeBJ2w4WA5O3AUPn0ZpPkxpVzuGBiTJDdmLa
U/5Du2ebqOFj0MbbsFW+wzpuZiXQQHTM1KONcbfwhJklo215NZiOixef5uuNoNaVgYP8HXP8IFz7
xPLc/17cwobF3IEXkS6Rda20BvsQDlJBZYv6hiN4SOhlz+Thxw4ikRx0iTkCivuAeIpAU1fAn2U4
cobzzmYWgH3W9qMpXZTxiXFw2WV/Ai38lrTHFepJwtiNy+HIHd2yxSOOSm1kRGIq5kYZKrdoyTdd
fLb0oBuVra2H8nCqtoUJgJmBUoodvR9mKritCnmFbrD0AGGcnr8Zb9M76Yrk2I5Q7+XkqNggoHO0
zjQfRx/X8Nj5rEssbJAhE9wGR3MdF3YpO342PiSP/sy0q2U1F8Swkz1ByLpI6rByozUib2kH8xHf
ONrokBpet3vHeEkAOeNQHmhbArdOxPVvUYQHoJSJ5ImwKYIgBmtcNtdbc3qlBCl6lXTrzBRG+2Dt
8p9kuaESYci9eFoMDpJkLWNCCviStIfhpPRz4nYacwyRVm0qnVO6p6tVnnt1Dp0sZO+wbY6wbsDT
9ZjclKjIsad6uYttjeHAMAXiSVWmFCVqZfcbYO594GKfX/HMRdqC1qUL9uDUEIgxuHnr0SZ25q/Z
QcUr4XZeAS3TTlx/I+DkMFHyN84DeVzQffvCieQj9xXotFnPoOof7jOk+lJIx3JreemsENjyd9O4
b9zl0bncH+AOWxNI02LbmBh2pt1j5VEAGp9jhShJC66Qx9dmOv82l2lzwM7oDCtG98hnD+ruCZnx
VcM1zv1dmiep7c2uStojDrIq2Y/b27h0kYoFphhTxXm0PwGUilQs59V6kF6fS89cvkqUmyY+B01S
ZArCH/crQT/BE+lXceqRXq8O07wd5B+yAdu2yoKNfrnjXL1ucun4xf6YYPIcVJRjXtF/Mft/kP+d
sXVgM2WW1CybU3NyKWWeCJFouKScrUuzgC3imNJsonB9bdXVX5gMTpEwpRqxvxaIXQr9dowiCHGj
3QvE1XgRdsU6rvA1OVORoVQzYTNOHh+nsaaFV+hJU+nhUBty5I9oHyrBHrFpqT/f7flvJ9DCkOKD
gLrjIshejaJZEGpr03lvdEXn7ZgUj/TPYkCxGm7dpYOwIUGONZf5DmDaFhoRrLqESHsLtdUfBSFD
rNomnWcYRyJkVXjxoM7VzF2AFnfJQJGzUkzbfVN12In/6r9foDwsQGFP4Gc/VVdaWuI4lgsDLVVy
QZbOO/TjrKTFk0yAg9fZ7k84jeHqhMBOGML7trI6P6Js30njny9Rd77OpUFT8AuyGxCX3+nAgXZD
oPYmP+IY9t1+buR3PzEaTzeTqcon3q4E6eKcDgqfEbJW0UqU8oTABDUmXhjxCiquGKkyVeeqhddP
sgf3U0M1+NJvn2Egm7inQ8bgmxPnXV66hDFL1Jqtonk+2ZBOB2+GBHAc0G3gTXCz8EGotYXwC9v9
UO4S83rwmFkIwquAIVsCd2TFGehVpmEXeSYYZ8mDeB8A14IJFedldmLgnxGzp+ir3AAjP8gTWT5O
tdAMBAVWoOD3waSIQCGZHyj9exEs1xQM+w38PPEBTJ38fpPEVz4aysNKPn26g5tUyd2Xdqbjdz/K
UQ67wako8W2MP7GxChKa87AqN+1wJWiaudxwsGDGn2uU1osfIOzLfRgXE80xiXzUs+9xOhtdn66D
M+FZOyyk9cYVNBWU0ZwCa6NlQ0Vx5PHTThVJ+C4ZJpdzqhKqFvjp2asSTCsCjK1ZXnKPU1o10usA
KPpAFYNplgqn1f/3RsAcTm/y1pRkF5WDWIfLI8fDPr2wSmUhpjLiU4uTsOUuxMIjt5ZEEjyFlZ4P
OGJQgOcCMOaoeYz4eh5UPebEvbYycPl+a1jt9ZMy4AtSuVRxahlO9ZQYFztXmjTeEQUw5cJCwgxY
u9w+QkE1USzXoW6SfdzsCjeGXNYYPB7mNKIT4yK4h4YIAJx+XGtNfFeARLVFZLdVeAWYitU494I+
rem7B90Xtkvx2bynRoRM4Jcs+2Sc07vlwfymvUNdFH+vU2vacBbz4dBqugjQBv9AIw1FWmnA+jgk
4wiUwRVHz/SH0xkNg9Al2051Gi6rNnxF809jFx69tcro2sxG6Hh5BHHA0AWzTrzBipLhNb4KU9Xq
61nMr2VqIbfg3y9a40EzDF7ZfaMoVehM7yDlcefK4sjqNV+I43SALrWbPkvKP1Xdq8RTf/+V6Dx7
yVzd4GcqQl4t2IU7KODzzQbnyenmN+uhlpE7m4atdfLDB5NU2V+2NimilJ09lw4jEsJkA9hrR3VB
9fnqqFTWxa599KSvtnnUbxGESJAvcgSSG4rBGQPPC6hC8p/GjzMvVQkYkWM6r6YMnziiZQGNic87
LuQ0RhogiIriqtVf4ffeIPdGIOYZOfuzwAblW8qeHMHyP/GO8jlUNdd7vr8dovlwvaKEu1p6oqPW
/xvuQ+k2PNF2yWWhIHZUQbe2n01tH47NkJAe4G6a9XA6mcOZ2FU8zifRHa/lcW12aDFInx6zBTeq
kqCjTAKIGMrqjvXmze94Pvp/Xnmj+o/2PTg8P0DBvtH7kcw+u7tPujivBFKRHvOU9VtJ6cQmUeSD
SmbNpg097tCXCPQB/BiILsFd+oGVxekaIYy6NVtDpElP7XtpmsyVTGeJKBB1jcE3PYUG+5BEQZBK
kb7P1xrzyVcMUU7rBaHsBC4oaf/3jZKMG93MsLf1DK3s4vRVi36jFuUPrpzKbDJS4xI9anwUwUZv
qCaP6n3onwhYxtme7r+R+Xfy9eu2LZ5/wd3eGSQfNV+946Yly4PnwMIVzFZFw8zJuLPFhIwdeWSd
PBop9XwMjUPu9e8qXlbpIyJduEd1vyICu60cOB9fbiCAfwzuUaBC8gh+ahms7fo1cJ7genl4ngdt
lse4bhqd3gy4FkuvaygVZLqaGRd0Shmaw8M1nLlBv/8rLNtbJTKX/4I/P3N7mAuxrGQqilnHiGwR
Kq2AptLi+gyF7+pPm8+qA5MNrNDnSbzuWhjxC1RQ2TpR8ZSCakLYocrVEkhY7aoZSK7n2EddRDiv
2nXxiYe1EuEdtvjkJpY+nME8YTlkG/nMexFEH/lhOV3gmitp8Q+zRRXhWTLOODWPwQhyAwySDXIz
DyoiqLnz+8sh+yqkuZySC1v94dCSPC0mIM1ATiQFu2IjRSVENlVuflp1UV0AI+djrDOby+AE1JhZ
AhhRZcLj7Tz9r7eud7+bnzhnzY+T8ISw84tkOq+No+ZwF4n70yNeWCvvbasa/vAvqAiLf+e5q6Dp
YsNQYejoyTesNsdeTAt53f5rWtkbEUesJjZ31sMu0Ywp6jeAtZp4O6RgkZKeMEXLz/Rxo0N4AyiY
XUySsLgYIZhvMK4YNdMQzXjoYNXXiPZfCHttoch23QoEmtQLbFmrD746qBKX92PTTwjhNt7oqk3y
b9Kd/YebOwE0gV8vdYHkUUjt6WLp/IRlCL2e1tBpRtN217whsoWlXXcUfmgcmhllcm6Ia3mXijQ6
YOUxNmXfolm55ErVSRka7xNFPlWqkSEWUzB56Ke+5v6AQUt+YhMnw2i8yPXciJ5+sXuZuu8WDCew
x0trtMo0Hv0Eo991tEZ7O3qoNR3bRoIoLBxb9o/xWONdKpizN1nsuxlSYJcIEsPG1kE/W0w1iVDs
JyJRRpAkVbM7RcTbTgCNV3UQdc+5ydWEEscNZ6GA/P0sRcWxoluRV0kfR2c5eL1IMAfZbq7r3DQp
EhhJNTQh/eqhkdd/Jx5ePr5sVCE7qt5iEfacJ+Z3eZ0VPwO5FOq9wD7yR+aOp30hrNpalPAx2+z/
YExoMBoDey9Heg95ptdpOLglBQ/vhfbQMiQA5Rx7/xEAA8sAtDz1g3KHv0tCrfAb9A7GBRkZdGkI
4mKM66UrAb76ZtGJ7Riyr1eXYQ36k4lTLsxQ/ftFwp+rhJJgUZVnMwE029a523ccXQtoDrJKLAKB
+vlhQ5snXVMk2znZ/08Vm8z5XfqJMwd+oPO6EnKv1PKg1vwDFfw71lEJc7ENATvC9UCALfSedZOV
rfIWq2liuBA4LVI2D1Aels1ec3QfwT6T0juQ53e4yoJajh/XwvlevRSb0UzOTIdAdQNxfNH5PHFF
ZpvpbnjE6jN6v0cxGaeszlbGxJ6US2nQAVZxSYkz05VzDdzH0Hiy90U9V6cEfmRL7AotR3kKSGfF
5GJAH0WRasI4iFcH8sHnl5roz9g6IL/iUUZrwZqXBugT8fAwuY47UZkQlZdvqNjw9ZL7iyUUSpMp
L6dCdFuGTQHfLBIrSbQKp25irU62xEVS6qD+gzeMfVc6d7ybQwuHcVFm+sYq2Qroghd6WDPBa/Vs
tBA4k43dGokEOJ8mi1wKfe6USe2zlLA0UO30SopRifffzP5lPgnOLDq59GQeEoYvpIqY5Ebm92oS
ZK1eQPu98y1m7RRXpVBzmw+FN/AwSxC8GNUJ1xj1HK78xS5NaLYsq5vWpfyz32IhqQ15iArnySae
X/lOyzNR1PrUNBTT/Ebk/Ufe+RyjrGQejbfna0dzza7MXIKNxjGTf2CL159kf6ClqQ+Z/Ay3UPyJ
EIFeELl9ydMm5d7DVdBXl5JlMOUBdDFnKKS34AfluC10WFpf7Or/LjvorMEInIcihqyysTJFaYpM
vW187cZ+D/g/nK4ZYcObfpJ3OpFFvO/NTKZKhRRTmj3Fli0LGyZgle/OgtRAM8csk6bIlNnomFCB
VBpCkhCYNdb0SLH20/Lb5j9B3COjZmQS3Nd06vTLnCvF+PO4UmdC26/SpeWX0G9auqSsRe59Xc7n
ikqzVlQKi86jxHIcxTFiz6doMjaxOMIgV+kxKGw/2hBFVlfdAeHlkm/PYnk+Ix+ZfHQnU8aJVhWO
UkLO9Ocpcs5CgZBz0ZLVAltOzeSeJRF+fPpb01PCmzMqMBTj5pcrVkd8LCcSMQAGuo8iIGU/Nva7
x3NwGc98XQAL0bWfFTt0oqb8ODIjO/E8PXCBZ+PfBhVnnhk0MW6VslAab8Y8X8PO8ecLA+hBh0mT
JRmOS2+Jy/XG0dAnNg/r9xy/btFGGREgWBnoHoZiLpZM1qRoTIUdkc85qqDml4s/ngm9h8MNipK0
ftZ2K+pRBtG87whdaWd4LuGcUkfZxjug8tAFdDn2ikQTqYOlK6ZS8f4U1uxArlGtVFb3D+QjE01o
h2sL9eZ6bsgwDLR8TOdV1tYTsXsKABg3raJpxsGijKiScvsm/lhBSozPYfrK4k81rLnrMqBG26qA
A2nMQXnOZJsQCc/BpRTvw9UVf+Cn1Ya+1KmiXgIE8AIhEo0giHHGVuOVoA7u+yV13qVjsmo5caRj
HvvQu8b0FHBIsAYUNj7udnif1mtR9w4TqJ/I4Z+advKa7qwP6EBshjefQwd9hMQi9g+ZYjIy37JQ
jWrsfyf1s/E6U8Ngn+eYoN3sDESvFnKXgls1OGSNv7VxRgFRHWGFYE7qlmdMwVjO0GWSm97M+3Js
l93mAD8Zk3/0Wh/EKaBNTGzjg66ES9FWnAdOgbNBl7gD4CNDY0z+r1nGZ2K1VnqIq497KNA3f4hg
aOVoIu0FwxO/b4uuWYxlAFRlj+5aqxrseZp6heT3jUFrmSDx/VS8o+CqY/vLfCqO2CjX9sq8+8TH
wLm1tOoFfaZYT66w2PC51CwuHwKmMkus1lgeE3zZYC/bK/889a1D4STIokPNks8srLB/veV1beAE
dlxL8pbznBUuVfGyd3/zZWXaA9V/mkzLpRBf8dbAVsOiYs+7B+VgHxFSVlTER/IyzEw9Cvxxuawf
m0xpOhfrhskLabmf0x/JM24ne0StmMT6NY1okz+gNaOzGQ94TJdeMtLVCLSkFwRgRzNwAJdhsldw
u0md1xm9dxO6oUUuhS30HojE4vM+p9EtRPGnIo6M678VmYjYzOeX/zj0s7gdkEuRe0jDdTegNp4G
6Mm+D/ULr/cLW3Q9t1NzwobEs5Vb2mAB6z5w3DuRpERBA8Da4COiN7oY5a74vToljTAl/eyq5vyk
FWJEBmq/399D9rlu/8XhJDqbbK75zQp8Up52ehdEt1sbUD7dq8j01sMqn75MFbUjd6WmtCgsPo5V
JwBQ7/i9fLGlU+SThnhkCioL5+SFasFRrspetZ95QPNiTSSrVS8FxGetAk07+JZiAKz3L3mZpogy
Au5L7Hl3iLUOrb+Zufno5dhkEjxrKBFncGGLYfsu+rfp8nTEBHl167VOft38X7MBMr8BTE1Fzqiv
ehKSOy5EMUj2iv9GrMmCX3Z+HfQlxovKLfRaoZIqjibJXx7u3YpuOjGsn+MOPESdNt5/2ooGRU7m
+JzOn6zgkPEiRwt2PxoBg3R4OTEjtI9st5H5cITbZD7wWGDsN+Ux7Ag8To1/T9tzCxKCwf8eEqq/
QMk96HvQaVGBRBzYB//lyG5umWN4uWpoKQATlIgCrpk07I3yN4h1rEM7Pr3k1y0+5vbsFAlssxOS
fbzRcbqF1Ia81TMfiIYqY8ErtRZ6fDUs8rjIxmZXWPOqVrx4jrG7GHBIuscJSJSNOZq4XpoeSEyD
Me4lUQxC+b4DfZoBsYIvArpbxZK9pUPfaCNPsECpODdgBDGUasPjZOPS/g1iIHuT+EhXjdD17gG/
2BZc7JYLIaWcX7l/CtLYN5KIvRYNmG6zRPLHnBa/Nm4NlxfQFnGGdmNVBqHpQr9Bht12OJQuVRR9
yfazpSKllS2/xxVz3uYzvha0KaAJPuBsr43KYJfZiZR0PmPasoPLy+5YgcxbmothAzsu9+KjzK3V
6YFqBG2kj/+dz2VSiYDRaNXdklWVDnJ9dPORJeOUB/8uJVH81BRiTlo8gVlTTUpIZPViqv49/w/u
Vkz/vpZVjRMRkgTyqj8m/71ouDS8Rzs0PsdXQPnYYknIGgSMxMSfENekS3bLxM3L2wyrM0aDBnJL
SJc2nlcGgr1bqKoEIl0Lhb790/AW4NA0gpOaBq0zmbFm4Tgm/MN8h4/ZyaiN82nxxByrjqzS2nc8
++zdWzse6SXszc1aNetlsNWT2BmotE++QE3jkPuVs12XKZFrOeI6L6orXCKS4L2gb9fBMKDvfjAi
bP8mOsrlyNg0CevesCib/D7tcXhbtCAIvhw/89FC5GfeLcoCLaObTJC526Pdge58iOLTr3AR4FMz
ZL/HRploGjFJyTvWKUeFNb2u3qoDxz3FWlW5GENEnHHg4r3aBzcdwSA7W+mMkZlHlN3/Ap5FZOll
YPOgwVrCei9+liw6N192OM0n8tkWmM9iKcaS2DXqNh5AfFcWlGltWUM+f3u/37hNKI5t+Xdp1erh
wPdDu59lfB6+3Ju8600P25cWV4UsS9kXBtuZ/+NwlLChQo57SwKZS6ipGFuAXgs46LV5gQdUi98r
DUDWzgVdOSJf5l4lFzkS+MV1t3iNJjdf+r02G1AKXkKzUPcTlTi7Wg26opmP0SJNs8ijw1coGChI
ZliiLjAGOK9JvwGvT2Dw8zgay06y5SO90+Q/Nrlr0zvpwigMY3bfuVNzyWYBBN/cV21t2/LIntOX
c5e4Wy3E8RiB0ETqVYJu7oYtnZ+pjcDsWPWtiYxCQkcQI8Tk03ZWWYzg7uJzhhnPujHG3paRXh3d
sfhzCpqeaTwiFPj/maSP0sIrfCEv+vVeCPH1L6x+CxfkvNJic0exzWnoP7A+O7c9cfjwOAcOIpes
4V2Ix3mygYT8N599iTXCadKmnou+ruNPM5ufskS1ClXbzUpfyr8fMex9K5DY2YJB3HTRPIO2yUtX
Q5ZdG6KEzSA5fCzaTiRdwF3RfSqxbi3exxYmEvkM/7Mc1zY9Ji0HwtiwgoekG84y5Wt6/s09TO7t
2yfw/03jqn+rCEJvpyuEN8irV//CArrxelUF7a4v7Ngjvd5a07ytS0ASVw7gHnquMuD6DjN6ejnJ
8/GJGlJsfK6EsI2DqUpz+AHX4a3odIllQiI8ttJDCqvO4NTMsGXZts3VNOQdmwgczlyybEsbweDo
t+mP2QUozaIPMH6Frx1GrH0qthIzHFxO2i+OB5qduM0jI0YPpZa+4fZ5Md5mAorNJbUT+emaZfA9
yOC0pgpHZsG7waSmPNK42CXxtwK5yDDTD/UE+9zTZZtF6MlnM0m9Pqq+fbvCjbYS40uEm/jyD2e9
jnhcDgwS9kN/ZDVK62czrDtaCEpWxg3kFnmP++o8JOl5kjgH0/GqHzJ3jSThSofRMXy2Bst+U9yO
0Z/PVnr39Hbf0FAsk3muwXUjod8zOFj7NoJAm8bhAla/uP/kUEmVOJJ0jJmhtBZ5zVw3sj+PtVSd
rqy8k5hCQonICjQ6beanRXNYX6cjVxSEOv+fh+LtHuFZXcJSsEU9kl0Febx6mH8zefh5E4CJ10m4
e30BAAReUJOpzyC18VNdc0LU2KbUhSEEXCpfqZq2RAkGG2NcrOGZJwVLS/pChNMgDGcl1bIfBQwj
lSpe9/5kZmTEshdRtPIhSbgk++sL9gmvEGHuVYHJUEb91MTBcu1PwbIKiJBkpqFq+j5dHfGflD8F
M2fq4cNDmpeq61hHKJKzXnmagBqTPDIoY0UaKZeZkUl/N7IcDxEymvGrMkr/78lgv+oRH5liCSoO
Ybk/9IrVgdEg2GhDFur7x+d8vKPGrSn2Z6SssFSJDwgnBIditHSUjSCdGyP8Ql0ztz7xmqfCz1Uf
boEo0tRTf16qj7yLVN4PyjMM/Oj/DtTAVl5hqjHSvvMjP8rZ2Fh/ZmwH7AR1sxJpyxTz/ZHz3kCo
hd2cSce9JKapGq9dC+nPUJt82BIUtIHBhqAOkV3chiJG8HuP8eYsKBNHrd0FtL87YdhkLbD7cJzA
HAjzd1wjWr+c16+SwSXdaE3bq6UrVjhJxXNfDc6RCKg/pTWuU0oP8n8TWwxQG+Q5f9QfpEqIFaFn
7MJ84aUr6sN+F/x0BHbTVJMjFkLZB63EItIeMlGf/5Y6Ydvp8F3drfrOzBv+mo8rGal0XKXdlscy
wy59Tm9AQM7aB8Nb5j/NL3tky5C5L9oa0JI/WSs7t3P1+3SjeSxhuKSa4CW03cFOTKy8fTrPGowQ
LfKkkjSMOE/gxviMLsLal+FT1LJQNM+MUhZZb6Mf/5hw+HNbpvkXkWSXMx6Kh07JbYK/DmMzDF7W
HwIJLtane1b+uXMdoX/Vhk8J4YXRuq37eAuRUcpAc5y0WjA30jlRHPsT9buXezxC88PXXd2448+v
z9zGhLmy7n7GaJQB/830hWdNkXHX7OP1LK4x7aoeBP8uQMQqAvNxMV5VE5wTgLqADcL6smZs7GlV
eY3b8sAUPX71h7e3ubTZsGIXnOUYGWy7RchGd+CSY9iZsZEESKOUbYqtUTebLSdaMXWY6yjNXvrp
g1Hx6COLrkSAcVpe2znLeGbQymKsjPysKopeXECyBzI4xOE6iG+F7D63uIaq5ts4eD5DxkURHh16
gLy6MuR6FF3iw6JssNxCvtwCDlB+hUthVzDAM6gM+9Izfa89mRjR4KWJqsyXDtfvOJHxEKsd0U8c
Ihvr+0triqE9tOYgLw8Zpz0V4PZot6SxQAUkTXydQJf3LaLTqGIAaZFtr5h1y7vtU1CXl1rgakcP
VGZUcXTNF2gHyhF8pbKiRaX2/kCL7PhrJZp7oF+NKvYORcBkQb/MuULhjy5vPyRU/uMtfYa2eR1o
eyOXXvxrLlNnbpOYHRpDy7eDir2ZXRUwtTXEnlFLz0w4U87K8Azw/gRkb7skN8MMdpwPFhQiF87v
jAmWn8ZROGRwO5W37QFEq6qqcxd3KhEysc6ME5wSdWc2PsN3d4S6T9UzLFhJuhhEWCtuYPqMoSiM
kX8o3Q9gZCDLg6FMvzlylV7OvwPG2pAYkW2J6+kDh+bUlisagzpep5oBI9xEQWVviL3nuv4xyykK
f7s/laqWxleS1M+wTvzVkENFQpds8OUo9BaKyDds5tkL7Lh4II+f7HoS06jlh7TGmwS5oJg+ZvQq
rEOXqV2hZPW/V0R7C1TlCByIwhb62tjD28dNnKwiq3Q89HLLW59n47U8ISnV3QEefw8m+gOxQG4T
Eiy3oOSWemNpaxfghX7XJHknTcyU/Xd9n9CM1RdNtjBDjix7eMFUVNkTINMH9XmQjAgQFtxZJ+73
7y27h0qtMdFBFABP0k50PHDEqP6mwgKxo4IGjCck0oAR8dxElfuVbOM8vmpIqAx2AFpUY9F6fAvz
wCslqByGXpauRH0qoxFqZ4Z3XYjiU9cVJ/Aelt3rApKpw7G25y7hn1GesXqDsWCA59Py949ixobx
xwu1i8KB1ehyJOUeSZ7PBPbEQkoXpTiA56z0FProd74IBl71OF7478pqX94vlppdGDuDM+oxEOTQ
lJltpZzNN/uYmRN2iSOP0HPD1d7FBztLzXSGL/kNq1sa7bxfteFxnimg6PLPvidEWLFs9pGbGoVi
voEmBXpRtfZaHtIO62mHD7Ama/rcruwGOQZukzsXfSPtl9FP93kVKXuRNz1hjXznPQAy5LJmifw6
sWxojC3tycmOc8WszGN0gLYmy1tAsEEEaPTOwp4iViS8QQOrgKaBnkg9lreSYUDubCTvCmTWTKnI
9/nLeyyKvx2GPsk/es/uhtKJ3JUMCJY/UNx2T2cd5IlIElaCV+ToGITfl9QBinyCI77lnmxLX1wV
vmw9SU6Do46IvWZyxMdDCeDJRrxhAvU+5JTphvOhNCWprOGxsIglZ1hJ0W/ZmePorVotiBWWDzWb
rAZ9uBUogrCBVyCeWAnTt0jfbVgc8VfiADXLmFhwkyAIKGnP6C9RDIWjVdksYVbkSQcmH04oD75o
/gGHot9oJUNJ0uuBJIApvieMHwM0MCkGBmPv9Ldzv4xWe7jcKKIcLybZlqcjWVYlm7cBw2bYERdC
m6Zh5Kn/FqKYFPJaIstSkXJOhgc1kE7gig736qhUg4GCc/96DTS054y1HB8Amwq1EwpbCGAJZ5h1
0WUHo21kvUYTgLTbjhmhQIUOcahgqphXMkPMaKE0JZD5K9+qlIMXNxd3rpzz9vpEKMblepb+p7xV
PTzTRV922/7vjZdcXFfYlNYmVd/slFY1+ZiSsU6B/Wr8UQUpYOu8rWjx8M7sa6Al031jgSsYkdeg
l9gkc+XrmBzrM6Ld2qRg4+N4up75tS2FViZlmj5g0EzidJ4k/8kjQARMFbUcSDEgdiqJLC+rLuFy
AowslCfgLVVMocRXMpTtBYfhLJPiRnJo2YAvWyHVnMRMl+gqVyI+rJakNMIdg+KIAWMJLFAigIO9
q7Yr0CHpK5KV5woOlBANQllj7tL+6AdiNvWXskUEdW8wdn64oJfGCWK9uyXmbRSGnP245a61Qj/3
ftM/33GAf1pXC7XkE2Kn92F2M4peH2pnM6mA8OKmtS2ujpgn65umsqamdbqWo4fPeSQ27tLlOYEi
kLL+9DawwyID2z/liwSpka7PkexKYInasskbSw7LfnzyjOa9cITVaOkBBhqJmTMy84y5JRyUQ1bN
n8/x//ikyTA/BMPuXqaUInyZPcXt2qhwwNSPEADqL2VljQuGWw8v22hUy7t/ClWrKAHG2UBSw+qj
JpRJFwlXmB8CUdgVvi+2wBHPjlKehMJYBjOmcWLg1RR+pXdqAiPsPOg/X77xRGqZDy+1B2pEjJjp
lX4K01wAuI/ypE/ZNMoPpegf6JuIy+j/uPaQ4wLZr4z86sRo0zgssg5nyGgyTL/yBZFB3FGUjfyd
lKGOmAY3h45QGVRnXsMvcyWqQbXxlxHy51NzpJ1ea5EkNSHFAHrYvnguVjJkl8i7J+AyXELZLGxH
KNRjyY/zjLRfSEp6o9zs3N3NeK0DjGYih/AKwoVAWU4HM4R3Apuy3mtaxxAofK18EDXCf+8iZ09k
fUjxOuEw23Nul2BGvdsWZNsp5mHZKgjvaNTwgeyvSuwAwMLcSOENq/F/o9umuHapjnf0oQNaAqPK
OD59e2eQU7XauyUe7dO3YRHbaWs+MgU1PBVL7VSVHz6Em/w4gthdx1QLdd0JtaFwotmR/XAraYoJ
6gmmhWxldxvIJpVCmgNkIu1v7FMCTeF2abYet6ig23L+XHsXI5pnBQ1zppyWqWYWucFi8emfxfdE
7kOzIh7QxTxjgIg0QoaabNvHMWqApGyvQluAcqzfeikKCekGI/5YSjEt6c+ss/bais2RydB03qsv
q1sHHnww4Y+KZFJgNqJwny05LjjDdHK5jdJvgkkJvvwY3quMyop96kURQ8Oi2jo7KfP9yV5IuBel
yDILr5Soin/k/ZhvQJX4OyC5fOGv9v6n3UE7+rMjrgUqJSm74enAIFNLSgZAgVDLzY4AUPpJAn0s
yKG4FH7ErKS41VHL3TMeY3XdGT/XBnhx8K9MHQu+X2xCpS7aH/hZiT+FsMGBKd/nVSrlHJ9XqHYv
7C2iK6gdzW5PnScqYFvK2F4AZHGlOTEmQOUbbyUxONyngdqkDV71eRij80W2dfWeHcKpKMYZpTDa
syLqlvujTvxICTDY7L7dDEFpd1Edmf8Km1WSaLX2UQypx7R3xGqoF0yO7jcOEEi6yUMkjoEIN/Bv
88K7Ceh/ev49F0fAehDK5ilv/fBVJLyrEwx43NTVe+m5rGl7D1iWrYfV111OdqdJBDIDwEA9Fhgd
+HNsuia8SNRo3mUeEEYgfwtmwi6YUpDhNO0dFulhtAHTj9U+FTy0J8RLEzP73YW792+MfNNSevDt
gBK+FS9NF4Zeaqp0QPUzFFIbqPJN3A4VGUuCOmgOOu79ApXBbp6BdAcqq30E9WS1VNqhwlryvlX4
954MoSK5xsTKoBPutpLiZ4u4p1ZPNMeLiaA86OfrChAcuPd71lzdXO5eDcDewuVkZuOlVW2zfo4t
pgrO+Bg1nVeAFM3zunzxpm+NNKUwbP/DMWIQG4YmJVCaPOTqm6HGjKdJaDRTRiB/omSGXDdGasPM
uYY19anfLaU4OcIPacRfNOWkhtpK0xsWVdUMMWvJu6ti2a8PNK2U46/Zi4nXtQl0sKEPGcDXrSAl
P7T8JjCFHuySu5YAG+B3kr1isyouT6u96XVgCQ7pec7p3oD2nHynzIfVpATtL3utkoyQkAIJ0U1Z
sN590vxEQEf0ryrdtiox7rVssvUh6ypkpOEBRsudL67U1onjiNUbDz8ymQ82mF5MqM7h1da/Qach
aTtl1V/oZw2Qu8MrO8hRPEe8r17jPOr7c2DBfK7zJ8zCDdyLp2fU60DtwApDhHz8oapaMmOhay9y
iFMacIfqkcflphiNkbps/mFYLWF/xwsIbEYDS46mYG2w/c2UDQ7VkdqdEaHqndBjYCCgZqV40++p
5YE0ZLd6HaAb9NblcjCBXZCauyJGrhp41FqSSjh0W4hE6PV/UnJY7H/AyuAE7X08p4Eq5gdpERfy
HDAODRcTxL+2oEsvFzdIRccjojVIO+JG8BPOA6hvhXw3cbEXT3I3nvZHQqMEU0OVxz8Ezo0Bl6vF
TiObECGgC7ezfjfhldJUGlXNEfNmi4LalobqAYX4JFInsM7ctUJNSJJ88RVx3433B8hMLc4Aue+M
ndHMrNUq3hcdMU2unRnSNNP29bM6adWFenNRELlY6wVz+jouueV2CPENsjv9XRq4vPe6fD7h6+Dp
5OyGe+jJL0k+6Utu8HbYa/Ns3KovdOzsBfUnmboPihvjykzV7Pqxq3M2JKlIsKuJae8Bm3nciTTp
jXBHgmc+6eDdUTtf0nDJWSmTzuNtPQxNqNIac6ynfyO8rOM8S6AHgnFEOmEIZYNelpaevwh1FQaW
U5mw+/337VP3x6ujZLi8qm27hBEmtWU6YOqVRhwmpcLORlcj+3nw5opMMpnUCFkEusdXMkKZAgG5
z9Yw+bT7uN1Gsah33Y1cfA2bZiITtO/huGT8s9deKFAKBCZkqc1WOPyIRs26OBBhGqyZ1R1yOSmy
8NiHzxaCDgoyQ/jVZ55rhdYkX3C1bX7cp9A5/NlZKn0TZOCLrVRjhJSZoDXAxi658cS3iKsyoQtp
+1kOp0Tlo2+kkARSsUFxmA8IoKFi8jyhuUXLmGiDDEW/Xzozd84LW6x8Hc5+oULRMckMCrLnTRmw
R3HQrK8p/AOz5qI6p0gaDRBsxibR9T++rwr05iprX5w0bTh+D7whnO7QipYtRtNiUZZ+TWEVCzBj
vBsqwxGXNUWHCIORz9ZiNwtrKdjX4USvnEFw7CYFKyEh1lkmLBr0LZinqNK75/zLVyhCBzuBNCeX
uAyLMVsk12ITfp3wu9BhkO0gascMkQ/dGApficE/qU01gbNr7pZfBcibvivj2fWBROU5ENYTVYW0
Az5KTddZbnbtoQZh0sx6BFBBVz560JNk7iqSj2NXx8jS85BLVlNzww38sJCxkzpdL1U2VT+CKl7s
h2VIvh8PGArQmiCf5sE0en47+tsm9xhhJVSWnfGMiBzi2cTPFTnveNlvudsLCpMxT+/nuxc8Jtpx
gN5q7iM4a47iDeqVFv31HciVlHPSOupoQYPRS/JLtSTTkTgP2T56UykRBy2JyZgl/UVaCe6GGYme
GtHtpc4xZJt1KjRSssg6SuSOVBki8vofCkvIMqYJl8fOlSveJNH0coRSsi13QeaIfg4wWKm6yKLA
r6V6jNoCqsiYl61k9CMpQhqUfVKpv5ukEbBgNIHQr0AkdQtPZ26/tcOa4crX8Bseebzh29LyZe1s
tkvqiiOT3y04SBUyNizskj+aPdEoy9Nek4AXqz7zzMv3q52KyGI+FxKvsp7w6vXxce7K+EyvSVtx
MW0/eRyyoPRd/w9MPkyHAkpevLHVfmVOSypLY2np0KzHKyVCDBLDAhRMIpDt3Eb1jLaMdIvtTSmo
DTrvAKOSC1Z14a3v/OOxIDclz11bbHfcYgtf/mJPPMDUMgyzZ7AinAftJQm4vhHiLsPzvsfVhZOi
iLELwHtEf4eBCInVGMkbHEy+17OEDcfrpY6PUhTgZjAjv4XoBFhPTOgZ9kBJU2RbqG1gVTUojat6
OLtbk4DGME28DTvtFURNqGwRc+wVnLSr5kCwSf+kjbgvnfHzzNKx5tOZECA3VlkPYd3VAEbTWbG0
40uasU9cb9IzDdJ2kztpMorLfqbjMJ3ACEXv7CwCxQihTHSWmEaSZ0E/SVc2vKFpbkgAXunXwILr
R6yrXbdR2H7V1YHTTikCrVdI5Oaak4FfChVt5tlh0PtLGV/kFlh+xEYVAUELLoeT80Xv7y3NfCAT
m6hb1Q72B557Kv228t0uAYgIOxoj2yZz9jI/6p5DX44Q+BgTq2wbtSf2Sg16X1k3RrBYc+WIBnVd
u8hifYa9CIULxFcIrpfnBeuRCAi8Y95M3Qun1qn7D+uGATCccAAHdnTf5LWCfi9ccBVFphEIhFZW
Wgy60XaepmpwQ37vFf39i7A3/NedC90Tbzk9m287L10HBNw5BapeV8dCLj05QFVaLnF9hTkeQS7G
Wo7/zR/pPcxbdQWWES2xrd/rGSd+KpMAALcQHAj+gZtr0L2Z8d7vO/yPs/dK0peTjBSZMa4o9Fqa
/sPb+pLdUIVXP9riWrMOmHFYMtAelG5z4FzUzHpzs0EC7EaU0BCIAcr3p46Ci34w0nDxzgjHnY5t
3TPBhqEvqnqgKqDNE4y2ag5gvIhyJ4w5bFVqfxdxhb9RrBZEI2Yn6h3+bG/VH0tsTnH+VMDFHy47
ihxY9i73HLnGpPbDUQUuXetYkOvYVpiTyNKJGFjURZYPUkjNrSCT6/cEnGNUB76zqBDb84BCm4ji
kjKRefiP5qqljW8uFanAX7HovT5IY5UNCavMNXdvHz8WZwrrVSkdRAG/WyshkpcXRyEKTZQutpRp
c69ovH95PppWLCtjEsEzI1diyH2RE1qwNp/r5grK0y+/VGKPFv/BOQ22Da0fwxv2zLzPWobITBCi
6YakCYc7Y8Pvw5A7rGVO/+5Jl4cYmayO+Ob+wUIWXdav6uQY6DDrzkiOqIROAKPR21alioDG6Yli
OpFSXQLsy+l4XgeHVb7drj+EmsKMuX/vaBe3iXF4rQEE71aIBiLmIXZDx6fqcrx9L4DHNTTCPYnT
aTcEn1q27yHC4JK/VjBkWaxtluCfU1qfyv2r4QMkvNZImhYbvB3iIWHIGW2q4qBTpbos4RYF6man
CWlyZoO+nexpPzCq/ViTGRvU2lKQAxH/v6EZNbV8wS5je/xnG4zZWwT65AXraQp2mf7G6FJGam1/
eE8ogvg7i5v1n/BSZ6tGtg63TEVLT+X4xCpLUi6ZYbZNn4Lcd9ktYLAsQPH5xqUYgUQHIZ1zzvwI
cxclqpwt0bQ5xtUoG/17wGWXOvbtjlN4asq8xFikxIGzK7Xjf1+BXzfAc6DO005lugq/AYw8ea6t
HG85wBfdHjAXZGI1oKl5Rv3aPyjlqpN/D2nVeGNAF0eULY5Z9wEIHQ+iJMfZ8uE/Xq7xEeC41eGZ
f9qhz3dWDCn2dVM4Pg1c2GAYF1sbEGMVu6ZHc384Q6nUgW/ztwnR0P4IAV9uBvKYZaUA+NkpTY7x
GCfUo4jzGc5YPFbvHxaJBD9oIzkQMs4eMKNeaF4v/XGVXJdO7tZgSaqZhnzD/9a0dTfD4fyOKlFM
Aql7zrMlXEgkXGVFZmLOINt1b1lQ8zrlGih1I4Nr+FLULac0S4/QNgKxwkKqZwXh3xSjVO5ZAh+U
3BwJJ/15YWjfEJYRccWUHx1YjO4yhW3majUIacCzXY/VesiyZshyouvxaiyj93sF4rf/sgxJLPc5
wnkbhpGOyRq/6W+TPpqYCjwzsKIPYuShVpT8C90gA3H3bR/14glSf7IPBAe6XQvMB4eY7aed23ff
7E0ZVYDAWMCM8Vpok2dqxnmh0TnFehlFbftor2QSryvZTX8rvDcYimgR1skwU2WUmDEiz18IooqM
pVipfcUanoK2IXn9Mi2iPwmXPFVxm8FeAJeTBgIPP2qJHzklXA/HaLPYsn5m0FPwrCmn3p2lM3ZT
KT9pUtHb0KlSgE4wDH+nnmbP9kxyB+F1xuOgEkkA6zjs/6iGOsXIOSygcjSqx6LhOiADbqphtrj4
Evk54XWd6u+EftKonONk5uLXFZ1YJTewg4Ib2SjD9ORwjgu6wgUwtOKQghnZcLsgT3oAE2zAubK3
gPh8Y4VAr9J1EDhgbBuZlQH8nfNe/bffe6j0vILfzSlX4Pi966P8qFIh2urSWqn0I+TzNNSVfQj9
xQzKjxHF7uri9mc7qh/ww3fmgyU5wSy2fnLwI20WDsXVgYQ94P7ZSoBlKEYSxomQHbQS/rCQeAKp
uM+cMtZ72OUFO+E/0v/pR0xxhTU1yCvZXn1OaCP+Rko1ZFgTkingOU8P/FQ0hjNTovQ5L5XM5DIV
sgZlvdnoxbUBVR25rdh2b73x6suAA4vzz3JF8h8t2eswd9u/+rUQiPxcGU77dkNPTkGBKTRS/+os
fEheA3wCM3lfoiejBGF4Y1bWSYe8T6ai6cslvUBQi6um2H9hN1WW9sZWvv/cp4ezdCrtY/bl2WcH
0SrOI6UZdQkYUs1COEIeBRksBNyCqwG7mU0UwA+54MvQnIRDFA2GcLZ04YNlfpyfeSqHv2J9a9Qy
wKU5+aPng3NGntXNDmDZQWVrpE+2ZW+hAhYfX4GAIU2fLk85J52iIMM6C0ThFrh/W5i28tQIlQ5/
eJ/5kPIJeWNDagTN2T7Tv3XI2W7xucw3GG4klfxax+fUW1CTY50R9Dvfm+TkMUbEgHkkXB/J965H
UGKafT6nmKrCCTJyiJHY25MZU6cdWhCjBMRre4WxZI1vBQdSGWOmNfGT3ySGR8cvsSdK4q7605Qm
RLFiU7MLpD0SJEf6nK0wTM3Qji7FElyeo6JkT3C/2xOp0r/rKcntBOPWNWII3AFDDRrpOixe09fI
vTDH9i2sdmNwmrAbYJoy7PcNmtqqm0DCL05rPfptEXHQIuP/dLRzMlY16DJsABVQiZYKqJb2kYxk
VQ6zBJUUp/oWKvl6zPxrnxJYWfBgbFlEKv73Tmt2osdCCBwEinPLszPFXusOCbyTzrBJBCHTRSkY
VMKg54YrKwo2Jk+mR69oompea7elKsjPXzPR9KzIQZ3CyvU3Au2eHrgm+jv/nc5sH4rOwQ37ifF1
0JEymJxQvDTvehl8m1bFC7SGVPwVoumGH0ZfYgkJu4uZ4EhYd/WZ5VJ7c23EsjNDUcjarpFukAG/
0Im3FqXP7XN/K+K+bf4x2d0Z9LEqx11jxZZXIuo3tLGQPKGRKlm/ULhJtJAHTSvyqBgxt3cG6Y9i
LFghIyJdAK6RsKSL6IWMXp/sSV4f5Uhyok7IRqqhDQy4k0oKKaJFYyqVxLrtr9h3njQoKql8eGxY
3Rg/rrzrX12Sm7aysd3IbyXPGX0wKqaxVcjLJim3bSnl1Qpnm+jP6646DTd1uZpDyT6tALirNAmJ
7oct8IFPhNydeFKfTkWFvYKSaGa6fSBaDi/MTxuZzk3jYIE7gr+4ivTm8+l2RvxIQrcrb6Z8gbVP
ecn1psMgPR3/1HnLGBJHs0t8l/fq5e9NA+D7wlb8BjQCrrJOPHbhHZPGUyILNzr9sU+VZwU46Mvf
76O3OWnQqfHQfdanmtT1ZlSFtCSY0U5aAYKkMvUfnFdz0o/OpRXGWj5RRRCaluqvDDC9wZBbCHSt
n1G/AUdvZ5Eo8yd8nHH6F+alCcFjlCGiruxRC0qabiUmH6oXFXVsLuHSRCY/bcBtXw+UnfitNPi8
OriXQQxVzx5pM9hHUprL5E+Gw7X7E9R+8/W3NbxUXZ5d9DllD1KSfhUxkWpVx0JGiyURu47OAGDs
dibW35WAYtKTyNH7ToBt8KgHEFQEZ7N4hCr0njlSFxBTbvIilpCMOKuDs9veviTQGWuSuaovNAPz
N/3XmyfIiK/wepG4axCMzIaUYPkoflD3KqvYNK/OLPOrRvdJ6PoXErmo2ZX4jjdA3P6Pzg/z8k+3
1W8e0GgiZFpLJStoBdw8DJB3eU0BOK1nTX6jEnc2prbPuDenwrO3Q/iZbkng7zPvb7qbtLJJph7q
b+mW3i94rXoVSKZDjqL42yfw1qkYrQtc1F06+L0TTZ79ypDZI4DMRJyPouysdvh/Yp8BVLzORSeh
L8RLXiXpJDpBgm6KMp8Pd7Pt0FAxi70zNixs/A0DcEoTncUbHPP/J5VVusPoc/YKLlVDc2oNdbfP
4zc2fYXhkhZW0OoYw6dnTTQM3M6UIowsSdLsHH9mFv/GiNHaxj2SHvS26XyEDCFr63R8lZZOIOMO
4FeE0Enn+9S1hvXTjkij9JL1BWkYfqDOsExLjJynVQZEqecAVVjHuJwn3oSoCUoUU0tQkgoPRFW9
JDX+PxF69aNqUrRKVavsh6xmg5zARclhAEQu7+T0BZBUt9G09W722EsrTOvMrVxy0iMgjpWlXyQT
MkXsoc1ZfmbOFPwRAxCaEo8ca9cLJYGBEvmGkGBk7OFLRTp6/yfsBd7Wv0/FMxgYJoPJRMH6QVTs
QsUtx8b6IVkzIn/6Bbr6E1olZe6pN7Cp608cBWn5IBO8Qc7mJdUPmFQ2ZuVsUGD1kB22PPuKhuWU
9hYPW7GwG1Q+yVUzzsnRafq4D2Rgl9bgvsm5ULR3IUNhef3BJT7XMJx4rdCT3MFWw6lYoRqLEveN
oW61FTSdQfAYp505n1EsQvv7Yb+KPSADkTK02PeAe2zwa/jJc35RJAtkcZ3Fma6X8IoDyJJmLxSb
hYSLc6cQrqP5I6HL5pF2YmsEuz4q0tMPg58IeYmY3EGrcIdqiUCLaKeR6vGx7yQcXtBIuiLeDQfB
r/U82PLR7XAgeXMaBPwjd/N0InbJDsS4Plq2w2KqsXb31WXCZk+hs3s3mDn3eh0lbAkB9z7E6kjL
Q9+BlZh95N73e0jXwaguul9BaVeY1Rpej3GbDj5rYhsscVi0GGTxPqbB0+a0Y6e1FLZLiiHQScos
0ckv5POMem+hy0U6HXE9G6m7OhdVYpPlB7v05k522//IUsbsjbwO6uY6JroLdd17n7I6sELvkH0z
KoCcDux4jusfPHi7IeFm4/28EnFvQb8/dSGmbA5/cDc9ssqUZquS96nvx8uKJCSQp0SLzBp1ly4x
QS7K8u/cwvaq/W4cbyP36d5Sl73ZknN8xCrKTR7iJRqq+PwlZUZ3TzTL5udoSfC5uREaPmEcTXt3
m8mts1cscnyT5W5FAwbR+RSwbZU1X1wwkoly0m7/ZQi0J3s6KhggjRrdVhQB0lMoEB8YlSCtA/dV
CCmKaLNsvRBW+3u9M3kSGKcMElH4YKqVTiCRrKBJfL8PPq9MhvYB4i6nMtaSfSXL9c4PIjOvkpPQ
1jXg8bSFibhROddxhFh0pKs7xYS7HSA0QROTFirTi6UQNVHwn69Mvd+XNKymygIDLndhlW/Qf0JH
tmGUSncX/ia6LJZE7LpHa+w9f0yxudWDf4/r0uABrA+Aiimu/CCCGsk96rWw4K4xW8xhft1PyQA7
fyZTJo7xvO8BnVn10QgKsyKT08dvnVWxIp9TYCpqwgOXQTn8QEF+Maj6KLlkByXbqADpg6As4hbJ
GgiOSwk5g2fp98EvlheCui7kfu9/ZThFI+iv+k6JT+dZLK8RDtmxgTv6uX02T8q49MHcenttrV7f
U8b2aZ82Pp47xEouvj6S8NySXB4BxDaSs16dgA4yjxuRpsmeunKB5VBr2eNHY/bsaDnKAaVaurB3
nwzu8nXvxx+r+TOyWMRE7RifwOUlNZQmpUxF7R6OZEA1X9b5xm3LXj4IeSZWcxOv1gUMYOc7Nf56
ZecWHomCd8SQ3uo843JMvQzMDQm1JdnpnTLiN6E89q7cChS0KQovA8PamWSmd7BBY0YlrV85wOWj
fnYr2cRz/NckxbJqOAQWpnmGOPPojWMjkjYqfpO+GP1NSjmP7M8WpaAaXvBrHnBSKTq0m5UqN82Z
2UmAuLmLvW+kFimYraaDrLvWCsIlEv5VZvcvAYgWCIrIlEb1m6tkrjGMvAGw4h8nzmTSsnJu8Ioh
e7KtCJNDyHq64AnnUgnL/srvoyDYwZmryMD1TYwva5xSXCwNsWFSpgZV1FtPcEETA87tFn7YWnyy
Igd0o3inFtXvKPh1L3xgL4JgqzG9n1HLK+hfB4SUXb5CyYS1+yYFaomlzbIki4IT+o5wIvprPMzI
SHy7PXnL7bXbjKjsFAUfiOVA+N0GdInk9xowQBEeDEtqahQEbF2kfRmLVRRaWThWgEuGPsTcQc+E
anxOi3Yx9mnKkphRoydwPtpxiPw11uClo2D6S5Z9H2UAQJHinfPAwWu30KHkPuQQyHZW4AOGvq5L
13wd11h+fHJcQGHHDeWHRSbSDVFsmUKC3CJYa4/FhoNNHf9xZQo5RhAt2z7lWIQxJq9KKf53wGWC
udWpU90FxbfaGStAm4bO5Kt8Vc7CX+nTUIJ0EY3IEiFqlsZ7f2SXD4i0wxsLGvbpzoHiYU9DCQRZ
jnVX6RZZjTds/ZvXEV51lSrYJfq3zxcKKUghoZ2LtjSenjxBrKktTAGbG5ZvOKTZrVOjnvSt39Is
aFNFRwd3IJnnazBqsFGKYGNLAbANZf8+Y9bK36NdYNrrowpb33O622uR0iMEpIkiBZ03Gsf3yN2W
YEwFrRlusZcwt1Vnu6ehGEkLd0w9P0QUX0Yl1vfbsqHSDeIGE4U/WeKZfYb1udFcpe/7RhQk0h6V
2grXG7AJZiXhBKUdoDwzJfut8+XD6jlfBIRWXRSXeIrwaVg4saxwpM53XU4WMBM84ElUCaXza8Xw
D7LPnZvNF0+P4mm6rTM2xMge9MqjZN9Ay5qEAV200FP2H6BOK2r0RTYgLlH5yG7f0xJ8dD+qHVjJ
0ALKUqjQgeFyhoqbbd+am0rhsxNQ4vOF8sdrjMr1pyZfE1OERYYHsCq1+gX9vIQeX57DvT9NXBNx
mxsfpf3R2ClhVPznoNz8VI1FVQiCMlkqM15JwnJQ8FgAgr5qZaAgQslquh7Qi01fipnrDShKhSKr
kWmG1tYgKxu7fnkQqVuZbJ2usqBQeYsYwkFdQt7sXq173q1ka40LfUXJXkoJsxG2xZealQuTSehP
UI7KfkFVr3E9aSphrSkOgPIV94ZJ343WcZM2V50OIhaTsVct9g7kGUcO1VggJ/BIL0dMhkIgI8D7
UeBIfDGNPSubQptumAOLV8rWFFNUyJBAnqKNTOWTsNnKTAP3H2mC8od5dFeM3K3Pc7FbtgQw4y8w
BzlF2DUqKG+Nsal4/xSYiAalil1od356q1QmX/SCiZ+eectkaaV/za5x6PSpTtLcthEvWFmRlF6z
mNU0K3Y0WDSRATOf35A6dgwxgcA5vxKiyTRQg9sctQJneXecEz/WD3RBxy+u3J4fwliTvrCis/FW
Ej2I9MdxX0wY8GVQSpldB5KTfUArI2olhHx12BK0CoNtaPl5/AnRuQc/NHPtpHSw9Vj54XfcYctb
SVt7TpgZuCF/LGLvE1doemNzdmtJZeMah2UmehVSgpb0r3sye/0f++F3/q8ZixPdRGgMCWDLTdw8
gN6JMmAqWn8W51Gd01ytWwZlpr+v4nN1IA3jx/IAnT6oDl3KwndsGnEthou15QWPeR278HAxwq4Z
1D8id2zdaqYSEpKHVy5i795kRiWAmLeHJEig1PIR4/01D9iLKkB/RJq9jR3z1qNF6Fez7WDIhpKO
OEmjo+0s5YMHVYpqNfP3zlXGkiRZeK+VVXrFmMzi1ojGTUUBS9TFmLoO50cW0uv/mZssoB6wP0Xj
czhRXkrVE8/CVBiidHx+FjG98chiHvI8lREF+5dMbeVdAFudH+LxVvMR37pmz8N1AD319jCWyqiU
bfijSk2EC88Tw7SVfg0Zbwba1mTkIlUuQZNb1RFPTUtirWclaL0kY9GZSnlRP4y1md0PUyAm9TeO
FMe4GCjHwiSOVLT3cR/B2lUmasgY4/PjUBPHnmpHz/t6CD5TKnbf8LTqDAD7NHagVbPiSURW2Khr
W05jb0OaGwFWDJuLHQ2nooBMRO7xAYjzxAMX83LJF2730YFPr/d3T3WFH4jHgO9WJ14RFZRZaZde
MXn4WfLveRSsvpuHbzqRF+J81gwitlhPx8V8ZzkSuMX1Ax8oWjZxXsRWMAQlX+1CPBwwC38AXXZR
mCPetdpAb1s24htuQIBc4HT+7e84dt2s3AR/PUNIUnRGbDKAiRS3lffhrsAN4VTTebU727FukCh+
kyvFfsgv61YoRfRTKC/O0fIA/AkytzN0brr063bEbnZxvwfLCEO0jVNpXawhSvOy+mLU9GGz/X5M
0ejKGr4OQDfdQ2gEgA8XXgQLdNQYn1yFTAVjm3gUGWb4q0Qft5qWd746O/84Q+FOxYO0YrFssJk3
H42kzCvFGrGhwxPm06fHDKKAhN00Dt6ZDp1LpuwdjKdd0eeLgzexZ/GtHwl17YKQsKcl/XpkrEQ9
7aZQ9TAQ1GwQiNtdUuo40IdEZNET3BDVjmDRXJZvJyMNWYGEIZpdh1ssfZNGZXWrMAh3xtbgkyUF
XxQBoco5QRTpTgYvZRJU8/MRM8FTw53eJRhHfvNHpZsmACRhfKh88y2HmF1Fk2RYLOW6tuk15OVc
zvL98JM3tsk69kYfoEpyhcu4EJ6nW8GTXXTWdDwjLm9CUQWsZxVSLAg0TchGlLSjdi8TnYlS5JOO
4yPggKpX5gEnv0sYSljreTf7SdN7R/5TyIeAzkmlMvcNDX81PdiHVdsNdV/ZmEmSsjzuNBhDx1WD
biIRYuGLSwvcJChTPha8WIRO6DrwCmBlAsbKmLf6mILc4lxQ64xgGAZfB8qaGqE1cucWAnlWLbPe
TIkRVX/hv5o4PUpqpGsqT7e4SfBihNGYnFDxX2PxKFUI1NOyMuBaj36BDwyvGwOH0kJkhMdRejYJ
enqC/mn6M7xr7GX5snAFQgXbbF/I+6k3Tz/0jEPla1mPFJRdh0yjMj6UwKIuy7Jjm+8TX2cv+e8H
ZfGUSMumhDHbsTe06HG280QogTsi9v6a41OvnBhaxRUHNoMkQoeapq1gXQsWVYqgcxqXkbQZwald
LKJUSH9+dDXKaVuKtUZSDqvAHQ+mZ7u9i57VhzIhzs/6Tm02KFFl6h7MPpF81sx41UdIbN2cylUN
4FzTWSyC90+ZfIyaD6Lxubxl4LSjIjdSVck7nHPdNrPdy8mQ+Cezt0gBobVxcu5wUKekbR6VBFuZ
bfXVn5p7Kld10hKC+D6BWH3XGv5378XAyC8g5Vz9B4LK3/3Pilt5iUnnNHkYnVJcnI0LLtLB6Q9I
9aFivRQDk/XLl0X4dZ9YKY+lAvtbnHO7Mb4rRY5oQV+TnqCQq8TQtBfQ5zYSKM8O/qKGTwi/rlYe
H4jpDW4Cq7lSDuj2xwwbwxu/3oGNyAxAWGeaYfsNVOsft1hw4KDbQyRClmCeA7XTayKVRBB1f1RV
5nWUbjP+geURR4VWRvN0QRaFB4ycx41ohg6ug0CHSq6XwADNdAF4PCLeptYU8ofSPuIhVdiPDBmV
lLNpWDTdz+0MN81LgBm3G9H2fJ1+n6NyImywgFsgMgH90pwCAAOPsvhlnMRn0wl+32WKboASP9G2
v2vcG1SV6nZgm9A2cf1QHl9HKK7p8S/eXRhbZudTYuWY/GRy44dC7ZtyLnv55TTHFA/OUtEhtCHX
nC7VG67pWtIShKY19TM+wfBnLkwsTD2mshJRmmrKVUq8wlNqeNzGwD7EzaXqC56V/hy1aWIQPCio
RdnHWnSzb2Gy66u6WDKm9xVPfTy9ad32ZKEUXV+JDhJO8gBg8z+2NWdoPqrM4ELibcQyLplzPQ2l
wKmHFaRZJgsWkYDhpK3povQrxyVb8LqmoGzEt5eUKcd6GoXj+AfuaiCdWO/S4+6OPOveSGPdmoev
dSyOssAmtxaHnsvhPN/a7Fhn1jjXTCNHDKrnz6Dzr85qERyldVV+XfGdvxJFmB7CHYh+BLU6m2hs
sDcAAadOpni1H3MWIg6tuY5lBEk1GGegrIqi7GL30qawzIPWuA91tkdq86T0Jo4P7b0RQvIrCvpQ
AVp9LqyjW5RLbhx3aHI1jKK6Vqu64icAE1tbH0gx49QscpwZNzOEDE73+m+4WkQq/EeFgpgKk+0y
hXAUQcC7i8x10PWtILQi4XJ54m7iSmNY6nrmZMYSN07Lq5in9PR+0DYhN4BcMhTncyJ1+tigfycL
ZV7fXYCfJYZ6tW4bx5CEbBMf65CkHiJq8H40bNR6h+BuCVN4OCiemPRwfiAH/TDSm0OjS1wTsZ/T
75P4sgdHO58uCV9ZJrcpIqSNl//AAQNxFbISAwXeo5I4+cBk9l/L3WFBRJTDmb/MFV+EpZXK8S0f
rVVZ82XN3ls+WLJ2zzujtLZNH6++lIntc8s80jDp/0vmytS+AoJW5Ftu+RZBftduczwXgZS50CXV
V8q2LpauAg/cUPo6q6ZmiJ5BoPmUcYIInEyoQ1Z8J8QHz7CdUQAZmeEVnN03uIz1WwyFAtjNRFuM
p/Yhpj39NJN/3uCK8GZOKO4LsuB6SnYS6Oompb3Q3QiCRVNfRjJeg9jb9fy3nWVJduzzBNnFiT+e
05mVK6Oqxsc+cxgjya201agcn4sIozOdwKn0vYNsk0lYKL+gz7NEsxKbZ2dETO64vsbr/bkaxzV5
ooCAm/WTS7qr4LiHDjul/CGHKAXy9OpYohE5us9X63NfKC8eLDIq7dnsDFMtmbJlD3lwmVhnTMMo
5VfuHa30DtKS9756nlzLIqeiWmluoCC4NdoacEt0AJUnoqXYXZmpDw1+D9lwwB+PtAp7QxEGZnfc
pxsoKJ4VeGoSYD91rRt7Di2CZC3rDkoTDwhUNr9+kVHB3Xv4StzUNBrp3BS7g2tfX3oxsNilUFTI
uipZI2pXvCk5assHXTpQYhbAgAp2mhQvGWmrCbmwghrLUAbtIbBExrRboOwh2mCWBgTCJqyCDkY4
hm4J1i76Je/OkIqySZCGLPYtbc+tHut8OfE/kG1fs+x8MT8FXN5o+R53WGlpqfTXYFAt15GGtUh8
drFUP43UKuIGl5fdllEZgNTWDpzk9rYEUaPRovErtKzqrl/Is3oi19A7darGGGQ3MBAEl4qWz1ZR
7sKC6MRwbEwjKKcbkUwRzT7nRyl3saHYCWLh9IY54A35RzDr8AuUKI5Z7279S4+jk7Eube6sP8wG
/jiMgNozjB84/eQ+Gd/Iu8pANeDABQBENDH74V7eA75AJyWr/eRt7k8nBsYWpJxrUhXGvP9Cg3by
aDjt4cCNRkJ8AWOCZ4flHe6BsU4FNMnM+n8JvOUqKJqOe2bwWB5xFG6qf+Cjk7tGmoHUg8ZRl2bt
POpqLVqduoxdsvaDg7E98eEpE+Pgz6swqNZ7OnsyJKsaH3u09jG+lbq+hc+E6CUTmfBrkz+r4TPK
byefnOEN13n02fTa7eoMQdOacoENu7CRSi1ApKjCYyxCL0euwDT4iOlW0UNpP4HgQjeJvifwtajv
bHpSP9BQuvkCQJvMUD0ewUiKJvlCqDg0z0asOqBAF+T611Auwn7P8jXE9xcxpkxaow/cZRKUm0GN
gOEXLmHS6Q913tfL1O+WEL6bC14Hbl+BPcuZuoYq9v70QSYrybZ6nMlLf2g1Z6BBVjlxVdAx6HF/
vLoFPWSyeW5XifI6Tgyqe8nnus1cgA9jrRRwrt2XCAfbXfWmmqe5rSFXE5DVh5sp1CDFldOxlGal
4dfE/0bCF4b8z5ER2nXmqifM6YO9VEiMoqvzHRSqKcndxwHPTntVcM4XJNBggQ23SnzwdG6wTd8u
sQCSYuHY73pXM6SNrG23yqi1QdHYU8dPa2KbGsdfXqE0wjjLjBvk67WaNEAqpKCi0ft0eOKVGcmr
PHSUjpvEdDnl6k66WtAwMiqlzGcUno1NeMo0KIS7Tlu6w3Xnoq1ONHL7OXQnXnWiQxIkU1WVnwZn
iZSfLKiuafirE8tbg9mzCSmCRXnyftttmrR5P49ilHXMpMjuV9NroNCqB/xQLq6I/UgWX+JLz9Fw
O33iICYCIN+7AOJ2V9GoD4WkQuMgfgy24cWaosiQX1NjkylHGCfmZ0WEtPI0uNtW1/Qq3jmcCUSl
6mnuffCbFdddpk1hcGFY6BgiFrkt1RARXffWz00L5gdXWu+kJ3020ytPToDaFdmZQUHkQnQfRoZz
KQspouWlc94HuQyK4PpoA2I7zZPbZ17JJOrNZWVTq92z91Rk0pB+fwxJ5bte2nkJIySy5iNRhAv5
NwBINsF+4W0MDuH6Ce1ULOWEXQfBo/MjCPaBsgcWRB+wlaKjJ9a3/OxHlM8MXhdxRU9qXL1uqYTF
Bq5IHW1B/rF8FAZTmuj1xRfFKcTZdt8qqFWvW01kIjqvYb0jOkaSWSlbeyNI711XB8z8CYbaEw2V
HSUwXmJYAyM0ETQB5V1w1ARz9p/w9zMmZDuR8PZZTb1hdvLRKzeFnVTLFQw9vUC7rjCZB0EvAqc8
Jd3yeTV0qd1TO85hAssJYlqrdqJ9xH1uo7IlnAm0yTrIjhNMu6WbVSAIG8M8u6wFVElWWR2bFkWQ
KVwRPlya7hWq/Ok9E0YztrTJ5QLZGjpjDdVPSqTe6+rkFcqftqHfvglqDtrqA7SD7BnkkT2xMf4m
CaRW9NCb9S3MSEazbgAFJDQ8dAg42nq6uqY0lTFvjN8SsX5fHUXXZqAuWCk3gWoyT/WLAeJCB3BM
9+QD8qp4ys9GKrTslWARKCGBoxjku/CZUjGquyDNQGlhDikgmUlqHPNjJ5sA3ygD4QSVaMzmeuEZ
m0OLLy1q5E93ftmiX7GrtD6apwKXHZ+mBy64KAUVWHS6erQOAUTgckHjCehMhkw4KjJDA5A7wMhG
4lGoD+tA3a/1uw41QabjGBsGznAr7OloN71G9ukkwT7PL4lFi9M9P1HOYOAFgUqYW0j0xTkin5IG
Qvfkh+GunFLTYqbyJnswdWkchLvvdn0FZgpmomt98OfydUbAB7ZDwxkumUiR/XuEgb3PC3jCjiGw
JPLzqlfMG7E7RL8ZP6L8eKDyVjTyqZy2qxIjt6ImJIedB+4o4sZEom9w3f+rALYPx9U6NasLaYt5
hT8nVJ6EUnImnhUzJvVyKcA/0MPKL1KM5xGaGGPoL/OpgJAtQAzTb/1BudYznMP4yoeio0TdFVmn
nkDAgWwCR4xfiBCDvb8Zl6jC+NDYK6NdvW+g9xknYvJYZMBd/qnTwhp3a7f5x+GVpCMLa+xOzBQB
tqTDD8UeymS+LCHc1uXeEDGSocS2/7QGnr45aiw0jNApOT7i0xuJLdLjBWiKPLhpkmfJXq7vA+PQ
qnNqATvd/8xjn6rAy3zvO620+4QVU42VncX73N0KC8nZzQ0oLobx9q61bLdnXcUqP+ciiq0V6PS4
YyNCpTPE43hrELAhsZoeU9NE5DHZ2Db9maqXpYDcfAtfmOl73blYh16ho3cm1CiWMieBN2fvuOHG
A++bPcfoag3tm/6dqsbsDVLN+MULxWEOTKU+98wmRPiWm3TAn+U9ydn6UB1+kKVOacVYjnRyGyub
0OT7E1j99uXG1F55tKpl+Pd4mAs5oNgCd2hKZ4GdiBMwEPja0bKhq1Ufwyx9D9iMfh5/2H/v+h4d
cGylJCeTshRXlv1/dtVZbi/iCGs4bvlghGn0Hy0FvOkuFExMV9Fy9QdPRPl4NDhLgRni5NF3Ppoq
lPLk49ouO0w6hoK+aY5AMGAiwFQBmDQ0Oh2PtqW1q/h0vDRa+izHMgQUM/vDBZ4uvmdpvG7WSD6O
2+Tp6Jk9ns+b7vyiy770EyLOKRGH8QEZ9yaZ922Kwez8r1wQUjpw1omYT1laAwWzfQnmv/3SCnMO
vvCZ+zWkVilvMGRqa+fS9OvjQ2oTcyM7Wk6dB6bH8HS2pZBXgsrAvbVR5sKJF6NbmiDbNF7M+kLf
nbgmZSghW/0GS4zWAJHo+qpl9AUM48aTWyskkiuq4DG3rSNNRIhv2JK1D3J7Mihf36opHBGxR5hA
la2OdMJkLF6cHeKT7CTPPshoJecz2pdtXlRb0mGpojgAs+CJzHo/7o5pQE8109lmgyYSlBz6wXSG
0EnpPOM9mNYL4THy0KlE8xEncn61ORaQQewamhxUp3GdksTc1tVqd6U2jzaQxRk6U+H9QONS7kkO
s8ydIQQTIMjWQ8apktEUt2l9yS2AI8PEmR/6LVwDsbPox3pM5xSjHK29vA/CnJSNOwkdm0YAk9Cn
upZH8lveOXCm2LzibzveI3XODigSWP6+UiYQrx6w9wOcH8pNmcM9nFRBwcjhRaAfSJworSUWCKEr
lLwA//0QYJihI3PsXR1sS5Hs7DO2fDbNoCKyA+XCGKCs7aqvsbDoPzPTZCyAjyz550c2/Bf2ff2X
bNz+RA2cY20QjZTMYy1/n0J9MIZ4rKJCe9NmQGSBxbaQnGAjbyVkfLbOPfaYB0hT4uPXkWDWXsU4
zgMsf2NCR2LuMoOuK+X7cXHtps6pEXNrb8YLIJj5VjOgc/18G8a8qN2KXuCLmWeIA842f21YeODR
X4opYBv+8xUfrITY8L/1qjppFzZFi7ZfvC26T4duqZpVK7fqdI+jcu7AmmmEgNTFWM1XVRNLm0v0
tKL3+YyjKY++v6hCRSpOGauUqwKJPh5ffiGuLgvO0GbIOJfVjrtnSpYICYfsU/kjalghRENvQXho
yczicMJF2NBYq/YwmozP3PcyWVv1AA3IsoZ77HECx7q0FFVxwxokF3Z4uuVoh41ESGIBx9RegD7s
8VzuUDj6LsufN56isBeeM1bIX0msamfx+F95XQ0/5ayUTo98Iw6cLFAq+cRd4WdVWuC8jwHIjVA2
XEdbQt09VqSBgSEmh8McVw0y4G41T6ua8YdR88TZ01X7Zj3ZXQVopb2/6fCrDSXxyNOodO7TCQIE
T3QpRIjSGJBwRldouM51W5l+Dp7ZOqRTjsbxBYZd5ULy4m4eJj0pU41vmpQLGGKnoBXGogth5ssh
QAE8Hga+fH6nkPSrpNLAz5PMafXKgBswyY0kEertHhMUfYAgUup8GXE7Q6Cu05J3JjCecym+SZYl
nDIr8xIeCJ9GG0P30iaXCOu45QcnugWO4z2OUfqIJPVz5f9YvsKashCjfvBPGOxYTd5xuox4/eJQ
92/+8NxDQFORfb+G770DYQ8ypyzdVtJ/OWMIwgwNjVmXP+mp6fItN50zJHFUbHwS7jMi7B5mAcC/
JEzbD8edNqOioG5QdPVG1BqyIsR+AWYP1PCp6rYIMwN/FOCaxzWIWBg35ZOGe5RR84L8XqlCDsyX
3sAT3KMMo3Ss7bgnkqprQZwbZZF+h2nspEChvBbyBC+0Tzp9+TzAxpMeQIv2aOK+PnAQlfzab+jB
xgdao5ElQuK5GeoySytiW7mpL8napL7pjypUncOBeguhIx0FOQLZnsXBPBWN3W80HJO6nqhEtD/V
BitG8qR+kuc5UqVvgo5A14OzLuzlkEZ8P2SlIpRQImB4AvXp283wLrmqHyaEAjrF6Pob/6LbI4Pw
DMcPndM3IaGUzmiGo+YMlxIPy9M/2CeERsz1HOMg2KeZUZ3E5t681tOtXPPPdU/5Xz9LuHcNkTYO
0Ai7KRonMwpvLiv/0JSSviyaKIDLTxBB25Fy/OzqB5gxlNP/iHq93dnWKlPsZv+oxzH783ctXrfr
5LYsD5eLn4EpEqMgeWrHO9JqPnIA3tQTn2czPlpbHPfFOO//q4gB7fEw6e+kz4N2um+73/zMKLKg
IpcycgdJS9k1BvwtW1Zmboq0wd3sMCrDe/MCO8FP+QNgYMFaXprlrL4PVSyVw33DFHTzZGtDIw33
xWgob/HqLu0/ic/Mzz0p9TL/9r+vhjYc5kl/Gnng9RNzGi7W3VNrUQT3TgZ3wxq9ZlDz/UxF7ToY
Psh2xzJSYxQmh1KgDWQQeR10xRAr7Y7KWGkaqDulPy/Wg5eUDz7jC8UbR4D0b1DJcEJ/veNEPfa6
QNoF0/kFdPJZtjE+6saLSD+PmZyJ3rmZxWIVAd9tBL6RgJRd3fslXtWZlSJNe6Oah5AjyFHeWtBU
zjaLdYg18anDXwty5ntyBmPLK13/2wG2SCaK6VzQSZNrtoHzfWx8D6vARe8+kdgLN14IBwMynrsy
jJ/wi28rzKuukyNCTHfzo/G5drTAfRqtSqyBpzQi9hYNTQu+4WeQoBWC0quAizJOEopd+kKpmvyo
g3H9SEuQPCC1vvd0ADOjDeXXHgfWUHUC5YBuDEAJ6kx9Txhrwc15PyQaFWQE4qTLUgAfESYHeo0w
8yIEgwZJJnb72slBEE5mSWNZvK2d1D6a1cSVd/o8NjgNGCpp+fqd7AXY8eAdFomeCUz0YEbEGlPg
lQC3ic5FoCvmzKKsQn9fUkgxmYlvIGaVEPz4N6LIikFlZREgMNIW4kpz83M7tMNxyRnAkut3V8sq
pnkB5tugW0e36uPxMlxnpOikYFZfx9tjpfowoVrUDPrZ9n2fFPxPmNC2j7l0ouDghoL252o2j2Z5
PEef0iTmWU5kV/hEtS3vn4pv3RITGVjZpWgTFvZ7QXzCnZl2XZiioLB1pMmKAJmDenHc8Z3NQ3MD
4g70/Mm1hm1ZqJWNh9ZRidkGL78u0hCwwVsgDEBaISJHLXzETcQQthSIcO34alLBhtNHF2dDJt+Y
kRYxcpUF1Js2IP4K6Eeu66S/IbeZTUYEAawg+idDnMm40vSa25gsswRcA4u47C+RiRxphwVwmZKZ
GKSg3M0ADWPQXSSQi8+8j4j0dc/3MWZV2jbYBOGVXYQCQr0cZw0pqVYAuwu6uJP+a9m0ULE8JE/X
rh2HGUVRtvTYKQW1dRYgsBt6CN6X+/+bowQYgSEkQqt0yvIk/Kajh5zvW2o3i7CtTVOGit6t3Q11
ELmFsMDRzLdxxT3o1FiOza86ozB57HI8xT3780yWznudLPb24fcXlzRMXMsdQzpoaVUYevqQfqXl
ivd0y5UgHBits/3f8H5sav/JLx7VqJd4LvUPILv0ttU0HQFHwhpE2t9W5pzwQML5DdRSrdQni0Iw
Ow2YZuuVUAX8kpkRo0PWJnsJuvW9guKbgZCyOY2gGzETKmxxTIE9O9xgEE7qJzS7Il2jKpH0VKf6
NQhZ2qKnlO1j8F5C2WdtEh6AU0FBMQxiTedtpifa4O9hiy43rqGPyuFvhmT9+i1hisfGpsendWYa
vBdDaqIgydTVVFaKVXDe51uPIv5F00j+osEzTIsEW1JW/2+ikavk2h2VBCgd+X0KP1jp6ZxhFfZP
Mfj51hZcMPZ1xREMo6bC4FFAnLFnWNMSga0OPQXKRcL8vCUwflfDeJN1n0zW0/kR3gyCEDwD5z4a
m0vSBA7iELvkyf09YCTAhDbLng9rPa5fTlAk8H9MWTzIFNGtBIGAsXHqZAgGTViEbsZwUCg45gfp
SrGul+T0eIUvWzcFc2ddOBf9YdRMJ99Vd70nlwsjM1dEh1D8eHI/PXY4RWLjCDHsmKqY38DD6g7V
bchF4bv8GAmaf4QjFq8RMJX2teFBmQFPPghcMQh4Un0YgdSVkEnS+skE8Kf309EArAdmbmMYwHs+
47c0wyF0RwrEteQlYt7TMxVJPetUUlcBT952AUcdH9yF0ZgIhlXNaP05NmQzqwP4liLIjwU5hUp4
TzTNFdBZfoc/aWK7mn3nIBe0s+OHocFkD54Hi5jX8XMStxHvms7LVJT7zZ2FNWfh15bZR4LWKw07
ykfweILaWNTWN+VvsGNvlpb1yv4uD1EUGkX/r9OeSc9uy6FoPlcKxTMO9jFYCoCxhItSXIMRtgmi
Hk4iEUwzYTUsPEvyetVkZcJe1erLQ+Hq2otgtHEGPguCjGpGMezfirNbm6dbk2iUTUwBSF7GPQEQ
uU3CNQg+I4q7TAscgnzXWo0W8jer00+THWcbqin9m4ftNkrCh45aPo5Oolxx/0XvY8nbMgUlFkrZ
DnLKydh8TF9ujipQecsfLRe2zoLEG9DL+Lhi4qRkeaFpwqQt8H2Uahebc+55fy6tHjiM0l74cT+4
5qk0nT6aaNzGW9qpmTxJn5Vfom+GaQ6P8xHynutGJdmm6VNXZs2/mxTnYMBnp7dRFYW7vZZJ6pdO
n7i6w1sPRgyfhcvpm98vtYVk7P0XLWt25Wv0QfRPw9xo7M/WKm7hVPfGvuCh61htO/zG+x6irChu
YWiMpkmsQPoJGXusGYjhtIxGPy/fkX1E6+bUL0I530XN6NYGS0SqIh/VgU80fzpeEHjuiClkaMHG
Q4AFAjlu5U/akMfu3GL8OJrxtgFnyzgBm0nBoCqVvGjKyswupxO/g/SFBXgT23Kym8i65T/ymSEX
KpgznZ0YHM38cNtPhusGCIV3OithF+SaT1U5ZSMopyjliDG35MISuz3ZsqpV1AG6m47a4G5XYekD
R5fTEeKvNDB3SFB2CoW1ySI0RWZ/6LmzOuK0x0UkfnkLUGr+1csQS6dIL+mJO9+q2CKOqVvzZjjU
PBUst4ktaAgH12NcKcgFpoNZxzbzdRXKdRpT2VRLG/+xR2ZkwA0uxiTXHCoo7iMjYbpqG7TDwbA4
ErPISoxFQ4VMsyzcnxPodSJChHTGprCKXeFH4+z+cxbU+JoTCF0UDtHWpQGbJLF6DFCG1gCVfKvW
cwKKlo5/NjkvE0tAHpoqLvLBOV92LHYU9PWWC5QwHlULAxlSYR3sk0YwxtlJXMauIu0FkWibMcjg
8p0uv9SsSgxjmlU9BdDFAwjyNJ8zDKwudnbQr6r0OIqs9WP8BYxGn6KQ3VRfeuZb0NrBBLyLQrOS
+2zKRBpktW5yNPKZe6Cw+gEftsieJm8ZiD5+249VlKnH0j8ib+ueWuoHuHFVJd9ob8hVMBnVA8ne
aL9bCuxq6qyARrCCFyfTGXaNGFq01s8G81iWomBYv0YgAw+saBAoHun4e5PYEcTVoH4IPI5NbYyT
ndY5uQK+6k422p3+EQ4mdYiBBwhsMOMAiG2TMmzgZu1zaY+pXX+y3Lesn0qaGbSB47OD10rTmu1L
dWZ05kCkeeaStA2uyCIomn+HS5/TkGMGAbo5y0CTtk/SkF9EJWHswW8xlukJ8iIrX+E9sTeTZjX4
uyayRl/yru5a8SAFkddsuUzEc4A5h4ZD+vliV9bDOHwTrUuleK2Nx5JzAouwX7P9TbSzONTBwxnH
JL4dpnaV7J1czbg1ZC2za/+8vYuoC5HTLwQDgxs0IML+AGtc6g5ttuEpN7dNvypEkhw+vLjcTLlf
1Zp2LCF7gUNWJc9XgTbhaVu+zIsTC+PhLA5Awbgja6LMcSYGOLAEUlBXNTng+lT0g5EOi4xCknld
HwV2C38sDbFlPUh4spFNlZp5UX1j5kixaFTSvNc7G0UAjkC8moaReOjSWm9Na3KbvD0NjJphRznp
ZH9hpPICj2xXzwfMi9iHqX7K7TMq43JbmnrJ8O0HmcM6vXd1Ui8jc3gSAJy1rs4Q9pih4I4cTrb+
v7IzmlxRGqG68lvvmMmy0vDsrOvINU3soVtlllpG8M1f272DAfb1GyXMDqeBYc/8Pb5bau7Zei5m
YzENaYlp09P4BlBl6fYxp6Fl4qhly+f12fBxZCyhx2KRxMD6s5o+yIN/6fpQgT2InRsaa5wEg4+e
xlxM9hzKQYSyyHgjt9rpQJFaeHfRSXMJATlK9nRK596N8IrsrD94TM5S8s7wMQ8NKo5QF2Md7Rt2
VTcoHvQbYeftcDo5eMUnKw/4ALsaIZhwczxRnWqbTWeBE/aVy4V+kF6sw5cc/CBPZcaSXoIXclQv
B+yxP3XK2lS72SqwCpdui3RpC7DCJuLNTvuSMR9DQTazq8vTQ9o0mEYdmWynruKHg8t4dDqXO7r4
mb9G9HFJ4Qhg361Gy4VHQs/3z1hCfhwxwQ8aD61bHqT/un9je8NaOWVq9HJKdEzscss+s9JfUCM0
m5BwJWqABsSe+cEp9IYGKdKyWG0JeBmfq5T7swPXWU3bihd9meAB/O+ydY4ObkKr4Nfh2Yc81TNC
6HJ0imzQeHM7WrChRHRDpQTrSCYG+8IsR6RFA3/m+9FAJejqpHVVvHbYg1zp8YOSQvYi1OKJbkyj
1Qwb9xkPWppJgX49XJvbE6BrEy7qYjgQvtb6J4Jhw7TRk8wpaGhkjW7s+9ymQfb/Sd1dnz4K+Dv4
IfqbFP0sNSGojk4ZAqlYEMURMxGD5kSVEnkjxYvBfnab36Ly2JmNP12F0mIvEfdNyW2xtQHhkyJR
AmYrluznwmveJ5kc29teJ5y59UMNZyolyYzMy4wmyh2TLn4QxhVgKZ841iYUADgECe3jah/DvMgy
ENOEpnGD7VS2Gq4pZtmQz8MX9NRx88nXKV8T5YiRhF5WI1qVd0Yk++GWD4CWHijxlddIZOjv19XB
dN9VWlABmewoRtLBmzOrCERQ01BsPifXFsrPOydgAjb4XZ8mOZpXlmgwj1RHOwrrKXPIeGr+XtrD
+8UaOyUfJ19Z3SrHVplVvwZcsnuAIhOefp/OSy1B1NUMcKjSmmvSy0KrNoLjoKc6ti3pH/Oo3GNk
su4VpBemcEOYWjhhaKBOFstvDkNL5fi4IPRlaWyrYIacNy/Ez8f+5rEhaL4ESWdYjT4aBJvWYFIK
+sOBI44UcUGiKT0fujHGlkCqBOeYybEBMFFQwmO73ZhYnizTtwd3eWrm7lNMwhYI4MsqS6Ub9Cpl
aW+f7ucQweW2yX2HxpFy6aasDsTIcGNHbL3KKT0hmHJg/6kH2ik/yLSdX3w+vll8Zhbu35NnYWAa
2pd+E/PymLcI0NLyHcZlgbNs5RnEiisX9uHw/FCdXmPpC/RTUNeJDa0ta66SJkpUY4O1uTPRb5GW
24EzPKe4zOfC6NxfCdxFuQPI5usCqj/1vBhhQXnWoSGYp2mC8hUxIMav+ls8G/8o7luAk2IfjzRa
eh/GXz62+qptnN0iekorRLxVali4mX0HToPg5y35gyY7HtZlOmnnnuZql0SZenHpqG3U16M4bGwi
JRSlIxpPJ+nfk+znC0HvaMtyQGvyJHslcUY2qevEICeJmFpSKF9yX24RYsq6PdZwtLPjeIhDjQfJ
0Xc41NL/ApUblg6Mu72QOOi4flwYjY/xuTHeY7H+JthiUgXI//07+8PeI0f4/wbVi53IZkgbiOQF
X4xPnfVQp1TpicS9ZDBY8g20PPfO3gKf1+B51uPtRNTUW8QEfRhgIC5dGzOeXWoJhJIUhPOf0G4Y
yAySGicAgcsYECXWwUvVhuRMP7vHEvXpQ59wK9IBM1DSBzjGQVHtAKKccrdrnrruDNJZQZF8Yi9t
4HE/lhTPnblFeRp0nxwDBciK/C11VLxNnVRqJs1npYkrJrLIsE+j/In80p8AdywJL2CwPVNXDtUF
G9sIRTe4dSUDNQyVFhufr+tbTjrhL4bj2h3UkJAn4KpUuRMAGEjTyg3zOl3yd0l7IdbNd7e/zXY9
Qx11xt+IRaQ7gw91bZsmMDLqxpxtcn1rjCXO1vq9h2bZbERY5sz6vbSLCEe6IpUGFGxIyluzxb8y
RXXSY4zMcZ5D2a/Tx0CNgSfpT9Got72OC7/Zr1LkcaUcx0boApfQA8nUOVKlRwLC0R2n8fXIFusy
oNVi1qnmid+Dq1fweNVh9T5j6b+FAeCcSS6ZcaIFzivlvatFSjplkt4+vzzUF/Xb6ieMZwZsJC2Q
uaGt/7fYtVQm7bjqV5QV5BznPBDo+kJcbQyYwkvTPoFjstt2sSqZqXGmu6GPS1MynVdyZYKJyiAV
TL6IWY+sONlgIrlAcLHzbGMoSgMh5d4Bn6DhYsIqo13Radv7C1XICjfPO/FyAmqzWR715ute8PJ+
rjJLX/BWMIV5CtXJMHyDMimjKuKWzTtyNCfAQsKlA67P5p0n8tarLgTEL2j6mE9IU1K0Mefeb7qJ
JUAb2KePIBGPZGLTgwC8IjGtp/SrWq5s7GYQ+Xd4Q/gTghUeWDBv2Ldo8u01FiZ3cJuKZZxa0d+A
hnbgwQ02U3zj6k74a/mYnJV7Vmuhp6s97tHo1flYeorNOENpJfAW8+V2RtJ4iJvaudEyLys9H4B5
IZPa/jC1qE0A5heW0a9uT4HC+9C6eOpWZa3ihTxqis5Sw+6HLdLyCwZ2f9zVpuFs4mfdtmwC32gc
uaS/cLJJLAvyvs0TMioeI/VEoOteO22uwBgvbkT3vTgdhqPoFgnNz3IL28UtL6rABiA4EzwN16PU
oTGOIO0Z3vLt4xB4c/rCd3CidnKgIB29K6pVu8ooHDxF60mL7HdobonJrhH/6q/JdjoU5nXKjH5E
L9xgkaE3954gykHr4mrfhuNpCGMbE4gG1BsDGAG80HKKmRxdZYmrzukR5bDSvSJyJ+nAI+UBpVt0
Zu/HO02Wg9rLy14EJrfx3lWgvWxLP+M+jVFDt5kFZSTr5yRRssL5wE/2aIdU+obxTNhvQT+zGw4d
3H0sbS10lCBrU0IHL73TluW5YukvBLKY9vxsrSHlGMgyHX3dI8q/e6WAvMS9bVOV8mOThXl2zE/q
cAXi4T35LL7lwyduUMGcXddiCNaULWL7x2bW6qMV9kWuS2G9I9J4qJr5oKeNSA8TrW7w1/wBADJ4
8QRUnh8ySgkW5HTxunQ/CV1fb+s+pwHpkrbokhX6c3M+P8zBD0eA1dCavymbyucEs9P0NP1//kZp
MnV1Ua2eD5jxmiObzj+EoeYdJ9uek0BpG54Ww4z4JI25XIXgYTbLgOy87jF0PH9pV8DWakCHFjEf
eZJDajg/lxBazNCh41lhjUTW3DRyJyfkD4wJ5CAN92GXF4wZnGblcEBlXV3cuxVjn6sRnnwN1KzC
zhhMCydgiEAlNQozxlWsddwwyQTTVIaNoibVZb9+zg3jPDumzaYMFiKdKkBKxP1222ltznWG9cYS
5IEjHyCeo5i9fawi5u9utVDR3LbCy9ZJL7lZP7dB6wHiBDuwGu+37cSsd7m+ylDd6rM+sI5yt4ad
P7Hqiyjtj5jM8wvJrczwq73Kt6riXAOTELaSJ59dZs5OlcZsYbwl6QIsI68x7BZH2rBHKxGvS0Ty
jRpET+Fc5r2TKmdrYhV3P7ZLq0vx59WP8YjIoRtLwgJ+61vjoDChocNrftA4G47tfe55lgJZX/jT
5hu5eYSdwwwoPSeAbxGlZrVsTClR6pJrqphfIrp1DDmnbbNOPrvus+q3zw/yf4SODN89mAZdPMqn
jXAhKC/glEF2v1SfEsB4TK1f35uLeQka8lsqM36o0p9vXDcTyiCs65oHVuhwxfRkz4d3vcWCCAEB
kPHSDQvil4SB4Fct7hhXTOmj3+FDz0Fx1Ks1qMZISr3Q1evqfJqRGO8zUgdepgEV7Hyt/FLFXpfr
omI/+ise4suMauVoDyPw7lMiD3ntoYyzSybDQLlJOv1tvDuZ/MqZ2KIByFsXOHuIVFwOrWfeCACy
ACR8C/v4z8FbsGE2aZc30xogshU9+ch64usixrDTMCqhBz4P7Jzd/F1k20nTrSkX3CQGtoc9V/vm
dzkhYgtPntv+BbO0Cfdq8rDgMHcE3aA41qWRJ3mvBIOelzjeY6LhPcNMM9M50qE5HKsK/r33ILG/
RyTLVTJZ4u25rgdYhJkuz2aO/w4b99FVJ4oD5lfCrtM++BYBVgyNnB0WN7dbnFj3JS99CbY5EvGh
N0cezujATpMNRXb9T35G26Q5b9D8fEQEZUeqHqOrOOxQL6gwUYIGv92QuqlV8170amQ6yjcGoEJn
IDXLMBHcf6vikdMg68P0i5bn1Og5qlr9G+kQIGusPVccT+Itt8atWGFfZkO5Kib0Vi51ZA+AMbTs
+1Z4MlFQQPFrepIinuBJODvEGsvLOOuUaWe3XJCdaYxtRej7k6XMaRaZPQ/jKmYVZcli8WojH9nm
+N1g09zjdVs/w6qlsQ0N6oet1/9JvC0it94/fGqxOvFurLP5v2VA+kN6HmfpWLjFAFF5DtAk0491
SXO/b/6immo4O3SPmFuDXJG2cXftHWhPziEpBg02wmO7qSySfBvmZarevXN4f+z4KL7WPXiXx/hp
eXERSqleDYLzCQS/Bj9soo6FT4uuzmPkbMHmMD9VafPPKxSo63v7/zfNLoravEr7KecGla7H+cDy
4i6VFfJ6fAe0VVwx0wwLbHyx0J1x2z3ycZv7J/o4NP/RcBYqdmBq2ryogi8OUvNdYdk3LCaGhiM8
Ivg+XLH93KwvM14et+L9QHrcm1y9DqnkNa9epgZPbBBKdXl+RFrl1gIQqERCtf1OkpLCO7B+mNq4
1YT+bOTHYVFoCXtD7TBH0O+88sOkyfelOmjvryFTSNLUst8iqBHI8kichcTqSAh7eLeawHYAXmHs
icVQMLbAmrRYuCYd6bBW2NUbhF0Lq1dAaVRmi9e+d+ci1/TJN4lFNtgqU8T1NOZEvoXNpTYY9bNg
Fzd33KeldtrJuQb47/OxjFT4++rjg1jujKfezdP+OGed33ZH42rrJ36S95Rh09yS8irxH8HNVcDY
Qjq06gC3zPvIeZrgI0O4PildjljAAGaJU6KjF/hf9UoqdBGofKkDhhdz2X3giD0JAU7FDjHKYg/L
Zb/CUbeXJs1woaxvOKK5rbJOVvBFYsalW7l4VdB61roX/8ldKVgpGV2e33yQoGuQbE6KnwQa5nN4
D6tYVGh980CYuUSMb5PqXa22S9lnTk5idn8u6l6uV64LZSVdZtsHcQfguy12rf08hOUqi9uSpVRp
YgRHPoq35dqRHLKJArlPTO4PEzbNRb+ISCe9mUkpJjhj3L6bi4i9E/PCxHphZIV2PZPKWkHEUH+g
9Qbzt55YXSoBsYELR4NDWUdjth2EqpizNvLOo06K5394nnXHVyGXB9O1d1nzYM/WAj4YR3hEOtuO
nQAKifVFUi365DaOJN+VeMfpjcUd2HqlfUSyB8M2K77hRRr03p9aqSD/auV8woLl0XOctldn7Ki2
x06h2sCfkNAXJBh+STpHYBTkZs+oGUhai4goxuBsW+lx9GojYwxooQsnbyJBWfIpetgrYQawP6by
FECKr/Ot/8KhrLtKuYppQco7bZw0B/L/emF+xHojGJMB3RUNipa0AhwOFE0M3RA4tEJyw397YV+A
O4UZupTZsxsUqkBuDg6hU/ysc8D/QQ5eOdtU7hDkZpusvwDBuX4kXbfX8I9DeuXTG/fMPguh3RUe
+V+LtDykQbASJZ7fUvd5ZgOF+MwTGB21WyUAdvQOM3+IMGcUZjFHFt5Bb9rhm6N7zBnezJfWNZuq
Uzs0o/bViNG90ri6QXmHM9wkPxLB1w7uuobpBcRuSQzbMQ544dvS0l843mW2KOHbGzk67KfxP7W0
AgDzmfbBQoAyvCbrDMt1mq76ygJWAPv5eDvkMJ8gzoCsnsyF8gHPiMXpsnQGQYfX0Z3NC74mBsFY
nBUaCrWTsnbnNyZAnRujbc/9yR0uXU4FNV9ymCSBH2iqdUjmwfLQwFpWv88YEXOUtqFRYvBK7m33
u4zs+jFq8NsuoY+q2jBrBJxEGYP7Hc8F55gX+5wIaSq5LPe96hhKq4rv/0Qm+n+7oV9lnxgiNPbO
tSzZ/+ZVLWBdIGsVt5zcRstlNhE2kj2/iW8QzrOMGj7vPj0wFZNwwGcgmSmDeieZh/n9M4KAmeQQ
5yhdmoqz0PC0HdZbaMy7hYW5uojRVOymIK0dOs9sR0MsEiiJQULyocHHXbwxBmPFwCB6jHEg3M18
y0AOaGUhXJX1jW0e5ZWFHIitZfdj76gcAt5SS5fBVMhbP8jBtg3V2YNs7jd1H7BOgWHAyan0g9HS
ki+fDqmUN2L9dk9RSzG5cLV1c0vZ1tHmDTFuVAL6mx97lZrjAdxCPEs8gWxnWJ+FdRyEJlVqvVDI
PhdHjZJp6d8Bt4U3R30WNBf7bR4SyXTFG3yr4q79rUNsLDmoWwNFqY+EqodkbiUpBAJd63KBv+Ii
2/MsQyQG/+VZ0YPbA1ri1GZyEvAh9xZWJU3cNWtZOSLQdLHb/efCHievvJ6zo6Vt/X7EHgVrY9ku
cgJBBsZYKADil9lM3p0SZ2mk9kjs7M2/30IREnFQovj66smYv30FrS/ovhbmUS06YL9bzkiIkSaM
O/ZWCz9rTFok3FzXsvT3hwoFs1/th77nOqxA0tvYF5stI5DMdYtQjp8wE8ByZT04nkf2PkIP9+yP
7YTWqD5pgF+PVNzWkBwzWDV3TvP7lPr9GfyiUzmLyDX+leUvUWANZB+0mbLhDALahBuFVRHpjlif
ZqcbIQT9SHvysbMZ9ItR8cjcKExfVTOdCZpi0lZ800uwp348jseEnY3V+uQCUfhrgpUWlxQ660Eq
Fsjc7HMKLufWVsNpJCLWyMDkQ+qNnX4bXF7tbcdE9VatEDvD4W34LYFCaErHnD8EaHRX9Ja3+tny
ToG/AQBinQ0MKA6zLMdy2B/hW1ry0h6qdMi6hqUu0WExf3u2Kb1Tqb8wswdbaIo9JUfRiNqYyhVI
5F4/KE1iANpMXwoGgOznd0X+hTZV8ybXuQtGGAOdw/C6Zigq+4NUtRE6FwAlUgskmBpJI0tNUeEW
uHQB4I5mmIbintPNWEYAY5aeY6kUAGV5bzJB6SmSfCPC9592x1SxeTlVTdUqgMXtjeQ30QgwdC5t
4t80z8NjB0060SOZoEr0p4B0xhQb+Yc4jnrEPOSdAqXt/vZW0nu8xZ4tNyJEgHd23L/MSJcXkl7y
VISPsCwbx3eO+xwjsIhRfPeXpzT0eCWijGWyWAlpFfpazxfW1+dWdj0y8c8SVw4TftjgRjvn8tRp
zxO7Xtu9THqso11Bi/Ks5voPbxJwva695Fy50o4xYrMQLtpUm2ZPnP+kF/DSMdWtYV9DHSbtHoCT
sZhCfCnh9fqdWOxxmp+lf9TwV8zeoBpn7EBVzAQDeVJBnO7TWQF7X6WgSxO3/j276kyWqEn9crC7
bI9zk5LkOjrPNJd0oM48pOlBDh5+7kuAQ3oPBkyd8alJTRAV01WziaaRlEjoaOi06xgI5KjuHuhz
jjSqsrB+qSV2855LRLWE3Nt3UYtjcN+8WP3LdFYymxf5Z/wfkDxbnKVfjl3b+LhePg5BnLJV0m+/
7w9XS3nKWRX5DuIkQVLHuqxkgqFKrSLm0ticinjB1xX+jLm1F1H19mylCQa1Lb/DERrs7kE+46KB
yo/8/8NQiMD5L+oZ8rUrQxfQDhFFF3l/sYumr5Q/6kDjvczRCDf6Eos246qz/RfYjA1XXc2TUgLC
VBqthtYyoSXNHrqKAU+mPu3vIixW1K1uOS09bYGzgH2jYJ2J7/IKW8VdEDKsK4g46fOhTc1BK9Ky
hj7aiYFiiHG6RGYRJhx0h9y52bPByRin2vFZL9rVQy/7nppfD7/emRyyoWY7WgvSzrM1c9hSqGg7
j0/xsPhV/joqM+PXVflwXY95rlslG8teNezW+vqseiVO2PF5xwWizzJXkmwv8OaWiQTAZ7CEmkTg
11/DLeQ7yZb4xIdgFMANsrIiJMw6k/2pNvwXrwg4oucr+6vVGxizUtO0Cc/s8NZQrL8RPuSf3A/W
0KoKmLMJoBgG8MGSIpgt9nMb8vI4f8nor9k0BQvwq5VG+Yf3pABdHIzgMEOdzzIFBlggg0Q1OZSR
2Q2u+60QuBNtOS3Qb26AiVbuQjbJR633sTutfxNQ0N1DGlPE7I36Nd6HqPC+3SSlt18AmyUg88Zi
t3B68D6clwc1eTx2nJS3AK6qFzfg5oNeZQOrBltP/E9zr33Wq93t7vr7YWbe7/g/K1YDc7aTfKhc
7D5qTYUpy0U12mAETo49klcUIPa9vzoM9kaeEKd1pQ2siR2X/wFz+qYz0cWRHsG52lpor3sfr3OK
d+ktPClEit4YXFu/tUT8ETQEk5owYQifN4QQPdLpG768p2fZ6Buaw1Y9JhFi4EbHN+5G7BPrtOlw
AjfI/gopz6RNuV0Hr0pqHe1XCySiam/4X/hc7kTdUzJT92n8UM2qO6259KjeBSQYPMNzs/Nw5zpc
9JzqGoHIiW6/K/gYRP8zyS7JQVdON2idn1hXctUfpYXuXcRlHQzdcoUlBIkkmDJaCpLFau15g7ep
b+OAhjUg23TsdL91TrasvRfYihgSux7plAv9Xb6587MIroC1IIO/6oS+LtWULfwx5VhyzDlBbfAU
OWO62ocT2Y/MfWCJp0x1XJTU788A8066PSfB11Vz2klwRuwTpNn3Vb0AdflAZAxEjIpAvL1KS7qk
WZK59ZxS4ev7NCJ4/gLwaqcIAmSpvXFY3Oi7fLRV6p9TM4jJkmMldBF64zvym2JznTfnUhqHYaep
7hyXhB7u+Osu68Hamcb5D6ZVRIE1fYRZQGGh7EKJ/CQ6W76e4Cbfar1brD3PVpOybAIMZCgU+UVM
QKV/iHOP0VlJKsUJpwCQpyUJ0TO7gsdKstn5w2MdXhWJtQ1XA/YE2w80O8ZVONsr0BLwQzQWhXtX
dCu2vVSvVu6foZCRS3sxCnufPpSE5599GmJQIJMdLb8yvQejUTO2+Kf4Ov5fo/EdLs1tn9ubKRRc
VsoTDsLS3Yz6HVjRWk2JSkrur0b+jfjQATuquPJBXMs5TPrJq0M+ee4YMTCTOykuUTYgDgkzxbCN
uChKvlz7zQPtjHNQdA/gATDCK3RZtEzpEfVXynK7lQ5z60OiqcFkcCkoK4XQoCW/7OOMIrqA6Hbn
Frmv2BCrr/UK9t0M/g4bbuceMJevOMeOEh3BjHpixdxTjRDSIt3Au4BFsED6nvVT9NvbBJY4AZhK
fWY9QOooCbGC0e5NaWt0hulXvpAdpUfvyC91nfZWrC/Ar049N8EHJMdLd4uLQ3Uv06jcNEHuwXVn
zfue6hzpaUZuHtuLs47h/VWs4drH2X86o5mL9l1SWZ1DcD3ihfftUOh9yKHS3D8djBxuZoWmaAds
1H43K/V21Ly4bNz7Aplo/hn7Ki/6Ax6NDGQ1XjTtLUQcKyN3aCprENpTaQue4XOqWgD5gpqOlYQc
SSh9tEzeL9PBOgxoAQU2RWwmc1aEqFATuPSKzJKny3a4TzX3gdBZyJZEvJpP7Ha2U97m3wAZmzmJ
HQ+hlfY8msguMbR0xtad5SFrnsvjfBRLfaP2b/S79pJX8cfXiS1NbHadEgIMH7sZhFPkUzjMuna3
yc3KpEV6E2ktDfrWVU7esB/dxOm5liCumvgNP98K5RAH2MmAjojvNzuyzxVcLKWCUKi++NHc7ZWw
+uZPS5KzDnn9I82/xbY5rMSdv6jDoJ14BPtqHcDiXvsGNrFK3aGe8n/G+NVnbbBA30OKYX9VpDDj
57x8lT9D2Mx1OuYk5FFbgEvEe7YztRaVOo3jpxUhBfy1xtU4suwFxvBUXvSpqa0fyv2abmfRVsw6
Q6b5/nfC8Ux0VSqV/zRCuh/zHciD1pocJH5hA3Gn3h3Xt+UEndQpAag4kP7W48Tpo+AeHJbIOIK1
VQK3KGFzVaEGubUiCiyn28ux+OWxehukrgh9piEMNu+KsBLShDwPz1McmJ7TVbvZ+hKsgGWdotKs
j58BsFM0JLoC7UtFT0N711y9l+DpNvOmfNSD+mwLmGL3KWsXQUrJTBmSa5NdjUYiYy0mnFbI7g7b
H/nZ1e034xQq/gqBUX1TBR6NVrmaDEWHOUDk12q08zqDbTOasEjZaXMyAjkIhohTfDXhv5smcujB
q9CkwS/FRpwjO43yu24t1DJghfcEGICCwDPhrGkjqXKIBOBYaVqcR3odTgkZoMwEuUk5izOwjy4e
BJM7SF9w5vDT+iyPM6ewvfkEdC8pWvBJLdopOo6L4uaWGJ+NUQhA37AoksTVvqsRbGVQqY2RfNs2
ANHKhwk5RtQFDxdU1zopgOBO5/6Ok0aMfYS/IDdlBg9qWeU2JXSyNG5r9pXCbtM7Nta0/623AX0k
Ah0nAfZUlXix+LzEGW14T10/lVZJdIILWILWI+dSbiQ9VeVUBdQdFY0Pgy4nNiCwPE7Ab47KMZ86
C0LxhrT043Q8BK5ibs6OQp+crMfKGpYf7/jcqfnREfrESZ65UCSfzQ7mPS0nlcW9tvhOkOCB3o6k
U911KTZP0zPSUj5vNVtMQfeJXVXRYH2uJjShpRrCDxemAAmz59wIlBGkJ5dRBfH4S0SZ9XrYoy4i
xBDoaNN9YMZcEX0a1st1tImUnu4IT9qcHg3rV5hBTF06tiz12Rer6o6o6r944N1SzmRIBgixp5Fl
uM/fkHoIWsy+7ylmvRqSEMx9D8csjdE9twXmkMurGzaue3kBzIaS9Uo1Ah7JpReCSGF6rel3wD4l
i7NGEZKnzpEmwBCXUMzvjao4IDxysDEXcoJcdSAqQkgzM/R8sTsqIP3C1w+vdEFQyBWG+uu+jMDq
/JixkVadBr2mNiv4nIlVGscDFSWZTBmXSITaO1EdDJIys4C3dU3fAwkp9qVfYfKqjdPPOKmVFelh
DVEB5PY7GyvOhOubDAJL5Fi8QyhH84+S2jMEH9b3EAglvjnFM+H8FdW4HZtF/5/OAgMzydw3sQ/x
BMvmvI//LyitYTKtr7T1T1BdXm/mDbC17vrfMUvz9nnnsxua4oUOM9MJUPgJjiXbiHzyJQPTRGBr
5fh5C3C1LpPnyxmAAE48VTE2gUR7Fwui9uVNyDW+b+JPnADMUHsJSxauyh7W8Sq16cpF9G4YwVUh
sBD+FeFJEhw6HFULnLYsCxsEmoLfSoTq9THp/172jjpVT1aY1csXuzd5j50KNzdxyk+ytlv0Hfbm
Jaz4bjACD3FZlP1CuiORuSnnVswR2EXxW5jTcdiQ1FEH9uLdfHRWoY6i4TU9duu8TGTsE6GSIWM1
9W6rsp984PWF/CuWY0fZ8t+QOnkx7YdbLI2LR79+nciZiKBl4T4YXVbs+18cMVH9MluDZkQnWtkz
tNOGn58sHSmitah7QRbrC6ZO6A/WNh0WTzCjs4qaOUNJGiSDInEXuXd80G9fQ12ra1Hh01cRVc8y
4rSWuTDAZREqUKxKkf1bNjb9kf3W5kgCt3JJlNXJ8dTnuomByZkJtha3os3PUYLESAfkQwdL/59X
3Lb7GOX2VC3AIi+4LQCin/Tt9iGeKVPHHIDmm91H6NpuD/aTK984j4iw8/0F8a3IVhzxj3Cxhbah
D51qlmX2b5fc1VsN8J2VzZ/TXPofPYC7h6YVfYlqH7fhHNhWrm6BgkNJvBURn2zyIHv4yLQT4jnl
63a0QhJ/bNluEx+gBY7td4TvpflqWPQbNdZ9q/f0gs9mihAUDdJNKFNcNRqfDEWiSY6LyOHo0c0K
sKlfcMdT+4ylG8MNBUrKhYXNNRoCnwuxaseSmmo4upVmhuC6aVA/377VH++DXC2+QCd5wYY1O3jI
8tKnhvGXOmBvhPuaLAAnndODSMwFHf/jVc7OgI3+EvsGHJk7K0WRZ77BYIe5wc/hU26S5CJ6yqDC
9+ucsUfQ+/o2OQ27lfnlajuiNBHV/n9CvQWnTImG5UrxahcgdHoV9Z3Fa1pFIK6NzAELdnd2JF/B
7YOX9avnY9BKJXIK/VG8adAx8DJ9dzmwjbO9PQ6NE+Kd0TZjXVlXcRMpYZvnobeE/vttSrCjyNoQ
1el2OPRftbuU9+YK6Xk0CCI8n2sfXw3XnXl4izFKYsLw95cvMF/OLM4Yy1TBxLPjpDHQVh299UOX
RcSv8As213gOqNl3SbsvohBvkl1h3cURzgb6eYaCmyCMy5C2bUvgz9q4Fvt74YoewUjuVh3vS960
tOPTRmwmQW1YZ/uWpqAIgINiZPamtT1pLkmXHEJ1a8pGC41EvinHZgDzUenbJORAFsiPyJl8iu83
i7zT9OGAQ4CC+3hpBhQkdazskxXej6RFLLYNRToXCaydwi3Jdgk6+9/x61ZcvFMwWmK4nE/mVdzs
turoo1b6/6kGAvaNjBaVnq/shi07PYC4v5vLaflSKgYpPhlWEVIHXgXF3jurYMyxp5L2PrW7tpv2
QiFLP9iG0w7aYvw4/LvEl366nlv1LlyOv1RHlrdbF9AcsYOp9yexi5ysgWi6dLnx7NBOENCAXwpm
KmCL9Jx54K2FmENmNPTZcIMEtxAyyqtkjjfpVytIhZ5BPPgxXRwdg90/0QziY86dzhKa1jzguRcO
H4D9hQRxWSfuoeIa4l15GJZv5fyXCtSsJYlsohNS2E7R/YsyqDw1yBRBJQqF3tP+8BJ/5E3/lB6n
cGmb5u9mfZHjk7gbB0RtOtBrqWvMlPGhjvO/RZ2OC3WyVoUCq/voisdm+CrlvAGJsJXqsGjHA7ID
y9Tp4lGXPGOoGuES73TSjg9w15NDVX8TN/QNEk3xec9A3Ra05tGqZgFcvr4pwXhI+RSTPk8PzILW
vNViEsw+bFGk2PsAHDfhKNHNO1i7/WjjW7hDuGZZ43BFVmD9zMRCuVP0HDAUFRJnFaqzNGkfy3bD
qeEFfrDTFE9oF28oBvwTRMbMLqTNd4ebenm2eVgEh4C8lLnxB6WT7RcBHMl/33UKCY1wgv2oAgeh
iBVhD63w7E4HZDZVuCWP9ABut5EE53Npqg6cZ9WOe2jjX2s3ySi80IhV7JGfk/eUZJ7PeUg59SqT
mAAszbbdDvoC7HCbGlUSaZzIe82LcpklX1+FxaoPfnQ2CFRt+jBxI9U7GFVxHMwhCDw+CtugepgL
rOY1oMsPAGBYrEIh6Q7+J6L1ezb3UJWh8k0gdpdlcuRwfvxB3KJOU1TVA/9r/84qXb80vS+kctwg
GRZ2JKlViMsODuT99Z77ly+58HYp3Sg5kjo+c+59Vxqn+EPfel2nmlWjGwV/0D8FU7o9iErCn4yJ
2m8X6PSEd4bwvq0rhcjxBBv2Fn8jPlWAkOO1ZO6YrW0Q9jm+DveJCsVNcmqODpjY9RhtD+JwhDQh
JdVQ8ywBCrMymO6VC2fHwNWj/K+jzHvFOE9xzY2UBxWcJJyLPkwibRdL+V/LVqDJqt942GZjIzCT
ho7BYmELpgU99B+edfuvv9kDKrC6k5nXOe0xp7ryyv1HzFLT/HBZdhw4qkC6nPZuXDt99Vf3CLeK
lRwMvKOO08fJMdBPC1QaoVxQf8BCXjAMz2gdbhcgKsRrA5N7+fYfvNhsSq6+Fsdt3pXdP4bvJsfF
rsOAD2iayZc34LwBdYHDMZxC0+9V1K0jZifAmjs3JHXgWA6urYGgS7TS+MjSlsM/ThbcQBlmNEDa
Bca4i5OSUnQGIx0XpcKKx5wmCkQ+VUk2htcy6SAUd0EB9eEgQY83/UDSMUvqqmjLbx3POpMOjq9T
JVl9hDr3p49sh1ektpjL/JQpD36+CqLGrqecD6dBalZZBkbeorRlFsuvREwXpWVPfyriHePTC3ED
wur1taWuX7cohdcN8479z4PH2stqa5aoZ3Zdo475BMQYxPlGdV69h5qVjp6QN/oZHnbaXKPOqOOI
ulM8sNNfiWJNF2b3J+fgWdYV4HlrrzJc4QVt2VyN8bgUgT7DHPKKxUI21MyYFe3yHDCl4paqTeCE
Q9HwXLeOc4VSSFtnKp/pzmlzLN0MHywhl0GAz7Ww3sADf5D47riBbxPlK9jBPBef8roApTD5zdFC
wPzpSWsn2HFANFBNgW+yi2Nydq4SZv+f8WTsRk885bfg6Qs1P3dU+6cdtjHe8VWvrWGoTtWf5/nj
KAC1alVNN0pVbGuY6EJotPf7zwV4/Vj9wFdeq7kJGJHmbAQgrW4irG9iStoHwAnDPKag1YAd5eGu
7wRUOdjDubKKzADEnAZ7t5Oz6VR/NoOUeOfspfiJ5rFtyv49ykEYFh4DRRSUdbvdhPZm8yz2TUEQ
kUnAzIkyKBnkExArDjnUlin/g12w8P/8jg2TuOxSjzOYH8WD1J/pyYhmOHJ9r5gIKbbE2oEl5Hrj
/6+yscvn7slMyUCdAd4UKTiC9QnT2Ob2R88zNXEFxaplQlqv/PlrRI/Ro7VAJXLSLNPXCGdKWfMH
gE1qNFzHjtQKSQK8KksYYwX1aLTVoNposwzMELd6WEScuAuBz35EpLSiIvtfNsgfn7d+ckh6itBJ
NLGe4CyFXUJR1+nBZZohqNQAWX9UvCJvE7R9giNNd6Dq/hOEbj2iL35NwNwkpBN2U0JnPEZQW8YM
gRHCZOt0KJK37B0pX4Y0Eeos1qimVRFUSxVUVh0Q+cZ5k3n0xUXXGvRsjRE9WVyrZWJavxtWl1gW
luIA2z4+n5zKM7wc56K8Cs8n4me8dlq2baozrBUuW8B8aGFHyjoWO2f5kp1EK2RVVT4I3snBZQ/j
Hvgt8FuCxztPWEI8D6MD3/2UJV1tgHsU4ibSRoPuw/dhRjqnoQbGmZzNyyZUM0wRPtNSDwczLCQT
7kV79LmR1Yy3RK0idFXs2NAmpSo9XujvzwYpZU3WFSgAjG8rE6wG9DfVSSQegw7vYcRQDfIhhK/o
CQQtwPXdckfpP/Z3ZfFSa23m3lBLO1O6yUq0kr2gQ4rraPJOdXEyI6gRbSVyxeydseurmSbUinSQ
VCuU1y591xURzngZm3RCq4CrmGrJhJziZ86g1LLDEmFY7RZw5r5HNebkMc4WpV38YLdGgLk+OuBc
ExbIdp3vNzEj9HelykKZ2qR6puiwGiRN6GdKtznABhJFHs55niFrpNiYkN2KDUwvV6BfQypmE3Ss
diYEf5iYSLjKrAt0B2jXgELicfBQEnaJW0eJgs5Es/1DXK9M/2/82LW9i4KfjyokWoWc5ciT90v4
W1hbG7wQvIGxsLslJymDxeuvBqYnoSRJ6cyXtO6BxfnzzPNuXEztfsBPC6GBdvidiEFlLqGGrkl4
4wj5dbrr+tRutERA0JxTrTznVPZZ/b+W415rD3qbUBas+W2ocwydzGe3DgM41Ls10d41r8it01Ac
iWus7iUSDHrvC8mk7j2Z+JsqSkk6VsIbmCb71JzgkBLuegJiMO9lgbl7TQA6W8GARhUOm6ES0tfU
60Y9YoM9YrmEUUHVNLpATCgv8s18BIwCd3P33f/A+9C9ZA39TxTenFr8DunUhklL6F0Pz8O5P9kQ
ttFXdhCbAbMU82lLOMbiuyuO8jPltE1TMNrUcYgOXYR3vQyfBUck6xIVaa4OWJrx3f30Ozrf2s1b
pG1XxmTM9GAopBZsE8pfui9KQRE5853GXDd12pD8Vv7CXasri4yPQL5JLI0SXFv/BDQVPYgIiyJP
aU92IhSZO9AihteMV7GyUop9buADU1jJoPMzyH3zgiMzemVkYKPyqfeFSfcLbfCLYrt7W0SSyRyJ
lSnocMTpWZdUU+prpJlBptnn1D3Z9dOyHyMghjFaAcSXB0dCjWV+LNVCLgUeLLr+99R5Hzbm9i1N
EELqibN1fDLo1pe9o3ns7thy3zBIvt3ihDjkRFpHzEnjnxuAxPpuMVV8PrQ5ETQARj9+BchUr7FH
jtWqtZyIjFvA9f0bcU2E4IEaTnpG36EOA5D1FgWC5CBMsiEQDUvoV8+41inDZZPNiRlT5PBELRV0
12HDOuecGlAEEtQddd6uUrf8N6jMIYBl9lrwty3gCnXfKaX9Avahy1tTYAWhyPa5btbJA29nRMh4
Gvhr5bJCIdnnKTgTOmhO7bNQUMdPTaGirEyL49yMSIWu15JW7AKDNfKuDnYDtgi+zsjTS+rSxd5T
JIEF6EKH/vUOinJR071yHnaxPOlOSR98ARau0eQ9dUlc5HhuGwFD6dSLr9Tyk6NCkBCk7oScZlad
Em0AT8HRYoTmZrqK/COY3KXVTbS5d6Yx7tcdUV/Pfxr1W9DeGDv2zUN3miCU+N24Y+Nsf4Ybg8N3
y3Y+Yi0HZrSZ6qMpzRlzL4891vEQlYdjfdLObXuTCzIkJ1HyeoBRJ2zY/ELsykL+XBBUEKzgudkn
rx8BgJVhvHPZ4yXywb/MzgQxJla0gXffCqWruOZC1OyICTrvj4oMpjdPmCYCbyGyoFbhIbSNfVGH
wNMHUVQp1fzwqZQo2PlhpKx35W/Tu0lbCN5i7P2pYaviU3zjTe7gGE56JLpA3Yz+2js/Y2OQvIp4
BRHyZvy7Ni1KdCVuCIDIL1MrB2DQ79PJOnmeh+rccQB0Sg++M2vFgyjSTnuDHKUSd892n1bWyc10
8n+IHsY6XK7lWER/KQr2T6vW1V59MlJVBhk5Fs5XbHXNrIMuMMHwlG94KCQu0iDB6HGCYyBJh4X/
6HxDi8Kgz+cMgfvk0XBpnVlgvEqSYcg4Nu5INUPslEeKTB0sp07nrIKOiYdbicGprNW0VTrLFgXQ
vISnocPLyzaAI0u891X7Y/GuZFU43ZKuMbWdWzlm3aS5TA4P5kHocbFqxajPCf5SSifUB+DBruWL
z7qWTaIVNljcLU0cc29dTVtG/uAEzSEg1QCPxMoQVtHrR1xpxNKiWGS4RN5g2Nz4YPhZzh6qmlqC
r9MTjNBU38QdV3auRA8i+IvXX3RdqDUgA9A4UmBqtkk0T7U2ASXMNQDHX8JEU9UBoZyrZLCQ29iE
oixQgsPYUw6o+8xBJZPqSYdK5XOF8A6003jAgAZe+0+hjGmbXHQqRKiPl4xaqxOiGSf7opqXu3LU
IKSnft05R+g5jihiexE3A68CVsoaOMKQdXDZ7TnuxIAfzf3vjeCfUe9lCytqfwY+1uFZ96Pf3iiN
A2rpp8bp+DU5TNv+fI287mAgFUb1eQBsOXBopPXOHHa2DNkCuSnP/9Wm4KFniZe78WBpzFfCsnAo
bHguvMJvh+OpjKT2oPilW5DpBgaPTjWA+ogeATj7/795SBwy66i+1mV4cYi7LHM24nkMou+VWjPx
fJOGzhVXQ6XsN3LUWMe7HswKhN0Nron3xCrG/YzFuED7JkDvJMRh+/XtVc0DHwZoJ+qR8xes06L2
cfYST4Qv1AYNqn/uoqHNIuH+Gh+zndO8cAFM743ZSLr+KoOTEo03tqVNXfPYUZol826bK8rbFOMw
dkr16RWJraxYYYgCbET1P/8Hlj18aNCHOyin0r1AEo821bpfG3Vgi3B86mf7zy4ZO5wbyXIn8q5d
ZQXPGJGJcTYQ7QkkUfC3XxK9gD8ockfYFCXA2yQZ4/OI+hCU/L+5ELimPAEs5q8OTTLbwWGGt1Z9
dUZDIB4Dkjnolvv2i7V7YqUTqnRLBfWBPVaaTYtznItA3d5QN0Qut2e8Zvba0zXOotMmsm9syIrd
7ARaGYDWJluEbH3KYLE8Qa40aDnJkx2AT2xqFdqpdlMjl1HVftPcOarKyUD9pWme3shrmlywbcLv
ZKheDA4IPg6kiFtwucEOvvKHsFa6tveQAcx3NNYBD0WV/+6JXoJyuOb8Lxuj2uL42jCgfseSmKJZ
b5IoC7ULIMCmo6VKfXSiDiWBE+6rv5ajPLUJ1ZYiljUkGcNVO7CfsqC0hShTk03caTakJRprF7aC
hIZOwnrS3JsmHqRuqT3rPGhddnt2rl1rBk0ZiTzAobO5QCJL/LUapojwUSoStuBceaZTu8UbM869
YZLd5NgQ5X+MBL2VpKnynW9uo8enJr4RaVrjetBpj1geFmn8bbJtauz47Iy1hzQT2pKjOSxiStJC
dsatVrWow9m3PZrFsHY63CcfCN8kdtbeYxT/NJmw3gnX0MlSq+U8k736ea6TjPCBukMztGyxycU4
EMgqdpJfUUvKdNePtL2OFMFLeT7XZccLXyhGj1a2wFf2xTKNoX3qJEuu2R+dtbG09ifKnNnPiqx4
2419CEPjIY/+3opwZp+lpb2hyL0XI2C+zwg7PuDpkFC1qhsskHu2wsZsbkjfnJsqEob/Nb7MUZL/
e6yw6evDw0qQ/0RKr4DxCmntjD+qNG8eachcjP9LpJorkNRg5NFHv/VAW5yNcjwn3dxOFlcXqRI2
EpZR3syCeIrPowAsnwNUA3b1TNdBGHok3jEsRMbss2lglcG5X8x5kXnIJD6jnadla9bmaWsDfuOz
r4SXagXgBFF1fc7zTqxkQdacGjH2i2MKiGV4caSU3aeEP017b3BWjJEsZqnse/PGm/xCBBVHJVmI
pk7bTwP0KfLH1BDM6Lp8UcrSRzv4L1u+Gvhhv2271/r5yB3RVqbmQNnxAXkl7MjCMUim4r6V+GR4
kC0xLsrH8YDkARyE2FW15QzIpgjrmCnjt1W5N8/7giub6yQZh7M538jze5zo6f/VpXUpsO7Opi9W
VWbL43XE1wU7H1+pFGaa0AZsSlznPG75aoIWdX+A063KD0TsZ8/hkQjFM6YtqB0LoLz4/DSZCTtv
Ej5k2EQXnVssdzaERaa2ElA4WenNrVYfrzyNyBCdiiBxDbETkzoLfA6ogwtZPhQHb7XCfJnY6uC2
JwqPcqrZORAnsMhu0KxTUiMO0I3uUz4evUGCEllh0IFeEybvXma0M/CIgndm6lMJaiqpUmc5utCK
spWMW65DrCq9aMjkEGvvr+I+ydJxVo6Z76eOjxoHZbv54trP05ELwygaMPJqJTIL5np3rQo96aFo
+UKjcww/1Ufn5Kua2q9V/yOu8gfMBJD+PtL7TVcCW9R5WGxCRLVowa+KHOV1exRsM+uSeV+1DQDM
ecRX848MPkJhbj8iG5JrUGAvk8F0MBKdrbyIRUDSGZAHqh0XNClliif11Y+6m8I/7uJ3oXGqSgSL
UPENLDac/DT7tsbIapVIFX/M9MZfUGegc/FBnY0N09NfqeU8bSHmrPMtdphjExK6OGE68xmzg+vu
Lj52m2EP4GX2klmT1T/TMV5AOoAu40AGPkGdF74LYwuGxK8McrID2oPNgzS0vLDG2r0DDKHMbw2N
Q//z6MhpB7GQBxQ468joIeLpFH87ncCOyp2cx1bQOrGptja9zZvLew3IsUSudJL9BHpuazKf4h56
LYGu03QTzdkkixhAMyko59GekfabRRI1V7w5ceWiTWjmtao5bnNA2pxplr3xKXiBeZqKPb6a/qRa
ogSIhzMPFzwxvUsJoFzng4UPVLk2U8u/72lSuRCiSx8NA7a5daxDTbFuof0sz8yw1dMWVfelLhNy
tRyHWLff5v5YkaSNOCdY2PxAlToUWaeo6+4dXAaZAPr84AJ/tzmbS69dQsnegUQwZ1LiaD89iDm+
bIbgXHaE5xrjHUZvmoHycB4DBQe+2a7O3QykgCMq9kYEfkRDYPnK2Not53R2RfL3YQEgCK6FN4nr
2BSoZgx2YRmD5kARPaa/K4biaW0WbCY6NKYSQFL7/R1WKdDA4u/MAS/3lJzTv5gyLVFRmTYuyjnK
tgl2SD9M3RcMie+rBh+mPI2CvqiXzFJNHOgSuqrARlGK8WO4uMruF7WE2h88B7XM2H/R3/hBFewP
igq55khDOff+WiXGVWDIPgk5GyCc12MyGCPej3T4vSsbUY7sziocqHyK2ifYgC7cq4VbWL2SCg8W
HZ5mAHtRPuX6RAWzUDN7GXbUu3ANlX0JOAuA94dgUM0ClXsVYjGgfs+M53hj0gCZ2a4mOldgk5xH
BJ5hrpe5Xf/6lchv+T/o6zZ5RxrJoyivk2CDZtEeBpNksKtU5imwWqbHtVXdvrCF0y8U+cwaUAeQ
LObQ4WviUKfssi+uV3SGZxIbTkfg9dC9f6ZH5kEWOR0pthb4wLqXq6Mpb4temdo76nhHbomo6nwS
dCBIw748Aev3M+nEmiKfbtgJJv27bAuFzOw0bCFaSGJyO7xRCkigHxLZWuJzHgJCfahPIPPhbTyV
afC3o6jNEU0YpFGhwKr79myOeqq/wAeq2aekBTS8VZmegtUStpQut8MA1kyrK0TLTwoShYsG4FQX
a1aoiV/iyUwtzV09ZRkz7hPdTZK0wwrFrUycB0tAW8p5u8VOwT+AQgVltc8WJqqb8BaTlLt1PRME
9Bbf35cOmKKz1rRmYK0AXjh/UFoiQbUPfxYUIJFNqlWBy5VAT89TViSOxjCoSN9bAiE5cWpQCnmL
7Oc73ahfhY5X3pCxrtNPXwRXj9/kQ61HKsLwuRDp6Jhlnp/aNkBnJ2b5/GpHVqrOtDufLwPjgAY5
6TFJkaThGJoDAxqHXkB8gfYfAedAZy/+xsIoiXJgw2nzsNa3C9BsbrAmGI7llryxpC+sfCXiSbFY
0JV4C7YsvPIOO8bchuip7bRjJ8ayw7lSqObx3MqsizT6ptsjJr/RcVTArbmwyk+d+sNCxRT45HDj
HSHG3+uNZI+cMBU/ykXkFXdQREbWd+fjWfOgXlxubMJZBYlZq2GQuWaHXhUb8/14b8Mk0CKnIhMQ
EIekX5mjr6ptE2tM4BpCZW1r+8E+0K3gUlqA99vRu01o2Hm+mc9dr48YSkedA4+vHtETxzsHe9ce
n59HydHyksAJmTIXvmwz9ozRixPrO8lKyAt+w33i0fntlgxeL5N9cK2XaF+2LsdCA0ljfavafa+q
VfoR9fOsPVfu49Lvr6OsINcRoLTSfDGH//GjUkGqIE3SMA55Lp+hiLPLd2irGfwut+YUOmXLsrCX
fBgYa0QKUqbcbg3FPwZL8wjFaUdh1WB+l5c+rPq6zuEo+m0fo5GvKgfs7gaEvpyhKoof0Q91KFI4
Oo7MLqgvUuiqB2uLzsDddAvvgEuxlaflO9392y2q04krwR2+fvWN04WaSG+EjDl24ZoQ1K5yOxXJ
fVSQWeH1iTo/uYt4EfKf7tqWfnLuD1HUPi2+ZmcFR+HLk466tuNgTPYKqREgqcyriTt/endSDR6K
jpmZaP/acr4TJrqkASHEM0TLX1uqmAPoa/sE8IV7Bu8ltkyWbmcX4YjNsf/xhpDeGDV657RVPjTa
Zm1tOgRio+10crFCwyrOsk1jkqGYe7F8PGwHpO73mingv+2Ccqnznw1v8QSe197AybC5q4oBoRsw
gTTXdFVNXZfrxaGcBUiPVRwDBvhY5C1HQ2AAopdBinshW4eTR/wER6G9zbLMi8IFFW6xFQEL/mkZ
XXDH9oC6bxShd21BkIBkTNg/dtLbVkW31rv/2MCNbb07PP8AejkeysqlkIDuZkrEeWhdMCfV1cCn
zSGXTyJgj2amvZn05J19+3JVQMtbC7o5bd7pNUejTpTFN5h+TyDIdmSHSx7uj34Aa4/Vpax4GsFe
+HfBhf4WfeX3RJ6s0vZUUABp2vuZWPVV0XekP0LyoIr7zNIoH2YQ/oVObyZc4ITdjOe83AbZTfwL
/wZTLeVqLTzk7sdnbBz5sdzcqoViociqaMfA/zMvq2qnnfLa9N7Lr3IgOuDoOVHTI4I43gTzu1ST
q2PBmBqaaJw5dnj+WfsN8NOABfm+LUZWpU0bIugz2smHHCyN95/apkw3tCoxuKRFi7TNHB0YP2kO
yWG9AuKB0dce6bTFTrE7sUMAfw3SDMfs4piJ8vDAAC8DOcRmSZ8W0ec7rRlSJH3jbQQawnHOzSUZ
wdNZ8q5W4rG5u+gdm6O97Jt8DHXTAvSPiM8/hYxfzal/BkNPDaun1x4qtNRVCAIquzaMdrQIFc7E
0phFOeeBkMhrySOqmModMbQZJGrsa/xkmeMh+mU97AoDgROU7V57uiItUZZmKnYPBYRS9NUu2d2O
X4EwEF1yHEFYqnm06d/75Ti7wnyl+2G2jTZvvz7FXlm0nSf4XAvapn4R58E7BjXELvXib9+3Fo2m
k+3KsxdUvaHmOQz2DibgTLgoXcYl4GsgoRlpAPxSHndEfs84Ns2vWdf0IJsyV6WRgXk+4+CVCpNH
itmkwdUyRkFPNxRlgfGTBy7hw+gWvaqJsQV2SxYKXzYl1T5mUh0Sa/N5eDpxAP0RCOaYgdkSJJOq
Szpeu7+Fon7ft58dAiuGzX87sl7T7mZl11MDXJ5YZTEaGCPFhJ0xmVsqSdybMCMvBc5NAI+kIWaX
6MPlk8czRPJP69R+27PBULhFgYMeitg+VDuEKSdA/w6WQqf0r7o1WaQbwcOLDf3i6NckXR+ZkjXI
Urvjb/EWR2W8+Tdbg/38LqdhTTR5NnwrkbKqepipMqNsZreTVQwtRNl63MTGZsSGb3Ein3GKwQj+
FerNTDZmxd6klVHkZVnrDmPgrX3fH0glftl91uMX+LtmnNKvpYoTUjNAct0kCf8JHA/MjSyzwJiF
8iEsOFnOAfjN5uIop4kI6tg7Ez6jJJd6T7ez1kw+4EflLJjxc/b5z4cZ7A12EZB4BpTY5wP96U8/
28X82b2Zy55XKr91Vcalte/u4SdSxVlqnUu3QZfat8Dr5PEo8sykjgU6xSOQjdppETrmYk4/mFmp
CJNgSgZD6/d9pXzixK+HB2QvHKWW2/g60O1amwU8Ggv8mw37SCS5N+MXH+DfczWuaJgnAv1OFksP
VpLuXVhQpVuNKQECcipB+37iJtBqsTZ9BhsTKW/MtvKmbNvLkx/GXvBL20KVmmfhnfIBGJFY9bI4
zsFYjOkGHvMCREig4HroK50arVYfYtc/tg3Ole/7ikwd5UUHvJF6uDxjhGEgaauxNHDT3bgJyx8m
MRJN8+LgkUCCQBvqKOfl8awcFwS3ZPlmj/58+Bs3CxYcdJyREWZsKHSxQbr/TIoO7ouoQ6fWmQcy
uMU6Fvpo4LCm7eb8Avz61C2a31VuUbs5j+5fN9TB/qPTIcxjes2DEE5LiKSQTria4PWQg9ZuCdn9
JANniR7Z4bIaPqmuEFS30a5q8Xdui1jkkwAVLwQSJCeU7oiri09BgE5YsBPoaVttHz1z0bcPvROk
zZTcpxRdI+CR3TThwD5tCFm9e7/MtCUu8diOx2tIt/emY7anQ9c29WthDso2bePaJ46+MyOKgjzK
ixJNTbyVbemWUnfootlBMiviGqSOyPo5vYmOCbTwZcGkG31PkM0SxGjgfUnSIplTxEXYZy8f7VNc
ANDmWkCJm9JsYNYugI/NPPTJgpLs6VsG4jf7yTyK2Em6OMEqTdBJ9GhebOFkkzfbgIVILBlJ1TbW
NaCbXsQDzRRu3u+LUASZFHuvlnlxzruzllRTAHRtMhmUFsfs2WHced0f2LqLMiF6wwjsOnOqV+iK
Utlkf1T4ebzLi4hwoSEjBQrA2hN/H04r/+hOsTor0E3LlSKDcRVk7TO0Lp1wVzcYxHzfRW44bvfz
9zBmVSjnMicxATCW4f0tE6D850KYh452tfgAI535yzoWc7xu0qf1SHTWbSlBfMwch7sgHHBKD7/k
WVytanCfDpp/DaXldViBVZ0tjgDZGoLMjBaRLzkF+1hdqSRl9UzoMtJcaK+9vqoArOL/pICu7CEN
HpKNG35s5f5vlovpstq6jJlkN/7RfRXgvRi3HdB4QjgwmBBUnFURe0Xy7LYJzwdK8o3Nlf7q1eNe
g3IAwz4SJIA0VIuyUpB6pa8uvPCW4sNMiX8pIMMBOoxKz0L+ZTOz8Kww+3GWaS8o2aDtnPppVvhI
k6uLB+1iT37pnhSTjQ1JwwWYAok+h6IrDeQumqBOlqo+VvuO+2jejYb+L/qHZYK3Ri4KyUKeGBED
4gRsRuswOtKs/N5YewbUWU9xTMyCPtKCqN5NoSMUCMFJvGnhPBAemzUfWBV2L/qUnJJpkfIcr/HR
X5SB024y6CAZKfImHAVFVtz6D4/VVHFXEOwvn4vF5vSAannpqR9GxFmBynsIM6YvRnvAJxiSxK/H
sik1JG0zYOhgYQdGeTNNYQtN9vPky6DFJ0GviiC4TtNp+fwczcfotUnNyIPKy7WvW/fyuFHcGMwY
EUVsHQ3bHzzHIPeM4rhVHRPYZUw6TnDEBQHcwxbX/LcdrXY5iTPM+kUhmh8p3ycRYs06FHzS3NNq
jBrJY/fZue3yXTd6OjR2s3FegLJTa+gQz1pyyvC7/hfZNmOmtadR0qDM3xW9r34b/uNOo2Z8HzeP
476VCsY53Z0hl2NUF0wBnans8gzx9jcADxNR5HN3IDt3xHDf2cdN3tnVHG6WMZdVcoBK8UsQDbd+
HsxbW5BDNvGtxVghTdKTiFGBf/SDZJn1Kw3Ee0SkmGA5YsAe+5HtWbjeK77pu3ROmQPC0tEsQwy4
7u2IhHYP1cBizYlObz1PD1HKoEmjrB7WHu7hDWUM4flWz7cQ/P6wF0TG9B/fGbtFfegGeBN6BhlJ
L+fm+v7Qjg+j9BSjot6l6DtAjsSM0xEVxkvR/yNjxhxUc3B9g8wG3F9MCaabE94/PXBXlD1rXsuC
Trm+IasF3zef74K8IBRyYVbOqaEOG69rCCYWGJCTcWTbO8tuRenOaDD2cmwQagrhXgy1xcIKw293
yPjnk1OH2CHSWgk6sDyi+wf7JDsCaQtKzOxXOFENJ/+nNPUj/9kEvIoKUrcowAS7jHMagaaggamX
mrzMfyylaqEgN+iQ0P2BoR0qwkx7GUrEVTaiPaZZoug0B8o+VS0uHbWqmuScTbUDJhvkda+HcGBw
osFN8g7y9i1qqOs6nAuCjrXX1hVQA2HHdpBHRHFcPfc69ez+lo1MXkYKzr3WAjoYspVMML0Qu+2j
WCstwdSvqufn551/2ICdfHKmppAqrZdEue/ktmS7GdPH025iFYMahBdc39A8QVuoL/fwJC1Pr2H/
U5PmGhQi5LZrljRTB/huqm9sWM3wgbXzBiqH4lX2X3+rRLsArzckXKe89xoxzp4uXGdishAjsfOS
1GplGxITK5U9E58orITfbE5ObusdNWAp8t/8N/OAQupM2w1Du0ylhWW6AYJeBa2Ivs3nrVnWk5+w
nte9oiBQsO0GmgWxyA9/QtTXBvPHuC7idRk3JvhhTut9Krad9b/4TqwxCXU4b/7g4S3BJxc016wN
2ofqHKNE5TeUysEPEcoQHmx+oWVBoL7sV0aPt+KyNS8UtXUfnDRjrjCmhk6YCNbq/0w7w0YyOs9a
ImCBpzFtfIsgMDdofUW19AoH2F/sq3bwYF90Z8r9CFpvBxiyFXq4auLgdsdM/HGC1Vf1tk6gwwfb
x6jKinDCzlagX8ATlLYD+yE7OA6Hdhb8O5HEA3gaQLhiV+sKc2GxHpM/PXrBQKMXyLOHHVg1+LqZ
s5q/56o/4ixtFSAw8sK1mfon60VtM9t0iSjR01StK264fmO857C3a1Zhl9HbmoAlED0JG9JFPGNN
qjwumO116Wu/lIJe7uw7h4HSe478jFYVMPSZimSA6yt8njxHiJMf2k3AY9IQucD/nTR9nRhKlnmH
LkDxV2AGLzo3s/F7raSP1Jbyid7+ZJGMP5lTPKwty/sfiAXJCdgfbuR4BHnbx6/7FWuyOuvj1Hbw
1fM+6VKdn8/nmarPgecQBaHH2Hz3WJAOOH574rgDx648KeHH7gHYxR6TlSO/rrRvIyq7M/ip86V8
iavmnvjvirvuYtYaDiWxYulekiubDDkl8ynOFx33hgEdBVSXI9CFcmmuKAA80noicDPmnl6RIfAB
pC4BMWP8VxaGK0ZxHpf7qp0p1xj+i7Sk6UYdGJvZ9+Ib8WQn3rZyO+3OHip0z1CtOeUOsQsIg67V
J5qDD8UK7t9oyJxRl6vMJ85E9uRNqt0hd2qmJWWc4DrhMKk/RoujlGHJB/bZoDiEWrGK4jUgpLs2
Rw8Nz1lyZcu2h6PQY6Wj0DWULbg3V5//o+C2KTpv1rb6r01wtbhquQtuM6zve0MdIgoF4b12nb8e
fFLMbjG5lAFEasB5rJ4O4IUwpN7u7n8tRELIEH1OsFtQbMPcwT5pFIlS/0Sr8Yrg50sE5fpcS8Ct
vjScYfUPV+oqj3XNME0hUGHhnHfsxM5JpeL6vHvolEfw6OXEY3/BpUKpQF0FVIwO6O/D7YA7/y2c
Aev2qen5zNaR6fn8ERfDnIRpp/WmhTJm3KnrcHtDk/o4vqPtzsNMFG6vZN4xjgwGTTDfkZGsP/ff
waGpxstZEOjZ9lIX5M+G5Efpp6Y8dyPlwRMKgj8H46PwPPx7d9S27I5+XKC7B4/tEv2SJZVEMD3y
c6zCSctw2D1OKo1IodBe+5bolV9Jo8Vbnn6A0DMwmNPVDzeAsXpFHKvzb0n9hvEV1ks9PZ5+iGN3
btV1DeHcPSOaLfYrDJGv2XEdO4oqwdcYxxVOI6sA+CIX47U8mPL8s567NXZWf72FJIY9okMiWY/i
Ify+99KL4lRPkMnuC3N3g/721jTTR0wc91OtOBLklg7/kjw7BMr5aNStWw1u6Vsmexl4qPNc2LNE
1ewL5Rr3IEVN0QvnyTdV4z4NbB2bGfoFm/pXXqXrRvJO3bN7UQ7wAPzBUTZAiv+TgqGHVFgnNDZB
D8KSjNkNGfJTFuO/g62jz1fyP/hnJgilu3e4e3mq7m1fVX0fu0v/gXSQyV58ZEbEa+oDBNls6LHh
L+evf8phZyOTGAeUvFwRjLkNowBx5l+7JhViD9F9oqfDpGRQWuZvmM94TL3nMP5HS9/xxKCintCP
mXIHEeMBknVsW+CD4cZri3Jt6ynOH6LI7K6YCbmG7985za81fRdrnohB9mMuv0OWWbOqD8eS+Z4p
WLyJqChlpelaRImNiaF8xKrc6pJ4WV79U7qn+kIBftIlA16EN7yedoxSv+5H65JkwVoyL4z3TAY4
ddhqIdfAYX4QftPEPwYYE6yqSryGKi4sDrixdmzr9zO3nwf/cTtCdtBHUEHjEbBs9bobl+EhFW5g
PGKGXsfUwmUngxlqRFiS5Dq78+jGfW8tzrj+r83xwXM4AIFdeGB43Row0vG9fW2FAeFCZhqctIPM
VW9QWR5hSEHlZr4+Nmg39+ouGXFXBkzXwPhnsUlYrEd0zo8Uec0Wfg17cL/UelTVXFDIL2q5oszH
8Favwk8xfwTL6/lshfQqHg60pOB1Cspd9+t+b16G+72Yrbbouc0TTWpnhm0EMDa3nd2yjAgpMJBi
942ryYkYUwbpcZ+/GbiIBsmkVw3rRgyE4yeXG5Fxj6JA1fjVFiB2nqzroy7AYPIeje+3nmSNGs5c
l+ZQm2t3L2SfiB7bAuW7dDhWgqA0Df53jtkD6iiNCBAkwrUwOh63Q+RJJPzXO3eI82VdUiVmXHQz
olPbvJeX9fEPP4kuL5p4BvxuOUA2O2cZektc2pUgEcKN++ztDNNpEO7INi/RDTBTzTIUrNXUAkDQ
eQWWVFhoT1Yi4nDmnC/FLCEKyPU+HWYNgSstoI9tfk/qiXmxCZNr96h+nWq8ncPa9AOiKwH37M6z
H8zx7Px7GCzlCfZyOJd//5DcYNyuWdZlu2WqRshzIWUZzzDpDhXTHfScqPc2fAznSUjuS6dcUeIS
Vm8ZTfzWEu0pDU7XNs4sSwUH/SSAqWFSzPcn5+BPT1W1ISCV3Xk5YfVVkyOjvnw88f53Zo1fSE/J
PoJ90r3C4EPjxVgixSCyF7HIMT8r/X+XhsfeOmzmxOjS8EoWehlYLdi2WKC/HwAYQbeUN/Lx3ap+
5kKrY9Vj1YdnyeC8qUTu3cXNAHdP6Y1SshOGMRIAls+bsoIHYjcmm/g8rpmYPCSldg8/533LbCoJ
OLLNlnp5JKjIXC9kCgxpA9B4fGy/jccpsXYJ3q330iD3TqvD8+sLY99OfEsjKb1c6ja3LMoJkQme
8sDsHfqNOP8AjoBMJ40h2sJr4lr9EzU3gzDMaL4jBmly/Lgm3937Xg9pWLD7if2MrgO/ZWLjHwA0
Wb2Jsr/W1xzjQBAxrTFcBj7e+FxCgOhl3hd7++UcdcIst6oG/yipkBR8oFbwILqfzDTLDQJ5reTI
GSkl1M44e115knBbpZ6hjYJYLy745yG8oSJu8nRr0B4vXbTOM06cpqiMoJ4W0zRCUlb8SX+h/uwB
9abhYv2t+aXHVYwvxcaV+6rMhHOSGJG8nrBq6SAuy7/F8BPo+QfvJtBv24jBr8h20pf+qQHjPITh
LGqXJ1D6Jtb08e6zFsfz5zu5u4ntmN4/pGcd5Fx5yH5Zri0CvKnEWGgSkWnwepVZD3wekd/TpFAS
bhPAlkAraI9FF3aiBj5RMlEXR8pPeDq6fI7qr+s3TzzYzaX0IW1WhGtgnYvhNULTkt2lVLkPA5eq
U1tJyGxNOBbuuLT2UU3LtsarVLDzz/olx1MIHTdDaBX/3VcmNnSE4g7Hd9kiBotQV1autv3cR7jr
pohfUkhJXDUi4zpV9o0m+QDtvjC58+xZxCz8YbwFKqyWAfzll/edHXwxtuWImJ7+9p00hO7opxFV
B+wwTM51iXfaq+CfpOgySMmN0qsNXgWDzb3X3KFPh42vXzdHzhRFfEdKjMmf/88g3F9mTWYtmdW5
tRjLO9g7Q5ULS7KJdsIKv7PcxcL8OSQZ55kojGd+d8X1EdkJpXNQTL0N4ctuDptuVt8tOWzo+k2x
wr7OLjvGkRse/rqGIXuDmQd4aHR9skui0gjO1Rv+Uotc6Rmy2jMydexaPlXvQSYZwvPKBTDi2mb7
GtV1TxcjeGixuNQ9u/zbGTIUZELeu2yqUuZb3tABY9DaxldZ3961zDDJ9MsMmEtGTG8+oQJNpeay
R2aL0fspkaYcNqqH/qDsmAmd5UNPlSmoNGPEchAxLEXf5dndQmeaoWIctDIVM2ROGk6Xt/yn+v54
BFE6kT6wMU3+uhKi24SsymvWtpSCFOtLgxvA2bSsUiBgZi8fWaX9uoJ9NglECC3nyWSok+8l/472
su21lt8uaUHackuxmjwlErGm5n464pe/gwF+Ha8myIpEtUoxG1jAOM2bcUN6eLb50Qkcm2aClbdI
wT5E4plmdSHJJ7lTZh72di5J5Q1bGc6TpUHjfUQY3SgDNKiH5cR3K9coE/4lkWaiVGLxe6spWvmI
EdyohZyj86kdeK6L7JtxrBWuNVStALouU2hOINwiZ78uySO4z8zcS7a6XXH+olfdaL1BH3iZmByW
aX5Pq53nh0AbI9ietNe/FscRhHFTsyjN+zFWNRaHSsaMfbpcak2EIzZaNDUml9O1INRzEiL+BKZw
O4PZpaf6WbvLNYSXQnRsfpOEYRv/nGrY2hRxlzKUdBbY5gWIz+4TtNeLtQOLlSnxS5jbySmjDl11
+onk7p0C2KqqykUtE8rDOc2wc77LT5EkQD0wh2BQKDSIYClnVsBDQr+a3dv6Q1V33hrnDfOBO84h
oUxZ6S7jF6ByzMtr8ABOfDSXQNFJtWzMhNMO/ljvE0PrRiDlGqXD5WYpEYujt63k4s9JlvoWSleY
b5cNL5mM9ioOX+m6IZbfmqwCTHCKEh9ijP5o663IyE85V213bKUEB9NCvnujyg3cFfU4dYdKbi3g
IfSKAXbTv/iD9AHg75PE3c/aR7x/Jy4uiG7BvzQ35RyHuxqPYAKQzMqLrKflWI5YtLd7xdQhaQ/j
hKOySTNnOSd7O+2qYxVmSXc3i0Y0lAj9zBBAh8RtwbNmH4dENIWEyDIe58YJ5JlG+LQjL1B7eE1p
G/CQcrft9jQM4w8b+JDCCFFSAG8grS22smJqLCZuBH25fn51y3kfXgs+tf3mlWHA2clTsaCWORtF
2xZUxL73ZRRiWRkxXvKCg3V7OWI3ygSIZ75wj0lf6pVd/xGiGSOicbG/ByMz/qLEXVHbmpfmZcl9
/HM064PKX+0wtMpc4oUTnT0cNH8ABsYlEmGxQYDq1gJ4nn7brHWM6nAhJb0I3oJazuFdKeE3Uj73
0gMLBOZhNoYEzOfCHTj6mhJxYqibUyQk0TSc9977AMzBEK7dZVVMvWpzb+y8OXsuZDywFqEuQ126
qYFj9IFs8A9Yy7Y36p1DymaApGtXNSeey1j4+//bmP1qdJEZ5CEEmMl9QZXaRVIH+0hXZX9LI7/s
5zorzvkq9Au81tkSMACzvIQE4XTlLTOf71cQ6P5YPUo56VmWq+MwOKRELTMYdcoqYX7m0guZnwo1
SqjBBpzgqge5KLpsp17qJjUlx3hjWSFuEDqX/Ja6VG8+AFvjPpSlMjfdnOc3Teqyfn7RqZz0k586
QUdqA/eCVds7OscZOb7ACKzO16xGYheQWYZx48nME0KHx57hdq9DS3xpYiIN/7XWPb32nWXW+3cz
35M9NPS3DKXqBXZ2poOS9ZMiqh/hsfOdOGIGIvlPr9mbppAFHadcNfnMApCHoBQE+NZatFHEAJQK
B0Qy4H3S6uupveO7zaWBdc8spvxHk0lA8ipzcjBeJegDH1/U7YCDq/XT6pw8x7Px0UJ3zKoCQc88
mOeoKXZt8PJTiX9SyDFq1Zj0o+O3ain92ebqBzIAkLQ/kjK/jr/zWBcedTaCshASlPOdqen7s/mX
8cQ2MoOw2vxefH6dxqFryHsvWr6lbKpiticdtgCbzAbL/Az/J5C3K2lXXGR8JCySrmkjgLGaJ9e0
ExF8NOHWu2+M87hemSSm/VteklUNaxICKM9i4C6e3y7Xcxnc+iLdjYQeIK5DxtAGqIPF0rGw+xLm
TGXNIwgZ2kyyzOIniYJ+YhsvVtw+116dsKb0Ih+gKUYuRCS8QCM5g+ELTkmz7gKbT9HRV0OftobL
fGlk+DRisjDKkYNp3RnrHp5fkc8L6d87GA/1Fu8TrT9TBwXS8MQmkSHb0P+6zRH+FhBKYcpcoqUz
/9QBCDb1KE99JwO7DYKAlNUdaI8hM0LsetB1MvjlXqA1GdljxfveGIW/enX68WJHzggozktXLDOK
DK+tu+3S8BepuW0FH6OAqWupDyZBTJCrSDb2bGuoJnC5XfO6GwC3x1dF2jt4XO8goAPf1MaWNbGi
vsaKZXB5tMCOVTE4ygSDXSvOQjWhDxiCw4zlkQyQRqIgJO9ZiD+WacqbcGBxcRRLRjk3C8EHchVb
H4hAoYJzV0veXQCd3M2mg0/HerkqDPAPhPH9Nij9aPy9BA6IZAny91Uswn5pL9zpDlhjLJJLhabo
W2UExZwhHFpp/Hvq9AN24PjpT+UJ1KandryDyzDwsFcIvzpY/RSzyn+F8eTA3+rB63Isz1Ax5/KK
uds1vIRkCvJmIrzpnbCBoHhxS3HaEPqlehvz2jKBmPYDyT7LVxR0+yc35DF0OO4ps68S9WAvHW8J
xcA1pWXAELB+K2xpg86KDP0HW0DrkQBJnuCDGtV09Bmidbq7TvtoSPgv+xWb16gOGnr/ixKZW2f9
Rxzb9+z/MTawFBTrSop+isewN/3uaAVEGG37TMvK0WVsoXPntxyFi1WZep9zNuTXhmdZCd4CJYek
22LgdJugr92BPgknAYx+O92GBiT04RYnaxJpCWdxyfmE4DXExEmYMpEduDzenziixuil84q9UEe6
gGxBwRG/i1yJP7/gX2C8Glt/8ZpVHDEro4bqjt4qmApCSqzy1TZuisvTf9O3271nf0bZ01wY6oEp
shznUFi17KLQxziQTtcY+DtF3LvW4Bs36XbuP6CeV2LkPR6bYozhfGI6FecNzYFar1Cm1D+3TXpJ
95XfpOH/7abY8DqFcKxNbLLquygk0Y0sE/80fLhsGVmhmOzZrnM0AS6i9p60Qlf+kE0FnEUDOTPb
06JBRnLsRzwbo7enaFc3z9Lo2ADNEHf2yO5dWOQTWSmGZ0sjKjSIroNQ2YnoBuYxmdt2PsX5jYaB
VJ7ki6dArasUYXzRzCjJ32q3nmY218uAyF/fhmOSYNunS2OuNc+N/oc365BDLsR9Y8I9xGlvGMcM
8l+S0+iEqGDdPXb8F6M19ahZXjyjlDjq+/vRK87bYE4HbW6/OBQSPZ9fAKr45PlsqHjPYHx2U6Tg
BMatddJfwPWalQs9U0a0Jt+nbBSVfB8T60yXKagws8yn49OTJs83Sxw/zBM5uJpGnPFxTLatk5fT
3nTMlzHNI9mMHdFCWKrtvhZw2BYW19F5k2JLYtooFbe5rY54+s2qoNV9njdbtTY4hkXPF+3qSNDt
yBIFOvS//9bhnAQ16URFjUnVm9e0DEMDdSngocBJaDjilcCvWO5h9AsQuyd7Zh5n65E2AUDjJjWG
+MQBsywz+xhF7xltk7hlYNXo25WOeoh6OwyusNS3b5dAXabUlANfZM8Q+2nXe67Hwpd2BzAK8vJ/
PNwDvGmDWwbXOw/KUxJmK/m5hdIDI9b2DCVB/Xnj1FcHx6YzmxT7GmnfEVIMccns/QLD5pmlzvsU
Yf/1RP/XkMraJ0pD4OD8VktYbJlXUwiSDk8331fkrhGF5SmoN4SGV7Om0bGgZFZbEW1+p5MtTGjy
mB3/KRe2KgEBm843ZOlj52KGdR1EXlagUiNcXjUDyDYrrLE9jYOjGgQx4ShalfErUb0L2Z73Muoe
efmNQo/ky+oAe0TXDR4nAjN2lxt6iKR8rSsYIZHMCYgrvKlYjZRYcLlOCkU8RaDBIH6vCZbHHZ65
yoP7FAuCP7mEszbwjVHSFMwlMLjshGeOYMFp7cIAtJS6ErpqMLdp1NSNMIld/PswnKMgTFkYioHK
qun6/eYi+lUII3QnHEh60RtBorhVcj2HutGdxxVre9+VMUeJ/kUFCcMN1htvg5ba8pnNsSvfyZes
XnDdJOuJ3XUtv0Riarmp8gmOwcUx3HqrZOwlkwEEvvqaZ8u+V9VQf1sjvRG0WfYDxx46y7LzF9XC
doCsa5mSZLIzF9a3lYzzpCxcOqDsQ1jOls55FqoVlThab9RBw6rTTyGlhQ7jtVAYf/F3ifHxvRk2
rd4z8C5EkG4i00c4WfIVCL4RIy5Xv46aupn9t+qLNXm6WH4RsTs6FUmmND4Bu9KIvCATofeBtbG7
KOZPiYdMgTRT2Oy9gcc7u2LvSkH+eqz+yBjIH6mW1oMMbiqWQF9qABE9aMh9pnTOnxTm8DLfhQ14
ZPLWp1gBDG/jUINJaQGbESqaqslZtojhgcp9MUHOyCTaG6vzpAbbfhZuMZIDo/KhQkJpFAlH0Akj
J+Mm4XCzwzpYknwupnw5I62kfJFnRFnBi8eAqczvCGAQaxgLC4c3sq/Vd2pgRE7Q9k/V7tUjFWBF
pjQCTqUYJ4QefZlfWqDTivOg+HCGd2KqtkOharJed7ovjAF61LpWUT4XgDjKaPhQ6g6R5tQsZ3B3
/3BEOZqudEFjvezle/btVeJabjOQCoKfdqnPlWWYhlM8s8jw8dRYnfzNOqCo6jcVquYuofSz1KbV
O/Hii8srP2q6FADVIeRtsQIKPAGxYLCBbPPAoAKAwplTxQfePbr5pqHVwdCNnZwqYStF1vFFwSV+
zJlpa2zsNqOldNajA1KbB16hHYw8d1F9F/HRloQxI7lWBEyQBez78F48SzW9coQ7Khce5CyH5Ij1
3aOghBC/p/e42kZ+rJTXlteU6JpAOqvzP0diALHQC++w64EBHBAgUlm4YqgUHA35CP1uIsGmMBpu
aBDhbAEILzMHwQ7GiYwfbfPzz4rV3MkrhdIGgjy9kjZ4STWLVvWm3htVPVvaFykuMjVaH9u55kYj
zJMB1t8pduzGGD9780KcBAwQoczYPA3DeKlQpjYj4wwwvRvFrShVkuxkLWHXorI4uiJvm1rHow0h
Saf26qAk4/+Qpwtqz1eLN1B74BW41VVpz+cUxibRET7VbMx+jx3pdUrlGK8goyKRs/qQy9jJL7hi
2oIgkvCSZ/oz+rUIe0qgw8JqtkaFttWA3AQthYv1d8If3j6sLsBeQl2jIE7PWc6N8JcQWWO36+i+
m++IrSxOSc71Dyz1BtUt+n/dOO66Deml4Yc2G7ei3Q2eOTKm9LJx5MkoLhlH4IudoEJtYzKIyhdk
tSEb4Ajir8rJLd7LzLUM1fteVJRvrS8gJCMZIOZPTgISNk/v92B+HmNKmyOsqZsl3T1D+q3eYMV5
niPUYX77JoccIqrrXdCMs7CZB0dnegTRK65EDd9GDnR1Bv2xq7QhUJnuGSLhJ1BHhFSg7A19SZfw
ENPz+h1UpyRv7S2WRV8gn6zAlywJYAug5J7GdnoOS7Up2arg7aIq7/GOC41FIJfk5YAy3uBtNb5g
my1+bYUo4slhe+VGGFoyh7mRDCPsG4twNjTjvoBu7tb5r0QLyNt0sn2jTw/fRLvJLT0vSifx5WEK
SmLs3ZXhu6XIWqGRh44qGhFXBHbxh95iptCm/H0uuYbOzchJ5mx28EDwT48M+xIo16Mtt2SW5Z1m
pY7sdzD8ym4/KnjlyE/aAeOiRcvkLEDN94DxqF8IE34f4bG56GrvUTg7X6OXtsRVLD+Xw+n84YH7
2dUuUaH4ctPNY/E1e68pjQlG99OPbOcoassr+xvHve+5jN/d45BmPGZiuUj1LNz1TCn0CL9W8ji2
dmOAW0H6a5+VItvvkOUxxj5cWWKhNmc9Wi/vA2El0ocYOb64erBgBpDxDS0jui3h/2oZKlu4IKFB
+It5ZpIjzRfhcJpqZ4yLUExtHlLedEb95ON1rxmEptsTTY5Lhv7E9x5OK/l+PZaBG+BDA4KFnUYq
dl6M8z2Yeml4ppXziVwzk6aZ6X5a9NQujLbRn35lJuJzvgan0oL6SOMd+Fw4hApdYOsHdHua8c0G
1MCIVELUm7TfyBJglAS6lX7C1nSnAjak80zt90s/8E6O0iLIYTX9oPGvOAcOMdw9BS0vJ160ugXh
j3yh9mVBNFWvchSKuY7o+0XHhGkZywFe4dIgoffQvLvXTG63z4zka8s6BPn5YMpdnzbhPxx7YTKZ
piODWBn/r/HvSGEluxO9upXaMH3hFUIQzRU4OgMdQ/aKju/81aHQMWPZUj9Y12WysEYGwoAe+fQh
nMoUyHd2ayu8/ufuB806Nv4YEqdIDENz5bYi9OcLibKl6XKEpJuo+X8ITHB9DAd8glpONRDKQiwr
Gug4UQz6JefHUxYHBg/pQk0+b/JVWyJAxUcDHZydV+w0pTG/YB0aPIbpbNwFq0KkD42J+RQ7fFN9
Hp0aEorktf4jq3udvylWHXA2HewoxulwV6O29hp6VKojyoJ/A7lvE6V9WxYERUJwktrCiSzYBVUx
+vC6VmRa47QOCuJRZb6DrU5mKUSHaca5avQjplILw+fS8QLm4eZvX2J040n+VFTx5E7EsHpqWCdE
ylptzJ3qS/XZdXhlyocQAVXqe2QGv0ytnsr0wkb4syZDOySkI9w+Ye6x6k74aLsYR//KtQ8bOaNz
OGrO9Jlg5RvtHfqOjBaF+TouDGPZ4udwO3MYw9ssv5fPLgGMhLw6hLppUiGPQ7JMKdLpYXWAixjl
rvpSSDrccX3AZE2v8fmQmILRR2GamYF1G9OUfuc+guYV69P+J4AnJkDKo8JwIryvA29rept4GLhN
RojwE8N4TRk7eVcHLpB/bl3i6bYrXWqsdyV89EYD3L98ixof8PoDtwfA3x9KYgD1v990pcD1zCBJ
CrC3QHv4lHW60CBnqBLaa7uEUOMtxyn7feLluj4I7jVQUZgu5MyQmyEVMqfgf4o5HHkjqFJkzbbI
oGiTAn0Kht8jv2h3e4QA2yID70PUGi3pNPybugR7+6MLIGAqEwAHP5dj03t7m4dB+fT/ZdGDhPJz
wsMsk/WAI1RuEXoMZp04Abu9e9J2CjiN2iGFChHrp7ybk60kVT6DX4gVybUHTO7NZ4kc3m4bGWRM
oup2MoIaJVeAvnISGvxG1l304vpQCw2izMyU5Qk93JGlgwkdFhW5Et9judRPYkb2oTcPOqjv2hoC
qJMXz5PLTF2l9oUlq2MK7A8wKWYoBqVxprmXYbzZoBffnhD7xQCLIfNLnetioaW9GShrjAUXYQuu
NEGTCgehzthCNh1tMATsuQrqc+1OkyC7mqf0RRON44TuvfCK9S35G+htOLrtS8Dc+MIHLrJIzW5O
HgbiJzWmgeo5WX41YzUbsXw/0v6HZIBSUd5M0vlGChwjpY5IGfhzpI/7PvrE1dAN//To1StzJ+i+
06LK43kEqP9aCheyrXAIXTCOrgA4f1u1N09G92/0P0vjZn9bo34iJBC/rpbWaP6Uc+AGmjPVL8eH
mFwhuI1DaYKDNqLOiveAQJEecK0Ttng/YgHnrAFY49sraLDJ3KKrmQo0EQi657ChjadY4ClHTc0i
NObLOuhF8fYjiuXB9JETJO/p82d8MTtkg6A4FLYfTZqXThBJbu/u7k/TObut3pfjMsdfPZJDMXMe
y+d/eUq/e2obKlxE7N46Upk2dnXFWHayI1wTvd6HZUEDb/VqwUcnANw87C4+bKhU2l9dApzx0OYz
Yx1YW0CpuNkLEJhVYwu/TRDJcHGSLrKo9uqN46WjLhnQ/hZVJyawS8QKrprchOvFtwDGLpHQdXU1
mP/zv8uJir0emhCkA7XDwtZhsJz09sEShttDVe1nBURO3fzyFKj1102DyIQ2Y74+XlppMUnRhWTY
nyiO6KYXfGV4PZ/rX+Eq6iO3yGCgG7QM9K63eb/q/Tat9JFWEKVSnFcAy5wJgmf3XpP6uCSyO7yl
Bkd7WDaptzuKs32KfN0PqhRlo4k/OuGpYM/JFyRGSP6UYhXZqkHcZ9vsV/4qXHfwOS8muIBzf3HI
eL/1fxSWbmMKEfmW2Tv3TNEyBJmEsCt8Cvjw8lsYVc0fLtsoZm65CtGtAJhDFMmzUvBOaqHkcyjl
FGgrEiZklcZpvovT6xFzzspUByRA+KBjj7IxXAn7vRvqOCHrvs0GtVG4bOWqQqFwCu7oWQa7b9PW
5nNFnoVTX5XXfwD1Tmm4e6kDsvDmbsy8nDOZodhmitLApSn1LGPgQx2dkipcnfd/L8ir+pB53uv4
+lCl2JZu/EZo5Aa/+PDio2EL+NO8ga9i0zGFTlsq2LpecTYqcQKtf+g1CFO9SeG6CIl1vmrtKYZJ
7UrUzOqYDn6yNUFzYKAWfxSGst0V6wQ5UKv9xDKjf+77UCFXRhd7zc8rCNgwx8wGl7KDaQcpDE8C
/8tC6QFl51R2yCJkcfuTS6AKiiG5Bi1RyUTaTf2N9BkIy1+ODAOd0+Iji100GC/P6fJideo5lsRH
r7FNyYWC7DI70qYK6Q6NBDnjEf2Nai/2eaSLFLFRwX3xNm3FX5N4ZpQ78Wi21t5Uq5BGw4/NajF6
O1eFE+1aBxdMsstGUM/8e3YIZaNToiBbp4NHHYuSpDxsLhEeCE9+GPij/GEpY1cOC9OfOAYrX7Tl
oQxt+sNemFWAnIAXIEL5z6ZFBXMsy8fSD6iSGI39DtxW52QOThXjQDaajR5TM67TlpL7yVWJ1vvg
dTYxTzVDCNFbvP1+8gvscPZVd5km0P9RuUrCv+YHXC/mAmvzOdQbV+DvUOEJUILVrmdaEJif/Rnh
mO9QHgGl65rO5GxISTQEUhhdHkFkYSB2HwX6EmymdjoS3VjmTuqnObJRSPvF/VGe109sUJwH1OR1
UQxZUM8gxWLxpE9E6FfzumUsldYl8vXfPwTQGrRgBsrPyc0tlpzh+yXS4QR40/mp5VpkrzoNES7t
yg597fZn3XkgNwBmWXpm7CGiREm9XGqXc2I6QAAyzSLlzHHOsptyYwMalgEhnHAmiaVOtJ/leCT7
TZ1z8yDNrfdn27ItZVDAirjgUAotWQ+060I6inS/Af6xZQYdoBGfJJ82BMCCWu/IwUu90iYGmIa5
Tq19uywu88u/pnA67LZiYtKda8RveAhnAIY1u7fc81FP5/GDbm0UlUgusLwKbu8LMpSw2N39zQN9
ezFAuXmpMvVLEP+ePuTDuct1uVWc0U0xbQxhCNATWpsOmICIL+/Ipt4T+l4Pp0T/hdn9ZNxqSwNx
hyx6P/BHf0LFscnP1HBZtS016V+M4eET5COiebh3vhNakKPNJcE9lmRZr9CQQKqoHEkjtn6RVQlP
ZY3AuFgsYLIgG6eHUERXfbhRl0N+xTIEovIEeuYQPKuxBzZjP5SfcYK1mmGKp27B9SdL8HOLALv2
ZnhsmAOqSJVaUJ08Huts+mDeMnA9qCvNXdpJciVfFpjI6OxBoLuAMLvso7qnloZcGwkoTR3Lap9A
B4NU4O8fyofZX91/Qbf4VGsbYReJLqJ6mO55f/U34/h7a6lGn2aWYb4vR/R74k3a2aOUZma+291g
cVHcc6ofSq5PVlvTtXbDHMvCzxOMvWDfZEUxERXDsAI/OY6B+yKPXkUOyn0fwI2PYXOp7VS/+ydq
ISYXl55KRbg/NgQS8RSeCiU8zKT/bV8KVrC5D28tfnS6GXltvqt7VQsJvBgfhiEhaM/01Y0Yqww8
vZI/AndISwD53/2DkAS4EwEgJENLlabV+uR0jQ7DcdidfFa6DRbPbzD6lkF1bD6WQE2UsiRoahyC
srfrWHWZfLx8zHsIBbOGI5xlzy3LLwMVUpEI6wJzWpurYKmM8c7C+tKqOCHTlv5YapJDS387f4FR
aBrOqDJ1XjjcJ1L/ht/8E5gThHR61/tO4uucGhBOgGy6G1eh4s02YPLvS7aHicp2U13Q5P+2hbds
ueToBVls0r7cIFUTutvfXuM9wm7n/B5dtZltJGMCdEVA4dPeusDmLyLHkM9mJGlp4MbhI/pYa8hU
6jzvDVTXjIiJ9aOIwS9MZ/SurvcBAJTyzhI13FPBi9Io/uc0Q/xS7f+Hvnqn6zAnLGtEvmyt7588
dv+KtA8ZaQmDuIhmq9x45043GZB8sCkoYPvFPyuwKHaTam5269aKyGWKydF25dGmEqdlnfXgPtrk
rEusOILgU3PIrTiyk+3RNuxpIrm7vBnKqWqju/gGFPCll+nsdaqQZRP5KSFtEuDsPOaNC3TGy1tl
EAta3ce4uKvfzz/FllMeeG6Xa94ok5p+eSHIP6kkfY4cYpkfvh1g7NUHMCzB+vuEgZBM1/7I76FE
HjX/rqNOMFyBGBOj60MaU4C4yhObfs7Segla/QilJOQrmB/l6UV6hXKnE7ZM7nNk83X/t/b4Xb1q
MCeJsQqMQkqqRLxiLnDls0ygL+0BDVYpAomZkc/cMfTx/EsVI7Cqm2gts5VgIEko5ddOgk1y/ViE
yvxCUoLRLaLFtlvTwQsLKHwiz+BMLGP3KApkuKnaEh76D0LyjfeSY03kZ4wJ+4QbN+LBjqsr4ojj
1MiGdkyMEMkx4d41G2vx4gLdzDwXaV8o8G8sdlvVZpwRGzeQUFU4zK22OvWxAhpDcBRAQA0yOaWZ
92FIRnTDNpqJGIEtfgAjDrzcV0kea74++yRSjlTRxIfqX5IIsUFqWMbsq3xTMZ3c5/Z0HSL5dZ9U
+4rYJrDwk1m01BzVOAOR3G48G9pDByMkeAIlCAniGiFNfF+66HKx1D7y8kjJ3qOFIiYnavpOYU7w
ZzwA6pX36OCdSYVVNm/s1kJlSI7jq247dPB0yJX6NV2mxsXdRRUUDAkrFhPcJ7I+Uwzvr7WeolqD
9vXP4VWa8Mj+ylCSZ9E303byWg1LLci8T5ILydvT6/73wdf9Fil7/e0NyIKzJUMaOqa/v290reZI
5qd7XXJOuODn5ZnimY1fyG+ULqsSuHGDLJmGrC5XrV9pDRrpb9u5bvTDWo1jvRUGBBxAt10boe88
teTrq0OT7iLJC9TukKRCvE1h2h3t+SocwRAkU5rtcVknYc4GbkQyYzW89PZ+2XjLxVEM6HNYl/7S
riWJfDJayEqwFYOEUtE8PsEPQu53RnETBBOm4Hx7hbWW6RG6F24Lp5wLhC2ARst5pCeZLtDEjBX1
Tqk/f1cUS6aRXyETYUaaMs62G6h37ZC+jH3iqBQX78+UN7YlMh4fW2iKsCC1te8CMdvesx5if238
wrd4mO8oAo3oMvyMZ0JV8UMXUs/9ZDeuyFmGXWRUpDpYSGxN3wvnV54OPLWX/0XjefMevIHHZdOV
e1VG/E3k30SNSeKcYmprnD5hESF04crl9AMqhD8e/SrZIWWP3pLmiDQ/1buWXccktHgtqLKThC+q
BDm/++6UZpZjjsOqmYx1y6j4LfnFKlCLGEY97a4Mcx+RIZuNFrYQbQxk0D1Nnhfss2W5eyF02WxM
37RTZUmaGPlEP7RSkAcJJyu8DvQ3hMCZZvg4Rljayk2gKvA3sJZI41DXbIzSh/f+u3yy3SRIseXm
QNlp456ikehLO0Rh63WcTlIQotKO8l3fGswzttt1Lyqi03qBIm646NJNIf/8OnKSF6zVudR6elm8
Zcak4xRklf0MYwOJNSgJhwA/1bydV4YuJxBtTkZfiyBzdsjhN9fivPJJL7wcuNc4pJ2F/ympC01B
ZfZkDUjMw1zusJ+y+sbAub+j1sDnlWHHc59HU2iFAjpJT9AnMI32KQ0pgd1J7cIWNtJHMZsco66J
G+Vwm5pnnUURrEppikgpFM/5tbA8mtaiF0bDrMSadSoxc21FgNJ6EYE6ozNoCPni5TQO22FPdRCB
+svNCJ/ZOn333sdZs5CsMFcqAjTMbi/gHAaK7Dsjq/+yJGgvvVqScC3z747oTDHrPvkJcd2F/cvn
FavOri3saoBgi6dRbri2Pq5JCjKk7ovQaazR0EOahV99BdaeaOf/g5I/qV80diraR4X7l/QwlDBJ
+CtEoVbOnQp9ESK2ysSfCTiXR0RPLBiYNHyDqCWhxItxXb5ZFX7zOwsl5bUW3S0b+v2aGp4TLVX8
FuGHh/vGl2dSow4kF61ipxu4XCjsAmWT9Cw27VuUc7n9OhuhAxQDd/1jDxJNfO/0D6sZdRKsQqQg
JNVALdtvSxFwRkUUhpE4ouWmywH+aUregx92tyUnaREzfCbC7Ql6r3uIwDQcA57qdJUX8cRKVWcp
wKdC3p0oYHaWOoQhy2sZNv13OTQGUsj9yhqTYrg3DyNYsYW3EqUgE9GUbjVTkvU+iW3Dd0libCPj
NR5mL7nw9z5oLit9HGwQS+KvA6/M7L79skyLVL4XhOuysWh3B6YWLCGxHvY56ufecwDA2u/UaTNg
u1VNsL9XZEXld6JXF1EfxlKqXijYGOInVYxjjH5wfGxpq6wDIeLmk3kiR9nGjXZ3ienN2DBaU6m5
ppwErVEAY8PPb4eB41VPSyJRqbtAghoZxbd1XpUkMipTRB376rsLPII4keZmHQZhr7nH6Ko2Q/ps
mL62PgIcZeeWugMzPd7i04E/twlXz8Kak9W8QAtleZypuJYBo2gaKIAV5oz5YKTIzxlk2rv9Sxk8
+yvqXhCtL4XYz3yugZTAuwKGiXU3JSSxVbhGRTQKKgb/pPHZuPm1Jj6xFGyXVxi3imx/ktm0cqwo
ii7sHfm2XIFeQoAZ4jgAYikOYWmxJlPwB/mmyFX2ABbLFLwPnpfzGylQOG0LCtcGlEX+aPjKT2vK
GjKmSA1ago3prSEfZAdUIfgJW5Z9KI7BDrbdwW0obNtLsRxJMICijPNpLta+C6mBFWlp1zxkx6jN
pdo4LhUXFQtlRhZRHTlIOKDzhcgK+pBSctpBXnULsLI5F6UuslXEHIOqwMNcRbNS5JWZZIiZaddt
Y57BiOMjL8JcVtYIaKfFatN/jgDPE1xClAiGjKifeh6U/X+BooUC83zgiosULjoA3Vwxe2AhHA+9
iEntbI9V2tj2PwN+JHjaQPL4WX9J2BXxr9Qfs9auAsks/qc86fMlCAVUZa+BGGks0W1gn9+hZVYp
cVwEGXFqpR8tk3UzGZM3/Sx6Zm4GSljWNwRWNyaxXuCt2jPMS7S88eyrUWQovsUo2Yd/XUhU1PzV
eIbQuduAdJHdi7vUwWr/z6tZ1VE8v6U4Ojjad8oowFEjj9vMkl44dcGmLZ7Tr+XciUaEieD0kHKV
3RDt1FShffLRvjokr8tqNsxJxNLCX9MXkdMstulHEHfAm9tVyX2ivrYRjLCS6J2sB0fkjY9iBCOx
D2+PvbErfYAK0fJKLj28Subhcuc42ktc3JJ1QjR5+IYL4zcUfjt4V5E3UqM/4FqJ73Jqzyzs45s4
7CPLBhonvyUd+Meb99ogSAVaH3MpWGnOGO5twja4xj+zmcpLx7avrrBv/nd8hMMrrl4m1n1Fsk03
VYCKEeH9JZc+sR2lN5RBnM/1w5VGqyzfSl58JLRqxEkWttRwwLoplQ1JwwMOmgc/FHuKuTWRNluA
faTFv05ZqwtAq7hl/Xl1eqzubudgOPLRCgM7zsS2fWtnA4Y6Z9mUwb7zqkbkl5n0traA7HxrFjd6
3SMc4mc39AIO1Pa5TMNWVHNDJPIbdVbvvaNcLZd+XXpdzY2n7CbuMrXdNUN0WwwDEhl93ab1p1Q9
8H3KyKILjX8mwoWN5ps9bofq8u7/wbTCo9dY8pEOybNRJMt9A4WjXl33eBNf+pIAgzE9AA8y8syl
XhR0WoWUMovpkFidj6PVG+ocquI4qy91J7uCaEKu2FXezhTmmT9wyPuk7Yz5I6N7yPv1rngJaCpL
rgJcNjSQQUS3ACl2LTwUWIz8krmBV27lil72+4MdYKr1sjaDbxw81YY+AbndUbgDRrVH+0NbEE+9
DfbFQgWhBT1+/k49dQ/Ab3cNgWnQr/2yGmCsuwAWr2ja2hqkB+h31cpiUfeRufBSijn0wITBemqP
dEt2N90ip85CgakNE+8nFZ1rPB0+kN4sFiKQxzhbuFI1q/YfVOP3giCyoXVymvq5I/j6jZHuYXUq
LFrAwLJxUyoNJnyGv2n7idUPqtI35RPPq+3BQ/eFlBzcxyJU0ylW8YzueXSBSrNRTxtJqg2exLUO
eT0RH0taIh2en9sCt7txQFizN76XxjdK4X4vgjH3NUbsfkOD/7653Mv0dv7IGrS4WbWZ9lFXeYqL
9bPSgjYvK8HrSXuYwn4wk3+b1JmPYTwnRRaF1bpnaQASbv2k/fY3tQCO2gbcBCCKw+JGeHZ70yMz
BAA5sf8pS7XsX5t1N3T/chn54kXoOCTzRkJm9XCjB+hbT5HUVMqxDt4wtmqf6wbmvRM1h2woIJMa
p9C6m3moyK82MPOk5ABXFzTJVsG/xZUxWzeBik6fqvpcUfmtN4qFEfZfC5dCbBflSWAAFH6Fx/Zz
fsMjIxiy2QgCmg8O2jRmvZM29AiLUHBVUzmuKpAIEgv65A8NX8/G38Hx91PvQoiKAM8XRFVcJm6C
4vSPaCQCp2UF/4pPaqskv/cG8PNA3cjcZc4rk4OcIFuEJjKrtqP72QShgrY87H82ciZvK+2Hv1dk
9Jgp1fnYoKwEBli/0xFzfIVZr0RQelAQsFksfAxZ2bRbKeeOkzw5bAYo9D1hc+XMYuQS7mu3DY2t
gMlWG6dip5nJY/drh1srSnEAkb+7bIoqWQsYdBG9vUbdijuSRQm7HdRRLhbdKoB7VDzzk9qS5GOM
LOjm7wAOpo2bWIq8haIvrk0zwi6aJCQMM9OVUAkptbHu5V20WBQV9yDweyRm7oV+MSyUvNaegLHi
A3t9wldZaDUkvDvA7zYPJOLiNwiFEG2AczJPa4hLcwrjQIVBiSY7W4kOq0FGfsq39vcL6UDsx3bL
Fkwytdq51Q1VGQaWRcmwUuP1SVlbkLCXFGPFx7FtoYmFTM3HZo7fObMdr4gcl30lNHZyGGH6su0u
ZDZdXZBQoJ9ZEyAGiAs8Zynb/2F8m1lXJ3idRXu6ANkYQkb/iHjCVuk7GQjZ2uzSyE6q17iXrlqz
s29ErMoMnFCokt33HnLcnVpFNwdhsdVf8zqOHL0gZFzByHnN7lrDLnaemotUIQK2GVJc0nolZ1Oe
oEwLauYmPZlBtWCf6sAJxzBFkeyJzfQxvjPHnpRfgnIlJ80yFnsOJLFPIBL03hkUnKWbmCGlG+wi
JYx1cLXAJuqLC6SZerlC6xZz+8VEGx768DIQjzG9/Zq7appoKXup8QOf1joD4YTgySER9FuEbFtv
/9t5Rb9HOI/Nw4ByqFKjvxRBMCmewcovYL8bw9rteoMnKJ/pC6rP4fr+kSvO8bjfuc3Wwo3qCBJt
F4BbRZpgvWUgN2Gdgi/G9DXflsTph5Hj1K8P2FyiaWkn34o5XUOOmrQOQNHi8lCmS9ILKnqHnJXk
zJHawWvG2H8JaS7ywL2eEAM1m4IXLohz67PdTCv72ia1Su/yeBMZIdBT+wJT+Lw+2v+4SOtaFyd+
kf7xhBP5fCY8zZ8N+NS4KXozWyMiFiGbC1ET+YRsqw/MZ/1ZJDVYNgw9Xm4mt6Yu1n2mwYU+C8W0
BSCokvmlI7bidZ76e+jhsOGmYSm05yISUTQl3BDpYVqtnVEd9+5sVrEG1spidNT+d/QVO6eqA8wT
+DZMilQ7YD3R/iKZYZNTZhUYXepUespkY4/7bZAGBj3KFLjDd4N1sBTRgCZDqg1V9u0UlKfLUDyr
LpsOEKlReFHzRn4GhryExc5xS4US74JtkNvTO0VwtVQIjhkPZ8bbNG1ADdB5T5XOKsHPH8g5HgN1
FHbRqLjXHEzB5uBYw7ytJO8WURkeL5hA7zoUZ9vOA5xvw6U+9IwzSFNH6zfIAwuVC+GuftEMMcBD
OijhFgkPHjwM3FYe9EuXpSJRORWm8qpCJHhGwUWC98QByTVljYGSmeVAfvOA7rYtsp/Wj0a/kBtF
AlfTFFw3YAS9Y+koj4SK+qMqxbsylaLqIFA3hvZ83yCTNZVaz7/B3/Sn8sNdO+nRL0QxFX5Ae2cM
jHIzJnau4CDDJNN0+EqHeici78KAfYtP7ELG9AFHvXadOrlHbTJS1dYKgigWfOY8WAuHpWLh8dxb
Snx6dys5zyC1Ih8hyb558cXhsAHZBXqFEZji75EgXpfiqspwPDaK21DEjMRvyiKXKz/kJ3qR1fuD
WVopCg7lmQ/6ME1mzMIBK3ld3ZP+uJn32KS3cLwnuCdh+Qh0yB5ET9ZKSs8aVVUaflQjEk/isyj5
ygVBXPmaw8irXGWYgkDyEdnNUIYHctLWktjNy59hle7eHFiODbXEXZLjqfvKG1bjFx5qldCXrmfe
979J1yieJeRNTlnoarhXfPdUxF09s2rhqCZ7krQR3+mslxVpw3gfT+NiWSFP1sv4pkXptZytekC5
RroCT1jLeAGpkcm3s3qVOniyU0NKk/uXijAP0l/8WYzdOQlYghImIikhCSQXZ2roxYgotrrs9zUd
8H7U6/fM2G7F9d2cPGi5hgzFExmelXUuB0Y8zec9kuScPrOSMHUy41BvvaqARNfIItMJIfNPp+Hm
8xgnj2iaq2CyqZQBKHvBwbPl0h3x6K7LUagn7MR9KyZyCijSjzI5801Fmo/ZT/mRtXVAdO6u7+Gv
bHWmNFpme5IMBgbBhM7laNU3Gxe4rAPXHOOEKMESGlaqWd/0uxMgvoQgBkDi2gbVOdl6RGkU6M8D
JVz9B416xe20RxiPey7dJPETIIf+gllVRDXLmE1vSOBkVxshS8VsDOY1QsKjyaYeTLR8tYPrLcvC
71iKd/1ZczAZPUOuPWXyg9ozTES9BEyvYpqFrws88RDRYchKoBHgVWvxk8nd6016hXpxrrMB+EyQ
DzfHAf9l1r8Y5xW7eESrU0fxKI9bx35GPEftJ0DxjRtzBfC17xVCf4pJItrrJGCwn/JDYhXtOeSY
QkoXWE3bZeB29cFF+paAXDYjkGawnOCkPIsMTYUc/ro7ak1RT6WK9vJ+FCPmPSUtLqf9xH1h4TCx
au+Z+rO/szqjoGaLLDElASuoEycMmnlwk3Zq3EvQSIm1DZheg6TU0oAP+IDMcL0TKSD9qU17J40X
ol7k1zBb8iQMB4ecKTWjxqBRz9/X2loCTWV2f9bm7cELF4z1SLtB0+6veFR99BDWymNvydhMoDf7
DQWhdxb/yiK5CPMMmskRhfP3VtiWHPBaTjTUEUkkIIUgEZbjtXTZytUsoaiQbgK7AXNOqvnfTkBa
pxdZHc+89AfqSyMPqEMnLX6GXP72y5y06y5WfgMLtHzRFAK7f9eqZQJT/kKFlZgJcj9m8E8NuqHi
VNb4eAXginRmFj1Lyc4fDZYDCEo8X+aEjCs4GxSL8c+WXMnu89zk05iGmwPecFvOgP2gFSx81+YJ
Dkd/3vuvmwvNt49QMgbidMfPBTwGuvjVgXe9/vewAJq3c4a9ES3Rsv6mc6EEBa6fI4Dzz0vIsON5
ufk5pXO4eJhxa/eaSKJiK0yYBCCcdhBYaWYLB2BGtP/IOrUx0cPEg7JcOHTfwAq66mmYoDZalM2D
uaRl238358I4ndgQxSLsv+4oDNWFb7tg8sBHBTxcO9AL7Q6JLZp0p3JGb7Ul+VlE+vGXaeeZ2YdM
+U+Rc301rIlGBV4XECyCy0AUT68Vg7vePIJX4d+89l7p6Oxe7KVPpLy1m5lTBG8CLz5prTSKCqfR
hDTXzCj3xH9WfjTxYIOt7pRCT56puwMYTGNtwJVYSrp9bFCUtg0O8f4qD9otgkiX8lrpgfLUwSeF
sOJ7TBlxa2JZu7quQtycX0/wvkg8Xov3ayo3jy6f4crkXi2ZQ9FTFvgYtgoQdxe7sOUKGfQZ4KuJ
R9taNK8IIAcIPt88dygSmD4/NGV7cnAefmPdn3Rz5ZmuW4MCSF9DrcgKD2JWpCWFtl7Evm2KR7tL
+4IfNUG3iTT97htE5WqefFnPLLx8bddsLI9GYgZZtCWz7VQnhw7Rup8O20hPUIlNtSOvyEvSJleA
3SMqBbb6mCwm4Vyx+nxyh5643inEqFj8COHNTmrpVGkcBa/iYZyh7tqaaVKMBG6jH9qI9b4lhusd
HosCHL8bylGOMjPRSZfBjwfuRl5xTcZES7bYyV/uJUXL44vJkGEeFjKAz2qP8K5Da7RHPnv67pkQ
4hlLiCKNJ4ZpD0qOZrhCN6nbJUJeA9e7kVjPSKUydzMUigb5sCY5ikb1HfkhgkUqdbPPS2EASZWs
0SpEJjQPJZKA+EdUzyUQMOF4aYjH45Ic5RLARyTj6fXBdqMJoU7RPIQQxKTRtVmKmts2o9k3K6G8
uTntHi3+G1TXHu4ZEGddDUbJ+VkRaoRNa48jlt0vxzYMqbwzMJmGxYNw59+CGoqNSkHtJZurYmw8
Z/kQKAKISbiLTJX8FwUCuXklh+sMUaILsiJldECJLQ1ct/lJ4DZ6tZfxQ582Vbkj5uh+b+4kYLaX
vS28elb6KvHKPOMhAAqCMu87bEHvogIKZoUDSYI/1D3kqFyRDmY/8Y812nIOWwjbaMIxrssaGCIf
ivW8PjvoQPbzZCGz+45KTSA123UrhTWVfO6MO4z95P13dDW2momfCHQ9cwM/7Nb+ncFNnD0INkLR
bhumrtwvXfPP3IeYVsQg820Iy2Ufr0iYR0sI0N/xAGu8QmQbnvPD3AeKLkB0poffY0yhuyVWLIPe
rz2BqZq42WsAQrYxt+wy87Q8k3qkRVVn7FnAV21GoYDA3+QaoimkljW27cHgOXASOZ2qABPD7Pfm
0pq+F908C8Fa6TPeMCgRj46zlIX4P+5PNcJefzeYD7y28f1lNC3/KKD/4DqfRFslUVzEUF1u0Rct
H99SchQ+crBuOtHIrIA4uK7yDbS1kstFXiWr628bhpupmiwlGdGY1nmPb+CO6TVXm4LVOmaQA7yR
fgZGiU3fgLEBHbLARc/41vPh8fciVCM8gKVhfsmC8VOAxsu+bZT9C/bAm4o3a6U3VG1QegpgRHf8
bAKUpy0vP8ZwxK1FL482LzJlZJuSE1W0m8oedlAD9WBiMqRFl8YCQ1vWpen+ua5O02GPTwt1Vk9n
bmtjN8Ptj5JHqD4RyNZoUlBePlXDxBefYUWU1R3Mte9ut7urRZcz++KRhPyhycU1sVN49EeAtblk
NRLQIbTOvg4Uyf65mYWxKf8zcjf6a8rDAqkXykXANF4DzL/xal7LOW6P7IvJ+NUqZwkCcCcZ/sTp
Vuv9bM18cA8hAICIJo/z3UfUI2dI43psgOiIjUUG4LpMkNtA7jQUOU6oOsxPRDci855bQGIW+oeq
R99nRb+xkZW5tzS+MKlT03kkBM+0QI3lL8o8t8SHSumhOCwscS/SUP5SrQZQ9rTFEZ7fYEQLISU3
uEwKZ0VF8Q0ZCoLMs+FhJSro3rKn4Eh0260Pgb4OGLsyX8NNgc6G05c6lOe5POmjt/7vLtspvG7Y
+FKopvkVtV1iQIhoBiEH5wQZGKAz0BrSct0+zGj3ynBEhTBxCTKcAEB5NQSLtKY2T+cjWlHwGHSl
CzVqOh6tnUkYGNXAwzFkk9iNMQl7LeScMWt/NkmMSIi/fTTi0uhsar7e/94BKc2qbZyTA5v8QydD
9JJx0lboQ7y/W1VZsj4BWOAzbSsZYkGceKlVreeRznhHf8iWhTLhASaYVspm2cvS5oDGSTpVKgeZ
KkNGtwUFt4UeSxa2KxkbUUAFngcUBObYmI73GM8/BWSXt30gipPmYYv7WSe8/WPE4udX97bbkLye
wo2mQl6cBRovzsk4YZfNukILbsJclNprZ4meQNcPot8QaXugij/t+gHMftN9d0qUMtRCK++zeFyx
/OmIfI3ps1gvGzt9ycqKW4GrxODvxl6r9pGfto8e/mdq1BzcZHLjazCJEZFji11Z1rb3j7+9xQzI
EGHNyCgvERCgVT9ydfSq7FQcqR6ufBNrX3xz/sJqIBxaBjbrN2GubPp46lZ0Q+493LGKNsxsmCDj
j5Eq1lN96GHXsHxVsOSg4k1JVlNhxOLfBF93fbsZu44davs2cdKQj/BY05kkxfPf0x2ie/KtrAFT
HKPlmGzkHz2yUnP+zSoGzqtRRvDzied8v8lpq+KEql/1Nyz4NQKkzuW+eG8Y0O/rgokN+qiDSMMi
9WCfvQikqouF94y5j38IkQucVNW4IohdmL7LMFYMtwE7Y8lAOfOlTlStwsAGanuilVS43E3WVn5W
j+IwwTSwR87SsQgW2BT6POgqe5WarunpiW+GtZ/c1+l1HSU9/TQSSJSchqCu81bcyIuvmyPXo3v1
xRVhaNB3Dkn06KN0X4jkrHBvHKJHQ2I0jPVwp+lHH3BPVqzX1yK+br4qcmEDA1kXZWMvKYK4r7LY
pxNC6jP3OoasZEtskgVWAmZIg70+nl2JNPyifo0e5yRbXSDVaL+Dkjjp4ULbwZELJCz/BcuZdErk
e6zLHEX34sfyYM8GB/2kGVF3MuSua4F8Ptig5emfLhTTu5BidpUqAXE/nJtgHm05XLIpKedrps9A
9Rcb2gSP7dC2Mz5DsK6QsJLQbS3um3kvEyM3lbObutQCvp5lgSzgykRpV6f9pp8SX/QbMdo0OJKx
70r7t1QM3Pq5dVFg7SHU3//UvjK+CXVQU+hNpdmmygHDmbUBKd9H50jYtslsiYiH4oy0UkpkK1Gu
BQEy1nfXgYTLIZdms+tAE61T90pXewsXX3tEMUTgNfBYC+nH75w06zdADiUWrAdnYyat/TPId9GR
x62QOzMh/wj3Z2hW/7Io0DkkwfNU0BzOvQKNmB9zy/ogD8hNyzapwjqhNP8QMb+RHOcSJe8SODxX
ASpvi63qYGg12t0KWvFnmU0t+SVicG+NAJJo0Ktu+4+zTRcnPSO7ZIDBLFPqRIz4alYHPgxkihFI
kYDeejtF3mCODu5p2p4T7M7ESx0QC7vT2y6ITREufEtvqKZOxA+fhcZsHjSZnL34sa+tdPgsL9hI
gRgLrTbgp65npgZi4STAegpiOwNTbT19WYbpyh+RwteUaU0S+127K5WTq6R9m6KZ62XFYXzULCmI
Pdxtsuj92jbLmEalNW3SrWzzxsxxLkxXv9SmRKDbwEyZuoUZV9uBKCI2VBVccPMfWvTrxmxKFifR
8rv1YbifRmyP/ZVlNvBdIfnXP7Av3uYnnT60pQ0T6kEACq+RG1NYlbia3p1O/sqL/QEfDXlldeA6
swdG7NppXIQwLLmcwrOzeJeUCMbqieEpNUIXHgJHdqKVr2BGyPJKQWgGnzMbIz4BRkE4rktO7Ml8
+pTLAN6GPwU13c6zF1g/73Tz5GYZecxjutmuI54JZBcTmSzmyFGO69kS5PSAf55+WZBKY9q/oy03
DID/17tAXQ/DMBmH+uiT5zkTbPD/UB0MvUd5z23s1iHNVpsR91yimaOX1IcLWBA6OHCc1B6VSaFr
Qxmgr2MJjp1uySrmGmcHww7gE+w9ehVS/TSX7HBur51IGEdZaLb5L2bMjYQhz+Hz3Bf+riqaxQ77
jiWZExGtaqmJqSxA4wD3sFwBQ2Eina1SeRb7iHqGWQQYdsS4SBrT1kA33MveIZXqCXrVfFP+MJwA
ks2vewIAnZDdw5LyBWZoLewkzdQF/V+wAGWUSstt9qXHc+G+5ohIK5x5GrbUl96dP/pK+z4XqmLY
MUX8p/p9//H7jTlm2Jb5TH0Qex5MS4zTHx1ilwr8KJiOEreeGW1Tkg8I12CSIBylISoBInqaxhVJ
GPC7V9/LJDMG7XCjb0GAgEQtFzceX2Xk+OZCO6Ji8bOjUpjVQ2ww3EEj5b8wiw6GOgMQANPxtRBe
G+c9jXcx9k0vPZvwOt9K7mmjc92KWPD8KSirWy/tnklI4ssNNB1YMmH4Wm7Q/yGLC1FtfsGc8YbA
INr2gbXlz87JjZUm4HzqfYbG7jWwLf9S75LdnH59Bf1Q+tHyLrWNnmAGu92qoh0Bet//XuPc1JjZ
fqprJ8dikksyGFxOG0hvAf+WLBqpdFp7dUdkcWo9ojEu/q9t5r/huaIRutSoDRzxswGTf849Snro
YCoDlrDwYkzLiyqtNM0KBtLNYc6HaSLD83nSdwqOWh/02Ox6aaLDOKJEPTgGPmtvl9cujdFuui6/
XZNzilQrmdlOpAeo0utEdNX2ZV1a83i9GoHx2TujILKtqyVs21CDclZxn56YodnhFM1pAwqrzcM5
7K+KjaTXDC1bCbKOrYa4gR47lnCcFl3+IvI466vPYc2LBS9i7kNlvlgnVIrZWg09t5UEwJg42/lY
mPjEyT91XY0AAsHHewaDb8j6ZKm7b7uxmfQkQb9TM7WnU8muSSU1ITZIJRjfPn7525uFBK9rTVpr
3EUc+weUlwgcGmxXNKahxIYFCv0BP9CYh0cF0o6rN0Rx1XeR5/ZBwZm1EdcHeP3APAxMGxcpS7QI
lKgHcKIPoL4E7x3+V5eO5Ea1oRf9IJIHXOGJ2Mxpu1WQ0qjDJ+jT6fkzM88IvdQEuXe/2j6/JUb/
2F6qGmDFfXwBkSj4292K9WQ5dzvZQNHx9qUoh1igEHZUFC7hGbTV2s4kB5B6Mw9l7I2Nn6RGucBV
UDe8aXCCVKG0MwhY49muElzU1caowDIV0YrQsP/uWimziPd8tv0VcLvf5hSEp2Y28MEcjeMmDhcH
4KCJfuwu06s/Jwewoa1znjF6/ZkOQNl2E9VP2nOq99B5mmuos65m0ivUh3hnSHbkD1xSBUBPX8Nf
1egCv87lJEteKZ5OP0QnnS8P8ok8PNV3mVoTHoebcisYXUdeqeLIhXumt+VdLNukNyEUULC3ug0y
MkvYLp+a42IGreYAowcqJxjIyp9O9tvAtx6mpjQOKH/588fRuZ54nG8qU1MJ/gyrbYNSCM5k/Sp6
la9/zEJz/XhjV0KhmBNeGUPdcr8uGdTjSAxpJ5T16tTPPIR8XoivGGdhbR6aOot+2Wo96WUaLUva
tOKs1YhqfRbFF3iu8ngCNQum+UBlJ298Wh9kdr1F0q1bz9FYfDXWjPfM9AscFoE1qDlcovoDtxB4
HzQkqVPhVZPTEe2cDZpZrk2vM5rFImGbrSzt5G2lzFXJ+rxVWo9jA4SYnPjsjh6rPkG23Y60vF9p
Sxn0mJ6cdZQOnSiAGtSdcFGZUZjUtrw2xjnYmEo62CBTzKrbcgcWpChrnMorNkJzBBg4FOfNsMpb
6qhB5TerIRLJtMeprE/2w0hUO6v2zP7m+fpa5cGHHCi+4xiJBatmWGsWBQNej8vqRJTGVAvfWm7m
/VPBF1kj2N92Yws5oHCa2Z8c1jFzSpt4jous+5mbs8tutt+JJ9cJtaCSMeGQCOVfUS3HQpx9rblQ
VD0f2BF6nU9Fupu7XHla3vxBX5dymLmV8b0fA/OG0ElsmN5Ci5r3xBvS8+dG9XSA2OiXGtuYeKjx
1KXrmIEu/SUSivm9K/KoyliUnqeJbrQARQ88lOD5ylc4AMkJjHHAm/bMI+kkUZuor4act7ObTZVz
++BXCBAKIHoavd7KuitCXt7L+Aez/0KsjM5XnNtlu9cwHbsAcq4ut76j04g1djAkWA3Q5USk2Brx
cMR18MMpPJACUrZkohVJ6n54Qai/SO0e58sUw/w0fnR6C1bGrVJ/LGPp4e7QKRIZ58yMRNNWewE5
QmYeIdlC4WdQ8FzWoBURMmNF9qM+XlvV/6kIu9kuIQf0ygVj4ji2rk6fcaZ68IpisxjyQ23t70B1
xPWKraTCin0KWEWGlcEtm2EQnv+HwgkYyWqzXEgUMbicHixjwql2cR36U1C5GVxwzCFLIQQMBfCt
DmFBUBPdy8qVJqF8DupvQVEavYSPW0ja0rluLdPP7eAx4S59gIfKBLwHvun2HTx+1ElFlfwDKhsX
4FqofVRV7yXwKzMlTw1/Hn8sBsWi7PINGvRXkuStAYNUPNOcbf02kotcTrXAGh6kTHhORdI/P+3h
CPGZ+bMkoPHeb8BmEbZGPrGG63luFVoE2y79PUOxOB4YCQH5SLa+cZtP6Gu5HxYH2DCNOL/OC6t/
UIdUDSxw9WEdErguzExoJltIX9PRPBuKjrd8Ww3nDpE/rSCYMDIuNPp05lDaNYlkz5sLoAETQ4CM
FNd9DJ9Tlc2GDlq6THYWRSvdk0R13FM7G0gPLrNs3Fa8vsq7agCAaQuNRlqg0JtlbKDRu48POt3W
WD5csu0mUS9+MHeQDqhSNUMVOP3i9TTh/7inmlAUBg/fnK9UAjQKn0hrZpXTzN4wnbWZd5X9sCFT
FYJWHUZMjkpiql9kHHYe7yMCFDgB/l/JAUGnE/kG0pWc7AVqNO5zpOm9PJqSnCcvQyIsSz51cTkH
F8fLOjm1FH1SaBhKsYZDbpJsSRZFkISAzR4qJhtgyYsiEx8MIYe7+G5YGHd84qlmby2vY4acvAiF
KrDxleW0vPcRUiu0BXzgx18/FsthkyFtqm64kkpIbZDlAyLOuqg961t7FnMVQCUwunjvFg/3EhxQ
JcqEzNgAbG6X5OmsWl6k0jseHqv4XTr5+0Ya5xIbRaUXE07dRFOKpHTHjLP12Tr8QbOcbonjtlCA
PNaFXpoSNQqajweC/ktlFQLIWQ6R8ujY5bmBWo81CSIupcpNhjkBH5C/XHHpwhWqu84U/LwPhhsC
9YVy+8TEGqD+vR2ozUbqyRnQHy+bRV5RLROR6zBrttk1LAs/tGsIekwnKedWk5FP2SnctNUOstNW
+MW5iU4dpV69ZrkpnRe0jEMCOT5JezOLfrgweNd3197mZ8Zw4+LNOTOSDr9n46vV1zf9le1mVwPh
v9qnEofYeGXcmi8KQWoQmgX4pK6eRY5BY8phRUlQ+lBqyBwqXUy18A2b7/viMYBDUCjg0joeV5wm
F+a8ZXozmmkJKNPFDi0sFDMzlQKtLYePl5Yu/ea7EU9zE4kXmUZewGX/1YJuDu+APIqpv6slEud9
QDBCkShSY9WYd8Imh0ERndVuUL5Q7VgWBMuCzrPZAhKJ1/Zc2nWtqx69We8fZ9/u7LURyPW/xCa6
64OK/ROfkZRY9tNWtpKbxMOxCwyljtyA0HGxDQM4Lc4O7pyexQbvgcWKCBqK/lTFO3NqCWW9487/
S6eIUVtQwXTCGWplKHUdZVei0Jc1DIdNZu/t2WJTRt7ez90oDU+6eOietavJhg3JpH9SofOdAcfu
2SfvX10DHKTZQboaHCqZKqPuJB5b2UMd2lQnQqpm2HPxGifV8r9+KueD1YgwmvfTLLUorhvfbyFT
B0kxOCtWGRp6M2aVIMvFJ7YNTJoedRCtMOrgN6j4sxTWX2NFK3aQilcG6vGN5lAUN8BIr1GnzKd9
DeXRoBklVBBiart6wtHXN7PcJ7JVMWu4CStMi3N3ANUrPdxPZ3Q8Q8BgwjDD7rOtu1Q6Hbvf9g0h
RCT1LSp634pHktCIZQS2Ge2QaD/iAtUwIRYEq50dlW0BXwO31nrYZiVjeYgoakkh2ke4aPH+Xi7g
abbELqNVYUDN1BW4pysVh1iO8qEqoEtr6wIfYCmRFVZMFqZZDk2o/Nh/R20RZxn+sITdeyBullJZ
jsgbY0qwXASSNUAu/OTZaXQnqjnaErx1VMdYggZJgW8CY40TYQjaw/aFkDBPdxI43O6ypPs3nNQ/
fiwMWQNYRngHdo/72cC1LOPwB+1QTiix6Q8TzPqzcw/wxYZxgrJzHq3Fl5L2qRmrPXa+Rk6NFzh1
d9OkRKJ57oycSxDWpR4rMiOZOJnatoK3GaV8xMNMG63+LsN0YyclSHd14FzB2J8vvF+4wmLO8qlz
3BJnSzwlSrTYr1PA6aKXMWkiPPOrLq+eWokirUgw3Z5QBwu6H3SkrkJJCyliUyJBdIR8J5wH3cZV
K+5Jj9TKIKB1SZkiYByqQxcTiUtB8X93QKGrwzQ32m0vlulL7jHyAmUqBjSyD8+4blH8uZ1eYrSd
qVITEwTCkcwsh0ZnJmTSoebfyVmvomYFl8C1VeHH3y7fH4rEnKp9R2Do7K+xbxuA5azJ/EWa9npm
+hwrOiv4VOxaSLocUznJv0+OO4oGw+v6Oq3rLM7mYKIFOihY4VjPgoSsPkMubY55PrpiYN4TnMhq
55hQi2BcppBxK9tngqD3mpdw1Vfsz6DTdN/GRJbz2r1l/cB3y4+4Jke6r3LHbLVLas3ztr9dVlN6
4nKh2SJ5Wkoccq+SPKoGzT/A5pNZA8yyQ55J6dAIxwIRCXslF9+eP5SbC5+kGTo2/XHRu87W9OX7
/OWGLoupJzCoUwOynOwSZu+CpRwF8gMxjGFYNq6q1Mz841DA02feSDnQtJ/z06SuUnLzrOXoP5pd
I83+o10yXJ1rfpJlJpOVQ6mTZawn7KUkLmiM4zA0dZT5hKpEHbuP3n+rXd07eva//G+6dkyBWbqm
DQef7MCFg7Vnot/nL1cRg5hRvev2aWF0tZ3A8t9JVw45JOZz2Q+kIc/w5qA/Hqwd+qDT1AIKVp5Z
F9Oxg5ArSu7TQxzEMUxOypONl5Hl0MjgNyh4Pnx5bsEncExeoI4qHdiPs6hIp17FIAQjJjygqg49
kGQ026rGW+a18yHKZF4gMznxx4JGaLP/HP98o2hRU3BTn12+3xiE34SQUKqpI1LSuojqAkJw8aUe
VZjSbf+F4nvnnDrQCTMno338RA8xUYMnXklwsKkJ5jCcCej2x9oEzFAwWLyyIC4X2y798IEe1vY7
XqMHqvpM+fg5g68m6dNsP4UxZdp8ZGS6j4SkazFKuDT0iuI6jvnPAPdx6o0DulEq75S0cI98uaFf
2qH5DGjdvjzlvxOJNtdpC1dUOexpAdi98TVodnmFpCsEOOZAheHJsKpcueUT5yD2ScX+pzpP84kn
qcH+y1TqkWxckkvBsnK9LcGox8/cetu0H4DOv5bJjCQpFRYRieDU4o9cOEN0rgg9x01qdYPWyDhE
nFzkFXQFhNoxYpcoPDplHiQHIohI0ggxuEkFgneoDLTuSgMIo170kKkUPiG7NNa565qRpQO6alP4
pgjKRujzW/cNqTGRqHWlQuzWRMnOWwab/xHaOZnlpHXDaJU4CRaUoOy49xc8p2uY78CdAK3wVsR3
c7mNdSZLqaShjLmci7ySNXt4PDkNaX5HBsjQgR70CGqLQo4xQx228Otqo6a3RJp1Urs0LMIs0dau
lSqwNIcXxycAKwUcGDEAArLYs9HHuFhvyMqr3RWzDdytnv1rCbCnfjpqKoKNgtQg3OkqJUZBMJjo
a5JFDB0WPG26+DL+B9v1zgzA+ft8ejYMBEn8uZhsqixbrdQhp+mAacjkBICzVogYXpGiLzSACKkW
egmapSAfiM0zXNtd5KvLB8cF8d9ZUvD+av6ZehfO+lJXg0A6+vMoAeVxgs6dDED8nL/aHIhw+xmt
2tqxYqIhsNLZPBYoB2lKo0aA6QYVxHbSD+B8IgSc4Qc0xKpsg3420stDTaTenW8xWXgJGhttoDBb
OiiBQxYu9OGpJvVplQbjc7OBTIOX4rt9PNNmU764o1bgIG9T8hjW/OnJjsMncAC7FUvmIKmID1o3
WlcbEWqDo6h2tV3VkOv0x36d/pqin77Bza0FZREzHm3FbwdrZBJQZb5TCjAaADY0Dques0hxixJX
Fqk4bQMT/lXXRAi5HB5ch8q+LMQGZn1UwM97ut+amzI3sJou3Rxkn0O6kKhhuA/u19IFfgC3lPZv
DQaw5UtcFr6hOKOWx7DHCgyg+Cxnz6BSFlXSjUcgqsZJR0mkNOkKl/LrNRTkqyYsx1M4FmT/3dEt
aQt4rV4TuwqKUEn/J8o6BJNo0xVIo3qt/KA3Exm0mCgJ7cOf9lTruqptD1bjR3WVtEgyDY+mpmXB
tSQa+crXKR7C0w2E3qj5GUOAEe/BBELZFMdTVSZZoTTzEgcKKujQUfMmAXeQ4DAzmpncFRZ5jmWO
SxQr+DK+2VE1P7JVqKuZ94ijKQlemBlzx8cYarOWwRGZhjVlC0DeV9dhbvFKrdFavRqG/l2KDgoh
58SxAYK4nRYW+3BwJCt95XJpg63ZfXeTIx+Ojvmqe13GnCSUsJcP6yB8r72af0iGEY88QSBHTyLK
2jMotdMTClAhlY3T5bWDu7ES0gs/T9HsKoJvnSo/cQlTtO3gwFJbOdMZCtEDaiwmBUKUTstnFUlN
QwItXmpFcGUXOr7BJS8hvW1wTYwJ1KuZFEX6htKmDex885Lopr1nSfYI6moV+lc0Yg71DJbwjavF
U3M+vVOGK50q6K0kln0lwCJXsjoXaWh0/5puq0PnFKHVD2ktES+zqtM1dLE9+2DB9zjaPdswMKMk
sNFhDLS01wj6CdHTUQSfUx/QnWGBqw0JWDbuzoWfeb/zomGob5wdZBSBGapOhT9g5fodt/8WCJxI
Td2MqbXYRRUm6SY2mn5fEZghzAxZ2Bb8oAK6yxH/4WavkcwFbILjra2Pgv5GZz2oBx4/M+NidUG6
CtjiraZuEsCPn13lUEP28zfo2g5F4reQ+aeC8L+ojATI5tDkGISENZkU+drO9oyAGSjnvBiI/jsz
cNVS7T16FlNqT2cSBuYHI2vaNknWJTEfCLxFwfTk5wbp959pYP2uVXZOZCyL6tbd/qLewQVfiekL
iQNlyrhvPOdsptIp81YmsqPm90ifLS5MFJlX/Q0t6iXzwYsV43rnYWYqSLVxndSsmzYWWjXDidr3
uma3/xUgyX1ZuGrX3x8oDcfUKk746CkMupbmWxbnG9LtZPXDfd9r0O2y5NYh26iHXYAtK+Lxpdec
a6IAujlpVRy4S8fqSuHuS+W6E6UHr4x5L7nMbyMgWskOI4P1db0e9odCQedLD4vJWr0B4LiIlCvQ
l/tQdxPJJa4wljrX4W8jgxvOhVFczG0aBTtDAo/EXs9kgk3E9TyxUvnobVijzFgbk9kcXYY3kUtu
lonQqrVgABL0Pd3giMKynmxdH1ts2eiS8UnZaWDISsN6SsjzTp+hXT1oxpmoOtKdwCMUUbAMiOG7
GK07NXlnyI1ksDRxs8pvtVevsBMxkqRmQDTByFE1j5+xLtPmQUHZJCWIAFA7fIRHY++R08IuVyEe
pmc+onNqcLoMUFOge/jwkcbTUzMJa8felJ55CVrA5WJPgBwJTHIgw2/FzR1p/tHy2Mlf0fIdNDPg
4Lb8DXfv3dk8SX9AC8MVwUmIDrHfZp5zbb7eK8ov6I3Gk23pHLsus1kQI56U3EU+jos/4RNqg31M
Xb83D6fVp/SP+3WK6bfnurh6MERCZeCTbv4T1HtHvXdHoBt2sWkM8VCZUxkkh7bVOS392r2JnLU0
CMrhXfU4VerTJSVeZmqf2eWdPOJOPxWfAfZXCDLaC1HfV3SDzLkGacwV+3DHCYQS+zpbLzTy510L
s0Fjtw7KLiWa7SiarbJP9TCR1pyt7PyU8gpg1VeL9Rjz+uGXVLJgPcoJrmBn1QGasUTBqmCyL2wG
hL/vjUMSjApWGK2m/DA8VTP+YbyK/dDi8O1Sd86t6GQyfKP114w1wCIm8Np9L1BtRuPggdxvYiX+
o729eW8r6euduW18mRT3q4Cn+3OIDuvDtGVAib/k8+2+IqrHeElwaIgOGt0dD7FhTvpxup0U5OQp
oe+BTP2/oXwnzNV3HXdZTbGG9BrUWoGup4tt5qgTG9Y9ks8YI2ItU9UvM4BvYbYeEeCao77i0HGg
dajNIlu5mm64H20pDbvVZzQX8EnTfpt4SDE+uIZ3Ib1X54bffMZwPQ8jK0aZQz3WZ2xJRet4kESu
arMLKMX3B8TCvV4PJheaNP+z7XwlmXFyj3lFGetkzpT7Yw5dj1W7tkKf7x91qomoD5ckOB2mcZ7O
PzbwtJj8WqFIQEGaJ9sO+TPP3q+z9By0dPPzH3zvI1TCQnng7ZHkdJxQ8273Pxcc25FnO5U3ptOx
pNbCa7VDFyY1A1Rzq967Mit9W6ShM5wp0PbD/A+spqnMvZtGd2Vt1e3MCt9BJMxSiZT+SfzA+tDE
jzCzP9JCTIvmTdi0mK1THCxJhVgzPZmPDtLIgaBUPnM8flIvJH7FHiC2vra+yeIL+Y8QKZWAUTto
CtQnS2j0nNRN3Ni3V4wNUwl10uxJMjYDfDsASm4glSBwHZW2Q6z8tHAAPkKTcaVKjugBjafN0DAZ
aBRbTSEevqCDWnDkQGs59S/hv2Tl9eaw8jdPQIPUG4Pq4Bary7GFTI1FT2NnUM/pPDZQLaq930MO
iOqcPK4R9osPjBDjaIQXXRNAHkKCK9/JrfJsH9fyCC5v2cr29vnlaEb15zbDhc16Vr/Yj/N14FzV
eobmE4yAt6+uJxH20cUc4k0xGAz8gOiCm/E+cugSVElAGOpd5L4qUM8m2j6TDfWU4yH7K2wKmT+w
vNO/ztteYUZNZExD3aVvDIlRQVuAkaDktgezb9oFFgOQI3tDvdzggl74fvFkHpRY/+k38Q2pf7Wq
efCmfgSRu0P5ERwJZKn44hEap99MNumwslxFEcFvF89Mb40zyr3iY2Ejbqqnj3S5z0326LlVd5h4
mSrVs7qsw/UB/fXJNPMsT8bB87VenwvrppFMtZs5+foxNy11fVLXGffljkFHwMFbaXSZkHzguCk7
3U8PVo1AQvIGBUBMAxjMujtSq8wJ0hNNy+nBDV2fV0cOkNsQg0wmHCkCvgIuOiAhAFTe70K/tQX3
rbikb90psM4EEqCGhQHpFj/vS6Q/sEwQp5xCq2tsVOmBkQDwbT567OLs4CCyJ1/4kfXeQk/aRSbA
RCw8ZLfS9Uvxqvls2jGbwXv3iJ6BqEuTXXMDNb90DadqtUQ/AjN7t0/ae+T5tElSSlfYXbDhTdGA
/3CTu1IS+5Tj3ovPI7SDQ26nysb8bXklRJBtTGouF1J5tnMRDHwriGNqNpatD9ycKlB/IPuY1RoM
Vyih9meySOmxts5hjoIyEvjvzyodCiqZUlF7ZMVIpVqMmR0IPCPe6nSZejQG+eOVqFtwne5wkVM4
lF2OuOGsKz5xwwzKN8P6Js8irzBiTDtmrv+no8urvAMZ63NQFmqW1LvTh4mg6NXTwSjvzMihzboM
Lt7tiEer/Uox/NafZyh9Shb8BmnPXMANjHnSXRpROmAk3GIWO8FgBDuFBvIX/IvCWXGmfajVDNk/
EFJaPKuc+mvlA/HTv7DScY+MUjCR2FSibhMhNGc54mg2lWtDSyO0Q7Vb04BNunA+NnQP8TXGTfPc
hnbM6F49qKWH/+okurYJK7i3QgzGjLHGerpXp+j/TwIj1XEXJKh95cMvUnd0PCrTjJEjC+iTvey9
Uae7HtJ4a0FZUFtgeXTRnAaBz/g1rD9JqIc3mReOEAypwIe9NbqFN0QXmZXuTE3K5zxOW3oFQCBH
RLGmx3ThiwEv5aJ4yF7Bkx2chTxSHgoE/E6WrKN6GlXQDwmqvHC3u8rtdDuelhip6yu+gU/zwts2
PpzkMclaZq6VyATmi6GI29KcejmvRlZC3+BPS42XPUpoZhL3rSTi0yCmHCZU3tv+rIvUCKokX3y+
2apGUpyaeGeQJSZbgCHBU554acgmineKVnZGu24HkglmM1d2VJ5WFvoZNZ0vppHfE2ENIQrASPPz
Q6YE92l5Lzs8f5hJZkqnb1h6rh/0fMH3wp0bhHn6FlGVhZaX+OhubZtMvscKtWy3VggKJ6bl+YV0
MnyV32hcE1kA2SU2zmnHCjMZennMCES+g6z2bqRo29BINLfGhvFNY+2g2pNoIxDh9Rq49+/H3gON
P331RFVgsLR2xL89Th0W142QXcwAc2x5+J+L3Fm7qyUdkHsuYzQ8KK+LHD4Lh0SCcN2tDAI9M1QM
crEG6kCm/RGMkCZcVKDUuC3l2NnpW0tHYvycdo5ppxoQzk21sGROrf+y6W1kmEEcXABfEC8i6YgC
LxQ+kC7cNG9yyJYXkmgZiB4KRFCnAhWwkvtURnNifu364T16B7UhhMsgvAaLeqQ41z2CWLbmmFAj
x8ZQaOzSEJ9w54JPWssjJCpBIBta7uJ5cVjf4E78e8YMb5scFAtgdiQM+svH2XB1kJ6TRTm3LqRE
rWKqq3QvosQwFRd1TMsOo8VfAoMBu9PVeTGsUVAfn3YnEFTZA+/OhsfHrUAKmudzPPHzh6279H5j
rkBEHaDTrUnhiQzaylGDmi1cwAJ6GSRHVGt7bYmrzrygFjo+jN/gCH+EQj8ZQ7jAKiUnfj+o1K8i
HII1/mrLHeM7mObP2g3S/QEeHzjjKy36uQnpm5ulqmeDIDQ4giAxQTJisI4OgPopjtO+yftTiDDy
Jw7xt8Zhn/5DOXHZoFe6qjBpOmJvG+F70LcJJJWLKhrOH0F3PkQ+qOTQF6uxsEzemxDUJ1y9uVD+
vWGiLzmoTYJb/rnnGbVMYQohBP73WndkjUX2GunbJqIn45vvrWjwBeiOdRjmYm5jvZorWJAlGekr
Jh23VeomW9uA0kG52au4MWlbQqzl5OheEpN1pDaSAVHNeI8IS3rTUMIn0kMh9ftqGR2zHeDvYCGi
ciJ8H83T9M2VofjgJzxSAB0/tlLjhb+SNe54Epw5fGH22urPyxsYmsQdv8HAvGjS/v463wr+lmuD
9c73oBL2CZnZnrkL1YSs6sVebbzHH5dIx2O08/mK+AWD9qzOYVam0tBT/iLIZz2aSN+gfFWhaR0j
hYsVy8sqvrSZmqM/vFirQnkIz5UHJW388QO0keV7RWv39fO0V1qXv6xgGZ7cgRsOdhyF1ralZoLl
+A3FimAFjmbFWyKYT5ALnXeDa/eKBtDySCsko/nEmsijS7vV6cZyRhfLH1bGdygRsUrMiMq8YmiC
TGbdKUezfog6U4IwV3KAMMtADnQXqGSU+duyNL8cQCTJzvVTS8MQAWkQVcR28P7AChhJA3BRWRSG
erHRIaBOqm/KGtwZJNE5HKDkAh2ywasMJ47py4NTjZyB2L39qCRMKzPdcBsLOD52jsxOQGFBCmw3
sSvEsSHmGKcqjZuQvfFicHCiOWNXQNEnnaMxmrtZ1axGPCNI7l6Zpd2Y4lc2+EbIFtS1y0pHdnoA
DUve7+VJUOf5Q58eFoflUMZYgPtbS8exS/xPOof5PqFJlv00366//uz8urrqndZq80lcJVRM21Fg
5Sl/D91CYwjgXjTUD+JJJtL1UKAkJMmCuuo/g26/fy8gNrZxGwCe7IqJo+rkXHjqniFhbVOn9atM
M48j96dMYBgWBxLiT/Cp9LVd+GwzXBvSe7pM79/vFsX7w/esA8gjQUVeQj8Z5mK+a21fmfIgG/e2
yA8AERtSm5qH2shOroYjJIciaFNA/xk3GS0K1vDXh/gZxtpgjneXpw21HLYLGfBloAFgyue9PBGc
q0u2zfLSW1kEpzuUNzx9o6jWJepaY0T2oL44XHhNIGsvMkQcMztPX4cYXiTZ4+rZYPrfqXUlhY5S
6vt5dpq50Xl2V2IGJ5MT8fGA6lVednYMA0jVVZ+BCyUYIfrH81FfzEXwq4kKXkveIvChsco8IWir
ehgWeylpY4xmnvy2s2IJcbsXJk/xs0sC+QaY+X/cwGmLwWDcyfHRd6yufy5ai5DDUCsvF9Br7PYM
y8LAxaWyaaf66vzS8Hhp3aw3sgJCc0Ajdmz/tQaH9cGVm8W3dNJvn3oSpQcfcFhMrDuNfW/t4GCP
AxOzwIHjySt0kKIsoc+qxY5QmI+RRFihGsw7JZdccbLDhmmm/nY6KxgymaafcVRW2EYyjdqJZEJP
rKIXxzs+YALBLI88FG0Y66/INZ9Ujc5/7xSr5mcIdFuSE0br8u+jCB3EiX+yy205Jdv0D3V0pmfz
EIzBvrMndEPqYkGMyHOJ7EsLJ2dK2jGwo9c+LiaCl35P2RoPPRAxLjoo0tfcw8qcczbGGHSLtM65
LwtAXP1fwUGoQHuiv9GnHHRNcrJ/IVEK96ouTwYCVGKYMjJ8bW4oiDlme8Ze1JYMlGMUn/zlGBq5
BbzhsZ6wh8RW/Oq4c0d8QisoDr+TjI+hPP7eo9LDXErDMtBv+Yxay+7f6af5OA8OEvGkEPlBRjg1
a3yaTLvALvb2YXwV7yX+/u1vFCpUhH4s6lODbubLjlyR86o0zYnZKzj9HlutR87bIA/EDuAkrom9
+Aq80jEkf3AK+DPTMb9TDal6d+HFgHRvNo0sbG3LZPO+IbWOQVinQ+xidBrfcmQfa1q5eXOipGkn
DmT5kaGxDs4KZofYJRh/yUjo9GmIKhwUTEBEoX+mUa0qfk8a5WhvZgNT+pFljHdJ4iQCas17JPPR
bCBgDEY1hHNf/4Mr8xn8nEuEme3F7zmK7LaQyfTppXFIktOgmM/4/3FRYRXysWLMkkIldwNby1SU
VFPSdHUF5p0eKUfllwnrnuJXWRSqlAYqQ/MibQdbBgNneMBzfP/gieEmeV5vXwlV0tDBVCsFjcfS
vryvED+lsWUVLavaIfO0NZhJMKyEh8PWI9bvLwT/Kjf6plwlhyikKop7EIsuptJ2jq6R+k25vuuc
Ox8oQWLqxQpNQ1k2Fm0pAmwZz4hMHAfykjOhFcfJX9En05X2LqXOeeJ1LvxSfml0NqJkLYCrYFTj
6VY1QAX+NjzLfXn2zV74euZzMCVhTo1pmlnZVyFenQ3jg7tEviG892gbJ68c4WejPTK79NqH7Dxr
/0XgV7PNTQ3V4LGr3vtpXA5JzY4bfXlWl1XZlK6ZSxomNTvUiPzdZ0l/Tab9TNMP/hct2TrCEX5j
oUe5PEtvhDirrZsWkVBrT/J/MLEeGxPZgZYvifcIgB2sGkaVP7avXU6A4K/KmVgC3cjL2OmnW0yg
hmp28/JcreXA+5IZlF2+CZSql3Y92Dp6+Vp5gbf6OX4qM4LMneY2Uh6Mx2DPr6f2j8AOQRLXNp+F
iKgC9qfgdguiCrQc+HJTPkklZVgE8X5QIFHe6WEqkUSuK3GUiOO+Hp+p9i++FZ6tJwEZHJhBRR2G
DYXpJpr7hC3YZ5m/XdfV/t6lILChfXCyZjNVwx5cyOPA5LSJzxwo2CV9Qbbygqpju8HPwmRCh1Rz
sg3W3TRD4JG0xoYz0LDwl+dmBQYV94mjL4UUaC1iGsm52J+1yzcMbq8fCkrYX7OM9BNxyib9L51f
ZhVbHeTsS/TyWLMWJJqtoNpfwyN0PTtsXcnPjxvyvmHTx7H9VWJPa1Xivfip7lT5S6Ncpz6v06Zj
qHUFla98b4sSJJuqMKtu/+ER8QWDbMfzj4SwGMkBSo4LwdDYhPSxNZ/E2L0DTwxfkYY2O7PNah3k
6JT45R6zQ9e4RfSDzrJkrCME3Kc3/ApzmFYOTMcZtdKjRjjpvjQ67eBkRFjy3eFx2egfFJ/C/Nxd
lKYVAlE5ooVLlYq36bRpXj5VR3v0w9CiQKQF0v2z+Rnj0vXT9UNiR0N8e+l3q1izjyrxGq27cNhb
RnwYtSloGQmpHeRR9sURDJQEduLxXK4dwbxL3OJlaGMImstSzuPSDqRGvfgPI9+O6JvLKyWMURpV
SOAKx5ipPnJm8cX+HoMbefLip7cyY31HEik0urTgxkUNI8jlZ1awEHvouXAYSqSFV8DPwoPZaHzh
eCfwjia82VkFSKC2yyelPpwzr19G05NFFFvguSaqvJjkl487e+vTwTkP6uHLI6W6Rm8R/xqov8Dt
eEYEiiwqU3bA4ODqV/Mp3OMOAmlGB7P/egTxnxh6g2Etypq0lFQAacnq89jHHmltvTyNMUSdNgnt
u0TxhhGA51y+uMXqDlJqZyou+RLX1gS35TS7Oh4V/A5SSoFxzzhgV2rtpUt3+Tl3IylACmYlgGnH
j6reI38Yj5qfK3/m0Pook/SMkpEqEuN/hvzdCqLYsPJsKRxAERVJSVYDS+aSs/CoC3WsufO/owJo
T/8ZyW6Ni+wKYIAf40CzEvWZINum0hY6mSE0jlVCNe6zs32/zv2v+4kq49XxD3ACbYDoLpU1CxOK
aN/0o/3m36IfW73JTtYs9TudFotkX/xDPGzpUmV+3A5rCM6wAJPPni0mdSGH6n+45Yl0yFl1Wq0t
o1v1/Z/cVVIrEOWagUTs7R/LM5yzM7DgBVM7aKYkG16WInp40Q1RL3wbaupH/KPDcIU59500MF2V
DhWc4ldrxALz8lHARFUnAELEwXo+P5MisGcpcKi05K8QWSPKVr0nlLcr2FNM0bWuv2tJaq0fVmZC
Vufr+p2PnobHCTDsoUlzUPO3gSUWb5uWM4Hwz8EwVKk5gsgdWGmKdsUTTfhtLBNOt4X5V6L2MNKQ
N4nu57+0OstxFNcwIMtcNlJXdYkRssPQAKqWBLZwqtzFms2ro9hbq6obqka03o+e2dhYNHLjMqa5
BYDFxY34TTKttF35w1VLRQ2YZ0/QE6Zr6JhmLxHOMNagKCb10T0vtgk1uPhyYpoxvEb3TjfCVdKk
Ek4QvPbkjNkBJotu08TjB5E9QMOSPw383yiHOWUouUZB/k7WhOfMKqF4ivWhiYOOQr5QTMk0dfKs
U2zExuhkuPrUfuLacnqNHB08INjGXKEWAl8CMgyljigPn+YNqykkB/oMGrn4w/t4Hg6Twte7X3nI
zFZws5kxmdZOLKD+L0SH0Y3FsmVIzttaCTO1PdZtS8+3Zhmc+5kkymo4HhTODSD5DGeahG4fXuzW
pF8WrJaZjZhTtlT5RexN8AwpGZslGXySXQdXvUImeZFuHhgTOSJy6o3/JVjExk3YZKVVdqPxmIL/
NTTaslykJBbE/pdQsN9xW7rHXBHQKTxIchUuwm+CND9kSzCirCNmbWTF0qJIYQAHiB5Ig3gSoFjz
RrDejbhAZ5vkKqX2MwWCzQlcz5HzPlHZnC8clqzRnjF0kz4HK0VZunaYzdDuzqKiNl3+wed7nZy+
qRrsNv8Xc0jc3D4VqBu904KaA7k3zjDjIrQM0vhbIx0Wp7kX0rP+gNy8chjPgVTx7WKPpZFIZ8lj
aTYy0YF293PboQcnwX/cZePiI8jtX58cUbM5MiY+n0F3UwOLxb2LLWHF1VVaf7fUWZjePGIQ4srA
lALyNidvQJNLH08vYDrkl+XGfKe+XHZn89/F2uFDFDqcyYxkW+fO2uXoptht970luSDQupRs9qPN
0Cir7Tax5IOory0mTrvZ7v1+Vhea0Pw+v4s7eXBXIL8mJ8hFR3sS13VRQVkdtzzOHnkXuU2ph/L2
1f0FYadQ0WI0hotsmfDq5GKJLogJuLSJzJROr//anYdMJEaJybRt+QlSJMarDUwrhXqMg8P/uWCF
F0IGSL103U2mrXFhGnvV+aKAAphfjh/vxoR0l3SznG/4afCZlE1If/KojUPCAmlTpjHNxoRPw+87
M3nZt6QBcyKEtirY3ik9vTHdMrcCYzT5+zxzwGeGy/AXn9zcYz3kqh0a+WOB9o7dlYh7YpaGnCSz
222i3SwmFHJ9QzUVI1MEuMZ29kBARIqiHo5elAuTey8IEWx4xxBuRKplfMnHhTpkWAc7ymMiXAXD
hDOgVtEzQ9SqH2BRPaLoL/8gszpVvrLQD1+E5Q46tpiVRE/7rzhUhgTyBDRf2ddGjck+hIZ082N4
yE9hECGgtpGAK7c5eypTAXrcCE1f2iU68L65VFGPB5i3Uyqo25eH3kmcEjQRF4yk2h4V8ay93HtE
snRpnywa7XYpexeP4fZovYtFW4bivl3DROxNWJytF+UEUjRGMn66IVOrT+ym5SId9Rsh+sC8kzCC
yIbsBRe5kl4kutzQlvyU5KSt7IAqD2+8LPnaRCzYR7M0MvlZPKd3xia1Our5+I2ruQwbJKmoRhKi
IH3LYTieHON4uUAt57CWCr8fZnypZm3QF3aR4Modq72n+XuxtNcg4K4592Z8kzeXFKOo1yS17kKn
xkzuXWkS2FctVnwaUHB7flCM2ZcLfMnLY3ijkAcI8KCY7HvObeSs2nHy2FrdszaPc3niU5G7xhw7
0DDcNHulpbPckuC4wi3VZQMSpKGAEgVfOf3hJJ5SPiYYCwqmX3osLDpW2xt3xe6WXPiI+VMk41nx
RtB5gyhh0GuS15/DuRBYv0H8VtupN4UAaPKraB+WH96NW8SogFapl6lZMkFvBWY94oCJKeFupOB0
mMcqlpeJy3tAAOjkMyWHyCph3VZzXQ6aiDaB102w4sfwX5bD8lXLHqLLIrpojuSzutVdCxraGxf6
rKS/6O1w2kLqPVuBAOIkh5uShELY+vASlc5yDZI1v8FyZC0xtwdBVjNBeK4XRYun95mmt0wa4o+x
4s3HZ26WNvqI/CWxVnOLOqMPinPs2abSUNL1rjSadlh1inK2HQS4M8QaeUE0o+sPeZLleZv8cefr
gHGTLT0IRlbIzZ5r7X/dEnmqGv2VvIX83MlrNePbjocwWBIamKrCUvMVlHFXvxoMEr8cPJXuOVgW
y0SG4B4a2oTQrZOiSudYtupn0KUDxomhK8wS2zafuQTb3cpCWsYPAGNSJNQh7YBL2M6jC6fDFgRA
Z6pLvc8yl4MRCCq1qf42OiFMKMPZt3Kkn40xakV96rpP4Tv6hift0/TERLewTCMdwEYNHHRtt13v
0H1zdgveX+/jrC518/gL+63lylf+HLc2oG1xHIuoeLtHQ6yrQZTTjXKDezn1KSQJ/fJPTl2lRvaG
TRmgJ++OWd3nxOogbpwHgWDokcfAW3yvYXTndubrw3NT9GKfbe0RMre601vPJEeCJQuqsJDzdJU+
2h0AtlLzDaXJcQiAa91MPCnsSlFh8h4GbSTfJ29ieH7riCjfk/W2gOgfrSVN69PcPWPFbBwGtrz+
WPoXlc7iJjJfykNe8Kpbhe4L222NFqdXPsSPY6MssVkdJmSUXRHpd7Xre4+VHHW5ORFwDCo51iIR
4iCJXQSE30OPEIt2aeLUkMJP3ExmoWiu/Ob1g2QLmp2ZGSyscMIP3Hb8kEuYhKrkC9tKKuxbUqi3
EDS1aoEC6zgaqm6OXxCRNc1jUUXbdVY2AWwcN05wJhuFg6U9sZO+JaldATF0jWCBJqvBT51MhtSe
WjNEQnusgovUlsmQnjpHIy+ENqGJqR/gZaLWOsKwIc9tRK4XDSzlMIX1oZurLsncZ3kuPznYZvjs
XyVNOZ03CgqWTLD4RgX2eVyZdrIoJtYKZEiViaJAfPL8Fe13OJZB9SuBuaepKqQ1RefIvI/l5bAH
LY4ghLuNx5AATlPeEHQpOyOPaUgdlD1u5+5bwK45IDIQmTon01+D9v7LNenaF1R2muZSZjvGY0UK
TX8b66Y9UXw/d76A4lpaFto1cWZisSdjLqd0ohQRAhAEd2OROv5soTOYlP4DaHsajlqz4JsIocfd
93wAMqyxV9KF+yLb8/8bTfhSJoFlCfVu8Tvl3AmmoJPDxdQF0hKOalG3VOqCICQj9/XEgA0KABk0
rtAk+C2njpkbj+H4kbEHPOSZ21/BluoKTHRICPZPITmcUti7Rag81AS7/gTudCw0CcqPwUtqJT2a
h2u2Mu5hSaJzMrjNeHB9JgedWou82aIo1tQ2JdXvGGUGjHNFl3fjO5CpJtXh6EdLCXmP4VGnkcJv
H5XxgpCx4tLAodp4nsPE45mXSpTGQjemU/g0cOrNFuiAWPToEE5NnWDEd7vU+7oDcwTQBbD8VE/d
v7KGeXzrP3dKNluFEFroboByynfjgIUBV3W2vdmDU+KnvQ2LHs7Z0uIm9V+YT90buMsjTAtYYUDM
iLE5ZPDe7tGxqGQ0L+J7Mfs6NHQBfgPB/uo9paU4g8M+8o85CnUiHJNmlcqTvrYHjTNlawO8yB9z
FMQLJGEhYtNp+1HozTuIYTyfGrVR/nacbJhDYcnhE3Sqm17wG63ZlBoCi9XIB5SKr5QgjvhY0C92
NhnTCpZA27wa1dqvnVDSsaYjCxL8rLM7uU2mEkdyigYEa+gPNpC2pszlL3vRl/QhAP7nnNikZRBR
tP54RbF3TbjyfbAgukPR1Rh0VzD7A4JqScrv18jGL2BQQ4xCrI3Uzncr9BB3j2YqI1sVnN66iWMw
cS0EZMLcuxIBS+OqZ92gMIkHZOfEdPpukZTHrliPi4Z4sR3SJsm6HTxQMwQNUF2/rZS/UhVc11H4
svi36eG3R0eBomGa4Afp6QNftxhvSPP9cA6GmAJR+FpFAN11y0Bf7rUWxjb90h5/P24PsfQ+1tsr
2F6zHgyZVh8/kcyV6agglgHpnyJqRCF/U56n7AMcqx7xCQJYcktguFEv4u9USDIflFvGsS4qoPOI
V0AKZuRmSsYeKbX5UpBvtyKJ+vB493/Hq8SruMxFCP55URMAda0KvyVDQ1/SxHuRLkzCixd2J2Dc
V0YX7N45ET9wOQWgrnYvJ+Vz+JbWQfQuQM6ZriEuPPC+hkDeH98lOfkqb5cxdcHrwKIRg5IlxNnz
i0gF34kglw04OKKEXcK4lPAEeulzysg4Mb/QClgQuesSr1WRRs+TiPuATmos5kOrk2W5eBllg6fx
KD+ESbyn01vs9xYLmNdeTP6NHBs6WglHW7egMHAadYqHJMswdkD1+yatGi0UgN3MoedGaEy8QNzJ
eptcRBUIgd1mHQvyFGg822EysYDLbYYvYBVtiVRpxN6exuORrQ/eUSQg2VFETvi0E59I66uEGMiT
yjYb3EeMamsussPvLe34MkyjWo5dgo9SxEzlr5qt8TjIHyMwis6zJ5KftClsxvrEFIFLFnypJWjE
Ey6iVimat6czdZ3oUDAVq0furTjGzfyCQ5CzD4DJnayudxZkviV5gl0OwdxkWgWDH9Ycl8DjjLyP
ppTNsbHox9hFBbX71o/jHwPLulce6Erczu0X5BjuJZ6Xd3vZU5keK9MPa+Vaq5ehxqGpHsXlJR8v
yIyK6NQCVtVPZfJKzeBvjsvdSqFqVxoapEwQNTx2FAqtuIfUJ4yO5Y4wxFEw/EAeAQ42Unxn2DnC
IfMIQyn/fA2VnAr42FCc/7T/VpMXsZIOhC+0ONeGJ+ybFqKPfP0BDc9q20Ut5TJxcfyhsRu1DjbR
Aty4cVFhNsocmOZPaEyFmScDPsaOEY5Co70jxux2nfKptGp4wLjZxQIFIWXctEzSES34fi9UpVc0
u9Ou7A8fE1bc7XuLsUCcpOlZHS51fRtz+5PUKtB/dQs5tpGxJlkN2tJqKH3paPKlZAdZs277VgoV
jig7k6VQmPezqko0JAlkCC4/d7r3qTJfkMoyroDn8gqbBliV39P0oRybH2EGSy9xOwDif1b/e1j1
mOmxKjD5D6X5lX/KJUBZgVnyonC54cb7fxzTTZweamgyXEE2cG8wetU5/NoN80D36WWkP9JYkAXi
f4Dqx/HZdG9dR2p5TQ3016VWVWOQCAnt3JVv7khYfLY53Ehhh2WnXt9GQgGcm609wRRWSsUXenDZ
pXLZWyPOlcR41MLnpOavlV3acpIIlkyTbEg7+K+D4c5e1s1VJ3Yi4zjfSPNtEB8Knk9XxYGx5yl1
GutNZrpTs28gPJ2VlvW0r2mczOj76fw+6/tve3cGAaAuoJFUFOCJ+RcnxiYDxQe6YNAWXETQQ5QM
9kOQky4iaMtkDJGePfM39k6kSsKRKtvZLeg/Oh0Ycx5kEz4yU0E8Z757wY+aiLtpcoXEv0c/LMQX
1TPFD2zktigvgIyOwlcDrBlh/xGM8n4CE00gFKHmeJ3+2/GaADi4wGyXbAgaI8cfxJMhHSfOlGnn
i/AT09vx/jubr2ivV6ibq6t7qRRomqLE5VVRLEilE/ChERgld86jO+h7jKtb7ZnPuRxc0yP5anRA
DGH0b9rYFOnwQc0h59hXfVD3KMp8+NuoNf3DldpOja0LrLGY4uw8vv4W/8WSNhB2XyYMp0LaIvUg
AYR6RjrTyYVdc2H2jL+EsGVGMjQ3bq6fomLR3ngsBX/f/czNg6cchizMgEF9FYIB+yJuqh0qfSrL
egbJWEBNJoLkTfaTLbUkKFENaZzhbnvCSG5De7LoO4OYU7AFvIZZ3i/1cWAJHQJRr483lQHOlcZ6
uOe40M4nVE2hYSMDCz7JHDAM6mF+8ixvuKupEN8NJmWGZoh3wuNrHI+LS0GImaw4j23Vxe1Okgqj
eFkJcgbMpBjhMl+Wtboe1zY5L+jigYEaWeU0e+nWhLP7pL1Vj+cC2RYMvWUsRZRX2y2ZR9uXay+9
rUfM4yDtAsaTWEqVBQCXEM0YDgMW4BSIQxeVK62y0xjtQRF/+UNvpQYIOYokyY+ytpyd5M5DaRMl
2f41cTocZ1Ryc+L1oUQOvPdtiaRRw9EowUGC2ft0pWWvDepvyiILCzPTUvQkxXGtXjsR8KAdffZk
TYv0ONZmkaKPWs9YjYnd2oATuZI7ZToKfLO/4hLZlHubL+EOLYebirNXtVLHMeUvq2zkIJ9qmUo1
pTr8Gzn5APZnUH2VJERkY4lLlKFjq6HCcDEFgN16APSgOqvwpnPepuuKrL/o9Ia2364JFufZGaxs
QiyVx5JvY5Jqu7DiMGYrY7UU43gKF4NuztAXd9ZvVDbdX27tWEbTF7AROR/zGonE5NqqckB9d9Tt
DEmYrY6uclwZHsd9qxpEPZvE1njq7o8JpWQRs+8yEFxXMyX/jqky0xE7ccdLKn0bnVal7dWZ1fIo
zxue0fcxBRXIxsUEWgs9RlGIHFUM9coTknMW+IKkiHomP5Fbzzn+XD1939osLOoDoXnE/T5snsRD
APGV53lES7GN4POBu2+JQvBfLfY0oHg57qfx1uuGFQqhWnxCpNoD5cGN/l+O9gAH8tfZ1zdsLbpz
HC6+JqIqBxsny9gWB1vSSgWsc7xvVdmjEdiM/9Q9tDRVTfHjZuHJPSQCg+8x26wybgjlv5eiARxr
f35f3Jh1/G6stubSD8xDsicFpHVNMBsM12MwefN8FWGk7qGyGztVZ2jSiESDLex5CQwMLYinoBEb
tFVWWFhQUW1rkgqyb7/LmQY8GiK+c9i2s4lZImwbTSNKIpEW4HvK02a1MpRuPtRXA0aZH7lj7tkT
MNfhFnlRgPeLv4sjqDwFytl+Upr/RmG2YwtQy+6KqJaNkkfdHtS5bXvQpmfRhdnBgZUf0E8pCFZX
z7jyX4P6gv9Ny3FUWorPZDA/kipHK+BYxwiKwpDvoIWh34No0tqRbE78vDLXw+mmH+AlyBvj6Dta
9h5jpvWo6U7OIHFogpLHc/dcjNwRBw4vbeCrM9nvz221DqeChGQoCKYz9lNyvgF9qTxFZKq6DIKd
JtL+WJIbG4oyi1X/5ojtW0zGmopItfdqf+wXMct45VqiUg2ZIsjMz1MDoQgt/AwDtS+BNfq5u0pp
HYJyCVE1RL/2DhFK2d/4imqEBBddbzrPfP44bvLAE0PmGtfCjUgQ8IP4Ium+mQCQZGVcK1ulIaas
3FbqRJY9IpPro6LDHktFq6aHSgykFwS7IVOlOAIJ0e/RsuHinmuDRHMvR4dSBm3uG2POMWx3+toC
G5EnNpqtnXrSqim4hUbasvcb3fMNbvdo2jUqiGK0xmUPE+Ew+wPDpTCSjSNyhV4nmTnFlwPVOPKT
CC0Si+CLQN0+Y5NDhvEcJjwkFyhxbHrNV9Jp5HvjPyPJSGYaTp57Cef+Fa2R8rKvy3SQaYAPEPKW
o9BabiaPMI9qw17fe0JS3uVaLXtQusINInFPXhauwbxMdU014RdwGaWSZd+hUrvcFL14PIWLL0kG
xJdVIwqwCGmf9+W+l0Pte2u4qvtsztnZ/QMft7FCfK4ckrIzDDKYwEvcKVGSHVodLTkv2gfZaZZD
nq9ZcScLhO21npKoEzPuomsDWMpA0/gzJnmrN7Poxhlc6HmSey4Ulux+vqQw4ChPJwTT8rHVsrYF
B7gHpJua5sD93/HKNIB74ftioXO5neJ8hBmSbeKuCWtYBuqMXJnGZivAmY4dKpL2JaW2UlyYuNMc
VON8UYFaKzuXo42MSqL5l5ag6t+2keUeqZ7g7PNZMCgJ4F0/WZtZUXt0CQaZhXcD6GBZz0R1zMtQ
LS4ezUgadzHYqaX8emcrSWgoVj1c94hCyYqSZ2GqVeL7BMpQ0tsj28yT4GgCFn0VIq9lcCu3Z/Nz
0RoVjzbEVGL248H74xUNA3eFVBtTQJuW0MlX5qdrXM8cJtIWpJk2HzGQzdXmQoSs51NzOVwBnHux
O+mXx/x3DhTDkBV1PnANF5t2ngVYT9wf5ee15mjYD3bsrW648E7ZvFtIOqFQuFWYykC9KgREyliJ
iA/hHqpcNAzTiXbsoELTDmRt+WlEdFTHh3BuAkFieOmI9rkD2ZVjKhdO1RHSfrbdFXzePDmFjFZn
5P0P8aH4akd11A6hc5Wl8Wct9lzspHeod+jp2U+wxTFblRrDULvsPt1twkGJH/ScQysS5npCYQaK
wIkByZYb2afGqTTrBzS3d8SevQ7QvuqOWwE/+HFGAgFwTYKTIbna3kLE5k2qPfrQUPDovHO2xI9u
97H1oPSYkbJSvsiSZ+cNxBAhu66NJcjCOKDJajjGXRLax4Yy7O0ArpMcwH/rSfDQzBBlp47FSmkl
RPqPnrPotpavj/cdAZXSdtcuoacnQCKdpiw4/aaaJXzS/70T0Tbrv361yuEB6dGGiA3E/DiWC6tL
AqS9ViAPvsS7CSEBfxR+OlgrVdP5seWdbm8U/qYLmc4WI/KHAw2cSkgtGIPtjneem6aS+pNEDFKo
r2DoVKACT0/+HnH4in3VFzyZd+p2gOLpr4HQMf2x9y9SUqHgmER1rhN4i269HZS7OZC7To3Ysliq
N6FGJ+VCJz/l0XPtJ+aLcckt4MlBJVdllJeflItGL+Cxj8z+5tCmeGN2+0FlsbKkO7Ofwff5qTeU
TSPxBOiMzwI/6+Une9fsX0p05ohH9hsufPAqrXn+hwK8Yo21jifXKSOraq2uoDKTAqiC1ZXpC1rj
OC9WzTUICfdg7Vco8FQ+XhIDvaYjXxvzD9068MILROKmRVx8QakVZflg78tW48yAyKQq4jSi24Tk
wPB1Xxy4rJgHi51e/9bwpC48GQDJQ2IAWLfON5zV4GLm6cjS80n3uOLBcc0fBF1HWfQQ/L36kOBZ
s4ZpzM/UyrivY6O7DwoPLsLB8aSxcItZhhHJRHMdBxxnIWSYZfSaQDtrMVGXU43wyA5Ss/Vxr6pz
eDcRBKEPM3BOhFEm41T+teAKjpVKuvhA3KA1CLEC4ZjbvhkmxrZ6+SIXxbNiAVsH0KbubETuo3mw
tkaGYgop78+T0D0oxw9I7s85W+us8KyoYb2NWT/3kUp4CN6zjl3jOnVcggvR2lkIFg8TH58tJjXm
TSPA29QBllXtMQhxrrTMW4V5dh0jefT2SV/tStf/Fiy/Gal9G6Ipjp+2MTomhNoZEKKujZUJGEel
9OiucZk7sqMS3eyUDF8kO5ABy3DL1CkDvgIoOuxpsBPRI9ICJYH8+uu0wFESaQHgcqKHhk4yYjHv
urSKZE7arbpZCQoDMHdXrPvWwC8DSu49NjC4G5rEgtmzYbpfZpnD371u0zE1jpP5gc0/f9q/fK+K
T3JWRs5jfQrXs9c13X7wNIb+2AXXXOvd3kR9+rGi8COnKrzSs1Hv8vP8wxT+Kqs720Vh8XE6bi7t
wCgkmmEFV3dZRt2BY9h+DjdixxMpzKUy4v5kMc6fM76Z1+sJnCnsi/kPYRDmdyW4tmfwEiskRIE4
DZBgTP5pcBY7NBvr4QMh4tFq4Mj8oZhsHJzxBjHALszaOiiZ3eXbYY84yVB3pJzhdMXC/z4bLKHl
afWjxWcelRWee9d+sZL9hNpy1AVOwzYN7XajW5ycNTEsjnpbRmZp1Fh45iZW/kTHjs6LhVPBUd7m
pb+3H28+7P+xQutAlBAK+qHQV4SCH54enCI+HAiwKQ8rKxoSaj+iqaZHJR/qRt78rTsARiAzn5GB
tjV/QuTpLLD1wZK3JiMbVd6RcoSXMC2BXVwn38MSpXbwp2wWfxXZRQ5fSOuAAHNbpURBMWE/rPjn
+j+twZYfDg0VRfx9rquKytpHx9XnjzVnQ4vhNX3xST95p5AxPdHTSEceEG51ZaOZ/iQYYGvERhMY
mdP5jWzL/kyhXXl7HvCaUPPKQNFcz0PlS24MYYBcVTDcIFzajLknPrFaoyQt6AOm+z095dL6IM8M
rzGkTsoJUCTMmh2vdWFEWtUwy7JFsQ5Fu+bUS97vnbrX7wmcmNkP6VOVBxVEA7Jv/7Le5YbxlT6z
MtQhLT5RKzuwMfbmfFWM+nGvNGG5z8C3snTHk8vGKTzvY3mQ+cKHNvFs9+wSxNhbkf7RqhU6K8x/
cy/yQ4ecHFEr0LJJESc7K/mgMwzivmgSyMpHL1Kb8C0O/wWmloge2hcz9nZJeCEnvNom6ZCLLXvt
eJN3DladYGxEZv2lDY1NUaYlK/DRromgLz0t8PKyvbtqnZHHhVAJHeJCIBkUqG5cPxKI+geFPU6B
5eQcWz8MhUMzfcaCOjv8BG9+GUz30jWUCNVtgJr7/3Rg2CPc5Cq/+jVN8v5cUIZpyzRZJeXjV0HN
ssufF+CP1RL+cC9StIcCjjKcrO599uvrPEe/e7D+tjyYYJfSyu6IxdkMkp6MEFIddCxH1U7mB1fx
OID45TRqwAjPTTyjeZ6ifVLmnPFVq0NXuPYyXDaDTDdmcoWyHtovmL3iXL/+AaKXhvrer6kA4Ui+
iz6VEnlMZybO85Pg2P1IS8IVJI1BffzM966EgfOemW7EB/b4d+DJ7kMqgG5aYMtNX2q+ykbkNGuL
0X7ie2AW2eGcQIco0k4sWe6Gk88I3rGG4dtO9tgPe369KxSNCR0sf8SSPUz7+PIobyEeh7KcFpaV
ATLAndy1vrHU9yAECVYrLAwFD8MTZSS4SrTPUeDd4IAVQgPJTjZPgvOiGf9Y2H29+Rc42dYilcmh
1IAOXhO3kgE9PCDeIgZgDU1bVYNANWLmYEKBXuLypqDiSgN5Gm2/QLfNfC2k80eguV2W4czfCR7f
/9islqj4McVJRI/OJNt1KK6kPOHIJCpLbqqRSOdemP4VqcYm2X2m4MO+TekLji2gnOa2p9bOWOHV
TCKI6dmySSahf+NvykisgKp5ffAYz0VgwyXjttwVvF5u1Fsm0UkFVcTi7KFBtjDc4+TbeXXzkPrY
pLZNEMIeWD1/ERJlopmwUdbWRyfnIOiryLhPSPXiUJwLOK5yip1zkDRRkrXUOUXb84O6GAwmrZs8
GJZRXIISunsdURS5B4YKcqCmgN4b+JkalBkZS+oUL+UFsYz9WQ8ehUwnYJe3wlkGze54d1/Rooak
wtguOSA1O1gKqx+CGKUFRku23+e1ccizLQgwUpSGXoFaRCraJMfki9hCkWayUaftGzY6CpMGQ0wz
OMYwWJHKNO42iDdh3PnOwfnsuzD7r0NprqPQD0uQ49CiKct4xU8UaEc26CK5BMj16FNCgHe7NdwL
ztjFlqt5M1wx77es6xaYhhlvMsPRYCIGhw+Px/bXql8KYLgfEpYAmhY+pZqrtdpQKW9bhixGBRWT
6rw0ab8/IF7C5eJFPUCUjpZl4UiRgTlIlMzZPbF194rOG+uEG8kCfRaygPrGBUo6ougOEnP1iFj8
BQ29ktM6Iu5btSQ/mkE+y8lNo+/rgOGX55zEUWoUB6P/F9dws8ogbbP/Gcm1vGZZtf0fWfM9Ajzu
adXAfB0fssm63w4R/15Xa20S6t3q+SIHuuTN+jGGC0MARJhccFtKwnPIN0sE8Ht30u1ctbQTFgBb
f4k6i0cubMDYMWOTe0kz1fI4icQq5fBwlq/zsB0DBnml0YQ721WFmkbiwn1ihE6sNb01PYkWPGrA
AOcMivSogvO66XQI83uPKVKfYx6Gs/GE8FCKFPdCoh85eDlsWQmJsheXkS3ud+k+gnLutWEz+i+7
ZgzinwRg3cl/TvfOXgUuaA/xqkYnYjHr3ezl0vJwV0vUtP+5jGiMGQtj5PhIPxFH7JewTqj4GSUe
wjmY5OIM2gtzP1s/K3QAIngZaeMVdZV0zC74HtceKexXGpP1oK7tqaj+aVjwVBQRfEXnGF+jmnAq
0cCcS2tfy1JDAmdtYcgJeyM+M9kB52986mFFLa+ngZk2n9v1ss4Fi/zSrvcBRTQhDE+0fCQP9BlH
AqMY6QVojSA316Ss5+qAgeRRpFx2tyXDw9gqNNtfXSrElZ4JVgB34OIPUnfyOBvNZXkId+o876sP
vQk1YGWWAZkgnE2ziQlRT9pbgCSbZSfxkOZU6Zy0dMk7E9wW4LhL+aae/nvNu+iZvE49gynDWARP
crw/HNKxYcgXCmil2DvMPTKbAaJZSbtGXuACrnHBVdxi1Awhrl5ENv62mTbauh21yz0s2hyaonUi
m2xx4+rGbqFPYUMIkFdHZP3HpGK4Re/pP7HUlir+ZRD+3Qm0qQEV4hN3GMONjFIkmsArvJIkjg2X
q0nYbrFXsNVIiSOdROdw8sbgaMqdCVtHtQuNLIygW9A8R+xvyJmEAiWyn4ne9XJ7L8CCWgjmh7JM
kCSyuIs46CzSsA1/Cp1r4ZwFzJFaWuDTelwlw5nO7ZD2QDL0tzRGvnioBKBr3L03KAeY8rdjdVpn
VnEGQvAEzUJU9fgztdHSTBjM19jdCTr33/eZ82dlzk+fNvjl2fe8nffMJ5v+0CygUKqpylxHT1HO
pf7lNhpJYjmr0Y3VwbavfP+nxwLRW/0tRxVPGlVxoKsDCF0g2BPd48z6BbhPmzpjizQZrlriPCJX
wzZTDoEhi3sFcmK+fUqSAKP4UFhu+t4HB58jCATQ0J/MeQ3OXfsWkkDausWUoYq6UvOuZvm5Ub4Y
waUVBr4jVRkBGs2zxDcDTQ6+nUkRE1APDti1XhlOMX0s3p8pz8DNi2BtbInn4Mp8p//RvdpmAfFi
wZW1J1jRpRsOTuI9hiELX0edhSwTo/9zMkEAC+0dwUPwxxKpFxJYAmg3TMF3aGe9QYeojXb6QlQX
KUjP7bRUlLcCLjzm7eYg+Qrjo/GVwYRV/5lG7dcQLali20n+dxCAgTRjMezRMBlxqt4yziWa4oFz
6dScOTB9ISmkMAe+Z+8GVyHkFTgaQhBuU1+I5TnKAYBt0fMW9l7XW5S2q8UU5t8zyaLJVrvUd6DD
FZk02wweEMHCVpojFWuhVSrczSqSy7Om+LJuoK/5W4VASgAFhAxZr/DJu/qcQhNOnNAJMb+c9P5F
FwWFJHsmYn+Ed0P68XA3fLgz1e0YRg/mSWkCBaOlJNzbMV4gNc+txhxDqj3mwOCtCu5ipu8VDS+V
q+InNlEd/Wu4+c9Kygoe7Ez9gMlKWhg+HtVTWbvX20aagHRzeoiOO+iFCJbX4EZV0L8S7j454UHV
82cPBCOrU+fOC0wyAOXcQsKpZ3JJymeVD4pLonvAKviaLQDAv9CRC0vU2AyA7QQwyrluRRSDrkPV
zUKFqRLcXjUhbE2P8GUM3oR/9XZqvz4Zc729XvTvhf1NIfJUfDmJqCbJTBKd7s9gJFSa0TgMmR4y
gEH5vZE2GdWb4Y60l97sO7FlhF3KSTBu1hiKrMLPz5n+XfD0wPesx5wDNa5owegtQ5YCmle151LU
YL7/wVOme5Ivb2DKelxSFm57Kq3rO4XWl7v7S1jLXXaVpA62w9OzqVVIbjYdauufJeyeidfZyUud
IqeBi4hdIiZlhPmyAjABzQ8zH8t9i7iwxc/geaEnYmVCGKDvJjDH/oDRPq4MQ/gVRbs7NZeLab4X
4CaI1ltgeKg7buc9bmIi6SQCcxWz01Wxi2JX2vwga2nLAfYViEJDSVaOsKYBGTfQNI5hUCJM9v0N
lucKEpZvapI7WKkVqSqG97M95trleAQ/QzXAnrzjswmljyw8cimOz/nH3wX2ao15prFFe4Ml7F+j
CCzQ73vVPR+tmoGDJlSI0yEzmGzXoXVTn0UqfM+rOFrtC8XQDVVC9EJ0Fnt5leWf34JZt9FFBXhV
hhosTsm9I2KD6HaiqtwpXAYCvl1wtbAmqsrEwtbaZ1j4YJg4yyyAeX992p9+fw6weqaZ7CN4/m41
LdE/xOMy8CyaSDdIaSWbxdV/fy7BZ4QU6EiJghOvaZczVyGDnN3KPIBCseZyhjhsL3suKR2bNrzo
lBTFwX80MCxNpeftgnBaIzG0K0XluD0jHcCx67w4dMgJXOdN4z76d6Hvg6z4FX2KaB9sfOcQxUxX
IkRuHyX7eLyz9S32N2XKhz9JlLnpYI7YPzxjhoBh/0CquqzsjtTB81z+/w4ron0GlpoSaqj0igpZ
jL4JJD2ALV3AqVOdHL1joGyieoy45qVIOCq22VOxixZL3tjNTzE0+imOoChhLJqegFkwnsiRe/qy
zp/yjZn29WPpLig0lT8uIVrACpwrDHkesWMpCYjO9Az2wZ/i8uDsbeU07jLc6VOA/9hGvToBUl0P
26vX5ImXoA5KZaTfWtKmuZUzk86FdQ4W73Yhqyr/viUL0yusGO44OHYH37/tQcvYsiYaaQgtR17g
yUP4uDN1yCbst7jYlmNcv3VBA1c0TIoNcEutK/469pJcanT9nRW1s2La1RNZ+cX+HnYa+5eNE5b/
MbOZPoMyjczWHiG4cArvOZBiVIU7+sQdN8pKM8W9Vl6y4T7xTBZXdoIVTg0i04enPXXaG9zhsy/j
IZtY9aJXilcf5/JPVXazWNTHKl9nQ1x7yOy7bdLMZYzIcW5Q6ekWAUp1A5fWcQ3hP4u0+TwXdJSl
UBr+c8XwJfaC4IoAlw1mp/mSSZuMGGjKr6HkXqBAHn1wEtwehQc27HUwpymTGBClUJcgAspufch4
49TEe0NKp0dBt1OfWtOUxVvJ0Krt7K7XDVJ2Is5ly2BKA0YtkytydOCNUr2fMtMsD21oJpJYOxhg
IRDELspupP0nfSUqU2C4v9+3j0t4WU5NDXMZJodmbDs0ZRSH/8yynf/Cq/R5iB96khdI1IPLuDeR
chp23fZk1v4gPacnrY6Qj1ebFAVqZEVXWtgUB4Gi9PSm60pz98TmyzT+dVYrduDSvff5rmL/Ukxs
Yo7SBJtmyOeQ5P+GwPLKPbdnpAt+ru/1dF1wcReDIzU04QjIH5wkb691Ci/Zh9IEsK3i3RLqozbZ
4qSijnhh9o26ikUC9HpXibTTGgJTMs1ww+O2ykm2n+tycQIaQgkFdvxxek1zZa0eS5FuSZ7ZhFLE
IQaou02JLvaJqQcJcbrukfnrDyVjkjyo5Sso0dLf7ujmahKSR6TqkL0VXvMZoMrJ/hHPODdGqEaC
J6fLsljTYfb9ml6HZXOhhtugojrtPETKVPSeUkkm8TYFTm53ry7Ku6nCSA0GrDeFLpe1RUSjqLX/
lgeKFS4PjG8aytNWdgva/BiW4RpMtGNdXmoLHzyadOZoB6MhQx39QfyjmiZ8SVy58tKnpriWFDrv
C/9T146CMD14lJ0PcCDnR8i0V10qsXdvsGaVx8D/0cxwjKTGAfqfbwdPliAtE9gQmxd9KaBMnPzP
So6Jrn+pilODkIovcSrtFEYbWhAbXFATnrku+N1duSWkkO0Zw9faL8E6woPcd7uF8hdRqAmsPxop
5F5671HdxCa4P3P5lOhlI8QiEX3czYUHAR9oF9Of4rK3nGRwaYXh7zIO0WR16Hi8GN9KeEFrwNHD
ER/yQEJd3tQ4JLtILb7D25L8V3ju41jwpG/tT4uFPihnlQDKcFqoiN49KF97WksM98qiIva7B7n5
66MfbdYj9qbNr74J8e/H8EPe1Hll83UHhAJVysxdQ1j8uvjQqnF2zvFWGClfkrVvaBU6hMNcv7+s
VYwBYcfuuO/KG9XH8DEQswCTznzyB5MO76l6Jb5ADqpbgaUExw/nMLA/Ue3olRTRny0kNeKxQe5d
0XI9QLm1kpdyXozph+QgbhV/DGSIgPqK4Zj2rvyPgcgjtXqGzjUpF4Sn3tKIGiWU1yksLqu6yxNC
3TPixb990BzakHke9rAi6bEvDXgnvdtXaX2zyNZt0cbw0BEMziRbLqbdEfD0jSYh1dk4xR9Cm8VQ
gWfZfj6nMaHFDwnP0K/+jryfwDpPkr/Uebp41rdGw2eBHTlEQMV/0Wq71UAsSKkljmdk2DpJSzdJ
wLG+yb97uYUI8F92TCvcSxLJEBwnoOix0E5Ln4XSjN8ioBikFSr390vWotLCgEYwYYxl8S9fs6HM
rehDfpK+dwGWAxQYXA5OjMSXRJ/F6z0clF7E4FQOUk/Vw56R7l9hiVX3ref8ix8BwCLxzDZjIzyd
GpqYBol43dWuVLkhPQWPGGDVwcnquZ/2fGF4+i8ciEJgwzjt4PgzYZZ/mqnmgdYoqIdh2P5n/i5o
2lgq7ySD2PHgMBpTAEYO4WMViqSGs75FTA4BmD2EK4bOYUfUyU04p6RXt6y1FCL9eCdfdECnGxC+
2HlulNPsegtTYw1aUY0fDCScnljBlA+4B3hdNqAQqSz5pYdeprKr8V8c/Tf7j1tNNpZqc2ThD6oH
L3Hyqasz5NjxIWFjFqPt3SC12BhNU4Cd5jPReCNYTjOn0NtD8+cTG39Q2TBNwaF57pdnmGReO1/E
mTicExfow9q3ZRpdyIXDkCSFU+7smu413ZcO8rDj1cx15+iAnp3DhjWDXvruiXlyJEdRFWSaNilk
zrsUofplLVgu+FllV9iCot2ImAL3GS7TWhxwC44LI67ZHfTyq2RKuB877hpJUoiHPcFYWKh5JmGL
/70c7tElGvuWmL2So+B9mai8IHj+jWEcgK8iJww3TsWxX3qhA9ElNO7RQUsBZ/tC76BxY7aqpXfs
ST5hoe7FpMVKfhuDmbXMDly6voZRQDy8yKH1GaNUFmfA5qFNlH9Nl4G1wefmiB5OyaRzhgTkdikC
zDfIDubIVw2ekW3EDaaAKB9hZ+7uV9fC3EELFUx336Xf2Q3sn8Lovf40n47O9jIZMy6anvPcLVF/
Jf23qEMzzvElWMFPF1pa0nU27Iz+24v6zxPXPva25AqQQtnvpvYMYzcHgSUoYXw5X4sfrx6qluYv
9j+0hhg3LRU6QIhniixcGumvkEkPFGHTGi7NEnsneekcTv81Peuu+M47y8ENNO9jtLtrK2e+Ygo8
cFLU2h5FGmlk39+AHKQRi/BQAC4HnRlgPtiKca+5WU4HxztiB0i/IP7BGXF5U7YD1sAXPsO8jrX5
/gdfJ8RH4NjMH6lhz34C5ffBrSGf5yvm3UtYO89rD7kFzMKoY0ORdP7cpPW67qlNpmVeRp0oyLBF
UoBkQ5renW3mviqB89ZD8nUoe+dtTinKgH+cnb7SuSQefHrpKOBamxFstZsHbHr/bVEGq8q6O2yL
P1lX57kJ0XRFqj0CeENnVkS5QrE/V1zyZIILmEL0WQPv5Tm+C8xmmgMP1GaQGSGNnu3A+U9Pde+v
dFi/FwNXVirpZZgH8uS2IW/x3S9aA2wnf8Ldqqe9LVZ0g0dXYFzIjLnEcItn3H77zfEgeC1LM6Po
FjtG7+YIrAzBO7fP67SO9LO6uuZW9y7h30DitBkLv+/aIQUIhf4EOg4JtudNbf5/Q8e4JksRcz5Y
PyhSETC8ZvUB2zhGuqL3Nc8HVVaWhp+9y+qqpwZLOZ0w5PjpGLnleWjTbaleZ1F0iQ94D1I5T7XZ
oKladfOa2JzuBVQLlC3xB5f1lFNPaBFtaM8FSi6wS/EajIVDKW4WnnJ7w0vu4OzqaLtJThJ+V+If
HiMWZJ+wKvY/1B2nKoBROHafyMyTI+2F0oJ9IKfGV/mHr15Gcld4YX3htjMPUKZ4b+ZG73KU5aJn
r+LADKzX/AMdw4AXjBahA8ydmtoi5GkeASxsp5YzrTx9leD5HjEZU9IndWR3TI/W66VHF4tDumHg
Ju5S2XH8zT1Z5t5HSCEyeh8Gl5JV8AL0jrbRfapkaQzjg2wHmKOc8m5gfQoZCn+WAAFgTsjPnPzh
IAXWjIwwVd6NejSiIEMcDK2+QJj+Q+39dbxii39uquWOS+qTf8z0b2tA65/j2rNKMBcCXqzVFnKT
p9LuciQDIUUKg0virKRJNI/uLmF3FgZkbO6Xl+Ym9WJSA/wdzvCjM7vd0o6fecuxCt9mZkMbFYjM
259poARlEt+ipHNouooiknNkIV3lgpxUIexxRlgXe/C5dXy2W0M6Yfk7lL+spKhGtSJIgGoPBg0B
gnj0MbfKugVWzpaO1/uT16RaaH+Em/o5oo9modbGtZ8/PnOPgzwWEV4XS/D2IjpHIfAm7Q/ZHFec
9E+D2gEWvcGaYVOqU7XqkmneTpmvEcs27eGFVSM6Q4JpgERvWmL3///NrGXQjkKqpUKuLlvjLS+/
Zf+DDKgs6Vq+jo7mZCoDtDvHQ4bfgRqpd5TnLu+n1KhOonrRsySKHBvkVc90Vtqbd4ar0Rki8Rst
jJO3CElxU+XDMbN99z6Nb+Cb/kQcrymPwx7S1WLxD1ycVuYD0/ML+RA2trzw+KsAhWv7G5gCWSrF
hAcjGyQtfF07pL7fHoIqIJKHZRWcMo6uoDS/vS9qm+yY98LAF++9h4mdyKW7bd2MAFkIkGo6uzIU
Jvb1qaKHG9ETn+BwMYHlS3afhCFCv4+hyNml38o8R66UeIUkstX2JrlUcRrbMsl7/kGNQRzWapS3
roMaHOc5oFJa+x89Zi/zbOMLFnBBdmppT+1KDrIAEwryZ1dshd/HpWDa2RhOfZbBktsbWgQu1vj5
hZQ+PFw6J3Ylo+Fq2ccQIxrvhKh2QGj1jr005G9fApcpWzXirzWBSRbaFWyHVBwCbabpFJTHMWzZ
geaItbcSH2fmhgHUtt4tLRdY3C5xg0xTGnB1/Fzg7fMcMLtrTLArZ/HlJ2R2LVZl7jw00R4ZYhK3
86BFfHFDr5dsmn2CYRcBionqZ6zzcErHX5XD8bY6B/b0IyNsBJzztgHsa9SoOwjbeGugRerMd/Mv
G3v+FobkhFzvKqt6HFzJaCJorx1jdixlfUhAnAQIp0x2eHTNgkdXhBUDgaTvTWKgyCs4Y3GqYYwi
HXByVGfOf/uyejYqXeyvu5FQYbv+KuUE2sctH0zkbWsJkrE86Qn5qAjwuOVhyJng08f8lXVRMPyG
1F/Karn2ZQmHa6YSW3cgOXsjmioA/WX6i64zgZiDeFYeDKOGiz9bXobzCQNiWFDd6hv7gFrUCZgK
UxW0tUKOpOHJR69xtpfRfDKdbJLoGE5HCaxeF6lYhB119JcN5JX8L6gziJzZ9wmZ2f5kee8nCUFu
cD4fB2GBMBv0kK1dlzAb0TdW7m7QpBgvnwKq/Ecg07GxDejq07sXwItqUrpRwnIRTHehIMOYGn1a
44QnC79zCxGsvdiB/jFXyb/2pXreWSnNRPlEDLCqKyS/uex85u7OeNLf7RiTEC7Wqfjf2IkmrQOR
tEa5r0+mO6DAmjL98oPCxp095dw95tRYPfy6AOKwu7ifNJV5hLDQ2TWASBuyBthBDieeLti4gRFr
gZvQmi1rz2K9J4/cKpUSBLg3vXrScLE8hXeP07Y4d87q7jGcdjO5+LcdIrArXu+bcftY3gA7k0SB
g9PiGwjf2SNYfy7sYf24eKfoyrncJ96hkozWbvhWpz71wcEuKaQv/axhQnnWVIU9H3u/leQ+llOV
IDFdBqiknQWJ0tSJWb0qBeI3U1U8tyuGEPjZuNsOPQHIAbYy0y67yiTZaKKT9Bdufow6nOVBAKJa
B4UlUxH6mA2PPmT0BYq4byklwLKcHC+NnikfsDFKWOdNJ7eotZEQ+zohuGaCDzkfybWhjUjOdtxL
UorfN0ok4BtoO/qGkCTBXD6lnBVctCZOTjop6zL1vcZWHhrHM1IlWb1GUOsb6BMuuZ0pBbY+sP6X
tx6FC1mfe1J39mTcDN7xD2gmFUenqojTxQPlEKB4Pwn+AqHsKxU3l6VmnnvTYY3uNiMC47FCSNMF
xRFX0f08tuz7O9/NaZVjtbTSOAqRZ/Ne0WUH0J/q4o0aPRpsQrctUWrA1WKJ9GQPulvu6L1bOIZU
pM4KgbjZJVCWqEDWvOGfDVzL2ji/96zhK2hvzi31tnktMTS8vYyTfFkAS7VjDgniDJzPvoABg3vR
03OgfrwdN7Jcy5TNr+FUa4JUxLroDhirkCJTIbZ+WAtsuV4+RKZJOI86uFHWygJ2RrE50C3U4kET
bZUscC6QNWRyt8pQrk/S4yctxhYzJotYpz7oaBKlBvQcnlz+kSWT1x1d2eNHqbpGp2JlRkW4XbNt
Rb1oFf0JBayoNdHafO2nrcDv0XLnmzomwzz5BuCfP5QshZnXQBCsV+6q2ZSgdNcjJbQeZgl9jxOG
AwHxqRXf7uf3vlyPlh0a5HfWG5cgr7FpW1bpQ1G2uWVRsSteGuPYQY3cmv0wjOTyg1KucyUBNwvM
kxnqnF0zTWb0QYGZPQjZ4Nw8kmoCiCYemPkRb9aJxyKl4pBryGUm2oO4RPSg6kP/JCL2PJGtAILy
EM6LG4eokbVWEYWpthp9zPVM8p8R9ubNzGLoqzZuu792fsBQFFZoTwUPJy1K5bimtKMbFgevdqcZ
3jXZcI9cSp+PjIdmZGMnf7Gv4bI5MojOdgKd2c3ufYVqh1BX3ZTzs85knALx0SJOljvM+paPSRgg
bmsnv0TkhfiDKnnkv5JKXz+VNTbBaAWcCwsnb7VFBZm6trrg1EKNWHG8nD5d2jguxqvtub5gYwqg
ViWoeKj0dXAQ2Q7B6WbQ7K3k8slXdL8KWnEida2MilSwtzQNYcfsR9VDrbDzoDZ4U74qlWsoI/Sp
hz/0r+E80695p1eZoI0DTXteBei/4TFrRuxnKb1+7QoxwOnHEbGuJnRINfsKoU1TWOJt10Lz17qs
dGRWOT/ZsXsbbSMUZiwS+f6KmQYbhvlW5TEH9eNmxHQ4M2rTpwOBqcOMLWteS+RXSXLxlDSaO47I
nPjcDL3cJ8hRHUFhe2tIl8PMThskJC3ejGZLbbX75a6Mr9Qp6KDgzly2nh69R4tyuZOloszP4DHl
AU2y4sAhjM+qlSHYRNGYOECqd4O7a4NdiNo0GZeuTPpn63ZzQWtmZO3rfwQK2l0naFE/6UJSED1T
zMm+268jKEdmPl4aBAReUG+ZZ1oi09Ugi8WEIXo7h+nE00GA4fdMrSddxOQUefhtARZDwmlrF6Ct
Mdx/TXaZHKGY9JXTdV2XJ/HRsh+mY3VBFhwI47TUnFmCHwjaXm5yIv/rew9F7qLizwaqvgE7dIDf
0jrQ9a5LNnVeWwyOwkeS7gYIbWGQi+TflM90zU3l7JaHHXgTVqEgBTU+DkU8CurfAiJQoHNlzxEi
Dc/3eUVHRkPWeh+BV3BpIaas3Qu+i68FzTHXVKgCu1xxAB1WvNiI8BuBA50dsXtFH+dnXE+Bhtwp
092qXkdkrl2kY5JWBbt4epuqHJd+AssQDJ01HFo8x1OMvHw9jPW8UkXjmhngwlCRu4rnFiFnkLDQ
jOxvF6kNlTV/l6d0WuWSxoDDz6NGtRngbKZxf8uVAKO6F0ou135otaSRanlFAgce8MbfiOMg83ca
T5ajX2G91gOueWyRoPVUeTQAekx2CN5wY9nMVeaoUzx/eSzEoDjZHp8NGvqCJ/o3YeIUEgWsP7mP
dUytEq6y9UAUf/5rBQt72Sbrjb5XFCcmTIrEOO2Fc002clb/UjpWWjQzuNU1vM2SNJH3b406QQRh
fzKsX25ez7wswdocfGuXY+0nGVJLviIiniF3OBfHyxk4u7YD7hJvTBmPpnS2Tw6D8zLAVPhP9snd
F2cwEAmv/7k/vbhoL5f35l3HSYH7C7AYv4GtU4zbUr/G+YC5JTB6ClMt7sKVqpIJ9RYylH8pMQ7T
eCnMFhKuwxCav+5Jcqn9AYnhkdwwZ3uFg12m2iae/A2jYNwjN+ibN69dXEUuEQs2rAStPS9begBx
SKFvmNPBRhKNgt7okE93M0Rc8m8Zw55e7jjAvfLVn4mH6jUNsq4Sd8nWLm0n1POnfEKT3eQM3QWp
8j/h721ZbJBB83yLRxMzH5ekmMwoz3VodWBHk4GQGkkJvoGyhRIbR+t1qlaNA1ivXOK0XD2Re5kA
qn/OHNtk/f+njHFprOzLBFMME8PwBfOWwPlZ5HJwHBh7gvXNsMIbaz1WTEYOJWVFKFAmkqV5IqXt
YMUUXQv93fyNQyapeJTPen8YSjNORwMH4+749nHAAuvMeNxBy8w2sNcLu5sVP3Rc913A4C1X513O
hmp15PxjtuqWF3Xf2uC02orNH3MrSepmWKBrNPMSamuwwJ1dsY0PaaOj6t4s1rWfhl5Df1GAe/kO
Zn66jGleAqIIIZMvS/anFag1t8VNCEBgjUrY7mSqUOt84zRTteKLaeB4OAHCcxSMLK7Z0z3k3Pcc
WWKNCcCahAFAh87seuZoWV/ItmU/+hKrYk1uHuTDmrkQoijLNfU55mAiiUCl+1mdvi5ol4tAaCQx
3zFDt10NwOUU6VTr06Uuqg9m8bd8EbLNem+r1M8M4Ilc3Hnjj00irPUOluBxavgsTdAGsmdQ5RNG
dpUMp7lk5ndD6kjlBDnhIYxqfvciPep6REI4J417E0mv6npAlW+c39bgNmEJsk12ziGutxznxW6u
NWrt8TsxjBzE26EoXrts4tWuJPv3EYTql7P5dXUWgI9sNbITigre6iE6ZQ6J/cBwo7MpPTyWIDnG
GNCaeHbUqTZuoX+/znP7k57s9ErDceGJqMTzlo440DWuMgDIPwkyAD/mIp5Pco2/uhqdolSXCPxG
+bRe3g1IB0WEI6qzbMX4DtcaB27P3+IR0yeqgV1/OTwZkPL0kCeDOQn5Er88rqX687RgJqWbnXsN
V1Ct8u3ghLqexjCm/4l5uzT+2phYjW7YTF5qf/ZCT731u59P78R3JprbeVyPwqKtOPmgG8/T8EkR
S4LGw5Q3C9W1JSyjSyl02QGnYCmQuShSKEYe9/mkZ+nDdWVK1A6G2OAavEhG/RUjrJgzJCSVcvJG
eBfvcrtMotXmfuTSWkxJXyUdKBE9I/fkDT78H486yqhSAk2Df8VCMlNvunSY6GhlCupnzRk8fu4V
WUdDg7KwF2m0EHCpYmkz7xCoyvbSMVt/NBqk5zA2njWDUXvIYBOPsiKZBaQ98KdCNecwZxXDi51f
B/yOxKR3nBgxp1HjzfRGkue6uMRKmn9UoFPSN+/ECr/P7U8yiWjTPHPdBtQDIAuJ93iVM9YxXpsR
LlWDgLdBFl0YAWIfs+4FlEhPlXI7aHMyDnte+Af291zDiT7O5ZKOa/GpKGht64ilaNTXb8n8uqIs
QIg6cjEQJfpnV5qAN0lcA0mtfQobSTNJL6TF9b9PJzFfw9fKvzcTIHCJXCfzkJnqg0tepmcvFEjX
u7S1J4Qk7noHrBXTuwYbz2szZ0amenUhqj7O8szaSFRjKyHlZ/nrOp7I1uY+OfJl8mR7n9eMJpv+
/8DwRGmWKmb2rB3zTRfCokYIICU9YY0RhC11fg7VrV5fQDaF4UfQ9ce7lUStWqI1GQyRO8diOaXP
kRvTS9LV6g96kH19lToMxL1uoXfTpllcBDSkt0cWJLwLLZd7xRDTvK+XTe/fBsk6orZakJZjmKM1
fLx4E/OZsOkATpZGASpPwHSzzwuxnLamMp2eTCVg+rTGZwGJmS5Mzx+l9TpMxNECLDgdc3uQyqvO
vvDHqxpFXTpNoLM7jrHATpvnDi3wcElMqid9466MSTUGlSL7Ww5ib5IYUcOCrazNtB0WgV4Q0bbf
6aJ/nXUjDk1AAJ6N1B9zZmhGQBWYKGXvOuyjYk5fbQpfsAbv8FdsY3dKzj8FHRdjQPzucchXw3Bd
TpGNHUFwtq1icqEdpI0amQ+KeWlrTHqYEt/Jl6QTrgqx/bFTOVJgDHDhp7fA2P/bCBnjkeyrMPe+
KijEsoyGJl+JUnbgnLt9A+TAv+wKubmrhAEvl3h0J+GmKxpF/FsW1kmx0E+o6fqGc5JvJZK40nA3
weAnD/bKApkvnY+vM9xhxsuq+G1UE/Vicq/wY+x3/Ug8ncmZ1zZ60YJoJ38pjO3iCE8qqTM9MVj0
FUqUnz24AfQMyKM/tqsLl1AuAdrlEut7syDH7uP9NzQFRkG7G8kr21hdaeohJ8ByjvJGGuL3U6ok
7C+C5OPIQTzBIcFzxHaoJV/08VJDCCmerYUwqhlB7r0ypZPxKTfDHO71NMPQ/jPoHrQwO7C+KPDh
mAUODow8Z/6h0KGBd+Ey2a+4Kfb2V5vq35ga77b2TSBVuBzNGdTJiXKWFUpjHLYC1sEyahPBIgSS
vAqPv+gPvHiHfHxZ6CHb6A/Vgjya5amz9TuNzoaliyLOcKa/OHGpwv5KuIkxR4ZT9z2/co2WAyz/
HQCq0FHhsfi57qpXj59MBB95Ze4xschGS1YYHFZni3Oa4pMFNTUOucUkXttrp8vbp1OMrBMvf49c
WZIwDb8+C2tvi0XnFHdUp5v5Dgm964mHCt1en5pyIyUb51C3nniUwiwQR6/3cLjiLyeIied1MSEw
OeC9O+I7XnIUa7WiWU1FK7R7e+ViqeQsfu4s7cbXiJ4RGFGkBroySJuubNfTz0yDvWadf8n3+z5l
/bax64id2LmY37EMEIxEHWFPgI20ulGyobklqZgum0kuZ3q6SFlWXMhCKOxuO5TKIa6NX78m4P66
v5+MLmN8R+T+xyqluaBME4RmYbe9sJtaUbQbwJdNG6DXaU2smRxHJ5un8j4eBJSzq4HbNvm39Ln+
INxhzEHo5qzbtJHqqkGXOVnABzLmoOKY9bZLD+HiW+WErVoyZkiOrAww+eDzdi3985KbAabK2fuE
Bc7gbugM0KLIH/cWzF83Lhg98M8A6v79j+mOGtyMIq43uc/LKi3Xp26gPrPdYPjmOMCWU9zuS51E
3IqSS17/GopRUpKT2w9JxjoDrgKIIBb4aBoXm9Z9OWCx9WsKze54dmCLQwFlEp7gpAk15u+Y8Hpj
dPA/INMN02NMVcCsAf97lNsLiqLSQL7m8/snevquvZ9U9C1AZ0uV6lIbMqE25l7X7qhEIUtmAmrP
K925zltlb2L2e1CACrO79bsQ8MviGjr66UGDU+uZIShiMlqEunDGc3FJElrtDrL0V21vo0IfyBDV
YpaaMb1fKUailj7iOhOdfauvWpFpTyY9jwXODUTk6aVELKc7xQSejWae4HHUP1utKDs7/8d6p28C
TtMrSIfgVl7MnZqkfHoFte95h+Wmh+uusxVaY2SSc1Hpi+7XsDqWjsBNO0BZWiztSd1f4LL3GQ/l
7/lPjBoAVWhfCZ7lAcisRQOsYckzSu4zQyiCyVuYN61t0HgXVb449jhwPqZNY2ov6PNshAizdhd0
boVAx6Jk7Y9IiDXBzqDoebrkM8go9GcL4xAeJE6IaB55Np4cy/tCNgmmbcZhRgsvQLhd5WCsh+U/
IaoHQtcR64UgDE9iGVPN1wkJqv3ELwrEpHn5ED6CPlAIFyIALWiN68lXxikPN7bdgx5DghihYg0Y
RYBpWzzTuV7pkyqpPEbQ4Cj92MN37T7P/c5TTwbHPoBzLYzqNc4Cq93nhRPVfFDADQm/zjzLcZjx
heO/ouShIOrn5eimcgm6BR6poBGVVfkdLYNhGZmFEtfwmLa0kOT7v1NvYm8ZYLUXqSkPymSm5TEp
hLmHk5e6A2YEvRgHTLx2etxYT1TechW7cHaloWyWhHpx8vZaCCR+3Xy3Ykjm9irKwyQ7ifHtJ5ct
9e8WKfT38ja7X5KwDexiv4lwoD1v4NYRTfnhludmDkk5mPo67FH3YhuUOrD3xPN1KgtLomTU5nRR
v61pFKamNRcPNW2PBj8o++AsSlxYaeKe4t01hXj23MWyfZkZUoN5in31kYnntwbUhxAktIe+73bE
9E+RZcFfwQF4+KmvTKwbOKNh9Cj6zruH01OuBYrD5G2eh05Xqq8UsU2dMyl7Cndb6BmQ/vle+hTw
jxEK3snUXKLRlQgDjK+mOCQHeD4GYtHNtTaO3QWroKBymsYz6+sUcmI5PtqZ+RPFMUPGnGZe2qi5
Nij1OryS/EOePfmfPxmBntRGHcOR4C6pLz+KxCcBO13oKHgRU3yws21Oe0Md1QfDrDM7+gD7OLhN
XsJF2vLsE7ptkkyOUAKAX6pCm4CLJhHZbHKAH6EwEURWbcssbtBvzB7OWwOCiiYiZoJ3DdCYMFbw
TSErSKPrtV5X5aniBqF9A+rzDPb5vvK32da6Goq+0dMAkwkT0yumfktO5NsFDEUzAx9HT6xoCR5l
ky1szso8XBOgsVlmjBNh5mrBXSb1K+YzCfHVsI5IMNQzeYV/PFc/sDRKGzqDbJXzsNXbZStIQiKI
0HLYo5sHFySpKQbMpz+SASn+cxZU9klRxn2sR834VsdO1LAn0xS4rAjkw7qKa5ohjsQpJTgCZ0cz
kHE5VkJTl2uNvuBTHT1AE48ocz6+vbaOe1opuOP3OmLHymsStTrF+SYfMZEXWtDdvAq8wXRaVsgX
22UmDZYhbz/d0nE2nWKsq3roeASnNrLdUvtFmI3+F0wLZMutAetCRYJDuxMab2NgTHyor5d8CMZl
TKgpobjU2zbQND1/cKls5aqnyB6hvjKg4Dlp4SnTcn+LeArtZP+pGkPEPE55zKSiAI4gOqiXY3G8
1tX54Ctml7znP+iRi8lM9LhcAzKTNm81lTI3WaZiFiYSckWwgfymcB6cipZRGjk4pM9rcXJNKMiF
hv41Gi3XeU7iNU3YaOm1Q9PMDeO6zS6xyN/K935tObEcjNGEqGXsj7lVTVON3hzIWOOHDA6QR2yz
G8EWjB2eaK2rplpWKIKlL+Fn5j+sMxsKLZH8NvunyF49Sw4CGUYCvKJD2V7CanD1ifwRgGSXksVQ
6hmRNyh9jsW49IDsiJV7HWsPqkMNsa8odtXAdMsZQWlSt+4tb5vzGrwSYW0CHfqsZdWnsNB56Xlz
6VXNCJviq+g3vyjZlIMcLumckg7WdcjX6iRCbKkvqNTzMG+xfUZeFF0VfmWANq9qoG34OKj3KShP
8kPw0LRRcawBx3QAMIoR3R98SSNDok9jdkLuELqdgyEYXSZcKzWEgeKygBHho8l+CP+rf1xVTWS5
g7hnuvk6avPEKE/+w9z45iEgihmdRdsPzkvyPKT1ztUxK/qEJ3IhqTXHfG1vPb7d0U/PDMjUtWoj
UHJ/6JxG5v74KCcsnpPGZ+GodrI9M4NmXAXjauJTYHQOivjipIgSTO9JbEwrRB9FnQ/02o8IBXXE
6U2wCUOUTy0znx84fdfr51IcjBIYexjfR9pRIPIiMmUUkCPTFUx4hfz3VxfSKdJrBZ9FLT87NibF
M1Maoj6vho6sVgOlE+/3VEcPebNUV7UX+Vi7M7np+W8xwluq9SM8aOLrVymubId/+twh0VaRdoNt
d6VPc94W4/8zDZDejkYKfuEdL7wBteXusMQifhfOA1xRVGhlycRCd0XGAym8My/H/IIOb2zxieSg
e1KvmhFN5SlL0LJ0+nb3Xl/ghUUVuPBGCZWUPRPGwe0kDWEISGaLsiZzfTbq7Ua2T9emQE042N3n
cTxs0n3ivDxCPCW6j12rBKzZfQxONvW0xQ1azxKbt9EO3sVxOOVikP2VeK+RDV2DKxWgf+ov/3/l
uw3tAG84357VCGzTliSfVT00Zvy6Y6TAqqyBB64eMyGJMWdLc4wCaNj4+9CwT7voNaREtUYPWCwY
lOfddID3RdnEZoRA+XTm9NJ2xQA7SAclHRMdTWh+eF6H4Q7nq17RZMBVrpV8uro332OXHv/W27bC
xF2qchC9v/lhiM2b1JNQm3dIaK3E3v6081JZElLDRqfhZ0uuxGPRBUxWLrQJWeKnQZOqlcnUdNYO
j5Tt1E250AfkAwMkVl/Ax3b7fMxt6T5j2V/FHBF5wl+tQzM8cHU7f0NfpsvgIacr1VK2nDqPfyqQ
m+xcAcgQmiOjRc3sT5fR+wvi38b7TGxBcKaecsnsNoYsDdmzPpdWRIsPEjExvvhQ87k1gKvyB3PN
VyHIalPG2TDWN2UfceJLbV1qgQo1cww1boVy4h4fterICPV4ip/iJGPq2NE7JXhwqhkJ0IMGxjTy
pShH7ho6MAWpRsVv/ZsLPw6461eikDYeP8TNOBksICtVBZenVLkKjVtg0VbATXxXBQ61HddsKW4A
rPX9WrFWKG7QKPDXMeQbqhOmkOiWPs66cNZjXikWBii4Oo4fSWhOynQDHfsLwBwoCKTuqLtqcdhG
Fjk6bbrvX0zv/W6E3X4QApFjQDZXzRqRZhf9Gp4xMXiwcohSIYja3yG7vkmpnzuQ5FknGu5Te5LT
5kMPalk1WFaxVrWsDHMQJDAlckmtTUXzpjZEQTYFbhNxVH5I3tueJHA6I0o5SMWM7Ir0H6jIruLE
jegLCF0a3IdepFUdWxoXUZGYwQe70gIiQ1xCs7RTB5b1udcPZrJnNP8lW7wiKk70/S6YOAvpmVnK
nf0+vWPwaKoBE4Yqj3ztg87n4Fq1u5VDF1BVpkU/u9OUulvPWZI0ujbdPa3g7/lZ+xoTCOIRoPdd
27eSjlH76M6GUf7gx6hQSPr5rZ7SYSyjt1Vx3C8wj4zV1Ds2/TTIC4XWin1N6CGEtn4FSfj6p70y
hYMdxlFuFR5FD0AaXlG67fhN1E48p1D/S1nz9gQlf8duoWUoOBz1BPIwA0rmwaOewRBtvkYOcjep
c790ACNv6gCCvoiwcNOqCu3viajrLpp3tvGSXdKETOPaEbmFfnOthNcvgg892matO2UUCyhRmoBe
HAMKK+i2GjhMbUcZ4iI8bmZkKWaWppaF+8R1kFUidZbLKcijDzOKbCBD7Inv6sChPhGLJkdegB4n
LdSJOpWsNQaEmfLnOitwtTklDp1d8WYrMg0jBf42QHMUsZ405XlTP8n+EHMN1nig1izixBIdCa8y
qB5LmHA4dYOqM97xe0ulePRU5hnUZ3rblQL6Z1kCPL+rS1BtLh7cPD0YpGb84JjrCiC3jA1RZ8ST
JeldZOQrooulmMJiGEEc0/b/22u4QZNEN3b0ANFWyQBAkdg0zb9B9lOKeO2gNWOJFpQtqA+wOFWZ
Qx+G6JDDkcH7gDVPhgrm6LqQ35BYPgn7dTwoVsM4dXl50pR111hAwn7UwzWGxswk3bnumtNC+zEM
i3AzgtF0lZKDclj2Q7MvuQ0wNGzh75/KSkiiXcjUx26KVpnrkVgMKVIXl+95QZaE7hW2KMAMGTGC
+l0ROa7Qbe7j0pKIHyUdnRmq9bgc11oc22ODKjzV7A5DHNLzF1pM9tWbdmVUqF3Y+p74I+nqTqn5
M6cxpv56aosJd3a67C1MfRQZAa5exeyjSwTN6CyGhL+/tEzRS3e++fwU20j7HuXqIZFGab+yhGlq
J4S2vSxqTSPRIGJTH9w2ox+CKogt3xfqCNM6+KKn5doM3XStqvDvtWbq3Gxu7zo276U9/CM91Y/3
H4HE5PhehdGCtZ9fp6xiX6ESVY9KCWfVusWcOnbnQfBeZKtj4oIPd7lgeLlpbgzWmHTA+RSyAkcP
g4A58sf4pF9E+IH3tFO9HE1cuBM5e42AJ7nfaTB3iHlbzUA/lBXUvBI5yWRV352SPQyv3OCU/xZ3
pvBK7+TagxPner1KL3PHmkWP5r1ciXEj2SYDxA+U5VSLiSwXjMX5i/5dpQOXaVwEty5Yp+3WGzXi
x3M805Ut89xCwlATKyd3Kqq3ntoIC8dGb0rSunWvTI/jImuiiuphFqwmt/Wn4gYVbxzqvoqvVqX5
xhfo4Gz5TNEwKeegcPnTeNksi6FrX4yA7HlNS2sLuU5oFK9E74sA8ElWv2JxaxYeNASNvTvGAcqM
LyBmoIbRWnn+7myw1i81o1MkrTPTnOjfdY/hYAYQ3hmP/eCya5W6fYsTICZvgaM7wUoVWa/NTvBf
/2bQQZFVFyd+2jNiEnnMUCrEWBSut16/OYIkk4I+g3/2K5FRcQGaoqLDEvmLPCznexqG5COrTczK
WuCHAxEkHScnG5xqAsm4uReYfQjADvqwRUhwpdWGJS0jvPVamlLYIbBCf3O43ByI7YI82FAi0lK0
8LKsvuI7vEJZ2X4bcdw/aQUjXVRdH9uaT9Y+DusRhQ76OAXBvFQeqxeP5WHYogJkao0BskktbivP
ep3PoEcquJvno3JthJHpBZXaWUAQbCbQTavhR0PpfTdvjY0LwvKUEL9TGUcBjL9LRkac4ACkP1dN
p3FcJ30cP5AgC9b4AOuvJzdhox9zgt+5lTzsGyVKL2Wz0ZZpQtgc/FY0jiTlk/DeFDGWARk2zbgO
tPfzPySMK/E9UOam0KrCuehzMDVZtWqcJQcx2eeFbKdW2r+Ha096OvLSMj1tAXbjJv5H9Z+WCJKY
1MKciNIBlhUIyZX0L5T1PxdccokoIJX1v3MlLJuV87lEZac2tQsAx0VuVFrYb8S3737FHiwmgTqZ
YGn/mHPuohak514s6vsIGF35PB6UnzzEY33h3lZ9XjV0+1Od1aJsg0QQtOt7FFe2of4gX8qNEPCG
eMVohW9Nq7bTz2Su/V3PGYKBejzEC+IhV/tf2uyc48ptEGWpYl/ii23TxnsHbfEXCuzu7qNVfyUD
cBzyywbQCc9vesXQw+FLtTsZ+JnQc9et/AdUBSS3YiB7SWstowwag5UJjv8QDMZwccZhccILwLwG
qEEYxHWAIBY2kiJT8oneVQ5Qz7lDXzte17kJ4xH/hMSgmKzeFEbXZVPRLeL8AMmLS1gPVmiTG9p/
oYi2RzjL3sndTIZO+d70UEZaffu6ZRqj7u49z0IlzJ69JRoYUSY7R7e61UkN7ccrVSqWtQ7cGk4k
6bRjvxfBa0HuUhHRjHbHDIfMSlDjpI2H/Tw6I/hUK3F8blRj1slgK7rdjk5GDfEQ6xiip8re2Xtl
SL+lDNTY5w7jcZtNu0HBh+4eLUkE+P3DpKUXPkTFCD28WE6X+u62p4r5NYEBhfHGskTFo6j/i1PK
C0NSJ//JwFBmnmZIIIkdd3PpMxyEEFnmkOFedfXI75BNrdo1shhIzaSVVTVv+8Hi5m804pbaijmf
/PhKhlZrG33jzEZsanfKat8zYgXCa3/P32FbddoCmRSqJZlonhfJZyA0J1X0VAKKsb4ELJHApY3u
jVEJTomVRHNB0EfEq1jJ5laJtvdEUVzzJ4a6u71eZ/eFaHMgMWnuwSThPXFl5ZPmQvxrW1PufrMy
jnLgMLCBmbrLi5FWNGBDqQXLtnKVK6xpxflZ00z3rppHcn1csl1Fkjdt2aygGwbqGmHuBE693oFJ
Z087ZlTOdOzHoZHGmDpKNpJKjtq5VVv7ZYkjnTE08QtOn7aEb5SEt4oOjC8au0lJpsr0IT8u0x2i
/q96vWrm6okucc4md+SRgUsQcCRMlTCT9+IUXYb8KCg36ul1l7ktp4hSjgBlPT3kRQ+Tm1PzNy7N
29gyaKRj2Z4BX+lrbecCcqCGj41WmVpb16qoqPMGYoqJQ+At2qaAQZYCUE+ylSjrfCM19L4790p6
vzcT6U7SG/q6r/tqIaG9wRULN0VRWRdm0Ypv6pay87qQUC9CXY5IdBd3bcgL+PFip4MVcSzyR9BB
Zq2U3qnyjk7X/1KLKUWw6cuXC0ggy6YN7e4lzED377jlJyS+KcgO7hDVjgWTF2uHLoq9BbV6tseF
VpXpcU9+g6xQKetg0H02yZkp/LNifWtd7Nx/L1T6J81yRWiY2TIMcie55L5yvpi5K0GyKDxWKqLg
xp+/Iy3B1aEkB7BhfCoJQY9fq5mxwNqrwAk6bl40VvKZAopkLDUQTPhLsmsQkzIjnvxUEzh6j01u
7r5IT3v0dptCloVihuterGBkFKPbzTkCSAeN4g6G2tNs9xpL4S1cd6bnkr7gJtYzs8FSdXtkZbE+
5XjJ3zSpDF0fyP0zaYMyVsogy551YOrQPR0eCkIdFkOoYuwql3bM43DTGKlDBGn3CqT4giLYajvj
oz2KmBuS5yxSxkKPAWYJ4wAaxi0nr4bs7bvetqwL2KCuKlBcWcTvMI/vv6IUzAK0ey/JNBEqw8p/
UYmcU0cRg5p4wL8t79IvmzvXs8NAfi7PqjjfAT0YNJu093jTSHO7Ug3e00XBhrz7/52NMKseRRBx
T/b+De+IMuxsGHWa6CGcOw3CaZu0gNaK+idKpCbg3OK1uyGIJMdeYJj6YteMoD/Ql78vASizNAz0
7yNya+5YOP8JI/I2H1PbgEZWr/QozR7j3tzkrZ9CW+3FdaCxWqybqMoVAVjgLm0yqkynMtl8OJVU
0kxIHmvB9VpN9HjPauLrSH/aXadDG7VF95H7bic/5hy4Bze6VwtMrY1MSKSr5GA31ZgVzsuwPYdb
nR12KcKZqmoria/Hj37OfMlPVdXtvuM5UqFYHBRuLwV+xUMTACRlvmmbYt/+AQc2ChjRJXQw+U/J
FJu9PhZNwQGNLIEbZCg0joYPUKNKA56+gtPV+GRCro4OpTdY1rv//UtZZAaMOHsO3aWOgiqtWHYj
ZVN5GaqdqAG6NF7zlUIU7Ki9HpjAAauQ87pZqG2Z46CBdZCHyGk1ZDtY1GrHHG+E3d/DD9hYU4YE
X/13P49SsrcPAqmFveD4ebMf6zadJ0l6HWeJn5Z+sta6+VdIybqx7gg2aSliPJ0fujZV7YDCNS0l
UA2iNfnrYqQeuzzXxvK921Wdi+O+C+AEeXNmRQJmL9WhLhXtLghPkKS2nE9rlOdzMlpnCOBY0OTJ
cCoIrSvqH6c7Q7Ce4vdC2q7uqRve8brdBSn3nV2QrPCQZ/apRby3Z+bKbWsGCcYaR5Pv8qG/BSYk
4ZhZczoeUQimjEOGO0uu40aXzFvHWUQ2Og+cVrwHg39UCyCfDJ+Pgk0SSkY23gQ0aLhPdLJmp/8I
42U22VjtMXwZzCANlrLlwxsXu2M7mX4gpH25DJYlgDaQuAcbpG8waj00K6+V3MsYxr5cL2rLBqZm
XGwIjAqF4ZcqEs2TscMnnsvWXZKG7/7NTKlAX1RAJ2Q6NWutFAE+3LXCJJ5royP0CmO4r2rkWNyf
dgJZ0jlm9XXG6iToTLvrgSiW5LvbQN0cbLGqB3sR0LkU+YpLTtxcxWzOuIvkggpixhWLPfDsLizI
mvidSd7fQ+UBIwOKv7cJMvzaZiDZCy2QBwPR9vSf/DMMGXutmTVBtkzlDCjEE9lbINQDUBbjgzTu
WVWqmlQY3ClnF5LPRPrLO/C4G6Ki5aUQaYLfob43/wpScAj1uFOsEj0oLhNrYj5KQ+hE3G3k3O7q
6VJMPDyaj0rsG7AGUYuPg1Z/vdpRP2T7GEZ/eQSLAulqqV56bMit1hbdE8qqv9CJgtjVE+H5/m3E
qLC/ai2zNgwj8C4qH2NDM9ujB4pJQqCwCw+SJHmuWaCHB8NKGLlJ00mrhqyrnHvzn+lPSxO5mobD
WJqG3k14tyoQcQX2/aHkz+Mc3dAZz62m+FSteUOOuYsrgIHatTmlA+VUvTfQH6NlmmnI86v5inqn
vewiHRhk8GHAJXXx3OQHM2D2Hsnb0WhP2MuXDPQz53cWicgxf8bmydkFCxHSIKM/u57WAo52uzI/
jIe6XnTVChJ/TYKFdZihPz7oAdXm5/t/kNMG6/nSbqxlLg2vS5qghbIFxxJGDnWBqsVBvn5uf4CW
gLkeNSlvrttvfD3JKGivlWT6RL9Lp/UmsIt/8az5clevEWTWDXrK2prJINZPH8tBPclixvgeHaa8
5k4xUMQ8a6zFrLAy0ujjbkKpqmpouQc3K9he671Gq89NDvN9bCBVPDfjn9R5XfLJoyWzqFlcG9xn
jGdWMG4pUwmXedHytnxJXHpJ6qqIfSUc2MfsuokXm/G2a9bt098pgfYqbF4YPYYF4q/2eoOKPaw9
/RZkCr7BPkfTudPZDtZeZlA3r/V8sv8EbANHGNyahJR2cb2ZGjsyl6j+Bu0DZywq6YKs1OvxW5pp
eDvD/4a4yZK7G33wobuxlQA0Hij+w0x3JgI39Lncwbo8AQy8IwZhAwbHpg6IDsKwS7G7lIrEv3pj
/zY+rz8tKByNR27wwPimR4TeZ1dmi+G8aYeiknFHQIz4dcHFx3MopjJpAplDczC4MUrFYIMZ0xKa
b/2FdgNUBTLFk44d28HsbAqC4CEVHL0DWJfuILwXTQy8WfvnPthFrCkxAT5ENlvr46BPi+SLxtcP
7nOB1TF7ZyCZT8zbYs2tj3gJtP5ldj1O7c5fy6xUsK95P0b/TElP3SfmLogTKcnBXXrOGFEsSDnN
/JdF6Dhy7ajbjfanbP6QTA8pPLKxF2d/aK2fUr8STafW1sTaIcVKtncB1holOIcqCmZuqlfth2w/
RZELJ7/ML4Th08CYZUjz83ac+OlFGk7En1T46Aa5bKHLcT9cDLmjCOp4E92MLSSNs1Zd9p4le+si
r4XaZ9sLo3H/NSMKtrPxLC8j4Z4VzYt2V5WlPdhaBbQPw6Wtt8COF7sy3KNPuQKt744YsJFd11u9
kURzprdmvarPUEbd4q7pVkl65X5rz3yYddhm0kLIuP83nYcGn5Yualat8VHpJDaX3zE8Fp8Yl662
rm73WPBQ1r0ZxD+G2H/gGbaSkgrgoYHxAWX0V83Jn6PZdG7o7g8IRL4ujEFdYn9xh4SanDqbviDF
6avHeOz/uPWGy+r7oLBRpEsIb6ZZwv8TrNZtDFiWVacLQPrKxRt9DKlu51L0U4YY5zFhw8FLXXY1
8VofQXXqUIWf/bT5o9koskb8T6KZa/CTL6VYXmu4EQXJd8bOBwwshP90WsPrrIjZRcZBNvh5V/sb
a5eVnooX4XyJVig1WZMWA6SowNw+TPqgrSPz7UQaAhnas0B5hjWB6UyPYUn9hmPA1ujVom1ftWzv
OY4Uzuq0sb4nKWHJ6s++BrHq5mbDL1z6DqRnOl1/RhTBw/vR8O29+p+1I6LgitzoF1PGi6d3kJa/
zGx8pK/YF5tJ1noBctyyVvVEhkzDMAkYlANqE11gYSH7sFkIfepS9oRidZO/JDSG5aDfEtkkTiu1
U48MgrL1M+w9Bgrq/LNfCxN5WSHHlec++vac3CFABwIVW0Vk8F4Wxi70EttEVpNgpD0smSoChqmQ
xa5FgaLe+Nxq85q8k7YOeFp+qi+yolLc3usPRwjMhyCa6g+TtKJAkanNuflqYdZMZ8/fSkpjZucc
DQffm9cb6HV/sfTny/554Arc2XIV17uZ5eWdRdHp6CRH1DRvv+9JqwG66BVWzNaOCKrs3sz9l9He
XC+J6ovJI/13R/jXcr/uZ7NL5mKD63y8NWAdtEU2CFHiBH+3LdMXaMxAHi5bp1RCnugQZIzxfRY3
V+i86q8NI6tAlGyiIYXCXDcDOegkGqRG1CIronVEIBhKiJN/l5l2usHqthPWbeaCdene9HKzdjfc
QoIWJ77equ+XbqH5RGI0WeXdPRysvTVDdvV7RC0GPiiB+5t6JKMjr9r8CAVkydrPmT6v827Kp+xV
ivaEoETWL8SSGESH5lcNujZVkbMy6gWmRBaCr4JrwrMuALmw7QX0jBPVcY5PLyAuJtutD51XviWU
6zQuNEtY0JAmdj0NmLagcSNlKH+bH1TWoBM9vyEs9nGITxg90TAucJDAIfePTjlVq+rs6ZLnJZ+8
yu4JnnBVlXr88RbtLiH+ZNAkJjCfSskuDRtWrbeV5n+g8sBgyISyPsXSfNh2+PCTEul5h3wi/0ZD
zO9DAf0SAkMs2zzIjyojOxJtN4mwMB/D6Y2EZDTbKzZlkW2KErZE0WOq+1c72PKqwItCs7wxK8Ow
OkGgRxszKutpBHsi2y6Ry0k9UvkCBfbRUhQngsFtGHiVvZkmJtr5rusQxHeb4UYhi6gE++uP+xlF
a0QmbssdD/K5amtV3/OqU/nfoJRGVBagGOgELP3ARTfuUZxX7sEHYqF5AZpecSAb21GM/sP29lOm
WJg0oEcw7big9kgrvguI4OPupOGqQB0Dp6ZqdMYybFDOPVrLa7cYmQRRdvQXN4U/GjSsW58OrDQA
rGYPZBsXs051IVwhN2R/IozE9mxr07kQWxQFUbHy3sdqsle8efe+aTyzNtKNB5D6ku23X8P8wLdz
a3WTvySC/mM7jwmM8jSzTGppmEpqk6Oogil0QpfwjRrbo3ew26LJsV2pV4eECDlIhU18gd9JtxhO
5untjEvC5PEClIDLzewB7Xu5z0tstXTFcl+yjPCQdWCE+EhQbXgzYmkn8WXP7GSLv30Ka4oD8IRQ
IZsN7v7QBKHzs55gOWr6b6nVew7KLU0db2Ms3m3uGE8ecvaY+Hl71qm7E+pOhYz/Wd+p6XtrV6ba
wWjh47opXO8ejDdhn640vuv6bbm53XgOr0fMRtFGa3kjSEOVQQMRmOkiDATemyOVecJZ5x5i5s/i
7hOsnWhtfi5QfMNNpw48M1trG/CqJIbr3+UFe0epDq0Kn929hz9dy+lycnALvIHWlq6D3jYG/mWw
7xFHrhWG4ACoJiNqJj2p0Xi4hXHZdp1OZPjL9VqN7yz6ITNa3nepv3pZsMNZGP/rYtSpgLIGQTvD
v144ru+LQ8SjzM75dmPFaQtH3Y4ToqKgXb1x48+4Q0EpHCeHeewxUmycK+fGEwUNJg9RTxOpbHKD
qG0x1CNNzrWBphGG1+zpz3qBylXdO61/sG1TCb0J7YtLrkKjn0MaYHCsVD54ReMpGA3y/9LecTho
9AzLKaKyBKbo491DDKKBlAyrls5DU6g/H1SC2MTTCgxy2n8mC18wyFrlmC7JKnTwrPs7qEeJjFAw
ZBwkAZsfiaYhfXx3Z2CiuEIQlVI0zwCyRFTvSGJCmhVSZm20OsS8R07mH9ivfah7O9emhrNGX3rM
EZq6LMz7pRi99ouS6nlyaDEVMR9HLnQWV+se6LttyYirltdZwoN2fOedkyfYFGHJu0QlflIpLo6P
2SdMBgLKEpOeq45eRE0wcR29ewQWsBQMhGh6bqvJikGf0XtqzR2xSz6/fiq7GEK2KxauBZPdLkr1
iZeUNTX0kzgkxiBo7etJ//lmzKpIGt1y9D6GMlJhVY+uIMCtEODgcD5ClBgImFuyCf5yxEGbi/ZW
sQv9tut0GbzQbU6jWg/K5JtpE40AAgvfL4mbq5VWkKCqbUQvb8pA+LJcxU3JbQi6nMN9AMbjlQkb
zyPsfbO4Z0lFGf5nsc4CA509XqrMUth6S/jCpOuZb7PbsQtBzmo3UREeBQUkW2bQ95DeY4m8WmE8
LHPqfsF9dPYX0L4+JimOmAXT/PQ8f2S5lcTOeJLLj8ives9RydVd0a8sHst/ItyAs0SWXAp7HXTY
asSu9aksUJ6u7LdXH+6ohqkXyx5nGVuL71laMTsgae4wGeVBjgJvQI79XstZ3adVqZlSXoXghaB1
doWcy29MIb4HidQiYDrQ3P8HClrFsa8xB6rnnZ299LKB4S43ynDiB3K/8Pfwewgw14izgAObnQh0
+N43uo3XD63YMqEVMbPmbXuWy8zDP0CxndRUFKOUWZJRdyN2+vlzSz6aX3cDsaj8CuSWVdzhR532
XHmXEU8bmKi8cYv3x6VKxWhJbZtrDp1gamv5TqiY3PgMaetDnj+Ow35hFnbXpQySFuc/L0g3UBMV
7PVRV1cgVw3tuS6Ja8250hLUl/X6R2WzxQGr2LhhFelbdNuvN/iPp5a5wB0haCa6/rs3LZJZoonI
b454X/v5C1ok+yzvhhWNzeKvnIrwWYsWMpTwtpoFuStd3OrgL9FGgvu+4vpXEmHmvob4wM9HG8D9
Z8IUnkuwt/rsNnXPlUlDS6hyoVtRD+PRXE089wihKwVcp0PzNtZPhe99VbZ2V4Ag4iGXYxT0JaVi
zqr1k9AjdjCgXOCvkYlnGl3tf8GiHGVxtcjZ6y9e3x+8TPHJer0+v4Xn2iFRpbVhZawVRlrLbNN3
vE9yq/COGrg3Ba3/TYfkWk84U/vLP3YgWdCEzKZhtvgdlMZdi/LsCBDi1JZhT9vmJlD0ORIBUh91
QzHpjR6MRxD5V+vOAv7IHYinZyDrwpwjq/4c9FgmF/d6817hultiz+tPp4nqArsa5mIJ69JKQEQp
GaLnNPlDQqQaEw7BV8KTl3efunxbmjKM6UdPxPhcAnA2kz8dGcnjtc0/XkQbxw9UFR8/gvWyCLPS
9RfWP1okJLZhZ8g6U0B2GXBk12riMXaQ94PsxHKAIJofw/xzq2QuOb/4kt8UPO5vapZLk2eAfuqZ
8zHd0c4YDf5Zff7jJDPTp90GYiX/bTj3nwpYGr1h3LHxvu+yGkXNJ+rPn6ircdw9Z/ApVbtd25FQ
faBJD2Uc7115XCtE3Z+GSSJSLgtSRy7QwklaG+Qu/FLxkj7mATKOkYYCiF2dK9orceJdqfGU/0p0
q7C2guP5ZeDs1+qcFzGpKQ4i9qcIFZnKB3UMDB+3ymvm1g9eD5xcmKyViB2dzFo2kdely+cq+PjN
svqZHsxY2v6HZHBMQBOMpxRD2zvNsqkoOm4pE2uVpQ7nAlHQ+6wuj/ueK+9PV7IWnyCW7d7Os3vm
RmCKTIIQOHK4byGIsxs+erDW5az1qNjg03QVLudnKPEQvvk7lMZti9VvHSl9UPoZQ40vs/ZD2b0W
oZahgmbt6allFY+Da2fQbnMcdKXl1scyHGqRGdzcXVunwoBqkAkBfPzoBZp/6X5QadfOT53An8jw
krMtWv+zqyqZPzP0EH4pPP3s5fcE+AwbxxMhgP8FxXQPK2qVCJehQQZBwSdT9kEPe1HAl7pFTuNy
X910e3slaCBaZooAo2bptnZkSOk2g4a7vaG2lm6xI/YQaSFXqikwql80PKDE9AO0vUlj/79rbk1e
9CTfDD9ud4oojZ19XhXFLRF53xoFjIcCr24OG7gMjaUp/xi+ylixQDWRCMz1Tj3WPL3slg4xC87w
WBtR5T8pN0lEV2OnVZtR9qgobwxSahUa858B6Q0r8MnroLzuiygXExFiOkyaPO/e9f6iJUjbniBV
/G3e0t+w/6m5+2zB32m8ZFXyntym1Yi6r7GlSLbITxN6lXssfCPWEneSDhetd68O+xwtKGx+QzRx
X0z9cD5jOQYzglk65JYkVvV9AvE3ZqzjpdlDa/BmaRA7C0Ngqf7xlykwQcxNUsKYceUMI98eXZoB
9GQB7lBZFKxW1XV83UO40JHTmLoTdG9kchYCztHN+HsqxLzLpgCZr3C/mBcAuhegqcbr9cUUmVL7
DkmX/m1UDB2sfbeAhaqfFCK7IF3GMiL3clxNnrsyd/VHfzsSOhBm2WwkfsWkR6u07T3sGJmpoRgs
zUbMecj3w6bXgxcPVWB7F4EshEDBfFSmXerN2KnZdJfgUtYElS9dhk64ZWKymyRKSbt3LXXWvNOz
p8WrHuleCG4Vuxq+Qx6OYFlYOwgh6DWshWzOOtJ4iyEze0LqAyTDPjWX9fnOFCActLoFrB9R5nDp
i6ZDfp0+1070cc6tmcmpYlz/S0BV1CTB0E3DdB5Nz4M0ccV1d6q9hWNzoEAdDrfD50T7kKe2kV0P
Dk3BFR8yRJFgnVIquK+MGuxv+qM/do98Ex8gp9WsGqhlYIKGfPr9XPZzo4lZ+LcIaLSab+XIXDc0
72wivfKvP3nb4vWkDaGESSeAS3HHg9a93bRTAjcV618mgFwJ2g0zSaisJvWr2uhGOgeN0qv3rVD0
hY80vcKNoSGU8Z91YzFCmkC08xP17L/E2jY8X77OC/RxqJlZfSWWU6Ko2gzSUBXcpJ/jUngIxliz
Om/7KXzKFX5KM+ZZVKJxdBWjN0qD5eSrWkQ0A95I2RS0wETKpjxD4kgBYj0s89t75rsX1kYhI36D
Fr/2Wq1/Ef3gaHupIbBZyZdkfEtEn6A2lYx3TyPMXptQi/u+BLLAdnWrCuNo/92fRGkaj4Kdj3Pe
YCXUU+ZUL0dMWBPG6wRMTlacgJ+kzB8dWguYvNx8jftSHRzi/f/7w3aqtyeBJFZCXxb4YyS3TPiB
NeTHe22VgYQRKZU/sIv75yDCJTzS79ax5v48Z1IR7ZF7qW6+NkBPrOmrcEqQAvefxsALomcUcvad
VeCe+YdtLtgBUe9PbfMRCowWG5RGyMNpg4scfbzoR3KluuZf6CWmDiwfMYLu23VPvTOBtRJVbXPk
Z1t1MkGsliiAVUgV2ml4yx1dgebJxbhegciWuALGse1Osn58DvazFCGvF+svxb7B6E2L0szMCpYg
4dlKBgvwfWGkPR55fyCGKhqSPAtIKV5aCumL1fGUMARomBkdOEdT7GOuhwVEEPWDbiHz5sQckxld
imxmnsM9VVoXTON1ZR0B1zYZIIRgROj2rnvBsTCr/xsGJZc6rJFOoW+HgLTcoxMOspVvs5JPgfFc
oJs9Z1t+dNUu6+r51tfrNhOFgZV0qaSsk0Qz18ycXQGVWHomOBQg3pLuT5hr+uW5zG1eN7yHKdZu
SnxoCSzv338cqbfBQb14TU/CL5ZrsiO/05H3FGp2HKpN8HxebPILTZ+LAWLMaP/Yen5YHLu1Zi7N
u90PNqCbYJB97pUingvi2FPtb5XtkdMWhojSG8mi7/g2RgY8lwseAUN/TEyG02KGo0zSsFZFfeY2
v67YuJLaASk/OFj9QrcwEgsO7P1yacuFoIITnjC1IMJTsi+ksYl1XiuXn/4WZa2lzlj1Nn3xvs+q
5Kw75lifeIgI+X8JPhHi1VD1+wOys00E9ahKtLhb8iqOtaaXfhPuCRDXvq/FDoMRW9dqDmW3Cbis
iHDeSZ9N+dzGNRHIbx0ERjRZyDtU5VYIocyjuny3TtSu4aqPKLJKDQrsPlQ3acPMVfGrdY+eAqMv
2NWr25QDftcf7hLg3C+DmxgQY9wCDxQUspn45dxL15NSWSrRW1B+6PlFge9mthKpcbgWmZ39pHh8
kjL+XKJQHl+aHdW786crAUuaFFn2f1OmpgQjrpqBoBmVun6ZPyeI1ASHgPvd+MqTUOVcg7zHyjE9
DwO42iOmwvIOgWlMHESGkmYTKX4JZ8MlsK9wVebYvVTt+1JNipPxIWswuQcytY56I6uLZF9sVc+Z
XGPi00zVHoemjB9FvQtYQ8Rld6fuN+veBucADXnue+kQjPWTh3kPyRCICXWx5tG9sxR85GvTc/60
5fPMEGw/hLltvWgv6+8j8S/fWQ2n+xbIOYaResQPQMFzTp5HdDMCFt9U8/4XRvVw0v5JOf+MDm6n
Ot6j5Q9gyZoo08sIorBXREn/sILh1+UeScDQ/GKdfVbGnvLfQ7Wa2cwtXxyMDfGn/cpinkj/b3GH
QZXczkfP7I9OoOEkzj2XQKe+8Rert6pfzJ0UwvHAFo41PhOwdjt6lXCqsd9eJdCH0i1Feek1Zm7z
lACHnSpnbnTPZKnwDGmb5oQunNXQg7+2zXUeASklEn/HF3i+nSsFplWmGWuGJ9rJnfeacB7YWKnb
ASgnCXI5zm5EU5p/vnYlk4m06vuH3Ajcko7l8sWB7Wc82l63BZkuKimBB6PSMTV8Jpurr0gdgGCN
L2yGkeA5oxnEFwyDi5d7SxRyryJjMN2a54beVhcGAtksCi4UpjiuQITXQzlrRAPMJ4ixS9n+m3XC
9SEjo+jjOQQfC/Vd9o1BQef/5a/Xf503EyaSrtW6Fb0G307pHCNxegXPe1TgBJv6GUajHKo4Y6FO
xkmdpwkc16UBN71ogCEc8rPkqf4WG0Rf2ME4OMohu5026BCT4N8xFbaQid8JTu7axnZVmNgLyUW/
cVa6cG0SCKh/l1s1QuasEa+iCskb2v1odgFXLAipqCjCO1uBnk6t3P9ypfz/IzIg+FX//n1TKshh
JblGZEdySba+7kZH6ETlB87Mu6OcZia9dRgPx4D1wZKuo2W+InSmfM4xwJ3wcP58zeezB7hYyRW3
OR2fTC7a4P2eC/Fts1jpa7YVcLjpRvCQbhGIi2Zpc9zE4wfXVKAgL5E3Bkru4xYUDntKhlR4rSNe
2rWAY/Z7ofS/n7oWnob4PXYhknw9SwrSb2NjhTkHpFH7ReCJGugxlfSEuFS03OMBhW9Ye7GMt46y
dIjM/+ldt3W86m/Xxsm6E6IDAu1zDkuE1UX+f8qFAvu1iHFk5KNVPLDsxjD1dmKrIlhyOwEuYaUU
qGKe6LmNo9KlofdBhEgBcfiu/2Ta/o/1Nsa4cCGjXHMB7GKZcm33ue+NHE61PYUEPCTKgTKtEyjF
o42vNUDdVHRYGII7iPWV+17VZllpt8Bh4zN6iZmLlSwH61xjH36F4ay4Ws25dGWTpGQSZpdye8vN
P+cVQekNylTwsuymzKBANeYlkqhXXdKcckYnzLIDZUME+KezmRVloZdjPaeQQseK87aINqmdSb/f
ZwBfqbWmqYoydiB1B6Sao7bwxq0luIekdugz+JqTcna9zE81VYPnnTDUPulkdOgJx5ipwDbFFvXz
teIqozqje48RdMGrZNX5Nt199kJ5MMm0A/goAhwyyCH5z1Xn5s7aPGRHfdYIC3L6qL+Gr+jEatfr
e9dxTCQEVRg2d7LZv+V2jKsGZApmZBPDRZ+kvw0WbtvBIaR1uIJjeAKFlGJPhLYl8qiQfgUex4Lo
r+N8buRBuyAI8mGYo7fEDqilllRgr6v5FbZNyozrcfLvNN7jyerL2CaHpXAULkieoo/K70AmVoEl
TbOPSJL/JqbAxTkcNfr3OnRD840y19zvrYGIQMV9gxKLSYh6Mch4AovNusLffug3YSE234hAD8Fq
5l962kLC66b3rhWFBZ7FJdPbo0DrA6c81KCkjb9Rjn7BbmRV71gncbmgSVhvFChnjC04ng6r4FV7
t1tu6V0PZB7ePlMaa5OaYHz1Z1GK11mTZJW8wMEwF/qkfDPCsHh0eBdFKSCbeMb/YYftMFZXy0Me
TW8Itlo6VwqAfko7/ps9H9UP4iUC5MHPxzKqwfina84vkT7W38XONDIDFP2KkvkpzSNGZALtoWt6
USEnxL9dBojQLpnAvafSdgnGsJyCsh5clPgz2w+Rb07ohQ9YaVbKbuNoK/9WJLGFk3zh0M35ROrN
wUkb5KVZfjgwUsZ6v/vfKaexh2q3kf7zcv7QK4jOfY1IyKjjUPYR2rdhqvok/ilJ2yTKaIdNoh0z
SltXIyDHpjbip1rVYOzF8qc7+Rp7n+rZrTGs64HIr7+vY8wosq3yuwzeMXKfOGxQf2Iq0QzrMGuh
ZSE0KqdQaZVWsbLn1a3/2iZbW7a/awAwvecw/ABZ5xg3NU8Vc0L5reZZO2THI/6HKi2dQ4OP0GIF
nQitpAP2GHnudclEpDR8az+dIWCShIuG2X+tmaqq/GJtZjnb5+nXQCEew3lx2NdCNM7fAdwv7wjJ
E+o5NkNL94A6xZVme8FHeJAfyrp2EmRl78kNToAZ1Cc0hlsBGyqNEiRlGfywxef6BSqk3BUS0dkc
9ADPTYg7xwh2d7gp39DZR9JWJiaf4JXJaZJeZcJveEzPN/pH/PRmUHZMC0zDVMprNocAZ9sbG3ok
Hakb5hqeXI5v7lArJDeh89zoPBf3VsDoKowtNfMYsHGGz3DDFvmRiht13REhawYYgFCFbPMXwyPj
xMT+vbdJMAGfnJkwiAc4UL+eYvm+b7tUIJlMSK1QHBy2HGHVMtr7UwygiANG0mVMWECYxNEnTqSR
hJg6In07SqWb7nCm0nmI69b9mp4WUWsV3YMksJS8DAzLyL5ub1EXu6zltfrk0NBSYD3mMFMcLtIJ
obfQp+Eix0wff2SBo4292D18/2jbPnV7ngINOiHwZ+8B02YR/RS1z6qtKQSHF5w61j39S1T19HZk
YBa1fUALoQAa55QXnYiYTJpA6UsbnbpRxGc1ALJjxCImbkR/1D5755zCCpSakqNh16ldkogGL7iN
Lu8ui+twuCcFmlSxaQTaI+b9MlFkLFy8Ns8MDJAUdFskmpkNC3ECCGq5n7zDmeMKKIm4dlLGQ+2M
zvHYnzvbHo8teTgsfqMWc8/pbh2TegpBwKQHJfbyag0GuMx12oXkJxptBE1xC6cr2ElkX97F64J7
dczEXjyWhUp069EkCXMAuoDbQeYk9CnZYujMulZc09pDLaJc9jgd43ZYx4Nhs/Mr/aOZAOc8rT1x
vei5OxPMrkGVhMmTSuZR3Mtiwer7LDKXLhBryoA1e3BgRxv3hyR7CUGu0NMDc6vsYJNUKcMNpcfV
z2CUwm7+uwBHFdKo8wMoQUaIXo80A8l07Ocx7tsjA41FihD3YTBgYcXJpROmc8U1DMEy5hxZpW6R
horWyrDK+1OytKjBUZpTFZ5RlEiZWidqf78QM41QPT/iYZaxwfY9uSS0AlQbbNoh69yzN4hTIgjE
+cz5Rj7aL4oEuSwtbncy8hU+12gOL8rqIaps2EbNihJiOblok4FFMWm66ou30ZxAZCy5aQeYiauA
FkCRJlItWcygEX4iDslUi06mTY8zLeEfe7Re8L+/HNi2b/ix0vBdZje7PfK6EEk3VlEvcIYg3jcV
r9NtTLHgP/JNRzGGrXcCDFLfaSXwP2RiZHCeMle+vM9ZU0AeyVyp/z6ryY0CfaPNhRsrIsz9HcBG
OgGxWePdRd8QramPGCp5WBoNeITj5SSZWZPL0lAVd/pVzfWLwEQuaHnLJrneF2pXWy1bsH49hped
JsSE5J4MHcL1LdpTlcHquuStbxGMhA7uZwi88qhq9zzNr44zcPhJGpCtua3TuB2mu8q0VOy4xbxw
V+tG2PPJbMCSNvO4deaulVSOyT+wSTaCuvisJaRDeVVFPB+aPvo1sXez9uGxNiSbv1gv0mwTg+oi
+JAtooGd+8V5Hpcv0AJjjYLffzvnks3GmLJRU4JZZNmkqJRc1mxOH+JCQFM0y/QPDfipxnrwFz8I
zyd0goyj8alHuh5ykOLfBzEWq90lNoADjWpiDxinS6/W7ekdGrjUHOMouxCu5BxN3WGIUG1pNsYM
G44blgqizWUT2S9UzDmlf8Tib0sqs7xei/9LQClWOucRv74Dhm/biaJgVLytqUmvaeR5TgVOA2wl
oWW61qU4AeEJ+7Gc/XAlfozUwR2IdtcA5h+nHs4/VcLjJ9a3fXQhr7F4HzGWYjHnrDLyVpgJ4L0k
AYRjpUoyf/1iAPZYoNlzZCswuMOijz0Vca30T66BcCiDapBuJpoF7t1n0cJtbXjs7xWECw60Wodd
qAnj2EXj0ELmjXsSxCHLEHgN1c9UxCU5XdIEhneRc9dPQokS/WFHP0Wz4/EKkdtcJ12dOGgdU29w
SfG3M0i0duD3RQC0a0aYbwG4pLZALZgsCyov2kziHm6GlUyKIR4Vn6tZVTHVvgYTlfoGNUNbOGBu
0pqEIo7n3mMkJWz7IKR07/N1ECzTmu4haEnaIJ7DB8RDXzrpWbJqhZIGW5pga2DeFyAtZKsnxnK8
vADfVeiptGPOkKcKHlZ8uhUC+DxiSuPsOGpED9wcj4BsEpYsjK37rwtP3oKvz5Ll71JLVyDcxNhY
XoAE8L+UPZxRd0PJPtvdAn5TSw2vzD3JHOuuFVPW/XyjIIZxO5dpp5gJ06IfAVphhMfohBPTmO8+
2Y0aL1L7OqbgOySS2DMjnC2T3GPaYtwL4m3W7TuSmiAwyMbnzC3IInqCpMTi9hVE1t2+Qbxi1cyR
e0MJxpV3/5m6bxHr9o5uVVI0JNcI02nIHf8Ev87b5PeEg2h9K4fQTuCGNvgUt+vr0FpfPcRboBzr
IpOoyCB/nCPLxTGF0f2My38OqEopgcwoBRQq93VsS2xgOTuQkv+qvUxxzl8FfNXIMCAYqFt1pKwi
ThDufu4/9xlSR5Jn9zLOzyWDEc1AwqfvLJuEx3Zg9hLIPMAVIEr9r2owwwGGAnnW3FHunO8L7FKy
SiMdP3B8ZhqNgHdEeGK4KzxW/DGb64Q/wVDOMYEjFrcX+CXj2uC9nHOKdfXZl6cMEWTUyMjBQ+cw
wUqnA/YjMIEys5trnRj6T6OX90k2wBTbyVimtzmdkO53wuKhNwKvnD4mXkJCLa3iNP8+8d0JULJN
7SWrDYqOIXZFio49OAWzdhV7sS4aQl/Ag4BjiZmhThphirgxwWXJCuNTEhSeUSNWeSX10eilFk4K
UqA6x530RY3RSoSf3U8oUPh68/EGV8yfqWrQKwo9F1uEYJtChvZSBGE46UlVXUOtlk2Gwdf6KojG
sq9X1CeavLPGsQ27s86AwGyrSKIi1CSdN1jHq3NNcBBE5eJyqn39WKWsunCwN7UjdqzpSJiV6Zdc
lsMeREYeWOVya/U7NsMRc/VoEHh6G40KPVwaot76NanvXDKN+nKxBGiO0mcuF3MtxnVv+TXsYJ1V
45MBRCOu0mhYFkRCzeNFInytKb5Tlka4Cwlic89W0NpP898PumnhOeoVi06IVGk9WnzCCGm534px
bQ2kJL/qgsLSo/31w0xyMsEMh02A6mrP++fpNnRwQFc4Zxzrf9GnFmB03fm2nVVBrSFPUHPuNDG6
qdPEePiMU7gSXe5U/ka+1H0Bl2K7VOboKF6LT8ZFbRRMx2hdTH32P/s0XQwhpdT+6M/kbrB9RNQt
jhXrooF0CsHC3wfzXYvfTgt3MP5qA9Uu4Kbxxi8gfEwGCuMiYH4HZ8eC8nLb7cv/aZ1fI58LVSyF
INs6ct5wApMKfxm7rDdND77nWjtfdHjZoiqLFxpRtI2UleQ88DIb2cA9crdWjelM/SyPmeD4aqr+
McdoggiAvbrhFpNSRlbRuNZAbVbplWIRRa1lz8b2A+hDVle3obhIiYkwGDyVjOi1AMB717E+wZNx
lL6/V7CnnkNfS3MBUkpZyOmD3AFA1jmfMslWR8NH2k/pmhgkfPTiqVC13KegI92oAeuZP+WTvyoi
F9hZgqk7k/ftubVvP1EHQi61w5y33U4avVIs3y6j2nrh8cWnUJ/vGm9MnU3jl7YetHYi32/xCzdN
x6R2aFLF8BHWqC51gYk8WW/j+ruWkEuQc5xw04gVXn7gR5LnaMFxlqJwr/i5IPqKIp9Ce/mLS+N+
eq9pPtHpT2iXLJfA5Lg4W96ZAyy5UqyZQqVUBFD31Piw2Pf1gYhvs/kf4wF3hc8kByblc+nkGAkM
2D1pcJ3bFsxx1mlHqvlxfxXioPBR8VoDx4J0iq4bNvDtIWd96fK1buQvschFmmFwgw33vUcls3Be
sV8YyqiDLT8pEY5QUoAVQjOAi4aH8lcmeME90lAbAdK7U4wymwDLG52lQo/hChqcAOGJZl3/OUOa
xQat19q9dI/SmdC0iuDpiRb8eT+nrndB1AGn6zlT4SI14F5Msh4RuZE6iTN8cCUL7vGy6txWYx2K
uu3dtVP5Gh1Dg2/TOJ/Qzdck2TtUJChMRRAbnSoDRNLcBWu2w0m41ILvZa76cWplJqORJc8PoAYA
QIrDbPNFeYd5yxo5fctbrhTvuux3YloWgUNWtERdC4YbhlWgLglEofhcIm7JOp09NQxSjr3qmGT5
R6SbQb/xPCZNuDHXSLpTzWmUVWlG4t/sa6mFZdJNu6hJNXIUMaOgxF/B7B5mQTfiqutUlErVf+R6
3ZU9lKcS7hPrPOfLDyjhfctxkGe5RvbZHMz4ZmRJKLqp1k7I4lLIBhG5yFRLY6JWcJ3gdb992gnu
FFR2sasopzLOLWJJkAGB5RVcYlzbBPF5lK/cjVKlbCWP/NR3KdYRiuqtapzwqrwgpr9Yo6D9ngoN
EH6qo59iMF9kfcEp+tEYYYhQMctBhE2jutCXcptvEdPHkJHZhnUm74Hpn2ERJUggFVInNilok5P0
LPUJ3Y2ILewvEThd8u9nz0pma49S1wlsIhuO+HgwZuvcqf0g8BmsZVZlgma+U5kQ7LPw9TU7YfZx
aE6d/twZggXePsNL5DZVencJDO4hxvSv3w5YsYKvl2+Jj/xTMfW92QqfJgDjwZrRNEZ5iLq7hsAs
RS2Yr6itxnASqKUn1tLXxOnDLD5oOaWxcxr44bvayL3gbjfAPkRUjPR1BGZck1o0gbX0HKK9kYJy
lx/6gDitFqOqREYD5FiW7ryu+Clt6Dg018EL9+D4nVCbMXfWZVIv0yXTXxG2V/lqSO4zcBQnnobx
a4Vijisq96oizNVNCGMN4YciI3eTiS5WLs2asEKaXA+8FqMpqMxNRvA7CbHS6Hp2+Q7C2/cBfIMH
fFU8MacLF2A4kpMNsNgXW4wyrNeqRazpv1mAzb/2yn+eSqEULFPjHfcgKcKf1+fcziiCuJiLFEPg
fkfIeesQM1f3i7dKCkUa7CdeDBkp/OB0nzYZlC/+J0yEyrdSG2AP8ofZcNOQq1BDBR2JnjsTOrZR
jlgxDllXil45Mh5xiu5uFYcHRa02VVyI5Etg1wLOFpxImHSJrJU9gkCNhuiCAvrKKzfFoYU/+aaU
fLDeRzEx6Y/OKbq7T6YrweqrALGs2IWWIfsKp8KqLJqZuvMwIHrc9iw1djUHIKPXP09oN1WwENrH
RsE54fpMPW/ICCOtEk7j3zBsN93GBcMjdRQxBf5KdlTZc5/WWIl0f+jaVOC4opd4VNFeqCNwBNo8
33qNkBF65pUB139k8XkLVP0CwT8u7cHd5LOXuW2bn+1v8vn3P5UREzNuA8cd3t22ZCdPXKqNKbDn
5tMzgNu4iNUg4ybcVgKBfme/gRLz2qyT7PFMA4CCkI4t7egqPTTli7tQ6wcwivM6PaO8qqpYWRbS
z42x5S6eTSPYtpz8ms07v0sNk3nhmd6xQAd4i+4f16hR3NgHkD7JNOeQnF1CrsPlHGQvMIQcWwEV
k4bq6g9GhD6tsvBCkXCuFCwj2z/wlOeUTPXu+406oGz7t1qmwkadpDiT9kgMqmrlW4CDtGyi/ZPE
DCPK9hmNN0myQQZ30vwNFnItw7wO9ZLYo4n6BpzumIRuCjYr5w9zbdyFlXCuJ4eaR44aJKuebe70
Ov1oTbozwpJOsuMzO3mN0ZJMPDhlnvehm6Cwk56+5H7nTWO2roYtSuXUuMf7kcgAWI6lf54vTrY2
us0Xdg9iVJbS65+cjoIfdFxNpiS0EScNxivm9Pjxs5UFA1CbciKP4PLngTKtchb21+TRwuBY8VPZ
CRSRlSMMpEaIALKC1F+zCIncFO0EXiJIHc10Vetq9rqFJ1xUyNwty6FycUS9yOFdgzCpmwQhvuXw
i71UAu3D8W2cx+zQeoDU7u91MZQj5MofdIZYSEcCIbqTLuCp6ah1A+fBElbwmfGaxVnYkiZhz5cQ
hRr/XwYy74KItdikK59Jy0XL+UviXXZfqk1X7yrsR8Lra/VKjgkBMzwpymo4OtAwCQKgyDM+6NR3
HR8ZWg463Oh925siadh2SDK0bT1jZVGwmcJ3roQMQ/WvwkfPlcZ0MWSOEZTTpuMLjCXD80hKr4fj
GwDUKy+rPTC5hg6nT1kotY0N81RKh5d4dzViplgcMgGoZATJh36mHJbiJiypnx9HvKlPZhb5CQRa
RLa8GTZRu0taDjHMM1f3SFPH9YZAki16fMP5uOdZb1yaalQUI56FzuBzBx/CA0s2GaWqYbHo/AP9
EbDtjlsZ7DIdkse8IHdCE23g0AShsr30qQkyNuK5kL1s0IaCXgEYTlnz3ymj1ken12/lurB+CuGr
LoEb84L69SH8vmsHCabzy6bno1dsi50WKjqwbAPuXcCfJMDwzbmDqirCMQbR9xpXq6tHOmaulc7m
W+CfrcUySR/rz7b1MgT5UtUxA98a8wFgZ9CKdMnTrhvactMhmVFsrBfeHAEb0NFBzvr68ltPyxnb
lmkSm5sHiUtaKOa+qOliPHYpKDcD9NdiRHyldIsgAkvazspkaHfE6AiWlhgaWNfrumoh2CfPRQDG
cyXwQ/JcbnM7taR9DGfF2QeJlVug4KHO8SeeGK1y3MVy6bA+t+WdMhIpGrYGRqCOClb3A5dYd0jL
CYkDMaD5+LcZ9Eo5CikoJIorRMSRi5bbx6IJqdytGD07/gBcz/rX3FRgIAmOv6EGlroxBVXyyk6A
Z7SCkLa3vP54OSLUebb64otqeXgLBOkYh5LuX1woWSvvQ7DiyfqhZD17UnvXlhs2RVqEg/6+Vivn
EdOMdFXXX1NokEgg4tMSiBbzsNSUwe0xN+5FmDlhtHEsVWdl9EXqNvmxPbkY9I+DBkvTDtLGfmhH
qACxKfwFHoPY7DWdjLCNJSCemG4tB7vauqhUuNZ1nsdtB1cCbVEREQ5t91PqkNu0plRAc7ebtxj/
pxGZgTJQeMRQ0fe00xjwasRbIRt+YzHhZN03PacuWa4NPg4MSGePvdJLXLdpieuzViVseQtxKCnT
twahEJLIcnwJMa32BEycLcNq7IRWHMAKAmgSVfccgo0HSPeq0MmuSBjyN9Qy+7IxpG6/21faP+ei
OIVHS43pA9IxHHgONHV9v6cxmMOcLMEmKxHR0BXTQmXqNwapRayfzSzx+SLd+t+fTYdw83Y2zRnX
0tSb31zsRav2B5UKnSHG6iLk9n5ujJXOvBUAHSPdYnSCl9VrOrRRxXD4KdfOPeRKbMriQOMFVVG3
8R8eVolffR6XfUcVrXtAz+FU4BiyyK9WNXQg4/XXW1CkqcVaObnUymDa8ygupxXLrgQw9efN2PAS
9xhyxRBsCfGtuHXwbNUWSCRGIN8pIO/CLjcolVXK/aEsaAQ+tcvpsmuC+CFFKaTVLVSQox1+HdDk
yzo+274jXoM9+Lsw7QNpF2APc6IPnPYTCqcqSRoeBDZkhNX0TrSXskFXPJl4mxSg1X7kB5N1hUDx
qUjcoA0NzZMGNBzntqc/L/JNCga+GoqTTFEkOWIp4g9UqbNU89teT1cClwcOTznmQgOIChotxKJC
wJEsn+3x/pqL7E7+CTKNdL4lmrY45UsThsCXVKHFxTNsk9azvqcn7veFpYv9BEPE37uTQtUv54I4
SoyggCKXzBix5r4ZpHU4vl7M3BChgDfMpn+XqBYi65NLBY6y5qPcfr2sHXUGxWPDOaEfViS+b2xX
0Ql5PlMDbriYhUWPX86loiOPidnzS6UcpkW+JhQp8hjrsKOs+13tNnD+iA/d8jT1FB1RENXVRlSn
2xJP7MxXM1LoZZc/GBkuqUzjk1RU6BddjPsgnrJ3hYQWO6p5U5enTLvJ78zVbVHD/gsRSR2sUUKw
MuCJzBCcEw0EmbQ97hqGm0C5LeaW3eCed+aWPvb+rcB3necC9lC5ztf2xILLLJ9p2TCeptV5tmiL
sEBnG1CPxZyxUih9SNnn5nJWdXYBPoaehoM5Cx9rkNJlaRFZPjHIKlLWeKOhe6Y7cv6ZdirRknkI
jT/7rXLoIRZkGHb7hb8GvXmZGgKc5FtUvDXvGY+hstEhG6BAA4CCe/waUNACBtFGuDLD4Lo2lzev
xQqMgnCekreNC30W9Emzp0WFtwuOBosB/x+9VmDCLtJK1gPXt4uMBQfSjWWRZmG8quIC+wSN48XT
EA4SuFYKf++r/T7cT6UNbWMcX05S0YJ64qF1fgOs9Q2wMsF4DOtbAUQKC7NedcFwstvPGV+8FiTP
aJFinWPyrd3PuSsgJQbUVLJWJT9BTXAF2RbXA1wTaw1lcpJUvV/927pT/6uYou3hvhqbWw1XK2r6
owODqgUXym88aDTjS9Stpcvgm0iE4IrFCcIbe37ju2WUR6wizbyStrhiIunXD9xMcrwhYxiYQm16
2vMUyiWwXj1ROm9+lq5i9AsyidWt2KGbhWVo1abAv58re0RZQjv0dxXOBfuVpfdUyQxCY9YGIwHP
5DJcgIyCt9K9P5sq769mXsZQNWUCfwU93I8EoVCFf0uo3wLursXBHBo1nSxu0zrJ5X7MjuQF3hTZ
rAf1EQKdQa0E/Xp27Rq81Dlv67yeH39z6+CZy+mWBZmj0od7kGwL8eSxniM36aivStk6+tQc4zFB
TrRT/T6G5safeNW8r/mhv0vgcZNwBXNEEVVo6fYCRfY273MngnhHooZIU/vRnaTSRoODbSIdZmJD
NZkHoe9CNUWDTiIqwedaesuxoP9z6cZSBu7yjDATUAR75Nu3MYFBQFfdMSotdDCTSET0cpp4YPNk
SYKMRd7aIcs7o60x/XvrzSNi1z2yh8eKTXzFvWcOLlhvLgD6UooHbhwqLicfKkUAMVFCZE91l+Bi
CLYfJgTnOYuIcyu7muwoSNKn/TZIzofi5cHzQt5gsj9vAgZZcJGnXtrkpvAxGmZZuJKw8wJbE6VY
ijTvUulVzODPGWmadiat38Jo286EAOkBXreSpFcLjBILaBan3naROyeNFDGe4PCc26kC3Abr0E/r
BBKftd9mF86zs5sYkpqVKbD/why05cvrp8Tp+8/LnTwjsI+JtHmrY6MmnBuigJWFsspBbHBeF68p
n3u3RiqkF17fLGDif5YxF7kovvJ0xlYTk3KhTqh0W0Xp+PT7Wv/u6U4yO+JVC2Bnz1rZFmjnAaVT
HvQN0wNkzSfHlUNBkBYR5bl2m1V77FdjO0lc3ojtEi9OyqLXHfYuuw3PixIZTOHBSWIGjjBUFdPv
Vqi/NK8H0e91Gi0UFG9XbYHOn6kR8SbfoZL8oDCIYXOa1gTSZi5g2YhG8ZOcwshIzHQTEtpu4evZ
//QGWBgnkGZzNHUC+wK8jXFR8p8Ga48OzzBte11axuzIt+5ywS6YtxjcW6rzRfCoxoiZgB4txv/t
7wWgdwBiA1gLT+7O+GxIM8ABXNfSycXWijbAbM3HHUny2foeNuqsbIyCOhGylz4QtS4AjVtQzKxO
O3XfKQCIoMcVhBOssy6dedbpYcKm6qVosNkSYebjAEDmEkzUvMk986TF41E7yO+I8CRYZCS+KUPj
J1UTf3vl608kaG/05x3xQny1VE4WZnYjxQ6U/OsBDxCgJYQr6GhLFAXUDj+/fY72VEvx6Dfc6HnV
varuWJjlJAI5x7Ue8KVl5nw5usQIqdgG+ISwDnVxMXsMG4ekX6uy5GE0pErC0XX4nA6nriKEOj+f
0qG+y6j85yX9O275c1YYE8UCc5RAsOQFqvIAL3KBDEm2dbN8Vjg7jAFYrG16/KxQ0lNHr1uawfwo
p6VQJnPr/5/vaheADszahaxcnBjCYEFljAf7+jSu9a+z9pTXAqOWROXs9cDsb2PAInpLlImrsE0P
Fb7QvJeNNcXjz+rC347m0g3744OxOL2pmP68V4vIi2IOj4mpqjAPfYMKi5HsNX9UWkJQLaoDVmaD
JumgjUgqcrwTx/Ud8i5UFoIFVciyAD1IkHi7rcCyEC+nBTt7IX7Q0xpURXBWq9gV6R17vvOWqche
GJd6HvK/Xk+Zkn4kf0xQnN9Pb7dIVuTtgEDlBNUYgq60n4TFzKwK5vXHLl5S6J5cTQrNZf/Ynfnq
EeSSlCd9VzusMR8sGhgOf22Hp1lig3YSS2vCLYWPeeu3uwA3puz8TMBsVdhP/zlUdrlFWCe3NADX
i1ga6a7SToB8mmUeJ/B/vgwahafNw0a4gMDoyWwJmXV3pQ4nGVkGXO0+dtGkxeYY15ga8l0c1XIm
PVr/JkzvqMYshuzTQuvtbS3sSLhWTiECGLj1jpXi/2S85CwlCMyKXAFGsXUqVVs4nXKB0pR4chcs
pnL8Z9/5KHVo7DY8oczkfvgLvaqPsrGlH5qfe3Qq1TM76m/0zEklmdKRI046RLUz9vl9Ln0vHZNU
k+eF/B9VGKUcZeNcQhhnzKuEO8JmLpntEodL7y+2Klc7lbQ1pyHEKxBBdSMEliRfRlXbezMSrTBk
6K2CzHxPCfPunI0wBWR3Sul+/udpPU6Q+buNvqqVCnKlRWf39pza113IE7yDo1yBEF4TP8mKNqVw
LSrQ0oIpwZrbpwNrqzwKjDzTW/1Oj46uxeCMabJJUnCPhs0P8Z/XZ9gO2QI1g5C/54YXPXlZ1Xlz
RXBb/ZYf2q0BaFv5FA8vrqIVtF9kqS2Mhov8TtP/GWIKAMkXhGo0zghYitJqGsTmlt2LiQ4fZrIn
jIepOcds/GqnXmc57MhlPwwTRufXIrPErLMd5acHcsTvfl+HmcDM57vz5+DsRFZ5yu522+fX1TUN
l/YObeDOTqOT+hWE3fK6p7pEMNnWm4/8LNUmi2vMp6J5ySU/JoLrjzhpEy6u3ehiUBjlF21i3KJb
eDwMY5XovXpl7Ogxs3Rn4TSVj9kLTNTn49ZoOtTCGLYLsFsODHvN43exqRMmVjpMUgAbNL3odg8q
h/TyHAP4KmjxQitmJ9LcgqcpGj/8TobUOa5y6xTyIt+I6S8XmoDPL1+nt/WBTanywnNEcuLKAdMr
wG7yFJAO8yb5SLnQjyZINSGOa9tRxAlOKwGUG8OWGEwC3pmeIR4Q6pl6WjIagY4ao9Jxezm0aa3b
yLPACNp7yjCJD5Xv6Jxlfy92FbvLJYPh08XmlRnUVZ8h2zsv27x6inIPP/DmrY2vLseO6tZKf8lq
xy0HB1u4KPgNeTfwzC1lS7Wq0EZaR8zGPvGc0TbfAOI0KJguPNvVJkYfAK92F0Fa3dZyMMX0DQzs
paRE997NgLvLqjerb1DGehxTz6TXFguk8x3mOHPf3OZxWM3fyS7sAMpgUvm2iOLuAMYJoL2dzlbC
3xJ4ZM/SvYajlP6qfJ4AuunE5GysPQYt3tBNIrfnKh/QfWxPvSyakElIrJLWUzQZVQoJPNjlWtKI
dPBZ7lZFGs1tBQdp/ky8qDCgDmz+7RSFFXMVQhBG5WWeKvC7tmCK64UF5tqsbuHAdGs/FELWVt0d
+gDf6BRW0NTFXekhKdk+d2bjPSIU6/oHCp1mcK9vcqDQ9ji7VnQy2J5wakLQgaHfwl5umfwzgh31
0Ik/hU87FsO0eIJ/mq5qcc2sAuKqynGKOMymQ0aSH1+pj0WhK54M3ddu5vvUZS/fs9V+M0NAH3ue
kU0FoywwGl/GH0wXhWTmrLOg1g8w98xITn52XY0Rvs6er7qrhiOhVxwmj8pqhjHmK4MwkvK2S5cG
QmAnKWolLYX3n3de/1sIEJn29JrjtGysLA6dDm91faCYqWirGrpHlnzcSy+foqDxMqK4Dw/crR6+
ZC7lHvbZPy/zgsV5nc2rdx74YT5Ec1klt+k3GTJmmddmjQkPAnMSw+BYwcd+fjDgV15SkU7Saw0F
/p/r+z7xP+ymUsDMnfsu3V9ETeRwhZwMS6yPIUpXZpZO/uf/tzK040zgw7ew7WPnAhnBTDeQIWIt
VsKNfbeMekXDw410GDLqWmp23KIJdHo73BFojA92tQsFo3VE1gkZaeEhduXNeXJrVaIV/CeahHiq
V4PQ8GEicVRRb6xmMkHMfqlYgqmwW4Kxg1fI5RYjF4XCXk1FCqgaV0v2k/7HFXcozo4mhrXO35iI
lEkA2/TJMnzfquxhXBSbwxIxqfj4q0QVm9VvW6Y/2u0haHYpV9rEcTCnqWX12cSCM3R4ACt+YnrO
iPm6JLT2B8gBC0fne4Ij90WvIfxRXa13uv+LOEeCEDcq9sTbASxLQ37NyJGmisvPyddyX25tvfkP
loDOoOtuiEMK+TQ/hyTZiOgagOF+t7JRiO0wjhu4GRjI/9R8VCAqWoF/gdAUuJyUUz3Ay7tpFd/Y
H3qhhcHf/Yc2acdDyv0KODqFYYR9EvI5ncAppAhA8/0QMwiwEM14pW1yovN0EVWFhbWxl64ZAptx
LBje/UbHqJXtT3VlSuG3fPYjPAOHBkT06yO+ou/Mi5KtnnyzKs4i0tEsQwsJ4+inFIcEDQN7tsnm
c1zVG1cgmJKIg9LubxMVD3DcDsihhniQBViR0/cTr8A21sStC56Gb/3ua88RbxJHrp8ZENQU728g
EtimnblXbr/RjdysMQSeZIqesUY859aMpQnifximrp8dvVw6rR5xW+GprRrV/MIazLkKE4iQo69a
/Ek7i4AgMN4OXR3uDagRjm/iqdKPLukQBJlQcQHXA7rsXwOsqgqlPpGhq+RfmbnWv3ZW7Pv13xUY
PNl9D7j5T4ntvrn10m9VS31GIlRip2y1dtVJRf8BfNoAAj1poYISgxgPsbZd6NFPaGCU/wfPeJc/
v7v3th0SWb3BBg/OuyXkAnDTBNr0mZwxerLRFyqMwLBDOV0HzydVewunbZWj9rU5EavhMIlVAp2x
lX9meRsOzVF0u71hQagRAGDoBexJeidTjmBH8j9TTefiXLNvoRy45vTJo3mvhM49O/jSUf3GEu8/
bwGBtMmQKhzXf9F18L7O06d3v7C5djS9hBefWkqb+CiajAj6guRAWOwC8Ty6TSpA5KrEKvl2kYkx
Xmr5J/JadbOt9+kqphKhnZ9tp6Rcty23cKigwrb4ySYnI8gj0MAbiN5bX58T/DYymkvRJL70y31M
I5spvOWMXxLIfNRJGCE+N38eKf+XgT9Bj1ZUge7CYLpu3yI9XVHKjO0GgcZzexbQ7D8/Fk3TVzvX
8ESRZelkP/aTtGYkV+8PKbxCWkE6D+3Yz+YoaqKVcdV8/DZzHZSn3Oe/rH8TGfze77z+3xIaAgrD
7NZjv1ymXWcHJ0BfQ8RtoNfJndalZRvrhGyyz3m7mOCuxskokoOAILtJsQczwxUinnWuJnVBzM0T
mXWrP5ihIgnOXKKWXoEzhDecsJzR9X22ZbfjDdg6j4LFlpVUw4hOX5TDrZeZ2gCjgn31aform2HI
w43mCaSeHq/Tth6AC7ojORIPZG9ZfvV47vyWPBFEvLEOa/25TZOk2n07/KbamttQKLbQIqvSg9kv
lTTWUIAUBF4SZ2+9p2PHuoefmMPZ4eIOoW+7LSyA7G8GOI4nXnq9bCUrI9745kC+iGylZ6iJursx
gMdRDh8gUmALLXPgWPFiu9f2vWdFO9rbW8MmSD8biGVa/uulpdchyT3Kp4OJlo6Z9r3fwNBTJ6Ts
VUhpZlSZng1hFNjS+QutXnd0JFERB2V8g8+Czdl8X6x6OL2ZokF1B9w9VH65LelAufDXIUYJ3u5m
OiWEojVLxsCd6RnLczurIi5jFpJcGZ1sLd8Mw3VZZEWc3eM/OlAivcvmV5WIpFZVvos0ZDtFX8bp
WDK3bzxXliK6LVV8DsqgD8zsC8ExyyWxYoRNXbbTC+KfKdakzpqE/6sKEpHQXVjxTubiKp7OgIP3
/87yNPIriE/NDUT30SPOmt6S+XeL9zKVLMOli3TKO1EkieCR/hiv3qEdPfbJ2SlXFwcgJp5kykUF
ylDOGsiL6PfHTfVtL2q+tNK+kzshH8AjoY1fVd+vsFNHdw+mLKcgYWem9XBFbh2ZaJaGmoqoLUy4
akWewP2oq0IMt21ig/JLmfzVU116eQlRBmYRBXBjwc4Egcf69+X+2lBTSIVdpVCCPG5jTnSafFrp
uwDznoi9DKgemvEnffCpZBhusRz1INfQCswnZH0K2k3trRW6qrbofm2vgLRxDNo7yZt4e4PquTzB
bydSP5TnKyiDS9UUV46k2llt2g+2hWIT3B30rSaWF0ul755jYpr1Iw3A05Uu4dakJAomJMTFlRuv
g6YI0MB8+VEn/l8ySorQa+8rbfQ/PhmDoBW50tgsWMth4MoBSsNbhTPXsDinhTDKHdhaMUygcRmN
s5DRu3F9/ERUvVJ+aRxrTQqKrpzGjY9E872IPt2Gt2YfhAmv1JG9oFtemvK47g19zbSGy+djJzY+
3/1g7qvVt+6Y6WxngUOB21fvFv7Xt+24GL/H+Zay7OiUcycaFcQjN4ObcLvCGjBZrOpxwBmCNUcs
jdLrWmVUFYgiQmJZ/EbK8BxW9GgwiO0US1gbgbXiVwBYj6Jjhc3C/bX8TzWkl60gu05WAZIQ0RM2
dW/QRc6pTlb/QCQRuG/T/A9qNz91ZzqcI0/dCEs2yd0OFyrRUdxugQmFcedTlACI4B3BZMUuJbX5
8d69whedEYvFQpkopkCzlkDvOM3I/ThUZqF+OYcaGYD+JNNtmpwM4+NbjFblcrtTrrbtljdE3+Wd
gj/FP+GsM09rCnS+/4PGRJXELvo4vb6NJi3pMWpOPZ5SPofkEV0UZHqJW5VYmYSKHi/O6amOkYtX
iLZpzEd2o/PcG8la/UmN8tdDCD3JHloowrY73FceVB+M/z4Di2hxyK6uxVFyY8jzEBoRdMS9i23j
htwrWRGdW1Rulh2vclUc4Vlwt8SOcOK2a3wbkBakxerk2a2bSOvY29slsf8EoNktkT/WCRVIGx75
kQqOgZQ3PbpVsP52aiqXIojlAujUlEf4+TAz22F7OyCYfLT6nKzZlgPJRlt6WhniHKngO+JqZDEV
pUPgySikNkBxVjw+LvE7XmGpxKKVyHAYi/co3Jr/mAbajG3/nmiKG36Vacyu+5gfCrVJFSJtzTfZ
jxgxlDgU+t0FYzXMry8dHaCiqFYJ4xGzC+GKLvlpH1orAIpKpmA3rJQ9SlTnkFuursofI/oPphYe
SC7bkev+Dmx5+Rn7s0xZvk9olHlOxCDKQzjOmypi4CrBP/jgf/YUZok4bGvgx3oJ+lxX4TMn5c5Q
o20ouGk/SVobcgkHKpSrEoYQUucGOyCnB51a1hMaTKUSDvFXRy9F/iB/Z8K5BhlzH356Dyturor2
oTbdynCcBpp5x1Th+9qIVUUKRvwuFLvjRA5MaDbn1+LdcBLlRpf87Ca4itT3AU5DFvUGoMbUC9NF
MqrP1FJK2tz0MGP7RN5BF/LMpWZOqJ5TwkdU+3lpkp4mdDhvMlqM83GbjvWKcbPRjPeqxtEMn2rj
86IMS6ru4tTxmuvYB4yoM8xVDVv12snB4hkpB1PH8C3BvW+hxGm3ZODunjQQ/vF6ckWa3gYDczmi
jJotNV0Vf+TnyUFrGhh2AZrsITyVm4tUqiNos4pnD6D2dPJaE6jRRB/8+VKbS94EQkHBstFJTwC7
+b9iIU2HE/JqVqA7cRLPfaWlkRur1cK5UJrtVcbtoqlJtDHmtCeHubcAYIVLTBr3/XxD4C3flt+b
DcRskx6SI7pKSYorSi38anR9IPPcGqwsHVpV7BKG8aRIOe5E32ofhIj28ikh9V2LBbv55r91x9aR
/dZjzllQ71hoOtHdd6rHdxvSsaJgk7DbOeRhtrAZ8JtxgPt+B9L1fu1s6bhAMenRyF/MJO28PK+m
aV2VhqcoiURtlDeGFSVktB3nAa4YYHHdqN1D7gdLE93+I+PQl2K1RIO1KAKAeRJACOlSH3RsgwbW
wCjeULtA9G9Fb0RHApy4JRbzKmPa7Unq1uQpuHQiX2XujSKhFsIb5AuYTrV+a7FamWW2wom9QsrJ
/24EsHxHX0Urv0qNpMBvYslYWT9UaQN5M7o1oAOkG64V2II7maJkU2TxPiUCUwkXkflo+s2kEc21
vI4pTJ+D6Bg5+Mh/spdx8oiiAehSB0C1xSCxHroQ1yBRKHAU+1bwcue3450hzNQ/E9XSqT4xsjut
1DXH4K99sZg9MYd19o03hAi8qETG1BXSlaQzBmiT2cfvdHDhZRwe+dQgXs414XPdoLFe7HuE7smB
zWFhBc6uFCOJxtp1DhdI6WLxhEvoa/557MDBRwpSaFEQfOt0BLJ4w4fdibUhSgkc3LBGsDkF2mC/
bAbTD/cmX3lI7b+R8xzy3Filo0YvIlheD4Hu49ho67EY/Ol2c7lBYUcxaSfZkZMF9oBR4o7qWF0E
K+/LCzPQaq7UhZwzVIdurKllrM1dcYm4x+mXkkqexhn/T+g8JR9HFGLilSRBgTa0wBlD7cryKY+N
E+r3tXyctv+q1mvbmrNF0pdv/QX/qFTaPjijfXvyQaxbWPq23n6vnAN7+tJjVvslyfz0TbHGIU7n
U6/XxlOoQUQ51U7nOpfMPxh6GA9ix5f7ULM9CqrYh5nPKEYw4dLpHV/o2eUMPuykqqYSlZl2aG7V
Ha/UDqj3gvbrCAm/PrB+7Whx0t30f9h01yMayKeO/QR4Zu89HRmlt3S4Zt47PQvr8KnawU3S9C3E
I8ciTxOrAwKu7JkPc2tSlJGQ1LpN5gMN2DmI78Y26bwAMg9tVqnE5YRKjwcyS+rNBwF5bkcOAbcY
DOzKnauRRRQ8iG3tM9sKL9/e6LZHjJ3OdBhNR3Qh7J4wxm+5Y5ZpMsfyDsmklzoSj19A1spJBiqR
o3dMW1i4N123a9x/Srlagxl+Jx5pZ0ohndckV0pJKzzipp4vq0ZvrA12qlp+bYtKs8za5mxhokLk
O8LN1NlZMguzvoFOsBrgyILOXUhKihzTqF8lgL17HCR8iKKYztMxSS4hPQpPWBKh3fisx7WGZs7Z
QtKsnJ8o8wnxweSah6gqQrxEKaPXca7eo9zEhCjbs2qHW86wMgc44xVy4j63hoR9/nPlqdqhsmu0
ZhNvVIiorKvBJw9wCAGegGyDiG8Mo5PPedWiZCYyV34TmjUcQTb2WzCAlaA046YW+J+GtKeJlPdB
EfFEdomXmeuV7tPyfKkuPo29eeh6Vk2OHkE5yHQVcBO1+il8vQBQHpArZiGrd25vXxpH0rpSMo1J
1L4fUylOoQqy1BTgq3ioI2glqK043Bk8ASydd9H+HATcbsl1YyGBfnLY/HtLi/xPoSnHlB638otj
HtTTKsDzqhoeDheMcz1yYzzLJ9v/g95Fp06br1PgGfwFZKjH7u2jDa+0fkwI6B2GSCtBV9yBq0Dq
a9q/skPVRQTsU3bCHQ/ByPmAppNcFGGMQl/LpiTwvkY/QTQjHH8bnR7dMQQah+pJ7GwXGP0UPuSu
3xF4utmI8V4a0Gijb4o3CDdnrBMWSw3tkiwAICdZh+mNbmgC37PiFQ0DmRTZSiMqGdeOlbhRimSE
0JyFN2tCvnIvddOOy6vYwxfLO10UX6uKzzkDXYHetPXrncDRRXVJmM4eJ+MMqjKIKchrTE+7ZL04
UkjGO9R3SbOLzHBp+yh51fVJ12w1wmUK/uqNL7994V9oGV0mve/gvmLRt/UskHY1eOnps5ADBShU
6s6Bx0Jm88ZvlTCRjvmhBh8VdG1KdQlsvmDDYtzn4ZTmMw8ea+3asIJx7lbzQCr3aPfaThvQsORg
zziUPFZXRb+6GSlGilF6iVM5EwAoFnApfOypYKiOtkjWqk/gJpWP2hlax2SELimS0YzzPoUKtLLu
wdzHVN8BXs/A4lbYo4yh15Ny1FQhImkxeoEH/bAyd/CpizO7ex9vjd4970LrIfTZsCY1RYWRbSWn
vSBWGCY0qwRMXQSHLm1XTBM5hfpsWk7hewW8BjCSJXZJqxcFlWhJIqVie94xDUIZly+q+/AT6Hc4
LpAVqFDSMGBCNA2DIqDVUBCng2fVfKQKzhfYaagFC1K5W9rSqoe4GcZWng7hLcLUIaHSgx0qULgB
SrFHk0l3rK77PWzQXuY5UkaeJkVDAgZO+hvScWFAbyApDD/jD60Wg/kyA8ljemWGcG1evxVEayYB
vAkWgFOsp7rBmogok07s/m+qFHY0fzQJgFdAjAovYmo083cUvZlKWj+ZoooF+Gr1VkVvtDBuHy/u
iaEXHoBIHnhnjQzQexZUiiJJ153e2PbYSvB+v7bkX8QXF9HQDblboCZP9HGYuLys1dBdMlLbPtvU
IUeMBArkOnDV0kELqc6c9hXWP5O7IKHipX2MizdNHm6mgows1tAMUQDoLNXfdBJWmRbG5mbQcyFH
Q09f0Ki1CAJmFqnQ7SI3HC6ysaG9Nm5O3ZdxQDaj16hyXslpKq98RGWv1oCWVluie1NckG6kS1WO
K0/KP0ADpNRJzivvLQASJFfpFvnUUWBelOExdPoRLbhgyUsh6XCSbPwokhZzBgLH8+QvZzfSEvLE
aNFln+rilo4AD0jkmsJvzSWBcYN8EiuNyDpeRT7VGoknAxp683b5yP8s0TfLRbe83gbGRrARqdZe
dJltxk4dItU2eZtvy8quCGTBfNZe4byixmqFYxf2xrL/cl4ZGu15hvOXCpYDmusMoAVqbJ31TaoD
ShM1kNqLPK354rTSlu6bXNqnibvVbE0GLITTQY/ZitgNKb9oVfr4UKqQdPZX7qW7jzo6vj3jD4YD
ogU3logYn9QHQjT0UyUP/vNBVBTC43YGSmiU1yoxMpDuto4PbgjOXE/Aqti3vm7RiwZC9ADFBxq3
csr2DeJRJfUmQ5GefevfcbjqGJeoyws8yuQb8POyh/xEkOnQNoGHJVbc4WPhlYDtHxqhUMKW76ql
Fs70KIo9lPf9pvjEPWwfB64uDDDMW9Fe1WOFPBwX9K+TOYeyy7jvJZKWbL3+iK5Aa7Sy33NfNbGt
W1QMdgUljor+g6BZIEo0xyo89+UPe9FsSI65w7BtucBBu0iBORUfsJxCqHMrQ/yH19Lm9YK4M9vY
HrqtBi858YDNZcMmr935MQ7bhZoRv3kO5ktXFvE2Ndr8CuiqZX5fbKuwYi4GW0Aa6mGyxe5zvXO5
M85D6KCqwXlV39sBJ9wLI8c8cUzAqSlcTJf+AepAlaphhJ2fFPruUOFzBy6wCqrpwWMuQVUK8+dD
YGXvUkUS+diLWGXUTxe3zNbJar351qqGcEIkW91/wy0dtbgMTvNeYFjgZ6oHx6XtahpdUaDP/+kq
J7E1/CLyqeHtMym1d8tuZ0i5oNi4LvZWtfoWkMFFWG0ZyJZIz+cZxIjFHz23g7OK83XSK5jp0VCu
MJRAQiBznzJ1hzFy4JEsgLtpIgbFVqiIrOb2dCBer9ewaJFg9vQ0H48QTIBqtfC45qcl+BJcN40D
xJeH5sxtPNkq0GjnhUnUenYfCkjY1N4O2R9+0+sVZPNAqSaFABeJRTL14u6x5JquNgUwO3SzjdTk
koDsxxfBpfwOejNgiv6lTsKRqUxWyqBzZGuWYiPnvQ3tDsqETIjJWU7P31wZ5ySDaOkhZf0hRVn9
XZv6GQqZagL+dqqcVe7IcooApN0MZFk7+5RUXIHjGlWCg+idmiIoLpqWUXLmrq3B+IQyJW7j49x+
qAvuaeAzTwgO4bK+CI9srb7FGYXaNXAAu2bDTsSN+ZqmIJ6OKGFsilNHcGkLzoY8HKvT9mSM0bBL
mbkVajZg8dUxhHbghZaENbRl0vJMQHq0CV7HO57g1v0QAMRu9FTuaw7OJb6saueqXS5NPUa38RIe
lGfXM8cSZjFNQPF5EvpxEX4SOPwm/9ohMG67NdT3Ai2tB0zWp+yKav+eySbzlm3+9eMjq7aCMPGw
mlto7ykNMP6kBNz8eeFT1SoEeGCWAqdrDwZtFxVg5+DFqxM7RaqIvwwIczWXdl7VDKNTc4/Tgj3L
PCan07105ckoOnD445Ef3gV+q8bHfIMXIKfVuxfGvnF3myU+2XjS8AtZ9SBDrTiuVZlj89lGKCxi
KMzEO46PF4uRlQeIOU3BE5fiGz9hycSCQnfseasgYEu7mgpcYa4zb4/K2KzjIT5bvNF3We4SjK3+
XhWfQy4Szel3paVLVK5fEhl4JD4Oqu6M871PWvWF2E6TJZdq2pIphI2ZzeY+v6iYt508C2VJlEoS
tu6VhoetVJbvXSdPHucNf1Q8fi0mfVFjhN9Rv61N3wEhYKHWl2bFzjV1ygSwYeQfXUIT+henwCPo
NP5oOkxosW+EKXT3n2Qyxm9E0RWa7p9nmZpZfgXLaJUMGrudiKq+qB56E686feX+2EVdC+OX/dfA
G5bw1VM2q10lzSaB39x1gFnL7CNy8P2OUKL0Ae91ik8ysyzQc4O6vTem+RhLV99YeIGUXx/YG1mc
0UudchiYdTrIv+NuUogQVBoZ4WzxxG7tWmZ/IMOpviSGPWCAfkr5KCEeKvqDzAdDjr2PoX5aRKmS
wb2U+TKCnqd2KpLwO0euPbvVmUJRv5J1udZUNYv42VSuvmoAD4yLvBcoLrq/uHDgwCQnaqYvJk++
0bhXGcG+TdtLf80Rp66Hzh39dLfQpBpQkQ0g4/z3G7hYGeHZSHJ6Z2clLlxoKfITK8GQGM+CConA
tdqXeWVGsHBLWjIPN/x9ar3HdPE6dh3HMeUR/QaewVxjaZHMshetAUmbNrPBLL8DvtkNmihR9zow
YJh4MFjoult+0IpO/VwIazcay8lVBwImZpAnKn4yRVXATAniua5l4H6Nnd/BRPpgPussuW4spvM/
xkprCWNXXoU3wC3MZxE/BFHKFX/WJX3gTj9svVQdp/yeKRtoKH1JJCKql7NpgIlNvmfHNX3QTO5c
0TlROqKbF2pcjA3y8SIhVt7jqYZ0gezstKGRQyox4kqUFJZBhSCWfXfNrhUZhlUmqWLLoz5eqI+i
+rxJBp+4s4n0BP+r4OeR0/W9CvvGQ75/3yABSV0v/p0M3QhMZXK7d+PjwiXKG6de0zFZ145nQQuX
VmuMaXu+TXyc+NEORAuYtoK4RsCf6JrqLj+gTE83J7NUgmu4oucY08qqZCIrkuxYUwWA9JJfS4pH
i6z8GYM3QSlBaKS6IZp6IjtOTgIZpbYK+lhmsA7YVXDiYXHFPrTt3ZTfAbRFPS3wEooC1RcL9iQ9
tFZEFIgaWRzgiDgONiDOm9ppMwKETTWYpKiqs9um+pddUy3wXahDL9wTifnAA7d2rgertRIrNpBv
1epPXXnkEr8VTsLrlgEhtbrrwvqWEHMC1SwMu2aN5WMqUFJk98L/8JwPBx2TMi8RYFq8dADLNnLO
7gaKmSlsofJysjOgHKmk1fNnKU4veMPKVZ+Bi8nJlZU164yAmMa9dcTQdJT8+DheIsX2C0kYzgEJ
BRj2jiNcWDYAnV53eO830P19Y5rNxWsQRHjp4L7ltmEVZDzxYZ75lODuvwi1XO3y8QBuBmVp5EKt
Or7J95fP20G+I9Mq5ViCmJlwgWZ5U3ev3/7reu0RvNCQWehr3ioNZlqvB+2JHD48yqSWSojm97kd
MztHsFAmrY9s8MqJiGzXKL3Be+kKCrYX9TKoFTN8jr0lcB7qjFjhm8FX06OJ/YW6oQi0g04o0s3A
B1/BQjBXuqK6rj7fcbTlDZ8G8Reg6T8R03UtT/K1hzpjEYIiTlfLfoYQDkJAewBrmaPdzKi51LP4
8aSSC6jg1PD+As57+XLSgp1YG/A8/HjJcWYLsDC1EWkAjHhiEi8XHtOcy2QZlWUMniR2Deaqkuv4
Fcx3G9PuxiuodWJnE6lfmYesFN0B34T5JbzpqrJUkpOqlgQ0h9vg6yr6DXSeo/toUJ5TJw2tgpQb
7S2PY6lnCIOLdBhqzIWdR2Haf1bTW8IbA9mOrUUb/4qTtSMuS95bjvQ5CTbjcErtV18pAQs8+qot
KdomN0EgPBaoMGdw8P5XnsWUKhYfCjrQ1zMUzSVi5EVVGE4P66a193aeO7wKCk7wGW3o7XELprkF
8JxrpzCHqGY/1es+W+SBzA60b+otnwPVKt+6Su5pgV5bkPRqji8vIdl3hDjwybEe4u6QA/6rEB4L
9MWIwAJc6di+3n8V0po12JebmzKJFEkM0Ska3jn+VP9lteG60l28pb2VvXkph+ASd6uI2v1lRM7c
WaJ2GNO2ZV54WJ5Z3B5vE0nYR53jUtOP6162dRSTwcKIkrundphuID502MCT0kyroykFDrhTJsm/
SLWxwjDTBIsAdZbflTXH0rkU0IfT2Yia8RDiooxwwJ3Um+uXbNS+jps/Fd7NQaVzYtfUfXuq+9L9
+kthco3jvxC6JftvQVBJehZZ9dpaLERDUAdw1MDVDM9K4Q1WZluh5/7Lw1O6h18Qagi9xPR+TVZ8
9mddLfiCdag0hMzidGEsT2lEp1w8lE0gZS67GGv5HCiEnN6b43JrmbKqq+/0H2JGiGD60dZmWmNS
jzaaXstrNHv9iaGpuUiHkPp7WlpWCcIyaMGVd+x5XF799xE4TQ7b7SsU1cfmyOKmi8vmwa4zTRHx
tYSEIGBfNXEzZXKNHCBrtZDCFxGwgcsrw/Z24ggLpsr5l/IPCnA3QuywHWznOGPqtcmZLgdTBccI
tYGcRi3H57foJ2HMYM82AIz79yi9vzdyf0nfWvBJXEDVhW5ueXBy/34UKqeeAzVI1yzRZqHP0XFD
7qiot2zlg827kl0LVElMSeLq6eNRFlQ0wh6T6p+kE72EFhw/rgiixP+b/5B3bErbl8qxfLW322Ac
DjfuAVOfFcG/u4dnvC0qZ8Le7vjWPV52gL3DbmO8dBWr3o1hTfP74qaXhHgwCXRV8YaRTvnkssSK
JjVXCaCNwCNNMQFq1qmF8EhhLP/UKq46HdmhBkKuH0HM7geqAw2dKdcVykZMuo5tGDkj8HvlOHhQ
L6bLL5Rc2gWxJV0L9ipklxVI6NXOQ5on48SCw85VQfmm/S1UDC4WHmEd6v4sjVOYCQeBvMHhJnq3
oSb5QyJHRE/l22p8kBnx/C/RHCaWh6d6AXMUGsMmGfeB3AcsYy5DVCLi4FOqULjQJQ0FKOcLsFOO
zhRjhJtzv20cdcjFx3dA06niW2/nojzUF44s5I0D1hj2l+sqSE3zngGnfrkd2zpZ1lqN2+EAhDwr
+m0wsCn+hgoS2MRYwuykq0YsAbVCeOnTFDeky7kYz7axt/SBi9Ic4tXPt3u8T8PhrNy2EyfFJc34
0Lp7/z5m1c5Hh0pJzWPsM8SdUWz9Sz24ucTZAGz+B96eg30QJWbJQLrLCctAmF0pV8ua0Mix3WNH
RNAkP6xgQfh3z68Ca+2Z6Q6XVmXQqiBDn40m1fHC6FeoG7OdMmmNFGIiaWwxTnOZ+wxsR1mYvESJ
YajjRPc6IDTgGKlB3h72suoShjRQN96v7Z6TMZT58dBpU6sbwZxV5jyrp6WOyk7ovVjr/XMoHoin
3UkxzyWTQeGt4aQ0DhQqnkYrIYtTH82lpKT0cpBVPbOTs2pSStuFThbactAfNAPLdwSDVHwHSGxC
Q/HkfsYkLBJkPVvmYYakiUB8CY3pntQDIDPjFyUm9Z+rMUI8k+3HovW1caOQ4FVnPriH63drOkZL
ndAJioB40BgMkXlE8/zXfDbQeicIfwNyXJpdzdgAjzZnHjeSMK6xeMiclZhFEnSIR3S0kUVHsgLl
y6jMjPgc5JcuryU8TDWppfNtjY/b11HW/vgq+8HfjjwZBBmf8NQYJY2i7o2C7fu6FODpxASE+HVH
UX3dqvd9KWT9//dRkt7VdVnPI6FeJnTRZ19sEjlAbIpKrsvLvulvwGc8j+RdIjV34Gzr7RGrcLC7
eFKqVaBMdDcjgHDmENsYA3LH99R28Z3AQ/h6LFR6xMecHsThxJ+19Rov/41C8iNMLe7k+1eqwPNL
0+Sf6kkqFQU0UV5/fTylaFg6BXUO3Ty7plhUOEoblUeJMBLFn2GaymQkLzrvtMn3rS4Mwcfg1HM4
cEMFyIBTuLNCbf4ii7sZHPcGlFrbHBqI4jRDAQ77aF4jR5bfZbaj9Uk0uHVGdsqFDM7Z/zbxjZ+U
ktE1fuqM2dbc0uVXvuHR7GqJFdnflJzmBSHi1wtxwNw7HkAzYjqi+SPHK0Q5oEA8yIByP7OLCReD
8zoweNs5xjFrlxs8klVj43+ywOPB0UCU9+lQOiAWZNHxMmcOIokdg/p7ZT80u+LVw0av2+WTDP8G
DasPhEVhvVCBC3AaHnqLddMtjQ6i1lFprtsH4sRv79yaIwDCn9wHMqWTraFHEhNyCMWj3c2GumNy
/UNbXtd5y65VhNydSxOKjNTYgaxfmN/5FpXrIgmzWPqQgioku6YSICJXgy+xmdBG8nZrZ3WuXhJ+
EWxVb9kbzomPLLMGrZFjnMuI1tIM2ctWAAO4l61YGGxnnFHStAcFXK0+6DvyHWP95m/Q+ioUbDDv
NPu+ROWftM+S3pcphvQ5NTdCOLQriiacpjxdmTtsEmmbYfqWHjWL9n24KoVlmsRjdd+jylNXT4LH
V7G0Pz8hb0Z184f/5DctVOuohaK0Z5QdIBofCvupmuMw8ysdA3PYOtcqLk1B3SHDwYcYRycgN5Jp
BoAM/lsHbn/35V0RUVV0MQ8El0nlGQysNYnlSE++CsArDNV7qhIX3xSuGt5CWUYE0lT0D3kj4JiS
D+kiiYUx7l6kyPCzOXpPZxOOuYBdM0N/kYYAshjUtbrwkYRNs7t98ZO24cRe3EbSyGdy9fes3NzS
EMjWs0wCS1Hv+rYqgfXxy2D/OO+ZxKF6B+jbQZMGDD/iGvL9H6kifqVeX7JlVkO5bjKpqH/SlwMK
kannco/gecc2vOxG68yBci4Jl0RS01sQtXcHExSEF9jVTI8cDYeFfau/E8ZgBBTrwjs/Bpd1o3Y4
1XiNjgD0gVD8K0H2ZqMTfLy00qh+uYj+d10O1JS0xmiA0Quy+/g5nxRtazf5QdQEFUywfr0v6I7I
ypEy0Bvnk+XaXnxR0+yZsqi/XDg18Iy9lk/WwmvSM/SE/tuAlfhNNU85/AmpSkue1rnvLSuL0WEJ
MUey6L/VDGbaP0vVbDmZS8Eh3LF0V/MHaJrwFiTBS8sFaWO8lSKMSFToj7YsIqJdh8znPqKvdNsr
dxvUIXfE6yAdEmb0Pw+jFqJEbpkSLlZTivSrynDZeZKCh9FbO9SIZgDcbVe6OSNhCzq0JzPnfJwx
1mOOC+BmXX0QAy4MStQnCUXbZ62Zr7BnlKFus26v2zsWScSPZU06FCuiKKVEJNsuji2iJBc2GFxo
vrB/kw7K8ib5tXubjlRyrjqPMw4suo9M5BTW0HSi21AFYJ40N5meK3pfgXy9VbeINamyHW3mZgOP
IT8z/3NS+u27mg0YGUdVO1E4WzN0hyun4zDCMp/yKA5/QwxMGqYg0UAPkxEvfTQ5GpK97dhN4UYW
UJ6kE0+vz++GPZ/nCIhtMrxGRtBP1+9P6F6DPuEuLPBL7Pm0EOP+vIXbyba67RMHULwFICSB6ZGh
VDWyHHNgG1UYsNMN3tIU3DhAGvsTnCa21MCpzlv7aaMQtu563j0ql1XsgUFfqG5xvYjZ3zLJ79pk
rKkmpJTzepUUwijrlrg8NL4TYk1KUhlwKlWqP0MVlsJllnQ42CypEL8jkdz8LZU5ETBRCB1yAnsJ
g3GK8U1nB3ETxSBJzYdm9hEIfCMfujv6yxnI+T1UqI5EVHmNtAgwGh6Pw2LDLiOfCLd2YbIvBdo1
M5x7bNUBL7PW7Vj85ETHxup8x0GUWFOO9CrZ65RizensUW/MKJQjWK4HYCxpHw0YX3h+aMKl0k35
LfQkVR1k8iqM2xD4lhf7q16aRItRMZYZ78Tna+AAwSEx9zK3Cdpp4OGCChIZ//x3Ep4yddKb/VSo
P8Sn4827OtLJ4xjIzXPdhAO+KBcVR8K9B+pUEaEcmFKMhRcIheYGXqxltwOO/gPWvHUE6ZXrAcjS
qncZ2qco9fp4U0YyVo+xvRMM184Si8EBzzMj8zwNqcX0YRgEX3FACX1tfZGNajAnMyVQ9K2JK+Xy
AR0HHVWRrzuYHhjni0JU+DrSbyAwmGLI3w+d4K+7VuEuTLfEEat6gyHtVb4fwuGvj8ju60ubH0a8
2ER7DQzTtLgeWmleIDqG+9a7ER6+xRJy0xuMVImLotkAkB0tNbpPBeScpT2nlu/R7SjBjXB+wIcf
Lpr1ksCetry3T15j1Le0+5csh0Ogq8He5pGvE5q3C35zP+9PMVVfLVUjKhvhn7NKhNMyMnPpebT5
wPNKbYgiH4nTLOH8Rp12nB01QnWiHSxarTqsT66sHDBN1yThEgWjK0fDWXnc6WgibRgtR4VFN/++
zdXT5mSYx+qAQvukecvwmHOj+z67XWApFWUat5Vs6UZmLeGSMjmnhuUT04vqryn13jjrisdxF4/e
bUVkj3oT4HV1/+lgA738stw14dwWjNnhhzfsGIwuceunbW26DeFspUjWVdMS7GKCJ70gCGXq92KP
IaqPrT3Hsk7hlrUJjpWaEZfNzfjbRMRrI9ZkdEuxV/Bgl1aPKpN6w5mNeBzr7TIGCiQV0HPJ8HQG
Hk1a0n7+1oNST2qemm8w1rNk65xbb0XZm+GTht9Ietbqw3RE9xz7h0DuqEtzZMRlgD6xXqzWGFMg
hurCCUfiW+rbBtYXDtvNx6M56gruNd6HnEqZzY47kfzmzDYVSFItOYrXrjsjM8MDpsmJ9/LF2DS0
72BaPY3eT8h6MH8nACB5PPsUFM3bODnrhtU7hrBjGAN7sHWCnXtFsUWNfubgmkLQ9GLjbU2MhlNk
Wb5yaXNAFpK6vBJFCQfQqiITiwIvJ6qFetppVfcm4xpoZvY0r+Ao5AhRCR6rt9Xccbw7p4tztyL8
sToSJVMRNWcja+yvEpwZ9eY1Zy54OgkvWBmHL4x5foNBGJJwVjW7gl8zr84qVhaXOqVRLjlUqQGT
hGptpXrIQwrrWr8ql+rdaBMvg1QCxjIHsX1DWWnxtgiVlFVPaAJt04mL9LTRGFl2x4zutoAe7lQH
9RqFkXmFdw1aEvHC1/j3YXNoHSc1dQcMGoe8TPXGyxsH7Ls3kNixDj0FMBznEF0MXdCAjX4bG0I5
vsNxY/3zcVM0kuarwKy50Yxlp8ax9bUgUDYuhNY8uPoj7mCKh8Xtwls6yaMkm97Wbaz6bEi6bkfj
HADNt2VqnXNmTDXBEq2vcrKtgjWJLLCQa45CxuIY5TI4tvAcQm4nRbHSf2pYvZaGu2S7CZH+gd+v
MqqYLVsXR5yaN0H95Hh24jOxslx6L4rEd0lzVY8uxjxUvwmULqCl88Nu2ZPeP4yCbuv21qrouJG9
JpG26pRrbHJs4tDvApKBVzMVOZ8JdnKdGfPtJPe2M+oByUzwet5R5TezVEAk7VeabdNe7PYI2h83
Sgg/Zsc10XArb+YjzXiYuHOWVWLKrCGlgiez35/d8XTtsdTH9ULv9td4sIvnyTo9tfhlWF6W4jTt
ZQpz8+rf8Op5SAk7F4yKkGI/L5oJPc1dMQdJXURuULs5R3r/k5sURpigLusJxzinm2iIm0hhuYoe
vOC7z85aytRxciztfFl11+yGV7HfcgvK0xwiPcQv8RezYzVd3tdTDmF7Xh63e+MOcbRbuTQ00u37
zZ3/oc+rNiplptkHJk0yMx+gT2CC0Z9wJwHprPGBKQHJnLamN8g6pbgULkrGdq+76+QwyK042QKR
D5Wh3ItBUuVsOvEt5SKYYlna6fgwxfJ1kqtyYroKT1lovAjvLTs6foPFDShA69kIkn0DS4Af/gJg
2GfRmgKen632gdxeYyNDFV0tXSSKNYAFn7CYu22GGUfy/i1QQ4yXzZb6AukVplJLhuHbcVSac0zt
nrjxswOQ+QtT1Odg7Fvw1c4DKUMtLRdweVYMCwGz3lHKZXJc/8sxM82YndKXHGSKsZg36wqx00lb
bLBC7lhT3Wvc9knYkoiHLVedDdL8bxDpm2ZQcku6gyfp6aeKJAa3yAR28PLJNaznC6RDjjo70xnK
W74MpH4cckrfmalDgtYbOIZEZkAKUzFQyjBXVnRHIgKXsyfVjON5oY3B4p/gH7+rZajlZs4xSE6K
exZGLWGeV2IGp5jDxjTwfFs5+p6XbBq4mFN/aHaXRbcRlJeYTKf7xRVvaXK9hAwx8C3gMBQGDQ3w
Gx2wQLp1uS0agdLwjkkNlHrPPbADe2nkmVzysjH882w5ZzoVDrcwN9Vfes7fCvb4j1qg0dWqwHb7
tq4wAxOpLxqaaRhDQd4KCn+Xq3r1++8O3H/dQxu6WaayEwHPmyWApn7NlMIFhodQY3xqNO5Y+MOD
GFxzPt5hJ5a7BGqrzXmXfXY53vJIU3uygO65LuJdriLD4yPwzecRtgLmJeoBYUQMQj3n8oV0M2UG
/EQesoqoqs4Vjnkuaq2w4rLPxLmxp4x+2T81ODDK+ICUFnlYE5FOWuoPRJLl2Aj4jPYVZktuVE0J
mViL9DTYyxq/BgwB0Cx2f4NiNGRbGHVOxGp4aEcpmgW8uRAfOIL2T0NaVyEFcCDs77EO6LRUVLtb
y6fprWzBjj3fCsKAS6aZ1lfGVSVWbG7c6On+Em+iWD1aos3BXN2nplzpohx6BUF/ndAm6ICmHbDY
SCVJsaFW1xIfrcuTQaijlAuj5LppGR4J2cxXfjCAkn/nxvKDENsCdEyJMZjO0r3vXZAnbPNoAxF/
dcEegB0P3Git966jbLtRALSg+0UJwAJyBw/Ve99ZIWsowoEI5lW6iaU2OW82jcDq0+CAYKggXH0K
gyazTttEcIVXmU0gQ70osuOg2wGRocEjn8f6nPhkgjYXbXHQ8TDDBg06nGocX1Y9SI4ED2wbxzQp
G5U4KOqVBOok1znIB0LbC4yiSIe2NgEqkaFBuHjp6ruj/mFTN+nYeJj/VJReQUNMARrqsNL+hkbD
nhfHBVrba6AZaBmczb88WSKISCo6WyKI8rAIcW2jipgIEs0URRarwVvsXrsBI29z2+1+Q/4fozNO
K2mBkiDrJzKU7Rq5B0zua2Ti/UNC+9s8edsIqAmv7uYmQwJUpqjjvytyQIeum6d1LcluBlPkznc4
h/eF8yUibs/Kta0NECnI6b7zA2mY0ICLfjRA63IZEzDks5caI0OtFyKioxkwEXrPQwAYqn1FzhMJ
sBh/z9TIm3ESAr9EjHC2uw/tyYo43SRt5+W8Kw3iUiQf+AVRnhhPNsvfUxqbbqGLy3+rxGnPkjfG
gsdQdQcc7hRfKGLVHSn4cya4jRM1DqeAR6U1BTVEqhR1cLEu1RdHq8cO3Pzh4v9FzcpyvTUdVI0O
QqQIkqa1Mysv1Diwia0StmHlwHIu3sChpyFXVM5wOcmlzC0gjcMdVqAGuHn4kIwtQFBuTKXlOp3k
PP9/gZKacokYNCXjQEn3m9JP8FA4rU2IXVvKC5Wwxc0ZrCqD29FzPWd2W6zpH+JDbpt/KyuVmd2m
WQaYFZOIzEsbiOS88aTSwt6I1VzYX4VCjq+apfsce8/TXiRQwo1EibITPOZa9MS0J/Kk3xBJ/WfD
3v81iMBoZQlXduFr8gq13X5tWDJlAsIEjNtssEhsdD8Bso7osbDEVEhA2nijXUclhvLeRVrQOg+D
XFzL/wUJlJOIr3t7R57b7bDwz77uWZzQU0YsJuK++KLylhDtLom1VyowpBIvTtwWp5bsknyBom5T
rVuvdCbeslrOfmfaXBc3Uv2CpxNijFkgGbJR+UuPRbnrFcZE4u++WK+FYDy14C7K4z8+QSAU7mgZ
z/DKIn7Uv+7p3EHOCMpUeY5c6traz/c7bltkTa8deEJOj3dENmgDJNggw4Xy3Wsd/2OkPEwjLx9p
vXumFamr3pTLuH8hNilRViOSR1uihrCspby6ZTy5Tkd5xdBNJCJDv7e+MZ9BlxiUX1mx8FD+yXno
JRcROYHMMCS4yKzNQieAaIAU8XgEer0tnR+JAMRMFxDwhPmKDnDM1eYnEYT2aDZ7UtqF/NYNByMS
166uMkJLgkI/Yylsr765w33HOqe/h5CqvznF90mUGuJcoOOTMD2fLtMZJTha4c9GeGBqX1Js98Ce
3u4rixlTd21Gkx74EtmamTD58a6jY2m3bM3/LeSABOwUjvbOxyPKzgMyTua5B7dpEOnTEmi3UYOm
BG4XEKHlalMTv3X5am05yBFHM7Khb0uM5DmPTOEfi0/zTK/JI5WYAgLYwdBugxvLAehdYd1ZtJBx
W9oAoQD15GxkL5Nd8nPLxUMCoi56P1GZ1Z+MrbkWswT/adrtGxhax1/qR/1hybh20kkND76yINqJ
saKnd2jbYwcza33J93OAjXheHdv+y7vqsFY0aHGSyEjvFpktTZcxcSQdd8RnV7kJsMWtUwnMyuD0
TTJmJipnbU4EQL6/a0m1zuABz3z4ipnNm4o41XqaUs/tIw8b0JUVJagXIs9h8A/8F6i4Evp5NJBf
Av9tYfp/mKsLBz+guHdbdkL96hmCnuYnBs2Oed/mufq9YeHbJjsrX1hTZot1m/aYVBxf/ksjioq5
kCv7LSuf2/gVargVp52sJvPjSw7vl7XYQHIvlKpjkZW+0D7a8gmlwPIQ+BEMgEoro0aS1DDTaJSL
xr0hUrDbgyFkZKVgQbmP5IULTxd1N/kBGJOj3EqBMkvOjkhWBHzGkckhRyyDuMr+g03rCrxyGUrn
VEenj6g0PzTe533v5J37Dcl87mRmft0NIu1Uj1Ezua51BQktsop8/qG65xZchIK282tntv1Qu5zd
TxWq4lb3QgPHXMKUZ7ME/L4NMyaDWSMDlS1wEAtsGRs5ySPiYqY7vzdmhtOY63qHlAotiMNyDIqJ
CQHBxP9mXAf6I7OYBd1LPA4HzF+xm2gezFBVvxg49J6P9Uj4Dx8Nm2O6qLDky/MS/UTRwPFWpWdv
NcCcAPy0zTW9ZslryT3MP2dtpZcLH+W4uAw+Awim4KDMnOqxmb0jELT5r006PEhxES8Si9+DlTx6
t0+/zeq6PMT11bqvMnuszLGN9owbd9+boXGaJu+3XX1Kj6ys8HQgi+HqJLy2ku6iWy+WW0oW26Xx
Gq9HXnuwt8e16jkxuTKWdCTI594kwRTLAJREsjxdC+MjEn68+CK0mPZsQbrvHdPZLsCODDoICWL1
76z1cduo49eVXPNo5La0oQDW6/6zDzXLOheLSLwQl6g7SVfzGE1so5rKcNpM4wXagiokozh4/zcv
/YBXoQpiqdX5uyZwWltbeB99N9OYy4L9VtDj9jMFVU0zGG3G8yBEupQDyXV/0ibom9ny8NpIF3Xr
ZVjY1TlUQoA9UCQWLB6N0O8/BOAuOSDQx/I/scpOqoVVCp+q0MENv4dmx9fR1E9OfVhGKFxAAzmE
jZZSw1Cb8e35GE9WlSa+B94LvKRiKjJ+8i/gixzYqjIqa+/bXUKC1OotU2vj/lBvTWxJcvzE/TBL
hUy13Xy/3tYrZ3JD2ZnrVneo33RfcV1ezlhNsTblZM+lStQ9dehvm3iaDY426ivhin62O2Y83vKN
gfniusFROWy1qAXlalydvxKvsxNk2c1ECbmhAzStXL42Y4hdGSTf3FjrnBTi87YLunI4YhsIkubf
X1Rtvn8E619ZmyPMYs8k9lQ65d17yoitzNIbUEFM+Zo89Ic5zi5LdNGmmJHQosmU8uVp8UPDh7go
BE59SVUs6w8GT+ABfFN8+E+0YvgDFhApsrFh9WUTDvK31L8rVazdSKMEPYGFXXITUEkCPwWU6NSv
NCyT++kqDWVVDDHM3FtGpM0SU70WMk2cN0ODi2lCEe7KLfMw5aSZkyNBzN7I7gm84bcgeGRyImvg
bhPW5fbcDC2+M41PbCIUFoUpCGKjmaALmyoOBPKDiu3I0L2JYVJ6L+wbWoV6ThzsYWvmoKFtqSeK
XZoEps13GeTUL7wCleTfhGnuUHvzJ2RV/zH3Gxy9E7JznL0MtKqrhF+0OKhzMhGXHQRkKjI5Vw2D
mX29PY1JAjFGWEB8hibN9PgaK2O5j4lKwC2tcivL0rPe7I3r0NMUyQ1472Fk7SyLK4iXTC2NnE1Q
EFvuav3DPagckQebyOJA+Aehyx/4pSC5OwHpaGjvABWaL8PiHhSDajGOj3Hbo867NezF9DeyVBua
osePIHtI8fryKDwX4IZ8/NbQcU2WHw8gLZZpuA/QfnzxehRE0FfNs0W+VOfS3IQ8KsnlmorPh95n
Zkzj0u2oYpo/HdlVwN3HGynbPpRbkzhMBVNumKaFCeDhBvqOPWIC+wP1tei9p4dZ0AeJwU+Z8xTF
j8MpxGN2Dcuk+yz2l70sJCpknFXV96nxg0o8fSQ62pmyCKL2DlsZBk+cNIeBeEl2y9G7zW0Bly2d
gypMwzBIN+q5Hb3K9h5HVf8q5Ra8OGvRPFNtZxro8Lhse4nfObaKwFPLYG3EpQ/vR6uN2j3ynJI6
2Y3X+wz9w2+sw/MtcYjAy/R4gfFUPDxbPWVC6dDCGZ+Rnl228yMrxh+quZ4lr4o+FjGGxI4yT2T7
D1/KfjpJfngBmSUP33ArvzQlSl1526JDmBgWX35hgOGouDRy9BidXgvJlR10hqbIAdHi48zEdyLj
8fHnOnwY95Inmgv2qU2mzFuTVW9MZMycILrp2KtzsesK+Ez5YVJevycrQN0AhrzMg7xx2aeU8GuS
7WwdYj6sqaCArRLE5ijVBfH4qtmo9EOzCmK9Kyh/8AuaWak6Ef9/ipmvpqZrmSbwbZVaBcHwLNxa
7QLGPBu1lb/s1TubezfHzATu0SVlFoCexVYRtPCAbv71wH2hAWoaO9OLu00wZSrUsd0TPfQ2v+QK
tAN/Z7c2CTgpWqzKfHIY2ksuplkZHUW0ETyVFH/OC9QYcMyMr7QTTIWL9fxEPuVbHQZKoEJbYJRs
HEhwBwCqjMmK2ENrz/v5BHvf65wn43rJPJ0Ss/p4QXxV0JwDR0sWSAogZM5ZLPFzxnCdvOxxUDVv
ab+mIVW6s1XkFIsg6tfwTnm3oNHzQSEnOPRk6P2VGUg6W8m6rXkCk1Zz5ws7srMCsLh423taRKU1
MBhwqd9dR2sUOrQKYLIPnoZtsdJwGvfShyOSA1Ah4x7nCf4XgYihOnaVgVCcpB4aJrBT16HHzp1G
pYu70psr7vGWUUGTP8wnyUxREM4PcIhoAzmDvHbSbgKNIsoFeYjmjdXapi0eK6ONHzcKcuvCqmTo
AOxzm3VAjJuNoT+SWEkevHny945FNfWKqdZXIvUUnne/G2bJbsVMrVPTR7QdOACTfyvCigdZIEmR
PWhK9ud89ExT34z8oM52jgeLTw8sxzgEFBsLUvxNMyByUh/WjKUupti5TppL4ckBO4rQyb0w8/8Q
qqUD8TvlvhGzuj15F7a6dw49Phb00Bm/PgGmwqY3KCVjIwFSvQbrqanwOIufAv4vO282Xhk3F+8R
BPQkbPTXcriRLDkDedn+mkKd1CHWE6cgw4S6W0JTXZzy1aE6YZ0XswvXteBwClZ1lOA7EVoLeFXu
5LriuKBAnByI/LFVdxjEoVDsv5itWHnrBzxhfn0leTywLzT6J2L4M877zB93cUlhf3QJMAsia90e
Sb0zW8eR/raY9NfoXDRw+YwwXwTb+eTNZalF0qycnwUJucTueMOpaNYEuZ7Px1yGjgltbxpU3VQ2
vcGebFFuMLODTsGfQ8YMpQ+rx3dBwSAYjAqC/oLtPkoP8ZHdTcFVNwQn9fZRsfyS8GApROZ3Punq
m8P3wrYEHtTuXhU4YCbVXsnrd8/QABe8loRMOUWx7xgdNmE3rfRUcU7UZaaVsgAjRmNS2k8MvKhy
xqBbHgHl/ERw9Wyem7FGE+4bymHt1QdTI6J+s3rj4qe0Ixv5P98jwss3TK0UeBrgdkVjeAcQ4zNG
SlbJpFA2e17djij+975C9/kvZWmXQ+GsFeOd1IdTiPHhZfWrrj6neJwp2V1WU0q4t+iz4Bim5282
e4LFne9B8YkJ+oza7apIGYEGiaEQUByvFWiXwJnVav9nfY7+zWaS1+hVhwLTBCdViX774/qg0uxn
5Y24NQZQ6sQbzd9YtV3KXdMwCH3W6dWk5lrBqA8gnWjCf6nFs8kLzQE3HNDK7fD8Dxu+JXrYP8bB
b7sZvQcwo5sYmdsQTNpfApAY8hIdGZSjF0jgwApV8q+JyvWuhtP94KOYYLcGz+Ap5ZX9FVw0NwiG
5HSE1YaQOCSTPogG7JRNvO5gCATRmo7MRYojUnCWEa1hturFla4To2xmfvSIyhGob9DmJFlc3ZKb
EXNV17rbJ4z1SiR3BVsnDR95tgi2S0y1aGJQHeMHnMEluDl2TZV2v+/wDcawmvpI9VkH2odKABIX
hAtX4k9Z4MSMUNHXon/FCDkBZ8HDX6SxytdzrANeGkQ3phAYaVljJukkRzBra39hmt+4xhmMDefJ
hBoBvAvrHQs0P9KYwUwL/a5q3vmPtm+DCebEDttClqTrp9FuRq8IzUl9bJ7bEaqy3ZTeJY+BLq8m
4iCmK451WbhZkjcVLzb7+7uaMM4woC7ZoLweMxEubYvvGtlAr3pD3Ij/yTB/Ey2GQvlN3975618G
a1+A8o4nwVaSSd1S547MTCENOG3ZR4QWtjzTCoQp3DGfsDMnePnmm8Ey+PUdoLLEZ+Qv9rxSiFLU
aYRXx3mU7r5i3sJIiXBfrZ3tJZC26F/Uhz+HuDDxFA+hXM5pNR82pE7cC+29p/qziswdrDqAhlr+
21hbLcqQJ3rFnLKsFdwxdXP+LMKmnqfbVFcgjWm1HCWFxB7sq40wsZmf6M6fCXTmRIImbrF8pYlM
h6BYsxkPrPI2kvoF6iAACqMCiAnWgeEjtLzvg3IYxff+V8UMw7uzSTQ4HhX1sZjKfaDXATxV0rE2
4ce8dz6opdQRGO7kITFpMDqIeD0BnFjU3KlD/ZJyAjbUQG2tXXx3GM0A46z+sspstfl1xw8cik0A
SoeKQpZxZjLYArfs0QYoAjx2sRr3cZtByZN3J/2nSDN/04jrx/lUX9oKti2XohXRluZbpHUY4wMg
VVU3A2TJbEXWBUaO70iWYKFW7xqnxvBIFlfbYN7kZfTIdYqjvWyQv7nGC1odlY8LmVDZ3Bj/t+Uh
PRdgmAepIOlLrEjSFsnJPfkX9ACJVbRMmLWv1THkXwusj11Do+JOEsd3pAyLo/C2ter22m/7X3UW
SCmuJ+2kAA3qHVCzm6AuXC8hidGpE+MHctPm31S0ovjYM5GSqbDPham0V2tY1y3RHfiwlxOEzE27
U2MrcfIjFi7CGJZ94lGYxb9Y9IutvxMoEnXbDU0gjetH9enTQj06jFNb30ensAuDOHTjAUYDlIeu
PL9pYA0wH20E/wy4F6Fg5AawpPzn6IzYlLjveZm8ANE/VRuJFLw9mJOL79xRXy/DKSmHYtRC4LWZ
E7qGmAdAtbEGQ3liIpg1euYQyc5zK1IfVaaw8W351MEyJR5oq6ny3m7BrIAAsq8RC2O6gvMi4tSQ
/4DbWiws9zYjkBJi7Hl21CF0KPO3gcoDZMMU6JpI1Ygt3iEAfQA+GCkOfm5bGG2z8KBIuFdEGz+P
BqXaUagPxKaSR7tddNHovDYASbVY7eVeK5BHjTtcxcZo2nhfoq0hGXzjZ2Jbw9Erfm6QrJliawUd
Bx/5I9S7TfqYWvtRu3u7M4dR0UZ9fnVZiqCbkfmkHN2yeHaSC64UjK0iHBSB3bFOktKMnIaqcJ/e
2kSKI+D8JzvlcInYN1gIL7A19DeL3u8olEzDfDUyx1GdWLi/GTE3CgI++uEs4w7FJmYjyVEl5A30
yKKHD4RRv8WAtHQ11iTMmDLMz7149//kGqqMvIB5R97nO5ZS/rHgDedKXOuUvfwulU2t/JNKoEba
P47ctInIYA0D3Cv4OiSMPo+yMJlK9RMlZEW1BT/UVsbCcFywqFojEGpl4fb3FzjXjMnYK0N0Wd8m
kOnqd4Nrwl1sH16aLw6ft7WUagWC2zHiK4wXemWyEQ6PiuQFRZfzoJqAdEPtYxKsShNJeFkYUbq2
sFyB9WLLM8DS0qWPRCyRs73dr5nbAYL1+O/8WMfoXRv9tg9Iyek7xiYcT0raKi6J41NjHCkVR18v
+VGqTxWGWaC/p4+zZjUGnnjW21WX+lbONgK9aDiytF5FFZ4Yj/StqBCknvzch4ILvjEeoplIryu1
5SuBUTOFNxDqoziXw8Ck6Hx/IgpaElB/gO4iUt7pmmr0iX3l1Z1xh8v1l4LMdoscxdOxn/hpTfNA
I45SOl9zHAiVtdniCTXNR8vL1dJJ0+5KHjWo3gfsYBexHmt1x/Anauq0/dnBEPVpVXxAAZ3OJbr6
rtUBoCsUsfwJXrRa64dBmqhI2Wdg2/RzRDZFNtKRDmzaTiHcGPiauNzpp/b2/O1Z/JK+mPjhTkQs
Y4OdUsg5+snSQSAnihqy4XTBwAF1UHIDFCCpChC7x4h6KBCV6St45s95caLaXlTxkOPultBBcsUL
vwu6YvEdOL8qYqxGaEYvIbAD/tUf/B6thQFuYvmMWyZsgCViTP7QAeAKiJyWj67srbJVwf3OWNsH
8EAIkgwaQzh721x7CQfsdTyNBLbI9zmBjq0zaTTQQttTlyXj/VexN3nG7aUSX9JRK5kqBshFNm3h
F87gjsPaNA3R82GQX4vvLeFMZNpEVgDERplv+TWTN8dtY9Bbo6tXMeGDQVWsw4Tqg1k/IEiVjSVX
fygmgjPIWLirlOGavJlFY2bZyK8s1dgwMyFvbu8WzKvGzVUZRivrIGzQs9226iuKlVq5/G/xKW5I
1b+CwtilzI7+AnxhzyV21s6w4/8EFqNmZt5MBeNhwGSp4guzgJRvosrf3tJvQCYxp1oeja+2u9Y3
P2rXlrj0H+qLTiEcOwOH0PsaNGAu9i32U4Atkj887LlngW8/mT5MxQ0Ysvjd4gWFGwmwiQ3N8HMm
zxGLV48O6nlkw3jtn9OENaSHnlyFhpXEw195k9uFzBEGHpZMFWl3yQuOQRIQ81XjKUga73Jc5U9y
Xhsp7aF0Nrv7pjPauRdehG1YoBL57fw7Jad7D1UxKo9whcSvGAJ4RAJPZttzKxwV3ayId8Lxxck5
73x6k5YmB65Z4FuNuNV/RQnmUcEjbd2Zj8WPdBUFdiWXIcYkXHrjk9OqTsZov6BfwHzYN8lGdK5l
39aUNK0doQiJq7Ujoll1f0x0omw+t4uhtwfYd4qGClLI/fYEe3i8S2VeWhLiEJ2a0cCSnft3oiPj
GbfLkWgjaCyCVJ0rFzW6caDFAF5LhRwBd/wRbtjQd9ytTGJ5SSZXUlA+KhDfCZIZU6+Cy2VMzLKV
l/fLw9jlyG5Fp17wkAXulCzyWrCUojp3vO+96wA02ZmcrdJU3DnvjQqmyul7wJsfDlCfPcaIpBey
FxjJ+gIRhPuhf9x76HkgBLzXILSQNQnSXhFd/us1DOwuGXx7sqtTIAN5H4Wf7wJ+0koaY24p4LGk
453Z2H4mDLadAKZhe2mHUkDqkuV37PozVYSieq39y9gwRps50CHYZoI837/KFbV75qA4ZnflR30/
57amnycXJizXvKjQxrRRdG20xadj0bFJmMnqnk12RN1dIqX810/thmSaJC56FQY01FSsUJK1mQwB
XYG1WYzUWVwrEroHqh38yOCUcAFdS/F61OThyEUrHLoXa0Adgry3T+D4MJHXgaNpFvxxrOjUjomF
E56oqxzv9zHR4553HLTXWpuD88JISsroKPvy0pr5l6BkMVjAEX/QzDkzigTkXuf3uMxqQreAlEyO
qgWrAii4jfkL22HYOpxaK050+Jg2RL30hY8qlZb4O+o0ky+puDH9FSm41ko7/VqARBibeN6eTQl2
TvRipnhHpQeiQNfM3xp5T6icaYdyLT7fBZsmXYJVp/5+5Pa3tQCZJCzVOnW9KYr5iTbyrLiAt59f
h6UBdpe4peAuCrjSHwA/+tP6IBhFsKwKSQVj0Duy7ckFib7y0ny4H4/+7PaDaN6ZoFw58vlqTuxf
t4uUt0EK41IfBhCu+kP1WgIQLXSSaRqOjrkCGMho2V93dOHQup35DLI60/MnPbZ60L9UXzOVtzpJ
Syx20i1sOJYiakPREapQfH3iTDZEOp+bdLof5Nz6Wy7/Mq1dEIL3YNClhuSQECTcqydpxueiotqV
0jiz9jxxbSwne2C1n3eByUo5Sz2FdUgfkB5BgrNjH98Jq/LUGO25ocx2txp+LOxeFq8FZF7IQBHE
pL8fsLjR2f8uyFY9gV1iXbAwc56fNga3z72tNQTiBiVLdurE6b0H+DZY+lYPBSNLOIQDdrtio99I
rW44Wn80dnfnNxN9NYydSMumlYRbn5l9fTgLYNN36jUwbHO2Z3RWqmmTa7dUgQS4AyKFD9HH+NGy
lKSJ/Tcr9cPXmYUIZG4MldA95N7QNvYGfwsPiwbHC7rsrfeooHzrER/ZrlOLEsGq8H0qwaDravWw
dQdMOpCVSvmetJYki4lVpBFPVOmD45nimOX+iPV/OV1re2D5s0nNRNDNCCryeYZD6IqEQ2Kkmes3
mhjHVKfY910g4tbhJRYabF/D4sha00RVsNJ5w19t7CUj7/g7+w1eyrZfvynw9+I4hd1r7KDXkpPk
sITnghkUSWnHcrpuDFDfI/SiFV74yl7tz7YmOEL3XXN/Acqi4HCZdhkLMG22/jQnMGWe/Uvzw9YY
ofQbqcOr1U1pI+n0J8XwuqYIpTz/ga6WR01giukzJpxl5zLVfj4ZbjUNU/eIiYYzdylKwtRRD1tO
l4SoB08WxfaEcZmtWJv6BmYon7JhTj7LUqhUpfnnuM4VfZWnmH2hXvggOilJOqADf/tCG99hkqY0
WAs/SRSxAM2aUksIcvFiR4x/MpX9zSTp5lgOzhN1UwHZDT8NK0SaPayCPK+0DoU0Fx+MThn6DK/L
iyRjL5jPNItQvKjhs9yNyFfwxWR12Fqu2eFHejHPT+GtBf/brAQEcwNiygACrsW7PDvJT/m1zMTI
1LdE1dvdI///5uSXJ1ROMy4zHJhZTU6PM86pzkdhsnSs9+zv/TeUtGxEjL6LAdbPitmOmmX1tcix
eTa054nd/RQNfvXglmtm4cX285lkjgX/FvyNnJ8mXHeav1G/HfBpNSB3eMopNMVn6NvXATKA9GT5
H0iqKRRD19/5h9CMmj7kV+tn04zwjMZc02LyOG4IoFQ8MrbXyVQ1771lC9fadgYC2KSsZ6PqSZ2v
Cx6Yv2Z1bMsOzsfKqtQF05FkxBpQNgkH9zTmQQtIIvKXibKHthGoEl1xnWAKnzMIni5qbDZdNg0m
7q1qX01wSn/DsfGJr++s/bBrxv5LCUFl3sSw8uYa3S3bz9LY7xUk9r3k5lc7whHB+ysiPz/iECOq
55dSkyx6gB78tML8afT8qPKPCpwEn/2dxQJC+FPRdbUUZV9DqSCORwNeoVRou10VDpg8bagYNmI8
Bo8EoawowMI5lLCQl7eq3IH81/zLzOjJHaprhTsoBG0LSl1m4d9QWVE3LQOj13nXAILTeSqORW+c
iiF1KNv5Iwi4tWTvyqoUHc1/0nBctYa8zlREBlk5uuEGY4pMUEQUzS0mm7V0HlZHUGqvIMEuOapb
HcDBonKUmriA1RGeiJ1JRGQ3c7UzTd8wPEVdlz45gA3E9J5AHHLF+AZxeQQNYU5TB/Ygi3O/Ax2j
6/AVGFz9blCMZDTJNPtzLSDN+L0MIV+pZEZIIuq0yyPXvn6oegXM+N+oEX3f+VJAOtj79To8sIQK
M/SwAga7H67hjA7E+Hu3dNqSG46PlNDEhkCQwa6EpvaKCppysdG+pKYI40TOw9UN/vuOVGO9P71Q
wIkIeUgA29WwBuqH9KcVrEDuCBscHsIyYqTow2p03dWyd31CNBvPgkWutvA/wbqrvA8s4JNZEbOv
r69sCfdlas7orhGsaZN3ykV+s+pqxMOe+ntmnmLNhHeQZDkliaIdaCDrTTgaYt6G2tt9mvWfB4V+
BciY52Oex9sdryehVn8nAQssF+eyzG4ZyKwaPfRpESFuiLhHundEtE+yB5axm6JSuXszyZyOPcLH
X67vtbxts4OTx9el9wX9itOJdrMAxSd0zEDvw3b8W1ti6KNs8K0ATWfC06/HWoy6mh4a+6wL9T9m
QyFdK85dOxzC5BlFpnWvwNcv/f+kQaGY5E9PtL+iZTvA2hzh1PZL4taGLKP2wBYTVtxjy66/+rJD
QrvXurBklZaOtvMrMOP0O5cu5+CHxkyelGpZPl9yhBKYP/4t6bJdlEDui5rzjdIpl4EG0xRgce2v
TbfaL8SMC1L6doBAcf5tFsV01Wp6tBGSU6j6zzfY2Cdm/Pnq0VFZaPD4YQZkNtVDTm4E6/EXi7JX
rVpx7iU8B1aSGNhZSReazR1zFo7aJZW3Pmabqm3MGyUHFj8Wdle4FkozOrbFz3Uk/ho5wLyCzTb7
Y6gjVsXsAl49VIKKlUld9/QDJghVQg7ua/91e5l94FxhZr+LEvBMoBgIZQMxmJkds3QBL2SrhZJb
YvyKcWGxWW8eK3v/gmoe+X5X6B+NAnMH1zTejY/PSyTtfHVBnFhfTcWAeqGBICriRGZ+lkKb1Pqu
qmyVDdxwD9E9pjIY8G3B/EZTAJlC8/cq0fcPz3cojHkDC31J0G+2G6m2UEDHf3DDTwsz/ARklXqc
Xng64IIxzRX7TtmgB3dmeN1ESaXoQMGtzuDAbwkFzmae0FliBkBMMQgYIQOvH2S2zfwQc2qeeupv
FWb+CWDIYMuegeSDUoEFJeCevvx5ZckrXGEzYDyd/97pzte31+0XSXeqHe88KWaBPpH9jnI5w6iG
ZMKjXg6SSd7HTKnvBQ5b30hvi9rf4fZikk9OweVxO8t+kluUzymEZuUWXFY+58aRZN5j2sr8SBjm
6Z95qV2lhPcvTp22fvobM3SU2W2S6ORMac4FT3oasNyPKY8IpEZhjVqcV0k4JHSSqhGYD0oPikJG
R57nPBmR7NCi8OR/voTLwDtoHx48ZlZdzUGFnrcOEREurG0gT0RQRzvEFJmzzW2UR/HDR59L91gR
ECzDf3t1VpK/npDDZtqTZJzhhBHNo1ncKEHPGyJayRDOQHBfFcuInP7nTuXSuV0CGXP3JBNLXdZ/
oFIQNr2FcNa/iNImgcfKDMzcZvgndtCsWEccqQQ+1TcHuN+XhELWW1LKzBd9/lio+W/XWNrrsV49
YzGT4AcIs7tN3+//L0YdkvHosd45afYeungb10astV4siSFlfYMKYT8VZmL1n6ea5TWCGxfpv3rH
0ajgngxhaCBsbvfAhSQgHvROgvVZ0KmiMvEk1hT6gYyMjsSLkJjCnjvSRvzoIo2YWLDlr4imhV+v
aFw/oFpwO5OF2bZNxGNGzE9CGcNOCw3lTUyGTtSUBAHFKmBARzad0lWZInpsBDRqeWJ/k+LdbtnA
1sj8fHtGjEsCPHVq1UBxd4p/vJXjED3d7gdGT860VS7UIUUAOTPtaLz3Zg/EUfMIhUCLNiqN0n5l
gEQ14n6kf19Fg3lk2pywcJD14s7yaqFDVV8twlIAuV5H7QRGNTB493XwlH20e5vyyyDC+td2CGYt
0bVqK6BEkyWUqy77GOnJSOOknVwdXD5dlAzv1umwNx0Ix5kkMdiubUMl76jqsvbreLKI348PdOPn
dX3xPVpky9lVDVY1kmxebcKPKppCqJ8QbzKEucIF1q0EXbnD+ztOkh7MUSxoBWjWnMY0xUvtBewZ
8/US2XdAbTKgY3xz09p5BBlOJ70KCy9yJYeHrFpSlSgBzuSuCv8No/wfFa8cTEPXg/y2U3cWHJDk
HV/3B59+DHfGuVFOLuUKyT9iBGoKQlok/paGp3IlBLuVh5JAF4fA4ELJgUqe+rqLoKO8OSHj/irr
Lg52fAMxYSA8OZtKEFibN2aTjZPt5oYFMnHQ+xI3S5zP7aXLgFKltLNvXj3Cp5qGDuCc6O7ycPQI
96TS8Nk0AQnToxyhSrEz951XSy8yiY/6mqhKVhhegeYwA2l3wbla97qJ8KZZ4I3+0B9cdhl2tHnd
o0RTzwKTI2zJ4u8FXGt0fldqZVG9wxywJnmnRyfienF0hWXNgH3ebYgKoOCfwgMtcHCw+kNThUzR
nLhOF7KEnt86nq6/JyNruhTUA8HRaXSWJPnsiu9NldmvN6YbrP4TksmZcc+wi13hUXSrBxezSeEQ
LgYaDS6PoUobXCMNHGQS3+qNMpScV41FtnOgModx2A9MYv83Bt1VFq5wYe+pC+QAPg1tJiHH9923
Fp+JyA1SoQzgnm5A7CLrPujTj79teFtniJrJSaJO+aD/gIVIDG4D9x7Dth3CLrLUKg/bk5/SdD05
ItW/ErJ8WVivZ6NRlb/4WC28a+so5PlXzsVjvy6lxJDQol7aeiHwh7QzYfLzhBPbIDkiGyW3DQU2
txJDr5XLSbZ4S0/JaA/RzYFTgnVCXWUhpFz30O6DDZhEKSMWdGntSDwukTegVKdDhN4nn1wHfWaC
Tv3nf8/r7rZkwE2zITsqZkngLHPpteqoOR5ET/ZqdILsOfBjBSehb773V+FaQs5J9DGljlXOWcZx
Baq57g3011MWkQv106NBDSg6Axek2ly9NGotXOiOCdtum1T3JFTFGo8MTdWwtg5fQ3DmTZadLuEi
3VfBMVkaW4Hnz5HJMnmYFdV0rFEdQeeSeeRblRTTUlOfsdRLvJTo1rD5Mnw0e8UJU8ZvQE7v4kq8
qCOtpbQnlhx+A8eM1rbTQSFX4fYKE/8ZRtWUCXQQ8DZRyRd7/IDRMEPcgYfMjmZ6CuoyR+WK0xAD
JyyZPzjZ8IYGXsrAP3rmv1R7m7Rc9GbKGdY1DMmuM9xe+BsAUg6cilMWOTX1J8TK+65Ybsc0M6HM
C5F5O7ylPad7QxK8fj0M2kZR0+WM2nSNI/sTSgq8xw0GsKHLiX9LRjD9a6Ffiqph1sYfVVNTDspG
6nXXQIWkcBS0LhcaNCJe1p9i/c2jDFK9ilbjifBLc/TcwMSWkkavueqn5GTOUumvyPZeMnq0UD+3
/Tn3cv3AvcBqejCypOlEb7j9EBUUhDLMNhUl+kLvCV3doqsP8rSCyHlN/pkIRlYYudtHEfpI1/Qx
kfqR/cXGsOJbzzW/6JkRYGLFZmSrE4+RQpl9s38ROKqW36TNuqggbPglvIaB+eqqGEfAr6moOhRp
ZPS7174zNFchzd57TcxcNb7RokCekrM5DXqMfBByn7Wwn7+cHavjw85WWEZ45gneVVvpztst6W3d
MSWZ6XWQCOJ1JTidnmHHGh/8haRcIHQFVbumQMFA480X36sfRwbSBcVZFz9/O4hZ96GYvu4E6Okm
1NoZhyZWTK5CpV0jDocEhSbNQa8VWqSPEaoRJPUunavlL4AvUBvnAT7gNEbeMuYi1SaNjJGUxBWU
DrhXFcpBnRdo5m27eETdTMzpn77EguAhCr4ofMjDKVn0x2WDGs4stVe8KXrDR1KD5jaEzIXi1UWR
xefOz1sHvXCMBJrLLPkKz+Q1Cqu9E3kqbYgNJOTjv48F1kcgTLPMHbtw9U2g/1Wc29kafI0ZJqND
vL0P/rw2GMgnXzHgT7+hT+drxzwHZzV70O5LOrwvQAtBYYsWrxguQw3ZWvPifuPKRRgXcV45r6ZM
71ccxHQs5ShKCE99ByX71e50kkzitHIm2H7fXcQjbeXkdOCTPaGvUGllAsfoMYQphPeSWwVKRC0O
TEJAagbheBxFV85ku6joHvi6TXkDNC0WpX981STmjIPF4W/grn82ynQoxwg3NMu+gMF12lC1rdjr
Cfu7+ebj+5q+L3vwEq4zWJh4vR5x85iFckiB5D2a3D9rJufpE798NFQ8kTRoh6VgEc6MxeCMfmZy
1t0mY1fejKTB9r19veF2tHmUT40hPL01u8/L6/vIk7leAy26g9rnOKppeIn71lMym2KgWtEQW7rG
YJXKdipvLNCy1q2O1gpf2cmmxBdwa50kJxJFrUW6tCufPmuzjW0OivRSooaLcm/rbGmpU5bVCV4e
NfuR36HM2r/ngNVedA0A9DpntSjF4g5Sf7AAqW7Mv/KbHyZjhvKm9h9HnDNbUbS0Ir0iKM8zJpmq
90x0s90xHIhAX4+YapazYOuj8BHIfmHp6cgA3a4pk5FKOJY5WuJZ1z1Ir+aKfAGkvSoE7ESEk+Or
vqaewKHxbk65aTooq9GLd9fERVbYFrwOv6LZdTJOv30Amlxwi4gc+9cviU01Gc8ycSLmzp4FCTpU
8OPqyBcFR6DEvtHdQA6uTM/T4HZFZNsy+lB8wM2/LD0v+KSvMusxw08OudiS5kxUIK/WegtBfeJV
wsWW5gbsEfUPqD+i+of4UN5kZs8rlmT8RCbFhEmO06SroH7sbOJRwc8iqsArGQRU8o1nhGZ7waOc
Nk+4wFcurpZofmBhh6zjYoAokoVj6PMIm0c/MYyjK3HnzWKwkwEDsFeUEbCRUBZzK678Q4L6JRCA
I9QfBPZP7jyPuh9gKQwXZZhWewDoKc6IhcmzWu298zbmtx7kX8NSkdriHtSdY7uU7uczKQQYugGZ
7+UITTn2iyyLGy9vHnQiwmAOZdagGzLazzrCjLBHeJ+EuNX09JEphfTA7vgzqnTM51f7ZFsEgWiB
XDMvq/UhouhjagfMbQCiYVvbtFxbILsRq3GJeeYHEcVvrChJAR0HC7YOfzphMHp873ossH+XPAJ6
n3kI6juEjw74vrXN5PzkrDtwpolpDmZnl1SvvOJ4fB36KbKSrZDRrUcyguoXsT4EeAG2PqbXN/S6
UxF3r90S1/Vdd34kGDz1vV3YLF1TH3ikLM4LRGgbq1IRVzmje9ysXP4I2uy1salqHG31AYPF3IoB
8QJ+1RV9jzucGsWptLGVYLkHaqLwAFiIlrixSwle4woH/cM3yiuJHlShSjsjjjDlxiI/HTc9mAX0
vbD7VRcrd8Id0Np9tt2cxDQmoT7BDGzNWkUMyaGeUNk9nsmHUCRVdEEMITiQoJc/8dVkMvuByZx5
dxGJPImfI908uJU0vXtdwf57OiWiFqGG3L4Rxtin4Kfvic7P1RD8Mno22/RRHzLcIthieq4+JDTQ
1N9W+nrq/KFG4qMFAh6QeJPtQOguYkmo0QGFZfnt6wMYA/K/wLLt+Gj/LxvFbfchQR48ViRcMxHk
wprzoDGr1+GCLhVn5ifh0j0a3XLzdeayBGOIo1jNTWWgxVluD7LbHD1SPXXVLB2Fxu3BpEEb8p3S
tUaaW3nFOUxczdK8xOfeyAFKeMa+Xpp0HTkmoWvRLqiQeK20eax4j767KRLqGg/DUuBzEV7fqTrq
1a4WDmTjOxxkZOWwAgt5lTQnSYEOWT/Z2zmcMRLn0TnGxcBw+bxoliYYZRfUL78pC2+wyyDXmQFk
xqLhVTi4cQrkiLfIwLq5DGvcy++iiY5jC0cznye6eLZg5oQ28LT1HULSnBiK04fvA0Sr9j2V9hZv
2myiAOSE3X23DXdBZKBwF8q2Ew/2rUysIq+aMGj3uSwH7h+3L4vRP6ZdQrBpr/gKMr/w1K5T4RaW
3g6yxg/I2BEZnpFa5m/4x6xBqy4qMk16h33eqon2eZvo3DwuqLaUbaT6Vij+78CpOigMOA+qV0gV
e1aUJlj/GZGfbKKojY0lkAI94sShpIYdhH2CPINv/axP6+a6vV67WgIvFngrotLCITIFLBYCEdc+
z2V1hY3sOEgPG1SsCi5y/d7knM1EqfdRIEiHQk+BPCur0wfJ6nSKkDwWa7lEHePrRGhtmO5+94xI
VvjpQI9Ipwl6GiCSSzOHRG9++VraBztKwl52EuWjEW60lFobNw22Rr8IRCM9MDcHKew79F1VUC6y
H3oZdXfkpaqUjOYcjoEkbcWkQl546EacqWMD+rAtaCffGTHuFMDU5DgiKFHj3KxjhTNxE1eXNLfF
057+RtiPJBjXEdq4oztfAsxE1oqn656WeJKs+0faMpcBYpaw9quv38/41W33lhkvic5FoFm2rRjC
CKhF+jt+VIU/6n5H9InTHB68Xgz+f+abm0POPJbIeKSseGes2Ddpudtaf2e7gVbZcVxoZKR1Le4u
JiHv0ILElwJtRE7OnmxoaaRDIT/AA7fliX++a+SLnUSGXwLumX/4SjTQ1/xdt6PlgAiNB+tAixGV
uhcVUxHCi9BWMcGhLHtk3pmfElft5UKQ9+491Por2xkvjnLbcNgji99tmL3UzGqJq5+rLNtUkcA8
vA2lUOBbEa8eFujxfZJPY/nHPOnmnYMeRYyzK2holqP0dniBB8fRcwRFAfO/Gvlmo5rie86hOX+L
poWN/e0cfkZspTooSXqbqENxEX/7Xg87d3bhGCJUsnwZL3QIMMqu7Ib9WYwHv0G3IF5U9yxcAsqn
gMm9Ls6zgGf/oa1c7VhQOBoIgu9bLgCVIZ9XEhCS089XIH8YwTRFcLJO1iKfnlln8xknmUULifaE
eHLm7bn8wX/wghd28EhmDKOZZejk4v8Ert/U+pM0pxVrUDwP3o267oYhHT5qTERACQed/K8lDwFN
47Y/W19DAExyojcY15soWQh78iJaWYDes1Ye7G2vsHMj6g6kBGJt3pIhGKHb/PdroQ4yvj/PYm1p
CbnPjraFPaV0gSoEtEJMsKfPP/lvT3lRPAguUpQEJfhqGzWq/0L775mO1MvNpoGEmt+FsDULOYpO
GEDtajLVMcOz/aZasCBtcTDNme0/n96fD4Ppe4Jw/Z7NyOIDWhRXPGXZt9YbBM9aD6rmedht2gyg
MVkhlwAaQEhj/xu8rWvCqWDODaInDQD5joZ0GzNe9TldrN9LL60nM6XMgXL5sBICNVCLLKIwAyMa
Lq+m7cWAwFrjyIFV3ajpZ2KZR/9tmRJb5KMSrR6jST5CVXefV5/l30R19FJsik1u4KdHGMtwU/ww
ffypMz8WqTJJ6pA+qZwnj1ANMoN9rYBMpt1yC2ZjC+AnWL4sJkvKg/YCMBNjGjQJTnoHwWUYtqSU
iWV7M1w9QhMFWBP0cjvU6scpd8lctcK+OanZD13vcmBv5a4iypTM+CPiDKcBN0TxcSMvKDauenze
Iz840CKuztpBxVqyk0WrxlygETnuuQOqIX6gD6qdYmI6fEqkajBNOAXCWac0IWMURjblysn74qVg
ndOdROXeKw+T3BgFap33jo/uVWeyN4lEo0fViMPMXda1vR8gokgwTXDmaqQzchUDLz4ixUKMaDhi
weuvG0OtUdwxVCZRjGVJRnYnuaoJanVq2DVtGAYWSoHrui5euSonePLHISeT0P2LO3VQvRhoC+vK
fF3CvlHF5/ZirYZpRkgfVmrWXiuxZEToRQ4fHVWKdfZcfxwUxO/bHcqsG7vF8wNEC1YaS+4EeO3T
TDjoyzuMm02GmWHUCsTVJiB9WTgY5GROEU7Gpxcbmq3JoBUTuG+r1pZQ9pLgROygemuFRikvJPkK
0iEfcu/CKRGwPJ3gifVrBHYR+8uKc3NsA2JhI5LKf+/JyGVnv+wS4krjX5kK5xQFyuPBomR/LJn0
+bd76PZQEXfHS7lfLEjon6mbzgPPlsSIwZi8F6Ete8KP9k3sou5zyqu7eVmUlpBYsJVC4jAFwXhg
/+eUeUgRlPTL4iurDSVJVmlkYC86QBvCg5R0ph9mQQktivnX4UUztAk1cRQbe3fIZQtB4Gq3ABKf
GJ4a53gd/7CWb/prB+Dm4MNA7stCPbkkpDxsrsh6FtRC5xZTtd/mNxpFdGVAzSXUWfiTJz8LqtYP
PhOar3kBMX0LFEUcSDM/rlj5Qkve3e27wakwP//GlyIeTyrbrsZl4jzy0SzJfRVaz0ye+WGOEK1C
zzo4mqB8iWxj4EAYerSFNOTI3Wemn6ceJuWEMoh/QpKxIAcPxGX8T9uocNOdDDkroH/n/6cgQCEW
C2BvDBdlGKUu2D/yy8hjx8O2bLNpyPj2JGwR7jb52om+t11FHnQj+vBAe9lS5dCu3oTE++ONG3f4
KCFU1WLAuuTaABpVTBHYmQWcmxGlvxkGDsqQ3LPvOgr4i5ogasYOmCYMhXifUepUFtOZXHwxlQUy
DtF7PbhwD8/QnWSQCzCBYnJQLDdxZUObUcmC9SHaxwbYcC49XdYUOwyNZXtnFUBiDSza3BQS3IGa
Q8xRyYzpU/z+dT+mCQZE7sXAclbo6tm98HoxPdPIJFmutsWxIfFmOjpzC354auuqP0n4mexoVB5w
hubxcxJ7aR0fi1k44OEVPg59BndmvuE4RGcC94PeFK7Q3GjyqxjHAbBRI+B/5rRkj5DJbi0jEwVF
gmRHOAtOKmTtGSiRbq9E0I7lCuvTilLGWiXS8VO6cGDtEhGDMH/o2KAHBZpI5WAjyJjUy8222mOY
S3qaP+CRc+RDZ6QO5XTgYNw388uWNvq08LTjzEKPVKej7dqE1gjMC+Aw6hcNPO7awFSHUdmnGLMM
fRkXj11Wjy4Qp2m6uBBj3T5xVsSBPBHOtBjjvnMVTty9Nj4Q6oNZhUMPJolGwmq5RSrjF8x9dujz
wub5k4/2ld+q4IbaYJrtYWQ2UDXbqsHw5iH8YqRYHBQuE2oGyxwfqR7u7Tvlyk2DONQFr3B5Ja4C
z7cIoZ1bbYcXqMewYaQc0VugOWzCZOe+oKqdSv8sgCNcnlleZbWA/jXvZghKSqFI/bcqWEDkniQz
Px/rmDVqcdTmUitqRE4YMBNXxlZl3Zz3fM1TyxJQyfBNjdP23dlZm+Ctd9WrGnuseSWYv7DdsZkV
MY08vq5RRWBRhOOlSx1UpRW83Iur3X/rx6zVwmG8MUjt92Ehzq7+qzKv22Ef+N+4Ck866a2QrLRe
3BmMfruq622oqJlNjswpQp+P6cT78DWFSeKZiz4QecWkERMOaiQ9Y7u/shG9sfcoS90BRyzs3Jtf
70YZ91TdUJFq+G6OIdHes3YnXzgJr87bcx5u5BxKde5uRr3K0aKZfCzgTyJvne1lcfSmau4lpYKQ
9nS6xzQJCLzQWdgMoWIByrS5wFkNlJLD5UmyXrcw2M96NT2K3n6HBPUKpvbJSsAsRpA70PmqDFmU
VTYkvAst6DKTkn8gAwDnfgNq/cEkBk0BvaM8lzKzgZAefRNK32o3Ib0yfRIdRJHzvdzrgfUirYVR
skdWblJ1mxZIjJPy61M4zo69VO7CIp3S3NG8bWcmVgo1j0usZL+pSL2OoU4GPf6vbS4H562msf54
glCi0+pTdwjnbGose71xbayA/Ad5219fuQVjg37uSTMw9Tv0jQbrTXeDz5vrV/oqS6zEg0JCm1+b
C1kEGhTJ59wu1qixdIct1uNOx/itmMzc45ISen2AUhIqQ5z+ATKO24f0jwnpxkNxHIB/Tw7uflVq
qqz6bpy2o7DkpeYY5tyxyxCd7Ecp5y1TS3KQ+GUMoaimpZmn+rpWTJU53YrfEFOnRw5GHsecTm85
YuTbnnU4COAVxoDPSRZ3063jUYYoUFniw/H8zCDagXki/mynVZwV33TTqTO7dqHBBH5ujnBgyu8n
897x1xBkYa4VSJi7KyGyJwQZJNToxaGthDTWBYu1ZH0HfxF7YoQ8upyoI7GbXC5oiqx4PRghF8+b
DsVHXn8/Bul4kQHbhZDQ7ZjnJdbiWfQhRO1W6Y2ugSLOqwBNnjkBS2hqL1J3brf9J+N6xtT1JJSx
tNudc7SXg3qafPVf6xjmZNvicmklGnhvZFDAYDahyeXddmNBu6Aw8rwEhwy298U3el+BKtCIfkf/
OY+5iRjwbVkghxu6y5xarj/xY4spKBe2lggk6m4Kv5AzbUxc/VkbWEHw/nC8twmql2z3+pZXqc2P
5qc15j5UAhqdXZmYKCEC7GlXyMHdG9sUTHnIGS7YVyZGnguhljVIY3TtJfuwQVSLlD9eRCfbt6gH
/s7a9VZTBGhHSzCrvA3Sc3W4wBY8PxWUVff3XkOW7fjXHMDresQKsPjzmCdV+SjYPWxEHjhay8dY
3lGTLVyG7ztBBC3pzQPnWK1TYN0gSJTE6VGdleNRlakD2b4lCJKJGL3cP8WSkINF+j+Gf4Zf6UvI
ghpjR9DCVU6tVVvhtitCruhHmmQLdmraKQocjVamSlqDHVqtSttXE+puW2F6q39gqB9posFOst8u
ZU77dNIiQ9JNYs7eyBkLr6/epuAglhp+VuzzF1T1SGk70t5/W7RsjXcM0HE2gCz2laeHoPh2rGXf
H8MF8PsF36UC2+5lKga/w3IOebT59xF1c5oH/jKCqIyrv6RHHOAYOMF1hSkUWEVUZ4z1+O+LswHS
3uzWe+lqm96UNL866h0UtkPgBiQsYYyEMyzeVe1dHD7Nn/3G3xE/CObfZisWQrKpZnp+QVAayaDp
BBt7sgl2wn4cq68sOlHyVCGnraU4ehSpPDoNxRERLkhandwHSOF6O43dZJ3i+jD639ydWxpTjZzI
VWexlVK99rnSdFIbUcsLcGPnCd2bWkAM3Qco5MCTppQe452EtNaTP3sIrMZP7pCw7+WK/1INZNYq
/SP/Y2fJ9JzwcAp+EIuJqiCPPZiyeqXPtzurgUYky2EtgIUYNOmdLZtblqwqeUzUxYqeP7hoSLVs
/jUjXiEVVG+LDX8Y48Gbl321T/04g676LPMvryFrGilyYxteYJPmwRbWiZlmIFdXyho5UQPrHCg/
rLnaPpj1XHDK4ZvWwwHp2Yzeo/t1qPw3e8QkhffEU//LK8JlI253Xv4ZoEopIh/NDW5WOMngxuiF
EgWDccCc8y13loofwTC0puvhJqDQkeCdoyCW0ut5FHX+8u/3CBvr3m4gSeSNVRldXDwU41iYxrzw
z8HbBLaKKOu77DeoRxKdRMJWiV4cac+7aXWDWXGmWHxS0xO/4v9xv5GtqA50glZ6dQ5ywFIbKep8
QWBSw44cDR6AqL0ld0ooRXfO4C/cfXsRA1idKIlyPRQVM0Q4ivWymIPd4VGCcua6PW4wef+Gml1B
UXCeJop6qa8oq9NLcyAPho1kMzVrhhIxMVcBqMua7DB2IJi7roBUa1BUaw0r0BzapdqrN0VBQpe8
euaNAeQMXhe0WXfb211kL4IdiGV/DFP4zWz1dKTep7FGF+3K3/HZOSpxDkljLHkpAzFoF2X8dcAh
qE9BOdbSlMIynupuzH9ETvC5M1yzkMR260V1dLNSKmxn2iUpdxrm/69/y1KsM23OVky5o6VeE4v0
8ClT4U0LWku+Bqw4nDDDvY+kJhiBuCjHIyyPoXMJl5835dHQtS9rXcw/tm2fVUUWsiDXyH0ifg5g
DjKt2mNk6SOni7Ey86DivNLIje+DAZYeqWQTQvcdNT5dIUZ2CbhWsb8WMXgN236SSs64UX7fqXqV
vB8+ka+wRpYP0NkJ1MZZfgfM1SRxMewZeZ0MGQGMGkE9gBI2mLK8aGLvMUDgMgn81MfTu2YRyjXh
eP401hR5T8xuSXqchgux4J6fzVLPq0Z0phmV806gjLUWRsMMR5m5eYsWnwO/A8UAjwkXPs3buV/M
F2BbBZr1FdbzkYxShLf9yJ0PdVfiyxed0+vz3q+l9AGcYCcngk7cjW3y76V64vC4n+Bqy4wh/xAL
A8RO1B16ghCLBPAYBK439emLQZ2tkHDbooGjMABwCtZaC4zpanOYUOKO9NI9DfEF7Q3WZuljkK4M
Vvic+E+UUFJJQ3Nkh/+pAb4LPMeCPpFuQbCPjN2XTY+DwDFHoiEQhiq57crV0An5rZuGJsz98RvR
pQbWsduIuv7OOpqUEb2IxXw1fSGGYtyOJenFQXz5gEcMcOafhsMMaWf0CFmmtIO0NtyhOKDv8m1a
mCag7T9AAvqybqSZ7IlAHIKn+bn+LLsF4AU0h6Z9aM2mQowULztBHKnasCXNW3k+Y1MFOvmEmWHb
jiPUm5wNDkUctLaeA69DFSoBySPfVXc1o6eO9Ua8o4+pkyw/iQ4eFUvBbtvb/pSWTwqW+M1WZSee
v0bB907Xc+nGinL4KYtluf46ZKJiuhYVNN4VKcOBSzpFYkoHzNw4gazzIjpYoX8ahfncI+/7taSt
fi7anAfkHYVOVXD/vBGbRA4Qq/S2QrTK77HNMaJHyMeWVGM9mdQrbrmY9RVsed3qxjq8VjceN/4v
G+krFmkaER0NOyTva1Q/4wgRuZ43jC9ItT/GlnMc/HLr7jDJcgu6uwZRcSXMOkm3WSGQIttFNIF5
YFSmQSLIL0e7PTTB8Bnkqm8hS+CtEbHf/xIohu6ewW89majStqrCeKFNtkBOrhRMrvy+AzP7BfsW
F8kDnpO6e+XTtZAQGL3grUtUjmIBbLrSIsKq6Sd82JyGav4XPptjTAcushLqF+4grefp9VCaBR+I
EMQ5qBY2GJ992wx2A42cue2Z6i2wnrrYOq6I3QrRROtdLLpxRyqCxBCJuqZFqOh0001y1rDzTLrT
WQFNGeZq/b664mafxaRANNJ6Z8+vSDtqQSRD7lp1WDwqI7QApxLtg+BvKQ3MLCylnG7dn9qKTRjt
ZN5JUZPSGZ7q6p2ApXwTWVGkX/0iNSdEOJbRw70+WPqGHelIq1x5FAy9AbU3P2oLWMIqNf3x/B9R
h9pF5HxIXQVaJsjvw/VZ2zDdFEWLfKhj1FYJjnu4n+3oFX0lAIx453Gnwebwio1jq2RfQsNRgmK6
vWFwDOC5zZC4BrQ7bf4fVNgqhX5cBipheri0AzBKKpeizeMJdtizvlxBN3dWMWnMN+Dja3UbAto5
pcc7OAfK/ltD+fqAo1PFe+vJTBZS5GA7eBNdhw/2O75a7ImfDYNZfnkaEyOJ9FnEcpbmmZ7TZaRu
WGv3B9TBaU3rJcDAaoUZLDgqM6GmEKCnKPOOe1LgPMSCHqRmmzhvxUMP9Oc6k+RJ6aeNef9DQgtz
0ty/6Pmsu83372hrWhbeI9eX0X/oFFA1bfKZDYM/vbUkPsvfcYd5w0xBmIda5+uzu3NFjIXLY3/m
ojvCiX4s/jnD2xFhIYAev3gqCIF7BsB72wr5Cqw2vFkf7cpK4rEeZXWKxLnlnGwuQzrMPEz/Okqb
eXgIbZcMibslQbejQnZsDxkol8++FIAfhuUvBy1vzXw9IV2RzoGuK1rqTwjMfNHVdYKDB8Zx8K94
Pfw1NOQo85miZ9jKT55eG17grCNbNhe/zbassb0yYz3bv3XhwGP0H2bCPub+P90RFWiEJFMcTl1g
cyKwcnU5o2JDkF0eaFq2P7Sypw9saOOb7ALK4G5K9GQeZIOgNzvWr4mB67sY6ZQdzVHE8VF3ZEih
xw3fUkwGQ2QwAVsqbrIFoF16vSc5u/YRZqL+FNM7mKdfy7f5HbU7BiEMyk7/o010lXB9W41WkRE/
XJPR3DD/wcng3kIYT9Ed48xMlKIAETYT+eAHe6SCKaecip+MbpW3Z05q6mhrvlFls3yEiMVDeFlL
/EgFkHEExkbIYcnWcFXn7en5vFOtQV3MXw6Rcmq4U1m+rPDMhodBe7j6waCYv5XNMiQ+G3t5iH4b
P4CpXUw4vlbYB+w6zzzwjckKOER1GkN4wRDFrFzDqbFbkxjk7ElFGRDPXbWVoP+ZtQSewRr+7Dg+
IHhfH1gnsbsdfSs2MmKiNWo49/WbCyTh8q1f7/5CxKqEOSpnqAhSwKKGqzkQfQSWWBxmj4DmpYOq
9v7RzkI7OK6gHnw+LbsgWq5NRyyNyZcOnP9D56PCgMMHZrAGo43P/+pDVXWGpNpgNlp9PiUmdRJk
rq6HrvIdx/PQ+nyI56CR8b1uFk6P0ym7JpvAoDsQSHqThGwD+UZ30Z2f0tqY61UKSn3muNPbLnpE
nvXzlTxe+uVZulm+IXAxcFcYo615XjP15W62emPaWcFM1mrUK/7ezdhfMZ/nmrTQyd8YtWws3Zxm
TRBodkMGdifsz6IfpR3c6LOyKCeYL5UtR4HmwWaKcPXBg2J5Bp1Kp0kWHRIQOYoAxJr3vEaQ6r4X
AuKtxInu5cUzhK7X+2opn1VSEMDrbBfTotZ8nEiGyQtFpczHB7ojha1LafHLR/jX7LPO2qOCeOCz
TcWILGPXk/Y5kIqO1R2g7NvuH4OBH62G9vd6kF9dmKCADfIQCLn9Vf1inRY2yMp3KsJR0CcWRq9L
YQtBZXIIACULaYWnob66btLJVryvhcIpYH/xAuFj8kwrJj2SxWs7ZvXY0jEoHWgCatvTtEJ9v8fk
HctHqJjguDiBadSxGHd2R5hTWNHQmfa3VtYlMSULltqVlOKVp7buMVQAUkvnek0dEQ8s7LIH0VJU
wJhOSUZAdhOZlUEOg1nyC8nU7qQfkJfHHhiMLjkSi6rQ6yuS6JMCGQNCppsG40Tniy7VDq8sscB4
Khi79fNNKZ9EorK7P+2V2pVzfIKzV7k+SSfZ7fIfkcsfXC5C02Gt+3bIsOOqE5nEYTpFVkyol8+H
V4HJnp+1AbqM01K/vpVKZB8c+czGrJSur07hgzi6pmNH0gqZXtcpWjdkqvwe8+g93IRdiMH5GOHE
p0oa65zCqTDF9352B5EMZrHzVQG75lwCWGqxlUnPxight7QFNpAtFqxsX6B5z+dOPBMYoRcqOf/T
Vv4bWVt0Tal7F0fuV85vlsyHZgX9VD7xedJJC41ifaW8tFqYjaHBPaNliduPRbuTNzSxouN6VpU7
YhWbp6gAlnJsSboHuDvqeGaJI03rFb2qCCU65NWnKTMNfWwryU6g3ArvhxkmedTcKgZzU/eT9v5X
meMO0egVxvlMe0JeFaYzh3T8om9cRGu09OBzyWbOFu6/pzear3eOYKsxf2YLr5qQmj2fZFeShfx7
J/rlK4ELO3sGV5GOsbQPZ8fF538Veb3bUzGD6QZE73Q8jJUhK5XsHp6reL+zQcJK+1LMI6LqgVmX
M/Hj2pIrmhwQ3TUWg1pgRfjD+dnHyFDmT0FoGH+xwiO0NKVM0HP1LrsjYgWFTHcSVnJzIu+zqdGP
Rf5SFeAWyoUUGQ6yKuidK0I9CbESnkOT/nxe/EeiLb7Z75Vv+nDn7+YQvmQdzP4b47kLexYdGOvN
z4i8LGKTdkG1XYEMAXU5BXnG/BvkcUnmmd9KlqrDtgXikmCRAz7EpvwGJ/2sp3CTCPJTKO60e/H5
rgnJWXbkNEM/R8bEyaAPyiweekJ52g5QHyA5MmZzrHul9Ymjq/1ZzqJ/fzo1PzUzvUFcjuQZ9EmO
GiNsOteOAeNub2VX1/nf3dAmw8bXLJIKDWm+ZD47QeELjqFefHTSspWltwSRgIUz8ol2gcScvVP/
EQd1pmEjkR1Vh04I4OYVhwSRfQcd7sSuYHlyXcVv0L+TVe/LzjDmzjeAA7/dkGBKSG1X4WwXyVKV
3GCt3YuEVF8crHSIFX//5RVAPPeGqjaNXEpsGPbsDGRB6hbv8rggTIFAL6HPlh2UM9DkQHYqsF1+
e2x7CulWT4jm8BFHq0MVUY/8dbBJ+YNKzbgbnbs9iaXFvSwUWNnjgmsX5E3InOcPsp8zaJ+Bu6YZ
FTUtqWMW32fnO6yNgWkofvKnGFFjVkEBTmD6fSWPSjZq6N4MjiGrCUKXvEI/XjZ6vKXiC+61Svnc
nsx4yIT02mhD6FowPJ8ehDXljUomAGqTTodxzd0suvR3sEnu2M1UE3hoMEG3MhIFUyEl8nWZ3Dr4
u3tjJoxLkzBRCsGh/Lq8t4/1RAsEBvWI0AwX6v0UE2fcl0EWfZTsidAR3/MfdnopMslwCx68pI4N
Px3TN4MGpYEM/634+IO16Mq4DQw95ghzRfdoJXpQoI5k7zkYSjz/bZTvzQdJXKlVRVmZvanKnrPJ
n/OIAKfoqweS15AT3r4Byd4tLTS8i2qpBwPEYPVG7FvFGEwsu0GK9fX69MeDB224jXUBXSrAupW5
1i1DP3+TyMAP/Aegfc8VeEoffZ1fF5ha1HuE+f+bHPsKWUO+iT6TNHQxIcTtww7E+ZeWR+RsSVcm
LFjjcbK/kIK4RLXXrbxCltPTQc5X+TBDK+KEahEWwG5Xf214OOGBXp+pZ0MImZL5i67vBj50ROyF
ePuScA0eJUR9Z7CVwfW3idZToi2FiLPJ13ii4wKOV8vresPe6Nk3hWa2qbwW2kLnXmj0KYizGdJd
5RbCpUCrGXVKhcZ8fw0ThHZPk4jtjWKWGFWakEDR130gMOukS+JROeOeDn+WFPF6+vlTrdwUuN4B
kXfvN8mOPi4vaQNxrmjFBa+ZoflCxHfviOv+T2KmV76amJQlvmUW8yX2oZbH/QiJpKzYOjdvhMPo
AjcqQotwrSyn9FpPtgybaaGt2HLP1dwj7xhHYpT4pPNxQCiHHaSuqB1PwEsVE9z6a07s2xuaBui0
Hfab/d2DxXTjMyk2K4EYeOh0HwLyZttJ04TclRk9q3fCnF1VLhRkZvMusRu5BMwTP26TmaEUePhF
DQNQuRdh1XtFKc7p6XLWZE3YFzwZgIV7X+wyr6QpUoroOkMPeyLcTZyydtpKRhhUU1QAK2d++GkT
Fdj9hTyM22+QKZVe2Xl5xvGR0/yqBE6PVufZsgII5O+MbPyvETzKvGvOFjVh9jcE7XM/kHPbRdJZ
71ky6JaNBhK/OhQnBi0KkcVNACqV2j53PfgB28nlq4FhQ/wSCNCX5K93Q6Z3VDwuwUMaUNDiFOKo
9oeHDDtwo5g+pydFxOHYcEG3w7z1Q9EGq8cL+rOfOAp1K8DivWMlE/sIWbV+iT/Dcok+3lY5XQ7Z
6Ar6t+MRb54ehFQRh8fW04aSpsJ3rfjYH+NNA/9f1tYbNdu4++df2Orj6jBBQPuo81sTxZdnIw/a
pAwNMmFkaylycWeVGg470Yp7apuambX0CH2tVCtp+3rgvA+WUCk5Q19oJ4ixCZqohEx6iSTFCms9
GXrf06dOS8FdAgAEnDtYWAOR09/f0IHqmeQxlBoOL7N+gWoU2yPqvNKc3Wt1YiFbCdUg74Y+r71v
zL7annjucBT25v2Uj9BbEEyO5tFsE2sjI9RxjvXelo31HrbdCHAKbQ/4I3vqXAO1s8xaVonvn7Uz
4GbO8R6+RQMT9sVnZh1E9h1x27SEPVwPfw3/sT2pOzj+wf60oPMECuJRm2clgG2qg5gMlCAGvbrd
92Q+8B7GgrVx0UGLnA1DNKg0CskRkaUPBwfuBetEuT6HmiBahaNCnOHQAESeWsEEVmhEz+UBpQom
vZW9cY27xX/oxsvsh0gRmm6ObDqXBshPK5m1bYlmsnkJO4gJJNdA5CmPO/O3ezP+cIrZL/ja0PVW
Iw98AxvY3mDPZ+gNj9dAKObSYHYJiWvQ2g5C8Uob4oVwkhZlTWrTPgZmkkSeC9jSz9x01xR9WBxF
OJYn4b+SJqepDuNBDsQdeihaoxoTD4bowg/ewxsu4EXj8MaXXn/esi/D/v/ZEHp+XCq/BjGp8MXH
SD8fuojF6WWnoFCGlUpj7iff9trgWeNQp9fYojElflKNUVZRrRS/25ZWLzT8Z88oRy1w3HS8qQb+
yWQpJpxmdy5/J9r8QsuguS4mfCyM5mFW6Zut1mFalSxKYwXaCKwYNjL6Ye8pmlYm/KEKWeDxpWW7
Y6JyJsAbFR9vpQ9aQ1hj7Z++gJTo+q+6LKu1ZlTBPT1kNIVxwukNQuPxJr1a6MaWtpZJ9Q80Cawg
QUuGKJKpp7++fyGiwqcXLFywFG90BXtMZsg5FOWf4Z6AiubI2MHXoMaQlxHVjEkhXLJ6qJfcbn4w
TgnywPgcy9qBDO5wbCgjdOxY/Hqa1U9bSlvEKCIzuIHVwDeyn/a9sc8RZE0tzxrR3iXN5ZcMUHaz
TJN4ZryPDv9AHut7Vxx0ieKwKEhyYc4ptIKkh7iYiWmKViRNPseVtjWt16GJtuZeAER2V8xz8h9f
57gxIjfCYt6Ef6fK+26BSd5QPKWZtpRv8lqXiuarrH7cRtetcWELjmUtyEQQz/kg96Crx3z7xCtv
pl4Lf049z9RwHYT9gD0PE1YnYl7MBelLFUVIkllzEZqYDowCnL7sM58Kgcnp6D08M6igWe/4M4/G
W83dLbAMPwbGd5zwaNt/FjVDUD/7aPJfP8+Dfhu6fALcPTNf76juyVpAavqikqyCMW8wvtCWy+NC
81q/Z0UGzesRrdUg5LBXpVvE7GFeZGmW9jb/VnxItdwk6vMXYTkc8DI5iWzRD4H8OZENzr1Y4tmg
YTI/dmsaNYQDt+NSqF/1u1sPb+mzl+ou7OGsu9gMgU7hjVVI895i1oagi6ojGceYFwW3YZEzE6gc
p6Gi2SpAMsFotXXODXCYyGc/G9OvGamqm65EmfxURbI3nMEK92UE5VzpJyibUm3T6x8enax4lvxT
Nn655USTE2e3gj9xvIGKXjIDFS6gPBZ1asxpbM5t2jnB+h8UK1hSEPBTpo6vcujgmbP7D5VlmwVe
lPszzqZdmHdFe4Y+8+2Rb1mCiUDJ7s2rH1U4Tdof5okbS/js6Xi8MJmKGnh0zB15fzcqvNni4uZu
1JYA1QLSRBBYheuYSLHWauCJMqFogJfw0z5QeY1wi6na+hE9TwYY2WbbFv8D/Cr62wIod8wc+53Q
oEH3X5sae604Nwjc5XwjmIrSP7+fff3jad2EVBJCjIoI04ZAShI72hqrRcJ/cPqXZ2uksTKnQkrJ
X+VkmZCk2FfrBao34yD2PTQIO3WBW8ror4B7cUJ1Jre2eEdYESegTkfnucaRZIibkeSph+TqZIe3
jlyCEk90CcUj4zbiN8k0ekNacyR+0n8mIRzeZS0ec9W78ruUZRF/nSO4rEpDFwGwSOKX28SW7Kls
8bogT7+i/Tu5PFnIQ+3XLcao7CGP4Ckw4vHER9i4tiIWc+0z9NiR0R72lRKcJos3+5YyNpnYnw/9
EL2jkdTh5/AoAhpghNLY30+Z0ezVe+BXCqD6F1TD24Z/NxlN6LjtoopM3cuzFEJthmdcc4xICh//
+31ay/RRHjjGN2BFDj90+tfJrZvHc4urT6tOLcxByf1sewASsMw+SZoPzxKVgpMpx8Q7GaxF4yq0
ijFI3Fel74Ddvv/b/itTm6Gkzs7u1b0pi+VR4tRSSqYRhiqGHzkk2HyT+cl6sW8H+WvgyxiESiht
krB8OYXrgSt0vQU7KvIdN2kbuC3V3bD6uL5p3IQn/O9gUvWgEvUb1hpquBsXlkqGEVyJw69cX5dg
O+8oiiM/KXN0RXAMyUb3a1/KoIBrB/oSR4bG7NXSnej5wJD6wGujrMon5V5BIVWrj+rqPNpY0clW
KjdJJg1dfIJiEfVEKGbcLjIxwbezd5DBP3sFZhhir8tHfr4flNwVAHtfsuvADNUtjHDO0yy/0rC2
DHBupcfN8lyotvtof/UHN6BHJqVhCN5OZPcXYmUsSnBT8oePSYNLACvuMQOuHAYx9OxULa065irY
5gBZGg+1mr8AM8ZRfzGY4rhIhT6neyezHQsKyEPGkwUWvaP28S+YkqstHR2UXg6WMRXKRpB+tIoB
ekT5x6eAnrOu2wFDVw0GP6kmpCtkZJxT0pBLH4La1He+BXsZOumt+bur8IXfcdgcbWeKN4KZgaQQ
6Qf2LQEvmAF7vDLozpBOLzKpTdu35Y1NWTY6gsuDJL1UHZMk6XIQlzP0tBJIRtNN+s9pWBtrLjta
RgOe63O1G/erMafcnLvmBxK5RFOpYT8KYP+ZuD6SpReo8DY/SI50sa54vFmCGBzRIeVclAO6F4PU
2bXMfcgxU/n6GviSSeWI1Fn2pi+MBODyuUiuTM7mcfckNdWA4Ke1Wx2EkByxAr0b2OacmA+A0UBI
L9HldBRREwDJBGfLPD2MsueDiw6wHW9lOkWq3rMKVC6JoAdUt8yHbjfMn12T/Amk2moOaB1bqm45
TlgpCdTvyMPjQUcDcLE57/rSuB2tIg5NPiW+Vcvdzjceje/AVdiUl9PyDxRMdcDKEJK2V0BpfpDO
GVSswNkjBimNQ1EFrLcCHXeQm5Ns6GERwLmPlNI9TiXVfjQiY+lqQJY1Zrra214wGZvtaB5V7xuG
wcbSFvUk6KsrrtOm8B90Zw3p5Po1E6vjSqOxfQHrzlOIPJekaO94WfXPtj723Cc62Cd8TR/li89x
rE6KcQoRR6C3siZp/XielVG07xm+vj0ZYaXx0cis7ScZpddcyV4q4GUU2pCpvDKxf7okhMCwmjFc
UY7z1lYyIGeIHZww2zlbQRTj57zrkafSqa5JmM6YNThUGg96gxwXZWijGVCltanQdOIL32+v+7lG
rN7C9uBoUcuuZPeWHwWV0gWQXsJR/bCxc0vjz/AEAirk40gTbQ/Ymuq87FuQKV0SOKZsCeRDB1qi
LpipKbPqmC9U7HVdBBrdqkVR8l6d+aMhJDk13tlENYxmQ1cTd2I/kI4V+Gh+wILsDkDLlbfQZcbT
1mQH09O5yJcFtSE58BU954QHR6angDr9F5K3Ijr5da6QjKs0YReFQgTTMBcsnKLR4vey5W8ipSxQ
cy+EupNfc+WVTE5qZwSGOb+gCIMvGbAFjjKN3YPxGRd4CIsTHqFu1QeF08zN63O2IrW0Z/MHyVO8
LLbxhq+FX+6MGmRx4HQdQ5FlogWAi9bHLtaDyIeuVpmo5PZ0ruf1S14R3+xFuTwRzym2RJnfNKsr
gqwNCfJEXf4vXqxXlG3eY9gB3lSw0Rn1g9O21YguLhQ05ikz/qQhc9Nu/j/4uxJMsGlDDP9SIefj
xSoFS4DjxsF5uLQTqqgX2eiQwucnRVxBBrethgCrTDlhckxWBq1Tm9c3+VxV0CDF3m25dXisHC2R
cJ8nn8M64MQm+hmnYWh5VjaMHWOBHEc2LGIshGt8rVBPIFUMZNbRClH5yRPKHRZ0KdqwIcC/VztX
N6prM+f4TYggCgF7Ipy+oflM+n8kIuOX63Wdkm3RqJN7sArCGfFEm6OCM8UeMbWt/JSxI5YlArjK
dOcu0Oy5PVNyamfPYRiIHsEd6uVgqDx6xoef0VDHlQyniYQrctSp2QzXKSkN+gwgdHUYFws6ApVY
NQx6VHqxHEJdiOgebKO1+hQ/WLyorkliYuYfyyBgVkZMJYo796M+b09mPt+inYYVnLBiHrNQMIJ+
YdfS97dLcCsqBHOLPaxkPTKd1+5/E1ckNEQ1BgSySiupQy4D7jBjSfyWrUxo0lu+BfcsO36CiUUl
HJc5ULeMNbOarnTVh3NsMJbfHoIIVQmWUYlRLVq+E7wTv5rUmOOaYzwj4PfwTSRHQrTdghPZcoVD
Xvul4vPFIr22JSzpBmgzLeqjSlDtKamuc9KioxH/hB//R1R9QnHL61B0JLe5tiw7qPHTGWke8+ip
SunsnLhoVz1qw2r+tdi3uhSTB1MiACNu35xtHm0XjNedG345IJDxKN7LkzsVzZxwceqm4lESmsIR
FozT3YR5XxP73Kfow4B3A4JK05PhjusYMNcKK0xIoyNCUDlStUdk3QJMbG5KebsiDwjE+O0QH/0f
sB3LSnIjevPouHZnxYhXEGYMZ/LjuALeQSA4P1PoXLbvkdOVwlDg17OZC2YfI5/QS4EMAgSO6qSW
42XY8V/lRJcPIF11/D99IN3HX+FMAkgATMPLPX4lwh32qQ0BNP4szpf+AeoVJCQpbKq/SqFf84aq
lXuN5yUwESGeM2hNnKDqVE+m2CK84M+4AiuNUTts2dzPi2nzyrtEtQ6999Vs/nqGM8nZt5xTURMx
l7I28bk70FW1z9llUGJCBtdcrCwy+yZncvd736GnakEciFg0uuxkVsw9dE7Zn86di9gCJIuJyi0j
btllofKgTNsI9FqVVRG/qqdZeN2nH/KulyyCqD8s12QrrUEnr7E9YAgR3ki9jIaV0Nu6N+ukb1j2
pSIfv7hlzYbLLJcQVbuiNPTJBhgHbIvQzWwfsTu45Fke2Otlk/ivrlESs7M7oQkw14BfllhzNbmS
hlvPskzSjR6S32K/eQIVUzA4JN4MLHzVPurDOgV/OV2UWGHnPrHblHUYw2jiY4F7e19yzYlC0wg/
kJYtIckEzTQwoEIaTztT2iFO35XvffDQZDHDDHtMuoGRwjMyE6RUBJqh4RsFlY76qRnUA0gBiRq1
8RJMuZLjzCm3+Deuf/F27U10lt/yOnhAtSDynHdLeWCnXtfOqylJi2h9cT7HvNgCHpdri+SsHMr2
+9s1LrPrg6mkMt1yQejhpHzOodf8Lr/y0rb2e0QbCIy8NfC3rTc6ZbYgUcsovEiHAYgJnUxKyAQ+
RnRAg8f8j5BKYD8IrmhffoBUndn9ieZJ8LmOAzBzlL2GHapLbPKy9M1kPoH3m9bo67VUJVyBBxbN
DQCafo9+DIl6zCJUHmXEmLaOhe96xIpF6ftYniKPRy++x9+JUHZEHmWvSSC4S8ic6LRUwq+KDvzW
CxDk3c7qsG1mNJCuvhM+QHrj1uXdszISYaRWh7TAgcoNY4kQJEy6agZrUOR279Ge74ute6BOileY
ZgqYhilG1QShRGoolFijicajdTlqrlidTv9ZXFFLD0THIbfiRu7jfOdywc2QtGfx0AHGGPysNO6I
SRF0/tHjUiNYggN02rJMEX6k2WCIEQa1SVs63I8hgNLmnBI5GHUpihzm3LTnFYsL2zbk3CbmLtD/
qkv960VQAZX+NQHiRxSlIBgCFQzFYx02EIn4+T2CnLCCeHBw3gXF1RaDqEYJH7IYIyhFBm0BteZa
9lmGO1v1Wl5lc3cYItcXtYIRWcYMjqF8m5R1jh1FXxYWQkzspNl/DbkM8fhwPl30vah9uQoh3h3S
leBxciOVZ+vuQpGOGyVrl5BXqu68YxNu3iCz8/21od5QScuZF/uPjmzX7szudnYt06mCfJnZupvz
qYhD+WXfGwGIpCKhDOFRCV9OArJaSMtp7W7yrMy+m087Ez/yKslxpaCsVuz1HNzEvmrgnapD9n7b
NZxht9/3Twi+DKZswxAfEthFtDzZLJbk0Ptuhgmr+gJFSL/H6EBoX9ImOaAwtZyXYu9MCrGr+eft
/xyR7eQB7x2WJd6sAHs1FLvteFS+F18ZL7hcnJBFBRm/GaR9MH3sItJ3zSGqUKk9Eb47nBT7VZg2
aiB+6QP0RgrHiBCMPKTXVxGjpBSw7fze9wekme8Ug2wpuQMeXPiLMwYqvhoWgtTT6KhkPYn0KVXM
GZhYkD4T5ECFDlI5X03/+ANAYuweA4g19G0imtKu1ZUE9wjFwoHAO47Mbe0Dgi6tV4kRcDR30mOz
1BseQ0TCb5hnskajPM3V7v2kg2T1N4x0DgYnGgF4rIlPXav4p+EcVRXPw5Q0EARvr7rtJ+MVSIPf
KttsGJ0fK6Frv/fn4/43qJdfxBRh1QRO4bIKuGks+n38UsckNZ7OiPirVF04Uq75NGTGlWU1cTwD
OawdxDfEKEf+uA/vgPJUu+jp+REAk6fKUNZO8c180IEs/DAF4zB3xkZMzVEcnhOfO+p0g+Jo4tHK
V/QaMxias2ZjviiFgwGosQVf/r5osfXZ2Z+ILHyHTgGOnzORlIjhr6sOTUnxVhOdhaaVAD3QK5aH
HWz+5jJX8Sym5ofYcssIsRWFO+cBu3l/cH0tyL0cXCV4NiYG+pCYJOiejpKJ5jr9OATA9PpkvE9f
QezsIlnzKRV6KD25h7gwbSNToOiQ416m2M/940/MYzOqHbYME+HYwzqJDKE9wXCsPlwPV9HkdOhd
uTTmNEGH6LHvO8iMMqM646ex5J3KyOPmHEZDp1a0mGDDimqCRhVf7E8sZeCWRPGgI+9qHc9Kgg68
GC4jnPV/S29JXmTYMxku1zHcLWJc2pbHyYYWF3UMkQ/OwGsob+/r8OEiAlv75nSDGPBaFrL/mEIY
rU/F+ey6Lf+7qlphHHXM4G+ZIvp3wcO7k7Q9XGZEEacjyU0I1TgOcG5ybeg2NpTLZ3N/708aDVgN
VB6bK03AV2DbqmHWNksLEKK4In6tXUslugifa6NQ/S5JOdko4auZ2tn0HGVeH1NPHwh5bF1y2oKZ
CghwVDDPWxh6u+0dL5zEkQrLfXKyg6I0/FMIeRB3D/W+nSHP746c89aX4DBT2vF9g9rnxc1NJanU
eesBrBF4yHxITiuDM4Rayh9T5GS3QIJ5+TP5h48NKyl0sF1IZxXvtgCyYyrLXXqMnnpF6RfyWf/Q
e3hzsQy4EHg5NuTjv8B+1ZJoRozWqn8fSN4dtVpdFvVy/pehFTILuZSwc+Fi4X+miHfZU5w5vH1R
x/xVv5WyS3pXvKtzDDviouu+/2aXEOZL7rcmZx0XOU1VlD0QP/xoM4uR4TXR40iLXYgkwyPLAtlV
1JdQue3/HAL4K5UAL4zebtP3xaFNA8sRJDv/jW2zFf6ksZkzv4mVZxzE7FqfV0ncAAXzTl7o6pc6
S+GBTpRY3mFEAX82I8AJ/yRaCWBJy7jQo/u8XBhU0HDZPLYgALES5NNQ7kzXp6etuaQoIw7p87dj
DSLSlmXJMfQ48aeciEDRJif7yYkWfsPFjEuivo1HYP9y4x3A4Ze02+JqnpGDUatctvwdjiVaK25h
qIaYYckpFNGqxDnx+Uazl9pPqYQdNqP/fk4w/vnmknjwMi5yiLIZ5VI/CptcQubu3ABulNCvRuUW
LsdoZaf0SO2q9MN8EI5KvOcIAfWo+rFI6TVz9KyRBuho9jDQ++u1DUHpM3+t2DFMUEsncLDDEqzm
qjQZrqFeiiGgL+isaLHWm9S/bzXSGX+qLxM+lhp950D1vO7Kb0MKK1jd11KtnhMCL+LsdZBJs8L1
fqQQZoh6HXTOJOFRdewIdClutPJjWfdeX1z1tN+0WxaVBtjNLBktqYntxVbYT85n1lwzhxj6+wff
RiEfmgLo3YkHsuuma6UroLMgcei/+Boz8CsE/5GPWIiJapAnGbWrPST1OFWsawhy9g5JRnNGRPaa
a1f8MXzR2LabWQaStt+V6+KgkDQ9oFhG6N67zRwoXUnsxIvtHya6eE+C3xOPhlEZgf3/kydeC8As
68UZ/t+hepZtyEbiVOJdH4d9Vq1HX4Gl3GFxxnCFCw6d/SGdxi5cbGn+NVchIKgnXIMYmr73YRvq
hKOauopaA4JOGdvgE29i18eZNOMJcwkrR7kKLncdind5rBRaobi6PGEyaGLCApdKmlXMY8O7Rykl
SpdsgVrXCSeBjKBWgLDXTNwTFeRWzXZdHbJRvEwXjiwLRPJKiDALWA09QYmrABoGjtMHhe0dMcbH
dCnjsJbDIS3slIs4bUWpJ/CfJdFGP68yF2Y3tPnZhdII4rahjStyV/LwPrHgUYywC9DAxmAMaJ9v
LAry5LBzwQxOMK/z8BR3QeevJbdrd5l6QaqO02AXwcr+2Wr2+FFFFLGTwPtd6+StuFnAOmZVJhPU
eCgo7mdGGhMogHnOZhToLcj/MijozMZs+3buDnpihf0c+F7GfoKFzTGGpyQzDJV6jKintphrXs/7
BfUotDDkkFQI0FayoztL11n+2iG55hPSDOhNi6hduU+HOpZ4xkcsEs+0pUht5ikSUnO4+Ge/smHE
gchubUCYOXQbHdjbE8eAr0vrLfuZVGlKgHEnuMEDpIZxtHNmm3GRMJ67EfPQMkTheKDUKjNdCpAB
IfC9Wb/4AYeco96uUt4qlqXQM4Refnoy/jP1aStWSM8Cz1Ff1m6FnagdMQZDBNvtW8NPusl8ubXW
BdtufyT+nUvKxlUOkOSIZZlBOk6FRxetzOEN/YJq3H0RqhrRR8K/fNpbCLhySDc3ZWdhCZStxkr6
+iS84HU6+NCvLqU9t6bSR10lWMz6EIf4akQXWwLPD6acqr8s4kC5fQCbP2j+ENwCoATteutIwcsr
R9TpQnYt9MMcQpoxWxvZGB+YKNJ76bGilF3IVVseM2fTscxY1P88OCfZwVi6PqyrczFmOF9uO94K
EijLyzqGDwHZPAMjo+TqelsP2pANz3Qtkoo0eks7oDafeleovtoYS1xfJXdXeNUer/L0uygN6tAr
Tfht7ccswLYHUdE7oHCDM1bOKfZ6McTPlw3FS+U510Ew1HYHisla3GIaQuxlE6PEdtMWOKQv0hL5
HOn8ndPFcT0FUNVK69PKDgsqaMjWuC+sfN9UXii/69K4aSJEIE3ZhNl4liCf1sppYiVUPRlB8o3P
Qq2FweF5mxIjETdD2vVz9cbol+I+Bnt/Fc4/M5zCGs7QCyHoLNUUtku+m102B03SWH1Is1p9DE7K
be7BJw+4TSdEp9sQbv3L/IE4JowNfFxPPHMlEoyqFb2W8C9ZqR9P0hAcH/7W8L/Wa8+WYxh4z2Gz
j2XXl86MoKyKBqI5ZR82+SMPQpxS7a1medE/w4ir07dfFELtfZY/cmBPWatM0u/3Hj+9dgS+Ww2B
yxaiaGrsx/MwkoYE6p0cQM9JfhwXU2m9ll6nBu3540j4sgssdzvBsPjcDfWktzHZ9JUeNdfy09AS
bMKGygqDLDokJjtPGNSZ/5lBF54HEoUEKymEKfNA1DmUdJOQdhGrauNV96hdLcdZrUrlfyVeICpG
hL1zs9Gp4alAP6IvM9bPTFX54GJLmScnZMFbJBkjos4B3j7m1K8ihMpdwKm/1zGwonYmYq1Sf/kJ
SPhXE6MBCCsyainPSlH7FQz3miq+4jPSiwkEKbN5ygw9U/Ol4khkLRKUAxWNqixSTrvJL20Fn4vZ
V9/9RWwfomo1C68magZvbxBF4Gx1on+jbEjX5cnll1Nqza0xs5m7Bw7A5k1ppRPTxp9oZSU1R40K
c/Nd5Y60F+cvx79RkshTLNvzr6ptRParWT4tTnq8NzCp6zBroWi+qvsAwVZXvFpeneWiPXfPDlbe
4c8N9RsMzm4n3rIqRHPdnltkhBcqbqYaw34+J3BMci3HcG8XjeAgtyy06vmv0NBASQ5OPMseA6eX
/WBnOdG9GpLHk3/rLLoXG4gYnfZZhOdY6ZnE9DPZareliNNDfvGqeG/H2HNNKmef1lfZqnO1UBIM
YzcgBtYsCqx3YM99jFnVzI1J/LzI+7P7GpVqs6PrfQmTr7Ax/CO0jNTg00OL2qo06G5H7hMEfnxC
iwMVfZ1jqJZBRORm8EZ1hLbRNseVc1H7gzDfuYYNHKJrMh2Ov4+6B2u6WM1fxfGDIePkRMZcCAVj
jRFlj4t+k6z6QfHR67CSMmOMnKij5CW/xwxSoL9Jw3GsSDADRbDaY0rHphFyDsj2FulHW/cn857p
Ng3AcjSk1eNVQcMx30SZhByXqzyDE5dzaUHw+YRZ75Kf5VFjbZCGMyc4HtNp6a+kPM/GOJQ2YviQ
32FZyWc71cj46FVEqCUole+8OiXPDsJlPD+wGnBBt4cqhDX4w3w3fZmyoFxwzFQPQjizR3tmEm5V
gyW822M0UJuxx48PP18wVfSyo9zmRINJOrDyLAvkTPsRtjQpQGVV0vG51DT7KgoYXsJUYuqUDy5G
sOJoP//kEi+rw4PEu2S2tLrreAVwraFOdQITMdkgR6dGuwlHB9GXW+ViZc1JyScHmFdX+m19IMoO
k96Id/tiqcuy5wAPbUUqFC4qCdtLg05wr0cKIuMJhoBF+Ev9rXXv4C+vliyAYMN2Q+SEsyeDEef3
62OfWcCdnRsREHp08j9XGveeODdebwQlIR1TkYsJ8JCKS3mS21KpmrXVnlzqUrBBEsIkcoA4uloc
x7QJGMY5+RY3IzoGVSCteyZLBdJ13hqOK72mc6deHTP7KoQGrTM57r0waeR9AC8q/0PgtJNjCZvy
LWfYDAoqYrZYhmKCZTJCmLRKAZk0VjSRLp2hr/e5olKgkYEVugxm9c7zwvRsfl3KZ6Ae4+7GBdP0
qnzUdXW+DemEoiEB4NVSPtdb5sGwBmxYT5Wp/GgompD+oKpSdxPRm1N/43xW68qeXtT2Aq3d5sgj
4J4CMBod9DZ+KmYQHVxONM2ajFL+e29sQf8ifBoTI/Sv8ZUGqPAGkS3SiZWZ8cwsaPsX6UULKTAd
xMCjbRF8YHhCiW5/S5b5YO+1uKWoLamTqUeB5+CpAUBhnmVXzcnXFmiBPWIDLNHZtkGsJvZW5UT6
f2DNdK+mD+AOSgtt8u1yERq4PDqLMd2rEBI0yNL3P6MRbeR9XxiCEpgM9+po5XhiKv+nFREHqK0Z
TjEUcSzsUwHhvo+M8/+uzBK6kTgQwn31aXgTtRvuD1K7MUd9N6BKi9rWO57DklEFlT29VYaQdICj
MpqcN2dWVSW/H0SFJ9uyx6muFwfDfRktMYRtwLEuMuQtnj/7+4dCtu6jFeBZUsUeCk2HZJAprro5
knHdM7b65Bu8I+qsg8aHo/AMUFXGWIj2otehPApmopPRkmTYi+b6pbqoxnFo3SdPdL7o3J7nP6Lv
BsG/Gu7+WFUc9Q5dHhnIIctA/zkO3L/3oV9hC/C+OU91qZ/KbajEIXmR2godgtkqB+pyn0RX722U
KzeenlbO1DEgZ7fNUSASscz/+JmOkMBV11TWlD+8sSetZlgeMTC3d/NaLO0O4cRnse/pI5NkUFc2
GJSSIjISmVwNh3dIxC34FV7gkEgppgA4xmDpPV/4f+wdHeWmcxVJh9ogGGnUhabOWQnHvzP7gt0V
q+Ty/mMXU1evKnm6l4lzD432i/R6Wq4g2YacCoMs8qGVz5yI6Ab2J94BduVPZ+IaWRMbMJVnmLnF
n+Nq+tVeu6Ks2DsstDsY/Y4pzrI0A7S+J9USv52P2BRqVxa2Dn7cXkq3sl0aUjcIhFtRZqGyb9Ok
RGGWJTN3xfd7C5AAZK81ZRi/X+sNsod4ObgL5z4FRprrJ2ha6QBzcMSB05HwAN0KGU0QBBwMohRm
TEBr1jKgLqAW3kFgBzDMb74TvyafZAL8WjEFjMicwoamNWWSPdQwDslELAFOAT9o2CEvQN4I4HKa
GnkP23UUlOOqhanULV22YYXueLTMdTGeKRXogwYKqxyDiIQdBgkEnx1pxbg0cvzFxVw9aczM2NEz
DxDhsOq/ZUIt76LJUUgK432cC8t2k4kxiuUh7UGJW+bxVrGeZCf3TWJAYXoprW/0P3Ydt5FlIKAL
rJv4WL1yWqXGux1YdxwPOwSVHxwrnP077lu7/JxYGMTxEHB0AmGqlzMAWLOkXD1QM/5baD5HCQ8L
GngTXD8QsgwcCu1bXaxd+665Qn91Ag/TptA7/zDVyh/TSHvtkkZeQ90WJMUnn/Oez6GvLvKaYUKg
Vg2LURxdJOD6vkDdhzeFn8j9/FnP3Gpm04akZ3+ZhxZFVp5JUiVlcQvhQhmlbKBJerGrHcTuDwdk
JRWqubF6RThUqYe5yzzGN66g6abHR1apWcWxu/qyCFVsdEg2r0V6Krw47nZ+gMHVBXihrduAlOew
XkZTwRwi7TmaSLzBl/rhMHfvD75k0gVPiNUQPJ5zyFV35LRD+5Np+76gIFwoF4GvMirV1kgaGGeq
3Icyozyl6XX+6UoBgu38PeX7oF85CKbPWvrXZ/1ROR4x6S5xjMjIK8VkWbuRWwq/ACoUKJM8r340
sYOyCbj3nurXtC+PImmRj4mdcTNmuHQw0i9Vj+b2pbW0akAnwnSGB4uKw5RZNQ0d+npD6J8VF2z5
/QUzNJCVSji7ZKjrIjaP9v2TQOie3zwugB4oH0eLkkLZq0TXYlUlkTHNkelhsj1mapj76I7fpZbi
5nTF2UMLlZOWoSYr2o4C6rILC3+7tYVwdqCvZKVsxpV2plL+pYUqamjM/qhXTSLjCEdvy6Sdkwdi
WopXssvDRxBCQ05E6013BaFrzSt7677E6FzePXuGZeyWesDIp8q8DGtmfF+Tj/+3sGxA9/3TbsOc
RPj4qeZHMuiGYnP/9cvU7K/kIAhmyrjqgVUGBNL71vIF58iShbvxZh70q/LAa937y3E+dEcJMu5c
fRchF5y3mZM/sCRGvPUvgcyCle5Xnw7EnHZBS9ztfoq+hjivmfLngupvWyz/H9BHCbyROL6fBMc0
VMe7U8vnTLO0aCy1gM/q4wJkeyB+jcI0dxFVGSd6bxl+0cQTvn0HjwHQgH6ag1jVImD+HkJPYapL
N33wtXElV2NBJ3itnRFkrAdvfgfS4uQVW85HCIUC73XKMrMvaHbYVRmNG7DxFamtUXI+4EjzXNCl
bc9Wnu98TYn87BN6WRWaIXqeWHKRu5uDJwX2StdxX8nkfI/QaYdLCw6tlO4E4nU0j0aMYgZuyCPi
dda8sqyiaAeAKolx5+14gS6lj/q5eBLiqJXUYiriCBTIQj9pRjkQtsCRCpICSUwSO0uFczLhPtf+
VoTSBdjP2Ipi4G2AX/eJFLYMJAU1SORpuOryAir2+eMHZgnqCiUiavBl4iHMFU+NekWqX9CT9SUt
ehRUORI2YfQCC/zooufoK2xeqcb/NEvhaWOaw8mL61EhO01hxxhrdGWvy/1RxHgx6L5oW9QKWawI
sHrKgMmcdjy/zTHFlkrwmN/5eDOfYg/Y6YAL17mA86Bd/pUlNBZy36qNjZ9EvG2+RFP0zbzgyMMN
5Rq4a2AB1WgvjAnG2liZsVNoZirUCCFvy878UxTWjHclmo8kE42k5ArLRGEnyfftKN/qd6KX0kiz
8As9O7IGohDpC4tjNNqt3m3k2E5WtYiBIokOtRWNslxLH+sSb4/mtCQOBcEUFkKzNXTQtOO9QZHL
M89VFKhr5+fz5pR6zeWJmK9pDrbe7yfpzAQphXwOaOKSFsAuCku3ITym9zO8ZV0H9ftdqyhud50p
1GQTW17pxiye/9W7oOYM7kmJcw5/rxNI565J5aZYVwMz4IdEdaKLDAdwMe+M1slDHFUuNXVxrTiI
iBYxhgd3qPJSsJjxLCGjPoiicH/UHnrVWOWZX7PToxHYEU0YFhVeGWYXx7qTU8G9SqiuqOsdNKmi
oRqvahTY9ikBGcVNl9udZN5NEM+XjBhTXF1BhBeS6t1BGtDTdDbVnTO35h8rmrJYSP6/SoUgnD8T
kI5h7hQ3qStTkx1rBOowuN7MnykMXbtKjfBWpuz/O5evlR7JTCrxas/8M5KL/EinsFy0hOkr15Go
GU201iq394nbVWfwCzv574GbKLoqhUDltI+C78+rwrRUC2rA9r+PQvbKo0jT3r7WeBsRiwilqJP0
4kdLqeq6disOgjcJZHObSG1d51gRWsT6nfs5DNe+tIALVvQXit4Z7sPMvnTJOvAEhQB0dpHS0a//
btBCHGaAuGVCkSZVCdnsY/kBNk+6vhH2dfla7dBHmlvZo9Y2xSnkyVSlWePc9U5TPpev8f47y6kH
kbs5DIYYGo2jOFBZZccJnUszhHjVDDrl8cxdgN6Du0kXLY6GmTZzRLWWI9aJ2igUi/1oMlcfzNO2
isepeUPTtgXaaJytyNcB0lm/6sofpDHuzfT1AFtVPsPNrSHEaomrd+fi4ej1bVJ5zl0QQiwlPoq+
/+/Kj5o0qc+WeqJhNOBsVbwuzT3kE/6czQEs/cBwtwCOU4oO7ERxZBt9ZHOpI7QPySH64MWTQaHn
dHyQd9g8NfWSWRlY6xtay5UcHwcQxCEPmEpWRTgChybInS3ldsiTFengmuwSSpRS/6uCWgipSAZh
YlfVFHhDT9+anIvM2Xg3UNjkTF3pWZ6GprWlpZMBUHV/35wQg8Cd7TpKbIZ8hxSJrYW7F7ac4bXN
muyNi0HaA0+IcmLSHoJ4W5H6r1pXB46mxcW7j+iFlYOCxrZKPDklUSA7vr8VQUT7KZ3pSjcnO4yK
W+cygjDhGsTL6ee5SGkkyJf7/RZalZ9n+YN3/YEfZnByDysPuuI4dhsh6ICZMJe3EyRlDWPeg9uH
sF5lf8ghloK6Ae1ZC2daUoYTSOcUgDCf90q6iKR68xfW0hMUT+E42SgV9qoGJ9e/i1asmDXtgGRZ
VcBsbrgjg3l1appgUknKG2V4FJEj5gGkUWZGzZ6/SBa0iZ99rs3PI9Ael3BcT3XPnxub1poU69Uk
zzhJT+frelFCk+6cLFcw+gMSAdGiDp3QAf9QUiN1yAXOaXuauprbMrJN26z3Zya05clcQnsyqnXd
khfyDD8wrWcqzPPLkJ1FgMVXWkEz3q/tAkJgw2miU9/xogRsnUVg+VY7WAMIZhIyAYW3ZZu+AYnI
iuD7VD6nDXgNMwblzlvZMwK7jFfMy3oWuZPY8C5zgnC3Rf/z44+ZUU0KAHs1ObspDA5lx4RbfRcV
tP9qcryNR+BYlW8/Zm1Cg32YZZS7QUUppq9RgPFYleCWzRai4Pjw8elNHhJFSpbr4GXGQR15NijS
rE7HR+eE70qvBOlhWQRPB1MSEIDVLrNpq2iQ3P5KKL+phEnNaJUlDzT2uz1Gt3WOlaeVzWMdApQZ
5GONyQ/W8eQffasByVSMx5WCjKhw+Bda2IfRxjqsxnPWrRYrlrotwUBBL8rKs80u87nK9mbDGLDN
2PQ50jHRqrrYwBne6o+FjqObbBvfdZF2aBNjupOULAhu7QUg0Z0FbQbcAH5H0cJeBRPWP3h9zTt3
ofq7sWRKUSMhFYj6z78XL8xG0iTd6UyvvN40DrljWwCVm+U6VofdICXm98lTjMbjgECXrDmcC0r4
iMciPKi66MYQrRcgzNzTJX6kBrM3/Q0SBr7DclXjucuzv84zTo51Cc6GQDXURMOrssqrC4UYxE4w
ITlARTWhHiT8+ZUdRSb32hYjipph8E2wmUWDKqF7EQZ6NWuDvPLbX8irNfUJjIoBF01zHNFvR1YV
262nir+2MJiw2xwL5WWMGzg9TriSTwAR+KImrj9J9sXLr3C7BM9zRZfXTeKf9K5i0qvRBpqZNuLS
XR1DCpFyKDxaQlZEbhnTluBfiHlU/PRiNaLDKNoNh504R+kia5RmZr2gn0rgoZuihfe9Gwq0B7Ws
fz/jLHeluAbSKDehzu81Py4CzYxm2QAfcCf4IHEWBXMIoJueYf65bXwCVsz4W3RxWMIB5clNZvrX
Jy2eot32kxlfVbMCxYX2Mlf/2pb//b7d/dKSxhzD3NnuQRJKh2uDeN0JB9yqINLgL4bFZQ9k/1RZ
U4gNpbJEEOS3e6UCeYexPe9RObpfHhtSpqTxCAVBcEKcZ9Pjms76qlcJveWPK0ttTL9LIptXVOuY
p2wa/7OK4YYR+r66m/Fu+L39bt1A9p5Aij84FZ/4sfJVVmifl3frJvvH1+yIugn5FJeiG7M/jpXx
tzI8pc3dKIGaPfVWLex31f5lrDGqZUkEl8LMOPsNJvhDs6Gk46kMdRzAkYD+EGyo+rAbXWVSnS5q
ZwnFQVoeMnIPVOO4uF/OMT/u3RNZz8HhKckpw6UuOt/1HSBvIkq3/t6EWb5GslV0IDSRVJr3NlXo
XRDGfMJCnYgpQhKUyrDvKcEbKCd9ASrFeLjLSRUlvC1H0DfXJ8K8LSsDM3uu3T2RzHIrNph1gd+T
2L0Hd6qkD751aWGmc6XRNnNtSs8ovOjhWqy77wcPjtxpXXHPOxsF8IJBzl9OysmHtoWcIpgC5aw1
ZQha+XwRQ7bskmOqLhSfrbWFFaQ5B1U76pYthwgZ4NLwAbPZ2foFMuvepp6k+nwoplyd9vTvVjWd
7BmPgQgYitUIiY/v6oe1rqrgT42RPEZp+kgeHXUmwjsU96pcjOjywE0z61MrJ6+iV0nAJSFnaj02
yBnaifHGz7BhUA1ZoaaWRUy07bhS0J25gR6xxXYG6ACHXw+W3Bx65JOQ0s0IDD+VrpnKJbVchuUE
3/GdRjW5AhOIkXZ3peskYPNahYxIga4jwB2jtSUzxnlTT7gpD4dTisapB4GpkoCV163vqMcEKQUN
DUFwLWL5c+rHIm+kELIEUHBF/9tOnSFds8XJAawWMQvbZn38sQ4EPD48KIOknhlK82myUZmWhlbd
99OvieeqLgeIcglNZQXX0RnA0g+F91x88bCYHQO41gfrBBEmntF6KG6jBc+wIuDSHy/0HhKsdxu5
orUwI99igmXWBos8/y+0ySsvIaFqXTm+sXG5jAX8HDgl1+o2ijFt6ZFhOER5O9cGQBDbarzTxFsR
DAqsyByDMTwkuo4/6T+uzRcEbiwq/MHOUNQQFOQp97l3rx/5eawd85M7UlJohRSN4QGWTkHsWQQM
130lexdBj9+MiTzjjLjdwSwXDd2TCMLba9uraPWdeqVM+UeL/m6XQhihLGsZ9wFA/etOwx+J3aeV
OkDZ81YExuf5FAis++6xBwlpYhSiIJHFo2DQZaGU2AwVgOfKbj94W3u6sJY2OZ5trC529b/fwSs1
Q/wvtM4gXv+sPXAAY8aDYzg/Gvjt81xtjGA1jOpVww2N4+XhjHkXSJBcjna9CSaTFWOi9TOgR83r
KcjZ7ldyDyX0cmPesD0vpjCCaq2p6HbVRiBWC5vy06OJHwrgIZ3HvVyr/TJzmTD6HeWyB0NykoIe
wbpUG9w/6axR4n2x4M4QL2LzbHcKmx9R+juDp0hBlE0HiGqNtST2xooFrO1vHcepoNfl7YHpq61j
XGYjH7+07k71WzR7RBpApAI2FpAbq91xpwtNiCEXgOIp7epqbi+r9kzyjdd46lrEJafHJubCEYyt
r4WslkmjyB19DBoJUbos8xnTCBciJufK6KEFIQaduHrhr2K22vS66jgfLu46PRzIu+hdLr5j0rTs
wXSAtzC2L0TXYTwJjAAHtYxHmAAB+sQaabILrXpA5pgAAfneNGrBS4dy8ZX3NIwuaQ3BuJc2SKpI
m+A8xbjOPN1G5OZOSqLbWSKjwJDO0Aq0xOuclUe8XwRil20iIgKiB9dot6Hs4fRbUFbKwi5P7fKT
7ieIc8Euzzg7T3nuryPgzVSPNP/RdXGpm0tv91dizYK50RAO55BT+9tMuTNfL8QpC/RtrrwcHvCr
RKz1kgtC5eEZmRIni4jEa3Z74Kewpnf7pJYf3ndv4OKAMvT/asdPMJKtcr+tqTuqYi94CfC+tPRX
ollcm2wF8d0Cq0w7XI/g+28XRTpmPZuhk6vPje3R5l5ifA7WOdQZvDN4eFZmGyaQD77mRWFo+Vqs
Y4C/aG0GB+L9SMBhUxdw5/VQ1sb7L+e3z5cJPZ38Ig+7SSpd53lumPPqcAj2fRhrKeWixoNwsY+a
WbDcoMUYyT/Rh4kksvfIdbpZ/bseavulvIkPi+X4CEyOHPsTUuKJVABiplFRwm84Ygux4MbxHPmo
nP5XtO322PHdYmFo15mcULN78odyRj53VcM+IfpNwalvp6aOiMfNQBH9IRi2zEm8xRv8+l5HhWwv
Ux8deJYh9ZGXfZkkD79WtduvWCGuTMKZ9DeGTXyPzoNDo+Mu3ngetHbX5e4/8bWXX8l/QV5Vzkrq
iQfuktWhl4p57p1DOKmfXbTUjw3nE9fFW1wq6KDSMBYc4Rp+/dKRlOYnasv3tmr8VjfVdkIDMH1Q
VEeAK/jD0DUZx3inI6A5lk3z1k0YJwJpg2vxtqKR4ZOjU28hrN4mbKp0zhFPQRT55lGgJhNakWx4
H1cb8f1z1UFgMptG9A88WgblQArLUlj/V38UndfkAunAXBkY9ew56o9jHRlJYrE0Z1MvREfb6xSi
0uOmgos2dI11kVENUrhSlTf+qK4RVlypa63fek4POdG3tYQkmwTsF8OiiyQdnxoirBZqzhB/39LV
IYqwAwAhBjFV3cypBLQtYvPRnG3T5Ku3nF9bEQc++7t+M10/wEpS9E4L/o5/dKrgHu+2GKlFpqnA
htv/F60KFxCnKPtfvIBYugQmZPTfF+m1jgU3kiALzDqS3IwTmJrSBolDlk1qNnv4s0lEvGL9qtqr
mGp6/m+/KiB3DbhMSg/EysSARgf6s8f1TWee8zxk+dTkIm2y9FuGMEQ/Wk95S57/sN9cTxxDAcI8
GkyHOhbpvyI/EZuRiOV0O49BFlempvKOuALXvyb4JnI8MxQs56+k5DvUhyGkq1++XA/iN3iJeKWm
GDs+89aGkCDCaRFz8nsTOiwGKJ+eIM26aiz+8D1a1LjAfqLhRCGqBFebC1nSZ89OcKWuViv2aULN
q/yIlMEymk+KMQ2ZW0k66bwVeRm2Y14FLPyFp0a+RpETac7HV30ULxklvEBfu1JKLLImDfwtpbdH
koohqqveDSrAc3LDbMAq2h2c93amnBTU9hZQrmW7dCZ99a7VKyIuQpcCitdRez/KnOBVPrORTsBo
vd2Qte/aI2jJo+RgXHZXJDZT9EUUtoQjLYI2WPK94vdjhWj9XoGYA7gfkHOPtuCbusIucNryXBcv
H3fqRXDO3iAZ53/lT9t0ELbwLDXUS7B0XzqkgolEDAqp9QUJW7IPJVJYT4pNErYg8eEWWshcf3BR
nVb94IYpAnjjSMIVKMYNLK31XZLomDitrnY4ok1VNr/HpvbghpMSNuTxpuptrZqqmYF3o7IXILSy
v2D8yaGoHN7DL/B7rAgOavDElw9vuk9n7b+93tAyLaFrLZP1DPBUxk/OaX0XJsqU9OeB/BoqPnYg
bi8q1yQFRMej15EPY0AiTKihBfETvVLRCiHXGa3a1u8MGpBUR7z3rTcXPExpSzUP4Jnoin7KF6UX
x9ybus3ADbacDHY5rfHjLeC+l9BABgWUxPpwWxKRBs/GuLpznE3eCCi5HYHvrRn7Ji3sNCOJNgtJ
zFCcpLZrQVe7umCRUvzRKeNFXc7dcWsHaZKbMQ+s8K/a0s1EaFSMRq1yW7GazSZwmNT22Fg+3S6f
NCfJromrfOy+Spw/YlicsPmRdgNWd56oOc6uLob1r2GObTnShCSDRUzDq27jkdIFQKeDdW8ecrfc
6YIc/y1nc2I+Shw+keWfE3uS3Ftb8ACcsr8YZWgHsh4tQEywxbtj07h3jios8vV9huyJSk87mJHT
b4fLuOfCi7FYCpds1vSBG9D33FXxIZM6Ky+Gm4gGml/E8coRGlDnXROPSam2ZFaVZVLlSQNHsyb7
2fSHWMA9aoYFIojACLOCWwJcZoOClvDZHfkRMABV/fJMnnn33/mRSqB4kqxIne6lKY6t5WLK5MoF
X5t989CYiL1LU/7nP/ibJnVz3z1bsSPmWxw8YqSaGltrWTW6yw9Ia2BKQviTa03VKch8UTVK8519
dS13SQzpn5FhKp+8rbhBGH6rMA2JKZJlbGjDX8yNq80PkJqgiP2ejB2FQaOulb7tQLSFzL7fSVzu
pWI9vT/ghMUrx1U8qYKjn/0chRlWuC3gK+6gehQ2S1Dhx3kyrqX5dsV9nAYQNoRX7xYxeiSwv0hk
hKKVLJ2DvmCQ6RA+u4puGUcG8TdH4EphiQ63q1ippUv9IdQQ5ohpdljuaZ4LSgzP5eIY+GbadIt/
dx/OFcRBqMvDamBqMmzlGLFAhelu+OGR7n1zRZq/Zm0/xwxrcNAmohYgCIQVt4LiBw6XvYHaJ9+q
22ozWLtzZGB1BG8oGu2mHiNLYRlnBO/ZlW6iai9m78PlABV0Bd3QncCVOlDGc26FkIcOrAdGmSJl
/cwnkKbK5rwU9EHix1eSvtLKWRse6YP8dX1wfSGBXIEiYYe04oGvGHhsoVFsap3jJFFSNOJDJ8Yc
P3k1YyQ6oBRXnOPg3rCOVuXu8Dyoe/NpyOUujBxOsOzfqA0GlJ+8yQMmrRDG1T9YWmusv9MHq80+
mEG7SKlmCNaAL8OPvF5H8UPNZuvMFw0hq1e6nquHi2uoJ7HONuhK4GQMWbNEyvbK52V8cJuWybaP
LUPqdPLHH4N1CLNhI5AcOu6saUXxkRovKnTS0Lum/WepT2zrzMvFOh05rBpxpe7b0x01xF/WuTC4
o8C3EYt10R2ccBiggdYWvya3gvrvNzvbqC95c9V5CU1ZqNBz92jUgVn2ZtVlCjslf6CiW0yScWIu
TFgLWzb4QHSXiTEYCw7tFc7huRBcd/5lBCkWhvqqL5vVIL42gs+kIntSdbjY8yz5m68ENkwowVvI
c+y2cF1xa2W6kIb9Yly8Ebgmh5vZkIG1w+zXe/HbWuW2o4cBSAoFp5m0w0QwTFeuRCzCZhmT7rJA
yMjdvyMf44cHeOUMHRLGHKjKimStjsVRy6RPmmUc7PYVS2j4ZHNoIkI63BxqE4IQUGHUE+RS4LfG
I0Ea2ueU3i0XZUTgy9vkiCDIKjYBjjemjdhVTXoymL1CunL7cWfgu3JHnotfK8kU5/nabS/iKQyA
DZEQrADPrwH4bLO5Ao6IfjgN6oUIeK+9+kBvSV+lhBiiOVibCdsY2nPAmOXJeBsoLVPbYTFW8tPD
eJOSeh+JwxpUp95HvURqiuqlSDLhovu3DEABrhz15Z9CSfC8EvGlabL8Ua43/U0v+s5WvjKDvasH
EjN4vVNtBDopYwNoaRdKogxtWnm3Wipd4KjYJep5cq9jcHHz3Ht80ZeIJdel24i+ar1Fn1YZrgWh
HBgwIPSh0XpHxfEi4+lmYNy3Rb+X3wt8gqGAX73T4q182KajulY0ZA65S9Z+fr7yahpEgDohSGBK
iC7zYfugmzHYI0vdWMvrEAAEYnhgxfASqF8Xka+kBSol52qqWm9bb+u0pdYBVty45V1havwa5slG
qeLCMftq3OpoSxMNAOL2Be7vSZurVLXgf25W/VnYjEgq6eESiflAo0a3qZVO0cr4oUvc8ajYTmnC
nJFEOdv3CWjgQjFmgaZYlqFNVS/ap9VB6UhKNAsGtD4furQnG5L695/AIXxgqjkoknG2YsvTMn2m
wyqOh2QFI04Fr5hbb5z7DeaRCqztNtzJgpZmg7lFn3KB1PpuKGw8a3X5K/awa4RMQKicHnqTFDx8
4bYALKsXJzvWOecp0/5IMyXPfwr4cjQGTjlEBVgYXB6YNFEgCVJdtSgVrFiqEc1wxplH3gtYcX9/
Y4q5Gl5qEyG74BTwyVddhrla/y5uLWivgCIGVLBXFJaJT4Xwd7ihM6vDIECEuqnuzfAO9aem1/Fk
wunvJHfU3QTFsCiFFmFXDRldnsk2qM5QCyPHTyBqBwhVCn8AE4kaReVzPOcZzKWcVGUlzAnA6GZo
fEaOJWN2w919zAFB+3d3sqXcQ7R3Yr8HRfeVu1SHvRphKI+P9UpoWB/D/yUB9XsWl3h27nAeUL8b
OXHgwVQRLoMFnNsVBGM3JjmGjxkQ32mgaeaQ7J1qOZHze1L0PQviFAkWIU5OzyVYmSsx9js1LvLI
jHaEYASviGONE4Jc6pSwvJiqmxtLLy6xYVP+xDJMoewkyJQkyTHLxva9139iWEeOUK3fRmidxF8p
0ZLHk3eEiAjuk+Z9QEtnXyJX6WmsNJLQYCkBbFTeexTlt4eY8lWVAXJ7PV4sNi1SWYVsYoLXL6fU
jkl7PxWIZ+nW7B+dNkSB6WjEHyLX3v7uzetu1pw1WOcgmFwD/YEPzJR8kr4ngpszfIZlzxHXxhNt
56mnwaxI+FOEeBbEXDOqCWEUdiJ384BaxSrJBcB+0ToEXF6v38m0PRBerAbQ6RvpzXqoWX23ugb3
bMhHTJg3+FiIyxmANDgXT9x1hy1Yf0j6OwkoEzIqC2kjOPTz8GniuPZRtIaFFwkfpZsCc+Efcku8
2SViZlw7bWS0jMuZWyiwJr7T84pTNiNFJhDAAYwXPkjBnr8OxPTV8rVdYQbPbGh+yIcK9VuKQ51i
5V3yDvvqEe//q0yBt/yuuxsOIWU7XAUzi3Dl1Ze9jZ+MaS/6JRu1Mk6g0La7KvWIqNBxwV04XIFd
DjdPFV3HWM9+SA8wrUHj5/kr1CMzq8DfzhkzbPbqQotWKVpWEl7FIGlQGTxCOSkq732gHl9lQJYY
TfHlvslpZHMtTY2pLVcM/2Qic43uWUkbh+9b/jzPVbz0Up+mnEnm9pokjHJ6d0UdfCpetIdKyiQ6
9wBU8fT1CuyESQbRdr8xfY3gsvJ5YBhNjUzg4BpcB6082cYtXgcHdc9yK/dY2r8f6cNlNmy3CHvF
wUr8KVbHcum9zUkoal3MU8nrhRi7tA6BnzFD+B/RkG5/nPHoSWeYDNuGyV8sCzW8tol25oik80Y1
5nTMcTenYEeKwzbEwOm7nYjhP/rXh5KLsT1s0UJm16YsgniDygcKYftgOzV3n9iOb1qeAhj8piAc
PCE+LnykZxwWfvzvh+1MjKVZ7JCkvi7llvoHkHexsh28qnCb3oBolyCV+PPu9DjMiokOTS/TPthd
AiOgBCtEM9KXfv57UBmPZ2WwEPjPW3zSzE0T5PYe54e5dLHoizPPpRs6eBRKfLjRPqnSfdvo5GoW
gi9cpYJeHwuH5azb5kBNjzJMQnBKi8ZxrMMnbQkXKXBn/cReODlS7FMRe02IBPh0jTXOAHlwL9HD
64hQLt1HApYJBXofn9VBoHzjTegAQBmgosEJsjGNJuk8x7hGzHs8zsIPTeMx9/kXwmCOPcFPg696
4tAyc3oYGa26CJmfbdF+fngiELmxcuy8nkTOweIaA8Fo04RNqrSFKILguv0MquXk/ii+UH25Rn1S
gjQNI2QvmFZsAfvSUFWXzO3mSlhA6qAqA1RnenaRuklq9izhYrENmhGIjQfFfMHk8s7yI56Cs+Zv
VfZpIGLmQM+ET/ZW4vtdnbu9tEirNalYP9z0Q1edfTn/N8/9YHi5msAEgrAeT6VUxQvGqgSUBlA1
gnGOhzm89kFfmA5X+UZvD6uX2BBJZA5he66csRknJHT8UNaDbAaP3I2pNNfwyI8Ey5+4ywyjngNo
Sv6HYrF21qUKt1p7T+pDOUO74Y3pWhozTj1IJTDRR8MiYlqI3/6akNV7DDyl9bTTcR7PC2FloCGC
N5rA3YM1bH18C6lj/HLw/uFBlTGAo3AlGuBliIrD5YRud+IFMgmNOhNV5RU4hs7dUUe9+fWDs+fB
Q91Uzxziw2Q6p01dtR4BzRIjP2/LiolCSEUlCOxm6zxeYKv3DmwkaJFlDDFRgbf/UP9/qWsyH71V
8xDURJ2Wns0jya7f5c7o3WMxR9J4soNeGoSSfV8tWYsvQGBO2a8jJ5atetRASLy6tD0ix+cDz1Tc
sIj9y6YxxwO+AX2Wa7o8beC2ldx8dxejHRZlNxreNgT/KqxrBTfSRfbO68BCerwEIErn01lwfKzT
Vfg1Z1GttF55gUHJqiunDMP9Jcmd5VFpdSSxyrZBI7Fdch4tMfSXYd/xHjO18xDOCDAbu8wR6HNC
R3+Qzb92sumw+vquN+yj5p5l7w+nycog7LUxTFW7Y9GHHigsu2QHH4vbSiGYEW/m9W3nwd5Y1Dr0
Rd+M9j5Fvj3Jruo5Ma03YQpGQTg1biY/FEYQ1AQw331t/79k8t2otBxuS+aW9OozPWApAYCinY53
1DC3f4sAM84bazb4LDHXe7Q1q52sG+6Fcs1m1AT6BpFqhMObA/cNgji6WzAVke8E2z4uRPerAUlv
JMWGIU92IZeqwB/XNhOyTXYO/SKk6YA6oSxM5ppUoiWNsgNkNMzBAfN3BUaFIA/BdlHrk8g9DonC
hqMKmePDUmZoUTguqLtSWrheKHHQGvaxMhQk6FeMNbHiXKU4w12eHDf5/56IqERroe5K3k5yNXY5
LnYrBym+DfGSLdxUByA4c+/SoAV2diamIlXGZNJuJG4uNdseOfkZWO3COhiS7sE1CuR4zxo0jTOx
830uLmF3gj+luxPFAiSHHjI6cvJ9PsNm1+gwBX2rAOeYK8inRusPZJex0QZ31mTiqsUHTlsOc2ya
mxHMe/z9pD3CsC5aecyyv03fBAFBkCbBbncihZD7N43Qe33eIXf8XzBodFzB74Yz3b9lfzPJzZ0v
Il+BrUoBJWXl2xPx9gc5kTYWenBWfqFfnFleetvcdw/FbmUzG3I0dg4ANL0rzLGfcIRbhbhcbBwc
13HJzjfLzrKsLTEl9qZFpDHGAwULYtAaM2VghYJ35A4K52h5a4jXWxiEe+75vaD78zRbKmGqtNQ2
17m7dcBbYho2gE2nC77EfMZOqosanhgGvD64E0f92x9kZOXHT4BaFE0ns6dpAQNTBJuhj0Gwtzpw
lMoBsizBnmX8+QQl/N2hCP3CW4ZifgzcmnfK+49bnSThF2gYGhlEOdrrESw6Rx9F2BXQJkm1O0vi
+uQqK1p5IBVYFA809MqPRJoaGBbvrMym7Hqgd3XTdBCEW4ITi/MPmd1CMnf+J8C4P4AspBLlg/fG
81itVn8cEE2+jRxNqFii3/XBYsJizwmICwJb2XrGhNt281JwUzrlbqMzbh2agX6LKkpLR73PQXXV
Uhnt5IcHcLGr9YiThEf/F3eseFHaDmRVmMbrs04ixH/kwDm5k5MQqr0+lzKd06doU7gne7e7X7cE
GpTsxzfvwgZ+oCCb9L1KV9rF89tVR8dwjbonTP8RhqH2ZknCeWBsIaJtXUO417xFPAvRey34pMED
bSWmme/6eqOBb8jdnwngZfzky7lel9BpCbh+H3O2X/OrcgRQE3z1obysOR9MqTL1wSf2m+LbvOZV
0ThjSm6s/A/luh4kH2nU9j4LrcdrIdeuxuhhKKFJY6PVQ8YWfmCuVuKf83vtqygdd8xlLrzkQglY
9BugzOnGMgE9fiTLlIOg/r5J2F8qWR1lmkat4oYj5umfXPw3E1PVAFl3cEveVpbEy9hkAUUSyt47
wmWfR1Jkic9eoQwpRKGYJxmwZnF7mPjbaV5iBic+rk+yRS4/EFzIsGZhmDkBxaOgrIfrFLU6F93A
IPIiaw/+piMLPCPpuzdxgAuL+tk5hompp7WqJFP+f/2IXpRsLw1dxm9XWSToUVgd0aYyJHyHz5yf
OawzLuLiTgBKdgc4Fh/kfGpouPIOBaqoL1KcU7mWvEt3z7P/zySGaCs0BVFxLQqhAgYjXbYCW2KH
a61Ywv/O5nIpR/PPmCqp37Oev8m0hQhOaXukw9PeDuA8YF5xPLMIedcCZ6xsOsaYOkO7CMJs+YWb
If8l+SfvN3/aTb3/3pII84StGGrnEGszG1BEitfU9oCmJJXBC38MGDf6AtcgvAzKpdudCdCi5WOd
MUp/EmXdkzwgtd/x9rMJ/zWg/k6zB5+4N2ahRqa60dw8kaYgNeo92RMP55YbuWSM4jiDW3H2WUgS
HYr1kXHJmQb7FpsMNVJ2QrwWGWnDv1KxY0DXe3Q/q4bcwjcsDgWiAQvjTaUr1bIa02IBdwI/2jqW
TFEgjx+MaLI0UjUFuu8ENk9QHp3JBAqsbqXJefod38nQP6A4zkeEEO3UeKXLn4rm6CJtWQjbzUXB
l25OJC+99c49McHuVbqBx/WpL4Mln2402hSpxifIW5gI0ZZZltBMO8NspBHc9QbHrWjvbVIEUHIi
tRJXsZ7IrVeBsQEfPGy9/f9HjhuNq++ALVh7OvDsIA0e93lSJ/qjmjYP3Pfof4ityAHKQbLC2JDS
ctMudGBiGVXw2PmZDUnPB4j6siSAqpPk47U+M6pVDxIsQfa9X2+gyy0DNC01HfI8Vv9VKncjG57g
FWmJ16a1SuVROxGzrS8MCxTNCHekKNH0MF3Io6MwyPpi8KQkWDzlthkIrNWgF2m+jLVwTp/yIcjn
roLDcsJeUb+pYJNuBcWs1Gl3jzL4gaQBGbRqt0f8quHHCwcq8F4buqobOfExrdcylIVS3ZXDXHDu
wZVJtQxrvRi6nBF9oIep9uCa4UxLUl2pM0lPo5F7DA5Mj8kiU7cppy+oBucXQewFSwBpjx9MF1fq
rG8YzA6B0iRo1ccq9XXnApW7oFgkrcGtc2stLqr0lL4RQabLDFq0Sso7WYzI/bmQU1/vMgYS4v7e
YiqJgC32p3lQj8rO6uUS6hCtqpOHIgqHZngcN9EIJANf+H0gL2hCBTjhGZHjQCIxRadLN792ho2T
N4dcDEk0uI2PHQgw9fopXIEwVOcI3njXSL9+HPnrBPNRfzrH4UQKcFpBcO+9k/ZIT25sfNCcWSJi
ZlaJcsLGtcDZWZ0tHzszvW3E1sMkv3U6IuX5iXtNb597Qr8hZpDGCYNU/pERQVSADcc0zT3fJ25p
aHkqfeaR62lknS3x3Pi9F3J/Iun9ZQeQ9Hj1G9m9ENQy9HbQ0SA5wqM3AknsAyZGtB2+qUfOP8r8
Ig5C0DszLjSrQULGaB7QsvwsvPzaG/m+7WLMr9OpXs9WkH1OLAHbO2yrM9eFKYvf2CgVr+1sRvsn
DxDvTPSCS6wFMCbrVoc1Qw57RFM3KiFg7kYWdI/8uPG1h+RS/y0xy5+1BdKWe2MFgxSHbfJ2AWJi
0f2KFRyeMAmcr+M6Dkxn869wj3jxuoaZKTP0pbL/61FWZ9wYhqr7PbQ996qzI1suLSjYsqCEtqoa
BZ3KduouxED1l0yE/Ji4gjh0Z0m9FXh6XY+cv8pnTyINCtb61fXOaQZ6sVJn31fxecMG+6sYjVO1
CsmTlqOjFtrUgSLy8luYA4VpRyoKkl5lRTWeghrQZqOBouzQF/GDXvSotLzCMn1l0Sm5L4b09Ei0
jQmBN0fdr4vmBPBksU2i1fmgYp67D3cGok251ttyWJIGuOBUrFUt7xdOCRxsm8ditihYQFnG1BeM
Jy8T6DTuWgMZfI+8ezJl3kIM1a86fkd1chDhdu+YBWn4XuqoTIjCadLXWXbU6jePJ7nLlGUH9CrQ
1CCLsR4tF95zpEHE6hSVvoV8xlocyq+8Inb4VDShvVkwKM58E+ArojyL6chnRtLIiE9AhZMKQ6FE
T8vVvy+/at7q/Qvtp9cmY2bVJ+53XtazIxGCazUnE/xNkTW+a4fElnwqTtPxvMeRVv2oY9UZk88v
in92664UA2JoKW2DTVxs/4a15jtR4MktR7hbvlKWQ1iIXXxrrnWIKGx0ovrICqoIP0Vb3uGaWU+h
Wt+rkn8ifbmYTJUo8X/laicH0qRI2P4cQj3AUUC1kngy5Gx0ZB/+lU2Dk7Idl/KmO7sGOcJ7EA4a
Ut/7MU9dVS4osAGX5QEdIjcCEdqbAYhglrxJ11Pv0gvaV3t9ylb+2zo4xMY2cSxgYIrIkskhKpk2
AKm8JWoiHxRTihEhNAoODYxLFSdCgzoPrrWlbyCvw9je7odgQKl8oeckq0ZedgbJSKD0f1HgyPIZ
nHB6D7OPP8rCCUQ4UFQ1pGOGwQm2nMVwh445hCD5y9isYaZ6dpBP7Qy3AbYPl2ynRVle/wZlknRG
tqxmpOv84OoOB7RdhpRRMBEDSwxWw1gqHy81Gt6OBSgpVN4YMeycViPGJNllXtnoa6tcLOJ6RGVJ
lnSsFISKtLuAIk/c3lNiFCTwwofM5gWZ0pS/+xi8M16cO0PPtFKdmtkF7l1+ABnvg4b1DSvQn7uN
OsMgId4xJs249GKnfNTEN8qlHrBLlUo66ULoeWuruKXviQzmwjuAC3csBI1AEHGuWCI0O82bwYAM
2knAivDdRjwJuG0/CZ8Plvx8P039eHlmn0gXiYWC8lHrQv4p1aA1ozWZ9APF5QJTaWIsM5nglXGJ
YCWYXfbtAsjauEB2HDAJHY0FRgIGQb4BDrIh+dIjiH29YaJ69kC4LQz2s5m+5aZvWvPnbJBtqqAa
THxI3PU4Bd9BtjQMQx0w6blJr3x/SO7taIFTQ3ENCcGFi0neJOqX/6KvgMX7XgnQkXvgj0lJ6gHu
ZfEO0mujLVwK57pfB3p2fqfk5397VLCVgCgtGjCTT/rZvwXePHXXnQQi8yp0+0F+8Aec/UE3v03i
qWCTffVUVv0KHCuh5FY1X9JYPfN/POfUaF4DSZUX9f4W3lwvaJ3MHGA5UDt/IcxUOZzydMjpwmMv
6yEBpR5Dqca/oqHjbYEVSc0GBYyJ6MrT1GfMiKsuMKlajNuCFulJhevjZFo3/t2IaDEedHQbgeCP
dEpq2bUkM6s9SertpwSAoxNSjNQvxPOJs3Tq/Zc/UijgVxBnx+PUdx7F80W0b/nxgd3ESulwd2Y9
JyXHi2+CH74fTx55TDNKxBrED6u5KTChEIE1sJgilJOnRq0UQd2M7zM1ugmj/YEQyKhpL8HCfJSq
YYHWXUE2QVwsba4MZZKJz6iY9Q9hLsM3dHvOz90ZGc4okBkxJOF7Z/UWOrBt6eQAoBe7UCGqaSKY
5JcitrVlF63x5PUNA9IoyaIbe2jTl7kzN8I9TueJ0Wo2+zAoDJiK+JcgiUPfXDstfLcw+nSvtaq/
oGADYS4W1mU46P0E1ucwSnYe66Q3VEpuM5OZNwe0F6WGWADr7S31t28pJ3VUgMhu9l9a7ozQyiHP
kqj3SfME8xgX5kQzPi0BA1JHfmyqLwtoQmEMV15PIKw5HU9NqspOBsNWJaLL8YCk6h4ziW3MRXS6
n5/hzumdnhqskSNUHL4xBwSpQr5kwie3mhy0uITd7VsDwOpW5QEKxYWxpb5GQcG+2PKeYfYK9hEr
oIV1culfIJ1lJOzzbH8hquwzYvm/C7kH+pYzW8+HJpM1NQOlYZDjqYPTeqdMdcD3QTTfnn1JE+vP
MOh3CzjA2NyRiMRApAjBq0b/k8AwfYDm0MOAdgeE3NvbbNr2RJ1Fnuz3rE4cX9Pl5lBuYpzwxcHQ
1mW1/d0cThOOa6CpOmzF7J2zsTR8wa6MuPHTN9xyqI6WTUG2meKI0Gti/70UWwPJGa3jReD75KrR
hjBKQDROKC+1Xef+1FkeOhh6M/xUOoY1a2yuyPOdLX8uWs71pOGcu+ZhPOwZ56xUrDh0x+4wlz7K
PFyotsNt3p7VJmwYDO//FQx92mqhzNBd/RvtZa06IF+lco+KPzuOF1W84QcXoGXR0a7PESe7gJSP
zqWW//+dXEg9T2lmN2qFhzx1VQVUIRQqPyfQ7Fweiq8ONdjRjxMuCrkGwdESA6SPG+guDfXhfMhk
2E/2/M1VkC22XilOEOLQLOFnReCRlWbEGHqYdgC+3xO8BSo+A40kl7GcUu1pNbYwUNCygTIE5F42
vo/tavWhUTH4Pld/vHxU604xaYNBT9GAE50exhSOlhUO/yE//r3ZVUWd9ZN6eTS13J7yZoF3lOrX
zGGFYs9Q/hai8mvxDnhwL6+z5AGXZZTnx69J+Vy1MU6IwS+/7G3HRgiW/zT/rmzjBZQbdThxnDTD
XfXqfwvrLm6DcbL3QMbNDyhKuEoJJubch1Z96tA3CN56TPsZ9XT135bPbId5gEniw/NN/YUNSdhT
qDbLK51SKC9Q+InGqcFoietpRWm+I6kOeFvE4QpelPvALcMc9nZWWKcgSyknpi4d00jrXXzY//xk
WLTyOdX6f+Z2oiH1loEml/PIQWC0nUNs6aYC5/wUsqvtNCSDU4dPsfDGWAJ/a9dSMkSIelOwEzh2
dfiMruqsfbbeATZ/C9YEskknIZCuVYMs6/AE26fJxn7Q4ZaZzHrt1atMa0/u9uqX8gkxZdGg0roO
MaVMDrIUFUa1shMFqdKOGi9Xzg/Y3XV5Pn0wCLK+zczqzCgh8+P8/w0gvGCW7hJq5i4LGCOwQgpj
Pd85LWG3SE4SRkd9hvQDg5y1o/pR44G4T1nZezuWDsXn2jrJiG9xxH0+b2//VbeEj/iaX5N4PGM3
RA2eUsXzRfNcT17MtdICVToymxnOo+Z6xBrpzsA6YuVleBCZedTkQgnIi+vWMNDUjSDgjKdrNq3h
G0ulK56nva5OIpToblgHTn5SFWD+iO2+2rDnu4CAhZ4sh3ARmmVwIci5d7FSubbDQz06t0XHJzZi
wxNyhc0J4t41MDXeZ6XWcfOglByh+FNwBOnwp+yP9+HKGJAA0OHGbeYbAySki5Gc5qEKvxDU1IRG
uA1DLaHPptcC+cbMkgCuOcZY8O1Ip44WwfotAtKkki6ER/L6vJG8VSWE2tdyEP7DOA1Coj3J2LwW
ZRpJmv1WfcmPNoGVx/HKyv2Ue23w1/Pvual881nnEeSGQ6Cke2HXAjOOHXdQv6a5jevRaEjYnb0s
bhizaMdEjfkocJf0e4QE1g/8r4VtSpXJVwQbJKhqd5WTS1LChoLM60CVsAmlDx4WFD8N1xjID9RP
j6Px2hd64gGjb6kjd0PY6RtWzexb8eXvoNq49bwcQflJT4BtG++x81axvOgqHV1ztJtTXC4Ria6B
kyHQFwnqLCp0T1+HxRu9jkU9fVTnHAeByucb2Pg9y7NSgQ+oa0OCy3xWcmUNP1oLpzNRxSeADjJ+
sZzP/ssiYh+fMvyfxPLHnRRV6XDUQ4thVS0yZy7B+sV+WZnuE0EB8sibJiknfi5BqS2SQtGMSfOn
cST15p0UpyjfyZ0Meoi2brw9MpxoNFRo+XsjaQ536lbpBcloVQB1FQYw2BH4HuRAZ/W2018brTd3
0X1pBAlEKwW5ZIBOQqlAJ9L6lUAQkGoy/Hd4P7Q+6sbunvafG77qT/69xrLbabnfCZD/q9aE6Pu7
nT5R+ezZnQItghPovKPqhc8iUsTVzMP79WifWQ+z9wx5H/YEWzogi0RmEaN+qJki6/sounQd4sxy
IEPqKkLFNifnNzjfoClBi/BRCru+u8bUUkOA6V56mP19rjZTzNbI23KQDOFzj4AAKFF85Len+Nea
aMtkXXUCK4hcvxGLDqHiI4e3VjY6dlBJcDNnix/EQWny9UpHPZMhrk0IN/TgahmPAl3t/so7PD6v
vUgJhiZQEU6Iy2KHV9EkFt0yEZgAJOiksqIXlzIYntXx+G+mSMJK3V7Q+qZ8VyGninhqU75gX5qv
cFQ1bWcS9//30qdaKQwylXJ0jddcltPtHKPfkK5pPY3F1dJ35H4mBAVmn9zEsO+ArkJtbBjkprZB
bXnIcZ765+ukxIqqyJByLquJsm+XW+lXOXhuyj2mm0mjIiTTnzDbwwk/DR307nrPtDP1G8lNQnl+
U2utqjl2AuQFMwiKi1TltN+KR3rkilHi2jRvg0Co6MQZLDA0yZNesYtgzukJRxeJHfbpd9hmYBm5
cv1IaNdKiFX5Ofr+rsPes69S0QDTaSo427ARXCkc5gamnx7Hv2+5SDJWZvMkdOAZ6VezTz+HU+2Z
SgwaQoTTpryVjX7n70o9shc+U3MktWXKVCk0dcBQ/uPyU7A3FiSdClPdEs6AfAH3bv3hk7EZB11G
9nrDYcu7Qx6s21n8j+dTCMKduojYHj68yDpPRFaIEfxPF248nYM7eUZkYWzrT9lO0k22VBbjRnun
22KGupIaI8LLaswO8fv6ajSndW0NAKCKyzzHOQqmexEypl5EfAlVfsdcgZaDaQ4A8Cx6yoQvhjQg
ae/HCCTLxKVrvKejsuVfwkyS0oisBVABWHolHxEbkgLL2LqVq3POGoGQ3nwaHpRbryH6ZL+3vVug
06LAbMTecNmm+jUJO0ErwFjYj9DGw8SeiVIeKmAitTHSLmsDo4JvpcagdXp4u5glzZmhookIPAPG
+zn1E+6IEd3gZzMYfJ74ISDBbD4EAx30WqlVWScFcFTmr5P1NXjN6cdWqtM0w63w3ESIaop7+JMU
lAaVVFEzi7koQLafiVjC6sEIWEx2SuxDOBTW7LR6SNndmbqLRHChx3/YIExDa2LCQFXdpTwLwl1A
7v12CX3cM6p4tk6eU/JIo5wvvi053wgHSBgpyoy8pq4kWaARdu7k0L3hEvEMzinXhu3ikc4nHAP7
ArA05vw7qmm8DQPb+msL2g6rSlTaOpn9QoBakaTKpro8zx4jZpZcCNHfbCAf+SmE3Z0lP/M+l0HY
8zKNMY1yCqPzMSWJXzhWn2/JaEeA1gdqzteXg9lNDkyqA4elCsYLcxVtBBgOfB7hN7UkTqZUJCYf
WyFeh3dFFr1/8LKQv6h/qAHCytraa0JKJl54C9xTuO/S32rJLgEd5UcjWsmMSyKqTUYVyeq6rFYG
qTACj73exw4YBULvwNzJH4UwxV6wz65pEaJbnXL1tQcISuyOrjazRrJSuXO4oku5SVn3vCwvE9uU
k8Fio/bRrVpeye40o2lZvxXIOcmvTFdkELokLBWr1vI9qYdxKBLyb6lDlgxUAE1HLGU9AwqPDS6V
QtUJC5QrWCwS5qmQlRyAajxNpkOLnXcfvrG6DM+eTe0fevT9LifjkU7AURftr1BcnaqtXP9GKcHO
xpFbCvKacTABG3JVAI6B92XBKVtwLx3NRJkwzerNg4iNSpHfTo6Psi+pyCDNOSnRy+OFYxOtRTXi
2n2KaqXe8C//n/Q7yb7g4RKKBeQcDIL6rzo9zitefcj0DzrgnE7KyGaEIWSkSkizEanCsYJQe5B5
JDbtX2onmFj/BgDd03LfnBXkFpVaFzlgpcpxVkbLfQhYbbRP9HoVF2V8DmGfYVgSzOIwGOKW0paD
5hdNVQ/LR7+gXRiGwLzmVpSGaH37AFTtFugGOur4HRqEtZf061NlRWQbnZFU/acdnpVuAbJ53/e9
IwbVMBqkNINMRZsCIkcuInEHCUkRPQGb/wqQVRkUk60CaQUftFVT7XPUUbq1fYmnrM4ZDv0An9Vl
YL1DvSA25/zZsTSCL85Q1Dghl3OOMJFjpuM2qVtD+NPdNtQwT4EIjsKdzyK7pnSelu+EK0ikRifJ
BNEx8ggshXyjQzGm17/5k9IrdpfLSCT59XH+RgikvFVsESXDSa6fDlmaKNJAXxKE93hEbZvK4NuX
sVb6dV96NFDhjn+Q/7YzcTprgF+OdL9PnOco0X3d8ramxCBsJc6VGOnVn/vE/kxRRADnwEfPv2Aq
70YO7Z9bjf5JZvpUe/LxnMBt9zkHxfUCscal+wrVgzs75RBYX2tcrXzhcqCBw1bqCDD50lN4gXuX
uyKrPgGXhf+0Jp/+5p1WsDJB/MSa4i97EgfSETQnfUdOyIp/CuA9vuQOdzL5HchtPSOdvlJn5+qG
MAQnm20zvHqtnjfW/8lIAYZv/IIwr7ICfLja8JHiviBly74NGxh8p7ZIEuF7fb1sW4Ga2LCrHTVU
QybvmcwHN62agL7Qi+PLObIYH9IL4X7gRgdecf/gR+ZwKVFe33XscegIuz9T/uvZRLkroweZJJXm
ZMxnNgY5B1YRsyddO8XillnJd6+maZPxTbUvFwzh/YCYsqA3oFWbcJv7zast1lQiuZGGuYeG/VQ6
N8gQ8reDwl4XtjbDZ0gD5vAjtabTPzgFZZVK9v/5aCSyV/fmNKpEQNtUAkFEvWfH+kV7lf7YZGu8
2o7kuqp/CXvSioOq4YIpg/7zy7Ka4esidRdq6OTTEnKtKhv2TLhk62X7GR+M6kQAClZcwrO7kKlw
4tN23AUH5PnEAl47WXnqT0fa+pDW/ZCBsoDcP/v5hP9Obeh0YF+2VTCduTxlMZnG0l5+TbFKAqqJ
ibG6/LVnwBUaxMNLGm2HPDXem+x3iTAEKeJgHAQZ0hfBs5d3oQ8Jg7OZHsWUQ7/B6KF0QCZGxaGS
vqWgk1QT6hzPr51XPo37C21fHoF3Q3UibW0wnDYQKnPhtixCUY2S3gqlzPgyaCXJUUnZK9Hq7/GM
pvv6tyeP+mYjeM8/LRz4dfbezLbcAShXhbR78wxSweZSoc7et5OH+5WTanT74PKTmX00bXMKoXrR
+tC8jEiTS3qH//VRKeDkS9SAiSkBfDaXTRuJDaDtsmQ0mXRdZeBMVUlEYQfFwP/FgTEpCq9P5Kx6
+9OEmSdy7VEdln3dNpcDDskTIElwLONa4aA2qLzyjiXRDHmnPmjLmlGXWgxMtFOT3M+2xWYI0GeE
I8s56DuI50qCMlDu/x/4AmvhUDwGdULcqZNtAU1/fi+ZYQGCw+V+8ohPNgWwqtsUHPy7VQo3LJyd
izE8y+4KXjxQkmbPmgjrJMR1rtlyGX80aRO0DIi+cKgCh4+e3Qd9Xsh5Uh0ngzeWww5PV9jQQWL8
tL2OHOLZoBGxBbuEtjJDdLLnvlJtmon7QiBhWAL5dVsJTyF+XfbVj0Igv/Vw2QJnlqPpzzxkPeS4
ZNJSgMhcTEAGoK8qBsymbinX9V8EwxvvP2tVDeF42XlCQRM01rwkosPN6s+m2+rJ2PkYZQTdXQSk
uCuHQbgb+//ZyQUeAEn/+lNVZqIrIIVSw4zYecet/n6CXJO+nG0i6t8pNhDUcyEgKwX+8ataR7wr
zxkEbgLWjOvfhBLOtSLVX1jlIdOZADQgGJisOzwb3j1dkXi0MPm+tx4CYwH068/cZZ65d8YkeoKY
ZuRDvlhFfWovvb5D6dkp60qFtA8YWuGIJpwkkEU833Oy9Sp+dzXq54L4cOsog1vbcCXJ4STZXoQ3
YwDkApDeasywp6HipHIcr1nJrfBHcBSz1C0Li+NNYmjiEzSFbcsDteng/HlKF6jnxIhhuqDZrnN7
Lc+eO3RJh/D8cn/UWo3TCIESv6MSUXbyCXy1otL4QCbdryB29Gceg2oQBPwvrVuRzFnlVBPz3Lbb
Z8pzvbxpHoV5Qj9aSXASvJTdGQToCSuhXi2LrLFtrJDyousQJDR6ocjB38dSBReCFuQD2E3mPSrj
rDajgcHg0A0qpE6Xh4VOGEKSYD8ADwI68w8tzEkQU7MJuboWjSLO8vKYVyr+D0Hq8Ir6nS63MNCo
Sg9hoqqZKB9/Lw3r1sAkwxFmK/tzxqwlavNiws7mafV2nNW20+pWL65nMgMW7DeAZXwfdvEl9FgG
+i2RyyMV+I8gVrfd6flzST4b1S7e876Y8h37eGT+cwyReRlxJFgwPK350WKkxYh6OvYMHw3yNfy9
wn1TjwUaZz5fSAmGpEEPXP1Rd5TMrhG9T4HFJ7PbDAFu8KB4Ll4xd2rgBDJN3YqJBMPwp2f4SNvP
j6d151NXARbSFp1pns2TcVDPNEgUq9bzpmmtIeI7Li5WF8UQ1hLgDHh3XChaSLlwCRX77qZbg2TA
iAXPnBSPBzJ4Lgufrzt7gTyc4dBxJhh0NkgiRAiHwu9d6V7YQVIAtY/SDEVno7WBnfPrJ2NjJiqd
8GaG7ITLL5DySwN02ARnLAiwbSct07XOGa/cRVbVRrF3h04sZa2uVdIzdBtHEAiq94uasJ7q4Gw+
rzOEqxCcHucPUZIEnu63USWen1ggoQOIYt7LGEG5Qc2wfIGvy66yqsDqyUrYLyf1qm9U404N+YOm
gYeSUbWtFz7J1+X6QR8u6a+LKmTsY5IjF1dM9K3Is+1r+QVqVXJkD1mzTrTldykoi3iHjoPjq+8x
g9PetcqFcUsCVcRILZupJT4CVoYqswabr3EkiVIWcBX9651AXLhfwjrUlDNdV34ty0w/oPngsgkm
sZpiHWwDDJhyKl1ERdOWWxYrjGMPmXmHQOzS/u6LB86frGgQon+voYAt+rneVEslPLhhvucXEp0o
Yd979RJk+YEw5ziafLnl92OoZlZpu4VV86eF7/SYD1X3b8+yJAKaol2BXKE/EfMdqILhrE5r4Twe
LL1n4QnujNra16AXK2eGJGlHG7FttStdv8Z6HKgtn2vSg4iqX8fZzRX2v6RcRJ/o86kZyjG7o8xR
PvYKApAu55Z7pRKoOPm8pv6G8CLHj5dfl6Q1lOA0BBwV96BaIfvuRLa9hGFMLSCeysO2HxW4fQQ9
3arveKD92JtD5CTl+Xzbr6gFPspYOLbyH7RiE39rVvJXb54zL4n3Qe4TYFHujnJd6XPBIpgbywhe
58lY0l/Gn8abV6bH014GAvVtOwB+cQHYXC/XEYIxlyR1t51CFEJyW+dri2nIRSZ2/oKZ9SRiM+Mq
lAARB1dxWeWwaqMwOg1uHD19twNcqgK+J7N6rX7nXkfkvOChF2d3iKFMGyDdxNGVpa6W8WIvRSIY
hF1VMsiCAHKEACm1YG75euGA37h19r9GhwuXmsgR3QYBuLF/eiIJ0Au1oMCySR39FdGEYzkETrAM
1Cq6ilFmn1tP7S5wJwalO9PjyIE6HbreI/6R7cvQv62K+5MjkYUFLYh/oKv6GvY6zHzt4TZ1o7jn
RlEauUUmsjyOc46EUxt6+bpLcxfZbrWlfqIPrbF5g+9l3OF7iurrEYquSS4BODY/ndyZd7nt3Lae
sys4ZHe7RXJzJ7VweK0UrUne1jsiWxL329dUd4T8LcpVwBYDO3L5CakLXPpKEx92Qtal8SE3bmb7
TpsC62pzZmfLsmtdFru7gt1fsi6eQ5FDbFDA1nevmE9ZpQSBWIQIUSkis8BPBoja7rpH9WNlNGd2
BeUMlMvsh78dGbQlGhLGTRJMcHrWRKheQUBlwPdjcUZfBznZiXG5z7ZCK8SxmS67rStMh4TgITbH
/bJ6irS9Ru9lX48i5lfso2ocJiiwflIAI19nGk2WqAPbro8s62u3YeUFNNUKffOAqYW59+y/bLA6
KUbFa1CP4A4xl+DlC5JCfVfcn+5Rfr/sobrjXGuUzhDzeYu6esHPO3ilvOgnyqbhAOLr0kKLgjDN
Ok2nL0cJCFgtMDn9t6qCATznlMD6G2l0pXVpvtfOGksuxatv5GSfButTtPcEfEdy6Rp1CEqf4dcD
f2EPeNAETm8qc/q51l0hz5BjTqgD1yEnd6bgP0xRXuK5NU6bHsHeQBN8mhI7DmgjnNHJnV897Mxd
izTVfjcDv/6Q/a7QU39XSP1wYeHd/OQb1U27Lzb0VbWzjwm6UA19CwKw9Ld7LwnbxKu3Ut5cK1SL
U95GXwP/DRH64J4nvQqVllD5BDGUIk7v/x1bhQdKiWv3t707KNsgZOSJfNX7pnxYGr5llU9XdqaP
b1vvPLaDuVb+6PnNPgEwh7VFBRveFs/Pvy0Ub0kQ8Bmoe1cN1nOgYCqo0axfc87K1+82owFMnnUE
ZBSMWQBOwfnKTFc6bj/EYBDBuawi6msVe8h75V0u7Zz8pWidK6Q1KmC34nljQ4RSZ1/9DllGkvm1
GwdWtWxSUnS1+24Ax37C1nOc3dPphyU39+jAzMNpeQx0CjPtIuPbinxFkRuiHkD9a7CVBVNKtLvf
7GuMfZciWH+XEiBNuiaR2DRys0z+QP5n18x1YKO5PlWA/9l+FTZUUEruTduNrqRFLJwrq0dyukjr
ZmV8WU3YufDP7WJyj8zA4/hfOOydOYM4CevZ1ssW3T5Kb4ig7ZNXFuwxyhZW9UIj8OHRc4jnq8LQ
Gyq9K851snIoRO52jQwlKq63v0u6Xg9dt8Pdp9LBfW5WgLYHlIvgFPFt5EDQWWPNhF6yd9SxjSK+
3YhCTnbO8nxluKReVX9JS01jQX5adq3LnHLqTX7l679wO3w21ACKUBn8bpGp8dcuQuIgzziCwtx7
0CrIkchWMmbzSbliDWn8vDq0mQqbyEG1354qJl2ESlX72JTIwFHY5tnZm+yvzR7AHwUkzGGzxgUY
km2qr/jjaNm1TPCoiL0hMZCxxhhNpOcExz4iooYPt7bIrFlChhUMGicnseFx/jVIzNQN4UFC9mDe
dMTW/33S48evomfhH8eN3J5S7xEEQcBrHZAT16XIRCo8gSET3lCeTe5GWKwrwhl7dUe/zMoRa97P
iomeEAnRKOJ7g8IIati385vKrZYs8qXHR86NZ3kegTBebTl26JlOBRSMOP6HvyS7KUV4BADailmj
kawnxcvO+YrlJQpwwYphHf50hf2tViMnyQ9bFO/T+8Q7hCZbPZV1g1JcPMGRtvUyC7MqGBKOwbUV
JNuApjm/cCb/44WDMzQxVd11DEr1Mwu1KiwONXAE0MkXsUQlgtxlYm9iI/H3oMhXmcUuGmCT8/vm
ExqczLaMB5AHOL/tRg24eZcXcSOYsUzOL33p+pTCEqp/aqM2zt/eyCgDRGlq5jZLnluXO55JqhSH
L9txf506sBP1i8dbqMnaeYlfBDLsyf90js45BRRXpQjUCBnM7j1630mDYUHUyP8I5RhYYejHhI6G
11kxHaL7TUjvnS2MiOpjyE43kJJ01x6YKMVd/vzJ6bLWpIjTsP6eZ0MyMVa8NOdu2k43NGP1VXw/
KxbkxNmNOFr4bwoY7H+y5sSBxscFDjlWmbwTx3rPgZys4xiYLq0uuO30yEMjGpdIudUYhAEA1Zej
K3I0NIvDoRsOXpAI2dVIwArHPvsPq8cQVz808Yg1iP69F46zoDQiXPpfh9ErZ3prV3faWJmSWc4C
1ZVKfUZkTmwFonIzehT/OGWjcxWzWQcY0xsQAs8wVsbUBv0RxrK5EPg6NIAN3jWzWnHybVOi3Xib
yYH4kj8E9o0UReWZayIS78EMok312VOfE5bqExYl3dDcKTZbSovKi+wkrSxTg6mdHICaeHzGdblB
SYrio6HdMIvtx/fZoogcOzFh0edOU/A5A4ESJpwgPHTNMdLcSxZOGiZkwGoclZjp2+jlurt7/9nE
QLnOD6xyx5TCrErFa+gXNvXK2XkMpJKlzrbpxevH9e/8NQ02kVbbFNB3x1xJkIhfj2Ajl3rkTQ61
oe0E81kmhlgRw5/LV8R9mkHjffQh5ppPQIbJwnmHuL2p8Lp08qUApsBaZFO3OrG9K+7R5Qo42RjZ
0cHgEx+AMaTgg9XDgYamiuxWUfLe9kzmb+RRiC8r8kG3sW6D5v1/p3iWNVoEQnmAhNM4qAtsuIGa
9LU/6+86lSvmNpE1YXEkD55VCVzX5Z+LyATwYrZhBmvN4E9pqChjZtZirPU8OSNBc2b52Mvb8nHt
AQ4USMl6iBApZEBPeC0F26WgF3tmbyp1L2jjgT9yujjBFEtnWO8Y16RnQU8LV1DuAtt6p8XzLPKk
yXLCrK/IgvxlAiGpvFcnbzIiDiXoq8eVrlYSZRYgecc7qeApJaQVWpsYTD3CgH5FMiRQSdsaznYz
TEyp71lDluX7QPO8hnZhZzPws2Ksci8ab4RuZZKY2BV3aBaDLzz53OgJ5cwIW0zojFBGwX+DsCTb
mnHnMh+dnRyG+U1Nx31FlNdNS6fFCxlveFyuo5/8MMrQER1mtv/1Ci7kb//ynWx+0x+d6D28zK4Y
gduT2o/UOx2bZLQ474aP3sC0NquPqSkyJUywUTjNTMEXc+xWAfWfE4X1yeOFxbeWYZEzhKqqAUCv
CoLXrY98OGiYWvDfmdzZBk7mBWhzNSYIGqDQZAI5zs87YH9dQVsyWnpiWbx7lT5kdK6drCheDobG
nxDZOzpTlQ3188s+hupiLwT2Z2sIHaM/mNdifwpOoxm0Ad4LR0qWZzODOWjND783MOfxoLBYscDe
F20RzpfM12vVE5F1uEscimakOffErMO8UTNEFYomT7Vq5g+Vp7zgP9IPiWtvMV2djuo+MDhUDNJ/
QV8bxPaJN2gtrv/IOEiqwh4KL1QSPm7EAp+BeCKM1GVS3GYqINwIXwtjPgDVVgu8bV0H6WwENoFc
lIO18bJZ3XLBLwWBH3he+8PjY9ha/6d84ZZWsTJsWe6xDpu0bkUsKkJ3wqNmP1vTJFV7hIe2T/ds
tNvumVcE6/hDRuoq1IUCUyL/r5pKApknZa64oIa6shEuwBtqxx0XYA5GJR1Rm3MA4TOzxFgfDrlY
WMfwVKNhV4BZOuVkg/E/zrbVUHn4ewfrvXA5lJeCEiSxGmIKpYXBl++E9BgUU0Tm9ZALrYT/G2fM
Gu9T4IxYW+UKto2LvMKD1bYDuekIgxMwupbqE8iGJ4M7TxiMrIrna0ozmf4eoNGateuWcq7r90Rf
1H1d63ofQ0UudXCHjAX1x51EiX1LPSEisu/q59oV1xVLgzMoqFh63rBTqKu8+aNjDCNSory8M278
ITfKlv+Xnm0fFbuLzPTgCrG9Px4t8C7snl9R7kXW0zRUuZX6z2qzcfPcorBZq/hfQvZnDwtDbw87
uqHoXO1pjtwQO/u5pG+XQJGbHN8dzere4ILMN6+tJhsdsjFVBjh+oGdqOK/6mOxIqHZJ1n5CO2zp
BEoq0bDHY74lVuVGqrpn+ZBrsz+1A985fNQKaSb20Zx2mMlU7qmfXSckr408Nc5uT3o/jFi9fnAs
0N6zbvr66+1kfmwyjj4yIWOeyoCztVOModvKugXwzZmnzjIq8SDP0fYI2I8Hp0sXeo6f6bBs25ix
ir7gMM9elcUUzIS1s5HJmp2rTDKoxm8f0k8/pD1g7BjbNmI6IpcSND/nM7uVSjL6yED6E0IVb+EB
LPYfbZTFRSu0YeOYAQ7Gh34Ot0FwSt/45hHjs6n0VyL0Ey9KnomuF2KG0D+w858BfyvkIw0qsBOi
BlW/jPibcV5Ylmx3T9cmmphxySf+xYT0CodP8CkWx6mR6jOzB8hbyodWv9x3vYfMNA0so6GZ7zmv
XW0LeCjpXiRdsjIpRFuTXcT9vci+VhYVlwt1u0VRpT75LrmYLE2MlHJCu8IOtjJdMGAm6YzzwRpa
2A8KkbZG8kefTVZq7u/8T0fkPkqaVHkktzYi++RnixvhV6SbvO0fH7kHFLMsSaQtI48B4whafqFO
LPZSCK8ePkh12qIAv9DYwIRC3vPb0o2z2681UXYiqGCQBQVj4iyRCzvcaZBgUicDrjSkA0d3ZlN6
rZWLHIViG/P5GsL7goNPJJprgse0PsVFGRt48R43OQGdc/7GEcNnd0wB/m+DmTKcPMK35mZV31hf
Kkj+lJbMB/HFqmgLaHCFrkmJwar/a4KHmCuW1Ld8fSHY4Xc5zPVfapaZdOebhqwDOguPk/I+t82I
pESG+oCfp6afawWFTizoGO5Mt5Mu0aTGGZRsLPns+P2CeXSESkmWuRKU32x3mB4MIT9o0UQJiBE7
ZUb8W9VU3Bk5HZ33hipF1lDFjzmJn9Bevz5O0QjVp7sdYb0BmlT0Uyd/XAU2Fna5ekzLe2ugV/ZW
KkeYt4SU4Quz1nZIJKNHynDnzVFBfK744Ur6+daz45/tzkAwYrwvPvjnP7F+JgwZGOEbjC/hACRd
WF1HsgbU8LyUK1o3+Ro3kxdNXvKjHqHj/DnmvovdI6Cvfu5gdTv4gM/LFxQxrjDHNNLUndSE3lMg
lSvx2ZuqazbI77yxDpENZRmsNrJjfNOW+HJpEIYrnAZRG2t3b7D3a/IgEe1dw8X/1lg0leScDzBG
N1w9f52ZjEAkum5+1s96ucoAoBrZSaknm5DfYxOXDvBXIvD+07BD9/80xwPz4HJRLjWRW8a6y4sO
MXFadVWKmJ5VUoKd05GFRBMkt8M1GyKr05XHTpzqHiRU1AyVNgMoZn/pgKWIPuYIN1tnN8+6Gt32
8OZTA1yHTJIpMoCnt90lQmR0qHowqS02BferGZS8p5lfR2WiGIBtwb5kSXok/syJo7vKiGv5DmOt
VA4HWoDwnAT8PudSUXO6WXU4garJbKkUYy6t45momcXHNADAeiHAktVSXNHgCTn64pnMb6BEeZ6m
w14XGVG5rS7QU1tYOLv37ZRVZk9IIBteEb1gMd2lODQr4H0pTWY5IhfxgE3L+b+2ngwwjTf7ILpt
bKjyfLtJLSdLY7is4r9/gQNMB4hvrgxK3nAz5XkDCBBGATsK2XAPgb1kvum20VtRx+TOdsNvzUnV
b+Dk/5OJgu6OX6G95JNW91ILMKZ4CPVmwmMo8mZoQpLJbyQxQPZEZQsFnNAKW7g8sjrPsnWaYSfg
94f7/FfTVxwVPN8/fP4DfNtKdgZq3Ly6HB0N0XR0cVj7t7V6cG/OjSc4K+P/8nHQqmPEGuJ2NU7r
R22Kf8Y8lEFqFhYb5Gs8VLfzcVYAqUbwe64Uycc+O3YO/SF06cd2tYQ5cVaMeisVHX0xef0zAU67
QWTwFiTzIfFQB8zDZ1IfHkx5x5w3aKzzKPVi8lchOuLwzahngkagpuMREONibDhBJGaN0I9zCC5u
7WjmOnAgPSDNVwCiiaoW1CjhaKeZQy9YvhVDki6MleV7wavjvVJPOur5sxMJGl1VNNO37VgfhcUV
k6qtVyXOTWld5MYY3/KbjdHRvQnLx5zQoUzwdO+A/0aJQorsKv5q60jXSA3iTeu4Vf/hbIGeevmn
+r+W4THkkpEgjdaXV5nuJ4/BGswiDdiS6Nz5fv8fs4W0yjffjsvd6v4LPsfIJa1m8tSAFm/yConG
IWIH503V9IkMpIA7TLnX24Q8B6rF7DW60N/6bs8ipTbOVXMLuyyBR+LGpPpbRTfak6fOA1wq/ARU
dsvdSi7cPSdVjx33WjyI1Xv2iYG8pBC1TO0EgDc7V+vqNsUscUQXO0WkKyJNvfNtzUll4ROZDHKd
mh5K9RLOph4AjRtmNDKC5g6Hjhqn8TOU74RJ5alMYMiPMbmP05YRAOt+8z6fvtZE46f8gyXOfsrh
uFmx6XZUO7D9UH84FNTGigZflmu+ULUuBeM205Gp9/CeyY4wuYiN5RG6k1R0iX+m0JfxtD2ZZtxw
34wxJt3d9cRWc0hf2IH9T2yQSu3ZU9ZXHlnRzgnbgMy/dakFpruw017uW2NZfBgGzWamHHQqjfkS
Sp6FrwEROZ0G5VXMtwPY2+wgEryzluQQKxueVl543DjDZnKI2ooqDQU9pYT2Hbafewvgmdlq/K81
fB6e5+wJTcdT1oc3b8XROfYX6iTLEvOMxqgHGILU3hnwe/tVAX1epekFAbWqM5O4kLre/ktam8jk
iKwU5BNM8fWp8yinLcoRjWWaeeqfbz2W0u44r+931kMZpyjvafPKH5HeMLMxSRrgJ9vnYqDheFu7
1BUMxDKBPhKIGG7TWhn0JP7xt47dobV+qjaYzIYvhxgCi87JQnxNw6/BqD0Ta7gWGjeqGxx1F8sf
dcYAQ9szHfS83OPrKypYJsfDwa6ZzpwgFn+BMR64nIWlY29LsjD1WtRkXKq78xzZ/acj7vTbHk/4
Dd3DYCN4w8OUgnL/BD84z3BdPdqZIjwWDt5SBQKrbTvClDoPsypFgNE1f0pImvCk7PCBi/FASLWl
zoMDawPHxC2SY820U3w8svXVZQnBpGiis5W6O2rA8nZ4gsotVeg06bEYb8TR1supQ0fnow8fiYZ7
oJA9hwJvfeuEENK+EU9W1sebiiUbU3g9SZsqieZMoIFhoIYcdjzeDD2WKZtQ+6j55KuT7Sb00/Yr
eWCX4FBB2iH8uaj7A+cPW8eg4eKRHHZETN5M8SIkcHfBEwIXh2tHPvXO/s+SQ6vYSCPMaoGbFoj7
desfXhqaLth520qjE35n01fF9bhO2Yk2sf7Fhvc17zw7Zzj+BSQ2Fvp6bEHipK1LQnlCKLlQpevP
wFAtq5T8wqLpkaJ1YXrnBJLabYIpxmu5gCJpzZGiw+2tInXDrTBFHrDPaOoi5WorY1hP7wKn0FII
mIA4YdflA5emFwP0owDM0//0J1yHkLSUTm7VQWRHOeYkaUZ5FdWEp13zv1tYAqfHbT71VzhAvWcD
1MzGjvYqXqhUzwju7rFQVd5e+paWBauuhj1CNVyaH7sNJ7byem8AtATShRf/OjJnf3aK0JA7G47E
gccu1nrCUIWi5bsDGuscB9G29rihh/3eNRiRzfFO55tUCbOu/g4yYguYhJK+GbX6esJi3PpJ8RgM
OikroAEodwcpd2UUOt0Pg/kB0o1JbUt8PLNTVXWprndmN91kITcXsRy13h9Hnm7yoteGLjmXcn2d
nFdXQPs2f7I619m5hgUeUGYNv4vtpD9SIUHqIePQFsvEVayk0/spx6ELzr8IKgUdLAgOf1rkNkJN
mdI+cCtqHQrD2CU7Hkcb5oaVpQoLHX8f9iK3ZfZDJaRoIED6VK51m0VTtU2I8VBiqCvbUc4KlVL9
YxGgix9900Z3t9M+HJwDAc3CPz4SqeZOxc0Vd05dfR5psLwYesPT7zxfj0BIv6SeVL5Xuem1XhkF
i1Gory3z1c/L5UzWpK5+daoazy/FE2OimyaUZenkCG/ONl5WsY2s0nQlxjmXi8p7HnM9En0WbGXM
LDtgE1EkxIO0x2BbEQghhyAwEQXKTnoZbWoCE9kjmEt1xv6bRjVTzu6l9AxpvA45oxbmE2xv1wvF
QUWhqIZKFc/dUcGIs8hofkWfylwWfh6C1a2lDSKevDhoo/antS91XnNKprpXw9CcIaJfhXx8C1YU
OjevNl7+OWSQUQtMeZbt9QpBwaWe0sLYs7WAStQSrqXHwzM0w+aJiWVG+xj797BMfq21iXLlle0q
ULW9VJRRnYUsOh01HIX0rBxCfyydO95bI4FBkdX1hvL7eA28M+wniScR+MM4HaJft0I5tX66GxO5
FqmeCIhSqP2A4FRKijWm7nMiqVgN7pdYBBajBfiYMEvlQUjfSUrrsnuvOVSbp3i9DRdjpumf1ROc
7wOU0vfUaMUShcsk5WBBePjQduZS2w8W+2jXAxF/MzlOiYmCrXRq48wGWjBQmmUkw74cKgAuVP12
xiN9KHRMDjB/lNZ7tzIjnyzVBzD0vlR8vXSRSqBVvgZzFhaZQkV629BKrnOSWYZnMueUrVjguoQc
b8QS5EYfr9CPaQKJTptMvdrrojma7iqeCr67BzOjBosv2uQgZ6ncgrmQziqraLB6kKx2CF4UCaPd
ge8bNlu1egNpx3oqYODNN7554h5o5jYWW2yOPjvvhsnpb3TG6r3MveA4vvQB/87D09NWs/MvulyF
bT+eeMWT/TrgBny293+9dkrL5IR1T0JEPaWkVmkmtpSP8HJreAwyYWQFIm7AnK2O5XEfwgxXpghF
RvDh7uT5R8fbtkScXTSXtAhYPP8P6nLUQWEpNWhEd1AJNDX54UrPCvccrECCcrmbl0gJljiqTVHm
yDQCBi40wrFUwZwstLv3t+t3+WJMbeSV8efvhuCR49k6429QRPQ9kExL8hy9KTyya41/osC9xunw
Br8iaurfw1SKPi6uqAl3LAq0owO48V86EXSWx08xPxyF0F6ib35rT0lU39VQ0PsRo3cGogcfr9Zh
YdrUuummdAHAQXmIKeYAkEHxMo8TLg21k+kAX1z3tPKCx1bBhNj+MPc/ScA8FnY2ScE3eqCuvAJu
j+TrmraKavoAWOCTIzpXr3gzhDE+9RbiekYQMdv8Ek8Xd/3ZavYnRtzkRY5+p5kz8bkWNvjYLdN/
JN4IY4BoclfK/uywkIPnVmqQnGmXNge7x6IG2A1bnPccpK00stqDnRi56WXAL121oygN/DS/QOq2
MdSvM/vMtrDZS22AAGs2gVXX8qUrU0PoCHAIhQPyASHjk4Wkm+nPd0+cMo59SJqt/1nl9AFtx3Bk
ofqoP/t2Zfpfx+3SQue+NfInWyaMgBkHvLVBIlNv9I/4xAApt2u6Eqecu311id19fK6vMt7H7DDo
obt4Y5d6BMorRyKx25MNpAy/DG706yASqm4k3+JM7pi7p2aQ4KfG5y2fPl3Mi9ZSsBq+uup1jR5/
c0ZwqGg5pQOV9qkZxk5YQq16sPLRkzUga9y+AsrmVcu2N3RM6yf33f8BL/QLHEMm20ga0c5qzAms
g3ReD0r/WTsuTlZu6ETREr+o3/bXeUbeP7GKHyY1/Cng6cU9ifferx1+1QIo520eCHtHnIqrbzJk
BEqZLTNyby4n4OeyOhBIMlHU4+IXQURrMw0vH4RknosQ3OnluefERC7Pu7R8cA/e2rL7LHlqfnmh
PISQ8xFyig7xsyhMEHg6le8eLa3qBNeqDa41kYX+vYNpk7hyVpk+Ma0MTS/dI7SrsBXKjHzzyXiJ
0z/8S6h0GX0PGsff4TYIFIqypVkMjA5SHnMbS58+1f5x9LLErYLUGOddP68Jr0suIOQp0+1FlbvX
EI69KvvkrPnuYuOP7Rwqmwldir7B84TtVNsmWXYvbHiVSYezyx584N4YJdX1xsyvA19ubExGkpli
nejRwtf6qDYhDOVQ6U0YkhPlOQvDHiV/cKQCo3fsC85lHgODsNRAtoF46NvmrAvgprXcZuhbbn8i
dcciq9xJD9MtKEY4fLQqfsPh1NMGSYsFXZCrCHTp6xtRkwuvGOiT/reJHVIBz5cnNEZ3pgPRFiTn
g16ze0Gb5m1U/1454nunRwayDAV1S6b1n3uDGUQSjqoU0qkWO52uNzwhnRbhG2Q9i93rlicpXChb
p4z6s5VdzipUnREWQ4/KRFZx4x/GtA6ryYuDeuojrG4ObK7Iu+9kJA1JLKwOOLm8YDOyh/d9STzf
P7YyFms6p2FwXitaJq1QHk77Yj5cneh3xSs78QFoI1cziOFTE5l1xU2y8ooTiuKGINSeFTxo4QTH
hZ25vi7GuPypQ2f5LLtP1Mm2tS2UBwhKE79uliC+NBrJbiqWt1bb9hQJJRKp5Opg+7DnAakqTkIy
TebzYncidZ1O8qNqIDf5d3R61N5iVP7SVo/WPx0SN4/LgFRjBgJ7v+mVuAQxBNVknzULkuiOARdc
UrYPEHWf9t6o1I0sw/pqI2n5hi7xwkmU7cZzKQhMA0DATLTqij2Edf66tJVQ3gWFRSkZW+s7MuUB
OmT7RfGzxmmkn2qjN2cPmQB5CDdZLIyGMvb0dfaYxNS+qEbXSZC5lfzYGli46P+/hTvDCXvGvFEU
L7HswVjOxa4p07SAiusWDtxFbsbgRkJTUvGDhn72yzDXP2CWNryktbKqOD+5V8oQ88wtCJsJ5nRE
zluKpeCo392dJcbxQn485OC5Qt6nYL4jG6JehTzcdSg8MnF/Iv5bcHgGr4RhnTi6LyVCxGItvi0O
3/QRHmtd1yp12cvM7X/eJyUNLsRbtPc6BatNhiRITMi00DwZJMqsGirqiFy7qlR0W9IfQWdDtvqR
agJpXw1wgHH6h3hpYMjLRGgScmE7TAS3aaMcvxcaPROHQpeUZcD4m9kKJmXtqgRksRqzzbmc31wP
8o/JwvpEluSTTWMneqtxm04btOCFo+hB19eapLEHhDMPXHnpqAM5jMy40LhNxLarKAdnrBp52pLN
vO7Ky03jE2UrrfTcmx2GmSZJ1osdpl+8lB0q1nIZJp307Nd/6RltvrwFEK2irlo89R3OPjaX42S1
SKysCCygvmvob0RfkBMMPGnJ2+Aniiff/1uMTEz1vIfYDKYsLVnIdLHb/y3JMXXnEoQPHr75VGwa
zKYmcu/+7GsnQlb+Lwu93iT0jLUKDNpRAc+i8vd2a9oo5KCra26T/AN+ueq4AOmKee0NI56w7ytc
I9rpT8b86H8uvs1cTYrsYv28MJEkQ320ijdBSY/g2yW4+1kZRw322htRiURa854Rh/4zCfbUuY4C
d9dI+ETXMV6EL5CKeZFeWh94rTvJXs5lVjo0uhRzreklf+Q0Gt6facFt5UoWjUdwNT3zXZ6bVdHR
JsMLPJhUL/H0ps+7mOm3GzgU9m9VGnXboNQKFAvN5yaGF49N9nkrByGqyEtVGug+/gMeno4RPYoh
m1AHxJA3D36WCHWgZh09WkquiyuPU1Ho1EGa5XfZ+l1aHq8SiRx5NmGcGZEfRWeSJwjWkKDSgknp
3EcjX1qGPTQaXfsrvTtaiouLtNr3HsMhqzoqb2AX824AY6VZ6R51YvIpRf4Tduri4wKwgVdQznpg
y8//MuPNkFX8SLqQ6MprsxFT7rIbsUYgRm+jg/zXrt1rYUFPXy75Uoys0kDPXsHDfMj7VtYyuA/m
sUwzD95drFFPRCUt6ytH0xMwt99KoUAywokwX4vAXGfOikJjSDEXwUPd+tht9L+HusOqHvhNumrY
gDphcZABv782tIAvZ7ZUwtMTdtBoB3UtYNXxowErMHmr5i5KfM8NpiYLc/GU7vofQqVGmaivdY5Z
VBzJDzT50GPDC61rruGIWJEk48yDOGZs0ippiDR+CY7iYPjT3FsHFKZZQUBdLgIfQDYPtiD49gYR
G4RmnEn95FuHqCJFvvqFiHIE0IPj1VFmRFVSOGKcmEE7ozysRybXlE2j/JT57ykQiJfPZNmR01NB
A82b4pXth6RO3jJrN2BC07W1TvcD3OXjWHrLRBMDJaA1gwCCGoWJx6suZjSsVjkj6Ohxa1d4NGTK
epbbi2rZ0Kz/Oo4+opmS9MBwZtTzQoiGMTU/7dRIqLXPjGmvIEWEFevduP+uVByIYErMnHejLYZi
GSNBYMr4ARGrUCU62m7cOiKNrAkB6nQ8dGd9n/Pq5JHrcRUiEKTuoSgLwIIVF/O9wV6Ic0cBK2c2
DRM4aVObPrJCChgBt1eBU0dT8ILOjv6e1HeQJdr5I7dejGMQLpttYBF4OOHvQI7/FQqTCvFNLCSY
O+7qUFmdbCfvz6vAVQbhw++v19oxIFltzBWtiUUVKxfZUoQmZNfY6mdGtKqB9Al/wK//vI3jTHqv
cli6/jqTeYB0VE+S/FzHd/7CyCTf+deegcjmGYnuJ/XODiOKlVDkYgU49LvR/KNwyv8DFJdP15AQ
ac6LBdA5D0Vu4Y+o+2BOw+AdwHva4cxGQ97gf72QpGaV77XiCjabgXlDs9ahSG9jSYYtK2+H8VI+
Xp3idMBIDsjVc5KOw/+u8oO7D4rJjAUWzF4NWmi8jQhhtBs99fVGAW19qOIwdQI+UyK56XxjzZBn
oWmLd5x0lk6QvYiLRME49PqEP8tKPzEypfVSc83V0ESX0Q0qusyntOqYd4VL+kbAZerkA3WHziMD
nl4rc3DGN9EXmynsY9ELBHGkjaZkGQoPn0fMxkQRtXCQ7qSow4bukDviCyP9nQrXEQ0RFGYaeODc
BhalC8DLmUhwLEnSksCCXqiSsPeVUF1JFYOFDJyAwlXcWaCM9Elx+T8fOdFTeNQbfuy9sLZaEwg8
hatdkt9w5hSOwNRTpt+mF81Id6S7v/Vrmy3AC5IjSVLOW/xUpFSwtptHkCyJ3BWPqn1se8Xeqap0
6R2BS49IO3LtPZwdJ0OEky97zWsilJ5PqnUjg+3Kvj4NtbXNdRSnAa8dTYuHlzRKdd/R++djB5Tv
45r8KA58AMkS/OPU/cw6+gZn/5rKoyvzJ/hb4HkQyFeEDl01LmNC+5Fn9qngZcemQnNI3mDpynlY
5t34coot/DlTbuNuf0noSZQlvOGJk/1Y95IQ7coeHXhtfg5Mop8KqpoiljXghX7erOzXd2nv5Xp6
h3FdyNkmoYweQeStPsUsDedabBDXg/sutNVqWBRKlH/x49II/NExxFjkY+ua5/iBXgS9tWMeMmJ8
4AiD/oCg36nPm9zmtYChlBIv8GdJlROuugZ4E2cYcbQuENTJWGlVqyBxqW9oEXIoFWIPceeG+xH8
xOtuB0uJANJTN260g+vevR8lCwF9ONBtZEK4AalHQI3MX3Rvunolh803smO2oSnObK58Roi0/XFh
7vB0qia4U32cw5rA76z8JiT+GwGcIX7dvxQx/uniZ0/LuIMK6uocHzumT0rpgUsWg+MSalreOMlM
2lw1PigPv+ZyoiKo6+YKblbz/6vQLjXaUU0myY1rxee4SPGZQ8loavwqmLRapG1WnSDRdAyqB6Uw
Zk/YMX1LF/7OX0xSOADoQaYgGimyvsBSuvbE6AQfHP/y8uOgf5e82VrqHdU8+B3hTX7DFl6N9DhH
WiSHXZ+jkBzNrFdQ8PdaxOL7Ols/7ITYC275O9g+1QEYFRGtnsPmfbib9Yzl44EwbCq5WFMvGAPI
T6VsMa/mk1PA3wD7tlsi7dnvoXTS8Ft0/DugoWoxf7pO0TyjwWOJ18EKqLA69JmMJVwk5cgoiwBJ
2lil+F6WqPMQ9DnB5OO5G9hbgEfBF74H2QHPIB7fTNS1/vnVnjLig17QKoTwKsJUbons+Fk60pjt
xLcC7nkctvRfmmJB0SSjQBoWi5UhXX3OcwV4JuQkelrTubXBRS6b2u2rKciaVs6N3oIuZKNU/EN9
DE6qRfN4Ntk7WpOmjFmbSaJFRhMTHtiuNsH/GbK+bWBm8XvpRFR/37pJuZVGGbw469jQQbvpNZAn
nU42vW1oxH0S5y4ZvcQt2w4ajOZrHqc61bgmADDxu9/jPz77hLaMUt7zRQYoY1Cc41xDH3ph0u4l
drQGE38rHnxYAwbsx9ohz3jgoCsr2/ANUOrKyoJuu/x7QQcyMEp6qeQipxU0LYolQXUzJObkLDs6
pBVN+LkGVdftzpD0p4svQcgNln1N3cEZXpC/6ZRB8jWVylQg4MiJFUDhKHIw0BREP2AoFdWBcThr
40I6+u++uTx5G2HP671aPqRhLN8AK/mI+EETgBXT70+NiRXHDJ0FWumnb7iXRndsTY84yDoxhQm6
aUL7VPlQk6LoMdVcRs70e46sPecXfPl+450Vwnt9UOPDHfnn/gDIMpdVU6iK9rbRMmIbkq9dkbHv
3VtZVYn59Y0ET79z3AnW+aS+OMYexQu7q/hy4pp1VjKzqt+DT1m4iyZIMNeYvYY+MUQmC9nXPPtZ
uUqNj5QWaPB9vbm7jX0UNKgkDYgKTEuFZ6Xt8xN3NwjBQ/laHOdmZ9dVKpgjdpSWPKNhVFDe5dbe
nb3q8xCN9ULAefOFr8IDXrpln+zn7+XI+ZB6UOmDq2LPXoId7gCGst8af0RzetndLLyCiP/c8xu2
2tO1DNS89hodzt5xGu1Ma6T55+mXgTBsCm9ji7sy48XwaJLIzzEg84eSjdiHGF+0ZPt5bRP/cOn9
9YybjtkM0m8H1lhNiu9DRPqSBwdSfzD6W0xxglJd7BBEN2wYXXC5huAM+taMpurMHCPq6V8cePDV
ST26xQL/NLw9C3DIjYgbU4uE/SKlkqfXPvGng5p5GwncUNUDx4r2xTLNje0wOLwj27ezUzMnBmvK
k1pBneQDtPG2Oblviaalg194WVgOOYrB7P8O6JM/NUzv1rq9xHvmqQnqGcQmvY/aGMCApZtMMcdR
pgOmw/sYheCbBx/JiswbkIrSQKZ+2NniAoZz0BNbjFFYM/eeGUa8Ika7Y4GthNbGnHV3YvZwku0v
Rcc7AI9SzO75gnu4HDXbBsPIkWG5rn8ik44sboVLqxOeGTJquJzHpt1JlPNXpL06PtPXEwijxsCP
X4sBrJNF5ONxIlz5fv/jZX7GuYF9SIGyBvdHf65TWLt6xL93DbGsCmiZNbkH2vfusXX9SpP4Z/mT
l+XChATTZiMnotOgpSvym4pyVBgAoOWhINtF9ruJa+sREaQa10LEZtynEjMhbZ/viHJXgcUWTUj9
bPqhj27FYUt/gIhkhkobNIboHXriLOGwB37GplsKPjfUOCG1uEWxlfkLCPs+7tDHBOwNGQcqGMWt
dFMj90RTTAldEnDCFJVQUWBirau8YRYE1xJ8ry7PLNA4CjemjNKyKTRaaugqOU31XbzETJudy5pc
ixXoQ+HJcnASOB+gSeKCk5ROVTe7A09jCic/66zaaZFwBu8DcNLyDqvOLxF7DOzRcuoJ5g2N3b6s
CPoE0eARdWGQTCZl1AEopYBFUAYhqwZj8mSbP5n7QL8PivoX8W8uSZfRV46FBSJMTyX9SoqfS3TO
5paUrm5lk6GJZaAcUhIHVt2Z/6SVZ3NVGoq6BrZeQACZa/ZKRTb8+RZ56f6yTdqqKvef3ev0AtLg
1v5mQY73s1ZSXfpnOoxMcXdJ/TNtYnQPb5/slM2ijmThMocBUXjebO16BRGbD+Yd+x711gdgX1gU
n1OFhp3r3ev4PJOQXWooERUTkZfZYRFMxdxD3G2m8bg2pidtinMRfgpSqq5tHix2AZYkvVzUewL9
I7gmfDA9Ds29fJM1+VrQChrOf8r0hS/r+cx7p3jSVd/NPmAXBHH3/F6XObOtSq605DUoVmlnXKI2
vRwHifKopdCDZ2EgoHWvjVZP8kKxxhGPWFj4FNyjRHHiRmpJWgFN0Nhry1Tj8gmlp6G+2mMhzUCi
5zzQzsXrhLOvsO6YgT5XD643w5z2+uuswkVQ5YpXVd1RPV3jBsV9lbaEaePD0UHV9A3a6vWVhXd0
dcFo2UsuIm0oICIa34hOKiWXIzLaqCq9Vt9Ii0gl8m/8yaFxBlHuX+KXIlche74CdtOhXe4UetUr
RP+ZOe4QIeKwPrHI41gCA/cyX8jgEl8PdmIB4kh/6jwb4GEokaIaWc8B3AQn6ncRomCdOFkh8PPk
5XkCxn9J4lK7Lj6WtJfV7cLH/SStJ9mD5clLeWHCWpbRZHU0l+AI0gUHE+M0GUBlfj5gIq3GMOf7
RMrrsu/gj09nvm+xaqvEyVMuI8Fm+ag69rpBbnhWm/mOxB3mXcY1njxHpch7KDShbJ1wb4qkJ3ZN
6DFabIzsNu2Wy9ZBzfQUSVss1zmy52F6Go6bjAv2UttyTqEgPmlMWMXcOfBROJhFXjM9PlVZMd7G
uTcICwjRhTqsZbge/JYJfBcJuA3ItHgzbJWbn375tiPLbeWE3opzNtuxPn+oQbqelo/Bi9+PotFA
3PpONl6+N+3poPLTL2Noj/pd2OK3d2v8wWK+tvhnhh1K3lgCwWyQd1+kw7QkjoZRBh37sGzZ7puX
CX2ZBYK6dTKvCwp7vtdoM9w8bbSLhjpKm4PaKTvQNNZjbIEnnPe4x/xG/Mv7bSQylCrsfiQIB6hT
RdvHitXO+DanBJ5HdkH0nXcgq9hiso2v91EgjDV1BWJoLaIALrmLynJ7h6bC5qu5QfOxxwOKSZ9F
5ceZqLVBpqBgimwNlVxDZu4kPBZuvw9wU/OV9kJQ5/C4Dn/EONsy8rhhrcxTbkMhktTfG0tzPDuP
NvIKUofvQJXq9bicRs8l8djEMHPkB8vDqKesbQtwUhEoUich1H7xzwxBNLgy3xA3UJNfWaYnCTtY
JAvkEtnjZSxgIdwICwCHx5dLTHgdQrzhIc+xRFuKYVx22Obo67JlgyjDAmhqP4/FpRRp9mLO7PK5
ozrkozO95KuFnbvyLwC74sY88weC7pv7vYjWVfUKYW1PbDQSbImeZY5NGDfipPXSwqyk9lNv0BG7
Jm0WhtJ8J7CeBwooaJZHIDnuHcThNqAHna3dR970Cok7hJt1qJUj9Ic44EUSmXyNT7IkXT0lTRtU
UQWDGBt/j8yL3AFOd/KDD2E8rDBqNnESrF4S111P72kwpUFiNqyrjrwTCT9o30qnQsF8vTThVWwB
lpNGMzEZUkpIXptCnpQjiX0X98AYDiIeEUTD4J/vrxuBaLLnkyYFT5F70boj3C8aly96VPlPs4M1
naBQxqMOANwWms6hXwA/HMTZP4a2jjR7zDQ0gboAIL/jLLSe0Lm4XV3zSSd4PxRC+ehbl5pt5mEF
26SPRMtrK/g7z01+OtfGqaRxrOJn5oFW666TcqaO9hEtNx/jCxi05rJ79OBd414j92FJV3MukBUH
4vv1jZSoTj9v7D/V6TJkfykDVfK+xnUO6U6S8RNUUh+f0TkSez93NDhAfz1sEIMFb47/6b43ezQr
AqxGsQ2EIx4w/YM7WExH6d0bwKLGdZcOXt7GijkpyCUtLNy/KtU7p6gD1Qw75sH0KUQ3l5rmTP2t
G0OT4LHCgWqcLoJ84h0rdFakJM4uikWphAWbpyGZt/X5Lxx+KacSZrkgkudqSI+K66c6Cu7JB/5M
+4xDgN+35Ssp/5jss1VQtS5WyJG0H2GGqZwRHETOe0h7ppmdRyjhltfF1g58XuyRdV2Aqa85cfiX
1+793xJRsCWpiEAmSQBXqUUx2eRL9rM0zoV5zl5J3xbuvEqkWT2ZxtpjpIqu3FPsTLVHqfTBInud
FG/ZD+mpSxkHW0akvE/dYxBQ9g+WGKLsB6Z+6niBEJxJw09PXSfyn0htyLLj64UCCqT3T2nn0ooJ
4AfD8dD/wXn0tZkjXAzrtfQR+beO3VOxshpbvnbdXeBsmdSIL2yLHiNEedt0EIyY3MDTUaWSie2H
C1iIG9DDeaQa+XgDHX+eMq0CW2YttvR9uSAOkwqUHGhS7DJKpI+m73A2qBz0TENvoX6il7qDy9dz
Ig7SSVepVQpqWhsF+H1dWpWxo5883vwOZSaJMzMFVmyDoTETtnARM9oqdGN/TtNyopAzCURDaoKO
hI74rewPnfMWz1E6KQLR1z9F5waHk54i6pU9c4fKy7N+uoHLSR3BtmLTZpbQrNoaH9YZ5314U4hw
OCvhBXfOUPPgjXwJb6UNBg/lQ1/G7oundC8Kl+qpiJYvvEOBUN3TjPr3kTSzgxxQHYe34FZ78mdO
bhIqc9i4wbIokOEXvbJRDwrrXEAwOtw7YMhzraSVjcm3otnljWkSmpyjQh4i2xozzR7VvNukyDRm
xgUvtGDdWwi1XmjqSqdl9dCiD3to0F08JoIBgktTUQXUTpxJ3jXBkUvHI7/44u9xQ1jYVr81bHEn
M+OTWJwpT3XHCU2r/908Azbw1y9ZanX1jWSz4xeqfjzHtTbvsXV/+vJYYu+Q7U6zv9z/N023naeS
wyUDEtyKS8FK6SCXqwRFZ8unPmX9JE8/pUj8jFo03MB+XPdJG30+gRx7tp/sOgP0jTP4Z1hanpJv
uhGi9OvyZR2ht/NRXGW+d3ZOfC72dqVhFIId5B2NKKN/TbhbpSEYNYeGnS9KSG695S7TTPDuEjip
aqOFZT4UxDMvCa8SpozS6DrYQXXlZ1Et09q4mH2F1M/YVEACKW1mNq+fOwPYc45afTKGQrHjCi6K
27iabfNPkf7JcLEikIQrywm2VPv9MROMbIKB9XtmOksmKr9Go4sdiHUYjW0oQjer9WMsbt7Uf2Vk
VBMbAlSS1BEwiTVUjcqdI2k9//0Wxj5PnUMeZYtHlxRvqBNQRB4LRpcmCIuZIF2eECTSljaEWTGd
RPauBlpCS/RweeWoYrVO97lsmVqm6j7Yfr4TUQAvDECSH73ZbUS7qskUcVyEO8YxkQQ/Pblkt9T+
qQUhkmLLQlMeUUECn6rpYsuXKVMN/hfzHJyZZm12SyNOmFPxoUUkTRfY6dEMBHVV+j8/P/oGJzDp
6xKM3Aq3icvv47kVIwrGZlRYy6nIPfQ73fAuDCone6MVrzW7SVzumNi+h9nRMCqfh+u/iVfE/eoJ
DbuUPFQrWcPTVazbCn73AzyEVorYs84wS+rkQpYgBYpt3+y9xWkUy2XrOf2anDl7t9EX2w1ZbuEO
3j7DAcMFLuF/WNkong0MxPhY6Ko3AEHU+F7pUzN9dJ0d3s7D/QHIWy86AlQu+rQBdSSHjQPduYq2
vZCgXUZ7FAVjhAk3VZk+OGA+yXPm7t/tKcKpgu0SWjDelweBPURGK91OWFwzse2xrpW9rBUs2GLy
6uUUVaw3DrKFKQhEZtnT+YDOUa4lC8fyYvRsJIqqLzSamdy93nkQjfKUtVJUbcpRAENJBLwvYCsS
L9Pjohh+2SvXSxAGyDCbui/K4kCWvbrXHwLzaiW1xCoTY3Vej6xwP5/q1uU8Fd1xsgbFrkDevMJQ
rvC9u+TqrKVAuDXo1slfSr5GfmzvPDcUVs0sMMlDOY6+vWbMo+ag1X9qAkRXlD6/OAxfgbIqJDdz
+v5169VWpeliGjRvPfnbaPL1KLd12aPqj+JiJDSdOu2kS3IFWICjL2ia3/dupnsS6pyuEgTfC9y2
0ynqqzWEf7MATOEpmR/rCUJ/dtqTNZfoesJiV0GPaM8y3ikX9Lbs7Jrl47BauXm0PFNswaw/RWrm
6NKskXe2FNx2eRWUbcBAoO095cESBOjsodUeOn2MrRFHgGPtUB4QUDNeU5jOr+DbwD73TyHWw+Ke
hYBS4BqNxB5dgKHDNHGzkIhbaH8nGRSG3mOGwPaVk6ucKttCgWOvhbWpenC1pJGb8DO1xvKEeNSe
nA9Z8HuR1DG1XNrs81/OxJuLiqAOjeWRy6aCiPAT3iRFNKQeMQsKsADNCMufiA3JK7gqvLcXEBpY
SQ8KECRRWkJ989Yg1E7APYGQ4w6u7hLol/tKYMvz9S05zfPr7btma5U0lvTTQ9dFUn801W5R1Phv
abnR6LAyGkoFBs9V/eFzlrsQ0Wp7ldPRLl7P9YxMVO4460avdwxQKTn5GgyQfznB11QUD8pDm4gi
ld1oaiUmmyEx0RHdpsB5DWPeKf7qavv5AZn4BDbBYrCL2nyIIyx+14WdSR83QqA1P9uTB3TrNFIb
Wu/WzY/L1B4Iy6olXNM9SdIFuvLRYR4pnf6apQU7zvlV0O0p3tN1C2LwD6QVj5hTjGtishyiDb4c
DYDABQHs+MX6WjfFBKrBinQcxJbZe9Dn7SbBT4W0Gyexb7bhuaHxNkkovW2by8ZUirEQQs43+jzv
x/zGa/ch43IgP/GzywS79TryD1e1Jym/AoRfV08YaoDoc0VUGqbWUuPN+8qxSY4tFf0X/dvJfykU
amsEm2j1kKr1fRuaydrc2ZiJb+yzVVDXkZPE55S9ZZMtiAnWMOxj/MkHnOahjKgGqS4IC19d9Ai8
q+aNn38IsjHq8XeLDV4sMkIQIxUszTmY+f/8y9DayGonlCSifpBRxSd64jYu9bweiC+Y/NHB5Cu0
VhXFJvdIWcM12cKLkj9PURm47r6XKuf/tB44an3tt5h95l16G9Lu4xJohfti1iOlQkkJpyTu/plU
G11d//1J3HJTXlxhdujr2WcVjTzRFGhC9fn1AoUB5/O7fhXJxmOedxqeguNQulhZXV/Yej5lzPiD
ZIcaImD1CqnwDnupM8l5k5xEQWYwFG4CxYvWGYFwKaWii4O+aT12OJZGMiB652pVvpXzPTkP94FT
EVLsVLnMybogUXdTrLc51sgahAXpvm/Xm1YiyhMdmxylj0+V6tNBMJEzO26t6wQSGXUB0wA89Mk6
9ixgAKRLtfw5AcbARYuVG/kwRNto4rGyLR957AdIAN1ktfXJAw4QhUjThBxpqm3fuXbp21x7jDYB
0LAvS03i5LjUhONcuCPcK2b7W8f/YS83zTDGjDEBijYS7k07zmEksmzqzu/jRsoB88j/RiZhTIfc
LAi0UxXqiDkL1z302RejJ7KY26WerBh1winipSeek5Ujg55JvCqy+2iQVvfNIl4uuHCq9eJdE4cn
Dcx32pmy34j3kcNjtqM8P4vvDjdHPnrG+nDVlbd5U77UF6W8BKsqsohU4QRVixdyCfcupZQSTuxF
DHYo/O+i7CI4XfurjzLNqsnzFYmJM0uGW3cpuT5BhBJFPfboMDB5q0GyPm3vH4NPRbTCGiNTB4cK
9FC/IfM0C4kyi4z8b5LOqrct9CBOgEXxSaI5og2qDvi5pHA7S+1T9hAAtHIVhmIk1l8BlkgW1Bz1
RbNT0PXdVy/AWOpaUhADOQynlE4OJdXOv0DF/dirdO+b2fFUBgzGvjwE7Eqns/sjDH+YHKmQsFcL
HUNQ3qOWB5HE53Gkhi+Be+lchsaODdadqthDUg142So/KZyZcDKWKM/V9oglj7cOXSOvL/K/Rnga
X3/RFq9nO/BEv6FxTAKY5E/h+8AaMQSg9CvR6Fy3AQQupPRC9Nx+wRN71PEeNp7Db3PvOm9c7P+W
NsZY8zssnyB2pTeZHBr4WPMEocTc9BNM5cpqhfSmeJtEOtvWG2M/2GcUdFPGMumResBmPg71fWKB
rih6vxn1B6b3WKaaUl4g02QwdD3dc+U6KhfHyKnZ6AeyXxCkDXaJFS5Ge+m8kDA0vm96Bc5SUVp0
G/PAWsa3jHJL1fDa244JPqzgFsYDxXRknZqp5YxFa0GC6p+t/H4U4KdrXQ8x3FC11BO+yJEGBv4T
v3Wu0ipzVIN1L/cg8PJqyhmwERMxub9qBI3nbaxFzDOMrJrJNc5neT4DcDRSlwexrtNtSYFBJ6Rp
afHbTjgu+K2kB/7aFsyDaXKjytEQwa/CxumvTUZ5EMc8UY+Yfj0BsmFhUvutGEkrckyviScYzIDZ
lAhfPP+I721LfdNICvKXprlt+HCpa9lA8wRWGCEMYYHSIeRpWtrZMvkz8EOG/DcWogCDGOBc0mQx
QOLnHToiq7bL5iQobmyZ68DQzGbApKDYZtBFvnoPd1B51O83Kz5IcynuX1f0W8pUd9OrY47ZxjE0
o57DznJjCkdlISVXMzy4qyChi/PV45tKs01eFYoXG9S3QWRx8SoBC8aPclXMdnIT7dWgqWRyJvfs
7d5hJmJYsKHabi3l6sFvgu8X2Y7eja1wStAyq0FMQXcz15KhLnYFVE1u9OJNF92fhlO6H9ygsg0j
G39iyqyVSlMsLkoC7XTJNaH9XeVCOFGzgRcWa5rbJRrsR8TqfpGnIVwPzQIj7PLB1ANPUdmFTHnC
H6qMimSFEUzeosKeebgHg3f5FXn5hgdJs9FJgxEudqbYxqIpvnLG+t3TYR6oT3zehik8lCSHWU10
UcWo3vzGEmiQIetJBTODxofuN7iz3vIbu/syIGcbGQCUgqWhH9gfnxfP6O/30kQRofopbdOUlg62
7XroXLhPgCFgJCohsGiynHPEUIpYR9hKtFsUypF42IUvl2KScMpwSkXXr3R4NXqL2+3YqZD9nS4d
7rwkcu+7qnKH72NpE8/8kHKha+Hogsmmpr5ojbG9Dme1e/SubHod3wIq1GR5nIUWwbVk2PbOj1n3
4KsSsv4HkJBOBEywZ2GcQvDei2w0l+922PzVgnam4qAWAqyNjFUYhVh1nKD/z3ZMpnIVXVGmRFcS
kbNnTGwRTNQ87fBjNu1x5V7o28OoXBxToDgJ20RAVX3UGC3r1Vuu/xReG92zrwAKp975VXiDp87Y
BkqMigLJeAgD6FyoTWfBwE/EWoHXBTAt6q/gjqGBcLgVgrbfg628gcTWdCSVDinPXeHI3N4B7sGt
yUICjIGyA3YpvXD5+W61Og0J2Lq7e9vCOIEbCLRot3voqwfFHxujTZBLrQos0rSpjgPjUUxycp+m
rPOoBESr31qdP24raO6wJrzZycVcb2uDzadfouJSZwWVyJlNUFWSPW84otwWwL/L5OSSYDFwu2Wq
G4k10e5EFjNl9HQ0V+Te9t3aBYJlLP4G2hP7vPv8DRKtVmlg/pevV3jesv6cVxgCTuFY4NJbfHrC
Zr5+zOCBwOrM0nNYqc9qomC9K61yv0i6gHhLIUsQowWboOlqiI03uqy3IXZPJtXHjdms+Ni1yzh5
89OvFN4phD/VIc2+71HXtNQpzzj4G/poQfrr8OgzqaaM6hbj+X0qdJblApzrR+9G2ZEzqZygQF1z
QZMvRkq8lXk1bFaDSJrudzHPshIFpC7TME3uZc4T2T485+09AkHxmd3FRj4GIUOsE++/YAfhHBb8
n7kOw+1KsYjW7GjT2U3v+f5/fUUSeqSpfdb4z54CTpqx/l26r8QwohwBLVbgTomN49J2BOGgtVr4
584X0UdtH7aLVPg3tF9XqDUuDSRLP9xso7zGAl8ke59pB2Fro9Hlxd3Tsqk9Z1W2cJ/TtpPD8k0W
i/0wnkxB55Pu9ug4/zwWCw8TroXNCFZgHfsMfLSz3jTQVxg7IrgoyCjKfTC34a5Dcmp9r/22skbc
0kI1GaT/vDsMOwA5VHqxWZWmXD2mrwYD5XauETbvI3k0VNDgCxx/VrWufKP5WckEoieJg0ChHm8d
eOToXbkj+D8/8kdSyKLRmYb9/65rkLCUmKhLAkh5MXW3Wtx0jPxAx/GqgtjvgsPsZmyttWToOfFL
qc1yVHN05hycSJWELk3Nol2zN/fdfNhMcJCsSsKz+eBUdV/bLFvs2a7RF7AWi+3QsgIWAwiL5z06
GcvfXWl2Y3tbizlbs/JlTNHDBr5o14YaKnxnKC75uQsiQt9otAWXsb/hN+V/YEa62NfjU4C9Y5oq
6Xoy1p/5xCX5Q9oB+N3Nr1JtwEMtsdD6CT7W2setP0nOSpcqDV7cscAtHDRM77CygBQgUWwPgl+u
SpAcE6pRURjRKy5fGB9/rhSYwJylGilz8Jbf84GVEtHhjnhWdF/5BorJ0S7vv5R9aiSyTv9gjztZ
XgLYShynPZf4RfTx0/s3ErnPmFwX0eGpcznf7vcNmVCA3MiHPiNlmesiN6elKpOg2ZRcbnm4PLgV
ftLoJ7dqzoYygIWMSCadpvpoihU/xH9UHC7qXg+T+HULa+PHgSUEyfcGPyT4NloB+rLoPLb+EURs
GUKrO1BLBPVhNRKk885QXXipi55VmDD9xywQ9w32txGcqe8gpY9DEY0924HwoqmgRtm5ieEjAbpg
b+6EOnzNeRFg9NGPW77CcaybYonYbjsJV5/Uwb4cWHgr7WpiDOENMB+kmEDDDYhmzsQK1S/JsXrW
mBwxEyWVKgtRWVBgZm5DnKzkhhAceEpe/jjTYOMq+GvDumUAj7gzXfTG0Itjicbr3R7YD/geahrK
DVYxLRL411UFxtN9EEHmq2Kac55uaqHaaOFqtu2iXcHkXor8km0vtBzvkfHIJ97z6cPh6fiyg3no
/TCWf8y0ufscqjRhzZI1gSHS2uYuCYsekHvLlx36oOCd3Lt2S5xLGosEOwCWkG3vISLylAajeUhO
YIrvBO19vaLSwkbfPuNHNLJKcLKTLnCgGpi4pyw8xA2NoPmpuG0B8OS7Db1aD5XsyCOCQ2HEWVF/
oeZjXcC3EGTMgjuRcYjzXN0PRe8Frs+vsy+DZeIUpl3AaWymt0+ZbHhrazsKXoowDEciTERqCFOv
LE+wXM5B/8FF9S4kqBbLNVA1lVFdzoM1JK0DJlDMxZ+7hxMYLA+Ez24qKqUVHFYgiLhQd2mqCCc5
l079PbzM5raV2R0vcPFa5Gi9nFr9V/pJpf9Evsidn87nuMht70vSRtaKeRrLSOx+vT7EFSgSq372
xY1QPV56qC/Gg/RBMHGBrcLYy6oW6SW154jK0+mZP+pDY+Wf+e3SLKEqOui/MDT3xVKYiI7s7ocs
uVFJX0fBOJVQa1llxyfeT3A0C8DS7MjcaeAsuZYHfqJcUnDJ+rWvEGJH84k5OVfmWvhe0VXqfrJN
g1UETEIIVB59YGCHPc7kzUN9Jzt7S74GeVIVyE2qt43oq/Ut+k1XkKWlmjD/sYYtkwG1cIh3wngj
vZ7rDI0m3LRNxsSg00mr2pve0qHSqAA7YV0y9O237IsSVQa+C4N7/PfY0UF+7ZsvK8fGZZR1kF8H
lH0Wgx9+x7U3NKuY8XnEdDnOCFhfx4oDwXIoD7bOvAR/JnQ+W5uFrzzGwCgMhaYRcJzRuROv6hxF
Ji7/HzQYMFQARzqSeNL+kKaUT+w5KPtVxu/url0LSU9HM+SjpMEsy8NeI5JfZJxjGK8UtrAeihRo
zdTb/1xbU2EHbclQIH9nH6ejVudMmtFbI1xAl+nBunl+7L56R38aqEPBhkB61tr5uQMrQajzbK/l
C8e8pMoBJp+BDWLgwvy9WWRx4S1bG0bNIzQMksoV3PoZbPBOB6PLBSVzcjCTiPKnxTFG0Tfr2sdA
g4Sc/J8lsHjtj8zPImiRaai1Oij+vKXe8OTksQ53eXU8sBVLJILof2dvyBKZk/xKBrqnWYhgOvon
jxPDWPuppYzh8lYmr8LFUWQHKVQ8ZBaHFIG97mtC1VEFCa/fvUP2stSUWWB+nzVMpwGx3xAW9ssV
5JuHZy7OYvR9+XLK9CuDKwqHGFwZ2E/5naoxQoXlQfU3oVMiAR1PROdspY2nnmxFs84XKXmVViIQ
oBW5UHw/encg+mbBdlCviIfXABO6BDuzJibpA7Qv/U5JXSNj+INLggmNPqsteoiiZ6tjE0+0zzNE
oKQ4abksApvnHWSZWpIl0D5RiCLt0IG5B9I/yuU03rXY7uEOIYq1VR414as3qPtQJaWTVvCym0ND
4MsSnnyuFzsePNzJLOeO+XllDUeJT26GS4VRByBJRbvKwdzZo92wRnXwksKrXvod84Zk5+wslPli
Y1tZnK+OGW7cyg0J0EpydiZKrjf1qp3zhhkrOz5EUj5CC8q+0VskbmpdhUGWBXz6IbJ6yYUiZmT5
goURxYkXv7dBLzW3mi8RWlXsMBtH5eGRQDa4hduhbFd3oDEVjY9rSCrDz59QeJdhbJvXJepW1Zvg
q9EXW4OOeKdno+iLIugK0prWRtxnZs7COnovU85QYkiZKBlurI1xcSWQmY0pyLYPfB1qB5xYWZ5v
shH6tRb+ONxoJLXBVXMQoBNRoybp3pRHx26BNxgPEaEAQ0gi78GukPOiOXMFAJxlUVj1SM+7gaqf
sr+JB/XxcrlZQQKUWfnAttJFGhxyLDZqsf+spZDrbnfa2iQTDlLUXy3FTHxynmHEVEqX9oG6UzI4
hZj/3jZwu4YZ3HrnjjEm0IQ0U+Pr7LQra3e1bSV63LohwmVwvEp3/1orNkmWaixJ8wfSPauKAGlr
fKA75oZ0NoSHjRUUZxrDDBggI0tr3VkID2dLrpReKQf9kzn0rHcu8ML2WvxZfU+brNyFLzhxNVhO
2inLjdvBPDKrQIRxtG93FA2AgvAq3dn8U1+tk8gkxL5UFtyoSQG9WELkccXXeOKPrfBKSA/XwxfU
SgbeK4QvalCDK09sllSQEHQWtA65Xpwt6wQqGTfHDJ0CHmca7LLqU6+2SpHTpbx5Idb+YR+FUpX/
0wwFJWlpiLF5DtBAttIDmbj7HhZhYHrJwktSTkFrOW2RU9lsuJy6xbYmlZsdekiNf4hMJoaPMYfz
AYv/6dzb2Fmf3KYsoTkqRMAoTyJ/yBR7dEw757SMxKjXoLXf5JIN5V5VS0kmuX/5WcPWzs83TWjx
ZQQgMJiRsMxFddpEGZxYjoBZ55zw6jdg2Ws8LOfmffFS4slpf+5055ziytE6UVUGQDKiEjXWfKeM
56w4xTIlj+8BAI/X/Y7wPaazvIP+UWTBAaaKHoCGNBIJDk35JEDcsUywtskIynAMtbLSFUaRkP2h
GN3xecRxjbzHmMk6op11YmVTBH5u0RpN69G82aEeeSR6WeLl2VJ3tHQ5CC/DNFmsrCC3lmz30yW+
zJeftuyPNwM9g961OQmykd7lJGMx0q9mnXiJ+LA06AJxZ8wL86AZTN2qmiC8XTFJzZoxOydJKaIs
swQXIV2PHR6z8/D6/kJlDzJtB42Cu/n9PsupzG4pMVq88vxZtSIczlFPTBoE8eMqH4Fpqlo+rHOG
ohq6QAmuVHuhHVomUc3/biSQEENIn5UKG/DGUKx+TUDWQlTcqBbkGucyxvyB6vCV35jS6EH4TK9U
pSBwNyOUsAjFXtbZiikBiWtAhPKHhWnjqkxJa7W88HaYwGvQNUbjVL3P9iFJycxAEQbr2MnWIsbr
YFbnKoVih7Lyu/OhJ6l220lMfITYlgxsVdyizZIkvNfk4QQB9dIz44ytAtOT6HSEPiu3R6Nf93AS
09ANOhkovFeuSDu/O6czBglSxtjZNc4my4u8BTXE4lcqkADedEIjUdchoShVMfQ0MCdA2gCG3Eg6
vTDy72jJtRZbgL4L/x+hNPGkUWGho/iwRrfdLwKXtRl61OYCBWtC5gpj6qaO3ih97le5zd6xkcou
nFTo+mb1D3v177/zgbAOtNcQec9bSwRCVO8shZvfYe9lVtP27XxW13rI1hjcX5qRH0UOvwAA/1VU
w5pdiCvpDw1+fghPbnn3ztyU7Eo8EVLa906UDRK0+zgLbGYoeV+i8b/3lsRCPp5/OVYlQmHZ0WYz
GW8l2f+KWceupFee9/MMSgXM1gfHo6J45ibTOXO45S6ZnXO9lnCccv/WfGHggqjuAjj7mY5vBmwF
QvlLkSRgUEDqpMb4DjFJdAEGbpSaSvR81nvbnjTJG7LMo88DuH/zMrTk0W/jH1P3nSgiBJwvuuqq
gDXaQQ+IgR666s4Yqsrj5Ms3DTQIhEJ+aXV/fe8b4r2Hv+DUGWfr1291WWLsmfI4WnbwM+BVo7Tk
SmCpSuBJsNI/B7koDhBtFTRvSgVGll8xktGmtWHvWL6kv3Fi17Gar23zbkQGSa5eH/XO0vIUz5N3
duS8L/PNvqKELCKb+lXuLAQajR/H1R9tYXvQuiB1psAZDCKDNp8M6Mg5YTL13iUYJhTXyYcstAuJ
uiLVmKNtvq5YDbBwwisijNp6IwQ4xuOq1aJJKF8blR4+5XPIvnJ5jnW4XmnjHh3OIrT8hL9ZDqTy
zy9169G5A3H5g87scBRkU2NVqfPEtzSna9/jo6MigvG2NR8qpyr+UYyAqSaO53YzzsLi4kPkw6xs
Ch93w+ub42CCapdf0p7ulqVMCi7SNaB+zjLGzGH82LYzEeswO4pT4lrb4ufi65ziQ1JakBvqsJT2
gn2Kk8oy9rTmZPZ54fd1OfafuU42Oafi8eNRiOBBgrtsD6lIzyQi8XRFRFTpXbL84/YZQzGi6N87
RX9kZliD9lyIzVQBuIKJIQQmXSdRezlJZlRDwxGK4kqSu/DVO4kLEO2x52htxpqpTZOxnJJ0ZGhC
uNkNHxfAv8ykJlBfMYgr7GHKzcbdDeLAEQCGIkuDp9ROi5wb85DiuKgTtugUdJZUSN7vXBvcF22E
XxATTDrN2PnmAikg8jzhBFAQNKNLFR8fjh6cju6YP85Kpkgc9P5WRFCx3y9xbGCkSfl2fn9+uuJx
RchXjpjpMYsQ6ymusoTt06sbTcepT7yJZKzQTWw/jlwlX94ZwgpObICI+g6jb90ytEiY3IeK6F8f
c7fU/Hd3GTbxRUbU9KYG02E8FZHLNH/FRVgoP0KVI48f5c64J8UySf+CouynJJop0uYUAUj/xCvj
TdHXRSL/HBNBG8lQM6opqRpPBp6KM2SLgoVSxItIjkdtKUEqbmn5RkD1uWQUjZYDVmip2Z95BVi/
HRMDyLpHY7+1+/UJ5c3AYY17Bx8q9zx3wDa8c/kOjxditDAcgdPkcNfE91cpQma5XcK566nDO5lu
xx60InYMOMB8Ct94icnhookTqisgfwqWAuDSAfO5MK5OjjfLCn0cyn9w0GMV6ZQy/wQyOtmEg7Qs
SNhzw6dnphGhRsA4DQga3bFL3TljAUIOHmE9sRPyh+94A+CK+aBBq4hu1gtElvOuimMMEe3D6c95
xxuF6ydxTrFnepE3CUQyoZ9PSt6Y7WEzPU/mEOBSNXAWtMwyZXejG3kPgRWCLMVPw5bZVJ0EiWt+
WjXas6Aiy6y7Gs9sDs/APmQEHvzUeQjOkJ2dvVpFrVT5c0R54bXTkDPePdCVUg4jLHFXpXe8Qqzg
kj17ARw6jxEOve/+Lc+fRp1O4bYYt2I6twi9jOEIGqhI32Wy0Gy2BmK5Z9jUn2BoZb4i1zY2ETxA
77t9CcvbGQYtRhPGoQmfUv3eYV8DOIAheopZfimIUfhIQ3nf3WhEuJ/0ZMz1aTGYYNdUgyEyfTrF
BaKDjdPwDTfAb2RhLvxnX9Fhyb7tO0ojwmv6ZfjQSAFcJ4LFePpNOcuMMpO/bqZy2uzA+X82C5uK
6u0MJ58axQN1hnMRt1EB86tPmBAFNlAnmvWhYDDr88BjDOt5AJ27cdxZuT4eNjKaDE/d5Ltd+jor
AwoiavUzfhmFGghnXK/VI4OhFQxDNJJuXOdK/9FvXIVePvgc4yC0DWOW8w0uxJY45eK3OFoGNnB4
PP0TXv0X51FIXydScHomMPYYOAOQeTTQGP2NPHfdxZW99n7NNA1pKe6Per0Imr543rLbCNwreMRc
aB/2lFeMDgFf34hINLzEoeH7CCBZpHfidtPTUXGxxE1BCBxPjVj79qwOBvgoRdb6U2YRmGibtqWS
a3FE5IgCRTz4wvuF1Ct1x62vEF+XIq2XuyhGpZNyLJvmFZTToDLmCgsN4xiw6KTKE1lGVFu2uo1a
FWzafXKPfJoji93bnWrU2Nca9gNYNTWSK8hevP7d61u33blqSRd3gSnV8wkFXf3Y9cBRL6l3vy2G
g2Z8VdU/ifPSYC/wk3oFI7yN7/RW7u215n86HMQcuyag5Ian4zmL88BQQUOkPzlTa00EmzkkhbkI
eeIvUnOR/9v2iZxOaUHZ2tT1ZGU3JQwkAkn79FJFrJbQ/WJH+gQa9CHvsMScQdNZOD9qzg47g+eV
asIv1vKA9nTP6rf7CAI8gkxfC+kCIoDlDFxFWxEd/NYm+MQjy5QBMC2X1OddV3b4qMmTa69wQyfD
OMjNmu3jKsRmoBZCaH/+vg5D/N+p9Ah1FPOpmyUUV+istnpDel/hMZlK233blexRUMb79q8bvNZk
T5uL7Tx2sYgBuHPyXAaRUbfrea8C9U4Q1vE6rsArk56eGfTciqMYsQl8mDOo/mxAnTnihEdZcnqs
QY/B/VYBza+9G07TW+k1YmRnIAzS0KZZweOywHgMq67CNZfU8Qd4fkcEnkc5+UfNdhhiD0DLn4cA
jOetWyw9nVSne9TaBDWgzo/recJFBjQFvM33M8lHAbSUwmiu/eOY4Ob4lY1PSBVcapPzXb5K2CmD
RgaH2Kwv/LEx2Qdaczkx2hNFDDNy7PMjElX5hllQeJtndPDE+h8txjIO2M3mMRJwcQOBjyvspLJY
hid/C1FJ0SR1Y76M35wZSlef+barjwXcdX1YVSaUlzsuGXP6ilLstKsENjInbV5iUuD8uEsXmW4J
pRZm5hRsj1rxWTTEddMx1IuB8g0UGEzyK3R5lzlcno8Mm9lxT4G/YYARV2VBeK8+gvivbFtni2jP
TrxGKMcyPLsrAwskyAxLZUXgNZjODDsNbNxTWxhwHEr+7NIwh/1kp+zuEzlAXu5tNemzE4s+N4n8
tukE2GjQZ/57WZg6li5lb596bVfRW65UPZacXAEaYcr/1kOTRNtOV0SqKU2sVnDqOE7X24Jt8/2D
TP/jzMH0SY0DU1/Bpp60tak0J5B5+8Hf+/WRQ6X+OhW4rIrsimlSazIIk5KPkZ3soIKMxPJjmS7M
4I0YOFj7xS7Jofzq14XYAgpCQBmty6yp/qiTpQFDrhw6oLVwHw43bH6SCH8QUJUGbt5Im8ExnGTU
uesaxfW3nA7TpdYT9ZCjOkX5HLnO+/HcRW3qJD+NyRkD/Ol9VJ2Qj29qZASlxzjh0K9U05Vp61zL
oU/mDkV2vVKpEcpL8KpbcPbMxZa9zrOC+mbg8rng9S/vfctggCGM7PBKFfFZHJo1V0gviFUaU9Wn
xaiJLVSTM0qbIBj7EntVbGIMM2urHkKKwo8Tof+G1VRIGfmZTBqo+ekeI+ITkdsb4H2hh9gd+RX8
6PxGh26TlLlIPFRFNOBRnmLWXluJqC4hGlpj+8soeiWQ6AiSJWXd/AUrSNnnuetPVQET0duyHR+O
hZ/KFScvGAqcAxt3ddtd8R5F0ZSHJz/5EAYSYX7VLvHWS6zD9PyU2U1x4qSCRbIUn/xyRBnBBsqF
oIXodCfSecEta+4ODKBO7bcdfmaxMBjh1BKpPuCN/yuuuaGMPXRqfu6vSf1UWpSgxiPFNXbA+4ug
Y53ojHYnEk8Q1S8kn6aXEdHWD/bojSaKSVXXteI4HyuVIQ2+glWbrql8EFy3DZmAkB1cdzoJRiLd
oGJnqAh0cnDDSKkQxOSdiXRZI9iw5e42txYUhDACR+LeaDodhblXQknNoh1x1Zt8wybWQrjv1zRj
bGKIkjDsI81YwOs56uC3bYY6aOyRTtCDIa0SIvTzM+0VFoRELqA62gVUm0sx8p8cMkpRwSG4XCoX
SNn5erzCAXOSG5C2VXmbBQ0ZS+fn181IOvtyadpFdhShz7TSWPhLg3DMDw2LhlqENldOHx9vVXAD
LFtjP9BM392evNLGbQYpFFnXwln2qFrb7Rjbo0vxZffpkWgSkKhjipgeHQhvAdvg2dM3ajVNXFnS
T+R4k8JGTakeJtawNf8XN6mEgvQr7PR/xXANG5oPuptAbzWszb24auOb6ulcJiJflIknlOuMgIaA
lpz8bQgQU9RF1zllems2m5mjv0L1hg9YNhALhwjh0Hof17Is1iVatAogA6IdlW9tR/iFCy+rMCNr
wOzEW5ycI+gYzWFVQuoQmf0irQiWAkF9pWVaox3vY5ReUi9/ySZOp+0sWkJjv3KGyIwhOE3ml5Ov
NpGLYHXMlnAfvjJCcBoPKc+ISVBNCwth5sezGzr0GaJv1FKcbthvc0QKD9UCtzU1o0xTQQLtpAd/
lKGIUW1W6PS0GJNohiPdMbKfbE/eLPQaNWX/oka9BerRtyzlD5bgbxjRln7urtaMvonZYs6kGRsP
vTzjL1neY2YyIFbK1bQl8iBRfcwQ8x/stJ6x5K5PKsdHUlavek6BePnxjT9tl6/Vx1qXG/qxPfMR
sXfvyrS+hOE5Z1L2YsHuzi6VP+1ja2H/BN4sUHntHdagodV7xCaHyYsmdYtvbTIAxzVq6qR7Lugq
Mua+IIgpCbJGk9jHl4lrHSBXQUEklOIlQCDyyE8MDe80e6ciba23FPetNr2YqzczzGNJA0wtAuZN
nFbYtf2s99+nN6vSex3cXY8aISkhT7WQGrTVYY9SLqrYAEAua6USyfC+gLv/lkJ4yOi0tIBes6Yy
LOT00zKUSLakhFpaT2uHz1SN0TQ1Oh6n60HzcbnkmqMjQI/fnJSmCApVZOMNVGNLdPonW0UtcJrg
eQBVaIplz2yx6EcTmpvO43T3o+clAo76+rFsdVmCO2rgQ/WTRuS5zMZZkrmRPfdH/pUE73SJUe1g
KlPQzCVtuyL1UBZh1RLVg7KFF0eH58Ovssm2Ofu5iOB5QTqvZGOzH4RNYAO6bFjGnGj7FtciuPsm
07vjGrV6mSAYFkB6cz5Zq1zfZJODOq4RsBkBI8IT9nHy+vSxKHANYS6DT1WHOGpg5R/8Y6E57FYF
Im2SGaBFbVG/GXqBlhznpQzwqLxiMs3pEP3+hLjLXVz6xJHooQPtiQHGMAdD06oj7w744jCPcMrN
HKRM3ZkjWy80sNiPX9dQPeXL+o/ikczYF4lyk85kw+e6YiUW9jdW8kws2eiBukr7cbQ6qqYySP5B
pBXnRI+Y9SEa69z5cGvrNWVqGhsT5fdIJVk/5HAM7DOYaBim6VVOVk+e61Q1FK0qhshW3uBy4jwW
RieKdnROVSKTpmCbYDG2qntTJbU85bTCaGP3ZAQkNn/MjZXuslWWuqknYiQ1hPn95caksh0tMfhV
CzCFqtO2mc0EcvMIwG53aaYSgYGH78yp7jApy3ch1AAA6FyUouvVHohVrrIQX02kSVkiomYgxEdw
bFjLE3tO6U3yeAIJKqNft0V0WubSdHgcpEGVjggxpn1FnV41iewfpgHigT0oL1GxW2CLhg6ZuD8S
X0zVHXKpJgwi79XunY/Chap3IfSSpFGeM/bKUK2rvOIlDZQHI29enXzVPCaHq4NTSk06uI8xIq7R
THK6MAJ1b21+M/29A/blbVdvHCsbHCKC9J91qS2tMo0ZpokzT+gj0u9KjsiyYs9gLGBKPzSV6/Rr
4+2mXPR/CdslwNNE0jV0NFzyufLcOc0DiLip0HuFxJ0I66t63dctrcpKYweGQtblBW7IzIFpxuBx
KEFvvpQHQg+4nvmgD/CJgzcRg4/iplVLtAj1BG2fOhxCgBxz8EAes4H3hy6BtKR2AC2MUoWVgAYD
ZHyW8alt/fm/hEzNStTTHm1x6ZyZxg/H0ut/W7NF5s4lP+xr382+s2XFeAQ3OjD8fbmN7cLPxe1t
A0zne1ePD/OtwQS02AgjYhksLbAPF+qf/1X0LaiCmx7IIcd2Ph/HIiwuhj0RjmFJVmQKE9lGE2jP
tWX0TGyMnvyxCKmbUprJbLg4RymagTrA90rN2i0jlg/V6GRyEoq8sQVEodYD5fajBMmLEbPnsFxx
+RQNj9ZpkJzskBWrzir3x/jYdbF8RCOwUCXs26FspKaT/wWTyUSKGbZQej73lMyEDNFuxP0TDmWC
cF7qTpgH8LS1XvvCIk5dq9Ajd123LC389v3zv1E1sW1clPaJoyJOTSe8ehTRBkdXKPsrRFEnozir
THXD2lL8GyVoM/3VFNSACdOjCHpd+12lj95YMJt5HMAhpEjFgkp6+Iy9mzqvfQlgrlbz9B+bNUA6
pY4/DySyuKtYoEWe29ljQlpun1OKVAu1jpc8DLM8mMY4Gt8b1+JW2DVBkrswGlCIVDIoy25Q9gDC
m9dYsXqWUXmc8dQ9NDx7yv8aUZjL6WjQ+ZvLv7ImFlfK4TzktxbAYSneUQuYZSMxkMPrTsG9ItKX
XRmvcTti1e2sq11yaEbOwkF2WmoSTMCTbHVkuZrpaEIsHA6fPFdCPFE1dl9kdYG5Yngaa0jFHki/
VnfgNKgI9+9p119smHwT5RnbDuqr2aGx8twRyuxBord8nphrUddIX0aPUYTrcLPo0dL2g7K3+GOn
+6OXZ+aMhVHfMx06MHkfrHlR3YVpDVuGnFO+jIUT7/K+EY7599+hj2wwh9gxZi8QqcuuAaycntNi
vYm6Hs9gDH86SQvBjJYVn+JTs6S63szwVKD3zdQmMGs8zdjYuMdKIUm7WT+vub3lv1fQbYGaZNDK
Rq+BipL6YAu9QGccw+++W+bfmIKtoKwZ26gH7G/4fRSFU5nOXXMrhGHe4xk8j7nQ7LTL0NsbjYpz
ry9R1emG8/pKF4t0QpiM58ZEXeiFB4+Njh/K2qa/pPmy9tgmWM1zVv8x7p0QqTFwQT18pFRbZqQJ
VFfdGIKR5qGtkKGrq+BkS1uk7/XvzTVAVj6kGY4cw/ProFn020eowFJV35FMf75vbnuhIiLSD2pi
/rC2UEQCxtvN+felo7uIZqK4UAHQOtqcb4Q5h8hwBxcVbQPxKe9n242o72aEVbewbVLTmxPN4A/v
l3CzQVCgHn9r7SLj1hGuMh8LDwwByIuvAeq0KqAOZOMafVok/9ESva73Y4wldbnWBxZjw7CTdIfi
bMu84qMVnxLY+LglSl0RK8v2h9BKOxCFJK4LH5lLHVBfV4TcAKlEjDgmT+92oWo8RiU+DHC5wuTm
F7cqAyE0YbX5aTYBSsVN4kUSZ8jBoMB3lLKQk/kQRpGMV2fzJaxjlzWBpzJ2+0lyX93y+zOKZK/C
Xq0qHMekFSuYz+o3s3eqq04FTD2ydw6cgEQrRzm6VaTXlPBQD2dObZgxZUzFwzN/PiA7lj0lGwCZ
xys3duxCvRMd0eAsf2rl1ctDuxECpW26hANvZ4fKsgnuO87dOyRrxDPTLUSQuN8dPkqslAJ2M05m
AToPJyAk0B46KjweuMfYDg8bx9LhKUxcjQGvyBgG/rudH9Qj9CakaRaG6MAi5mxUr5Nio5zE1cVV
Ox9G/Oa1+oilJAQKsCaOiPklWsc5GAmEzsG9320RrYEP46UJkwZhDqtnc8rjXN75cSsS+tcK51ei
yDem6Jr0lUjJh3sTLbmrQMM0xIeC9yHg55X/M1AJLccsaMSPvGn3MOCmJdkXDYwLFpiTUyoU8k+z
QjbqoRBqTLguXohAei0Y0V/BgMDQTUHP41dvkvKkIAWJKHgvTOmVTs0+lhpT/LB78Xm5cLScohKV
24a/Xyz/7KxRhnWsg3h/6QZPeeEl5lMs20jgko60NjErQodDeksZZv65aqots53GskpQcreb8vSv
7iUinVRWgMLHCV5unu6wOXkcR9SuAj12cO+917YslSB+iyfOBXnDcyULOPdql/MJup0IFjdqB3Sz
C0vb32F5regQX1dgKRX51yCRebOGeNe/EYeggxNE9JIPLhs7vbYR1bQNsVyv9SjUjdfjytmUnoWF
h8B3HqKir/pGB5h7oEshXQvj2PVtV/DLQBXXT37DUKOaqKEcfGtZ4PbeAFVcILJRuzdSPT5C8XAM
w+m1MzJfTyFVqCBPv4NCpPobMPe7IWCWD0KCkU1+7qLUJ6lEj445HCqaPQPXtsEi2afg5v49tZf3
l0t+8VCSTYA/7bpB3O2DGaS1kPhBOnWpid/dRQgniKmgSXtmpLPLA2l8sZW7vg0Vrs3fplPwdtji
zVyT1XVOV3h0nCHWaq6tH71lJMewEMF/LFJTCKCI8pecVRWH+u8q9Nzal6c/JINF8Te8HXPo0gmf
sMoZd++uVenm2NpS02PgJFD3YDyRIts3D52FiIUhx/h+JiZPnWqq33LV98WEyjkWz8JOiF1FtFoM
tC8Aee1eLX1tD/9SJUNto2lkgydK5qGiSizF351356Y2wA54dH+IGNBgR0GQZDvNKl6mmZDA7241
8tgWeGJTpPH1QbajqOagA637h8DoWQJKpv220U4rXKVlYmheoQU+tI4Zts9ITeAqNZWL5I224r/7
ydKHIVG0QpXK1murGKe7H/z7pDyh/3KYN3+Je4S+1qlZMuRKgUkHosE294pWN3DTBgWoHb2BYkz6
iDrxBozo22wy/4XiT2v2FdQpvEBxPhoY9M+rdR6Pqg72UpkPu2Qs9dA30j0zu0Ld2CUTwx39oq+P
boOk1BkJDJlld5LadoWY8+HZT3YYuFE4M80hsrGCEmvqGXYW//33voF+IGFzmcEVuy7XZoKSXYjj
XPOhDTue4GTx4iVw0qIsEcbrRoGwk3BxFTEvpFCzJSPlvrsm84tDsLvYdVcB89wPPAH8CUOmrAFi
HmG6GfHwYjTkwaToWUYfQIsiVwldnbZqRkfSPdgul4334DyyoJwM6tqd3H4MGswwht63gRjKPUD0
1AadicFRwC1erbibViTpHe5VkndKpiByuc0O2agIVKwbrCd5ZXqN4HgAkKNAoFg/Picdg82/bqVN
rNTEVKve47o0tu6VaoYFhKdQkTob4yFpbbqd+JTrNXgvJEH9J+xvLEshCe8croKipafLRx+jlrJ0
U5hbuvYn1eG6HKx+EctHbgtzH4H68YQnvT3Cgt+GeNEQ4617wbLtYYw5X017jvExqghzb3cXrTxy
1Bfd9EP+j4h/6aCud2R8fqvy4rGjFqxpoQ4z42SLTb8zJD9wsHfUticvG60Xit59R4N+7b1+K2T1
WNsCZg8pJL4PjXIWKYOea2b+hRqrQDFyYL0aHn/MeKXlUkB9EEZTu17kWquCC1kxmOBS1kXlT49y
VUGU+dHac37Y8CVS9MOJO4fyNY9zJ0v2qBOTj1wGLIPES/JhzaDFmFjcFh+JsBBQWPP+YxvnK0LP
DsP2y7z0osD8B7p7ZGyKIQcsQm+OWmTNp+SGpyhdVo8HGMhkFnbtfEBwH8hU6zXZPeA2BoqC9gq5
0gvfZk3e/pijJKrjUQKxFsgxZ7TrZqGIzMipg8CFoi08X3Pn6JdMO8M3cRqxxAhv+gEj2+WxFzC6
0hJs0Qdb4WzQW/iflnL3v8bKmFNRFURi1XHteDAyUOPwSfxbvVkcLj6SkQbjWk841yIkU52A6zhS
mZtQhkWx79zq3COOWmDtfww7YOt0yj/z/osMUoVjoii09Ag3TZvwBwpdCSCxYvDGEY3KENvFUfRp
ZsnnfYl1lN8HZEF6AVQ3TRknZxoyEvSNnf5YBgjLYgEUmfhsp9YEPyRKjPnP7l97IA03vLPEuYMV
P0CMI+f1qdzO5TMfDmEG231hEntNtfBoTfjRfuSw035DM8N07lKCjBkMNzJktjHRZWc2AaNSdo7I
FuhULesJpezwasgiXstMEY0idHzaCD5Uu+N598ZT9R7pxQlB+0EVF361LfZu6KrLSiG7ESdoR89w
3lvwAssU+kVyF11T8vPDtLVIO47UDAp/PHryF6W+Q9L3d/4Po4QKiOipz/zVFdHXV5sWQ3e1km44
0kU2/+ddHbYAY46zJHbMy2GZdMRsST20edi7yxXdJ9vTgR/znd7dihwOJVzYH8cIHnBFAsCWqYKX
2fxTAFTzUYjfc+Fm6mvaSITDSHGvS4pB2Dg3DipFk9QaQe6dGzpk6jEBOR7l9OT0X+HbkrtF1GVM
nWAF+do3mDEbpcP0LP6dSXjQwOvHCbo/oBlUMIbr3bgu9axnYxN9AtBfRwGbw1mKO4BwUP5BSYlE
e1ApgeKBZenld0zx2LKqN5X8xzonAaISAqs5dQwYN6N2XlIyzD3jLpLYvxlljGmah/0A6XcC3JAV
UHY6rHdkjtgtWQQCMU9w88XDbRTbZNYabGfgntqmLaiVls0P8I9/aVhAf+btYqHQxt7z6lnaYq93
fpnd1gRhKr6M+mzgkGjMk3JGQ3P7tGml93C8aL4Fc1+spmyPBEjw3Iq9gC/pdsoe+TFBPuH1yZfe
wUeR6MGA2oU+DM3GNdC+Ct3xnmfzBcVjv5fnR8bn5m93xouJwyBD2GZasOkvRrISSQYZR6fVWU5V
Sl8mBazp1cksHPIAPDOxGf8Eg3YkMy/znLn0jORTxxhDOuaYLps2O5y40UAckmuucLHQDBGHmZXG
vjLaFGLjcJsUkjw3/Mvkfk15ZNhQYGq7cK8wdbapbNdVVi7z/L9wDki1IsvD4gC+sGgiJUqi99hy
8Z0LiLX52GTUIO/d0c9OQdfPgnAKoMxwcaboKNFFlu46L/4v1dXuphepTChfddYd1MyRsO+g+m6L
KJrqguFhV4utvG76YQJdI7itOxJROP7P//wC/Kj32Y4XvXGhB42lAGhhMP8f1Dzayi/lwqqXw2Px
YmLg09Ig2n82OvtgZ4Pcmz7Y1M0zGpLaVumSHiL6WwdDfPqZJEnMTfaybPJJt+7479P/0wYZwT+U
rhr6HvzDr7xwW/Syutl1bNfXb0dU3SomrDfubGUmfjb2lk/RirmiUuLzjTI9EZoSYFEHjyeYIhxd
d5zELkdqaNQVnRBEaM6n/z5J/1lwvtBFD43MjrwzwMsWURpzSYoq9YoOQTUwTp26B+hA2kgLRXTY
SjV3jbASebTHYWWwEaF7yAHB/rYc0WirY6TChadCCWjeVqXIPvHL0ZAajS8Mz/6bp3tWeKJbl0YX
xY2NiXAGD8PBljpTaVm/nr2NtdP5hDL7zAv6e8ZxdIjFrwfXrXPBckW5k4qqhIEGO2WoeLpvuD/H
PP+JHVNArnyZ0aBD/tdQxDLs5nR2cMQg2FuTP6R9vSQ74RlOS+1tcwlubWzjYU/0yyPlWy4as4MN
5O4Titd9xOLQ3kBEX5zBLJFXqo29QAxOHnrxQz96ot1VCSOiRV4A8506Urro0VMwYuY5sfpChvmT
vZ/DlFd3ecgoWeDmC0rcjr4P7+l+1SH7w6uaEhh/MYP4ASa+2CDW8ONdRx3S7m04omq+eImIBILj
+191kSOB5zHFvCwdsfxsCqtAo7wmuHR0OJhVdTftZoNWRx6Opckv0F2kLKuubJwJrzgl4A9iTHeF
7cXgc3CRdp/EbNWJxUOJSLdrYpe2VFHcOpoYHmG9oNs/cQF6xCsjO2J8M8RxPRo6Ljxn6m/9VPCS
MbxoNiBexo1tcx4eEjn4yBvgXBvMk77KNmcVoU6dVfIQ1p+ObqwYIWO3hQZVMAuyAPwTD2+oCnOS
NnfhlGCH/35mtR6QwiXNMsQ77lx2btLv3THiidjxGZaXm80RczhKglu6UI8uDegDWMe18oaA0y6+
sa/uOX+cuopsRvFlVmcGcibc/OA/kkis6feBKFMAQXUfWXbMWhHR7Zz/3zKwxAbhNaLoN2az66G2
8QpYf7czkddvxQzoelBnTUWTHglRQGZ1J66BU5sEmR/9LuOcT5lPUExcVtpGTrc0DMvLwLWZgANO
pIsi7DE/ZQ+zhGO+7bS462obBZw6bM0ZyXL2/xHBBSDa3rhnz5j91jwje5lF0ukcFisf28P10Vh/
IDjodxV4xsItbJKFgUzTzAUumYAP8DeuYRZqSIuxLs8ZB3IbVt4gC0BL3k8cGetDcan0IXjbopEU
fru2xykoUvrl1IZ11eqczjnmTzTbJ/xWs7kWoKZxPlRDQOqO+wvah35VpJNMwCeViJlBy6cPiupK
QNQYaX1it5FtVDCcQAQKZQ1LJ+FPaiX+3evFYolwaknkQULsvIN3t7vmZcYJnIatAz8GQvo3/+Um
WhQKfuO5zFUfz5Yd+IOk/V6YIEJYHJR64UPh1+qDqv/f+oG2Z9XWubKcuGdK0R5h5IZiUomZz4uY
pL9DJZHuVfTMe7RzWqefdWz5rc0Q7mL+nU/VugAA8Sx+26Y7n9tEGImuI/hcID0TqGyYRzqw9J9s
0cNtwvC1tNsoOreoHTPtJWnzBwd3SFAITDDLMeOLMzOeDwWDzwTY2+14TukoQI0TNRhxCLHZA19x
p/BbpIIfDJUBfXYvuTpy3RRSWYnc1vhC+eXAHSvNjK4IMOU0sp2d7/jG+vi7gdosUqUEduwusrBt
PhcDI/kXPbEKHCT6nRzkbStnqA8v8sOrZfykMttuTVtBogSs7WFmG86ohbNO4+GPcUx998Pnjv9i
7xwdWtRMPm4WQj7E02gkNumtdB5HXZZDbu5y648Qbjf2bk5coOe3ZrqvpFlv+M+Qe/BDGpHFqG0C
VinPN8rU2lMbOfelhMyBD5QgZT8NFwzP5r3mWoLa8AorrGx8QfYk3whYXl7XNgI8u4zp2Jf+FpAQ
X07nmQVO0SxxGeExpNp5mt0WjfKoKvXcVpTAC3P9YDoERDN2N2e+0BsZQ8Ykzd+wFB0V+l5CSxlF
SUtcw8e4/4/2FydXAO7rzR/GMr60RC6h5FKPhvYJeGWBC2d4oe4CWaMhXWWuS4HctqEAK4eBNHaA
/W8zeE0cWYsTTE5YYpNbModlA2ZNF1ExVO7TxUuMNsABhXs/5x6HibraMcNfS2DlnWaoFq+HwBJ6
l8Oef2TPwmFlB7LKGAbqEQLBJHOV5NZ1890f8Z3/miIuP20cohpwJdYsg3et1GqJ17rPXH4tont8
YfURP8TP/5/8UARw8uwLAAGk/k4rKHZ3UbHKts3KNUd0oc8G2IKwUL8yRi5dj4WVhFFJjsbXzFwc
tUMILGiuCXh+oRfENSmgFHJvDjDgrAxifH9qgRSqo+TA5OUVHkz4yb1WOHlGqQlo7kra8JEUq7+Z
KWYrO3Qm26H8kUFaThdR5wZVLpT55/geNIzzFl3Lj1S8LT6ZxA5jHHArxT3QpD4eZQHqBfGHTPZu
VcNepemnV1EkXWgVdBQbXGehNFiqrsbHSvK/BI+uyX6NgYj4F44/Tdg5Y66c1Dms+1b3wowlFF20
8F+Eer1u5HUdGN2LbJ54Ef72scxDae8MTjMVSjJgs+n2dX0sqdh4xbqquOPsAYq2XrIcmKauiDNk
rjUmiMZvfWiHUNtBs9+h0n/KAvTyK2tjO5HYb1GgYKNfUi9CLY9d5PC6Jty3qwRf7/PU05KlGrBV
QxKBS3UvBVhoWRIeJCAupZKP8xGQRl15Oj2kiq7nHT2L+cWau87hKEN5FlrtkmhMpNxNkTkB43X1
lfCMfr1PHO86AaeOqKCvTlzft/W4ON0BdCcuZNBz9FitLKyb5vkyNziCyy8QTY5LfwjWeQ0x93jz
xAmXKq10p6h8TSyDd+FfR4maGVGEuOC6ufiun88+3Xl6GvQvc7+4W9iDmaGIdSuLRP55kNbY59cE
GLw3avzDGB7/sQd9ZParKgkCl+o85wF0rsTrkh5mRz08cqytOvfZGnjHSOG+PHomruuahlYetVNf
mYpFjESjyCuFico2dflH0Jowo+6RUQ1Eyoq+HFVjmCjDtFrok9QhdCW3Ljf3OgivTIGihsH4Ya7e
9gdmNj6OKOnV74BBFSA44S1MaBsfBPMtEDK17vs6MTW2sECgV3+7VSaevdhdaLlQCLZGvHUTxA62
8Hk7oy/p4hEErMX/yQ3Quq92w5aRfcGyx+lW8M6X/1XllQIX1USxPWBxQew0prxi0nu925MIIWE0
+6jG5wVZ/6/Uday0OKjvgkXfwx1wwFIfFS41AgNseJMG2gLNIztUkkuvmAXIb/FX5QyH1PH/3Coz
nf/aYZev0gNnhsK9+woaTA4JPfj3DpIDVcVyS6a/XkEahzjyLSJj6IbtrKN1xiqN8FMPk9iAqST0
OZyIuvetYVvDuz4qAC9zdwnPqg1iZME3GxeGnB8dxMIKy5K1WlX+20AvIkmXi0k/YIaPIkLHlulk
IjgZn0OIs6PSDP4qVl7kphIBARPwcaE8cUmffHscroJKwYd17N7pTzTya0VHyaAwrC70l7fNAEWW
YZ65A9PYVhohdKm+H+WIeEMWEVW3jK/LCmTKGCVtHTcMOLN+evy837dQ8AdVmImOhA0PXxkhKIZ2
1YW9UhBo/xoMCCrxioAqtLaYz936dESl0EikLeYhVnp3D/d4KCT+sKM3jj5hP6NKDxJNyCx5UU57
hEx2W+96clJZmKkLRRPuj85jBJqUp2yxUHh6+6KZr23PlC1WiNadP5dpvc7rh7qyoqOWptcx/pMS
883gHaMl5yBTqNG+EfeqQPdOwQitZRBGRzkWeKF/8H/EKhoCX0GpRQVTAUzlnnYvZQe8FmAK7Vn9
YB7YzW+ZCj4mCJ0mjSGEVyOKfGtxFZI+RPxd2acGirAjfjjMP0GOfR7YMSwbRUVkQzNVATevGzA/
VWAWq9wtJ2uZbEf3xzzH8I6SlCUG2e9KxVYY4Hn7sa95FccGi7fJitsEtC+4mFlKIXU0Sh6IHrqf
da/+WhVrqxK4beLAC7HnknosYY+eabUn2nzk52gV7zIP8CJOmiKMfXJ4C2o6OlkOz2qBPn8KkLBR
6gsFtTnx7TLhgza4kKbF8UocuK8YKdjK61Yy6fcOcHfPWMTsfgf5y3IaxU0/ZJsl0U/Bm6VgLqgN
wTw01vjiSk/qlzXjF/MAu9iH5ozRUZ8InsexAli+VYFtKO+t+18v0n/xiDNOK47RAsMtlYZgXQ/q
HD66Q62d2Yr4fE/pqmMJqMDGXGAX4jpe1VlfrzoAlRynmsget9/jTsUvZj1mBksWZGWdooP/EWRP
j+JIFiMfrb7XsT2LzOBnqsIlbja3/shpD2NpoKY095X5ONT+Ou4uc6kkXz0eXI4ZsK6nV6XUk9aq
gcbrl+sr9LVSLmmaVyz3ZoP6BAlBVHF9TPFzbjt0xt8jK2K4je/9iqJF4tJAxLiYZCxUppVfX5iN
KG3ry6PXBAG6d/4/FHnsbXt95hIOiamd/UdcYq3UboBXC4SjO/gV489kFlenssc34eMSMM2/Hj8e
FZVjmg3o7vxNA7Ovwan5BzGs8UP2xRnzMtAXHKH3+pF+xDH0zPBd9urgYII4WEkc+7OEaN39g2SZ
kJYEXDSruWKWH7mfR9489qDVgmz8+FfCQ6dWfbHNAWSAf7QmtBLmVrq2VXdkV2CPESrzOLlNIZcr
9Xc6beRubqhM4ZXo8QmG7lNFrO5XfGroYeMVXvYCs/T+IYEL+SIhj64piARKJnJjbdXMeZ+SFPr1
Feh88X26gmWZc0axWFj2fbmrIKqC1kQgl4ulWk7iApOR/aGiQptRbdUkM3iD8ykbqWNtXp8tagvV
XAqQ2M8yL0lYBheJG7PyxLnvlxc2u/7D6s+Z83fAW2C7d0AwuPo2SJNYpchjlQwbT7B49mHRoIUI
C5tPz4nfzMt/JXDq2x63pwUN3+M7WV32GP0vygMMHh+O5cu+93SXmumFawPI62ZX16xMGC47Io6Z
bCwp3uOqueyJrUETDdaDSS+zV/CgJ8fSgpWUZJpiY8756ItWwkgejmk6ZEsSwbZxwShs1gG8glu2
nfk+m4Tfj1jKhNixUPibG0U11YEdjeGpHa3AVb775omF3eWttbGqYAvpBkI7+VaV4/ZxIuYfJpOD
L7GI5z4ek+Vl1WDQ94WQeEmGoVKtQhVX8vzTvPzkd30hqQhwfFVvTjFYC7v4odVTFkON/jF9l6Hz
taTkaiHQZ53DnTs17qO108ArpnT1JNRy2MNzCJk5Rf3y8WDcTpB0eeCDRCAN4uBlJPseiX96t6Im
KWwfZEyOcjo87RYfE3PeS2n8KDGKGzHEPX2qJ2zXT78ydG2lmaP8Q8PMKmeYZxmZPr+Y7APj4fVD
d834SaUYjYtuQvlFpFS3uxW0K51IACjzslcmBtW1+WgoL11frXqgZwVWWZ+yH6TFxOD6/8D21oLB
M6iXXgiiRSxQRWcB6UNsILco83VNsOtNXYT/rxl0s0woT9bX7lfsks88TDFgdSSCC6jNDqYFhh7b
ziSd3HHgSo09B5agQmNNnaj2FnO/H3dX4XWWPj4TSMbohvIlLlYPi+JjUCOyOjRWZtyP/fgiIzJI
DZzC01cTZiLs4NR8FdXiXdMoH7lfaTgrUnSvtbSu3ExX9V9XPawQX6hPbKx9fC5GnCXyQT5y0rrA
bEQK2lHbW9eJa1JiLsdgyLL9IVoHlgtIzvsvpPJFOwHcsDW6u+l9PoPzt6Auqa2tCVzbqg3bVzhP
E+mCvy9ABT3/oJOxChMTy7cXmE/OlGfGDjBZyFgZpEteHNFw2mWJShZi7ANCKlbPz4G3EbixN9JW
uLQtm9fJ0MQigY4dIbsAD/hkbgoeT49jY7OBG2iSwoxaYEF8myWk96N/oVUavCHiZVFU/4PznU60
HbBxKG/yATMYu+M2RVgSdaIiP0SRGlO50QTJc+2vZjOS3JHbg+1TE3tMeOeyVS2LpePZfkfWHn+8
KDuzm4IEIeP5uQ+2gioNzKWSuqZmpe6LeqbKlkNdqtRgS5BldSCv8rJIRIpfFFD4u7/mARliY2on
zl2454U7BsTC19evdfb0uhNd5KKj+Ab1KqS7X09l9vytvlIxxxnRM/i+hZ21jZVa6phwZxYZizaw
NlFVlAc1Qf5GdkYFV/lLR0Z+hotiLj6UBtFintRRiEt2kL2K14iEDZMg3/zfYgbNPCUcQh6+m3G5
oZTupkV6Y17Ik4RkhsGzR2GUWfvXMfK6Bhfa3qOVKK8ZoPuvvZqLza7mbzoJoXsIILRAh1YpA7xY
QNcKg0zoLdrgyu+MaMrHK0E2AEC1ihRG30DDif0Tah8OUF+Kg8kzVz+mymFMuLaOLCOVgMnIZ+Rv
N3Ly3GvKjkyeobcQPyMnOiethGaPJjUTMhaSzCRxL+i8X3b1ogF74B8SwoAIC4vTI7pFEHPxyvbl
8ibbVeR4oycr5z61SzYoGeumJi7LTGwsKeIERvsLSQ39lQkO09NPUqch5BBZeoDjYlVVdNU1FEuL
ZSROWoF+6+Gg8ST/EBvtq0ghk5EPHE45t4vlJnemNYP9cT4+d+KgJwdf3yRD8kBqEwEFnjVAjI6V
OzzGGv7sTcTbShYWAkChFCNPl4uTfI42eC58/G06LeB1QUgn+S4EuNG8SQKaYHawvVbBsFuT8A71
qIIeafMBP1C0wnhZo3ht5/85m7QyC+OoxxB4L+fsdZa/VpTcdoXsGHpBWYJdxNALdyuBp7Rkn2fR
AbxIQz//6Q/Bfs1G3HAMR/B3Ynkr9knVTK4Qi6734VShRj+ysa+mok6a6BheJwlFH/K1+p4u3ED6
SMw5ThJoGssyr2Cn2xnlxj1MYbaMeJctpk/A96Hn+hroZERAjhxSCKYM9NOGM8fkd0mXmIvw9L3R
UBASY889geAS/96lRoDXxNLmeKudLokVOGrphdmngbpnnsSAmkP8fFRgbd+9SeHe+GPCzdK6hE9G
e+R1lUSiNfQKEpwpZwj+UYDoVAM8V6Y3HNsV4HERPu2khSW3r8rIsQNg+GtZ1A2srd5Vu5AorGkb
149YEofge+MQK+871oZjOsh7gLke5z2fozjPLVXo22za6QKU6gc3B53/nWkHv7aGSrgFgYAND+VM
4d1l/ViQNfNR5qIREepqDyB7XfCQqZjjsYifupDOJfFUpzWoknCAIOeVihroMlUCUkOPqd1HRqEK
KH0u6rQFZHzZHcxREDgfNPLlFJJ9xopO6OYAt75bC/XUuunhXy6d4XpP1BpQemcX5h8CALrFCjen
h+0Dh1Fr2AeRDRpFfBW3qM2h77uP+z/zjLCdy1ioX+T79qfeARX3g3b/ZNe6SSQr+jJTeP90WfDg
zfe/ZXrNEYKefNOO7deVGQoCUSnMHmczxFvfISYqo3gie4KJwqfBh1P0TwXZoOVngntqkVqh8WFz
sWKy3ExPA07wFBFS4LBLgjDAB3DtuQBzELPxK6sVWwk0hfqrmZUVh8dZlY20xIV7llJDh+Yoem7N
qKIiTvUHlUZnPoKDZuf9RMBlJvM/h6BZyDk5vsoFPRYRKODLom6WtCT/Vg6Q7LlvidhU4jE1Bm7D
xlGgqgGfUiumVUqxEaabF/n8/hczXTBU/wyNAmsGCUFwtlvrd9pNfs1U43yBqcZL0nehHGWpOMY/
cXvRSl1iS07eFJhXlKF2J4NSI0pf1P7Peb54XFH8DJjr3BU5Mv1oCxPqO4/ymSETW7O7StJjvJhW
ky/O9z5XhNPN0sGXIj5ErXB9WR5WBVYZB3nYj8ni+/Rw3IjSMm7CM7kFwga4I/4zDVl+R79cR8iU
gxLux3G/N2IYKrNg4yAbsNt0NEfPlK+THJgAOgOW83Jzvpkzzc9ydG7fgRCPHytOZWQYAtM9oUYx
C57TvLrEUsqGWlkNqb9gxhNSM3Wxynj4rPZZ+fAFGMV6CFEqx5oq6Ys6/GGIIaHx779MNnCfulNt
NG05BhQ7LHsu9leVIMLSLawsuGCw0+0j6hvfJh6lXXUOkD+xG7bEMTMUc90KRzs9jkPvCnseLV3i
RsNdjuofsfHFpS791ejB3UVs9mIH7IKSG7qZl6NjOEqBCE/kvYyPwHkXk6Lhzoz8jnUMKWU+nU+q
0zHtIl09ipVFG9ZE+mKcw3Tkx4A+RuM/yPJDPsH9XJIOrZQExf40iUdk54Z1QBXxRlJNwoEz8sqS
0Qe4bPmKBJJg9m7o7C+m1bl91qSF8g474vxt7eGYGB3cRp50wBAaFpHFYYl0ByRNnIEgkGlxPkJy
1qy65tTUFurcl7D4j2n1jn0HkfZ1thBlBsTfObKWLjrx1KXTWYk6kEq4FjnNan5ANp8kY2cUhISO
YRQA2ELyKB53MlHsFyti0WqqZPrCMcli/5L+GjR8JDv3e/9bmmNidO/u2WCaDyCiB3yXvG6Srltt
d9TxMUC1OzllquNRQ90AYOpEu2MtMP/uvpwejVk1OZe2MdXhi69uEaIuCZpyZ37onFp3QZaeL3Wh
KhzzgKJj2IUprj5YRLXaQTuSOXtu0X00FPRvGfuiLWuXXTv/uyfv7Jo2FV3SjuyF7opEg/Jkz32/
V0Wmqdbt4O5MEZA1rirfi68PWd5LJlzsVKr1Cwio9hijX8VzogdL3JDEnjfAXDLVXeVAzFq/HsGY
AhFZtDmdApaSnEl1vd43nVUOPUdVjZbPmd4C37c6phHCZct+UHmkULcZvK9t6gbD8omoYPJh0Xed
QxQ0xzD6km6nEhsK20WSACGGhSFzsEthfUY9C6J2I6lDVG/76AqX9LSIxRs6Jro4bPFdYhr7T/Wk
TJDY2+GpgD/e36E1oFLuO33ZL0vMI2nmiaufljsB8AJnxYhkhkuOhbSEZ5rkumB18lAkxIcWDNgc
1sHM94CQF+Z3XfSYgehPECkv4Ubr2bs6L1MVmPic0+5vzRfBNYzgVM5ejPEJSdTiVZf/6A+nPJ6w
F0XrtT0UetgC/bRY5GgXlFpR9KRFz7t5YSLjc8eoQk2QkE3rPiv92LawIBcuxzyvPSVUFWsEBYyR
+kEDR1hAw/TvhcAoqiX2fcwg1avpxFPeUOUBV1Pzou50zwf3+sYEdxhWJhl6MR2pgqzN/fxN2O60
pEYNKRf+nXaS/FioGpJfFLtjbhcbXbjE+jmIcmcTRJr2MEeW6ShHmOQIlOLFZ5CNup7cMIcwLA5S
Wv65ro69Dxb6I2vGGC81rNQuaBO1Ha4LtD7Z0XsqAwjd47TH0jtsWl/Q+rk70DSXp8J+o/eLG7wW
LMLm6OvUTjgXOzTQ5wcrXdjmoMaiO0ZmLdfH6U3hwJmWQs+emTzcxT1lLZ4uoC+MFJz1fkPOuu4A
GOyt7VBhRY6DEAn9yZEixSk3oTc21C1Yg8QrbH7LDxWIN8AFuY/gMQX7ZFppn8B7sTfq/zMiwMVK
clD/R1X+tL+5Kh4mXyKL2K2fInuF1KupH0Dk/ib5R51nc/kpMyiy17pGYwbILjDK0HkfJqQgwyf8
hI4eGyQD7MrbXrLIU//R0OHJelQTXRUZ3+VF+UqB6fQ4PLn8CtH8KsPQOQYMsEp2FUIN3avk6WeS
Cr4cm5T9plnPbCWzejMUMteFQbxDa1BrFeyk88tg4uuWxjkusOTHIUN1bZzTlEhJWkSW2UNULvKW
5Geo/JoAtFFM/2eo7z9w3E7ACvvK5xUnMTuZe6fQvlVWyAZuLCFCy68kcex8wOIJzlLZLmVqaz1C
AcILPtMWw2n8SdOa9Gp2GWFKTSqBrffxs4nQGdbdcBcvp05PsziAJSlKc2lFBmFDOK0WBt+hAwAs
ZiN8HE9x3yCypW2KBsWsl++DTl9d71PszG3+Ja5JXrL9pmyAKexn0bhfbbNnOBpCF+k0mOTNBVku
ZmEzSE29eaBbdEBMZvmW7/gpYh6bpbC781v/c9lawirmXr1koTr2LMXkSxUjPW7NAL++DlOmx01/
rZLp5z5Pjp0/1WnhHDxRIlcIImuG9um5M4QKxPvEoyhlkbogTbx/rmCCNV1H+bdfzrIJDi6KBSIS
jCi/g6IMrEGwZTT4iy4PoM4n9QAgIe8oXQ+w+xzidjUffX3PjGWEyyYByx8pJkfan/RQ+gXdNDZh
fequ6KRUv4SPmOmM28HIjq9UhopaukYGWRxOC8wpjaNl6bnWJiiiDva1HBKzpteW1FGEPW6PcQ1T
+iWo23QYTeY8FjKtNyvut40j+VJ2dpVxaK7Suo4qJlMr4ngD0RdiwjJ6JRLKV74pmuGJ531jC23A
4ykpZ5hq8lhpQFIba1itMVsp28DxTxl4+HBdw+MUE2eqUzS8pbKAngY/oGh/FiCTlZTqDdqroior
wKmWF60ODAx30vEIdq/Awg1T2R2vxoJKhNOHJJg5fCEl9Nb91qeDT8ybU/9joEoXELKS8ArcMyOO
CwmFnO+sgOD29TbS23HNlw680tUuBl7ARQ7rqQyyc+twRbkfL15+X2ZrJBJgq1pXukziVKOxn6P7
Jr/88vdaKIoo6hqY3WwilQR/gyg3y4wMlSRsam0ndYUYByJqIlRMsvAxToUpZ1DYmsPBNViuSTzC
UngtbciL2znn+8A4mrphykdMSA/cg+gd2HcQAipY9b4VyFZ5XlaFy6NF/aBbOW0Q23X7/YM0Cza6
p7C91cheHHnH5CSf4k46UxFXEXSka8zUrRwD6z88LjynZMlBHgDE87YFrIJYywbJtEEP4LJeHgl3
upHgWx4aurvXgTp0S/RguSz9pOP/hELBu55apHtIWYrAnRuozqznrFcJaQcE4lAnyzTjWIu1JNLS
9Y/hXCDsiVc/DFDCitCjKjtkDk4JW9rtx/x0F3YG5KRoXHvqA9sjsJN6h0ujvhBZjuBruUg8/zPY
eA+o0zDz1Vk6BfowH4pdtPWHxiaOk5etelbkk6ZNsq3IsiMsSA7yefS7fs4LWfop0oixLKNWwk2G
/Af9TgrHK2qP/cay6nnvQE/ElNBSuwY35fQ2GGQu86+2TSUVaHFFQ3L2bbTUdHHLJwV+lUuQW6sL
hZE+1pdHEEFxN3Yi/vHdXEiF1K6PMVKbX0d2g/ABV5ySNOxyW0/BbGXjgepmunFlDKgzPWaRuvvh
pD/eTczxqjGkWAWAjOVU4lqa0EVksneHvgTyttGS9Bv232tApL2APmLpW6dNNwLlJiQV+Lx+3Dp3
49CQ0Ofk0YLsvjL7Khxvwz9i/yc9otjQJTkqibs6Ri+tB1fhJGbrNY6Nx/TI6NMYziFLuNR6Jt04
Bm/CcLOnDHcfUOon5LywxTiuaKA+DkUc/uxRaHn8iz6LUTpJH5UmQE7D41aGWhgFAsir83hQE7aN
CFbtoYVPvzLqrZ+zH3ctt43zd1jiR8B+N0B9nsYQDvUiIOAas1GzveefVsQrgM3QB0UWYoQNV6M1
Z05fcIdR2BdUWABlZlWVQZ+KzDGEGK5fcN4tNZU/MUJuH/sCwD3QBTTGt/o3WJpit6K8SiSzmWrB
VKN6qcyByMsGNRpLNGa8Dp+yfwKUXXdmPsgV8mHfURRa/9rnYjyvoiL+iA0oKd6EafxgvtxOWnkm
PGroUvvSwboVfNE0irF55LBa6gWZh+fY0YGiCCT+ojijYw0bWTCDcKCC+bkgrAjYTM+3KReFG0xV
1I+FuETbqmBrVgxLfaCF5g61YwW30rAFE+38PzvA8K+CeM0Karj0aTtt2NoWLQKpNbV72CY4aMMZ
yYTbaVeFJubPVrL2/bSL1WwYkSXBr9q0q1uNbSIMY2xakAjD2/rvw0Y4+Xa+lxL5ns62TQgvYOSB
3GvDimpFE1VF7JnPfK3sJxbIDeNYjgjjPXZ9cuJ5mlZHn9CKZUGkSYw6kxdCLXYWSts/+gWYhOBK
hpZ2w/rfJW1ENEmIxWyMZhzzsL+We0/JDGJ+YZz+E5+Uk1tyB+QuPcekhEVAn497wSbFVXCD2SHi
DN2ef/W6vtnybFOiVnvKzfxSRYdmtAoXMxA1LJDSgFLQl4F5OFkcVz5qTQjglVX4twtGwbwlU1vN
aBmoSJS/xx6rJ9RcwgcCKZftwM+58GPQnfqoAUq1AyiCFRlAgho0WNaxv/OCfSeUFV9hzBTqgf1Q
2SNPHxC9NKQC8ODoB3jKALMx3pxmXrFzw23xgw2XpxdMSOOaLyHXZe5pXrz4a+dA4wheWsrvXCcm
/qY7bkZvUxq1AnHYdclRgk04kU4YAEDeTopM0PGChC0/0XMtK4TLbof01BDzyj0mQjtxp9c+qfXf
uxN2BBRZyLw7Jtp2W6EpkFmE9liobfd45asfqyp8evcFQZu2uQCJ/QpsBcTquAteGfOOX+q+Pj0n
h+cRVxd9/Z9v3auk5xGOov7bnrVkanAws5VBqSi+STtkRcMNWpsH71Hhp04pyIWMApx5c5NcM3DX
rj5mCPfFwLU6WaP/vEtM0YfMksF7UaL0ha+9hV7y09FtoArkC2OTI4r2oHw988AdgBc4IVF2TYbc
ZWVzhw2B+NKaBAlAHhpj0/LCdD1hBs/Q/B05MoQI4evg3LqHTnEOgek6WPLLn+1H+GucL3dM2IVj
KYkZHOgG/9Yrx+qgqh7IP+hWzNWf1ScZFEcf0jJBT17x2uiNyuMheVT1L6LnqSdNTNo2wzIAwa+g
q9Jh2AvEFRmB/mI8aOQTuRQSIwSusmnunaqdzVPdeeVxb22ssh3bA9JC+QpwRxF9L+Cco67NoSP0
q3viXprM7RuFFMmfLaWCjte0yjKF9Rz5tLlnhtDLziaiCpXjcPWRnFluXi6XNvQWVf2MNavm2LKx
dA5w//wpxtNXYU/keSMpvj73PqzodfzocSfG0dwISYB8/h8O3GmkedPa58sc7iROluiYBrrBXbpt
JIKFW6w8jQBfaC01yBhCsFQwbkRwHI5oXM/MVeMWjOtSTB0XEdhBUtSKN4yRHk/fh6AOJiqpkKRH
Qw4YlUkKxYK1GiEVDtCWaqnTLtywDijrm/wJaAEBvNK+4skllqDWKkvkY3keT2RCTLk/JEx5VEXE
g5mfXxdfypKsFzAbU87evdoTYNXPiUuCOuobbmk56MdmQuj2ueZgWUDH/EYLBnPTGOZhZDxsi4gj
FpLOvye0F2cIfCnpPzos3KLba431cSmqwfbq9qomvH1pqV5qkkH2cb8do19C7QZJ+RUl18I/ZHpL
Ivf55uG/vDkXK/BL0H0QboinYhgqalxzywM+g6JGxVXE7EZ38+25eh+EMoFPm40ouwRC8uMe3to/
jnRHr+s+kqoKsPPo0IZ7OhqSDyXdL/4QTi8g601KPTnIU1ONLGkOtURorBBAByxEILKgYvN43NIj
YU9HGcm2mNFhr4UwGaKuPLifyu0uhc1d0lS4o0C+Kr3QCSqrOhZ5eeUtqipo1RC/D7vzE0JV6nsZ
MSA26WQuIYBgewia1MJQvqanQzAQyYKPEgkr4+SmtvPung8aFjW7oWB7dfxhXtIfKKRoEbNJoCmr
OGUNrDf3sBr0RvymSHSm8OooZ/5ie3hvcJiasfo8ra3z66qHIYG2mFeq+VAFADXhoZoGGwyKBWWg
HLunyd/2T2ot318xm1XWLMSR9xULKWM1Q8gInzDRWAykSEkoLxccS4Rc6CNb1mljjZb3Dt7rKFDk
J8JuNIGTbVzWeiYSJaGWh3GeFMrGZVzwIXEXTlcpovazUxir1B5l0tEMqUoTXG63wnSzmKqgdCg4
6PqmeSATKa9GaNAuT4e9l8/SIyFImlQHIKOQo3HFfdCJiJHG5MgxRsExUUnu/1Hb1VmmaJfvrF63
GD73yWyrJduumlxyhHvyAiM4oHYa+XTdFHs+7yQh/stHD9gHp9N1san/Ti+J7SMYTeTUNWrB+1Jj
ebWHfMUs2MJWyV1E+PpMrLreDPT13ao9hGfWP7G3+yG89H1Kw9DE0NN6xwP10XHJWjxKWCoc8W3n
e9k5PnuGpyxBJY/H7uXrjpL3gHYZrynPwM5FLeWyvvR9urSeF/pzE4m7m+O9H4hbmuagv8gh5Iym
KALPnLT/um1Rzjb1cADtXcbGCDSvWqDyG8tnrAevl00WR/0vwpIl15WIgaefFBmijh9bt5LBlzg2
aNN4mxtYUYE+j0ameTb+N5g9Xv0hUO+qkxRLF8GbryDtOx2MWv/S2qLrU4Llb4On/3OSYNIP+u6h
rV5/oIC3OwczLYr57YAW+A9Jgi3qgL9nSDFcURWb/IkgBRzf3iUK+6VtE9osp0SRCvEUAVisxCWj
PwMPQB6pwCnEFPe8iUVzno0oExZ87IVb49WkUJp/4Uc4ARzx6U8nHRL4OM/a/6gnEQh+mhVR6+OU
Hkl4YtqPlnIlrdnrnDRjHzNgKk+mwCw6W+jzC3+5l1GAmMRmfSQy3BpqRWlRyVqiq4hRqmXO8aFn
c7kIV8e7pqFgA4xXSwwT471GiIyD1et2bR+w7d7BBiRcuMDnUhBjcUQncqNY5TaFSotuL6BfY3A4
R0TmzlOghYLh7nABryiOP1JGgUMjxPYNmroaAkKKEd7SEv3CQR2sb8IvrZG92KriUDx3rPMt0mh0
M1iP55JVwFczYbpul1v6Yl5jdAn3M8baTrHOAGc9N7huF/XWaBHiMbB9sCMK6KguP/eh2f1JOosb
G7ys6qPf9X1JAZr5FibjtnPdtrPh/i0MwfaOwTi2mI4cWmXjMIw/UTdC2LpgzdKQJK9vHrFZEP7V
SWxnrFaVN1VslZGmPYn7Kb1u78nNZmClUvvZ83SphhIES9wtPyMTRGf/Ti7T130wgmnv+kvZH9j9
uyVrZgC7cVjHi0UPn5uwLIpFrHnrzhym/4fg43Gm6bWwgs4h4lLIZuVPV18QbzVIgjbw788jr1YS
vUjGRecEJEEcIikpx1XlYVjOioTpjsfdaAUbQlHaU0gr15sP8VgFyAOPL46QBoMTsatdjw74nIj+
HyfetmX4NMsTHBa3oUeTKgaYUp8DaS/Ai8KNRCCekYKhUeDUJc58b9uqPmQdWMHsNqUqPs+zNy3b
qxCqnRNimW6WD3taK8psRUgXsF0UXxXJvHOUBEdAr819IP31sBHuukP8XtP2acNMxEyQQMwqoisp
ls4lydSUZgN62jS/5/n9YI/rxi4KFcq4B1DvLLhzp7dsFzrItOWm9nNDniVO6xHQTSKJPhUV/o1e
CnC3xFza8F2InURT18ZCUj9esrsHvpjlxZ8ut9kXcOifK5E+caMtDp7N8qcyEB/FociDbCJa4/4H
7RL9ooQqIcOyds+IWUiy+o/nUwzfNwJNKISyHcNs+cEMgb/ABktqHmxfe/Ww3VxFMS4YYRsXLYOv
2N8KAlgTU9NGYvQNKj3vLWq4lFbXffPWQrfdOLfbpif9BR2Dray4F8KbSpKcaH89ukuaJjly+5xs
+f/ygCULXAUH3E82MY8H486r5VZmWQAdK7Nle2x1zNzUlRjfNUK77d4b3HWVN5aGhvIOEDQQZ11j
c20UfeJZhPZr7ELMrPC0tYQqxJ8IDDSd6KBhbrX+0XYTwZYswI3HJqDM5qFKUw3qHLquGE7A4RU/
nQsTxFHHkFMF8Sf4ipblV+V0yyGV0pXkdjD0GYf6sV7WkcVEkU3zUwKSb+a5Uz8iDio5ZP9NpCE8
mpJQ+Ivq9ExvhEKim3AwtNk1RCOlOhir3VythIR/oTjMi2nzm1nwK08yfHNyu4VBkVFYMA4BBJzs
rL4Xpe6nv9ysoTgR546VO4fH99h7QhkBidkC4wdYck6pT2CuYOUWSAp0WdglcbvOj87s/djKRA+c
LDjqZBwblJnKYxNPWB/y+cKJfTD1WhQ5na380hNNFcO2p6Bb6DCMIAN+R26SkBQKxd/1TTE1I9yy
NLDgM2i64zjIGnYbdNh+Jid9ZPxIiS7hirL7NQ1lLJA1hKE7bq4T9Lw1o3tgJTXU3C50avMVviCv
3bPJtWlZbPHsgZlUJROBymH1j93uV7AVfAOjsl7Ow7qn3HXlfwfan/2YQWloWk3d8gPHKVsDquPA
kkG9Ho6kFiPi6KXULGQMZ5tDHQTLDzfvq32t6mZFBB79CYPYvIsTSJTpUqzdF1hz45+dAh/ge5jP
hHDXCSK2nsHrHndpDJdsaxlNjucFhqIPEJsRZXnWoJYW9wTvUwJkrgNZweiwMBTcdd5ZzVEc+nB4
tDQ7TJcUIFGxmO9slGVPJHyCaWn2vKjKLwiA8T4SxsXSjjs9TTN1gM3uX2cEGWt4ncnR5FeltpTN
4n8hfw78+cACcDAtz0taKgclJr3GjVnUGg7CidyXFNcjULJkHcn2J6WxtbEUbnjK6fGLxf/GeqJQ
osNffaXMl7qTTiWloVvDWHhdzZhocginutwZQ6Ey2zstY0a4Trijj0avUJv1rBUuXXyJSPStgq+8
FUkq8+0Kd+TI4Ka8LyQ9QqtFcFFc2y7pEWZs/V3RkH61/ZTMTSZTZkpecrF5dkTsZvMWGlycPud0
cLP/xB5+w0/pDUjUjCxMaUkrP3SJU0sF/KaHmopVIBHr9nzYkbqDsAHY90DdnRaq+ZkHpPdTA/mm
OoScCTMb+KWWLIHjenUWI6jzs04W0m4n3kdpAuVy6tInvMi9w23yWTYlc8kOAPizT32653nh2gjy
B/3OKeRgiyW0O8IssbgiLsP1YTNiin4jaRi7seaoGFQx5nKCxqe/GeaSZ3zZYwO/16hwJ1XGCpd0
XKT63g8lj4pjfFjxY58iKWA1RWjkqLqeHAdDluSLXqvVqjRRS/dx0Qrs6j3sz+kCEmlK4+yNkp05
9rJTFR/KfgEFEWyq648fVkOlH0f9731on7HgY4rAKsrdVVwwok8CU6muf2rITqBwWkpDrLqYGHwd
2dIyf+vTScxpYuCuqDDoF5Ecdf1uYL0muL8B81EwJ98Fgg8Dltt25IPsgAZroAlOK9dyyKUJuXJx
E3ewkiOGrDDKzc69vyVgANG+H9fTXS4e366Y8db/jcG1DQRqrS5Cgp+EI0o7uRKD/4o16Q+IoV8s
5HV+q4k6DR6IVdfS3mneIvr9TvV8ffY8qhJS4b1z7VhEPcB0VqaNC0m7R7ZFazox1lYdG5HtPIRu
KvOi5non5CZrv2HfLv4CuNzgkN/4pRV/ICw7sgGCiEV24evSAs4FvNCTfEfIzCmleduLRNqVvglj
t7NRb396Gm8k3vp70DyXwiAuYTTyArWDjQi70E5gWA6Y3aLbo0ybAOfQFKvJiiIHqeIghsYy17jb
MQ4XWwIOUGwSWmhs0vHyLEM1Fc0roy/r9g8JpaTqQENLFa0d9oEGaKTGxOO9qJvtaTJ4/W0TF1N+
Fv5GxJ5h7jYaZGDExEAnROKJIyrT2SKnQQapC/+ko0q1hvPzR1G2rrnR/BbetwPSKKdMr+hK+EXY
IU8Sk0pVIRCw151h329xVm1nqYJoPBbNtMtbrmJIo6/TZ/TNKPiPnXq67eehXWyWlVE49bjlIYGt
FccWKkcc2IRIDN24payW3KK+JPZoWmg3CquOZQySi9TeC26Pd4mYlgx4w/KeVvNliln/3kE65XOW
dMHxJJEWMco7MKyn/vASBK1FDyd8v3dLMXGJd4+GHgp1oPMB+jxjNbzi/qVd9Pb92WUJam1OFk+m
80Yns0ynFbF0rFf4/sD6OAId/Pu+z4F4o8AddY8zhXcfzlYf+0UEcin2igux6IwNElx3wZ0Wlh+7
UUH3YkwYBGYbjx0DBy83XUA+e4gcV9KDXs1l4W7itZfbpnYaTA2wXRVPcMFoef7SCwcYzaRGn2d/
1IVg34bfWddYK0XN1rkksS107ZwtWA/0KgkhtCm1bnQ1Usjy92SlUdsRmrVX2m3p5mGBIh5WJ1ip
5nizWaj5ZyMTdxGg1TTDrri8FmnwZN/wFqPAXU9jP/druwj9gYn4jJjKRpQuVnbZ+sbWYGVjIngi
cOA0Hp3cQOfsamkXY8Szq5H5tvoPatSEfu7/ZEBdh5Jue0QzEVHiVnjVaA/0crSSmA2mobL+/uaw
R3MGGFGVpoSiaV4riIt6XsG5qCwPL47lXFF9FR9i/SyIhRDe5gyXc0+7rb9Uo6+cIlLug6Xscu2L
9vjQw9fMPCn211HM5nWul97uPZpgK9B0QsNHSvNl+gTvCZUAw8/E5FJJQi3LJ2hRn4rPr+4HHoP4
n9g7rqvWaTb7G532KmQqFscRllv9jHECxG2rc1Tikd550i3yfuo+x2WmYdW7G+EZ+tXV4qfn/7aw
zNpP3geYjP7/1h1Ben1yte+1GAncYL6FvQ4e8VR9IhFnHUzjNbGSwU6YuxyU3WuDkWdDbpbE4Ivs
GMxAS3d+0mOZ07dB8S52a94Msss+/s6MbCdW2+Zi/pCBn52AAYRl5sG3f4w+rb9qFRpaX+FZwnCG
YLvynrZ+2kWpvPaCeJr5dNnr2PRX9f5IHn/2sXePHWq88Jcp38JMAfOWwIxcqo4INQ7SrRC1jGwp
o4pie7FHqktheNu98jCq9JKcNU1aSWhVqB09k8NVzTpUw2+3JsdJRLPgoexLGyd4xT+luX3BMdqO
ZpuVsy0IBn2ZuIdBwO/+mB4cCc60gz3YRoGJ0kxob7ovSEIfPPtMFr3jLoabt4wOXAEzzsb8gNNC
Mt4SM6Ep3fiyRw7wG8CQjphHAK/ZQxko/HUn5lvayGCDRif4ORCAPl9bUo3bqYbT9FwvGp8A7lhA
1kOe3qvBA0K4bnQNlXywo+poVdqhuMuxfiFfw4HLFW02ueU1YuPLjfsg412nUhpPvWguj+CN7d+w
Eq3eiin0D5qm6Qov5Zg/QmPRvfwtheStku53Jo/gDiddBvkc5LhJqIpIvNpW8DuTeOH03Oj6TdZP
Kk9tOM0fQCznpB+SzLgI4tWH665RexEUKCtfj9MylDGWS69hmvUMfS/mJVx7f0ggi6ulN+v9TjWs
mWeW9YBCQ+Uc7uexgA2O4wMJ1BJ8wMBZ27ZVI71ChRF4MA23NLEpb5xdZFWLI9TVRMxUuXfb/hAi
uQiuo0OEp1ptHfo5zctkHkFEeeAR1M9xbiNW/6qVgnGwZiKYRq+sx7wKOBiE9xRz75DqaxdoT1ec
YRhl0UEin65qwRfUAlIy9qJzymhuNbpDafFUgYOH0qXZJVW6fDgF+dT7Z383aQA9gjo6g3HRmJfU
5XfcNyOJavkg47HsPNPVXa6DFlvAw2KUgITQEhi3I4sxtW4cE6s41xy9HBKdsOvKYa0oSFlPKFLa
lpQYKXWdBI55iHBVZuR18e8Mmh6NzYobBjnDcJ1XMRzrIYvK+a7QceEcM/Jwr1bEQ0Pbk4myL4Wv
hkP4Z/gRxc1e2BOg2ho84O38o8hC2x8SMvrut9aXDbLJzya9vW0rbFrlsxzX1TbeyTWY2dC7e5Kn
WqS/MHgqv50KXpEWsVdCyWqBpfUBYiN2GiOUQR4W7H7dEz4bfwmp9c622P5yWA9UShX5sdEO+COE
8KCQHu9hvyfWzDxQFdVYHp9SaqO4k9Exhj1/OeTWEr1o+qo5DHFjMfIPemi4A7WQuKeJV873madJ
e4otmD2wY4x77HhMtz/MLLZhKYrS+VfNjtCrSNlqM7WPBsplcQ5nr7aO4ttacrLD8KVgA/Gm5oLi
bngOMVTOFzvs9Iig1CfGA3O/K9kvknXK9rWWHjNYf3mKwkRknGYNNdtAt6J+tdKr1spQvTRtoVIj
OpeWCeoBFrLxbDkktW09Mh0DzRWVvc7dMgrg4X5W7DIQhJ6F9N495A3lYjR7OmbXBzMGiuvO5Ngq
m04nOeuya9TeuHt60oBPfB5C7mz/as87ZLaaM+r2EXrpet7rnrbkUOwTi7LKFLFVZZkXJ759SVek
WioSui+hG3jDhEheziAavWf/I4hdeq2cUJhnqIXLst65TwqOIBdED22bJgtGTW0cPAz1vS/+SHIJ
raHEMKz+5yCrAa5syuX/uUHA37XkF4iNmQbtFNKWm+KyZ1Tv9kzWMqqbpvYgNQ1rec2C/fR3VOuS
arlaDZZ52iDYRFQXCOWmkf8xOZYEnz7h5Da5GPlFQL2qDKvxrl6pzPMbfxoJnTc7apvn602aFmyX
wgkbRwsXvPBapuRfC3z1ISGOB2yfRZsLwOERzLPjawFp+Y3Y9BakrnnmQdf3DnMq26ykchtFMdt4
XN7oh4WoJvf0+dFWPLiKbBoh7g4wsdUQpy3FPLjNUqDcca2a+Lg2N7einVJ/kV4Cb5kn9ty280cR
bgRNq4n+bkDxIKFJ9nB4q2PsgUVoxysTQ+1wk3vWXNPVEMRSPdiiwZAHE33iQb4IJ3nInTdJ25qj
6ijq0Ti4MDSecvrF5XOUSQbH6RTx9xRGq9FqeSb0Bdy82HYWAZD1VgMFO33z8snwVgDOqdYmLmaZ
45fbuUPiAqHuOSCb0KOSCL8cLc49QMISQEdGtrWgZKdEL/+vTaqmrouyI9WHLf1FoEyLEFF3XjLk
yRjtKUkB8tWml6Qd29KPTkdfqUEA/LKAoosx4/P+aRrS8OiaBsQKo8QoPRxnmJ293Mjn528Accjm
0AJ3oT4AQtevopfAMblYuZsgvQCN6szWRemPQrQ2ovAu8JWmESX6kLyMLgGlgkdshpzlUeRt/RIs
Nm4d0jSsEGAZb3Bq2dz7YDUjJ8hDYWUy6sUcG+aEPr1LfcL7sbXDAdZ517dom7qHuPpoo5BEVUXR
m5HVj0X7FGNvwwOQpIal72X5RiPtRkcQPsKnCDEK/9H+vWB42f/lpdAFtjDmFQIuBsxLqriC/EKp
nNxdNeVbn+Dpox/fkmZPeI7bAtqQHKh6J12g/ooVSzeOPj2iuupCvmE7DbrgbmOWTHEgp9woOrzS
FTvBRQJUeVUIA5/admv8S4KkWvGfdWEaUZUVW/jO6lXAgaKFKRHHrwBGz9f+i/24uiz5lzehmhlc
+5Q5Fef9rPvoENTgyZ2Eq+BaWfT+bC5AIhe9933cVKI054PK2e8kUQcjAgineuctxINcBTwn4dGy
sOqK5kCF6h8PgwnBX2SQCMbID0RYr2ymejb4aSYQwqZecPRMn9DKMWAN/yOrefMFoNQjBDGYKccU
hQWgbn+euyi0Q8peSrtoKBVtU/PDtNMDT/Dfexatx0/dH7O7EpG5X8Ivpc5i3KC0SF8da3upMaUv
xH5Vd6V6HBo9Z4a9eLyAb1RjboYmmRmxdyVfsytQoql28f6gP32vtrm+qO1i5++DSaqOWkXwXQOS
uITKLeu5hIrhF+VoMfdBKeqhfpCPbDaaJjfwi6w2Q02WEm+I+aJ+TmmanHW0wrn9Dd9xKEd1sLGr
c3qyMPcvmjNVARHBmFGTMOKaqyHeOVhkB4cQOtN12jTJ8xgufTQv1qsag3MGFmcf6XeZnYTtO+Cd
C1pfzazqHSgB1MPiDlKRC6gdTrGlI5oTg6H8jLq8EQUDKnChIa8SBzVL/4kmaf1UfDg4Hb+0GDKM
AyOsA+qn5uVs5fA55dF+9UVXnTcyn7ggXS9Hy6IbaVojXlTdkMIR5+vCoVXAxvMXVcNKrtOyWe5H
QiI91kTXZVQwrQ0l5yKZ1IKa7VhPxvrBr7BDpqCVw9KKEt25MssJJQbXlDlShsHXecB1xISaJcGL
9/sxvWBRUkE2l1+4qy6usfpYmy4rRMzhy9nqTmyXY4TgBntsYHNp0pG4YQANStU52IDXfd3nqatc
6aHU84moJWTT3YO0NLKnh8atWGsGwbaOr2izNXuuoQPJ/LOu/E/vH7cWhRh7V7R6Z1EaAA18+o9R
yYdbenou1D3M7J9q76tAqA8cvQKrZjg0wTieYFhV84wfoy2/z5rWFJj+irCpp+/lx5ozA7qAeVJD
M1HeDh6tNGubWGAM2qding7CLzRmr8y429Ex9uGbOqGFrkUAICUvw/+vE8eqe+xVjkuLseq75DBd
yL+TPXqmdvSUCGi5gJDgPEs9oXRpn+qdBjvkByORVwdbwvGKFopVDp9SeOlHCO3SAlqnvgesjTfk
a5dpEFQ9/6FOg/8qHpI5Q1NNKXIkqOV4fr8bYn3C+C0lM4cYkT+hzJ2p6l4eGlvUFS975PKYkcsj
8XnJEnFNwqH0yzritXJLT4kcc4vW7eQZc0czYh2+Zdnnoz1h0rTuWEQ7/vqUiLABcUmjGRbLsKMv
Dx5y7rKD6r1MmV/uEijcWomsgHQtKgJeK4v/9dlqtMJLZLSaYQJ0aHhAzLzEaClfCz5pjh5hjvQy
FOVm5lnDXNVBT6DEBNcBh9XoRKC94TiIec0m55F2TKZ65Se7/AscCaZKjhUSU7xL9AC8J1QUJOUM
P+AQLfUYRbOsWnZaXGKvYuaTGvB9Jphwt/0tdJGdSGXmSykN2/0G2azycrTAA7RgLM8WrlyC42uR
xeZiROCo3q0Ppo4uVOR2dD/XuOd273DJ7hkmrwTMZFaNmiAWd25Yf21ee/CJyJ+LAaO7YBWjnFGS
ByaqQK2gkVczq2CXfRp/L+XcO9EAn0Uv/teHY+/8kkyUG87A+dYwufAV9sv4jvFP0gaAfGxCbDO8
g1Gx9YDPJi3JsrlkedQHomZlaL53XVjeHR+ZFLFv+m+mz+cojSw3lf6y+14n5WEpMbWmya0Th8IZ
oQteban8aur8XrEeThfvDlD8bcGX9Ssb5u6W73oKs0mfRfucC4TvNyf9nPbUSipo6+m2+Y9+Ey6n
27bdGyQ1PScEomh9Si/tSC1WIOPw60hoikEcfc9s50xCgG9urRL1+AmedHk/8sHAl9F+1ZVK/etv
wnA8L6iMe/SOUzGyhir9JflzjvvgnMrf4CxTEiGMVYhW0q5iRFKgsP71N6n7FNVVA5XoPwbc8iDM
3zWPyLE1PsS7jJ3aslOABMRrpb8zwKX0pvbFwOKCPBoXpmeOLZxdxM9O2k8lIEnXKiR0RSrI9ngb
RQKxlqBMDx0Jap0nInwFCdqMYEwy8+alKQSEnaw94mLGlFJ9ezE9RBWM5EYnpVpIILvQsjT4y0dp
ljXuv3cRgzHyfQXlkQTAGHAfn9Ocu90TOPxMgt75uH8O9JDs1U5n5pzFbBMUVhUhxwz0Csv6NNp8
iA4ERz51vAhbdWZ325shuU3NrMczZjH0E6Y2bHq90wGDcca4eZzn0HThx42AfJCGgxonKE9knJPK
1hTs2Gt7d4NPK4UpU5Qblvb/syOHIOQ94JZVHA4Bhs4tk5/fR/2DNzL2VTkq/k/duYvKcJUL9kWM
ukfDDBu9O0jM7ep9wuzXWH2cay8au3ibJygaSwhy8rtGCxEOTHrXEorBnk4ZECJGjdZgZZCd/b5z
dGdxl+ouuTpBxIBpzeMXVCcru/tcpqDN0nGlkYZY6hc75b5FwJJYEY916hN0k9+TQITjbPODR4Gb
Dj3P73IfYcSHMow2ZJ4AKNZKI/h+pCjcxv2LopEM+euXKaKemjEUF1xdFJnPebpODLejVE5Ap3eE
tTo+qqo1RAQnZsAET92iOA3ppdb3/D4LuyThdqy3FPQzqD+QrrViBgwwaFuPihTf/RGzH07FpMO2
FCZsj6T3cjselaMgl3hnMeYNNCEplw41tDOMYh9u+z3uhTkWUpwCWrZ+xEGeG8fEVqNCx8UMWg7B
LaQAgk1ohZGKOHXEvEYiaOSxGjw0l5clxQNcKOkCFSbQOjuWtoPTTGUceDINAVOiNuHjp99JCByu
K0mpLasPP3DeBAz8tSg2X9Lrl74vXI1qu1jiwFrrtwxv3Bo5GRnai6xTbQo8JwbttVKWlLCObX3Q
Aq5LYc/RHmq9+zqilwwM/zBmn2GhZ0Quhj+Y0C8FP6zqLbMKoXQzKOAPaWH/TNYG9E4g6MGPo98b
eMBycf8TLzxLrGz1TWbp2+7VMA0rotOMKS+eIuYZYA5FOFu8FxGI8w5baLtbhBCIGsMkDPhzVQ1Q
H4kaRn7GoSseROOHoKcWvTtjxvBojIjTYPwJhNpBf/uaqS24dmoN//BzeVgaGsPGi7a9iBq3mlQW
jl6mAAT4UI58/VAGE7SMjo18PDE4vpP/zItm91YtVyRv/kQ2cPPhSuDAZNUffKobovB/GEoEFUwd
pLmMhNYjOiZWsTx1dFzh3EIXoMXrsHjuT/5sbGks5bcAYMv2NIwka98qVXdmwYZkQ9tULx87Z89d
uZtaHHPmcDzb/J62zQ+RyIZTMyRkPy285sd29Cuupz9d+5Ms5KZky32mkFJoEIMGPyi1I+h+WW2S
mUEQWTk2XSb4c7nY82KNg45tbou8Ze6Kye2O0LBya7Fp8RqKZpuOBulD3cQHxM9OLqQQsJPtiJF1
fXOFiBaWOf5bl3RiT71qiHkuqObNyX0rqfj/HAH58s/h+wsk/8DZnkefW/Ce+gsrcEf0OXMF88//
3FYcwy50eaojduKN5jGXi7kbKIzvrrhnmFC2ab4imRWD/t/7eTKKjv0CLl4SOqD4fu/vjivJgry9
Vt1Ae71wAWOTEXOdS+rtKiibcwG8I60OYU+m7icfN6A1dBsOsoJzppUJ111mFpWF/+yYChZ3mEcz
wQiPFuI0s6gfKv4GVbUgkCFkiSY1aZ1TgWbqKbTM6q2V8fjnYQTO2upWtW62PAkcoOy5e0HmN9Lk
LSj/PdVksZ4DMCqm0G70u8Yl2WoFG66pweRXcwwobJlt/imF3k6iU3f8JGhU5XsGQpb/ee0OPMDa
n6L/PEUxnb2lV120Ov0Y7HlSzEu7tQOhwWryQH1JcFytGo6VeWZcipWOnzFMpFkRyWtIiRa3bf8r
7A1LdReZwrj7r+BMek/mzUFlDuAhqotczbzBh+pW3ktDgj1i9MQoVRjJcuSptSqdNhDf7Ly/dp+x
cRuA8wEZbmFs2keCepRXdCp9O550SivDeJsTtdA7ASUPnp3DGIOdppC37v3Ior0KTE/EmBbnHlmi
YqwjnWcQgiYj+OxYsqrea+OJ1bHwZ0s3WiFPTXB5F4dse6mo35bgdmXNS0atw3LfU7qBlsIdc6NP
azhLC0xAyuF1LXklEbCxjk7IxZhcxI6Wn/b4GpJW2cV8FJok+3NqmBxzmrQxSAXWppi2U+WHjzgX
IkOFDeqBWhQVhmMtLKpIyqf/aqChTCFS6z4LwA6GGaLR6sA/jFetMs09CUnz7Ch11CqAPv8mH2P1
f/nfNfvzrmtF5fPVGMnUOtCXlxFM6lHbVWp4/N37nYcyfyMY92FDDmiss+yTVeruC0ajGS2Jjn0s
0aT/967gl2u9nYNYJa7AcCxi288n7ZhTZ8BXndv6gLNrwbcfUS6WJpEQfywphnKm++jUIl4N1dvN
CUYq2LXmQ2HwFwmANHK2g8NJ3rlwH719V73u9i8N5VNlaCfySPriIYGjaYwV5hD9bC5ChyIuNPDi
EHslp/2UfrYDJixN0MTxHidDYA3dRJZROs0Cnsel3ScCrxuckz2S3/ofY13CdMoYORS9frpB2k35
q61jiDvfwome3Zv99eK8MGtZU6b1Qz2lEcEmRVltyCbJcYj3dL8M4WaTBw13KrDdazpWJCcIIUZx
fnvJCMWLh6GlzGyLr8osWURsw+og4+VJGdyOODaOOcUMIIOMFLPttxsodFT9Z5LT/yC85wDtKt7Z
vHH1KHio5/+Cesyj2iG8Gfy0T8+2+Ssp9njAacQbf+VaqGn7t5+b3MwqzxZIBrfBRiqUZlOYg55b
DTumNQ+aVOkqWpgC/iH9Rt2st0QgyiMSu4bat2vc7TSjExKDOAacQ6cJWG7NoUrOD9ttEovmKPql
ReBW9hqFM+BwiuGAW7N0cy90JdPePWolQ6HpMUY0bqYIWcDoT2BbFIflYRsn1k4BlUrsVau+uDO3
GDgHput5DTXIwTr4s4syd9jgRNqX6E6orRM45H8Z4fInTD+LlnBou6YFAznWxPf1tYLfVRPhxz5j
VfBq2CtmUyoR/9sPg02EM2UJVJwqMYs8xgF6DegHY/vhpeZmAE3Ywk4uVJFvC4jag8DWUJ0KvjYL
XU71/WCM5YCRpdF3lYryyStJQKFbB24nivcuozyDh3C4GpAQGWMP14S8Ki9+GKgjdv3jqxDTTEGa
+5NhgqylQsHwScrjytuftjaj7eUbWK2aaKRva2ENapffh28HkSl5FeZYgz6eUHxrtnrCbodyi5Hl
JI5xpfjVKIeidyH4Ps99pCLxLfFEwi2EjeL0OuBj1ivy+oXO7x1f1dxAB9zGBD08TcX4il95ryDc
2Cv57qO6ipmRhosx6g/LRHSwsKTXuxbx/PLX1aGlu4LGte0OZvKRlZvzqau9FeamKVyjYAMM+XTu
TwqPD+UqdFowj7pqinFokI6rC3H4QFpLJVJbNqieOuBGJ+dooTsYmQdaaM+kC7VyVizq2t1jDYoT
C+Wu2JoIxnlaIbISASDKAKGDbiNjyHB3TuHHz9Cp7G4vNKKLoKDUy2dNTbkc0Ha0PMYZInz0a9Z5
DpNqxnjFtZr+ixNjZRht2nqUpxkZtGBac00ww/r6w1GsVxIe8vHOR10R/eTiLSlZndOYPPK75t6H
U5gQMW8X9EbwHS6CKpRYb4xy+D2udhhYwBwu3d0k1ZrUlVr6ngOqOS5IprPUwwaycftPFjTI3ZnT
D0Xj523f+T+darh2+Q5numxFp7VWaQrNnAaVUGhn9sK8f802x/QXByb4+lTRKJ9QUoYlZsy/akVn
wftZKrJ587e5MHiVmEtlLYx4Y65FT/wGedQTWSvsaBcdn++LiduTCxGXPf/zi6K/KclNeGOsAff2
CHupdgSJ/E/cXodtT23P117xIaj0DW3RBjq/jZn3JG3sGbQCFFCIH+ggYCH6GEBgqT3Gub4u96bK
dlpaMGb759yI8/c5+uyVsQ+3rctXyA6kf+z+4P6MgRb+yw1Nxhzxf0ECqAhYKerY2BWRrF2JHbLp
CBVPY1XluXL1l5rs73ujV2P0MmQlrWxT5eHSybA7YiCZ3nHbWnr+7yi15dWluk1ZoiJ1EdtXSJx6
E8tJhAwA/NzwY5GqRw91hObavCdZZmlh8dFhnmJRLbodDPF1p55SoJtoaKrRk4eBzkFe/ccnbJU8
3XLGhMUxiA6aeqzet1AelgX10gpQQ2v/Nq+vIFEDykpLQclM5FHEiJF+XhbYEFP2hO6Neq9NMqQc
WIRc0tRYdyoWVsn346YSM9GicQmX+P7pDR+3vkgObqqswfWfzZpW73L8UFwKSa7S0sGKcFOoj9ZO
kSpUfd6Tosg+AV8YH3wzXKztIOV+FfOMM1xNeYS/jcis4fCqwnyj7iHLRJyI2SK/PH80stCHEjsb
kNav4wC8LHXhzKSo5OyGmlTeToOmIaoloxrlLjIAvWonZSE3h+tL5Wy95vYRRiC3P5j3YEOvJUjP
qzUGfMKoa4tRW59V5SpDSEalhaWLWIqmRo0W2EPnCldaK1wNh18Zr4cUY5S4b0TahEnjbKVb/QDJ
Ji0d1WV8IJm1wvAz/sveaxVm3RYRi2aGhZnGBsDJQ64C4Nj3qRZ8tJgS+KECJcaD/SvRMaTY+UXR
4u9l7iBBfDAYTY5XyM5mHFAPA3++mbTE7VROgp892OnxdYbSeFHnmjT32C12wDNfG2MFcGn5DyaR
ylmDm9L1Kt2sUlSalgk/iOyIB/ju3SAMsDbDAMNJSOVIgzQ0Z5BBoE19uFnmvcTLugBfvSr+ZsEB
ajf/jIJ9/lafKb1OE2InUV4ZJcKZg7tmwiQ2YxuYsVtv1Adl0XPzzHNH1hAOg1lIi0PM1eczsgLu
cCqtgpqxqSVJPSRKjqboockBh9l3pFxVP9GtUb/Qh+uYX6rSXVdBqeiwPlhOV+Et2kyeU+AmLxQG
ULmj2WTsC+KBXZJsTKo1TiaKMPc0axZttadbVnAjrw5LeQWqTnISoW3qy6MtjM5hr7ytt22vpMEj
pIEr+NIiW6dAISgv2vz0bDeG/amaG0fY8d917yhrVNrZdOgIfqRkJDdUYekX4tA/MnSmmL8FTHXq
OWbNM2/pLuR0Sc0HSmPICjLEz04UbPWwCCFqr4pMEv2NnewNd7klROvkJeh6JLYAiK1Wg3KdrODN
VSCrfnOTF0xEt42LRSrnuLbvZNAiVoJkx8GSqIQdbxGkwIReoQ/082mTUB9ySUCQJOfcgLBVudnQ
5J8UlBTc2OxVU6kNtdZjaWQCMm++9kppwpZgND1vGkw0nvoB3OBrGwyDILZkeCt+i6wLkouQrvuR
Vcfr9Qg/phfqhhmZ7d2p4cRFA5i3KYH7qj1XfDmzKZmBwwMq0YI/aT+OZdDZRFQMA2QjCr94D3Td
Hm1u3Sy8g/tipp8yDt5DytS6uS98X8fyyIjNGLGcTlOCC6553WkB9FMKugPwTwkSmqOiVFD7ssNc
keiB3wu/Gp6WJBDw1pB3UGcUpnZ1NwbmfjOx14njWorgNhgfT2JKsK1GgJo3YPMHcKeiJpVaua+Y
w4aHFlOXSWS58WUFpnZmf7mnIOjYPoEwGppMJeUgUiYyEv9KVEywdft/lhPjkloh0sWXda6VVNkj
8s58dW3oOkzQsxEvALq/Saz1TcZX6I3AYfj+g2Wm9IaTgZHZM7lLNN6XnN4uYC/N0PhirFTFW7Pu
Gs1DQwuuUtOYc662IdmrCADfaO0IW/FKNDosxQmk5tck8JACmdV+OZBIVhf44VtzkwNrj9zinI/F
G+0FTYAinpsPA4uxkM4w67dGnShBc/KkhXsC47nxfOW/sv46TgkyPWJnj3Rb1yNpxcyzUcPoYxgl
+mU7VRee1kkiOoxQvBZjbeibBgnnFK5/D8aUm5nb06zG5SJZ5B/riafa9oJEpPu1xUgwVzxExAnV
AhOFXHqVfVrYDoYyjJg2rgVQtZ1c26/K3tNjHU9+kisuOAk+WQpFPQ82q08JBxLadYV8KgPab2Ym
L89zA8NqfJ3fgUbataV0JRoC8yL0/n6FFr60bNS0a9HyL9vC/unVYLQyRsa+YvybF8YGomZ7PUzn
6vzDkxekzS+MnQLJIX1NFDQGtlYH6SRR7FZ7zG4gPyDyhLEn1Ue/L4kvUTa9XsSntNMuUqFxPCqm
/Xp02wyKCFngSJ/9AcdgijYPAZ45OJ16FlQNsPapjFgDdA7T/cSN5sTZpGzCOKTxpJlpfx3wGYXj
LgJPOGzTwXaAlEFzqGOhBJ+7OPA4ombCtf55BwCpoz0jkerpwAi/0OclEK84RhmEbgCaxfk+uK+4
VP4BHiTYm7NXtZLXV5dG8SHxmhmNt9VTQbhjdPevV7N7Dn1vCJAAMoneKpI4O/bUJZCIRE+ZsC3/
7ENd6T5wuiCACQ4nhapSt/hPz8WU1Xx+uCkkcro+OLYg+c4wlo6+QDdEqFOT1ckKqeCjHw5Tx0LK
amOacEr1B49b2QA1cNiQ5OqUQXysl8gLnnJjdEPU42Rdp1QR+YJfqGU1Hp+WB6MpUFBnbyOndZzQ
spz2k84OrAKjyYeX35/P93sKwKbGSpHneZOhQ/O1dsZ4rCyIdzY629SodzG81VAFF7cy4EMovGF2
AA+gEuE1VjCblhjUSdXL/IYQw1PYTQgVwflxWP0dknioVbA+xUkm0O9tTj0pSVyVi9xD76V/yJjD
lH75f9/oRC/ckI/EMivlrMG+/Q6gj43UaJ2FNhEKLOvR9hPjQ4XOpxUgt9FY7SoWMKfBb5OlZtbT
IfzM4loPBThi1mRsyHAzljKWu8iiZ24aZeqLlxFWkqWmCU4GArQxWUFNkPEfAQgXuEKebbnWjPKC
b3BbzTIXH3e5YsjR3wmInt+2nPYGDucMhul5pOjJsTlg5O0mI1zuY2Iot16yKexHjpqS2CjpR1CT
lGv5nbe780o6qGzDcmSIQFKnZVEFDwN4CtVR4fsM0QbDj29SdOZhJqfoSzADf9KbB01+eCflffM/
nhKGLEMDitGbHfRhp45G2iDkBpdAFGkEH6R9OBHK7sEqNdY9O3jg05Yc0JP99q8fGEtZ9lxHR6zR
1IR4Vbc88LbnbSQNBuzdl3lryKBhWZhYo3gTF7eYsi6qratz9AJszC2w5T3/kHVLKD2SYyVWXFUS
Zt/tNGjPj4qkg7EN/yWldIW2z4WIXEEdYn59TnGB4oORz/B74MdlHwWqbRsEZ1q+VO34I7veWsvj
ZchPjuu8p4OR92s7XAUw7qrDIA39/x6qa4hy5Uq0ewKEnQNpdbNr/LZWS5fZSnGV1v3JA1mEtTRY
rMSA72UYjrxXS1wJcIJG9bn/6ZoKZy+xCWWhwDPqfbMcgWZF98aysfwrovi9OuIhBcZCV1Vsiieu
0ahUkX9KB4rwavy18+bjE1te+MqSfCt7/YfdGR/7DtRf06dV1VINpLyJOSw765pf0S1m2WW3N9uV
G2dAswRIKlQ5DgyGMAF+9h1o2/TJ+7Yyk1eXn048ip404m4R25aJTulaG472ol9m8qQj/G+hvhoF
JRvhVggZgXv85EsW9X0eP3ro7c2QoRKSw0AmZNzeYo7Ptukv8s3W9EW16VP2tLiBVXLniaMC/mjL
BPxmVZYbmdXRTUI/5UUTDFYzXau5Z26dkmqhl+23kigtqYIbX7ArNcSq+yAFIA5jqYaGJeGCpsDL
x66Mb+K2oF1vsAQNUxgZ60nKEXFrij2jckU+ZcW2Qz/je0mQtbhdeWWQv3HUEldXwE4Z5FjT7G+L
cxEHNv+OKNsNGzSRoCLGgZlQR42rq0zxbQShsqooW5njBY9bFmAVgi749/JBqPDCveGmQZLEZlWQ
yrKYHQEPe6YGXpSEjnoZeNzxLBVr7l8I0gAmOWKjx4v1LZefrFhUhCa0jjpIcHXr77wsQ9en83TC
XBwaLM/Jvzb6K/zhcqcaSu1eP6lY24UThqQlOAHUgbGPD7v+qazlsBU31LL1NeKhl4268+paGjVI
AyqcklgoPrI69XGNo1+u1rSVLhwgntzdFFZHO25bvC+pm8G52Y0o0qFeERH+KRt614wd3twCry1D
t9EInEChb37UNsjtkJV9ZuHNEQV1dwezTXUNV+2CEWleDG0u538SrZ4YaEfuXO+ionY5HmiPcCMu
RHcln43zKsD14whD8KUQTYhkRkb4efUUwF2rQ9GKoci9s/Mmw6Vkdia7aQr6BFei3IFpX9FLl1DY
gPM2Aw3uEM6hqWo7zX82o8BM1MjuG0+/SO6BxtIyt58ESwVyYpWdibBtS1gYF+oKKAKaRp5YOPMW
O8CL1VhzS31WCGMW/Uc5tNjUAbY+lEbPLiTe2j+MDjOxOraUAVBgwgoIgvV1j8VoB9t7SoLNeE1Y
Aj/IOZlcZ+MLDSDthKYWSgpfNHi8A0ORbQVz84OLj+Nzt1wXeqd9ziaew0NPklaRsZcmo8HmeZIt
5gPUXWB+bbt5fCsLO5EV6KdtJr6TllYVK3n+6hsDFreUsPWBTvuBmasaFJyqFubKs0IBG9HoxoYo
MfEPvTIr7d/XVLLysWZPw4s9E5ygJGfIfQ5islhuCRCDT2SgemqL+1WbPj5Nr5mj34ppPzo3XVd9
kBlVS48HEk5SOqA5zRPCwBFjU0rbYHpNMsNAZBPiiYDWLCXnG3JkWBahSdmT8vxdVzFNwsD2zCpo
eZ57KB7Wrmbc84LYwsOPkGyBozxmt7SeUlqqvvwG/tUQwSXeh/FcVES6MEgie2tMxxjaqQWQjiQ0
qF1waHJB9PUdK4zusfIjcTs1HD60DOxjf1hxYLd5K1GoRuYFHbXvfKfHDCwqSANvLFPFehqX+ayD
I6Kzdk10SdKurohhgsMroQksuF/GNKrsdZ4zx+X03Wxel84Rh/7Xn1jsN9RM0YNEPg80ieIkAZo4
BWAUIz3AL+OOSDeM2HNBYlSRxUmPeYG4SCczyfY/B89+YPTREURkI0dTA1dFW2iZxskk+Z7PKcNr
8U8RZ9HkooqY1nNzu8drHa9bt1GHnDsFfMPLpsZRUk4HrLvLDZTfeDkfj1uFKicz5LPSDCD7L0PN
P4g0wBrQKy/UV4WC2K9npk7PhhhXngW/fVUL+WKVrjYmbxU06UMYh9GEsrBOTCy5UgoN4z2rAYPU
oU5XJqn1SbiyswFOFaG6y2EvJrHfhaKO83oqOAo/Fv4rEqnDymxaRxyHOMnkoIYZOv7jGc8mih1V
f/n/xm3ieQD3/ilbbXNgJMcJc1U+MEfxy3jncQIdS+gdfnt8Nn3qIv51FuigPBjSxk58QdGxZaP8
Cv7Wmgg9BHDoBydX5rshqihc2u+eSYd9xUGbnRqdg247NAaSKP+mPAadzM7wF0CwjlnJcrhmdeun
t8DRYvdhiXBAC5L0uuGcqJdsh0IcQqhmarvp0EOjC8LcFfMYPHB5N/3EhRjSv+0eHhsT5NR7bOAh
wFW5NcvuPPl/XKbb/sQolEqUKwgadQjuL6peKgsjtMw+mPNTsZYPfBTYZJd+/4ElKvTAqz5728Bp
Y2BpvOIXxlo2GrNc6Yip9zaT+AAjcKA5DMOPCU72YngssMXCYWY34OpsXpn9PNyuq6xAjfm3dbAg
r5/5ZTeZ0pg9wGT+RNFz1OuwicmDb0xZzGutQ7FwrIpiCj0+Ze8GOkEIH2NUH95dbqYWWROioX95
CKD0pBIXzJFz7ZjAMRR2ohEjP9tnGk22r3HlrhAWtofgt2oB7HMsyMqJcMed+ZPGj0GJcAZQ26OI
IZ0nk2yonoWZMJSiqv2a+HfwuKSOXDPvZ+4mot/07SbW2RZ2ercjHN6gDn0Q6Ji4j8badrqwfqA+
ta8+FgcIEmNdtTvsVMFJfvLqmF7hJZBfPuT/aR9wYEAyqRc/zgXUYHd5CGG4VoR6RYoJBbkvkgqZ
cCTKUS1NmyOFXDz/OjIE5pLtqsaCCJX1qv0AzvlYu01eGMqCt3uI0LB+vrHU4N43x/29WLBP8lL6
LnOPmeOYsOlmhBKGNSX54s6rNz3WVR3aLDDBJM99RIdLBo6A6wmQoUFbHdyt7K1bjyQbvywWiJdn
lE2mmNDZ8fP8F6qn4cAs76OB9cWe3a+aHDkuM7Iqmb4s84vByqtEeyPJ7oWfTP8jxg+/jEIwJVHE
Li6SWcNRJzsCw3mBB0LZFCONsTfCy6aUHEhNmy8/daRdWihG1Ks1b5VXcbupvCEj98qQxFmeJJRg
ktgyBxdeiNsqP89atCOuAIDxbqoYBAOYQTeqULmFuJQ5G4Ffx05PMWkpPlIYfBhLJWquHMyMDgG6
AzBN9Jso1Y88IpfEJidjeAYjtmKm0SCES9LTeTBwgk7LojbdDKFJMfuxEnn5co5A/EW6aV4T0fbF
7OkntqfC7ZodBoDAXmGIaLR2vIOheCDI3m4fwISxjOqoTPuhjT+9tVBZMx8yAQ6hz6dK1LcJhXnq
5I16/mrHkh3BihvJRu3p/oJ9BAFcxHuw+Re1TKRgMgHSdjoNZPuF9vlpnc+O6sTs/EK/S1V4+M1r
NyhtWXGCYABm5VNvXWvi1pa63wrM1/k+fS1SHJd2wBBj0WFc8eMZkJcUK2Cwm8N++jRNwnSClMvS
fY5N7mlNPPQ+MbWFm11s6I+iAHK6wOSM88PAWbbBNR9P9eHUX6+rK+FAnc3vEAwDmPEEqdtw3UXA
LcJ9YlyzIMJqySa6N1cJEnuL4t0Z+CuQhgwWnnP6c6wm/2jjstILutpefq0ScbaQVMsq37aC8YLr
sCxdiBuv7Nmr/xfB1iS4RazHkoeLlGxRVmRO2wLdrgzlZZ1y4Y03EPzfBb4lo1UTuyh1UPv1kCPr
TD9Pbmj7bSEzF1Ijz+IlWCUkVzW3gw2f4tYWWggjouGgKktNwppyv1IxRKmTVV/XSpSgDeMkqXD8
ngB3zvideaDW+9DwAeeQnvJY+a31ghfs7rbyAZIu/85lyqsfVK2Vapdl3QH4WROlO05VvsYHwhOh
y1RRZABotcYjbfD/n1O+qwx1cY/AhrJnDAdLn39e1tyOf15K+NhBDPCxyKwTV5TgCWsL3kPEZS7P
1xlM9ZDt7oY1sjWcMLlD67zs6YR7dQwGmKi7opA1GLJmaIlovr7SCE4O7q0mYNZtTw39DVLfXqMH
eHULnrFM3DXP+1PrhbB1I4UPwy/UtkE2VFMceiQSMtpo9xkwOIabM9R80eeZyzmXshqOfwFwQVLp
UUV0CZAJJkGvYJYcPvhOtUrrvHJDRYZjVTk43nDD/+YMZzaLs/S6ka+AzOCO8+6kZOGmKz2ur9ro
Xe1RTQVTu2/CMbnewP3KQ2WUhGRLDlGiZplZ3SrxjNHsKwPk2ZgS8Zu9Z2AbzOO6Q1gOPnyxB00L
gCrW9d5v7DKvi+sng9c05WT46dDS0BsM/Auu0sePX28gnlyxQ5/IAkx3uO6uvY9bOHnPngz+4qic
197JdYpVroMlbD870lhovO1RYCRndQWOZd5/388Lsz06GGpMHXb8F7/X6wQ5m+HjggYlY7uDvtK9
Kve2lJiVHZGqRkQpk7zR7263sZHn75umOKNllg93VOIkYvthqGr6cLd/MucHaKvtWDnu5rAzeYAS
p6hq3l3r5m+WFoXT1QTzAU8mgXfEelv7NbuLlY5y0FAkRLIEn2dLQRbrWfRBn3WW+vbBxiNbXhEV
IT2tJxyPZXaP4JLuYXczVJAzc10TkHkrOW9UDSuQCfuoh3pSaLXTUKpSGYAsjQdngBtEddxrCHK+
PaWEtkG/jZOGnCH1gI+bxZCvc4dm7reIwJVXZ1YenSD2DAd9cT1hJefF+yk6oDBRQ3k7vPBGbg4O
dScZTsOEfSBptf7bgfd7O6s9DQRc8ovxRzwSYTFARTVjreYDEeZJbVTpFj6PPXw7l9EAqmVn2Ysz
6OctXVXBNM6dx8b2Nw4mZyFmsRz4ElqjPRg2ilASX8jZ69pUqVdS5vYZr5Cqvj9p9QzDbEFj2FIM
8tRnrp2wMlgg1KUTAYHYwRpfGXGTmdTZ7sI5CjI2uOI2pv9dwGsosZ3mD5RplA4NGqUtBweMVL2i
GjvcfI7CZUjqbscUqRSEpelA0D0U0RjEHOuz/cYNTMsGSmNRlTonb9hf0sPsMBhWnggvspWZRm1m
f+VqadBBmCurCXpwVjwSqDegRaAVK+9MgLQQvT5L42AaWhu+KNXz+VBgPTWX4E6UXYb5CWEtxuOV
wWoXdwyiqhmjwKBYdJc8+dvhhHkf6YYH9NJ845bxmsXcCa1y2U2qYWQDd4Y+t/fVYD1nrbo0fZU7
PIuDQwbIneC4JhtnuGBIWCd9epezltQDFKjql0R1i1M24he1GG+Y5VHT55nH22GDH6M71Zj20gYl
BqekcRzTHKaZ9MYy4t7aZVsTJDOnNjQNBMs5N/t26PXWB9BsRYRC0TjXZZMy13h0nhNvpyfECwxu
rGXK3aN5T6ze+uakwSs4pGV5xk3eN6dAktn31T+UJJS2J+PIXtd3Uh7emv/+VnzRwy0rPjcbMAFx
VQf0rcnAmRX7O6V/PM5UB0tQ5s8iKzx0j2d+9Fdi4/el6rF6WPpxTnNxvVqabKiIcUEG1s2ToI1G
7MmOmp6hbk2EN6MIWcDIHLSBwloJK1501mkz9l3fkbcgKliNGkIUI7w7D2CPmKGHdxOC7PJKNsx/
XaNXIcjzxrZ4oya1RH7eaN4NViBGdVYlgcbrnsSy2MNQPMnK129txeyCgeYpItd/+DnFDA0zNb4P
qUZnP3DhtEElhdo5w517qlM0iELOFg7+N1932TaAOY8d66GFH7sRXOcam2yhqrbx1bZ3w4LJ9yL2
voIOWB6lcOByU/KkiLgYCCdRv4E4NiAQ3JECZ9sRJk3YgMhsNZZaDokZWOvzHli7E8ZTwdiJ8y36
r/Mi0Flj8FbI/xKFZ/83rxG2zpSSQAVHr0mLrRspTuWy4qMbSUbIvSfNheGFZ2QO7YgKQnbqvTVl
e4z4WmXjAtAZnh5DgTxgn4xMw5OVHQTdtgNm1TZjM53+Tyod51ca+FaQmQcj/c70dB+8I1SHhtcp
XbZc+xjXzAUPcDeUe5qHkldbkSE0j8SdpV6pBE//Sk25FMvwQhzOP4nEn1yz0vs4FPjM7O+S0ITG
/vfpSkEDOlRhSxFpGyVSWA8jC0uq07SrRBKsgNhOWq9RM89SQmE+3Md+7JTz8N0wk8ZBQMlxzUgv
kHTGSsUB9wclIUBuFmjeavDV5If3PfpCpaWLD6l4tKEu+xfN7+OtQnZWbySfy/7d7BkSTHTcK0Vj
wfaWXkYrhJBh4ahZE8UdQpNJWE/HOSKRvUdnw6QY+bte4iQPMS7tBE5IVCD/C5S8/VaUkMiWb4iq
rIzcPyJ/F7mNg36CUU5PUIpvktpyLNfwCKobw0KFdcKVbAc34uLH3x9GP9PhThbLdhGc1/2Ntt50
xqL1xV4jOJGDmOEidAwBTQYcw9cmoyxBpkxzGdbllR2SJta7Wm7nI3Xqo4p+VL5C70b6qQgi52SS
aCg9QK8FcQbDOBKTgtqSjOxpkuZ+13GAPVcruCNKrPoskxy24ETDHciaZbiT3wQ1RQkSNNLhsA/r
EmO5Zs9kK7ehEknC63qDPnockViPZCtI23j5vTlQGldxMO7NTIpJTVWe+nLh91STgZVksAsmOUIX
8oefv4mJIiIxjNaPtOl+FfIYxZXwH/Gbq6sPjkJILJ937irrpCXv3h+Kncd5hCZkoLqJTn9u1G2r
giTA/PMLqiTFCvXV8Ora416ncLJh6hCayII3wKvyJAYz9Rfj5n9nSBlX3UWE8yFI+Cynsjxy78Kd
G0CqeZoRVPTFYqKth1B6sNHW14+DqWnnOVSOIP3Q3wFNt9VvGqOGexB1Y2c93fenwEAfky1/B/1q
skqPbBzZlFwAhZD5QLfFbDIcTXuvhPAz1fYL1NUmwWcHc/36D4cdwpQPCW3r3zByFpHPSJiwY/vv
vtS6h5Vv9sEy7Ay1i055m8q1u6l7iPaDGPtFLB16Asgv34pSl7O9r9X0aOoMCJKRCmUp+6dkFBba
Ycgvx+Mb4bYf56GUIWW/jvZVbEB/QwqFTVt6okWYOTpKTXk/V1PnPZmjYO9MI+Qplc//IE2QaDYm
CdW69I6UmJnwB5JYWfpRvXWhodV94Kz5x5flIyag5EgOdeh94t7Ii6vezrpfX2ZeMT2VjMGRXGs2
uxvacfxfkys8P/sDcZ0VkWSCaEPXo3CffANgJAnJ6tdRurAhsyrY55BlCEQweg3yjVcHYt1e0+at
s3w42kFEw1nZDOSUOxHQ5YmBwzD1QGnbtsKQyjSFOT1YcuJv3FwZHSyHiAHn7/DRdh/Pii7nBQYt
QASz5HLd6T7U8BC58qKyYW4Z+cx/7eT/EeEoxCZsHi4E6XTQIpXRw6u5PH6wydi5gbtJSMUhkBdB
Lb+gZMlyx5Mz2m/+CVk0Mi9a7NxuwSSCrVoW2L7EsLQ9WLzvAZmChal13XLlbiQkccO7LHxRU5+o
KizElk5xEWc7XW6jEfG7VUBObEhv4BvbtorkvjauxcLG4OZGv7/ag8k20Jb7yxxQG2a2OKcdNva5
c1mTLSloC7RhsnmpOSV1RyQ2I/wUqZCrQJBb6c3c0HXxuM77Mcx0KNWtZ0zdy3yI7ZAc/iiTfby/
K8ubqJ5ZSON4mXZ+uT+eDHnPoiFDjV+l5fy42P+ENsYsU5OrRXQD68J3XOueRLskS4os5aFrm1e2
WP7eIe1mu45jwbUHWiMjh6AL12q39FO0RTBBgJ3J97ssnYSLD1JnByOfHupBA/BBS/x5T1OkpUEu
AlvXp11G6EYfyFcNDItOlncVbPGtXE+jke7e6yvKRTKbe1m+T6MGCawMtR4YnuPxezcF5oydrEf/
gksvHWdy1xPsxDmxk7oJdNJoy+Hea2RjNf6JNysaz6oXQYVzPNIZurX1dKMuihNHV7z3SrU4kchf
OCEqQrNfPiVhdZ0FG6EAqPDUpY+evRcrzIjvkM47ZMQ8clwsdrKFIK+4OLQjQghmcG2Ozm1oBqi8
2PY7QKxWXPzhaHWrQKNGktd3Zb2XRjZAPuBwj5DM+NvdY80+Iw8KW6PTjFW+TyH5Qwcf5yZ4YYwn
DGnUJ64udydXxHEpvOLeqnb2pkOZZi8DhP8VQkcEJIOWuvSEXZKsdq4oSLc62i5FoMPYlQ2G65yX
WZL76ER6l6OTAqdID51/0gc2FssmP05iwrqdyu9zDOFQpzsHB5byvTSrTP40RMesSHG9Uh3OQW/X
42I/vmcqv06QA4eSLgnT2K54xH6uwv7xyKGKFZE7k+BUmmtVUp+O89mgL5fG8R5YoJEjw8be09mR
fbiwK+CFzSt8f/j/i9CkZrxfoHNQZpoFnOy2P9rW/obo3RpC+BKIRE7O1WMMRFrCCrNa7es1nQPD
Ddfmsm2ExkhD3nes0Lg2GrV5NnhdsTJQ2ZTs/IMUWSjcYUHJ0xzn97TEs/2mShz4aygYf+qtSIdl
b0/7F5zIYCoV5v1c1SixJJXkxJqvQYdj03soXG1hefs9pCKRnC3SU8wwCVoBZQEPsK9X36BzSCyi
8niq+C/Q7+jsShX0h2SEUUP30nRSn0Pyve6NuGUwOqG8XQwzwJf9IIIHJHB97A3ZBUsCJK4GYJ0U
Dn/Ud3YthILgdGVDnxAc0QVKRQCnvzzHKismIRWdnU2nykY5DiS0XQnqcw6McD7mqYN/L4+AMDFC
OQV62NYccXG5y5K4XLm1QEUA7tf/DwMkHlI/JVHQ4tD20cZUMnqFfBdWJReYVlK66oI9dWt9lIXn
yux0UIzVF3ZEbP+iYtFSf7XkTItB+vZMj0grblJW4OF0FIzZmT3ZUt+2uWSeolMdOusWmeDoBjve
NwAsCvTUva0/kI734kezrjhF+ofUr+aFGkuT0tT3LUza4JxhuHR0iZJWsk5ApUjKvyGeu5SkTTaN
BZ+wm3dSHSgr/jeugmneKMg5BGjwgnJVammeuH3jqpRPdzmKmp4VBGHlUM1o27EjLE5R5WQVPDzs
FfFdlaYHM1fvRvdj4x2H4hbl7yraVNGFn9wwS+zNKUWFETS2b7ieWmrPprddj/jiUKljAdLNzgp/
4VGj1FObjHEkfHuqylVdlGw7EvMj5Sm+jl2UDB0JgxFZ35/+PST0SMdE8LKDMnkRGxDxh0Yzkzzn
ilrxXdrFnShyV/2cK5a7mvNckTj7stWzLbQxG28jTQm++qmEXNwz2dMyT7YFsimMae6vTrFZYXTG
8EObyVdMCHh/pmZ0qH0ZOddclL0Cm9qsBrdxtHzLTunpgT7TGeD5CtxIE+HXBPywHDsuZFBQe+Qz
jdf7ole3udYBNhOzccPPDTGq1X+21GcRPJMuu+YzqAKOD/BXYJYi1b/310QTYrTqnex4VDWSCJkX
5/Wp7RYn/oNV6h+RcQDDFBkVXnJGztvgkqRpHsHIYAWaDPXjboCZ0z6jXbkY+EvthBWzW/8n8jMs
nnnxMUvxC8t1kzYu7WDgk+Y/H0GOv+Gwo+oy2D/uXXg2vGz6BwGHQXBX5ok/rPKaAHrkZM0qHzdO
p0UTDDNWZC6BKJnJlgaExHNfHy8uSnI8Kni786eUzZwu9tY1B1iTqZFwMgFehHefCew4Jreq0ftF
nkEGzC8frSZIWMPGW6NoNrxjeWgETumrIMbnhdJSTpqtqgW6mnq7DaDL4LbaG2uhqeYv6Xuw9CeL
ddEoi4hISf0bOcKYXYe2fl+KYXR0es6gctVj9qaFAf8wSki1v7Bdy/MN7iHYSr3RwlfY6W6+BD05
FO4AQNmWKL/rb+B7BL64rEx7isK8HtvHqJlN963Geal4rlb1bIH+9Gdq3Ra3SQasB3fBRVxU0d+a
mlfQcgagnFOQ7th/HaqP55J+2f/+ouT/L9Ijvfry6ewRTCLT6nBKqamR/H/JOXNdOkG2/PXgmhrl
zGFLefZKFUGRwFQtDTvtrRt4NDBF31ARsmao5C6vzcEVMPOG8P6LxRGCrsR2Gfe0gaDWIb1BSk5L
v3cZrQPPMQXOB40vvkH8bCUt4r3E4c0TIkOjFa9AtZv7hHdHu/C27jC9BgBMyXFAIj6TqnRqrkNR
kXDoKPmMM1VXbga3perIi73oJvPkJqLSS1Slgp06NSUBMKFlgI1RjPQlORGAPciaUZCvl7bQmloN
HQ0eom41fdosXixLRj13Ik2ok964BPIfevbz0NTT7/2U0/Ennk4mPw3Ma/5C73PMU/RxDNd1RPpM
Yp15x/pkCNxbDe78IXQPQEofyeFRHokaOMfRkhlarPYVKg7F77EzN+T+6AgH+Y99ILpdLvOFRuIq
axGznM5QQB/KwXW8CRjikQNg5ons3GVKtzGE8Bz+/Eiep36yFi1ay2btt9yMShCiIFCXDBuvlnQD
K17YktbihMSsAjvT6xpgSQRXbIfHqMoMcvi955W1FywPlscMXytkN2AAKEFEwXrNirQQrZhIU3BQ
lHhmnEL9TCNgJ1ipmsG2BB/1arSsPCexl6Jjl98StjITOVqPVCTlZAUTnoYBI0HoTCf5jaosUdLG
LG47JOOoXK4o3oD4+Nfpw6ah/KQzRapV4eO5H2C3O9kbSzoS0cSGRC9685z4VGlW4iAijU6dktRV
H+zke9F6ghfk0oYXMXtJZ3W7wSoWGr1jOXPCwAwh3LRsKnj64wRLOcMr3pfAKVArjhDexEs0HZXe
T+LlpkNYUgfDuwfGpQcoWrRVE3ky3+Ds4PdnoOv4TVNPj9J7U9He6ASogNA/D/HxpwlgsPUMW/32
DeuoM/CFVsud8BVXHs7lUyCctHIPjMCurSBccMM0K+cuyWz2CM0S2SMbZHdFTbLwgTqQvSx4V2+9
GDCEPUkjzVdn16MidLPlkPZs5JMw/082v3kHZpRxz+2XskAsWY00PZXgj391bddKi74QkvMrugVQ
X8LrZsqyUiyeUBPbrxpZEt8CGUz0M0FM/bQUhf7zh6b55oXrpCRAy+UwJ8zBbqCeMjDKD1iw6KNh
UCIB/5vHJWEhdtx5UQzX8mMyR2/IcKNE8UDCKkgGjsDo9RRQ+BfAdgSF+2Zyd7tzPbFcaKVHWKSM
rAI5xu0+E62RrhlppWhQjhDk1VpxpGcJ42REby2bu/rC2V961MXyxWvF3a+/wX1d+4A29q0rIlX7
8UCGXyJo2XiyWmcKdio2aJEQOe8V6E6TJOaTd11/oQ8xSQ4mVDAi2qnb9NJ5CulYsNrZtLJ6buoa
/fWJ6Jk2InF1bVLFvyBszJVNB2GT/IL3UwIKLg+DaWwvfeopO6MpAwcCw6zjVIls0k9HzsM4892d
+QV8NeGKvR9/qq/Y/VNbB8iYwN0h9pamm85JzL7eepRpyfZH43Kk6iSUsp1GBEfuBOd/fEJwnS2P
qGS3IV/EZbewM61BaFFyITIPfBWCM7YVgmmvGXM4i8IvWA0HmV7p/UJ/XG6iJd+hR+8KnshuhEDN
q0MYZgyqCBAVLFKaVTfPbakAkUauQMgyE/LsjakyQpQzNkPn2KoKGf4KgQzzdzTzaEgxugvVJ3Vd
c2ppRF7yweL7tw9qRnk7gx1yThudRaHtFtazFC4sQS2ABFXjQbF6G10YejyLY5KFIMA3mSekKJcL
oZ9t0GTuht4CHxWf4h6en5M5MbdCETEl5tU5b+EEO1h9YiOc6+Nrbh1NYhnrpV9FoEhSbdL0NGwW
p3W6tsmye6hhoJ+Tctsx1LG3cFgu/iCJ4r6AevBWkAXb0t2k1pFhEJdDdg1Bl+yLDi1eF+fqKEpS
ddU9PLHWoLfFPaAI2RyMDiCBCpLJ4Z2FUPlxnqDILTwhG2yu2PgdXcmm2y7IyhjH0e5quYReBzkp
maMGQ5XIEv79Kec4sZ0g9OF+mvF0tyYClallxkpyDOLWMRO7I3qbWoj6uSlLLd/RSOXJhdJY5MRE
2QeacnklqU4BPV38FnEfB4+pH8GHckmgA/VHzMYiW94/cVPdrOrTa7UfV9NYzkb/12t0V8GP3C93
KRZE95evhNvqsfqKa+hwVR395wmD3mB8olfahWWAQIOPs534npPoUbN+5wPuyJYaTICd+9zUh4cN
EjWmPRy5VohfN9zZNy1j+TIXFb83UqnpAvWH6Z4tsOIMlehJUp3kC8phfq+ROpQy0MuhzaG7y8dH
1Z300MkywYmtCrFe2BxRjNhVvqXlD3ScDfspYOk3sqA1EGOcAP+Y6WUIXi3Du18MTcDpUgXaRlko
p3pP0iAYyRNlJ3DMY+kbdN5sivkUqW9gBONPWP38QbeU9xagV9rTdnwFw+E7nURDS+ePwJ57VaIZ
eeE3MDI7AAJDxu9O0E9ie+Jg4wIFtPMJcFJlfFMcYqccGju8RNfdfa5dDL65XAySPnEW/bQVMoZP
U8awJ4XhSN8FwvXRsmlUj4AUdQB/MeoAwaBt8KmKmli7cvWGzdl9SPfXKeQTgEeIMBc7EF0F+vnN
3A+fVWejrKxqlUn49BIJtXF5Luo92nRzaUHryqqtdIecxY6tHk46zGzNr57+twH8YADYKo81dJJk
vbqdIyNQRkuoeDrpgNK7L0v8ZQ+KvWX56xzUUtNXCf0C9LZH62JMGTB/OOAdDN2GIKIcq4OpnE61
887uqQzFUy3oVJFD7sMbcls/Shy2ofcUh9A5+SJ2UkYFelwJMSD34y5cj6sr+doP9g60aGIwoMuc
KHjQoHPgQLzaqYobbgX8mV4mnBu8+v/zjGsyBpAjjx+fMoP+9PnI7qOO0PKBdVD0uknuNWAgIf7X
kCABfHjA1clkpTV6IFOB1NQlWWZJlKYRj8cds9HVK4SWYkdFU6DNq0gCVxPCtTAENa1UxpGcOY5+
SRYJ/bedVEY3RXLPDrnF7A2SIsgnFHTwThG5VfEceNmUgDeXiXeeBPa71PND8fKeRECPUGWP/fdP
9vOytjTBUeJEjGmxRGEG8ktysq7NCE0vjTBCNA+JwxQyu002nd+Cc+ieWbj7VICN2MJvX/QCZlNz
yfOYjZoNY3OgYOMIq+VdfQACuZe6LSchYGTEYUvpDlvqvVpksquKoaDpKydVQEEwap4UFxKTcCsH
+kjV2SvJgY0Fx66M9T5OsfmhXKCYnFPd8JPSLw49L58Ec8PQv85FyKNmbq1VKKh/s/nZZ55lYtIk
vfonlxlyNc0R4Z9u1FkqCPBnO0MNW2r65GlLkWZnS8yrIQpM38sMPqftk7E3668Dw5Bpa1Hk119B
UQpxTbXFoVsAkXO0+smDuSh1oLKILoiISjArzTQvN7Zbc3DbVoQNoVF2OVPPYiJEg7nR+MkLXsjp
sovyaEvU6zO8t1MpNxQ6vI5Z4hh21aCjcXd4LcxvG++QklVbPKKPOPJ61L1RhM+Sz+qE0KuRthnc
kobEj29F/fG/3feeyyukDufqPwFNpdHiqqGLYyudilY0hHQodbLnrB12N54eAGMvPQPcnZI4pB3F
LpASR2zvv6nXHDxAF4MOxff8wSqYAP7ii/or5DjVNwx1WrhwGiD/357fYTxZ/93AtUsHd1WDwgoP
m/xR6XAOZRnFk/gIGUv9UDzS+6gy/MvGO60HajiPGCOvy8wUcPTeKemopGeU99/dtq0JsOz4lkTZ
eDHw4a6JKkLjYG4wL0Hn6kQKJ+dbgEDi1AJWmtdV33oX/N28lLdUw+i0jlCzVxu0yKgbozyBVzvr
Gh6bud5LW1EKlavomUnYC3omNoJTX6moLgThxtT9gGKOh9EHA2sq5NdZ7+BOF2P0WcDy11fMSD+R
pDEdEoSY1yRxBDVZBOtESPfK6fDr0stbOB+X48EutrBNFCy8tEkTVnXt4GGIA1fpkTbefkIOJO/z
oYqDimwQ0sTtYhV3KBkqUJk5vu7VcXmRe0yhzfx+uELBNm4NR8uqB2XqV91pG69bF/r6UUYmJzF+
SDjxwr4Y+MIBGFW8Un3VLvaZuwYbOZ7e+niCK0/HqP6mOHJvwfzICzRfKrJWulQHTBbJKkQra4qU
23Xfgbf0tVJQTGrtWyNIb/B84Ynu5p0xuUqb5GCJ8wmQ0nfHaTO3izfILv7n6OfDPtTNbHY6nM4M
x0v0GF6VRxlDZFVaSHyF6SVIIXH4u7SFtHFLSK2SIuDF4lQINEOk7ZUm+6+xYuPwF7dEnZFRuZy2
9I0OQOz30oSTvhlUz6AYNLB4qQPZr5WLe/57I+Pkke3pS8Yq4E43giYM/nGA7gP+r/+tRKG8sh2Z
JkOr1oKH9Fz6DKlOc8PhzZxlQMxC6NPxMbPk6C7bAOwayE0gjU3oP80DhneM+sWrC4caiCWyjy41
9I3qB3AnCI8rdmgWr8p8Bxh07tgNGmeeRbbzAzhKpSlgiWRgsuqyQwM9MFZd1QAsDNURpEYnecCy
/zRaZ19KWGuQ78NVjaVP1EL1OIWovXYw+d6+cTnjnz3nx7D4yVSHnGbW/2Jd9ZkaiWm+01n2v72T
gb5vG2XAg8Pu+5DpiwykfJc9Xd0aDMF5X9NWVMtE1s+8WBTkEv025GX7lBjsb4uHrI50mvVCzQrf
ptrI0VPxPtvmArJpHBzZ3aBdY8vuaJU+ruBzBdGdexIIC5fxYuW5SWkiOK/ssGgRB6urkryRswmO
3WQL79g7vxQd3kgwC4Ib0fm+o9cuyz1zk6JJhSGzW15o7TR9EdB1Ckpgxnq+LYPpf8DUxCs7JR1u
3IHRKrWoy/TDW4lv9j8B3qBpOgz0msAUv2CuGPrbXlatoyVlupog1Yo5Z8uKFIDJO0/YpVjbSuxD
Syd3AyIFURcYg0f6cokSliKZ3PQkNvgx9wMJG/uWEtwQeXyJi2dfbRA/UUhpxp7F+7LT2WMb/GZ2
18F9quLxl5eLQ5xb4FAoIkgS9SvmQKAy2oqZRZA5Ejo/wGVPnIZvZ+kL3DOy1nzBpdwkFEXEZns+
8KIqQeqKWodEXctmXTMfYQMFXO/HYotV9Gt9QDxGQpVDahkYuFZyonKk8/xhFzl9KnJ3khOcklAP
OQtmLqnIHVm8mVQ/b2ggfwJa66kvgGCmRxL99as9w5Q71RE0pE5SLQs9od2+nDzEhwZntsc72J5E
8+HgpWumSedbleAL+LMQWYQe9qdz/afRKeABKJvM+vsEQjfRVrp4zgTVj3QM60+6fh2J6/lDq5wc
HyfcpmjGiQ6NFc/+RFv0nwSoue5SA8RDyzYxVz1lYtkGhVBrEFACDRvZ6jo9GcNuGs6z9/8iYR67
hHiIHuljEcZVCwNCqOLLrLpCQb/w6Txw6Naj9kwDMbee0X+m3CGBG9h32EYKy2waIR4g8H1L1R5r
oP1D2rxVSsTUj05I51zLDWrt/IAUgOPF3FBlGLB9jSGgG+y2reuhtTH6Qn78yoM2LrwK6XJaC7W6
4y9qdRY4hO6AcLh/9JtDiriCJaw4jYgMMarVDy6P8KWJrxQFZbtEBNhMLc/4oX8p71JRYXnUnDON
CpNFTbqGzVwxJuw9X3WnSdTqNge/9bPytuIy9cF82v72loBkX8e2irw6xpGxvC+IT25glsecQP2i
qfgzsImLAXaSdOZLimOlLJyzpFIWPZZ8UiFm++ymZ2/XwnBsUMFTvpjUwam9+4VGPzj1pE1KrBTW
H3VscPgR/2IIJJbnouM+WO41BeqHJG8fJoGeomQ7UxKx6qDKIKDSehTwBbApZelJlQ/vWINBenYk
/xNuQX4Ch/Z5DwI/bGmXflLlOJH/0lYs1o1w6dCdTaKIXqhOzKXYeRbEAjUsccjyQ0DRBI6SfX49
l325l4xB8NQww3ikHLYUZ/OMuoSwDcgEO7V13Meg/H/xsZuqCAK52JwuCU7kfah3xqPUR6joFzNq
zivrYkOUVjhu9RyfvLIdIAgI0vQ6UuCinStZnCozDGyrgcqiBAEpWvXWnDL5l6Aoihqca72rTNsC
n6er48e5OT/OTNySBGe0c7dQ9I/x5RaJufedZY5FGpvL3b5hLMa8k/1ksQ5qNdmU/Y35+iH5gKRg
KOyXWw3XwkJc+3MRFJ6D3U17xvZeYelF6cWUUJaet/l6hem4Kpu8NTtiK2mSYw97+13YFokd0yZt
lGFPEqyqs/f+XcZit7BCYuurDWkqBprhWRZEh8VYXyDH7wNco3VcA27V6S1ZizibN8/iCgv2FwNF
2Gyux/9I4GE9Y5P9XJMjtxsk3ZONprGa6OOTiYzKhe43F09QZ2CNn7qazQvkFlFWZFdtis4mbUiF
m1OxJkl5GRzvrWo5oN62TIwyXpjdkSoHX0L3/mJvMp3IWiA4FpKjtw8ENxsCrv+ndh4nRtXQ7f3i
PzqWYqQfrKK1t1LjhLJkR2LoHLWqyeb3iEBB353mZ/LoifSSU26L14Nn8oL6JxOQL2CkkcazRJvd
XssDK33F+lmtbzi1fEkpKyrhO8bht+h6LPPA2mtZbFixbAwDEuwLVCv+7avD9TR+iQeYziAZEFRk
wCFjGjrY1+ERCFSJGcj3esAwxxFsbI7LnA/xq9Y1VBqPF0R++ISBz86JXN4Iff7ed2VnOqcp/ZDk
0LjwXfy6EmdnQegr97YVnBEHiSZ0xuwmgZDChLbmuBdB7sU4b7ww6urWl6mfGTJOlpGFRwg3XhMo
EW2PSomEwE/dFeaFkqz0XGjRYyjotmomFCZRmNSn5yTFo4LJJUo0IWfSEN98kUnc5zAgMiSvpSlU
t+l0qcKsieHWiTTNSyfgMkcCDbsc+J8hqPHKHVa0YVjx6EOeAL4REMWiY7Vxq82WAA617RMsjUkB
5e6SyAI40/diApLWmxX4N2Bpnr/Qpg9OMPAkKJmXBwXSlav74aNWa+GwMPVGN/1rUFar8rBWELpT
f9C2dEOBG1vTNTfhDmH79R1hePJ8u07pcAP6BNkl25nRBag3xF4iuvbI9Trs8yNb3jWyA+F04bpe
i1t7b3GtDn425APz/X6dXxm5O7BQsXkMmnJE0wWmnwaJ8nC6kfxCtOVPj0XTpS3R3zygiU/lkSQW
Lub7A8fYJxeAnmYLwkUkA+Xwg16DJ6IBoc5+Fx9FYxIpYiZQsVbSSxU1BsB2kQ4Jun/QAbHQK670
HJhLTa8/rYobjwr5Ppn1IsWMN8PTRX1bohH0MzGUsiaLg8JQC6rpQ/LIG7mM9ue9O28HyYLniM/R
iyrs5PRcfYD98oy/BCTS08BDzNy3D5D72PdDVOyKMU0VsDu2U52v4//eor6dqUzrjMt8J0NJQn/W
NMeBQwXWs2Ow4DhuU5lKB5PrEEtAByzjf3nkW+11C5xH5v1/0I137Mm1eqDf12Q7eJQom6ox+JnK
oy21/CMVDKT77vV4zKkrPNlW9k3/aBJCN08CDzs6FsYBpVFa6TfDMUYkWcTh7f4/Azz7Nbdwa2H+
EbIlLA/N3c8NIO+gJx43pKFhPPFk11UUwuaoSM8SLkywQgDyezEIO5JZT+yvvVcAn2uonWNmvMGJ
Fu4a0D+sVDO9wWkaSUTQrZb68gIwmcPt4Rq/ohwmisg5JvkDNPLK0EGZec88Y0a7ksJ2t7TEJhi0
sXYLy7kSKypW8dfHze5RPd1ItrYSf4S8E+3YruHOv5IPGki1KKIIyXxWCFRhG2/v1YiwcEt6a57v
auBEVo1UuMzllmxMsv8W2rDPIaxZGYiYPRpsw30M7eeYCos1AgU6FepIngAi9B/1dPw+MoqCLUT4
uM3cAQJhTE0wBBnfHwCOX4M09warJ/Vf9VD6KLokpxR/js35e16ZOLlYbqT/qG4wM0VDLln4cvGF
+BpInS2ZpldkSVTbLDMjxDw2gUEx1dqbbWmlVdCUADr/mLTtQIcDv+hkuK9vskebb5fBLs44zq7/
k9YdbtIMRARiUXtBWWUfmY0R/05xth2IY+7lraSIjihKGKfTToCMm4x0I3Zvpm7Xb3gm3ejXdcZV
OIdsdgBXSoA98oNGgl2xNryRodOfS5DFVz/I79V1mN9u75hvxM/udrCxz+dd9xxn5vppSYTf6o87
toD8+0/z0E229bwGZcg6OCVaC/7cHngqc1ScfblJ571ZvZrKxlz9uTpWaeDnVKEvXxlG7aRn9lbx
5JroQ1+cBqfvDwb6m0UYLIRNh1vosSprumNY4N7OkVgcw5QxzaFJJowXENN45S8VJOsuEC0ln0Px
x6h4+6Sxp0ft7pvoA8VmGqOcUqwtWjyvvLSW+mjWjImHCdHZAH0EosZauRWGRqMh7w0jQkDQnIpt
hVnwj18kV7Xvu3eA7iZHRowCvb/GoS3OovoFrZQwTnTG1EA4eLNBhvzK/4E6sv9Gfh7uJH4AdK6f
WboSoZnj3FKmBSDIDGmJ1hHNlractfHdeelZfUMmQYc7xR4vbkg3xuKTJhzAShd9L91gzw6TbIMB
w77HdRcESJf+Ap80EmpX8HFTT1aloVwQ6a9CqHqWmAHsmv79yqsz7T18GQo0yrPkpBox69SQrV/Y
e42yX+AdMSsaMB85z7QP2Xr4huJVvh0CayOX5YU4oX+OPcGyeNTDortk87F6ju/sQHBe7QSVCRTJ
Rah/jjyax6BbnvMgngHftcZPg5WBYsv6aALNKbxYGoog6waNurgYtV8Vv3Lm+Edlw7i91LE1CjUD
bcAso5MWoESFJkR/QzRvap0ZMxH6bJHM9IbGpFsOSAErCuI3+jaFi2uwbHFx2YH7toaMaKoQMu3n
9Sl/5YbsbbB0V1rrNksFQ5TnDXuGJOSCnwxUOpdrQEwhbhU15ANbgOqNu6wV9MSZhKxac+9pBGT8
rZgbAlliflzSu85AhwAmO8gXTr0gIgzfcTbyo6dLKXnzVQGm5VjzCCLqhsCn2VMtSYK8ZiS9DQ4l
rgyrzk+swx182sJF3WDU2WWV4HuF7iIyd5taZp+h11TIRKq7z2EIz4N5bHyE31QT6ZkP5knYBYBr
gXhTGU+enxTuZOZCNWQhC8+PTIbKk50O6UAfXhgnFxwOl34053pgoTMRgWSyNHe3L4+FPmGWuTZL
69dLXjf5jDtYUXDPUJhcsISjYuJkXWFMgaLTqny9OBwQApkc+V5zHx5fSr5jvKSEqV5FSgo40GPT
K4sVRZpZ8s4YkSSG9SlBDG2WHgqsHNzGio/aMTQl/8K0rIZacH6NClaLS2qjRK/pNAKUE5tvn+1q
NzsbWrTSANEgkFkFNHbweZd+WiYaJ/K5SnzpqF0rEGstSCz5W0e+Th1kQ2wZ1a/vAopZyEyUUghs
vcPxG3H2Rt56aB4uXqVN7sXLucs40Zh214eKqp5Zd5+gb3uWZfsb5WZZwyq2Gx9WO0uK3a8q8GT6
fA9BtqVP4xlTyGZA/UqcWvpFhhv5oXzsN0qG9gTn5ruTQl5Yg4LoSw5mqpVahO2sy8ACK1pPxiYa
ZvUtpOG87fFu12uJCwcZ5VN5RlSXUHXRIvguJlrjIZ44Oartwev84bjcVNYcbGTObM/3WyMkg+qT
0NjLsveEFayT7dX6+APUfkyqXPegoiG9EdPBe6R73xst/0Yc3AzHV3dINFcT0Y7G81XqQbp+dqt4
RtDE4uZG6iBBkUkDitZtMCdBIa3VhpiXVJep5zN9i08VgqqwEiZccWXor88ZolkPLnhu+S+X4u9P
rKQgN4D0Yt5T243ma+ERivr4VG3mf5KaFCsvh3E4VkrXsVAPnOWFKL0MUxoW97RX+wvseR0Lw60V
OWcU/OS2KZRnhqPCmo0HYx/IcQzciP/pQxqL5pdMxwM6M74Bn8sCwEi27Cfq6uW+4icBlCJBCniK
VmHxdD/2vFfzM/HOl9v47Cy4EpHHHUuzePWLhQNKvNUcESFkTf2N225jEvJVu+LyWqNd5SvYtiUD
59odtnI8/puexfHkQobVaShyYCyT/5CmLNDJqlTI0eUb1HrAq2rSKjN8aYBybzPIOin3VglHk39h
Clp0UoRdSUZdrPpfd0F3Vb3OovTyQpORNaHEGXkHawqqvu1wQho1wj+2fdx0/kWkSz8uHwxeqkzp
GhPHWGzP4NnXKeEoD7fkz/l/mfHCSJPWi035aVTk+vSFI5BqG3xo5bPOsP6cgsEczv82oVCsGBfI
tlFc5nZ5bAaZ/8W4HweaLA5W8HqjWLw3nqLVHG04SsmjsJOkDTBUC45dG5V8HNty9tUoB7Dg5+Qc
GHvrOiaoROA7J3IUZzCQ5aYpNZURsicpq8vR97JppIw6X7nHWcZAtTqnDBgJfJKaTRCH8KLyZkiE
8HJTJTVr8eDmKdjO1Q/HdwyOPHsMmrJRbrZGnupqHBwJtNyhnoOSyCaqENaEV0CVC4ibJrNvkFH0
l13z8De0qGy8QRvijfouF30maXNf47muXAHDHYYLvpts8qX0r/aE9U0qiapdQfNZM4Kt0rSCl6Lj
etjOkj+srkJxZakBt0xuVBx2dEnSOnd1ZbNd3PWxsnFC+e7531KXu3c5y94Hntl5HupwYJom8nbM
YepqmHBlYFx4IxDRF6oOMY5MK81RHpmSVAQw8qIa8P9Jh9usGjDigtNbwsPiGcuaE2EP9vON14aR
s+yQzBbyM5PggEhQbfe9xI/rwbY+75LbzGwjwm6qoK0MdgClS6gTjevZNi+nI0KU9P89G7e9+IXN
JRKWPfzGfldLb6VPkJlui5K+6Biz7CyNA/T2f+vFA7BaEvvhxdpJU6cnrEzl0hzxDKV8ws1ROkaZ
11CZyHir1WiAbG/KThIgb2TrlR2RGxvnNTMCARjVp88lCJ2IJJL0OIlTNe2R1tNjrSlTvsvGUDOE
3NJ9vrU+duHcQQ40KWTnx+EUIXqn4GsMQEk+pqx4TN4Zck6Hi9sd1tjCwwjeYpygGOvWyVpN6tGY
G80r7U0wNX3OVpsj5YkTXzbsQo2+pvNoyoSiE1mscESZzxIw3FOwq8iTTiuXNQAWNxwsEEgQx74u
Jo8BR1/KcjKgM19t9yzFe+23o9tyGpy7dSNemoImg7qXvHCJf765o1J9NVDhiuSvO2yvH7Lg2NYq
qvo3m7l2DE34jSHEIXjkJSVs9tCJX/+Hiw/UBdND1vBUXeXPNPuakMKk4ojcSqnbRb93g6tlV3bW
DiBwXFNUu3w27jqy8/37To/UTap/wxgfSInN/nP/lpNIxmQ+QnhzXYRfqXJY7GCUeKtbAJp8WapM
Eq05q8O8u4p17U6qf1E7h8leldndSw4NsCQNoyLbWfFi5F8UpDoadoh/TI4+SEaqm60SAxEkMhGE
CSuAW6ui3qp/ZricmEf3D8OhI0v0qdFTHq0GxMyPI76bB26ayk9z3z0ivj5D2lBwQPun3wHhRJvQ
dYaNbAWp9BKiRzwe4TQ7TBQwt5IYGaPEhDhLejQ/Cnb+nY19iSQCbxlyB/bZcGqxMMgZQbvM17gb
by7l9oJBOfVbWZweOOqih7i7EaM6VrNYzNR44KGqPufSVSEpVevxjSolyUwENhx3uf86/e/uDOgR
eo2sQ5gF7FTxz3m80a+PEFO4KP7FCoO6OmcFOWS8K/taPouk5F66Y5wqTNNZVoiEsgGlTXLFj4t2
VLpUs1Fy64dQw0w5P6OaP3KHLgXRwlkYNm+KeO+McWJpuHcaFck+G8NYhDzeSGcD/5BfDZe0/79e
ReUCqS+wEetJOMGYnOIBe2eZhhiqSDVO3j0pCEpPK6i3HEhtgT7BnW/TuCdyzN7ju4h2VaZ0fbSt
ltXDiplmbcxfZMxHCkXsVPMXKLkUwrnj1oJigr8NQZER1RShRo8C52GcyIKj/YVFAWoQtQt47QWc
cTFHas7I3zj/b2aCDFdrprLTvCe3RyPsl/rVMEi72KE2Z08c92Usr1jJ6CVFK/b6K95DVj5hU758
tZ5AjEWv5xsdNm5/HKWp6WWt4TPzIYULSTkIf5F09D7vCevkLz3XX31287pIrayyNH76BEFsM/6d
lYEN87t6RRH0MpgLJjPAIADkmsEdDZnfS9AGBU2/5hI0nHwCsT3uQVAfa88ugSUDEyZ4iSvGkX1w
/7r/3P6pLd+nCrF/r7YRidAXi00GKhO7Bf8TAIMPCiuslBOOFRVFBl8/cGZxkwZJGbFLuJgEFKnx
aYYvhcQK9/NIL3FbJTeccnK9BSchsamQ7VzmimYQGjTdXGDUNHum6XN4IvK6CPJYQwTNmIoAFCS2
jCNq1j2MumxJqYNFZZla7a0UEto1NSw7Gp5Jb3GsNw7UpvO0VEozBGRTPAcwqnQwRqtsBAcVwPTQ
1edk5CJ4rYx3ow95AHD5Xzkvfkz1dqfW8xE/CtkckPVdFupoE+FjwNF3wxOlc4s1tMpK4nbhbqlV
tPUJocl61Eb3JcDSS0BjJBR8EfQtFOvbrlIe12HeeMDlVGQWp1V2ZiGRKascsdVReqblscnoPGYl
10XUxKlq83MoXHBDY/h6jAAI3dPkrFPoKz8lL99ABvWmcJYd9qCZ+s90sytZJvAaDhsMAh5cXfJD
MwhRWWHYpCooFt1S4yxNM8J1iP7E7mjSaT1zoseuApPSimKgidjiYjUyiVzbHKB9N/YWOEtloNnF
BatnG26RJNOsBidTPtiQqE3iqJYLsAMqNl8r+rcYeT8pw1rfOWUdKzp/Lq/b5l8OIH6uU04g8vkh
RJUBQnrGb39pKb245AmHCgpB6Pp6SrfHVxXzaw85xyECVTOHiTqZY28FhWEjA+FdFB5qhbPYZ4v2
E7GhmpJp6KCd1a06FZ6/fAGqoHXW041qnmwY6l29Xa0zhqDRBEt4A+huwdIPKG8H4xn1TjEhlVgy
ql28fUj+govoHCnQ+PGOe0FMsQAKlnWzc2alf8Lv8g7VpZUyRWNkK3kHFoc2Z5EzhK39IjJb5GQe
mHt2CFDIchJWY1vlRK5aZKk3ZfBGfLJ2ninnwhOxwOmLAfxisBpAU71+LROgWWx3cF082yNN3qLH
akFCXKWMw0RSyK/e3lSJikv541hdEBncjs0fkqeRuPp6FyakFb5ehjoCyiZMVY618IP6v6CW38nZ
C7LjKlQE6TdyHbBVOEBR/LxNsvjxaH2sM1KQeI2MXBJPgDTO225VA9K+tfXvgyadb2Qc5zV8KhMu
kP8TQKQ0t8B4IpIh5uf2n7eBbzWpl+2KjMwBaWwK0kilMGSnfmi+LlM7A+eM1ePzsVZ65RW6v29I
sWqvK2DUkVZfN4dCiOPZlqq16OWJaG01CnBGAi1V/gVHJiYQFeSRjElz7IZVGUFk8/e6f3UZS8Uf
QMY6CZjyUEko1J7kEYPpml/WjjuL6TQRx3qAmlas82vLjAioR+YCSkTGsBvmXORQJ6G9MT8aoLp6
sq53ADDD9dlADEkIUdjykn3zRJ3hYizH4/ZSud//qfD7+kelyV2KNBsGeWyDAjYESoBJZxRMjpFb
ITiK40xt9L7Xef+6zJ4n3AdpMZetp1UK446IATDF1rXq92/JazDFY0WIo2qIWQJVlN5V/iyQi1L/
cxtnycpqhxA9NocikfgBg3U0ke+kfJzR9TN1EU02fQynt7JErX/Ps51wTbd2Nj7Pc+Dx3YIKFgsL
9+27vAPhQ36C8GZzg8Zedg6oCq5uEgXgMC/FOA7Didb7yPjdGLrNrxInfjF3haPYF8GlMVjvJAhh
99AZC0ZVVcp1dOye1FbUGMh3Q0B4ti1x9ivLEr55mcvUYr6O/gS4nGDXI4HqT7PPgnJJ1fcIduGN
7thA/HoBvwwnE6UgXUBN/oanf1Q7nD0HGYwI716sZh4nmLS8lvE90EJEhfWWm1PORS9SDR6Dmh6V
aC1XCvd02QnBjMc5igCw6Jn5ZNenJvsAwITvaKxcBouyyhJY8a4VdArkf10+BeBGiPKNWbLfu5hc
a1/y5nSmJzUTiTRj16ITbMGIXBR5a2bpp54cJ7IMNX3KQN/mUYCYm8s9piz8mGFLcAEFSeHag9W5
eZPAD0VyfsCfsNjdsb5p2YTd6ce2u1F7tJCvnrRaUfoFGi8g6bASZj8MheEDva67hep8s3zlR7rJ
3lsqmB39rWqGa8YmG5XX8nzFxT2p/f3vQ//isUunzf3m7TLbKTBjZ2C+L7S6NB9iN1ukhtApAIOh
0EvPiG9kA22PJwrkWnWlyfgtzvfQDe2pbJrrmmxfBsQCNePPgQMS01scELsK2QIkItiLCrD6swhM
p6JJ1VqjXCQwP9rrD7yqzMUwjSvA0UfYvmL0j5K+nwUjPm5qiaQI7Wr9YVDwdbme+io/JYfVUbkF
dNHjtEMhJU1ULVxVoEArGCVXej7bXnVqrAd70joa2aXETAEgUF+sy/4STsZz9BXJEpp7GrD7C04F
J9g3WNp2FglwyAXw93QiMuBIPTMud7qZNKhBzR/8LLCTvFFkc12n9bAqi5mcIewwL/8mKuf7UZOD
htjyKzwDCMRtnOu8VEEWXUFKszuAl+30dFP56LzcFy5JBelfVMHYgjfOC9clWMKrgoOUy12vEm3v
1rKtJ8qfs0YbY6GP8pafWDioG1WEMOCIXzVKiPwlEA0mP2Iq0JEBebqlpGDGMXiEE+41D4Duo9YV
4YmOnxyJTvt0HytOwJXZzRQ5KekIORpm5Vse3ESocAndVqCemsNFXd/c1IPzBDn3iu7nM0n0n3bi
yM612aMZyFYq3NZUyk29f9sOmu19OCKZEaq1hglBW6uIFs7aB1B2BFNoFC4Kbmzy1mBbakuoXJuT
oKb6Gv9u+GAlfxF+X9PBPhexXi/DvV2pQX/FYCd8r9FfHrumzv1BirkQAo6FvL2Nlha57bXU16jl
NkXaWvHUgzp+nBq0mfiaTTlq9m0NoLISzkb+yfvgt9QmpK9dpDErY77KJBm4Tbi+zMD5g3IR0zln
E8IQJ6pEnydctj6uJooNdMzsPJeOpRG3bsKsGzgVPSdomsZOTXNOFjfJRuDpUskSHdNwjAeDNK4m
4UE+OiHtZ3bl893IvpbIA/pC9nfm8PqB58AlLWc0mOGongi37/ozpCfbtvkzm1tScKyJuDWnrKYn
09ZgKyToA4adMpbQanVCkQuMHzzBRoi6eBjDuEvyLKG26iMdhmYJu64Lft2+1LxViP2l4Q8qmA9V
+Kak9zQ5rUe3FjmPxjUN7FYxJBeNbiK+/yguvucwDCbLuPZdhWjp5UlXNEh+8QdtMjor5JMA/By4
OPVMzuRE4JEnJn/JFWj2h4AomGC6x0PZ63dVD4ROshTvhnhiBmVlT6KXX4vdAXc2jjQ/ZNDGiiLR
tfaziQLYzBgFAnapocqxNPNNPERj3o+wa0xo/xIit/1AO/uPIWTnoFUZgC68EsG0IWWRQGIcUytC
iPl5V41jgAGF4ukR5eizxHA0WwmbSZHWNROUhC8NcM5Cm8FGwiByZcmL/9Dh2K8KPwYZzZZuYHZI
AjRX7Cvf0Q7jEOJ3eL9f40ZHukofN3T2ujg1ONm40qkMceRFkYOBpmq3ZP5kaKsaT3O6aDkCqj/+
VdipD83SQYIAF2NQl8fhEnGXLaAqb5nr/s8FPAPBrkt/DTNkSY8yaA0/6n5NZBTsH5qWXZzf8OKR
JY2bwwTwS6pQaVNw+jdsn9EIVN8uQw58x9H7vvsd24DvM8lG5gQ6MaNYQ0PiTVeDF0Pd5BSxfF7L
iUgu4Btz58lFW0u2IScHNVJMEfw2UQV5bfhpQmNncafMCxGG2jyxqbTLj47Zz8j/1dfgRV7nZBK/
Xwv5mCBDddZojZCcsQtZdI9BbjG65gymmsrKAojvHWMtQWDHd6TwlToUX4nny8aFN0PkFssqX5N2
W0OIha6nTCsL0rzHoT0ZScsvdVKIDXT9FazLO7xBr/uXH6xPznTnaLOGvDcypPDsk1NoA1na+MjF
gOwfiCNqwREszn+V/rRIWs9oqeIJpnr1jYGZcFXXjj0JzWnsVo2ZAbiz3voukOQvXdCTnVjHlHEI
LadX0MwnHcZqt1zvO8JYPnPHjT0g6L+rACxAfyVIfBBHMrUDG2zYM2OD57xoGsSVCPeTOiVLMbh/
U1ikqTh/fIuZbnWI2YJWDzibz5+GMRv9/pUlbSou5APKnr3a1rhZFbsGTmkqsu0LoTEsbdwzgCQ0
BbXt+rvLnkvJ+ENP96/omyXz1K62LuEKQkgZWGHkWZmrXNONDtZoNoHeJMTS3ocwn+WPFkFxFLe6
uTnQqJt9l/e9Xq0FL+OtBf57k/mGSXMNe70LoakuvblRlR5KRjAUd7lMpc50MhgUVRGiVPeFt+N8
KvbIYAZs+xL4oK4IiIoyPuBSnkiJUD5Ujmd+3ZCe8CnZpSGt+OYSukeiJZ5YXogmk5ILLqM6/CyD
lOyfFPrj6inbPEub4bGY2zsySo5QMFGp7n5xf1cw7hCkon4PKotAtWDdjJ5V9kAYsdsW0EB9AMh0
2xvJRX0UOiEsOI6Wc5aTf2JvGr9vxkWaEGSuKqlXmMGRY8icm9KgaPQn0oQyGPbprOv/SDLfrMpK
YEWtilzbjjn/SWYy/XPN5Q+1EdMs3Xn0aZHWnTA+k4iu4UUZ45mZpw05ggSj3AI1xlQ9daUq2hXz
hFVYie6CXvF0kR8S+vy1kU4L1uwuIqetwqOmB+12k9aeUM1mmL6+2A12qE9Fh9R+haw//yuQqm6s
fXwiPg0nVPH9JmGMq2+CAyaKRZyPkHS2zS/9TnUBApcVPREzzJ1aABrVfsPnjaYaNWbDFcLRnJQi
N0GuYHWufky8bhtphELkSYIehKbj4EI45e2Z8F9BwU+R4QIiEXF06IAvYU0REh2io+6dys/ocKVC
nijiIokD7MfbePRJSCpexao28q32CCO5XqnE11OL7FLR3F/p8Uq7iejvrHK1ejbeVYwuLYTXqjca
avqXbJQ7Q4gYhytCgm7dAD0V2y1PMV7lbQVQ6/XeA8avOp0zQNAYkOAUJ5XgVQK+CD44yTRLpQ3v
vKYazkYuZ0lVKXnUHmEq+SFEpgSBb2/G7pjmBzcw+QYG/UJPio57VVWkQHEMiRunj5tW9pDDJuz7
R99LyBL42eCwdb6lRABaxh80zT/ECHs0V5bQcZPQ3y8ZqS2cWVV8eMfEMyLcLh+BQkQnG4mt3ssH
lafTLH/oYJOS+9zI628yMVZFogoiYQEETOdURFXBzxjDZseNEuKEX6ZxXjctjiF7Z2kc9cQatBAo
aOTeRLzizGx3xtwItAgbHDMQdy5WT9w2lyedznhkSsZUkkZ+pLH3EuiIyqufMtQxLVsksJHNKVFf
zZyQwQZ3y16gz2J/B5228fK1Lp0p5pp8Qp2aUo0SAakuLHdM5lCJUU2VLQ0sU8AEOD27cH2qlE1U
obOmW3o2EqA7MA8ro9LsupvWKL/PyJYUkutCEKQVDmCGr2Bq7gkSksVfWWAhJbYAfEal76kWO3hi
tLw6HPI6Q8wjMCkEPBDtwRyJubnDmQcK3bnUN+B3RqJU6RKN6yJhnqp0Z3YfzqYdkmCpIpNxAE26
bh2N7gzGiWsMFg8RZ8ILj9cldM6UI9TUl6pm9Owo8Qipqgynmr+OYNks6RTm/Sv+5N8Ba0TkCT+m
Xua/UXhfynxvPPklUXWCJbJW31Sjdrr638CDPRX8K45zipGPE6zq3J0GLCa7EFzLrCc2yA+C2qqv
7Jbl4cqewppxKhHGu2nMggsIssMVPErOls7l085BKn5oBn+yNFtnPiWoxT1egpseDDrT4JcrZr95
oaNFzoZDeYnqYOcdKekfBhCESUvWpg3SD+U3QRiarLjnti+Bu+2v0w3p7kvZJrOPLI992bAH+OaP
muQyrMBfU8uDucHsxpx4O/KZ/9DwM1D2ESkLcxjnSBUlXc1vj6JGyLcrSeDvGoxKWmW8VbVfZWG9
Tb/GNfa8YAdbiKG8Vox/IW7W46ruQ8GrHl0RDQGKknq5eRiFBn8WaNJwm57tWYKsSolf9C0L/bRN
jETsjNV0ucH7zFpXr8y5uxqdqnJlxRcSKhfiM+bSKZsLUQZFwFGwQQSKiI2fCGpVDFXzEmctt7nc
t3IM+LPaFpyXGX/SMAy1ohohfBcCB0GONrx2HfMWW+U0Cg43DPzVLJvXNwjimfxKqgBCvDURViTX
XbwZhQMTaTpSadr/ICKmu/8MVscpGb0ZTTHqG03iXNgXLpjrsoVkIKwCaytMWXXKZd1FBfJbop8t
WfUwY2XZb4wPEY1SS50HNx9PsaOsSlF4EPgEIWops7O7I/JUOY8G8Dl7cd1q6e7PF3FEyjODUlbG
cts3yunQetMRvLH62m/b3Ky0Ln98WjIcjf1E6Kqul++iGqaDx+kiXGmZ1A1i9zYSrbioHgWMtUBy
c2TVxsO47YzwAJ1JxJpS1jK2ju/LKppWpux3NwG5IoJfaQ7TFgfx+SzUFWavrdrUf1eoTHuazbjp
sZuWIuSVS18A8idIv0S8jolNpkt8h2gf5NeCTPf63Ou0WMubfij83+GCJ8Y7V4i5dRMlo6SDBkU0
0IbRHTXPqZGLttJDQdb+tfOGnjCrnzlB2k1yIO7EsDcZgPlnX2AIKEBGsHQU6em2C65mhQrJSHtX
XcJ9jmNcQR8KztYlU4QewbUYli5f5ZjfRxv8a1XymPrUtQBIjCdzcCMXfdOPxj175EoAW0P509O4
b3NBO/XZYlT3AJyKdtUZxwS9WrWlayYsF9MH9JYVyj/Wvp5zDhGzyG8ha6OzlamuEzDDx5fzqgOh
R75BTjfvPaCGbr3ipsTZjbbhhqY3RJDZxJzP4P2PZ9vKY/YC+lm5fNXOUx+lL0L+5isKBHC9pZ+y
XoJV92Gg/9YCIJ9+22ZZhZKmzUXMwm1C5WKP/HRXRi3xfG/JLzFh99pzVAuhBS6kR5fjrN95ccHX
PtpfaX3+wZx7z+mNPok7N7BmIN0stdVq6srTpKp0WdQZNr5B642ShKvDb4xfkR6K43fEdN4iza7j
TzPxw94ng7CL6tQYFY+bt8brvQf93RRby0rTW9552F+SPPx3fVq7gdNTS9Ul7G9dI+4xV7bFnLmz
9LrnoJEpHCTAE4MSe2aW1OKQi05KPjCgtCktDEGvKR0z5+xJfep/gl6iUhkZlBhwFfbXDkkUqp7U
K3DPaRokMFiMW3qcmtR7+reVO0MBiRl3sCxwqG3SlBA77lzzs6zN9oyuyAj1/FUz1XO1+2bSpkBd
Q1OriYGKDI+AJlIxlr4/JDERW+nMsUpmQzt8pk08x7k3dkh0gizdRUNGwZB5+LiVUXlwkRuPcvxE
qKDuC/j0lb+apku0F/s9j+nWWGyNQ5kFHNe/yx3n9jMm8cXPdrM4TynU2klgjOZ3TMO8tJry3jb2
HoHebRSOHBGnUlEhr4m1bVaGL+8EZE1JsvSiY9y+Pnfp5qgDGaZUU09vcNmJJ5fgnMZFjGlgFN2s
IbgaSkAsEsS5jIUfqQ8Bui/Z9ZYEZzinEvukIedJ4d7ixDGT8PUYdvNFFGH+bDLr6fBut9fI0nFb
IdzS6dcqryq6yWd+aFePFQqFuYowc2BAC0Y/V49vn8oC02uud2fm7LCdqlwXA2plyaAT3ftKPBX3
xDbPZcABq3DXB5mU2pY+oWFWuOLRoi5tVaJRrXYVag2T8OX63p0qGH069D5DM91UQktBTtumCPYD
7J8+qTox3xmy9bsTtvHrjkMC/ovKtvWNAzxHO8XvWGsRCOYLjCWSmg3FbZqaZd92HJb7UOFnQOjX
cJMOaC+hTVWmCGb9Re+6LKYX8xT6kcRPeaRMx4ayWrt79fjR9cmmRg8Htp169oTyt3sVehQAZMlL
Wjkes7qLXgSIhbvE60VkuxG5H5CZvj9FWQA7RfVWaF+p5WaxfVsSTUKM5aZreJXDI5CkLOx8T9Di
uxp3x1c6uhYb2pDbkpEeU5beDqx6Ucu+WcG3sGziyriAYS0HQby6j8JtvouYULNzMW6g1x4Y0Yd4
ri6otJq86jOzxQkq4H8if8dLhFxvX1KmVuScOiK1UKPjddfpgC2VaxnVeOuil6nF6Wq3xtxr35jC
XheKaeFtgZf1m4Ry4MKNBFbfieT4LJHYc4cl6gv4hPVPxKWILgE9wo2ATz71ZWGhnjgdJV2Ltz/h
1+a/vkv+Z23ooZbTWyzWjd2OJO18taWhuSQwTpKM+QQXMQwlDM3P/9eaPkjLgN2W67rUczNznil1
dyEp5DKvV1xYvzS1kJK98tbiMmaOVXznn8Tqd0SHtFQ+9Lk400OpquJiW8bg0i9rTH9dbARGSFuY
cd0PU8TmlecOIHFsURgs6PBQoDnCldAy5fjMfvJJYCi3Juo4diIoXV139mx6ugcpGggV/uFWlqxI
ZSjT1UFBnTHw/TyDsozSedVN01AEi6+KDc6/WpFPSX672Y3HtKGipc+kGzFdzUxXuSOuxxb7eede
c6MXqqDexWl9VpkioBC8B9u+blgSEFMEDR2zEUsVTTPUGNTGoqXxbdxGZ2PRGWUnD1Hs3tOYYkfQ
3IIws5Tq4w2BiFbjLzTRYa5QSBiRyYO3nAdugmb84nJkRlkZkHZL/4+Z1EMxBnUdFq+frO5GdXz9
6qA8wX7EqnDbcGxF/BzyT7qkfiD5W2gy6Gg3/poLD3rbSie3KSnd3ulBuoaHBjAuMCZ2TGL+qK7c
sl7PY18Zlagng9PdBcWJodTrEl4P6XH/NBDdYEspsRtybYq8NhhOOjZ5bo4PwTxS42wSCHL7F+Pw
n+RIdFKzxfKx/t8d8uee9chORxcQfkJBKiXYyB7kg4gnKulbsTQE9IQ1fldZWJBpO0QfoGql8ZAc
QciL4b8Df6zTQN8Dlx/AJnhoKr9cgDCKWjc0nViLO7Dvi0b2RX7IDNVdi0r1jLZjOpsk0B2PsyWN
5VZhnl0rJPjh6geZBdL2LUcBhk7lGT2YAZg8OzYMpknnI8LmWivDsOu6uLwUQ8hwGmzGj7MBE+s0
jeJ02coKAMvkzrpAKE9TBMvA/auk2qPn/jpFuyuzmyUZZ5QHfw6G6t4CwC1ZoezHK1MrBdPUypf3
6g33SevO6D1rGQMdRNkoyLlo/YJMBf8phTtNsa9PIOSkgxziABoLfLkp6v5egDakJKzwxe3RYVqR
0pt601Usx8H506wy5PfFUnlhArV/qdMV/B7CKl7wOZ3LQj+Go2VXBbdUVCpC2dY+bGxXxUdCOM57
KFjTHllCpjGN4XsQxK2ClJVtY2oylhRK08cpqsgPzf8B2uqWKkXk15cWwCBevU1+K7bzy+yekIjD
Y7Jp92Jik7SOeaK4FWsqjBpPHm04JEfxT8nTxAHOy08fvvCD+kknpoAemMfL0e/1LBqn9uXeircW
5cDb9Wcv6CVEVTIp/tNnVGNse+RWsRoKBqMUrteFc+vTckHfXpetPhR5ebpmRRYSrul5pQSaWHgK
P4Dh+YM9oBFA1YNt/pRWGKn5upYlu59gn8xmhq7+q+DHnlm6DAlzZNuBkhSNLJOfhfhTMoK6qC8d
5LakzqXYuductjJ9T2bcvw4rZ1qm7r3AvoKLF1PkiQeETBJptt6QwMt/fJ55eeVlx+jxdq2G5tZ2
/vtQwnsQkgmwQX9rC2KvgDHxctVYYZZBhjSDIcnEgYQcSgn1+Ua6avxCA/SoTDEVgAOQlZiD2eIJ
VAmtH/1850bT9OY3y3TpbB8Hfo1t71jY8vKySJ/x/P6yBt2Tv15J8o8TBWrh1dEPCi+lnYWo4agx
SqFt6Jmxy4HIMmaTdjnAEDMK4J+MTcIjsKAVDtDCtkE1MBJCILBl5fQex2XhtIutpa+OQca8Kg60
yTHnE4gQ3wnfcOZ43n4Pb3rNIOu5xgDz59rt0cQgBfIkCm6W7wDgl4oMRit8KP9g3lXLV2Kz4lYo
f27xqX6n7WnAS3KeZPY5h6Ju3YRbQJX1yJN0A0ruCTZoPpPSTeIFHCYv3FvacODj3xDrJT+Jgo1i
myuyk2MjDuqE+wdXY6OM3W94wJKZzUjeIdkZkDpoNGCEzXzPkOagAz3Rld3srE6JX6W6Bh8so+uk
tmfZQvQZbKx9g6m6YxxDDONXJ2Ea8dJCL4S1r5d22u8XBxEJVNZQwblXAJArEF+5bThRccWYoiei
bZ9nCpSbKuFkhiElKjWYLOOyKJl7KT7K1Trv/CWe5VGG4SCnK5l6jFyG45mLVsy02Zr7EFi4D6RQ
8xnxRdWO9yR1XMWFOWfxO+7u9TH08/n3IzTwXG1AFHEDK9pE93nrh3mos+7PmHKTA7z3msqxrQlI
RxmDbPOPcnwJ9o+peFlW/7ozmA+ccWvfVW7Or/+ygmhftoSWLGaR96FdsL2Plj92Dsp5OO4hIBTd
LhQTYaEBEwmv9u2Z1zA7/F8pfdfAhDeftYSi8LlHgDQvNDGBpvnSaIM2E/N2/H3fWqb1kO6tUBpd
2UjvKx1svcjuAkUqqtYX+Far4bbHT60tyJ1henRD8E9lEbXtdtWKhF8ZTVMMm/FIbiazlvX6EZd2
rGIWl6RwsVriKMa/HxLo4T5RFWH5701ZD0N8jCM/kLlJdSpRaYbUv0QoDUESsgpABMdYmv8RisUb
sFQRvMqmCqulfzyJYY6I1JTVrzFZpQjQVbn707Dm8r3N9lbKyU3U+Tkwm4/JP2ERpF+JHSnuD5TN
3Bd0Y1z2fY9otZRDsaxRhNNSFKql+TPrmfDNJBi0Z8+PnS8TCefjAchGBDPxDgVHKcLqteTaNgIW
2NLPRoTbAf597PACklUrCFXwJzRS7VcH8wIox5J2NmUv/5J51QjO4L5v6MiVXPMobuZa2SdFqvJX
tgtwcnNNCDEqETN+1qkPvXL1OSEfgVU7yt85Xb3cH3QH2xp57Kj8EeUv8aTRHA4UqjmNUdy5Q0ei
vkvHMx6f3W6CrNMcD4/IrfV5VmHbX9X6OjXe4WEIHfMbDtDKUe9Tclz6v9xSqxJJ6Laz7AKouLbh
CZkhWPxUioKSVQ7wQwiLbMRwSu1489hxXzH/8KoIVPgPmNgXi5zxxzF5aRtrGKlKnpyShFNe5yFO
J48EpWvCJ3sLu1BAYbQ7kM8HNjmCXzn8jNwOSaXY0NWIWfPwCat08hE6rVsAxTvLnE+4n4uzudeW
2Dr8fxATUqOZXrNQPrFyYQjxX3lyaZalRV1wOZbqGUNIVYH61Mvql5JbNfbN6xkF6FRNNWJmL7aL
RTR91qPsTkgEa99Xw7mhkyvHTWFUgRl/VjZI7Yo4XxxVCBhpG9/ot0FySSOO7XXO4R/53v/IHQil
XL/vYRKfNIREPFnmQc6io2fm7+WsoMbBTbdQTxkIaN8gaG/in2fU2OpIIVQ2thumrP+2R1OTOar6
a4z9lVydmiS6xEP8yw7qMj6nt0z4q8KF4TJs22TxyAPu9F9NAmQGlpOcN6pmttywm7dRwmiudqEx
eyc2d3lyWIbVSMGCxtreeCTDx7hLnZdyLCPPA1dnTD8SXDXP2WTX6m6ipVlitrMxkHIEDmgUpMLs
SFQ5KYQVQDWhWFTCeMwes6eEJ/reROhwNSoVpmzho++PvrUMqLB2KBC7/RG3YHvVV9nir8CIum0B
xD3xnBgWvZM6ygnsuCb7MI2Vq/QEEL7leCn9e/grWJKqwuIsl23xH+f6nsY44puEXTyj6gBRyf6I
4UPEJkrWoPjG9ZN/LdTodZ3WPVoLXW7jUFwS1VLSz8nsA7im0o1LNimlRwQe0FdUTaGWEy8slO3g
HUJZ+tTuhEPxRjrHD1X1M+oa+50OndIVtzMjROeoLrBlQJeyB3Ojk2k+bnq+PPOSO8rLUGIjEMa0
QzxTAZP0d2O7MF7DBYZ9ETAUEFHK1QyvSobAuGypv8CPDpelhUW/Sbloq9YNUm2r0d4S785TqGkS
nJWCpHvgvdrZOwbJGhFU52CcBYSN2gUJHTrDN3KFSId2AiFDXmfQXryo88O3VAIGEbvHx2zzpc0U
6yUiESn6yEfLPfGdjeJcqir4KXHPpzOWzVpZ8ypXTd3N7ZUYQ986z8dJ2e/YyxNhHmbGkGmD1qyp
6Lza41z6f3fj/2Xpy3HBfDBZJr8WhjSc1AVpBNPzdOpwGv7SUhm8+ub8idHVRRHbaCUaXkuGnHYO
dosG/+50f8Z/Pcq56FzeISrbWfDjcYbpmZBRCBVC+mRW257nKgXrsmmwJyRYDko0LGQpF7yiyQzL
HIc7o5k7ZrgB4d2KtHumIuySTqOMBAa7j2FfKXIxoRUE3K7fMIoLhs5uTEuvVhLYfa557c0cpJjr
WETYK/G23ymNSyzAtQC0Nb8C4w4ojyvgeC99skxIRfW8fsUKAY6fI1Hw3715IgL5PvmBxG9kYeT0
DDfXQ95kGGR+yYtzJZApScZfTkjS+4wR4ggt3Sq76eOrDsVxJpvqRYFh5ocwfb23Pr3FeUkwuP5m
hk6oF4RlkkvHG0Rbposjefh9tqsnTQvmh9GL3GDwKX1hv5C49Ln1gxXD0W/9XpvweuYdvHRDkIh4
dv6MGdF3tYCemZJcpncuiTCLYUECOJ50dCg5Jh75yIdAsD5yWbDbzLpDG9uEGUFq4/VUsvuS3mi5
7m3MKMjR247RC7soxHRDTaPA2Xcb61marz6RlDTVlpsth9Rw5Yk6O5hGp405V9mJM1LPfbkj0+SJ
/1Nj+U2HC2xK3T4gBCZh/DMHMNymrpWWsAo0PIGQBFPka6RArEGsvLXnlDrB1hMlvnhHK9NOfhA1
m/kmnbbx/gkJRzkYPa1dOZRV16lXuxjaRR+V634WI1k/rDSqokCI2U/vh5gZZ3hudB2XstbJp6BZ
I8EUqpqrYZcYxDnH4SyCE+Mh3QjeIi7O4JxH4v4Xsv8yd3z/84ucZjt0G61wcYEcSl/NsWLTN7Qd
/QejJO/iACxio1ANFncl3xi8CQz0sBCa6AUmssrLACVdcSUd8xwxLbiaAWt4SoE5h6voKqJ2nAvv
ojq9F5/zX+3wOKBYrzk1QGe5thl0tec3h/b2nPRm0QR+25iE6jDAZxGCyCh6f8T/y0nJ7LuTDb+2
Dt+UNIVpfMxB1LjXGF0N6IL+Dn3IdiU/o7fMEIrfGM0edcR8rPL8g/ZEqLKPuocSD29q3dnilkLP
f2VXPqtnVAH+439HjyZMHFaz8gz/cWOgUYowMu7Vtxgn9FzEqN/bmoViAzXblTPoe5XiU4O5uEn0
gUDw8VbtvFcrgYepU6ZOgdYG4uv5lSlXqLFExyH2+DCZqfEeOmjPzlMS6W3qW6UasnTGGuSXHDrm
vlv16wuXuDKeStB79yTPe/zEzeNYvzCwGYPp7joSl8vUV2E2/jF0HnsP5GXEXaHAWLqP87SR0A3S
Dolwf9QFrUFyPYN9teYtlafonlxcY92YR77ghrdFAYPYhjCEdU3z2pPpfPvlsR3L4d64yqSWHMuU
eqvRVYoQoQjHYTtb/KPaDJb6cHiOGmht1UPA92J42Li4SbPOv/ubIjOPgXgAt4d/wCnOixOL/OjT
9Qf1zPi1pLFt+MhJykfuGhBJQYjTlbVfcA5TTsB7dMQqtkwhfRtdshXt/uTG3AF6P4RqClHUckHG
1gwObPKlZtVhakPomikFNiUJfi2PlA6CJzHotLZheIc+MNZ9fklSpOhJPQDNxnNPxw7Ntw85lXez
i58nqFfkQwOrN0YvVXtKG6gV8Qwo7fT9G5g8Oe2hCXaMevcBRrGp9330hglYzg0MtYmLYjV3kYj0
TFG6ppFk/YMx0342hvYrRI6K6kjp0fAeI3+l9qnMW7ao1N1q4UEEfcuf8xb4dWek6L4+y9KoX4u1
h5tyX+U+hJ79023XWH8zIrdmtUdqjHj3N0HBBFKKYt4t7yzGs+9d3JhY6Z540wGkEl/hAGhdP4l7
5swe2bSbXEMMVXKq9D6kyZkyoEOVED92ELmLGpoZsDD2GjJ+pgA3XSWSlZl+wNegDTxq28hSZXqP
bG7p1PTX7YOuaIAoGDl1lNUy5w/xWGeUEK4gX3B1JtdQ2a/LA2DmragZAAYEKZv6Rvjc9SUCQkU9
Ughorhw/4PrH0LgwiQIyVR2P5aUTdV+tk6oxprq3IOD8lHZR8KWW+Pbgeoi7khTqmoyeoJiPDgQv
QnCH3uNbuNrrI9trFlMk914spvTbw4b5i2TYbmu5ROdjGPO+ZB9AkfWKCDq/VJjo/roLAFg2/ZVL
GFgn0Bfe/sUOW9ZNk8Jzt0OBXlDwEoY2uVaSaRcMr5HEoP5AHJnTZKXeabNKz152rsriygOyIVw5
Nwcjd/s1AaYjY/VKITz/M3+dpq4aSVQiUajzF9Mn6LOc41mZ1VHaT3aBzCgI/UshSpCfGMVTjpUn
wc6tS9S9atbkfrarqN/Zqn8XzqxVrfRJ9vJUqAuES2eZjc4Ep881uQ9t6jdXO7FxUgu93Tcop6RO
qA/y08F9zMcKJbtjIbeguq+FgWLw7GIoX3PedgGsVy509ctYctSCTbDnEAd/vVtq8dhgogQ5HXDK
EID0oK809bpg6TCFXigHy5ELdIEi/x37u02oSigvqwUHXbmL+6mjwr5yNgkUC8vkHnyDs7jhdRyO
lMnhBpC2y96iudnxamlJJE4f778zsLNx3KxRIgxwGYwoFejEPzjG5KkNCyniHtIWyVi0U8l7VggN
e47WG0o1NPmpDXHE+O9C6qmyOh7ql8TmXXsPeNhvWJaM4fjHySKYOzeRARWlZUqj0FaWaR7WcDfZ
fHNN6SKnvwZKTOxD1rTXgy2K/qBATGFRl+EfDRAHUDY0O2kZadSDICu3jbwtexrgSaYmgEFS1r97
H1wjqClBCIn9VtRh2r+hxOAgwGVixyT1+eYl9i8law9LKlTqSnFN23Q16VPbwaIMIFQb7oktm693
c9Ys8b2JhXJ+A9yFBXKh7q33C2ybcLgLeldioN60RK83ZjgvveIj7zPX7psI35X53wV6EyvVWfow
vMOv6l/rNIlRvdbH3k9PiMwMS2bGCgnnz8chTLRFJIrGjEvZpB835zfGsLKrdE8KObej88a7Hzv+
MvpLFG87Z8SvS5579oH0C5a84Simdd3bTRwWofOQRUmKmQdEUcGEs8yJCSi0rEDs3u3FsraL7bMp
OB90Vef7HJKIJsr7u1F/4WxnQG47nyWNoAwxNVE5JZgQqLDNso0szrKsBdFZ/vapzcnM3VbUp1ba
7SXYAFR33hvqhe6aGNYOjrYnOp5poe0R4+FQztl64XU807h7oqyZSvVUJWyJaVF9hkOktK9TOnsj
A7TT3dWEijUI1DcJ6X1BnCzkihmLh0T3jBbC1pqbUfzHv3S86a01kmEDgm7Ohk3dGel8Kngi6tOC
qFU/O5w11YZFXYP+aQT8Y7nlU+Rw4QP4Vcns1wAk04kKX3wD6xmCk1L9/sMTks8oKai5qnT73q3D
YBsgC+voSbDg2GNLUAHRbyea4CYJ8cyFcHCtrJ4lrzBgdO1kS3MtuidTtIiENkaKYPJgWsCTlTUr
FCnlA9ueOOYSUAAJcxvJCjBZin/iX0ooDUXCuUdT1b/zqa/03cy7JaA3vW8mycUN2j7z57suV6J0
OgOhQQyWhPfOsksWfAjWmJrCSR1exs9mnJoHt1/CkZUwwJcfUmDvDvP5gBKqEa5N8+gG6Sm/cBAq
dHQpOk5dJpTjrQvxF51eOwRAqbzy85Kjzgh+fnfCfCn+gVwu4bSgZA2CuS6kAHOxuuKoEWmlso1Q
/8s6XSHkj7/vvLZflFXpVVADZ0i2ao9BQ5S0NuQzeETJRs8Pxqp70jGPU30SvwRBFfUM9jMh9vHa
KynNlTHMThO5ygtF7XoKqPkSIJz4Kzbk6D8IC7WyOPg/OsELs0Vja0eHtlTjZ4CT7G0Kx7yOp2Hh
3SMfszlMKcWRd2CwCcEiJIrvBxqXs2xGqRBGp1/L5JP/3yk6/Ktp+xdcZu04Ri7pfoyQVL3Eg7yH
arhTT36owYWZ7krw0/Fl3IcWbXXsWwE4pS8EUKrnn71qrARdecV67H9lHtWXmw/WCZkMN2Uw20DV
BepaPoXeWDAXCHnNqRp5al+AKCHtSjcDdQ9zdFq3IfQnHgNuYakpSmyMw8XwjlLAb/Av1rQ8WCr5
/oKgUUxORVUCTYQpI7nGp2ztEcr2C1t5CkHKe8XZDCI01spLqmva6FQPI6qXjo1AWGyJuBNBwBGc
irR68LvFK+MY9wbZGftiC7s07g96W5LuxUHAygurc070YL3A2l/DDw9d4hkq45rZjxKBz+9MbrRY
qlkWgmQ+VupqsEYygHXUIb6Jm3ypMDz7pfhQpN3fNPcfBtleVkOdaLE0qInquX8blWM9xuI8jdwI
EuwL2Y35rOAN2vYMurxuxcaGJHd4LGqDXfAXkPkVem+H8BfUnQwP8FW3bBr1sJ3RPwJdXMh20kgQ
t9BDI2FP2mT76Dxbs7g2AhmZdgLAwjPh8mnwkbTfrrdKpwidBOKgw4TIdv1bxCHUvp7Oyb4TWjAt
qQBCxb4nrIkXxcjUjaIv4i3WVv7E4ZJem5gUUQP0u0A/8BRYU9u0qh+hq1akVlYEH7O8SXg8bb3L
UwhFQ3aWepRPRk49alD1UNgrjfltAufLQ2moKrqOURfoghyxmBuxJ5e4FlTqJN5e2ue9SNECRHbn
j8qJCT7y2NJcn7Es0nC5S1ry4fFDPtI79fbWBBXLMtFwzuJ3IZ/0nuVWq1Y65YhA+iMEX+6SBUnV
RhauDzSMP2A9vxShemqrjktUnrU5497+Twubz6f0JWhgh1M+gINLyMvxaToNUQcnNocWt1a8TJ87
JDCBN3I5Gl3pp15v9mkZ6EHxilupgMMrGqmCa/xt1Y5x/+EDxie0RWziuz8lIeRmTCrH61hPkcxA
EmoEMj7dP7ee4AdkEMi5fRsrGWdGpIz/T+6l2zKx3NZcT+fbtCaxVMGP7Xb+PoKsAFttXL9toYQH
hzEp9jHGcklelriX2bI4iEgRvpZxm6wjIYL8aUmClSmBMG9gRmYDgn6nAAHEC8Wrxyqroc9kAClk
MRNpEpsLDrtCQ4BHMp0EEME+EQ1W/nyOMwO/cw1N0Kjzw99wWY+AdAeiX9yQAS2wMZUi5bDG5m8I
sR3omgiVmWNC0r2/ddkaz71duUWNvTZhmnWorH5q53lhhcBBkSM03enOCwrSApiYVMYAWYUoJell
AlOkfmiHcxfF4qMFUJEdgOe5muLP0Bz1PQXKyz9iQLEKL1pggad6Enln9APgodc2hba6KYmEWuIi
XFSmxN9voW80SxQQrGNtQg7lMAJ20LPV0CSrHdoaUIjdsF+A9pANfQpc7ep/8d2ZV8pdISLbkAdp
NQFYx+fPH5hc95uToNBFQmcA4/GQna46qPCdpE6zsWbDZAjWkTehwmyM+cM1rzsK+gHF7sRhe6JM
Utu6yOYX4svYdxweYFZRDq0ELaOrH9HbY1Po92faP4pbIbTArEyD1z5YM2WUEkGxpbiAxKyMtZTd
UjEUpQopz7evPnv5MCehkVg8U/lmVwvJzAfkym2UV45huUQkWUc7sG6Xippy/jwwtCJVe66UtUZm
ZRMDAi3fE9ffuFUJUfghBYdgHDkkqLhvTKrn3exjEyejrFKJKHpdiiRcjdZuyUjUT0xlYqyvd8bQ
MVuJ6GiTt8fn5fUfF2by86FX2Rje+rGzrEiLiTagVNP/x0WOrIhPq9s7uxhUsRywCcA3+d5v7vwX
aakHPQNvOSBiVSwBPZRJmP1ZS5lk1Hf0daNiuDvyqOl+VP3FpVDA4nX4D13oDH/cV4jrIOyVTPFF
n1qUn9v4pHIVx2Uq0P1E18Mr5h/iHah0XRxOb6hUZU5jDVEeDTOVQcyuxMZFf91SQ6XC/pI42LV8
t0V+bWOXf4S582kdW2DN2plawF0kJWdsiOh32s0Vgn3SD8V4Lpdy33BoHq2whdUlJ0BBo65EYwMO
8DFiqB9lDiQ5SR92Qgjy6IyaUVoGxqIg36J9NZpJTPh0Nr2T0oPJ8LqHOwbMzbKny6tZXSbweEV8
Pa8NecQSCBfK5DxHA6hHWWW/VYbDw9iI7/1/nZ0i0dX07fJ3mLNpG5joIz4QV+2rI/O4hTzpUX1d
S5GjML0ycNe+HinSIck3wm40dDHvY5250fEDAmv5NPw90SSGhldcpWbu6H+DizWyEDwJoKRViVi5
3ecix1CafynTe/h0mMRITasacZKoL5J1rkMXIJEajOO5rqUOEos5lBJBqE2l4NAzp33Qw8Fi007Y
F8XJEjNrZ/DcWdEhe3OlU+W5uzzLhzyEv9EusmCvFK46qNhBASQldQf9hr3ETqw1LIjsrRp+CEsI
MrRnETBKKFUIgZkbYelRU1MsmID/uWV9caPQxcx3UhGIVycw2KXDcX6bPUMDx+lRCLdW+ASiXeme
zJzK7aJWPPX1tQiZhD4PkdvKrR+bKKPpiojcREZVsGLbU76QziL7KHumfGsVR0+byI5pF0DlDccv
CA9qQ3kMG8xwfOX4WiSMSZCI52/iYlz11/b39k4R4Dmu3JIse2/hYZEhBWjON1osJOKOOk8DA5N/
lKKT/AAq5qJPDbBNFkC4ge9uuCREJD0I462o76785O0IyNAyOLvfxVndZKTfQys2Ps5NLyWipLKW
qZABGK9ZFqVmwv3DwrDfCEhnzltKdy5/uYy7WabbnbZl9nvhxG6cCpWQWUsWJMmq8cdMCMeFqbJV
2KC/hav5IOxFSbBVd+NyDmxnTgHLGVSzQeXnDmaiwNPV0vZEc9LCM4NojDwjUzKpGm/bV9Azqme1
kmN2L8eX+JxOvnQmI8daK+z2Sc5ve5z5T0E3TZxcnu+6V6BzfOAOERVJ9MhbDQp44oelwjBrE0nS
gr3o1BIF3STohtwdbnYwz2T5N+BW3jJfKaQrgJPXLqpEiI+wvWqEqo87CyrLZWsXP0Yf5/D7r0rK
tj5KXAnO9GB2JgY7M+sG9cSFE6q6NGvAxGZOTAqtJUoBHw7uYXu4799cichlkx1x0kfZqdRKC5di
OaY9HBUfEPW7CwlD7dNLsqxtA5r24VFH8WQlCoXxbMtjFt1E2L0bS/ivxE3t/rSvyqYRc2fVk7FN
R0L/0R89bRGdLSsij/3NlREFQQwHOb/djSsPAwoKA8UMj4c7W+kCG/NxU4v/fsBVz/56sGXmk8ov
ZcWiZ5EX67VrbGOKhp3DQe8ML9Iy/LVAGLyDkDIy5hlGi/n221cdLPugW3rvfNNTAU5mnsfAEyz0
RInhD+AHBmZPFbpBHK3GK1OoEg8V5RrLJUZ6+cQ+jfEMAtyVwOsRY4lLCNNf79X3n5DtMR729sEV
EdXTNYsXY5OppMdLTN64Bzlaq0nRw7Ei1PP/K4w/Sg4wTH6yJ+PAC2e0WjAujTQc9qtQXpHUp18L
cTrD9cGiOgqDYUinKEDNgK5YKbr73/3IGNeXhCPEG74NrYqoObKKpJ2MrVtypLw4UXq6djRVXFCB
XDwdLJ8kKqjDcmt3uDGl7U7RXhOV8VI272i3LIlkiX71M5qcj2HTUoz0I+4Cmci349WXvZJLWfh5
KfnGSyPOoowRJyqP7JmWH9BFT1e3O3+wUzguFPNlVfTxAQu+mQKo0mg6w6CVwEqkAk9JZ0EvWABw
oEy6GVi4dtmDutHyYGaCETmOzw5lscf49Lv0VybP9iW3CPUUK1d9ar/8B+UACBDoYwhd3CD8R9JU
xueijcIpL9kERIU5JWB8KFPywt+3d40eZasFzdHF54AohxI/Wy1v8sfOYGf5KiqnFCB0ibNkhIk3
EUHgXMikKb6KCKdyGNdOH50bGUNIycX9j6CkEp5YVAyuUz80w7ifFQFaoHLy0wBN9xkx7EAmI3nD
VxWzeX4Myl/L2FgLuLJNbEdtoLHEmJETv5WKx4o2ogQNGGWw7GvgU0vXIyputgkpKJ2QRWMffTLc
U86QviObJJMvGcNN0l97syfBgVGOj7WWYnJ6PvI2+Sv1rtMhW59dg/N1aW01n9sHyx/RdX+V/bFI
Mc3ysykX+X68zqW5fMLZdauWkpWwryWm3EmGpXlm+VQ7tw4JQDLSMxeHifVlCckASQODZwRL8uGG
a6sp9xak7uQ+DXjxpFNExNTk5egA1NMIgiIC+5gcmO6h46skwddho86zsOe3cgrv4uGct/QKOGiy
1IdrCdHXDZShpR2I+vUbZbgg96pjnF8LgAg/bsMWr2KCm9NzLlJ+BuJCnN0jtMXnAmY6mii/1quU
3/XO2InMLcnEv94yd+BLRR8IdSc6Fwc6lMh06sKfukcoHi2yVBr+xX4ehMIqLg44ovB5abLL9VPW
bhvZHr0VOWoCfGd0k+0UaDSfIv4fF7CIy/j7V+2JtGzYpN0bQ0wwHwPq9QQoeqo3W1uVxv3UMqA7
70qVyNaB34kMAoiw546ucPnqo5qUJKYmAQJBCGhZTiAjxtozbZgY0zgOumpxAi+nYwIPAtxXkqw7
64xsecxyt6Ph3anHiGReNHtcut9zksSAXPAZnWBs+xIaHRHbvt7eiqGqPlPZrNcYsqgxltGo9K7U
2Y+e/Jn5jn4mwBY/ME2/iuZOIgvHbrkwwiz2BUoBJz/yDqoFmNRTTbSCpG3eiY/XIHifmdawz8li
HpE+f9jQodMh57T0urEdrC3NyM44eg/Ga52gaECb4rWfwQr90Y5eVnk0PrK00IzcLVL+U24goRfy
djDCpp0T4hf1Qa0QpxUsrMO0qO92q0ortqniXbE9h24Ty9/risbNVn49P/poe2KW2Sg0okf4/PHn
DrXf7bmY/jf6TUyX3jwMjtfKo9V6+w9VH0i8Ivk/41fqhPpFKneK3obl4C7dTujU521e+j7pyYGO
cuAs0RRqLXqY3Po0BDU432HaV7Ix9RdmgRVS+3KzSU3q+MkDcyENcIaWTEN7OCpn/BuPY/NIPKR5
KboYM5BG1oOqqy6JChIkZGTiGOQbQ2TfYNp5WWG69ZaR5rAEsL1ih3XPpnq7XmIk0Aki2+1xXCK0
fL9CvWNwQ2b8ULUf600nuZELRuqyWH0nBuSI/EIY7op4bYBR+oiaJTd1wuePJ+bwpbpp70s1QrIz
yd6WAFbGh2Q/CYbHM1A9zVoSVu8XfU+0puWbnalVIsC1n3L55MtBo9K2V/EQGeoDZZrApgyuIsQ4
Osiwyl+j9DmALgqMh/erX/B5M6V0CpZAMGC6Ht5h9dK2C6x3sBUAXPd92PKJx4KR67/CrG92kd0W
8lwqCBOgSvgo6OcDGmp6atCgMINElVXwORaVB6bKXwL6SIkdlLleYjBn6WZkMcbvWgApTDy6wxNI
B0eUbhs0nnnrSyl7/xDmbdo9zd6dbD+BcQQCcIFmrNFo6aXw28EKWzc5sU8ZGK4CLq4C2bdUdvTV
8+WNEUWTeiF6xO9BzFy1ewuasbJU/eeaLgkdMDFKiImGxGgEodwznambjJDmUC7gjLUYUHZ8Ue/q
AAhubto99P7kUah1txptBx4Q3vdatjM7M1L14adAQ/UcI3ZsSmF2pO7ib4z6v/o0Y6Xf54nUDjOj
oS7FyCEeK+RZgdXSKvvoIz87Mdy08v3pAO00MlheeR+XODW50T+h1jZblpkMw4cPlRY7rrzf9w3o
mPiquTOBcs211GVjswB/LApFHh/t3TWItE3USDcP9C93o/3wp7OjRnfmVjVYK145xdBsN8nqoTbO
cfdW7s9sc/bDnZy32INCD6bcsmBTt/W+FvtU4ERMOOeJFbiPtuH53K6ag9u4F15qI+ZPLU7H8OMP
Lhl1MGrUOs3bX3W/bjo9PDBtx8GnAaQFk5URkGFQj1nJTVfj7suOLQA9LHhLBcbJIFRPnTQpsa6a
immX6fldwhPXgwY4sRKsI8h+gJhn5WrOVcS8m4dBX9+JY59qdI4biYJQRXvhfHnGrPS4wiihm5cW
PVzDFjyqC2fTk9lUWDUmG7fX8F/UoHPnkbp6cbrogZi+cpWxa60s2bguwls0D/VoMCLjvXSrJyve
eXfAc/cnvZ6k/3bk8K08JOFbz28p/Vc+lXKLcaK8Ebn7u+4Qh9TYDxv1wxMCSDWmcDWVKL1grbzI
mxSnDWDZ6HERsMuwO0bkhbz4EzVf2f4xtv2UavsvM488n1eNLighS1n3Uey8G0iZYPQaV+hojUsq
5DQStvc5/cf8/QPrs6vv7O9LwvYBRjEATf3gazMActMGA77RSu+1wnFXxfN9UeKXSEXgRtwJkZus
5KXpqZ05utfxzfQyQy0ucMHFz9vkp3tAiSVPBmkQ4BAnEzvWxwr0mbwevDLJ9iM+4thkRGzjDRjD
zZjFRV2DhIEWM5dwsJvlomttAkIU03Q4ovQwAwOCr53dh6o9TvzUKMyfstQlK0uKe/a2PIUX8m7U
XvXkEeKLcEmZ5BY8vaJy/b0GhjensoCXX3sllOuQr7tTRY00zkZ/IOSW5OzmG+RANFCnUG4cnDNe
UtyP75VvLBwQURWmt03GlBkmzyzOujQd48n40LMuJX0pKQXuXHsNj8OTSo6sk9RXqw3L1wrKHy3N
9tvgkNO9lW1N3xo4J8ue+WupmecuZ2tZTnO8nf+ljOsHZuWFyPgJbqsZpWrm6aKkpnsrsKHN4WFW
1sY8/mbskZv2MrF6ssc/gl7OAKpTVLMnoENkRnZ4gw8WoblWEXlVfe9yLwYOJEcQJC5LwzJceMxF
OjVnpV/egEnTvmE749RtaVbA5H/4Y/zwquTmfJhJdJUR/h4DAmxhbTi3rqAQBZmH3C4wi5VB1S0r
47nGW8HlusEEakbdAlyH6hXx94nJtDpZ70yqYbTDNVR/BhL6txDP2jc/JWuGjv3e3N2BxjZa1HJO
R7UHB7khL1O3wKGMi3XskfsBGNkehp+WQxB5z/pma0cLX+/NpTo98Z+NM0cReVS+8QJ2RcYT6XXR
2TEceUG8CVtqrTKmgePYOsA+hDgKHCSbgdnXbg84YzSBvroNOWeE0OuBa4ja+DAtu9euCTWILnbh
4pE7+otgsyL5kINwNlzUw9+lfdNPTv2jSm1OzCwgu3Ac8jsKscGfNBjdBHAEElujMyjvcdGVkgib
sY/ke3aJV5VXCohZjxIHWH3djfGi/CgVF47fSOHGFzDI5y51lopW4Ox7jHc1AX40SYS2RYA0liEU
boisCMNGmi9jdSbw9JOXbQWz0jXUg2pes+53VL/2tRud4dquSm/rbyLnKNaQ+L8hJwJEQ9wimC/L
+LgsILEnILi0qSYaqILZXbKvZbQvJRTdxG0vwFcWfFTCIWY8Hcpm3+C+BBdSgsEBiAVq0qCyCrij
34rADCeAytikVQghxXc5b8Elyn3LC/Zlb6hF+NvT3M9XroIPD+JI25jlnL/8YUp0vN74FOd4oJku
gjQ6G6JPfEU2ZoXjVJEgBugG/aGYaoTrnUYKNZmty4u+hANGiraYQCiFwXJ5BSwjWytBQzyIlc+l
k5auXXDIAcWMU9EFDrfyjpcWTkA3khY8dPEYEwNZkVqYH7ZECUZz1xyv3tUje+DfP4KhDOK0oJMm
zajsrVamBJFFyApyimGETJxy8HnKa1VY/Y1lwUvCejk/8DBwF2tLUsu8ijLcqPOmc8yo66Y3Ebd8
dK/EnSYOVyAUKDdgyCvtjoOCHfLROfwzAnuQTN6Hr1ajAAG/ouHJMvRRVkl5lcHsWgP5sHdlrcJ7
fQ4EIiFk4Xa3e5R+/NdsGGqLAgpsm9qoBlx//KNELk7UUdaj1ecONE8w2jIzgTs77xv9JlCLD9Ks
HPwnAKM4sWil9wqp1wmWJETCi5sdSd1ps7Yl54gqmSDo1iYTicnjJi0S7Z3ro6FwKwZXzJTUXeWE
eg2bc9G87kz80XVXdogg/OXcxLu/UnmHYXipphZ6mTLBRNJ2gGjcsdc8wPzCw3Tpp3emeMKhMo8d
hhDfQX9hK2+6oPEk9H/rcynlQIl7e4URDJonK1U1tbs129Xbrf1I8Iz4A1nlzeimQl0UsK1LXrCD
3JhqDjZ8g39+4QgTtc+nZLjvoWKOnNFMeBsMnpzT3Uho5r2guW6sVTs3h0TOuFqN6/lw+jVgs+p5
anbAR/gkhaANfE7uhisvkGO7gGgHXhixHnbIiWSxC6Ulay2sHNu9jfod4Q8o/zlDi7Hi8bwdnp2V
PGFamh0cLZcX0m6URXNuT9xj/METRsFLil7K16s6WJjBcLRbNFhRfY1SrgY7PtmscqARrQHpfXus
QubeOmmvZ+YBjvLBlIcMig0HHopBb83qnP2CCmld0MxpgwafGLQ7ZvOZ+L9N53EP+Ve3Ek0tAoTp
QXWa+rIrVNj9A7NkMVHTOPtGPcC+eXngZgo3ilg6Dginej+eT0HG8S6DepWc3TK7QDNDxPgo3yhx
YsoDZm3henvQ0Ynd87cgJBloq3Z4Bh0OrkeaJS0+19Rf1W+eHCxfExWbIvDqU5wBuyBk3QWTpPc/
CGb+YqsjYfSQH55y8X4wltE04bc4pJIDH+HVTpPSugM2C02r32PnErKayg6LCd06z0DCsj4hWSuH
FQ2qLf3lqayKAllsQ0Hg7hlk2Hvn7Cpa2jm9DNBJHsNnAj9tufkVTAG4VOvxK0BBXr6nqRFNlRXw
xbulSUh4064hlbTXu03DbEpsOZB26HuEKC170bW4OMWD6TXIevfOnVwQfg4B1ewg1+CI2l95aKU8
cN2tGm6Pbd8r9crEzORCb/hnH5PO7350a1UguhrqIcJUQHfP2J2E6MGw/4B+tlcAkJi9aoqyziF3
S56alOBpXPJclppcvoIo8DjvsBWgBOLMDVs86Am5k6WYjkkRGejyVS8Baf+ih7vk/KSVB483vRSh
e0+b6tDhkAbe2uH6kE/aY67QVamh1P3JZsv/VjBfs8HtKfitPlwRs6mLDXqWsEsFt1c727iGnqyn
eSnxzxoPVi3SIw7D2wNwKfh6f7XtPLfQbNwdSQY7nhyB8mqVY8mo27Lv7cncHGbEz1SJvJ7qr4L2
ln/O1P4E1ibbjZLwUfXocWsIxEsWP7mCcTvxWDSIRLS0Xi7etbfyiN9M9eYnT7H9Vx9A60rJum4j
GJ3D5BGmKCY5txwQiU7hGRqJETiHUCzaQcfQAd/kfCFfr6yauhdx+GGyel1myQN/qbXFz3Nx8qiH
zc/SlWuP9EnM1CUpKpsCA4J6UeXEsRUZIDp0sPJng4fDEP8tAIQ4lzkzl+XI54V8dNbATKPmT8lY
SmXLy628i2C9uJzxggeLO3kav8QGHdhymhHuY0Yp8cVlwRBnUSOsWM54bMz+P/3VIIaNBhsG9ieX
+VXH+f69aboSnPNxqC8xKippKdp7VZADDQ3IFHIxzdCevBgtrtbjMsGzjIzOypb0TgR3qO9lG+B8
rETFP1V9Dlb2bIJ/kqCWinsADL5bN0n5NZ+TKe1b19UIgHyZ3xdyekYEqxmP6zphhXmUu5D27MQq
4kXTFisGJH9hIotY2ZHvG2QCaniy0oVrFbqeAhBjGFis+iIs8V6dZzNmpahjDg3kepFEtrFL3EaV
LhnN0AhaUKqbqXd4m3gktJYr7sCX6qTka3fKdeX/U+FquBpcCdYmhpLBmw580RG1SkilDZxEqXIR
eHDKXBZ89y4owtw4YtwZGxIRlLev2+QrB2S8DT3Nsfetv0PyZgzXcS9ywQ1oCiwOV7KzRcukpnSU
x3qhFVvd4JdiRW2jfhF4nK9nnI3hJEPkSjm9zfG2MM1so5tCbK3nde8sAKAauDBaQ3YgVVktoTa6
8ZzAbLj6xfE1MotJgLJDtfYYlOGKWdzM2JPezsP4bUuhUHAlLklHUgssqDaUEYlKjTsGeWT7ZNpa
quD+7/SRJ38CYktA1ASan++Ztz2267aV7j0H+qyPVFDXCms2YBtWKMhR5BoMiRuga7i2GlqcoPjO
ilg6zUbS8kLDoPRkaK/I2HjHztlzUD55BrR3CmxHk4IpllLaenQiQzWxjlUDCd0GBy72/X5iEXpa
GGSLWR+pwcCV6ufz4wPDIi5r+cAExRjZNPht4LaII/KFinMzLketuda97Q0yTWa+Z9N+4IdpJQ4j
rsxVixB1DES4nEfJWgcF2FY3NVPaqo3v2lNhlCGVQnzKJIRlKhE/33sWDHAgrIyhNKGUeTz7aE/B
YCUBOwHKwVuRgAQIJhv/uhAhClCxBahTlMlYuJ70eJlTSU7oXblzknl4Yx7OwEprQbUhIERlHxD7
ikBS2zE5HQFDYHDlr/omFF6+FejGX/ocD6I+Aog7NYxF+fK3/hO+L4PsWPyYM8oqf6/dgDUzYVDd
iuxFz0egVG7a1/azE+/s1kJn+CwAmLeFDnQXnE6FFVzNL9kXnLR0mxv3rYfhhvhah9qPTVt5jmJP
9Q33TRV5tjgCeZupQHD91QbmTS5Lkzx8yjsXcjkXDcSWW/jHrWTe7ZMv8O4JeXuhqEU7M5lJeazF
GjG7yZB1UxfTO9l7xluuf9ioGA7emxVFm64ZpbNSD/5A/BLmU/9WgnxIEtHx2vvd6K3Z7yaptJK+
ZZmQ5el0LACTl3j/AVkQiHi7Hp+B8LdDiDUasOZSFJBuctpL8LJNTSNQaMheEok1pZJate/x9Sfz
3NdFqD8Ew/H4cwBMOWA8Qt3XK7jX1EO8mPJp50/uc1AEM49s1gr9We3yIuxr7UUJRK6JNVHBmqhO
oEH9Kl9X7vnSY/MF3oz8DyLjQVvkM1EunOwnISc2KYhUjgAgjx8lcyBDMdrMNhbDZ6i2nC8xpuGv
F1HKD2409vaJx6VLoI9pWN8dIBJrQTOPbcT0FFhE6CGBzdQTCC+yR8G0wftwvR7qc/qBuLe9uI5B
MDpWXl+1kLS/h7ZoddPiO2x+yhmjldvSsf/BjsaYu490yvLT9T/NJUMRDA3f4lxIZQmdkB2U+ZyD
5KVbfVn4Fvbf+FgpRUV8ouQz+eVWSKOSSoCUySWoh5ABQYafjgNSfrLcaw+TfARBXEPmiabEb+/b
dnszHeCEvtm/WKchOJnXbKvgYMboiGi/sFGeUdpqYXm8TZezz8vSmOdnlHXVHA4r60jfO0zRpnwj
xGutDzhTeVSswjc3+0qA7KbioNJv/N7GwJcrXpv3VIMfwSpGK2SIfhm+ChY3HF/iPO8diWFKbRmJ
uPqOukoBo63oKb0BOhJX9rAOi7Mhu9Fz6nNX0YHt+bozVT4CQPz0hPNj3bCsR+RRItgq7UmcDGDy
/0GRSNPqKryiiCXbrugb8SwvStveoWOuQA9XnRyeBkSaoofJ9YCL0+0xEF4O53HjK0IeyOZgtij7
YoUE8dlVxGAzn7biGFgHr4aDHAq3V8I84Lzy6mrT/5QaoQ53JwHbf/7H2eH/X96CsEdHriNXtCdK
zmeCJASDDySrBqW1EvLvCew7Clpbm5Suqhw+xAXwEmFz51VeU7IFyyyvdg6uHYQFbJgv92sPACLb
6LAzI5dXgqXomSQzr+Uj0D4hIXwhC5Rrsjhi7uHEp39nfkMi+WDCjHpQsvcD6RDcfiKBOf9jreV4
ERWVSLoxjzVkts+AoTz/LPMIjtGAJDi/cBSym8EVWimjYsl0LhWswC1HuOzX3an6TFdQ5RYti56z
R4gkDdLHkC3s/csK0wxQ+NGq07NRribvtrsmcgNKL8rAIXz1mBXSpdKzKpPyabAA//M2qpVRM71c
uV+PACWyk2gMWR3IjycPMj48X9fpvSuoG4sssHAb7zqDYp3Dj3CCbL13lTc84yMaN4F+yUQIPfc/
qtdEsdYeH5iEy2Dux/LJ2AOio5PofLczL5vvA5+3mvFbcEsd32z3UMXTG9xA1Deafamtbfvq0t17
IfgtghhDSK0b40tcjgGbLr1ZXnqZ8IxA62RaCku1e88vcsMgqWosNcUm7L0mlYGKsxC/JYhipDI6
bquvCDGCpTfVz1f0QqdTMOhBmB6pFBnOicKSVNuYns5aPSyf1z/LGsXj567kO5qC2j62mB02VCpp
mRzd34QxX//I23RK2tbzA5lDApfIos+v/mbf6jawpwfWoTxunF7Tvs7bSLATGVs5r1FyYcXxe8Ug
zDXLRvMlDlaenTEGIOYZSZ8q3fVkiibiD1ER3Jf3whqiFRoSTh0NgA4Dwt6v+U2KpcROV1fc0otl
CG59NZH97kwyIPJ8vOd2ktDQIPNONsj6ZxFACxD66MRN0im0O4sInmUC4dvoDSSNbwdrnBzd2HJ2
7/Kz0a2UTMknBa6BCM6zEpSf0E5gwszvFFn1TpOJNnFD8LQbkBC5MxRBnN6WT5NEjFyxqskNUQ+X
l3Hh7jasOiU4j9lUBW61G0qaglhF1UGRZXqb5YSZ1LwyQIaMeWQh9hDtaHe8BIsI4BSHkC/gJnIh
r80nCNJmAxhudgvv4huWnKv1qFgaLoKNIBJFg/68NnZPBvRQUsHKDdrQS13srFKq1h3X0dyI7nSX
6fO4U32Nu1QVtX5KG7i168zjxsRwj0Kvv0WeNonlN4yRQqWxyeHjsO2z7H9z22D5SuxEjKfCE+FI
j8tJwgtQF7jzgQG0JRX1e+Dxi/iIrtSbgiesLkMQaJhGeGZH9DD+SY/dUUPzOroDoUucD7wzGLOp
CeZYaBTVNTX0hn1ihLqhzk+TKY/Mwp9xZzAQhq25MKvQMBwJ9yLV0kQBkj/x2JtKNSraXh3yAWUr
E3x4BI65TgmqZVzsH9X7sfKAUgyuakVuFlCFUR+q3AI1sNIMCvsCAFqW0GR+C7aegZRcsa5J0fcH
E2tzYWWW/PI3lY/6T3JNKanuC9lutExmYXIMlUdERWm0PTZMPvtGWR3s4qN8U5i1W0Q2G3cDY9R6
vX8kbDTzC6TN12TfUjadOI4t0822xoDisqVZHBFVbe46YX1V975ZZcp8uBQ2SskgdEuJ16b6s7TI
FNzDmEJBYUoqL/gjZLnc+1fwUiwabDWBENS+z5xaBxQU5xmFOd+rMANDfoG58Xx+JnWa9wv5t+8f
4EjOX5ewBtDwhKNUE9ly7ywwaBiib5pCG/p83vZabP1dBnO9VDJH0PdFuAygElpc4bHAsmKnQmDt
2EYpGyBtoLtKbR9sY/PB3WkpDeMfrc8CtNX1vTT/dDhnkeftjdt1w+TGYUK402cHftmDtHOY6sVE
LUvFrG5YRh8He2U45zHCH1qEIqwGTCuWJ5kkGAqm+ohueNJG2aN50ExiZxjydQAyOAWvdIBcR4RF
a4NnvMLEdVHhalFhpcb82Zd8u3DGou50UjbnTDGB3yp0y/Pu1maTUz49gtA66965jC9wRPv5LNum
5clwrNv36zfKpgR+liWJFRCp1beUBUwshMkFo+KVO2RLFvYw00eGGvZJ/ym0eE86o1CLLHBa/u89
uNM2TbsbSxcRlAft7dHZp1a5UwymRXSVxXqa9yAgxq0APLBGq9qMyTuw3n8i601POrlznxscxdGY
XJE9WTxWutXPvPsAg1ec9r+r6XDvdnccFn/KyEShZpeboIYuXkss2rgySS62eI2zup9QpRZL5uyc
5V8o4FNjVn6Ke5uvlsy2ssxkpa6kKhIZ5Va70Z9YWbIU5furw+D3lPFWqfam621WQV2n82wfhH5J
23YpIIlwJigyHN5Noh3owfO9NVf493OIgAf/bXMVEDZhuXwQRk4fG4aG2I52VUr2QKctJl2ZYHQ5
+AHVMXgyKmhyJ/BC2t9WoyKAUv3GcvpwUpXOoJ5ZZczbTxGUcneN32jODNtVNd/qrcXwjqVZYzz9
a1SKlIX2wO3jlr5NiihqwbMmQxOxKi+kdSzP7lBbo6C3fvpVq/mUfu/y56l1D80wez9mo3VMXCFG
baeR2UB9qURGfaQoNd8YejhgMe+gn39ZOlRSPPXYMP1EzgJWU+j5Sf1vWREWQyjxdLRXqfOkcAPa
DHdkglSujun3n2Idx2jACqFU7GgVIbfMIDcyUBEbBNWBiKMUp7AZaz0TMBz2WfBQSxbVU9H8sGAK
r6orGjL/DiQv50Xf552XPfF2IsJJvK4bLmWSWIm9kJwuruBT2tNjmRk6+8pBIf7/vs93Ovir8/3w
0J1mt4qY/C9d7mfu6e/AeVcfpgqgNYlBnvXjNSh5y+cEIegXrU6ub4YhPFIROZTSOf3o07WZMgRk
g/e/gCm4HJF6VBX27Wrq0APXe7bUdhm3XLIoFEverssBi7/keOFssPBBM6joX4v2WOubdx5ZqwAC
eR7LOGdR8p86BobX1yIKLKLzj4nz8oORZcNHkendew9Lb1gXyk8Is7l5JHv5AOaaSnQoOYsIiHYS
P7+KXkr6WBj9axLASNHEgGtU/aBTkMCh/C7Qa/vfsPXdo2u0G+KFK1AL9vHdzxs0hZO5e8Y+1fCq
F3jGViL9tE+GeXsnaUk/O14B3GFDAeRpwleiy7LndpRmmwOwMNRajeYR+/QInhbAYp438K+O3VsB
8V0k/ydIH8Qj5M0GkqUo1CNfQZgCCIBaF3P2UI21BzxgOLlsUfllMO125euPDp3GSB3iXhNkCgX6
xbrliyCkTDvSZJ7gHlQ2iawU5NAK55LgeGk9WWHp2l/Q/W+PA4tAx/iFNiFWXCYbm+zZ2793bm/Q
lEXOujKTliOmi+tQhHikrUNWtyyK53JbNZnxGt9+07h20KJzaTxGxcBhyB1n7zJPLuMSYWkdHKyb
DxeicE48BMvsX4Ul4EqDnKUl4PR1bLDk9vvJLqOuFbLblcKpK3EfDUXS3JfRGEOZtnYb+JvjYVQ0
bC1U19AueeS+hjBUgN8yHX4aU4W7EQSo2lDhD2rkH4ptkVH96hDW8SUFjJmhBIQgXk4DaOykGYMV
keeaRQSqMyBEzFO4zymD0WsOckFsgBCydKgatcVTR7bV4jHLE77AjQzlGtbP7qXOD1o8cRZapXkR
C2mfEKuHVYpTxHmyEwri/1XoDaplUgqrXYXBC8s/a4Xt0TAdZeWW1TXZJwkfq/tOB+wvZzh/uvPm
F0f4yZ9poXoiMR/XCNGcCWuK+v5X0v3m51BcO/bM3in4i8nXYKbO1dgEYMGbfKImqmA0xC7hJxCj
O7RAaun0Gk1yUh9btyT7K2HPzyIzNES2ZGkm1pR4BmWAzgnJFVzKL9g+1c5uNlr9qKsPyl079kKa
vc9Ek2SBfatW8WdWq4qfb1RCbJnu/R7qr835PntQiWFQs00FkQQivBM2qAkbxn7PRg2m/KT+k9pU
XV7XDAfDZpnyXxpHLZC0Yqung43bQf+HyVQAJ96ntBNjSRlNvnzz/FNtDQKXEOHBfJ5vnzQ6lOjC
z78KxEJi+nzR0IK/Q4vEF1KJ2Dfjlg+DMIz59eAma9qD55WK20SnoADbyRWlyqgx0YXp5OIDDP79
4m5axbCQFYjUxPX9b24KowIsfJO/QIwj7priER0alfnPI6Ith4ERtoz+VY168EZOBob7VIei9CyG
vR7doslqhmOpTzlLn6443oKUtydzGoJcr7siMYNT2enj/+GqJoHMj+sfY7ymPfWyhxan4IXnoW/w
hWPM0tz49xSbfK80bSrLJyDIY+eSKqX8GsAYRnzi5BV4ApIoGRAqzlunRduiDfn0eANTiQH+Ugq9
/ir0GkOKDMtaicTDBBdyLSfSjqQLGY67CLeOTNrj93PfUhUJzOu/KdxxK5R5iVyncEIY44wpaebW
9DQonDcPYcZOzFNBRrD0prL2CtY+rhHzhGCeu2qaR1Z39zUu0RAJhojk/89YMO83uI8DQeA/t+9s
FutRMDQkW1c7BP8/505lT/DWoeEaHXUfnvChyOZOiN/UkCUx6fIxQYS7a0cE7eA+wS4JUeV0x2Ua
xP4tvm6qcKrPLuILqw+ElunexLFP1VSAp4h7OnOQ3oMHYoJNrM2okVRvp96DeTI+273+bYTMomXf
6yF0lt0fHklq0TMK9TjWp8qqsq48vd9956HY9UPfhvQFXZp7qKpwRVIuU+BrbOpY9FNio/ExbVTq
gxWdXsqGr/L8uXItsWEs5fiHvtkknZL1KFbLrs97PBtMRFn9QL0v6PssVVTilaviNjHL9DwlULpC
7GZdxspa8INvMsScQshansly4ktX/At2aFGJ6Bo3ytqcdHENQLvxz+bRjjpGXee+pgHv8nXLJCOt
Qu1Qsmtar4fv95hscBG6tSSeFV0mXOLVPTQDXqCO2S7BtkOAEbeX+sMhojo9RpjZFFPnSaCC9uAo
t7niChNRTBts/eUWv+H4JMpjjzLNj53OsufRuttGdzpDoGFixdWJUxNZdGUcngEYXWpYBL+ryh/g
q+ZSqByXStdSTQxrqzGEHJcaiZL07q8UY+6Lty0MbICGDGb+BhIx2S8GZ4a+zbPfMLBslvr+x8W7
74H3VzZ1Bp9H5UmbYFg2NtYfTiTWaI0Npvq3v5eYTzGBjhKBCfHLKOuUhyslYPTapJjGmHlc5K5+
T+GkVdFvfTZcwJEXAnYaclgB32bpn3Lg3fDAMURo7cqbaDjVmyTLvWG5rMSLbpD1TFhe15CXNAh0
kjLmWM0UGa1Go48dCFiKL78GOw6lsv7NriuoMrANZZ/uaHL81MmI6Z/8yCBGG5i3xBUGrwnDFWLU
1RBawKdmlwOCoLvmAwHdCjLI6q1g90kiD/kyp5Ib0nOAbOL3Gzd5vtWLp1k59zmBiUrxijxqDP5m
3g3UJdjjRaE4h+zW650cPuLuQdVhkVH2y+GGn5601n53QbIhp2CaZC76CM/qFZ8mmrt1QPEavqgt
K+7FUryoP+CX+4bUTAa0u5UC5KPtb3OBNOmd39gVg4ufGxZxZ0MiOm61zasxcYOV4cz+XHEPuEqK
xvtX6XP5+dl/uwc38DP+uuuZG5TLbny27Um742V+B6j/d18W8ljYTBAr2AewclC+GbmLDqCTjAGz
qFpbhV3QnGw4CQT71lgCcVoPpqSeP3e92E4RySzPlgx9BtUPFqWY+LQDJLnvXnQtv6+hqWCJaSnO
weLtBCXMIv45ZdwP3m+xxgJuO34+Bi0RbmI8hoDVP7NPc3J9P/8R6/YBy1AfYn5OaypZtlmjjKi6
vhYZhBGz+o+kr0XlaQS5ICko/L7I4/Q+UajckrgSen/AKSxDBXeMtK3Utje1c9Gkn16jPWS5FTu3
bTrdx07ylstGPI7FSihhKMlVeq6S00AvA4H4+qF2uy4QllCHbEzLYRQQ7kJxooIqz9cpjPNs15zb
p5YCQ+HuRdcfF0OiMXBG148rtl92TqHz8y6VmKjpqZMeYEWkt+688cBDrjhJaoH12lstWvG1GcxE
S7nFLpZ2ng5uk1ssowhwiB50R8SD4S6fG0EGcWvEwhTG2vYqVpLQgHL8iJ2SCQKtCrljY/PD1Zm2
F3tV9CNSLyKM3Xo6TR0CLLIDi9vtrmXfufh80Hpg8gpljagO4H1tq+AN9tsTA6j9llrhYHi8ar4h
AFJAiIDbC+OorlTqNR0e4B4VZUT/UmjUac67AzBfYmtnz7tOAMRnpDUcfnzqUSnwL1VBUXCNmr1N
NmHfQ7RQhr/BptX6XNmYiHjM9UScdWojN+zCtSj9ouSBuCoh5fz6aSpvGciG4MhC8XKbC3Pt0bhG
EzmRW2pT0TWq5T4cFv7YLzyn6Z2EiWQs6noFDfSNMlJQHyNr1YU+eaeWJALv51clpq+Q+MSPORwQ
oK80nSVpd9VR9Wd/+4YrVJzm1yQCDIukcX8XmDnPooTbBzdQxbsvIYdO0AYyFdMaTSzkhw8nRDji
kiF3wStN2/rv4ZNjz0gJ1YGDUhcAP5NVq4EK5qzZghFuyWBL9C/KrNxyPBlXGR94g4CoiqpFJUJr
0rn1HRfqPS5PrJ/9qBmnse6gCPAxrS/lMBj07a1pHlMRfEqsDsBpnQc6qXiyP8UVD6BXSveo3SEJ
dRkZbZaLhv/1HDOCQEoz8WODQiKbKx8rKr1DLsXRBTWW7TH3bRNgl2/oiMMKGtCsh6zsLYDrOqL3
N1AOBB9sESIKu+Jq9nJU0kZHSeT6+qWkm7k8xYE4nDbv5X5UqCa5jQB6zL5arzo3n5XRsQr5DU7m
xIYLoesqbb719zzFvrsbFIizSrKuBlYhnnyBx+sfJdgeHawsztcjlahipyzuZyx7lHEM00HPGgtC
XluZ/YkuRT0WJWHmV4buk7ruStqSlpwBmJ5CJgtc5oqa5HU5FwgLYnCsKjOJXv1yZR22X+yQ0atF
SPdrjAZVySTuIxmOOkutxHnbvmVvckhy9Tq+ij1mV9FX6EAx8Hm/GUnYd585zSX+sSpQUly0HiMo
IJyJRETJS6Bpxfb1IrVVzvZjVlDjog4li+os4KccLqX2z240fDhfkya/5OPSpKo401Pzlu1KC6Kn
lVPNx8D+sWjrGNVLoxdDSXxX3axTEiFxU1+twJL0Aw7HK+TRMxkQrKJbQWGsXNpvJGTlB9CgU2by
gE1FG32x2kqFXSHpeqmwJnnufdRysNb9bpCw/fXdFdmEN8q2S+mHUOq0e+EnLZLvOeVwgAYjogT5
hiFfexNTkZPxm0l7PkiW3nVkVTEdxArR4bqUTCtQpVYgtipLqw8tFo3X1rVknDB7JgXaVXa9cGGK
WB5+hAl8Xv7X2eT11jHA943/q8KFQghNAqjEAT6M8L7Pg63Kl8heZSmFmGZ8FzKIFKZMWdBcA40+
/3HJA4LrB3cJ1FiWywQES1y5c8S+4skp9+gXNUABjZaPj8KtcSOfJHeny/+UGsoCfAmvH3L3e/Ua
uxge45cergkcYEIkT4TSe3qsom4VyH346YkN5DlhxMxQHG/qvqHVtpP5ROk33a9FR7vihIdV7g7r
7/JOWuc0VEiUDIgX0rz9C6FF/jVQ0olt49YUFMZa+z1He9A1Bu+Mn6Z76fKZqQz8+HEUOgBb47am
EKGmmuzraTWeSXQBOHzJcjJdgdHZYEyg1n3VGPkvRvR8Jl9G6svWYrn2XcbKMPAjBA/4X9sRoklc
4eX2X+qBgcnvmlVMdt1JKrUMV9NoEXGGi+TuWRzPzXploOCihWV1jR9AMvenSX8mrkj+tZMyGgzY
iheErx/zyYwKSwpvu2G+ChUMXjGAnqYVxJwaBMa+3OrfwKxSAt/bwq/d8VHMMgCUfalqWU3kGie0
Wf3sJZltRM7AHNupbpFSj1Y7Ihe41+cdAIH2kTKTN36Wi08DiOVMoyY6kUNbMc3CV9D3Ym7QbU8A
wcTSkjXlcScbz03/FWIIgjTi7s+ZBIRwqdoIhpzIA0XwECFD5l4Ij+YfIb1R/o2knvhTgeBC/fEa
+ouyDHCZ3GoSwTBa34nhb4g5CoFhPkp9berNPwbEQSzecy9QsN6t5JVwlxjDqEEKUFz1RFV134RZ
PDf1uG30Tnwk85s2CyLFnqygsX4XfqFjgiyks9vIt1vCUXd8W5fC+iYb5MxKtbutLFQsuDG9Cq9w
Y7jxhuGW2/v8ynMsp/nh917Y9PWPoP2mMFT/ZVSNl8UlWu4rs4VIqZ5VjRcxb5FBCg8nDCoLLnxK
iJWKV6aHkQFXg51n/WVp0C0jQMx2gwiW2YLBTt5PUNjprR5cE4gzOta9NvYgMScAE0s0/feaEL6Z
QhN1MVr83fx34ZfB1X8xtLSVhpRbZMjigngicpZ3A8KzKHEbpSC/bMvOpQITCdlLfpAFZ/khjEQP
r0zndwgFtTzQCsyoCAG9dwMJ10gq1NgUfC026WeBSouf+tbzEr+ETJFEvYF+4HmaBkoaOY5pKpZV
tYtCX4zUzktU/jmjhU5rp7lV51OdMMcUoh0gkdD3wae49cB0T/zCrIduQLsbanaq2hCBr4llt3jz
brfLF7LC/UqvT8/R10yQ/QVkDDMRE2RnLd/gUowJQDsvbfD6V6Ce09Vjdo0pRUpidApBHcdzaUb5
zKz8tlp4e6LVfoq4C97bOX3jIYG0LcvZpQpj/4cuXN7Ggg+qk3nX9c4+mvKFgTKDZhEUUFh3MO7K
3F0Sn9CHWpASpfvtQvZUx/tWwURaMRTY3ZbAKDRhbS7brEGARgn71QUlI1dXNN8qW5S1mF5e5gAY
Q06YZP8+RpZLqM7kXip9B64bbdRrlSEOruLcdQ146rj1As3cKAIkAmcXeQRKWlLd0Ypk9fYycYng
jE1FgbCNuXAjZBmcvyQMY/stOxXX9+VMq2uUdg8TTal7aRZPPIhmklF5iUU/uKhzt+r11hTX/nlc
22NkJFdR/+TfusdJz2wBR50keXRAB9XaW1mZQmUULK091JQwS4RWl/K0zlAsAvO6Wh8NguLqFiB5
G7uYzxLO1A470/8HyGFeKjXXhBECtuF8i7uSNo1Q4BIg+VSBUeCsU8dqWKiERElamyz+rRIkL6TK
mJSjmMe/P254UN/JqKCCSUp8e4xpabYAAO9wc8F2D+N2nb79PIocjB3aUPI6q8iRc3iHvNKGd2DD
5uZ3bUPVUYyX5t0pF4gZYcSNpJqQlHyD4lA+Xi+4JxmD/q50NRpfgpvENd2Gq1iaNuxhW4UbW777
9WjP4qiNVPNRNBeCvx2ieYw6cBzSFY2w3lZgoR+KO2a+epmmty9EHZpemVV54JOaCu86uGiKqM1F
yv5NjWJlO3XRN7iG6WU+6tMZqe9X11inwFjhzPQbs+Rn5Weee5OFsiFIAsQKatTJMWynKS8d0plH
Os0nbCB6UAQKg7iDrprOhdraCzf2iz9Bh1AJuoJFmeIgCciV5I2UVSBq+C2ig0g/oRS7BPuiepMP
WwduGAofceLq9eT0bS9lRrGFbDzXZIPtAKsATfORr5EFe0oEQM0htFBbvr0kv/InDo9w0yglj/hc
5CTvQxOAxoEb31bfFcOfoh2f4Ls0+hrdLVn0QPCy6tK6v6yzGHvrsXJ+oN8A+4nVMmd0kVez6lrf
4ZTc/TMZfjYDX9ER7vTydNSXMd6XxCljsLrEzYrN+XNF5kjWLvKpcXlFn0AfM30/TBdbMv5Hi+it
at3wxVpHlNDAyC+FsCvsQyOTk/3qiPvUXAhKDFk7nct6SKLhXEXp4Pso53gIFMcY+apo7NewMQBe
0deDIMZ0WHuBiMuABYDuUQLcWr97fNLxoglKWV5m4RIU9invdf7UuFIT8WpCV46/QV/8hSsoW/Xn
c7uMwNoA5EPuIIJWOuJK/mtpILNYuoZvRES3Qo7PHmhaYB1Jvi8U3oQ/ALfDskzZTJBxvU8P8E1U
lnNwkaoSQ/OCe6noIWxi/vb87k3WEMqDa0fxj6Ag4WWk3pQct/2VhXsJS6uFde978okKCRvFnzm3
BB0ACPQULT2bFm/Y7wPiy1TZKsvXcm7LeD/CDigwnsM28y7QQToVAB9RR6C4tWbgkap0AZVHqxFb
UE9eHbAG42jeTkyCnOxNgVWjb1JyoyfVdI/7oIyZt4Wrat/qtZRcBH0sgXjJTF5gp4rKR3gscZuA
KjFXHlmYW4TNGLeWaa3lWKnWlnHf6N3yGVJ/yFl+vWyDm+ihZf4dg390xrnvWsY7DSBixrB/Yyhg
y4UxH3wh0uDQKnV+VwOGV69ii1TiJ76Zz1xkls5+FnJGFLJwgJl2y6ozY0vkm0IdVeCw1MZrmfm/
5Hik+Yc4Q4lBloB+qHTv4VJk65Id13sCX9VckaRAn86Kaglw6er93CF1V3hrDBKdiQT1dFV0ECwz
YvkYSqO3H0GDdVsGeBRqUVZ3B9XcK+wELAH4LW+ERBi6om/oxhhwLU7mNhf5PaMa/YQykOYqSrE0
phwBArwNvZ+pFrzjlXyfPwJvZkbtBy9b6VucjMzi32GyPpGQoBGSnYxU05i6m7wJVHWGJc4UMTjN
xLkNAKYxtKXw9mCFsn23liNgdvorEGwBEsQh4993TgmLNeoSWCBFbiLF3cN8AD3sloxJ33G1XJBd
k68X4IobbLzaiSrWPnkATSEXSpUWPxPekh1Oyp234m6Zxr8EVoESu+CNlaW0ewHFAUNhWlHeGe15
u5lcltb3dFLQz3OuBEVl9k4EapDnWJbc6PZLr5mEMlgXbGu9W3H8CwxqY0n0SKjOqn0PfvgSfAX3
E3Q3U45Wv9buqJjkc2INR68k49xZ8lVLDG8UhpgnUI7pbSGhlWMKpDHtP8PvImVsp4KNV0GYH8My
DnutjowKkex9zYoiCoh10vu1DnmI3xOUowH+UA2VJgDU5VduJOTrFTJxblUfbNKz1FphRX4tjfWX
f4CDUOUaqWx25oGuFST38c8cV8E1gsB6JlQbRXTXCs7ugvY1B7HFMFqGG4M/zjeJR9x6k5YecSMF
DI1g0uwKO0Knqk0K4tPaPc6g+bb+koXuv8paZenDfJqxDZ8NJBLTroFsxwP/kqx0jaRG8+miq0zQ
iJGTuOFBquJ5VhhCtIprp1bSuvdHQUeVNmC5PjUByt9i+YMFa1bfCWjuL1T6zbeYEWSN6NSx4u94
l/ReCmSQPTHOfJ3k6MjGnFvT3AYs8ZFu630T9JGtQNXGihrxIGY1atLBwk+2OJSqRzNhUNg0q2Vy
PwPwoT5R9qqBZHxEcWoFSm3juVM7pUf/ItDkNYt4OdYnQSgDGrvGs0KwWUANqj6wD9LQ5WssVUU1
9dCHIQK+Y0xDgrYpiU+aub11uzY7VJP7DuQBTj9Ac9jMKBQPFCklPEK7wAm2sHw7ghSMAN61Py0P
qjTSMSHkXqqkv0mlua35hOWa/R/pzm0tXCnL2M0rilUGvnK5R+TldXn+lJJkV+w4oX0CGKyYy90t
rDqPi6uT+gzXSHO7Nz/OaMUq0OuDRhRVkgfwjPtXvW4St6NBnrHTOK3IaXuT9nlNefJBZUofo+ns
37O/Nihd09Y/xG5Hx3VGYNgTm1Ju1M8ADR8IZNg50Z5OpWCj+ilHP43ewnxr7cvWlHBqNiAyVA9q
HqT136F3HPAKbat7e90GKA6NHRpmlwyH1n2rNpeQLD1DtYxMAhnocjow9wTIu1V+Gshw39bbx7Dx
SDoaejpxpMCFPBC6P/gnFYG3psQAWjg//EU/oMjwnEsUNKz16WRiwbvqO8pc035fuE7nTs5RBF4A
dxgkUzKLQbo6RYQigOTXOFFq856Ve2l63f2ZsC+kNWkt4WuqfNFWb6vFiKA3NoGM6YYuFYeoOLnm
4Ameobj0ploNKD5X27pLOEb5uXRWpz4R1xVdMKjLVRpmUr3JFLkv3moTVq1fMR1K3nOc77JExDA+
c7oLv9m8sQJJ49PGclV7h/+pjgvSMh1NidpCH8JMFTzkf2V1bXuQqqqSNZMbYuTSe3gOTWr8/2fZ
1+IQld4b4CLSrdr8lpaDBzoCpDRfL4DxdPEwDFifYjfTVcI9elLqLdSXiEf/Tv0Ytjkxd1KeUXf/
rdGzzf7nOKACMvrn1/GHVHqsK+Y0zJOKTHG9GtNnfcIMzjMhE7kNaXFZRBNohxux8H740+M5EOl2
V166li41nJMEAqxr/1AIqGunQZA4xWbHi8SGiKq4hWd5I2/wwM81QmR/Qg6W5e8UMncsclA8iF6K
JsZ3S0UUW4ioWG8uJm70k8IIKYGxBwknftoVqX1pbkFx4tq8NNGp4+HoiK5t9NmA5SuVUwVhR+JM
Q/TM+lQypy/Dz0KIJmu6rDH9y//HRGsUvOfCGaVYKKdnVf95oVrivT49RO2+7nYZEcLdn9TRWuXB
1KXG6Pd4UoaA6VemD2p55IzKoFzqSPiohqV/rCC/IyRXdBxP1aF9LfpPUHRqNSjF8MPe2El41akH
V0lwHwEVBMtY6Zs0tkyGM6vhdWMf3/536sMmEg2TlDe/m7gw/REJp9Yndkl9xTZSlfz4l2fBusAS
ahbFaBVV+d0l0NH7IYnIl2jGfggCLM2BL8iHG7/p8N9CbMi76qLAJ6ZvMCT6p43r7Syl7+LnE+aM
BqS0Y+vagDBbGXILz/dWT8T0/rRSBfcT10CIvavQW3H8nX9d7sB41qQbiun2AA0xOtfDShHZF2b1
LN3DwawAqDdKMIEG+Azrpu3afCpHCb3MwqOAYCvwheA8cp6UMNfwFZS+ysY61jS83x7/6GtZB4+l
s8XjWbPl+jo1ZjhhTKRQgE8lneOqZBkfEe7DkLpAH41uOJVX3Bp9dXiwS/tD1G/uIk/FuXYLPQli
gAGbtxz8RUvHZqHlS70FDPhxZIbQz9ZyHdJ5kxgwFNMphxYgw4rwjyVdGY/1qvbR/lo7E3QOHzbf
ICE2yFwmYP1TRIEsuK8noEf2oBzcuneVBw+nEbTQK9oZQyacxZjJvDT1mSvAj6x2BZOCQ85w9AzA
qxPJqfwsYcp83bOgLsM5vIFiFhCRzPrPUI2H60hIEt2Zu21qbTFN0lvgLLE4Zl4fpXwmoMoRaZOT
QRYphPmFT/ma4RB//RrCU4S2bq41/hxFHKsRHWGKmF6LTf05IhfUxvbNlH38dMiSMG89ZrATffcF
WT8M4gZ3w3Nk586YQpCjFYRuLfOQP6pIWuCHf9YNUFbuAcXglSdcsjCCutOgagY8er2G/rpIyv6U
m1wxX4UlUJWjJVnzVsq1Imr82axjvrUZTO3FdEvFd+OvldbTcF36HuWcAt2PVYCseUG8JAzYOtiz
2cFbSmiZr9qQuNobl7+WgGcbaYlZLpF7ZlT5YCMNOWUSs18UX3+J1vwqSa6J/tEoNVCbAJqhEMDz
Gep6N8cxmTkV1DmoDPCeWNONmh2pTffOK5jyhC2x23q0OW7TC3MBChloPSLgIbyi0l+wAaKQ7N3X
qMChIMDN4bhagKGtvmygrB1EKQk3B2DC4Ppdzg74ymSzT69DI7F0B9dV2slGAfv+Ni/dv8UbCr/R
i0noOAbExf+e9YUaK57UTR5Qt1IQ9P2K6YJPOz3A1I4tBH+KUQ1kSS1zMFNf9E3yVGj8O/c9nUEe
FvRfJsDAKX02h4KGKSGgWf/2AxU062Xa11lJoNWE3btbOnAvpXdT/3mAkuD88q87qUvLpp9/U7IU
6i/Rs54S8/He3ZAkyfRpJCq1NMxYwRDMGj9d0f4wNXl7J9w5LCDmBwTaYjWygzsJkQ9ptiLowT+e
AROgcs/68kROLp6/A0o+6wXbivsOmDzYY+V+qac2MMULUfGF/vzAJX36YJ0qYOcaLuBBrwX5eF++
oC7KJp2W5ET8CliTLojIP6z6iUkdVaqHjp5sjhoztH0e6h+tEo7h/PLZg7tQ/KMrEewunOYh+D9W
OCjDJP9YrwUtySeo/8iiIsw1IZTPm60vfI/6hdzyBqkKg/1jSlZpsHvLVFeES5WCNAb0g01KZpKe
c7RBmBJTugnP/QIleBU8YJk7kv0AyG5R3M7UF1c5emyguMevUrY7El7VfX2v91eKtl0HWWJgCUIn
FcHPIRh6Ur/j/XAvLWC94Q7kzvJzRy6o6Y29iQ0AusO6RkFlcXPmL83jxWq+1fMd/ayB4htUNDHx
xSMjLiD9tuR9NxvTRhtgI+k+BXFfjNypIkSfQmLciFWY98h0mm4lL1ZjKG0IlAloGiMVwqWCFMdO
JcWweTg6E60uvVI1Aq/mLmFmKBRvrJ/KEAUDQJ4FDI3gKcVM8iUrl8Qo1SJ/6awtCYe/oBBeYhvb
brO5sXMn3FJtVeFx4VWBA50KBBEeD2Lfr44HUwhocYro/rBrtEU/dzmNX8K9gzP6oBczWBE0Z/P+
RPc1AxnT/W4EVbVflr39F0gfcuYqyApdYxZFaIfNosNmZNWRVLKBgTTUdeZUnTHfuQ6sb+fuvA2X
GUyZi1BmR0PZN5lcJ9/sJxWjOCs51wgT5qhV9sfdG/MvML6ObBsDDh9ThjVONZrBrZTl3r1moail
IjrXXvx8FZ2hmG/97emziZ3THJLnujIi10jJmBSxUPPTUfP1fCvJyNL6tP7f5NHJFF3kLjnxJsgS
3nVtdVZ5n0Xy0GuJvggkxuSTPHpEPqvO6qPLpXgJgaFt+aJbfuQjw8AcrzsYz26RxlJurNVjJbcR
w4AljjP3EUchMJwZmgTEe6xn4yDwyMCjlMuZHxvyvCIGjgyL9vaMqGeo7akvU53ks/4hH5Nb7343
m/DE1sNaZ5Nm6YR9xBiZSr8eNfIWiAUv3F1AXGbbggYdCpAT9EUI1DFlwg2uUNnIggl1KnIMTkSH
r1Mp7gPEnaie05gXUMqAFRVxguzwFRyyRAqSxau+sMSwsj+X+SgToor1PUi6XWyRO+v6twNQ59WX
xfEfVoFv+XR5gTmm8WcSryZa93H+P+ApcdR51OgrzQRlK1cjRkmgWtMHmv3mfJEVnkStAnaUyTqG
Hm8re8fC+D9B261cgiYKjKIEBHvq2tGWeLZwfShoQnt45rAl1Hm6IVzk6SeUf0hlVTsyBEt0XSdu
ucNBwYRzCV95PBsGnpPB39vTbDTvMcpokxHF+DR4kJIzCqhG+TEtBZzZMlMyrB83egAKh0L1CyGc
pMvJ+o0e+Q6NfHei7pLbLp8HLr40vMv+Rpest0pH1pmq6a3hY04ubtZBNUlIgdu6RqMysRwd1bfC
72wyThWprcTu4o82Y/dK7ja1ijoOh/a3X15r0E0gla4P7Fa8S2/BwimDLeN3/MiiLFOnZY7McpAq
zyDzwMG72Gbo3tVzWYtIzTPJIA6ZQx9i6Gu3idPGx4iSfAJVXsI+lom+OhR5Xzsp9j37ZoIRx14t
iU40SGv4iqkthMEiDvvdt1HmdQFBA0O7LVulAfRFwgd5xa7OewZieMBSiFBdzLaVcmc9+rfLzMna
UWi7+xF1gY4ZE09KdM/mbbuwDo6FEyJqEHYGwtC3rEo55+Ny7/pR/m6kiSMtTmJQEQwIbe8f3wU1
8pKTLqTg1TzpJJy/MatEFEECiGp0egwfGjK68rGiZtgkGElA/ui73ow/BwkEpGpxZPUQqJJmSJgN
5hM1CeC8d++QiEN3Mc4u5vdMUjW5qn63AT59wb+E/62TQPWQ+h9UM6TtYgUbgYZwGk+i/1MoN7zn
9NJfw6JRNYPAFQtac8sXBDqFfMe882ir4aypiaUkBljJAuNiF3m5QjLHKNuUDyMQ1GbFZlr+Zqze
CxYgA7DUvPUvTV5sJ2n2dQ71gXdlQebNzQSILNToUszgngWOuFYgoEzHFQsSlsE8pUHBlUrskbuQ
0XeOMqpCWi1x7ID/0JG2JBwGXd/zX6HUtR81AIrWXd4zG9CJXI9L6KIF2hrWQey2qWJZ1EHMk4hF
yp54g3iER3wS2mInFCcck1NHy4uM321STtQ7jdqMhWLH5RusnVObg9mU+rVScmsQI1FxFNIx7nlW
oi4zNSvDFrRTSivOQ/C1IMtOR4tASV9KZ4E+bEDFGcPvpN96tYBxDkHOQUJzECl6qwuXkWRdTb9p
ZAA+zSwiYlFF9uYNhUfgMJSO2P5/1NapfATjo7/5D+t4FSMMAB2Gu9o39qPPDCoyKUHkTYIzmwjy
wZ3LyUrqnPVssu/40T0wvWMpf+HU7EvD5s5fj26MnEJNDPLufOiwYbCo3kfwxj9MHKHTLmz+sN4y
2FWlMEJoHVSH28bisv6oMQLz/nt4Hn/j3jGOaxQ1BgbAx+WbSo89Mt0OYBJtPiXJhIXq5AgCJZw+
mtBIerk7bWIc8vrcLdcBo2MCCo9RHlFMCBkZmPCZQ6LYEODwQjjy6w0fPZiWSJ1F2/cDWKgd86Ld
2EEKc80ngB1h8/LRmZX2YOMnqcg1xeD+zo2GVeQQRfu9y2RXXlA6LZEt0BxA6xfgz3pRm8DCYuSd
X99r5CG9vS365gLsFj3M8l1QqikjJ2h5TvZDtnJlwQpK5w3IKNFWHpsVBli8CRrEpFGSPcWi4rbB
Xs7SU38FxfELYdBTkb/PBOlpd9bGZzX+83RkvVEWyF/Cd7zyU1gOuJCS3v6Fje6/K4kpVi+89LR0
sEc/ctyXrSSkkU3YsXAH5veASOUJHW0j0IJ6QlDjfbUKiPE0pJHJw/9daSCfnPd/T/bNSilhybSy
eophp43ItRZgtViPrku0/MO7bGhr/pg864gT0H4/mtHBAIScvLHA1RIXsks4TJaDJUF49Mq7zo8o
/Y5aNRR1CT/uXkZ4Dj5tSYkjzcPzVT9ZIQ1vJ1TOAG4zbE0aSytXSykcqQ99VuW3ZfpY8slqmn+Z
ou0zFlAQWDu8bMxDvod7RjNqV22Out62Y5P9qfjxPU1ec5cfAvD7NaWmArSV7RQXhRjUzH3UZoY+
Z1lSkngBxKVDrRv7Fp00BJXOU80ExMks4OpVIcZVl+/ekwzqv9xE26Gg926QHbBiqYizdAVerMGF
DfDOk7vp0/R7XxanCCdySD085ZWN1B47zFfYhY5CY8LGpFkSK3RPVW9gA4UoS0gutpAQZnKUo67k
tHjAcRGXVHxFsfObruh0kP4y/rCmXXpZs13U144bJOt2kqkmVjTemVBSqXMvM6y6yhMaOCbgIur9
9ZYMcOw/7aAXMXj1erLSicPnK+Bxu/w75o1HtaenpBjgiLmgyu7PnH4CiL6hio8//H4ylOYB1Djy
dSfEbSVR7p8W1ykebuIhbDs+2k1Gk2RgKjgL1HSRSvEw9y/K3/sRyZjTUZoj+wIP6w/8bpi3caKW
yRpoDtc7TWpaXf+MLdupHUv9BMvOFAhOEbMRrCj/vWV1/3IB7dSjJsNRi+BY6WjnoY9SJ0Lo5amM
Ot6+lyxWJMXgWYgBJZpGRGcaBavTLUy5CF+ecpVB4pxNbn2pNXJQ0mQtyFnokjVa2qhIywQWrabc
8SI327UFS749DCHfwn0GF/NHbpbZmWLkz36o2NoIRyz8wZe8s2E9ULQpYW4r/iUsaN3dKyygwT1N
aorpHBixEctqH8nJ1djRvfrP6rzuthupIY0IaSvIEhC6p6oYu7DkhhaEBrsneiT0QBv+tr5xdXpH
ArUon7/ZEYiOT57FVeZakvWxJ68UvCzLy8UqnzyNs1eCnOhwcYpYmeEgwUBb0XnMsEMaOWlmn2B+
D5mvoiBQkPIBkbjiGdAYvQS4d40543B8zcpqiFLveNFUHX99mxXxEqWPaRWRLcroTmNh7qM847mk
RYvzWauNfeqU719EfWaY0j1LWHEGx8tPKAOuYR7q3Kxk64Slg2TroMzVD8fvUfgqCwrwooFusHeB
M8421zstZLQ8SbkohWUZ10YU4/Ac7BzRHDr89Nz2dETYC0wwntlDvOw1G9JaYonkWqV4NIdsfXhr
KnuLPqZuFFRe5DDuqzAJVxYCn8xK5op3Xl4asC/0ti/c1YYIAAUik4LsSUvSI1uMmg+O7sVFGjWu
omGIs3GxQnaIT589+bbOL9HUm1oVV8HVC4/8KGlyizXluoDl8CAMvB52c9bF1l23EyQMDTZNmbpp
gB/j3Ottm6/pW1ORwjYxEq63DQcqPJ7TOgVNXATnDylG9Linlz2ySXnsql89UXcn9srRqGUU3o7N
cVed0f9nsN7UmBRZNtbeNnF3Nz3FVSWrEDDnlkOzIuK+V934GlJdPK2OPB/VoWYRiwRT0XohwMCe
sp1eMW2golgtZVHYAwd2TlCe7CYF/IqSOmNwUW64dlyHC4oAP+UMpxIfwZKAjM8qvUisLcJiY4VK
X2nFG/BLPrZI1p5PlmfKF4ivIU6YV6ck+xf4VXSjAuheG3nymyXAhWEmRyYOkiyDlGNtq2NClRym
YkJ260ZE04dQ4cn+b7y+Bp8c0yiIPs0RfL0P+cMjaSMJX8z8z+EPlYY8S/Y0qyXY3lQifUfXv7XL
dxBni4XPOK/NAF1HpVaraGfhymzGqeXRH10MUtNKc/h7lHVn/jAwpZabVPJphJYBfYO3/BKnadiN
LpjcWPmRlGbI7ZEInBfhp9c9rUu7YakIp+KJQILs2VYY83Xf3nCaDIoMl/hbPybly17Rvye2jTMf
AUuJWHN9k3X9wN4aAsaW+f/lNQ3oo9sw2zFVHrbaSimQIYVPBqBWtexRvdCHyvrNJC20hjUwbJC5
t2jvWKJ2LT7Fx5pSLRUqS54c6ID+S9AgfoRbLnplcLJAD6SMx2KtE+Obz83QbuBckNU3X4aYysCa
b6PWhxuoK1JIYgeUFCN7u7yZ7q1n2HWiHAEYNEhoF6egeXrep0O74VOmp0ugIhe4Y3p6oSoFuKot
OSgfJq0Qc8KoYEETNu9SPi0dtXkPw1bY1zqMZeY9iVYnNLLi/AUs/12q8wJKRHwFaENPpL5/7OzN
iJ7YIGwYlKF5WUBJABRxCAiv2PHd056s+ldKzhSw7WjHH3FcebCoar4zRucRy7nGzcRHsPMIVg8R
gdw4W8nNPIXP5UINP3niUP9tOcpwIdIkSNFOVYgeCCgEr2KuWQg3VO78D/3L+lRs7qLMGII6qLUD
/lDaSVIBH/YUzF426IF41DRR1ndfYalEuKg/mDLw+h18k+RuO37pF0PJH6T9YzRMcl9RPoww3yWk
hS/TD5aWMWP7l2ZAJ4+p9lpOn1VidotKx/oCJeZBTUKWFzIpJNX1c1SW3hzZ6ZTedqMdY1/B3245
igUcCI1iZ8kTm9wXZSWNPKkn4EP1dl+K1rEooIqCh/8QV+AWOFZ4M0Z1so6DHR5LQz9Soff1PMnp
3s5dTaNGrFYp1TiHxRmxjiOdCY4r6JFGmiGsxd/g3Xi5bBD5B+jCeiH73XF+RtdtlgQizkhDm46Y
k4nOWCSSDzBnS2fqaDzDxtNYbNcisYp9cetvkRyDO+Laa6szCwazRnlWkHSCDRGlp9ku2RFF+EKf
YQbpoXUbAdi40bf3ebv4Q6TJrD2JJSRW0sSkLwk4Bd+l8Ia91t4xXxVqJuu5xEiHfjbixESiJyS/
uSsLonydsjsvBWXyxX8hFrF9ZUClomSlnB5KhLqxKuJlqQIBRLsFyuXhg1PlA3+w//RgREOocf0u
4EkUeXZQSJ0/fchoAV6vexKY/Bz98zrmk1Llt0dREmPbBHBiL6V76703DTLXy+rIlQyc47qvheqL
QBmdftQcbCjkMOlXYZgemSbf3BbltJGqyIQ6rZ+JckkhpoI79IyOMWpzsyEfGaT6CJp0oWoj/ptS
mf+PBW0z9m2q0aeEPJzp+ETZ4Zd8trLFV0BcCGw+JCeBzZsLMvvg6cvZizI+ouMOoZMCj1PBcMbw
fsAJ2DoFFunI9QvdPCR2Qx4TqV6KEmyTk9KDduUMvoe2zRmAI2BMFpLa9alKwYMu0q3JsRoKFKhT
nA5UIkSclMYoJ/QWLk1oztD/+3HOxR3MNUoT54oBk+PfkHKY95hC6BYQtaUMeYwflWjqAFUlEFBJ
EYz1srWjllBGsHCVkU9vkWyUVBX760sn+xamtf/st8tzM4ZHCWf9Ii8BMbiy4AOHKNaDPX6iT0Zm
WpUhD7pCEdW8vre5yLmXecHEbVeSnZI/28Fwr8IkWEQzeDgBpXZO/fsykkqMKVH5tWt2csEMWeQY
Ou1s9WjrhvvkwgG5JBbq5rYtl+pg/GUjgor5KBBfKdADoQ6LQUTLRLR/hyTm7oIcbBRuV8rn/tu3
n0bymLvX7VDvOmi+3geJIl+c0cEDteS9fveT8SCtvziQ2iSPgHZJTJsEPnSFjJp95Q5FkMJca/Ot
gFwQqUpJPlTHu0gmPedGZgz/R5ujHMkY0HYdBzfkjhhW8MyulaalPp+NrPxo8Udz7R3sREgQXSU2
oxMpMG5ghjDTWOkY5d6gJ+bngTUAep3bpFsf9sOgWJCoaG5d1s3NVRG7ihfOcz4OM4AsX2afHCdH
gZXKaxouMLDSnrFs6za1mr4InBFrC1LgPCD+VCt6cK5XDNi/9rJHesKr5pD6dnMa5zKL/EkQGdLD
/sUm5II/IBUi02w6Gpweh057Yk0SM1fWdfCV7Aqs0mjoPBEcPjmGmy7+u9d+C4wrB3v96J8L/S74
8ZwQVPQvsYVdpyyw654QUhSEpYt9HcTemfXnXECdzCReeFT/q6/HdI4NnQJeSqwDOrjXWk8Vo6FP
p+hStuVFgrv+7ZoBgL+qyxfadftulbpr9FoGRs5wbqLI1WmxkIV1iIAmEE/5Q/u7zLibGhbkGo3t
bhYj2o1PJ17xSxJ3JqKPaWcBVvknwj+P4GdfzDmwyuc9P31n0iPxENdemf0w2X+MhnhBgiZXN5Dw
tLM1/OCte5jm6d+3WZ0+6CH75DWItwn7XO/6XuVmj0MZvYoiwHASK1ULCEAp01cEtMth01y6W8Zv
s8/n5DtBSGfI9Wdvej2uRPRzvuyH8mc/bTFMkwExz5Wbm7ezUDwCBRUfLZyMaZbgFqqgET4g4/iz
zRjtP1woiEfQS0Bs7MLnoC7z9+S+exhstqHca0oB1x4pYoHN8Ccz0heqUwfSrnn3q3hoQFnCxMSV
mGmkZdQ/1iQf74GVyD2IKtaUYICPKqGACMdo+aNJ/dovo9MvCCykCrGmt99Dr6gR8y0xaZG2Vc8h
kVgQggYc4fCVa0ABAYiR2KIAQHNKWQm5O1UAdI0d4Vxp4K6bjV2wr1MilBn6JkpJDNzWr8gQCzor
zxCbjhBr+r8jnPUCr2ZLli9Nrn+Ok9NMis3lIW2wNQQs2NoVqT8kxwE3nWjDUGqaSAAh1J9jmvGE
C6E8WWCgoZLSlUWSTe2WCcddk5u+QkRfAmSch64wTcrFGXkhsbHnKH5sorvt8Q9TYJMjlWQRdt7T
CYW+JxI385uMkMibyrz4EZBSmSi1yPioW5Gw00qd7Hy8tGJ3tO6sIqUD0T+aQiFcmer8AmQoHKNF
h3IQkmUUdd0fWrBkjjkJQfvztDV5VOBsOB3bjI5j9RbUXzRhNhVQpG9ww14Bl+nrUUtmt3ur/5Ei
zZ500NetXRnGLyeB7ZlmeYuerkjlv0PpVPxlgC7fP2amfwEas6xtk4WrTST2zQP8Fd/WTmCshX6G
geLp8TNj+RZ9ZC6eLXQOwbcsq1zi5Z47kSXyPFJKBclzBdWgfz14e9/foaiOpdqW2qljrqoh8Diy
Su6nT4HynbEPLswM2n0/gWV8OlyoNGZAvuRSmENBC6sFJjP3osLsZMShtKKmc42+HAtQI2N9mTMX
s6NNchsaKC26ID/D7F24y/xgUrE4oWJ4pM8UJlhUwjOXT7aNZ1wE2bU+OklrRR53LSc85OzEJ6Px
8QI5nq0ikx75/IrS3je0kjPIHVd8TDo324krCOTS7XfAZTTh4G0OYK/UEZ1QMYRtCCuuvjX752ml
8erAheO4VZGLxrIZVUG4QqKvcSP8olJJWR8AGmmqRw19TVnbye1Gh6TweLYFAFd8sSQp0FPZDhnY
X2+mgCtxpvqoSBuFhGy9CQAxhsb+lF0kC7z+sTwjOMXu3Ee3vUoI9HxVWnfq0Sdd3pns/uzHF1Od
S01p4TLDsFY1CF0cY/l9uAkYgEa9m1DAfGCwGdmZiZDl2WG1d+JitHkHfTSIuXCsNIsIsTN7h6Po
etYra4Dw2fZxBHZuaI6+5SbG2xcmQ1jm8P1nQIewitwAjzpZ9bPa6n3Llhq5ORRrn2ZrebLK9d10
NeDtRkwKG7mp/g9Zn+KKPdQ1PJtXo2EbPFG5mIgMK8jZeWw1XZXVhkjFAMeDxan3AXUm1exhtPQ7
l4b07I6MGToBNEwC9KeCdwnB86Wd+zrMGzr+ntRkM00/NqxjAeVx9n11Esh9B1cSoOeCt9fklq54
jFJURkrBfZlRVkbMdn/mpJTr6ecYmY1u+ila5Y+7m4zdkagDTrBm+CatTvKN6ffZXsSoMOk0e3V9
mhQdnPMtcaNIecjC/rBnLXYhiqZHK2TJx7wXUAZXMS148BxPMpNqvEHzhVygnhsegZhZ73+oaalJ
uSXp36z/VtvOknSWpqWAgkfkaY+tWmRIfiw+RSFCFkztSmL22GsH+9MVUNn3mBwgjZvF4hIXj8zo
llQtd7E+6BUR+VWa9JPqkSRdnRkRCZmXXah3+rLldEpGoBLFhTFybMd5323HQIRhw4vwoeodhuht
TnbvDlO6XnNVeUCQwOUEFhDMzRDRphG1rY0R2n3w2fsSgHYV2z8UAp7hITp7alsa1SmRCpMQrN2u
yth4sAbaZ2SMyDbZ9GUjSQGoJt023apaK9grzKQEJuftq2eGqi14H9/Y8BLq4h81yp5zgm9uuIn5
r17rFzIM4SOtE2fWnqzqf9/54J+t1TPefKLxEiMjQc7o5Y6wA+kfK5i+KkagAb/d1ViUEjCiiRGK
jxY8ykmjmOH2793/ngD+xIXYV2JbPwotOrm/08lm7dchrDKezJ2YTjMeBPLnulefwCXtQXGUImok
DqK6JNkLO84LCOOCvw2k0JU7vYdnZi6mcxEUFEUy6Ql4n+omZr6opvO09hBiQaylgEHEST+GhQeJ
3M9GGRRWlT9ciaTh+8ovDiAsXazLH4wdn0AhVmS/k4gchQrANL4fATXRHUUvsK5i0uKkl4ECENSt
Ks+gEAr02353PJzIvWjeOSqaHbRb8y16jH5IABe3fiaDZdZcBxMd42wSyDj2DOhrBCSCPz7nA4Rh
Yw8OaZvUJKzfOKObKBsr64knpFLvXtUACGPZF4kcgPiYP0Hk1MvEBUS4cvmqzE6+4cemqaerU5CR
Jyr5ex4FaFN09Y1fRmqUVqPdwaOcwtCfizIwbFbDH+9cAZ6G0n28bvR/IB1zEIJqNAtf5WjKiZwG
/3jdDvYJtHNbpnxlcT/G4XzktL7sGR/5vOWK1sLP5CWC5Y4/MWygfLfYZTXVva+f+hSGkynxkEIH
QJFlG1GvabKcogjtAegBFhpF3GibXgoNSPbY8BYPHOidVlrv2yXFf+ybYCv8S4JqwlkFKpXQB0ZK
GHdagqANaRqnr82MGn1rd5qXfeA60DD5botts15NLrgUvgyK3LpPdir5qbt+Iwyn3UYlgdroKe59
jhO5xPomYLk36W/3Qb4aw6eb7xfce/X+ZZsu7lDtM3q6TgBkNzVGBysQqNBVfS9fYdkJPMLk0bwG
mnWJ5JhrjDOpgILmIt8YalxojGD8LwfZYu8Ry+ymDb2OAfCXwRcAxtVNZDqwWE+3hK4psUeat4m6
XMXvURoEy63CxsFREsPCRRLzbImAmWEzS7EixJPDAvLGs+cD/9Qk+xPjF8HeJIJ6AASS7ZSE4WyD
FdkW4XObo08fDvYYnkcqWayu+q/cZi2X442gf/WJPnHKWLihLDYo3UMF1HE2hdrlGzjrE+vPTogV
QRgqQtTq6AjdyS50dMH8HG+yE6shteyKKuAbJ0MhJ9tiSTS1Mxwun8RHoXm/s8v9H0u4lF+5gpDl
8sD0GSUYfK0swV1qHnj+9NiYez1TJ3nJlo2eqiPZLfoXxtZytdjeWbwm3PdcmMrWGzQ2qwt/IcEw
3mNiLSqhCEniTeaLkYcJ1JVm865P4nIerFAymy2Q8oPOECiktsFu3sphLNJ/zO5Ndsfz5mJOhpSi
AR/TuPC8GIjHSsaN3Bi2ntx6PiBZiDjPwdXS0C/Zfl5C0kmSxlVlG4il5J6IGmGFjHaqIvdnOEQw
ct27hRREczhf+GT8iWdrx8xZi1ZFIKlCFNDTG9Z9WAvpC2IHFkf3qERuo8LZh8QbaP2RqA2AJ09j
hO71kmqMpXvqVkhuH431x418kILo3W7sr02G+xU1+WE2xoz3r73mtoG5FICeoUz0utRK+y4JQ8Ic
nYK5Tj40N3oDENBTI5AE97ZD4ziIJWg4XFlKMxrtRUMIWoJo/ePKjWrOW4qVPYNslUrMv7Dp2n/u
pBrFHj47vNn4LyoI3dfP5RKedx7d/Fanj70Ky24J+aTE+srkC0Z8+o7aBDCyqnYBBcFtPW/HV3u+
g5QSVYJikRu+GCq3zkHJVAXmcaXJ6K06qFRZdl8zfQoMYxJl/y+5srR8iAqh7PcoIZKgXE+W0Jcn
Hxn51n91h2GmTWoXX9RyZzD98N1FFkBnWXGYqQwR9GH29eg94B5MZ2YUYEWscmwjcw90lZDnFiv7
+ksKfxTfY4AGEzrEKUu5aVydXu1hWYLROVi0nYGFc0XDUMBIRhC5k9IKsEcKTtFPnFi1CUrsLNik
xJ3r/VoUzLApAmaobrdiiI/CmDZmnYqxY6WX5M8pQ7kRY3j7y5yv9arH9x5hcrVPSbmqECS6xcNw
pXHFga4xKabX1IB2Zhmq/t8ffFxgiNyLdl3vKtlod5m3mA3fUI8hRKBywF6RcPk7KOHMZ1J7c/NZ
7G4y7UMGzoQ1bYFcWk6CmD+/2wMEY4eBUc9HGBqp7QcSU//fvEyE3g/sMC1nxe+gzbjOAMGq4YyI
13YKeGJc56Ux13O9YsmKTMHnI9iXhOKwhhxJxAzAeGuPTpFMGhKgfvwdjB0paxgbfRemNCingWvl
bCeqH5vpU1miyDvBy+lPNJAgyYVxMpF8SikuYxIxF4GDrw3RwDjJELkRERVELPHTRTlx8lqCus8T
vmT/TA8jddaMjTqFbEAph7NhtKd0C4V4fztGS5e/306/O8oqGC84+xrD/d/eJO6/R5APkEI42KqB
BO4lbRn+EclC1Pl4sfILsCyVj3zfdYbTeQr/J+A7DM52bNKeYUB4vx5ybeH8hTpVgNL2oir+1PnB
XayNfhiZc+7YzLzniMITrA9zm0+q+qLwFoOhHm4724bwk9j2nnHxU9X6iiE5rZvtaog/WacxvtxW
2XY8oAorhsPGmENeHXXlNcEDMsci45TCUlXlJJO9XvzQvpzmsO6o2hTl4JPDGkAxfKSJEf016560
TF99M9cyWi5NSBOSlC8R+JRc3BeFEyoxh5K2Pl800S0i2THozBUSj6dv5UcZNlpMoqclG14rvN+u
75/9DlnszwC1RWYUvLKubG74CgjPKCxDyxsQC2Yrse/CWptaaAwKMLjlcO5A3Hv+ohW8kfByOexI
HMAGKT9CrsqpB+CM2//5D3Kepy6/U78qNHX7W1Z9eiGxQxEIdSLBvW5j9RYUjo0e61zpO0WqUpP7
+hk2+9Pn5SnN2740mqvF51qK3OVyRnZm8Cj8Cy/x2Lo8cP56Mjv7SGPPi0ZOuzabzFLyzYUkbe2R
i/nvHUmpivlZ5x7CJHiLfEC8TzAjsSrBtC/Z6tAYPgkjLTO4lCVoebNtEPKyflYJjcgg+RJiIQ2n
3qKhM7/0nWKFQvxEJLJtcYvXe2N+5mthspbf3w1zgx1O2ZfXnLo+bAydOaoMsEaJQFsXZCeL79rK
xVRXrG5wysg6jFPJrO4bUA4ny6I42JjDveazcAzcfIG5HI/M7nqCUYUqF92/L2yrO/o3jKohiArc
vm7A85OjzMi8jugy0GFJnociVQBNs63OELadgo/GQ/FjUviGc+XGFGZs/nn2qKE0SoZtNmm+rGG6
3map+79HONAsBWauc2O5eByeQPphmXFdl+UEhBNXLOB17L41KsIXGRjmhzrlXB/VJExGLgzlE0No
n97pAPjIwRpDHN2co+SzcVodcyHCU51SGRVmS4elktgxZEiYKSuaQugJ9qscLlg0UBCIJvYgshzd
xXVRnJ7pTvJ6D3aQueaikDfQcciyz/+9fb5I+MDReWV0MliajprRcJ5Ho3BCd2H63ykpyWKX+OiW
Bsm5cIO5W+fKptIGevfCkQuqJHL2GnXDJf2bmyLaS3UpcLGMSAR7cyxVsErKf/CdmhgSa8E7l6PM
Fy9pl6FAKTKp5oaSKtkfPWN5zCfwo/7DJ/NjBXYumXth4QxwvjSo8s/vt45MQCkjWIglJkS/LSIH
fOsGAsGg2z+ZiQ5xN9bFplrurpBd+47jpFtSGAGR9PncFH+A07sOHqZ7bw1kzSf0cOxwdvJaCaLk
LHgQiyh4pFI18thIE5lh5lToWbBaECGmNTlYkXBMhB90QF0VpNfdAnU/gf7Wr6bEqMcQTPIhY6h0
l9YZ1O+yLhAiC0rmWWxsSo0BiEOvzLlvIsD9ntUI4XCPolMIHkUzTtqqAROURrIBRlwEZBKYBb+j
RsIdRu7VK/FbGa98aZ1+3PgCWwoIL35g4dw1GzYJcCYXtnp5L4FR1P9DtAtYAB3Hn0whBxeZGpB0
r06xFRsgkenlp6Ldq65AygJA1fYKvE7+JiJ+AvdBWwPPbb9if4K3+QAjFtDf2pCjF/VUJnU4WqeA
lQ3ZEWWwWWNq4fZHFycWxYtt9WtJqAMYyfYdf0y6xYOUg7gN4xRCMayhcQYNG9JY4iY1suTM60Sp
1gL1QS9I/B9WIu420A+09JZ+n7arvYBnLd7KDD5SzK4ff/hCLkBdEargxqrRfFDBI8KROqB5oxcW
Wg14sM4R0Pkj3uB24nMIArHnsqFl4/QaBJ7DYnbRfDhx6VMGPNq/b6fFkZUU0Cs6gZDVNBLDHsHi
qaFZ181k8xR3ai/i7X27fo2CEY0ikS2YPaJoh28nuPEnCt1AIav7vvf7kPw6R6pEH6UrCxE99xJ3
40idmg38cLM6PfEqIOfqgj7bRQInX/RoDehWj8dG8aRbZna8PiDQ75dfrl/MILD2ysy44rUddtRW
/kHC0GToqSzx0q67CIWtdmTKzjPHT+krBhE91PL95oljDSaJQX+VrZZbs84DP5b+vS0NdaFOtViw
6HKZWU3kWajcbRAvAjuNZWDFAV5yxHGmZU0r7lmF2+e7YSQNiFME6/sFAUdcAkz2juuUR488jNQ1
z05vjNnWv4scl+ud4JoLxfMv0c7smekmo1kE0pNqh1rUKolneSzUk0PcY/BpLx9vo5bZglAHVKLv
nbP/OUs86t7h1E2TTDEkZ9eEmajGsr+bjo7FWetlAMXZEf+qv/jb6wxXKZcUeU6c3XahZMKT/PAK
9425m9ccAj2Y1uPXB3UUmhRXCO1lPRRu8UGpsb68aTAcSOJ0cCmlvrwy+Wf7Vsuf2LMD9HtmraNX
OqLIrn69GKn7mzBMh9lQZye1gmsFEtbw6fuRJtylEevHZeGyfBQRHp0/GzK/qoTKH1dIkntKOZ6k
Q3ZcJ38RtgftZa6a2KAYphH1U3phsaiJ5dDq8s8HmQDWoH8mVEk+MvXmxItLOcRy4Y6quqhNWr0B
qAQH8IfRC4RXftQTwpTWENEv4Cd/Q9LDt5MjNn4u3L1QCp8TdO5kBdZ8dsiBeMUeQZ503iOLOWCq
rHDkL5MjFxGWzMsmhTRkEqLhvQzJW+E8qnyIR5xuQ9fuaI+/Ur1ERa2MWcfvfnSmMAZvLoJXQ2TA
9H2N5qJM5j3F1JelpIp5+c3ztt2+AJ/X/ZSYWE72YORj/3WWZ9XeYoQgnDDmkLnpwCPLPJFWM0na
R8iC9HLXXUKYTjkm/Zou3aq99UvPqMlgQCUhxjxUyK7d1H/92P2YsqNImh0iv38zTEbD0Kc6naDQ
FINDKX98/n7tLzGGGKor79ncvAOSrcXUYpKdIda0Q/kb7g0CIBctPogphiwMOByiARq2R73sCM+B
gLOTsHqsMW7VMGZXOOnH+mZ+KsmgoM4r4vgEpN3IOk7C7heLymP7/kWcC7X54n03JgmDSaOfQ89K
4G6Psc4E1BitwNDVFg9nixOMfbEu43m0EE3qsU4IP+mm/cjE/sf7kGA3bK3U2ATKPVIlqCaBfzNj
N56bR6Imt/jZCWOtEE1+9gNejOrg9TUh0SxtQHHBqlID3xZenHQ4+gxD6sBzd3ARxsCBvdVK+Lj/
EnZzPZ7qmnhyODBmB2RhoQLNf0ROeHjg0tIGJFXXX5qb7MsPHhBctWUCQFTZP2RNLg5LzJljXCel
xeTWzIZBgzg3VWlrCoVSulHRoIM26W4AXw43YepNbAiFpv3c4iu8yacgXNFV0gx1RFTXQufo8vlW
ua50lDohY66N0L/0Cxmk5kwTA3hqm65DP6I8iD7Y23dLcx71bI9DMG7rJG9vm7EVmDDnA7iACNQJ
QJcPnFgDBKyDOFvcUsnEvpd3yCG8WxPsJqa4QUOpP5+fZFg71+gMWvOVs/tTkH9BoVAuw9MBmrjB
p8UMc3ogqVK1iDDHb/V5aTUhpHdWGXjRoFlDKYv1sM4m6JbfoWIjZl9pnJU3KBsn8l7CYnD6QNeS
jPvSLIgK3NDoLRNYPkp39xx5yhFbVzBGCsh7S4lKLcuIdLy7F9m0gxA/n5d3VOrFxDxuCu0FxnD5
x/iCljfSyUTP6emIOCqFKJ8lLZ53tZwriTZ7usBDF8wFnFiaZaTDFTWqAX71YIzGxXeqehaVGtWf
KOcR2pjHoqgpRg6vQ2ilg2FCjLLB4oOxQg5ODwZqj1w4sjNbMdKY4V9SQGD/2RkHgA3MxUua7ntT
7nCYPnSfD+r3STlaDEt4i68+ZOc85OPtNQ8AzVR9DRSJ/FIsmlJdSa+grfpeJy/51BNgIhZcb49q
XX8u/dVuC2bPc7woNLavAj2j64XKmm0jmlTzfdE9tnWYd2CTwcErktz1Nf+8bPztG9wyTMg/7Nca
ch3SOPbWhxOIgz+Oc3+AMZHNLE1+2yuRvDfUPvksCTpKE/ztUXysM1Qk5zmXyX9XLzGe9UoT85XR
yvEsXzmbSmpErh1Mh2DtEfRyns0dVnp0y0kiWouSiF7WDuPPFwf8xjh3Kghn4aluh0afSAFsSTis
+VnaOQviZPbXkzKn1Lh6GNGXAmvJjO/deO37kiMM6qWdvkl2EkHBRfzBs+msIJjIZd1eUGbJyOMM
OKpsRJRcWvE5Vbt5PDO8z6C6NRvS1kATwa+QIxV1uBHl8X0865+gntqlvrLfgBM1FsGBsohp1VjY
5z9O+RXmIC99aaNY37hHcvw7qf1F0tVzYGo3M5gwc6CH71q13x5puyKDvaSZXdGHSs82/MzA70yg
/q1peHN/7SxSxnwstCXUx46+1yeXSnysFIjYrLP089UkpKxpnG7eaN6BO0NMeBEO4vNC/j9j0FDa
FKrJ+vEMzKeckSqW63w134CGt9QQIWS7SEfLnb2R3aC19ELe0O6+6lVn60GDnuSYqRz/OMNhGJPF
N7HSElxhclXgBMQkZaZhHe/Gr6q7s8OmafThPhjEpcG7jysJ8yrgrTrALlxfzyRvoNgi9dRa7TmH
covVxu2+5lx1W2S/3RkVEwnJe/FWmHHF5B4q0LWyfwN9v9JK1eWOH1sqw/5GqERn/7HisS94Mxwl
vy9KeXdi5inMKpMEalrS8p8V+FolDV4XyRfqvltToW4Zb/t0W0LFJBqsVlUBG682pBl9RP+6x+M5
GdJLkezEAp3e47h7yd4OTPW2h9imbti0U5pYsnfiq1QS3xxOAPZ8O/gHu+B35IiY/m137a1NdP88
YxQGuG23cYDPPElEHmOnSHfkgamNzqDEKl2yvTzyFJx09iJmfErI2G1t4imXjClVlvrE38OXLRFP
caXc29ndAn7r2HiiunazI4GHZjq4y7aNE8mPa+1jq9zHN6H0jS4k4KxRkC5+DmR4/yZuNjcqD5ry
zRV/BxfBPwLM88lHqE29PF1N9f1iHqGKJK7WW07dKsVtIsVkUToFOUS34u/p/eAd8DBHWdX77CDe
R5IEl1zxiqNQREvGof8MxnXBqaaIQnk7v5cf49/Fu3TS37CTb8goERbXrkojoCLzAB7vqniwh5JG
qyiAk6ULdugS3p5bDtvOa4dSPPkJhUTyvB2Whjl9gixigDLfkY0swHd4KCqj50PCe/q6d8+g1CIt
Hs3Galal+b6WCKlVLl8Cos4owESg1NpPOdBl482PBq9x3kDDUGk0v3IEqgYw/DpCxfZHJjZ1+qV3
vBBsnu+cyExqxRVLqp7QPVdb0vO77AfZxsuXyUfCfQ3pdgs/vWaxg5+OvYcyDn3HvNHzb2izh2+c
YLilVJA/JynNzmZlwQLWuCziNwgeaeVTNlmT0I169ZgaHydFUxefu3l5yO3GLyAk9K/9Br43lI4f
YT9vMi0s1LQBbeYVLTdTIyhXEMMXWlO0dNDY9S5KmK5H+64hJd0Ep1lhx9VwC0FP+J4XPlEo2DD7
Gd8esBzvZnL3hCV3HjqqEBnJLycIyl7/vnkboezMm7XMSrVW0JWf/wJshJEfpxjwUNUUL5VgI4yj
97HQlzJk66ap9REWZRz235yB7SWUEjX3/WVEwdj5FhuyX9zmIHwI/FnhiCM/b2wAU6UvNw8BXeMG
KvZEiXiPiuiYGgRJifN1rsV1xi4jtyYqxjGN5qAMl1uz7UOP8yONYX2Ns4sK6iVKbA0r8t4aIQSf
yjDw3esGkOiw/LhR2bd41SB8O27VlJ4gfedn8FDI6NNYjZ9zFBdUnbRlFeFF0AntcZpq6i5EXb3Z
DNEbGFL03Nk5ui7BuDLAwqObh2eMuf1aiJRyLRF/oc3I5niRIzd6kiW6Rwp/oZ3gjxVaT7uURe8A
kWY6zCkPPSyHCb74j8xc8VHxnYRzXdTlyefNjDDhFZByajukkOHeKMvTfSkk0Vw0gBUfPNka6j2B
TYh5v1IytFVFZ2+js77enVIHOwWXm0jaILmRIEr4Z2AG8Nc1sQvhRLGmDLcxSDIDYgEsg8CC4tIn
dtUsCv/vBM3UsWJeEXP/KPm7Zx2V8A8r62+YqHPuEReGUnscVtJ4vOgKLrpUladfqzpAPZg/+KZl
e2rl7W7Iyb4ZwSEsmCzSX8MvYN0KCX7fseY0iBSg0B5PPPvcXJPkpK7qDDSSZbToN3yrn912H093
Y2ecCUVJ+qcERVqQmA+3rUQDYGe3EYLb/lIKUGF+Y1F3nFSkmba8BVPC5Z4OawWBLJDglg7BeOKM
/s2V4JdGq38GaBBCCyFLeO0EGyjVTK8d1rXKr5cpgzA+E/xF9+Vzz9qx7xrBRRSbrtVixxHOgrGW
HTrMaNT0mKgsrg4+Vs5WrYvfgsFrD1D+nftN47G9MEUk/luijkcUN5r91xiSgPqDaLl6HDsBYw5K
3s9WEvDiiPrHA24HAtMdjQj7oXHvQqw15gKy1VL2rBzNVpACG4FWh8Kj22FV0DpKi/N0wfm+aVvI
d7xXi9kNKTox+c6b4EN3mXYKxcQ7goD2ndHrGvEEHTrlByNpN+9NuVsNBhEAC9sqIN8Dp4b2QwWM
uv0s5fjFIYHRkjWBVdR7FUdFXw4+HGLnYf3Gxtbch6DR67UhoTJ0noX4TQm+1dAKXcdfpLNnIbRE
/JM+TmkUlUyqeWZPPIIOdauq2wE4IEZe8QQYg+jbz5hVfK8tAhDMDAVces3fwbUbbBzyieiBRDI8
FsL0BJ5rv9VVTxkBQfqDvKYZHTh//4TP07HB+HHTbHSZmZSa5jLsr/AUQcJfXUq63VZK17SQhWWS
oOUn1FqTeJ+hjagj2B2mymwcBsSwPnzASlNM/YZxstLJtxhZjjrwM1ja/2mFEOfLgRJcwQAgtyFI
F6K0dldXuw9rs88/xOkCQ4kaLPEWAQfa77t/9rYt9bCdQzNzSufSeQ7L3jXE3w2O7SD+WUFdYwra
IZXes0iOG5XA8s93lb6AJYTg1hFZJ9xCCJ2EzRAbsmVBIpSuk5hOCMPQEOXGTkle6+tTXBep991y
VYan1IsjaSAvDqZkV+oTGPf3IP3dC9x4uBzQ0B9FUHQRXgnBq0GbCwkczaMgckuBjoSbvmOKv256
wU0NFwTgMNiwX1+9nkrNRJA8TtG7RPSalv/GxiBBhRRqLMRT24ajjEtnzWmK+werQjYIGRqw6eFk
VXATF82uDBnLFuzT2C3dmJA1alA7KDi7WOPas7/ChVhP0K2Rui/1tJxEiZ+jvbr3ZSEU44UoR2dZ
dzxir5JnU8k26I6CJH8/FprDBtBcUZWDf3VrQ2d4mGhrAX/zulDz2QHwdVHHRrzD2880Ikh/tKyb
esHrZp/VdoNFf3+lgdYO+/tXUYF4ZXJe/Pxt0eWzMi41OAWEkivPpt6dE7UcbkuEigRh7RPrwoCB
k1HxEa6Zhbj1vZaUEsb7Wl3AJbgjAu5V1Tap7QMoUPQaOkAHQ2lYGb1hNF4o1Isvnhz0dvT6YHkx
0Ql/BDJrkEJo6lSnplyo3GzHvmWgQrFYvdEapMV/6phI8ZvNqCD6S4pOYgxGBvc51C7EIviSO/Tb
MgzTXrhm8Nkowkehmos1dHBPm+5j7FL1iBuymAgNx9tEZsG7qY9lmH+G1N0+HiSPOmEEwq40mTqE
CFfmAc1g5hEH9wXdMG8NPBBbGs3FHI/yciC4VX/2UAFr7LLdw3GyJxgVTQxT2H4k1Zy3QhCv7LKh
dwuRJNFkWO/77te+Tl8lkaNXRkMN8b2lK1GtmMUeq2H4912d5vADYEaSWcxfycGLUpE8y59nsn0w
RQIpW/M691T3YC5rB5IdnUWfxFltHOccyesYBfeVv9VXw7LxTNfrfs5WlvuCjHll47zbijwkYJwW
wQsBj+Lra//Wk/kqxVpXPyKa1CymNDckwOcfozFWD1o5vs60S3W0mIeJiMyNt/LKHO/uPYXmkJiA
o1XVu43+iHVugKtoHwbclDm/rGpcuFHPY96nOvVxAyCfRD+woZ+a7afaWetGKsR0y+OtBBtWme9Y
oNfU+gieLsip+L41dnSOnWPlaf40nK4IJ0agFsg68H5MAptCX0Ax84Brqf9ozEiWDtF/Vpu0Z+vH
dV95gj2QhjtzbKz70z4k/B8nt4xuveworsEJqMRRopMu6i9SsztvCZCsc/dzwOR4Q0fbRWeF6cUp
mdeJvIpKCUSzquLuB4z+aOZOMlYU5jhaXf04uuDjgf5b71CzDpG4mSYpFCpzJ2VXj6sLpDZehl7K
zLTOK1vdLYhkrxys9Iv9zC2eNZlN8EW9DmXGbZBahfe5x8DF3FmQH7v5C/iba4UvqoRwCGChTn2O
y7fQ8PZEI5BTTs4Q8oFGEJnYhwR5VFxEKLoD44X256dFgmWe+CmrqVEsoP7VTRpzzpXcDxu/xO7g
D4b3MAC2QxXTp/AAjZ/DxFy0i2cuiANijYGyYG8tMyV3j868+oGo0hhNtHX3gqckz4tanLc8ul5f
BbkeqAkY8CMdd1Mhx7+ClijJPYaNBXei4lyEdCN3BxXIwI+sx/+bYkBe3TUDVHOguCMXdzxiPZiQ
3dvB7IrevlKCT4Ph2r9G74UIjOv1tJm/drGqd1VKAXHP9yUUoqWtwLLR5NQxfg3g/f8ZmyXia4LU
bcgu0pQc9yUx+lGkYaWUX4itzceRUtpJX6wznp26WFhMcynI9cD2Ncq+8K4zqKbG9BQ2r4zSY8AN
U/Qmi0PzIuWKs2fBvE5VWeF5sqnTfNak1yZ/nA++eyFu9g1Jf6gpUN8lLNL4H4TLACn43NGu1SuP
aPX+7kMHFESr4aDX72lJvp6KqYlv+7/2IYVkRK4X4vQqNc0qEnIYkXy3veJQGNFDghbm+y1/t8aD
V4oiCubF3PY0nVwYtJ11ppyshVrwmrgw3LPsxN6di7aFIiIUhWe/J7Py1qxeuI0CZUeskgNAxyyK
yP2WmQbLynd7H4bLjyi8XtvsVHhoUtZhgGa62tepvXVHeOPSIiOKM5OuWtrlGjlZz+CITsnrJ34u
4CkQpR8PvKhCa0zlMdb6DPFDI7NVqiNCpSsHjxBGZ68NrdD6iJoX1svzcDgQtvZsEbwFpNjiNS16
MTaiQakgmmOa8GiO1dtJYh5+krU2nXhMEv54CaBH9tdDnO6RF9E8Dgt+3LCnDFOrr5iW/0fWfe5l
Z5emws3f7Zq+2qpsp5a2jvALwpEKHQF/J6CWn6R9DoBmVS+qh6GNDobosPG+MNk2lM7n1425/pot
csyC68cTe+guS+/t8piWuxuTLRHVyLHnsgpY6wg5gxOpgLriOku5ZukfRxR4C20xk6Gk/vSNuz27
ooWw4uKILt7fKlwffZm0xGSdo3T7xo/+xAkMTkCqvS+4EOJcQgnSnZ0EvOAgKTXZ9UqLlYeFI6Mm
2SR86rc8R7Y9czy1HkqrNhg04J6SMMmavV324/CPiPEa7hGPsOL7P0fqBSPYyOHEdbSlgDPKS3oA
nEnvedc9RCCsNdqXJBdeLYR2a8ER2DqaoLFABcfVP/h8FbKCPKh6el5C2+ySI+JM41+bpo6hw9CQ
XcjsIyhZ/lc5Ah7eFCDH96VMsjy+eSPQu6bvk9Bpc2vN69EVWr43n0TZkOHg1QZ3pi0k25t/kEPX
Wag8tizZUhgfYZPBCrewXLgq3HRiDrXhgfF3hbGfaQq+gcteI5YPwXOCL8SSJD1aazPm1plHyMwQ
IRY096vAv5cHyhMBoQTMLecSQ3ZaeoNGLx589R18Ld30UJIL6A/XXglKXCfgPg/7jJ/R/FZbOoys
6GjiF+V72J2UczlfdWMAaDPdK3o2GdSrWocg/KuOD2wzL94zMthP5gh3BKfryu01eENmLu8oZEwE
SlWhTXNVHKlZZ7siNevlJwy9rEr8mKa+xJWi+VXpPNJhDmiXuv/NUKsgIWREqdjPWqocY6hrrUBB
DyH9KcXhwxSaEcggbwamMo/l2MJjlFJL50ndJFqgi3h9/Jk1F7IjkzpQH7j5p6O1Y2Ms1xRXq39W
HV26g0B4VQgUErhG+k663G0LiJaGTkKIzK66s/Nat5psf8rJEP7wDlKkK3MwTeBMUqJRkUaoW9YX
0rE2QDdZvuHEaTuB/NilmJpT035POiMv09n4RlN+MbLvzO/D7y6GPLH1d7ONS72qHOF2e/or9DVn
wFVR0misBAMxTcOJH27YD+JWgPdhIn9hR2Pl0weTbsUSa6deHIyrFMjl/5Ot1zBQqu17EmaGtSP0
tD6KYzKQxlfCdjmGH4WBuA12AsKi8t1rXeDWh+8NAjwwreqO9XHKzc4elilaKYqqJXuCGa9VRfxD
0eeoN+781e4zxYyUXtGGh2jFJ9hEBHb2IBIwuSIC63q/CQNN7jJ611/7tjsN5ksIPmkcgMXjB2XO
r0xBjzHECdqr8rsPhLCYnKGJGBYdyFfT1OPimcsxiSsCqakiPr3e+JsXBtyYFiGtI/fxru8mRe5M
Zuvk6ZLNNzGkS87YOpO9og2bAt8QdCBw8XP7hCwC+8viRlT6ZLV/yapqMC9uk3CRh8bo0ecbbmat
z5okdqUG9S9EfAKqIUUYvyiGO3wN/dfzqN3YgjVfEd1kMtn+Js8TuORUfEotMSuUHpfKwH1IFfWd
PUcW94fIKR2FdinT+F5OuNdPKRiIgrLrpa0xRdQndzhTJKjhnLPIV3rL8kjtdSYKI3p2uYWs6ILb
joG+JxuuAhLv1urf3uNi7kzfWcnAN4sS4oGEsEH/lVUtYkzUaRyNic85d4e/vopl508St9qhSJEQ
xkcaK/k+BSNqwkb2w5pK4l7LUlJg6ZDp33jKKqDiP8ZSLE+cSPGfUPj/M6apc4ExfKqqZdvvcS7S
g78VnS/Ho0Nar18qjgIGV1LB894AXS53n4ccWwmCpdUlVAPgHpqh0JoaHCIzHYoSeMIyve9n9iJJ
v9ax1h1hXIGkNUeKwP4O/otKkpq+SuLOxjWR4ttYMVD5NcWJZsvN1pwBzspE2hFUxXyOL+GN2Mm/
4zxv9VhxtW1w1bmIyBan9aSpYDZDT2Y6oGCE4nRJZAU9eEA/vlbT4WWq/pBZw2G3h4a6oTTiwPQ3
O0cVtKMgsrYRBfM9+CgSgHPKevtFrMiB1k2AYQA6g9XLlQmV5KtuajJyIgB8fVCt7dxmRGmmOv6H
vPP4nrI8TnVCflbOXWF4mACrMO5+1PVjBqQo8CrgrrK037rc04rNawVzoWOZB6HcnqN476PTuD0o
ZCp+gJ5CfXbSGLtBs5286hoqlP8VWKsdZipiUtWpkkf/O8nKXDtKCuxVNXafxa28BDldSIwpux9H
YTrNyZVVdrLs9E+uo4LD+VPOfYj4Erjyc0mpwgKS3mAYjJcszZGXPYRzj6b6Fmf8b4KyERuuAwBZ
SBYCYcfOAZeejRSh9YqVifNukWouC0mHQXDuDCcHO2gsi+YgkWo8CELr9zC5YOSDln+NqyTgGLRx
94+z3ZvLVXD/td6/AyNOK8Ve0UZu6wOvp2e804eVHWq4Chnnu8kqENDCQMNZovFartRkpb8k36Px
T31lR/7OVP6WziowtGULylFOJLwrfPAU6c0V5j7IIjk04ROS8Iawog0ha1OgdJ0BELqnfuandoHr
vVdrSdabAq+JvhJodJeQrGiDHZEofDk5IXpiZzt/cT2k+TS/pnvgGy7e0V7rg015LKTkeimQy7d0
++xq5BmmMhGkc/6wamIWg4wIDRqmCwGOJYyxrMZAa0mEWl6MZj6HyCo7snAMkMETZNrUsPvTMN3u
oHU2jsA6di924WTRspAnKCJ+LayxbHW8Mu54wEArbb/bHAQBTkxHd99d5YcfDsiBx69WidBCwEpM
vtudOsS+C99wDqKRcOuZpUZ7zXWvVx4SFRzCY8DqdBuyJFXwQcxEeNk7BCov/BsISH8TnBD1txmP
vk/Mc0Y51vaSz2hvcseipFPutF9lFppzAR0CNJAhf9zkG1HKM2AQ9sLnsP0BMLm3Z/0tTdIIAl4t
zTC3NwVjdzVs+EZLEMQCiHJXkzlVL7w40LLI0EpGR1fFrW6blRwisZMlipP4qHTCjIgkupzI0cKh
bo0PLQ4IwEO4oMgFCB2dKBNTX/ewEXTYX2cL4h750BkCxdzAMQoUdtOQc1x4XfdXfVeuuxb8hQE4
aT4z312jClM1f3inYBa7r011Q3StglwCiuOY1cnYRn1dfkqDJnJNw/yqE7zqalkc0CIanNYLSnBL
W0O3RFjvuJSwem6ieu4Jc6eLhh3auoARtqFRZs1eT5e9DVc+oV0vzEPwYwBeTMcShU0RjnMmboM4
T0n283DtnPwT9TCI2tW96G2oq4ftdtLgJ2M7eNMK5BLGGWqeRN0P9wHumAKYUmN2PJxVbh4+1dIG
8E0GBPIuBuMcokRRgEsV/96Q6nOrXOMrLctHrVNVUAkpMdrz+IkVMkEK7tzyAYqtDmtezpFxZ92R
4ys37us1SM7xvVUrXwWzAJMhENVz3t7JRedp3K2pvYaBF3OS6+UYC8S6XObW5h0mSSk7IETGgg5j
WcGNs/4+Qt11dF/mKlPq16GEh7nKjwjdvbQvr3OXuvM/QPMM42D0ZbcXWwUqyeruuzWO6XdvWEqA
dLbPb6nOVNZaHdbVtl4jTMDdBVVqBZnvQr/qmpIftTv0j3OCaCoh7FopOCABKMUtcHhc+MpOQrp5
81jZRIn2LNY/0opelESyzPDMw5O3qva0jOJXCRA0LoifsxJSQi1GZ/ukBku9jiwreKoEMsYd3zgp
J3iFeBTJIBmVgd5yNrq0q5BioXt9y9UWmqnqsTdailzJ72Ar3U9w0xyInzNrOgZW50rriAACl5w9
W1vI7v+xI4WBeRz1XFQNa9s+KkMXznYwfLsjGO4RbuZh9Lsv0gJ+bnBIaMufFRkd41rCiMUqbQqD
nY3zFcKycMir8FarV4lLK7tLMv0jfiExwRDHn7TCcwuFauHGcDVLd3XH6FtHKdmPPqTdIGA3HRLN
Rn3u1zXdPaNNfuCVgzxj4LYdYPv3ILR2qdRJj5w58eGr6tWiIYkxUjK+qBPMkVZSiE9x/CBcbVjy
wd6SnzBD79slfAqdl8A+u0M5Kd4RXWgO/T6sfLBnsivAgbiStr4KWKjX0Xns+ADEHHxcp9E/FID7
gVRIsvNyG7vm7MskUTjCOL4uEBzBCWDs4Ih7ct4o93aBV07MmnxsIm59HZ+uGGPzN5GxlwObcl/B
2AvUmnpBluc/ltObrmBM0deGHuLL806WVPbadPO1GKa1fWZl9us7NgyRbGfPZsC29/88MXyyWaQz
hxeQ8a63zXPYUax5H28MJ3hXrXMtVxtAaj5PGfD921nXXOPLzL5SWgknr6aIhd1IZdAKN7G20UGn
hwbIVELbuuL8MT3AwSr3+CxUCWrMUdVV0syYkSbsZClWn1h4TQB+uqFoc/FlDj1GZ4EIp+7+aoFQ
6fzeiLm7ka+2rhkMBKf4NR7yZrqrA+7ifGIeBvdOYh6tj4LS+fJtsJw+QBj98yTk4cMpUkk5vZG4
AY4n/L6NEq7jXGREC9N01ALMy7X+EGNKbKjV81ePtCyHjDn0lChn2RfK2mYZPK2aYoReqTIduZBW
O2Wvl1zkjHYkbBodI/Z6kYsMCZd1apPasA3iSxD1fegSs2Z/YFHxWMS/LiiiGFxabOQLvlxI9jwq
MyZsTiNTieYjIGWCMdC7bOsFMVrhHPA/xjOLBC9ty2YZ+ZnpCELPm5WiXChFfe8QrtQ1ghCteCUf
Tq4+/2lB+iOqO7xcRbxeWDmEFbWxLAu7TCoW6DaxkaYzeSE2BB25NY40X4TRDwGxUqFJ8D0WD/u9
HxSg/+ONAw3slVi7EMa4xNqcG4jFKzWc/y45I1CJ9Wg/IOFHBruhZOx/qFb4heBSMjC40JGFEyqo
KJl/coYBd1mf3ecGzdwKS//5VirzP1qvtTmmDDfCfbeDmQ9WkbaR6JDZRGoaNZdJvJTuufro2udE
8wr0/8ZzSN2hQdW+gZThyizP9xPt5KFARjdsOJx5IqljU7B6ZCnKPqil8TB43tns+jK2GyoHxHIX
XY1116tOH818gYfrnRUAOibSgv1DwuOB3E6Oq2tealf7zY3vHEjYhHGHT6QiZk/BMd+J3wnisVm4
GDq0DPIMB4Q9/RG4k5rbqAuIY2hQKcUqqEXFOroZUBA0EuA4/JUh/ygrgWQPiv8iXh/I3KWF4pK7
Alq5VUJjCse2b63F0WivD7EPbnT/x2PSyOtTy9kkxEeAyIsl7YvxaZDJJSwW0EFuCedO5rJ8X6rU
7blbIRW6X/2LuORzUvmsKbkgd/h33fjOC/LP/Oo8LDG+7qxQSN5Ng2ZkD6f+LLjYxpPrfgdLN7kL
ej4EYEYbmei8PNAFdBE0wHN1bVL3Zb4q20Z4MxFbGTFO4+mZ4pBsBlaJIJVfL2YUp8OGursYF5cc
QUhRQVibKHOs6K8cdTI9D22DiJhokaXcuomF+2mmB/iLcU5tqKa9on8yd810qVjow68Q5Ov+hZv4
d/aFZ9+BOHTrl8OBvIjQIa17N6WSkG8OCjthMWC0iCMDc6gGDOV5sqPs3qDjpS+NtwSENHLc/lZ/
6+M7MwnFyI6qjVK7ddlAMGI6vmoBeJweJ++iYIiAf52osRhjId5rT4E+sWbRNi7C2C4RxmSYdpnI
2XFexzPNuEgMxHyaSKPP5Mkjenn0pAQgPv6f/MbEnHamkqIXRZuZNaU0oSl6Ndxwaeb/W0HlN0Sh
ibiqhxsBOeNZyFVkrN8/7c94y4vg8ava/DoIRRizRO1HI13qnrGO0ou0tjOSWon8py5M8gwxNwb5
Llx7XAk5kPyPKBIeYCEiDAWdz00BAhhovrI7QtVppORrX6l/dOqcwlTCBvAwsHcK4tvuLYMpzSzW
lgYoLF2OsN/EgJ3fgvQ7M5JGvakvF+2YJqyw3+DwGMMHFeatdVcwHdnKRVWjWhgGib0AS39/Mrzg
qJrPA1WlsoW/T5aDcq35EalrokPTfZYtv/fgBr56raF05ZF+oTCeiAb0l0klBHxt1zYrMu7QAyUT
Ks6jDBZ0atqa8k2vNSUy3ufWpwA8kQJpLTsirNnS44hql6FlM4c2sG/g7CAPohCZivZb45vy5yDD
LZIgS892PM2y09LfsfkH+XlsgIQ/jrfTd7qbXr+761YsCFy1oSMsgRCQCaBCR2ig0Tb4w659TZ4C
KLRdIohDGnx1PyL52p/t4gupGqCxJvKgeaYPILpTMKDvnFMZVwCAHKi+3xCJ3fCNPqa/rq5ItRbg
BCDS0VoVw5iQw2jAjPo7xHv/eANnDB49BLovcKzl44JkVF3Bt99VLlP5go6SrH0M0eXg50aT+n5/
lxNUfoYrlpQXBW37EubAPF/q1HCzCjr6XsQjcZIliDwsoz3zgPJH3e6rsa9TOjyuOtIh/n/L1Do6
sq4UiJpcNoIroRZcdv0ZPEYMQty8yd1Luphz60zC90SvVx+zh+8OQFVc4Y6jaM+cvto1JfgAvAS9
cl/W6iD/IEWSCFGUfltCi4VzIY5q+OJJBK3qx1DNn+sNAZfBDvyvCKSmzj0qQOjSrviqcFEUDjoD
W049r7aN0CmvCmQjrysiDcP1brNBdBqPIakM6Es0hyleCSBfsYpU5wl26kEs59B/LJNAuEh+as95
cnv++FC87ZqD1PFwT3R4O8pxulgEMVR0OFNEEj3IbDmahwh90nLhHCAw3exLtGRYjVhma8djhbEw
+591RAFX0PqnrivP+Vy/IJPYQ3xwcEqQgM4Mw0SPEXDWvHRU8dDGGhHS1HfdD7U1YKo4vVHNzL+v
r1f4SAMZn77u1jHFSHUYt6vlYo5fJ2L9oxC25DjHbx85KufQ5SrBOXiAAVIktUuo1w/S3xnkieGH
xVdp8PSJ1aj4KLNDaPbkEHprAY06IG6zOMq6hO3RuBslwofkjFkXBBVeyxGCRXDBu/mGXG0GZ9fw
eetT5yj6ROnFot1bzh3gG45SJyqbKoRUpv93PWZMkmtE1EcQeg+bms81Pnf/q/ZamCvixEh2cMZ+
rF47bBzsKG1gdEYdgs2cb6EdFKFGxM5QLt5KKQ2uUkBxFZ/r1/3ZPK2XGgj7CTLf8MRxx4Fq0Of2
0awC9BDHEd+v2rgdZdg59A1o/hLZ9RZzpZF082U76l+TBeIgOgrTV0mOFb3mXBl8oHyR1XvrLOUi
wc3kn3BLqczV/+DFBQYpy3KVRsTQW1eFbCNvyBls4w0dfIG3Rux0zWPK71N8NtVhlU4/DxHW5H0l
p6NIevpcpPwk3EX6AJVRAZPLJwf0jQAGNS1R+0LBcoVya9tQPbI8KjyK3k0CK/zgE6i3+/exV9PO
BClgY4LTCPfVTZcYcx6nOH8yistliVSRztrQ2cYLmKi377rmql5lfSCrgILe5PLM0j/b/eoYxglJ
08NunFG+bdd/JZ+UHSJ8Y4hfgD7NudB3joF/AMbxNlmsGNT5MxAwrM4pk7fNaVVEt2jRjl1nF/dl
GyOHaHC4MHu+QwLfeVkLcF7PiNnvsz6+l0PfVBgQR6VzpvKjEAtnWB+Xm6po2064/YTPCB2ekH6S
Ui8/cdD84RvAxkt1HUAGRuV45r6L47Ckiyj3yNZPX+w2yEN5LVFj/xE9C5l0Dzfkv/IyRf5R97zw
opYNDgThDJcuVIY0uOo5XAaUmBQI3N9SFlqZBBcUN9m8PRoph0odSjmF8UYN6rgxefzppPeHyhPU
tc+dvVQ2bzzpmC3Vj7n807N46q4TpLiV1oPejflkyrdjqbxUBdX+sgCNvA9lHJC933C+yfF/t22E
HA71CJAzeBV2/fSayi8tFW5YD6mtmACdP8Q7sxp3gpPgcoUQgG641SuiJiJfJXUqLd8b/Wtgddsg
QJP7INGd1xcy1gXgGjsSHdiwRYBph1pOgM3rjxKajYUvovMQBvzwMzazKjNZi+fvF5KSf2OxX8zc
G7om87q12sHJLAlXQm60PSIiRW02AChFxvEgIQGqtK1ztv1PI/7kT48E8XdKP2Q3A4lZkBpKoFnS
KxIJssz3fbYR1TngtFKM5cWL0v0FTquN3zTa5BBOTzKSyL8FXiD6zer8aATAqip8OF9k2+3x7aSo
Hj5AuVFm2YDhayHbwLaKZE6MDJOivyF/ihmZ5581Tx8+1C/gcth4MGEzpwqAQEr8MgQKm0Bs8yx0
EM45KMaQtgUfH6+zWJ4smQBOk4hry03+pBa7awslu2fTHXIhUkgYGv+GMSvxUTCmX+TzpMEKYFeU
UjyNoNTqQnkzErpcWa3czDdtZqtNH08SFVtBtQluIe6IZgR/gVg76CAbqmNgtjp/+dpoWOAbRqw0
j81LZ1Vo0sVby1aFJrbq1NRiTRkLoJhP8fWE2nnJu7bGY2wu7c8Xv1IgS/wpzFj0wmSkfdD8TMqo
3OCgJbidCmcvxD7mhAMgXAuM+R3wRUFZNQPA/fwzOwRSYtx3rb6Zl6tQlejdT2+LngHi+a6NrFZ9
OdJPcnVgSWGsx9gBYJYkch/Z+XW104sKCQg/qXb1DOXyiwxefcMqi+k+TFXHUzUoVSeo5vVZd1pe
M0tQ/ZnOZFbFJyLkahvYC1uvyakrSXJW97hAREZwL3MI9ZcK7+/u0iAQY/HPkYpLkYINjEBK9lmi
4mBxVdmFxp6qIGdIuJu9wStjKxGe5LqrYi7X5MPz0wesUrF9eTUWMMmDgAoGsjYFFPmkyLPiIXrr
fyRsH9oucvxzcf5oe69rZU0lfke6tNs7MPtNt8lYv8K+iClMGXjchybDmVKJ829XtNFSQBdyjwTT
mJySaQ+z+WFdQQUkXh0s5NtHQgNx3090oMd3CONVQAjkhciRz6pIEYZr6qT4cs0UxpaCXTdnKLza
XI0LLsh9a4m6IHO/xpW/QA+B684ssYMonOsHV9vf/fCXNWwSujvZ176Inv0Oo3ryu4kznQg7GCUx
GkPpr2VwI9Wrp2rGkOM71OMjgQIWTSyuUuZMfAylYJifT6xZDypDHjsSjRefiZJv6OeAMS5cFhuk
bAwbxVg5FNcNUdJNUDYsqjpgUoXFALu4LA5n39D/97Pi73+4KlVDXB+2OHFwyvh5lOYmW/eIA98f
uBLVb4U4v8rN/wppNfD0asSEPH6Jct0wrt3aqgf9uFmeZDUQI30uBw+/0g1WbuR6Rqu+jDpS8ULy
Ojj857ccINzbQezePm1VVAHvCCryW6oY225Tk+wVGwlBjszuWrSDkJvnlK+1jFV8s2jIphFbPDtw
PGN2joVLb3aDp06K8NmkqDl0nSO4DGGx6+BCNtMmLMKKw+PAQ9BcNQV1ZorVuqvuyDChlW3vTfVk
zzznmCLtui0O/FyTAq0ocXg6AYbC9gje8Tnu0XLxR4KOMi/LIwTq8h2b0sBFeaJl5gJ0UTHVwetF
nVxgXG+605ZJCykJpjgzrnZIBvVqUqBMaMFYhtv0dIgZENYzA9yxgpYPEkhCMY+yB3nScp16jMVa
EO2lL5R5bT+8tdvzZ23akqIqiLxdwZ/YEf8RkGlITPdmkfU+A7edPXJxy4Vlm2z9/GehhCBiF9WP
mQSPk+UfzDIBd+hHDVKw7Xyuyos1lVua5a6uWFtYc5oWbb19foZKiMwlj2opnmm2GDVgrK5uMluZ
uazm61dBo+Rl/lfpLWsX2sPJObZIoE1gYnwn9oNBz740QtS4cmdU4NLSZ/5VR8VF20OSVqcpcudV
9wc11XfzhW1ySvo60vEdK/7JsHeOW5Vnw9tKl4evZ+6Mgezk5ap/66QWxsVAqEQb8UWkDC7Pvb3n
yT0fZPEzhFZZ8N+Q4m5VInGH2qalLput86mSRd7+W+O6UvCUuSOVaP7xAv8+NLVFSRulC9/zOJ9g
8yyreRoVL3gmH672OOvYoArb4NVl5IxcVGIz9JY69bQM2lYihVIFQK9Rg5/80K0HMQWXT1eUoetV
AlAJ2N6Sa0+z50B5VNXjW/LyfblZjlgas1/c2oFKEiU1bsMQR8IDsWpognN7D/2OK3GB7VSAp6VU
KPn0JjlyCD7Egn5LMFJFSSXz9D1hvWjtAPHPd05hAVTzMgUs5ojs3574Y7SW/ZRSRR5Lo8e0spVY
L7liAlego2rKFW9V2O5N1KFVzHn5/4zb9S2mvNayyONOJdRgciMPm1cLzrdKMoBS3HJH9po8v6sb
s+RkOpfSrOG8rIJTU/Bx6PDPdRdDFPYhn68Sp9d9gUkTKUHp3ADEIxae2ylSq08NuuOM3dlNSnW6
lTIuwzerVlKU7IOWefjIZdZtY1gwCTyvstFW3xgWkDiC8xJRDUrtOXM0eh6KlkJufbQlylKYY6kP
oYpey6lE+yLheOPG72vNsZsfqM3liOuYNU0lnqLrjNXSvdHXfH+ah2Ye2XQP7Kn8V3o1D8TEjhVI
tWEGpHPVfxMRzMhpXixlBIYCBW4d6/FrfiU4L23Cpq769yNPwSzVVzUdp8UMLkmtuvxNVKt96NMm
Vg+Ke4sXDV7UTIq466tXPzOhOiRtMH519c0E/UzBAu3qlszP791P52/Mt5FcHMAT/60vaPlk7CP3
3/DFhH0nG7sm1aTafItW7/oSEWXgGm3Wxf+XBZvnSq1qt/VWLTjPzy8LqJIUHPu4yOxMTQGCIf4F
2XpbXnAgJvOGGUqKxFfEG4WE7sPcL35AqyChDvI3M4aa7HeKXMN4Yme+VOX4VPO+c81kd0jtaxM8
aY3odpkJNmrHBUKzShzLGg++Razd8575EqBTJsLeQ7KH6vyS2RapdxHip1VzcyycCvnff1V5jNW6
3jxv3tbkcjNadJHwAnz0/iZA4DhqoywaM2zFQP4QwIJIHuA6qmA2bS47bmKDl1HBMxjcLg9w60oY
ZreANZVkyXv8G/geZA1mkn2YhmjeQqj5RQamlrXnrJYGdWO1+6KBBmMJEVwT/qEookvIjr1JO4cg
bfnfLDFbcPnXIqQhRXjw3K8aTz8ZutNmMzEZ85Big7JTL7tFU0WoeGHRXhiLEwVJZKa7zhNH56PX
/5dvdVhmp2vDxK7gdDMLijWDBH2mGopiRbfpUTVXUg0vQxJ1IO8d51A/5oQcSCymOKdxSSFDgTbE
dmrmmPDlFfw0aseFIo154PTBskvrcDQ2iv4mI5IHlJGv1v0X+wqZBwe4trpYlPxIK1lfSZlSK9W7
Lg7Ounb03r5ed2H7jkLqyiYkvY0LrAwJkIE6LE2bdyEx+TGVNjXyR/pRTQnWqJe+nHYMpFS0Eh2R
1F23PBJr6GAKIBbFTnqIlqkIDbbxAGaH9u1CgXzKPbca1+YMZKH2G117hrjg5OdSjMVwqB+teAEa
kncJXJEjyrthkbpuSQnh/T3N2zRALqYOSmI+4GZHYHSC3WkzRXw38wSnWMrNpftjQl4j/1N7O4Jb
iz2q4EbwFr2+O+t+QxmN+AU/pMIrFp/LFuVCEUrjPs4tF/96yE89DjmGWNM/vGjBkSj6snnN31i4
q2UtmTEt3VFB6/8jMjXzfRfaYNSOv67j79+57vQ1QS5S20PydV6oaXDY3IEALJiB4pbDFCDHd46a
NP2BZFn0WiVskfoFqmP2cpPvrNFQZCgDJ+kVbM7aoO5oDRwbMtModVVzt3TJWMTDr6WqAr3O8H4Y
NsDkJlWzxs6Jk2sVtbWL9YT4ed3Usiq7CWKc1KqpUGcXl+M7KTXQP5/weXKFQUyuuABVXLB410Q8
FNGIM7R2/2/A/h+V5NWwmmgxAHm/pzRhqYDLJcJp85WzWjomRMLmXV1QRu8fevmwz+WVLX0RLDfs
7CBk0ItR/lKfXTFX0tNrNvIPHegxDbsgzl34FYc/q8V3C7Jrm4asyBdJxukdrcJ/8XCHPxhASWVG
Prdt64XxM5nxL2Z3Yi1qqblwpjlEQOU0Y8wcJQfxHvHyQP/clqxoEms3lsuqyFN81xgR21drxz/h
s3OiB4rDP1KUtogtwwj6kLpsAYIPfkneMW4/cEf5RFTQNdZl7LCZ6ONKMz/Gcz/VuV9jP5q2xdYe
RJuwOs/2UHiKBQo5Hci7uNmIxTfxijcGbkGonBCcM4x5uOREAkBy7ryP409KKQuCiEBn+5gACLZx
kuU3Jx/qw7a3NwLPLposcGw36KezwCyJPpKL9iKCXD9QoK02okrPFVH8pQlRVAnlgSwsVAhMTa1d
tvSaB7al3/r6AfrhPwS27kZl09j0P+6TaxNP00E3v94mow7r52rO43MO8OZYZdJoYU3HX0ymgGAk
u5jaf5iQcHA1o585NKYX8ADR3rj3lsVXgr6qKG/CZRAQfwvK6wzb2bOslbWsTegptS9x6y1DOnU9
B+THSEO90MT7sPMlqDkVGUFj8SAcnUiz5pOhXHaKpb/Bfonw3Nu2Xx2DzFYjjv76ugbWyFbMBqNs
S25XfEg4H3TUQVu/urW9Ao76GzcL6dnjQUdAl+8FOcZro4BjtuwD2x9aV87QGeaUihiAl7YHDHpq
e2wuJdhTYU/83xVfFSfYBgEU6ER8zAsbVoazbO+AmrDeNm3tTyuGc+GZDkvczqkT8sC/xkLSKOo/
7IZGd/542jSam1565AAFI93bLfGbHRMz1C25f4NeQAuQrG/IJL1IrKklyZAz9H3E30m6rp+ggSpr
uZ/v6hUBkdLgXwYjnGdsKK8vrOmXTLpimwbp983xQ2c5FDSZIfRD79yRAmeLbYLWDATNQYDINdXU
uFojckOy3z4t2+24tHFNSlftdsUWeV/pI2g5xbkergqwUuldhq/kJF9uzvDrs08A6z4vr/jHXGUq
YRAaWC3lObMiz/JESjqNoIQd/mS2Syo9r8QMnsCSfQTO0iKmSG4aBjSPlJZ+mKBVcQzNh+amQqY9
MQyBTKr55SU1HJgU0fJaldiKw9sJJU/HhHKvh1FM2WdIAap5VAUuMnjNeHugMo6tALJzGWhM6BHw
qWK+idlyyWd8c5tP+ASZAM35vjM9NBK5SWPa4lRB1AuvHWpqS0bPyRL5ZsaZ3s8WpclHOFJvcxwe
6Sa/pwKPA106dHubqCReO280yjG4EMOv4kLedfa+8yziGdEQX64yiBeTf94wNZQJ1KnsWDw1pA39
WmcqGu3TU1XIkE30om+LyrcJRAOKIIINlM1k7cgRlqv5baAmrN55WgxCrSomNiz5HQCZuOisyDCv
rwCW+YpPMZF+tHr6V/COuf5YQDgy0VqIIL6sznunnvmXuMb8w8Gh7NUOGdQQ9BX1E1t/a6Q0iY1A
DigoACO7J62nIAUy8mutcwD4G7JcYKLMuPv4pDEEvnr7kWMCn/UMYB5MNiYE4HGqyUuWWZizyvmR
0XzEUUNotiYpItTtLJCWStoKu/5iBUQWzHT3jbZolankqF0h22oiLi/QA59tC7uP8cq2t5w9QjMm
kYT2+9pIh1vOnWTtgzvNTdCrX8JI+oEVJ87vEeXppkYj2OctJfgFuzJPnuUuqcAHkPfy+6eB5woE
JoVwFKgp7qfx+Kx/aRDnVVa8q6aqMInEW7Wa38NkJ8GjD+NZzJGaINfy4qhdH7IwKGLwujRE0I5l
aT/HMORfjeFOR+ayanOJze3e9pNTp6I7YziPcIVTsIyuk8/KL0BhSZa/5TTPMeIBuBDLK3fnBeCI
fe0VsnpAFthUFvdx80fBOEJBCR2Pa8jqUZCfE9BtGYYlZLtiEz/17bLzj7oKufeEzyYGwgT4aILY
3cTz4QYIUGEgT9JRiySeJxilrzgstjdOn7vZb++fPMmIthr5mR8lOo7I1snENFgBwDWowXyzAFLh
1ybL8agh1/a0Gbim8ToY56Of/ilx3a/UcfRrMcB239a+Zjh2JZHXfmC6lcCx9564leolsE97uDw8
HBbWNYE4XUNH/pBti5pG5qXuYMG3eVXQcE7323q19djFaq5Y8d0/ct5qmyZztgOFs74SaOW1kqOs
86hBYfOv9j3XycbU6CR7+5Psgo7VLpv7c9huina+uoMZwGdekUrz76toAiQqWng+F6CxdVtDXjqY
5CZ+qjE8YuDVqU0rsnQ7ZE3WZwaOqJ3l2jt3DB4/kCXHIVSlTWGVlikB2+VAN1ZmS6yP8fxdxVVk
LS+llgf4j84XZ67l7tmnXsCfkhZPwvZgzfU0b3/6Ev+yKMNWgz0XA8qDcRy65Hm1Y72N6wOqKiVr
te3PgpR9ZXwkJ6nEWWWKuCF4tHWZE+tnYJr5cs5+DdOqoKK5YAS7eDqTYKrLZGay6qjcIZZpAKbZ
XABQ4qWikw+ovoo/UX/iCxl3Z9GEXnRewaIZ70gHT65/khKSrUjWrnkMdHy7mmCag7+3lXQ+pWFM
fNyt09HFzX6hQewdLjbtzbHBWsKtrfo6Q5VculHT0vaQ0Eh8zlUJjGwcPRd6LwMKoM+eX2RYBD3z
LACs4glatAZcfzJ5VX6isgxE497xY3ILVw0KYqEw1ffiD/JKjrxHnn4qPm/MF0IF/Kz8jgVzQgKv
vEzZqmdPOiNfN1ZcvW8CiEtqQUxVD1XSMIpns7wIPbWjVyT6noM+Nzeo6Tnibxf5rEXFV7t6h3QU
MYee5NbO+y9IuJeaJ0GL5fNmkbLHg3cU6vWZBWBo9s70ilZt3+9TGZid2VxGzCmj7sqBtlVzlFmb
gMi39IEnqr6CYAo+lHFhkV5eYJ8/m2idAF7SiFVh2jzllFyeXPxy7DOPgH9bvbgP+6OVblSAhUvf
cbWZQKYjkEOB3vg7WsJGAZBkOxmfseZyYAQoQWIlKeL0auowrqnUGUQPQwuj9FVkfPkUD410zopK
RDWvbBEbWgazvcXvGCxuKT3MZB57Pa9br9KX3hiWqkVNzR9IIh1Wo6mGLsWNS3Tt5meFmDbFxFQz
cs76IYM62bpjbZCLbWUPljI+j8qLiWsQODPMMwOc+746xS0WLo6HDMG5KReMbkNbn+29w742y+lp
Tp3A1RRL19SzeA73yf8LpgjzKlqrvaehZ30oN5n/YBmr4Fz8LDDUYkJTbq5LbtfQT3czL71iaVyk
um5X74oD9lAK5Q1q7dY4bWeBlU7nqoqZB+4mA/yf2SA3cWbKJVvyd58ZNocHrAS3EfcQ7tpNXqbp
BIhXB59x/Z0N8ajliclYkl5Em2oK6QTaxsRW6ErXG8YY43J3fAw2TdTOjuSSC08t6DnCws5+y8Ec
XWGB4QsGZ0VSs1k/Fq0Lg7+EtIgbVuLJKMU0synOORl/IiTaKclwNrLUi4Di0CoXTN8Pc21nZBkp
POQT33tzoTRjLIpLPmTEcEWbLhYAobrolvY/erwlPPTeRJSt3FmPfMhPj+pMkWo5h/38s4OrjeT+
zl0OAGRBLr5K4QqcfRHkGQoXZWCdFgDq9sw1Ue3zm84QZFKTXLeZvEvtH/hTejsvaXutD9qlPeM2
0TJLMKnivfyC9C0O/NIjP77ePhjhu3C2JrZ5HO7A5WvCpBM8Bhr21oRGblzcz8KFj5k0Q6GYOG6x
1hzgUxaUgl2O/LzA8YaTVZIM0HvWgZijcU2r4HxlcydBy46Ka0icf6GDBOHICDCmd7qdSTCO839c
d7PeUaCLPvSMarcz8KnI+KbZZTcL6jcGo2tqfBGcwUH6FAjFMxr34wg80Te+6blXVp5wUjh5syBu
BKWoXjWk17pe4SxrDWZPy4oDqbWVNlc9rVQvLExuXomHER11nQSD9zrcEBhhZQpPEWSf3/CJyMrV
hS5k9KiegHndDYeWKt+j9rNfgKPU0tNzeHf3Och0llD4NiWvmINdSb34WIulezRsWb31zmorNIZL
FPskysZzKdCXo4ECxMJJ7bj740uIQE4T+fKT7oa8N/SVYkr319Caccqm3BXKaUOwEqqdXLd3bLvk
CURPWPy0ckXgRCloMB8ayfwzMj6wtaCp7dcueXl3Y8HW9yKU282uwVXgH8MfeZ45iaasgeRevX5S
URD6X/kHtu5r7BlSCNrsuMaMiKrb9a9PvW87Lt4FnWhWhyYfvseLxrFWAmaUmGRH1LXnZeh3GBpF
0AY0hcELiO9jdutuVuKYY41FHoHXWQJGDffGsP8eun7olU0xD94/T67BIp49RfhYiUwrXj/eAwMj
mib3JY4CG69a+unK2fh9mBoQ9Od2HHOmrTLB0sv5LTu8n15XkPJgiARTSqJXSk0LWhCVEKaBCYta
z0/yBoeg9zfX413FwO5UQH1G+j04mvkp+gI6Hnj22negF4r2XRl0SKZFNlgdNzVvwl5tnWnyAtKG
Od+7zKW6XEE4FjkrrUmDIHKywRB6/u6rADGU7Z8WAoMp22s4J3SnHiNx3Ok/YpnKXMdJ9oJxLN7V
ShwYatDNYQDLMMLBdzcjwRJ8Wy4Y8iuYPoJiO6bIZNfsYtluqbZmoo48NJPdwbidYgSIMUCzYzUQ
Yjvw89BpDx5UoEVj2BONYazFrnn0WS7v5R/fe7IzAAvsVyVPZOOm0WPZ0L0BbKFwR2lVxsDkQvb3
wvtVOhPKM92ZrSeJ9B3UOz4EOjzjIyFj3EfqDGLoPnbfppWRkTh7oupZPPAuta6b1yPEFKh4aLtU
YtvAnY8TJNSY3DSJrCq8NmVbPdw0gQ1Di+6ZKtu9NHebKoQKfCri4jn84ZWCwW4uGeRJvkFFG33z
/ecZ9ABeiz2BWf9CSnotVp+qaGrNsHfSuFoDFbIAJ09lcb5l8LkwtWipjsBed4zJQltVergAWE4o
kVXb/ER2JsMvATFPyvf6DHECCXku473C3usSgJMqrNqzM6laOV9nhd5HumdQy5OEiWjzSuSeO6Uk
QPYTnvzf4HOZDr3b8oimbA9tA3FOczB7Yaa/vhvLrEAz7dA5JlJ0zwcV5/NZQSiRDe7Nr5NOKvpG
/WOigI4nsmOzADwT4TZOf7ItQL8zKT0HMCpdu17m85GxKQ7tnexJUGGoUhnrOrNEVmedsTsOsqjj
QGmWMllZmxBp9IbdK87TPxpeT7LLPZiO+F56HUKqfuoCvPaDA6nB5nBKS1aSg0Gd0P1fwBd11uUE
lNpuZmSmc8svUqJMJ6grbYuqEbB1k0ZmyxuGGIXJ3KzGDXtNMEce0O9mxvRVMWuFJOR6+xxhQEwY
fLrIHE807wnSHWWGKlvlg29qUnov7O6pl1ZwHTMKkNYkYs4TO9eFupAsexmhcX5+h7xXWGhOAFB9
OGVjCmwk2lHz6KM6PHUdE/2i9G9np/1TEDmo3w7TmWXCisXmNmGsdD1pbWRMhs4i1YU+4zXwKDPi
Ryl0NhoJlLUVKQyfsa0tZ3BBI7WBTDhiLPQMAQxCubt4OiC6+IUa96DxxC7dPB30Rof3UDhRd//B
M5KtKyCSnQKPV7uT/3RFtLVXowDSwo7MBb8aEGAHFwCqyph5OEHp6ZeCNH2HbnqfpjGFlEYW/AiX
afdLicz1gWa7N+tNBN7JXqg9zTSaoqMW6jqxTb+m3ixYOh6HaE8+AovDLnOk9Wi+MEtLehSe75E3
wCVmDH9Opv87eT26js0i0ZgOJ/7Ac7kUXtXDD0WRX0IF4yzeCDIrgSdjnH4QoD6rZiJZIf2N2ccs
w8vVHfnMzlIlrsFNZTLOTDrhSLCWULAY+LN8py5GE4KgN/CZBt+s3RGUu4VM5oYJ/aWTWb4/Rh6F
9ENg4few7ujzM53ioCPh+B7oS4mu2jrfV86xlpLZdxeVUm6R0mZzhO7iQdPnPQrnjIwUlcm/GXb7
sgjL1Z8zOKCbir2nM1EyUM+v1BFBXvfIHrQm7HbYzbf7ZWy/Ta/gSjbBdg1lNDDtjFWRYC+jJXKB
nJHVg745+QMSExBYHFkGhywqk/jDfDIBcQJkVlWanR98kcMkHKkpzxHtRPVUUe4u/QvyQZ/eZbyW
L/uiSOjEB2uOw36Ah+c90BFVjOOGk7FTIo9NjvKF/tHgnYkeW05uHcm3AzyRpIArORSL+sYtV3Nw
fGRoEsLYuKUNerRFJxOFWDwE9u6ZKqDwxQ3FMgicV+YCdwGEz+cpFyXRfhTP6ziyl/vxlTrRdJPq
Zo7x98XzPglRWVmZxPzh0AmdPL5QirmGILGsmnAeo20CPyNwHbvOKOSbDzzxirRLlfgeHPopaUNf
1EgSN9LfpogVBbuatTSFl+na2BR6KRQgn9bazHsnRopQey5/OaSKyrB0ndbueXaXr8eymi0Us7zl
b02yXB8wOAu6MjLymWxskgxBoh9jtDhlbWeFLQGL5hzlCdjcp6xnPiFQ8CBIkib0rJ4PdmtTbhZH
7rx3Rmbh54vwUicKkPy0ydgAjSixAWneIdLOvxWKqLUOy/od+fviVumMGukTaOo02FSaOLt7rHj7
R7bmqmlh5Bp9vZWcwBxPMjMjbkJ4X+x1GHG+BZ6xFcOGb2lV2pYRvIt5B/W5WE3uEO+Y57FITg9x
1Zgf9Bbs/+67H6ebusu/1ZGFGRtuRvOE11tptnkDBij6HlAhCVsbimPpvrmn/EVze75U83jIuXTI
CNw9Bt+K7q0KpcCCH53fM2M9hBufBrz/RYtY94TEXUzimwhbfWKE83PHXDJk48SkbVkmGp/fSEcv
qPuCXa+S0LzrjsxZm+alzGbIlHrkuWQXRqv6qTH2DX8Imqck0saSrOcmlp2QNRbohbCLd0ahNtHk
I/UnTZcAmbca3SvuX8s8Pdpnk/qJaDahmJ3REVIJDRy+vOfn9hdT/CnuctB4hLnJNbybBcTTAtXO
eauVKOZphjsYqMUOfDEfV6dYxcXld3BZo2wBg+4TgeLFthMICjwLK4FrVkJ1Rv1pm+xanDI5e+IJ
YxFvuj8DcuMk6AiBog7Uzxib6jhlf6BbUX6VgsqhRQUvc+QwFwxq1BC8NokJm+NxHIrAyqA7BvnD
i17Tr0A3/zyVNEU+1a8gO+1/SMiuM7WrXj5shuOuAN11AS9cwiMW7wKXIFKJKZF2+ilolmn3iU1H
6exgTQVex93FJ5fPIESlQwAhZybGNkTl+VomEH2s6caMqSIAHATYwxWoDO/apoh3AqoovdMiZXWl
F2ifZRvAeSGlCFETcUGxhoFMQHtg5bC1/NWzWkekNBpLn8bbxF8fP42GitC4gZNZeMYxtnf5PAt6
ZyTP9Sy/ZIvoADWSBSDOac2/QaU8bb70XzQV/hC84uMYglm9IhxZ4mrxAJW6sY+SIJrkiiwqE8Rn
OVr79SrDMkNCJTXIUAOkJkZLDGXy1J9vye5qb7n/hSKhBlwUV8yZ5Cw0cNikscgZVsWnDxzBAhtp
wAOdI2l69z91Ud6+CzyjQ5eRWndgkGO+SB429MTjis4bDfhiZLw759/n0IyWRcds6LpmiD69SfGX
Qky3nrQdU5xVvsr99yGU93fGXAqlnIJNq8oI7H4prX5MBQSRtEwpCCfTKrxjX+6MnUDkTjqx/Y82
e2+uwhy64EAWTc92F+iXopWgOCWDahM5p4vib7pM/xIe5rMMIccGrYcmBSD++2Oeck5fUmUUhWyi
wDd76/DIiyy6PF+ic2+CyQU7nOMFLV3REW/AnhHWJjNzaJLwBYIh0LngWI4HhNCHfaPqwNTGiWQ/
1AUBmtI/qpd5nrMAw2POnfbgVeb93Ct0D84CRtlkcxzLGCfOtoVgXqt3sKUEcm7JdUwNRRGTVVSV
2zBt+o1h/PrgXzJPm12u+FdyHo0z/Rprm3Hp3lOit0AdiF4dcBw8LDoi0sZI/p6kVzwUsAwwtGKK
R2xNpe4e22jzngWT5kolC+hLzwfXoWJmB8lfSj53lA2o07agHVQsmCPzm7hw6fqjwmLZFuHZwi2E
dgvAz9BJV2Mypzx2WOrSM8KNFR7/W29RPBwHklZGXvl0r77eGDUyJb6jXeMfr+77s4wWEZJhzfRF
1Eu1j80SRH15+TJJtSutk5DI3FIUfpg8s/PemSGZItBH0jAnbctk8jMNgKvDwUuBfVR5VUVrW0Uv
xzbLNgOqgA4iVuZ6T/+VcHEkUYHknKz3BleAkNus9lpedYWKa2TexS0idjaPztq/FFR0zNF3BMqE
k87wcWvhgWMTCcVR7NUwZhSF6RdDUeBCTletimnPkC16kQkNVVafeDyNIUj+t16f2LB+mQ+Oqpzw
oFb4vhrxTdH8g9s9O9HMObqL/cN6+tmq1rUPI4skz10tIBoPTPJxdv5KEC45k019Gq5xlSY3ZVOD
5VKhPZpeOhPqooefxLFXtShoEuMGiA7Gbh62pTwO4hDPOrat+JjbsH5wu5asZgGu79DpmcSJ4Nhb
N1khS668Rk5J6p33qbsE1lG9TtyuzMXLEJvmnXnxh0LNC3VG3yb7ylXpJy7CiRspsR8fO3fbnFe/
6LCA9+/v4qXMvosdf0D5xZ9J2rsvd9LvH987P+BDr1RcWkNvTkH5tqeEA2IBweAVSlGvzegUSzJe
V9/eGHfx10DQRAOii3+an0D32ZGNmSsDMqLZa3vkd1ZhzRZyR83yabx+nMADuHdMbKnxgQ0V0FSf
uz1ADaTYS+tnDM9sU9TcWPfU491pFaVgS86MBIxhMxSjwKrhxeRdpWNAav6sHTOKYrDvF0UJB2Fl
DrfhbSzUZ3UhrV/fMBgNy+LdHDujgdAjB5Z4cKaQ44wJ/zVonjakjKhfjRTRBZUdtNU4pdG1hwab
LWI6tJyc//uTC3dDU2P/vYUrFSaYlZifK0IHZ52DKzNt+aeQJO2a7KQMxBkQyANVMEAMiYbjipWb
vu36qqeLgcdTgeMBRsjB7LPmZuk9QNNNuFW9Mg8h7ClbBQNwXo6RxOwoX+ABdaVMUlW/e9dGzAR5
8GlIKAtzLXFhOnlhZDU2rnSmCT0EZM6GOLB88KNyA7tlbLTBaUGHKRUBG4LtF7PQ5KNmrDV8rbPw
09EPCkdYZKvBRbTNUd0aR0WxFShTY20qzLHhXdAdbTtgmc6RdCB8GkELsCfCZKAU8fWaRJ6HyEqZ
ogeaz7Om88OBKx/yLdBCNAgVEIRqNaRWZRQFrLi5s0IvOWVZJFLWFBbXVsFVcmZ12kJxnnDhkTjZ
RBcxk5nuOqiXcpuYiLgZ8xXWNFfgkWQEbbvx7Q8UyoTycZbrFcLOAczmKtFMfStK1oiRxbkzMe3u
UU2HTa78ZXYOUNuckWck1Xyp+GAi3vviOOt8nELj8ZfUraNkq2bksn/YZON1j78r+wWAAHh7SeLj
83F2fIp4Q/ECI7cdPfnlnXQn0LdLMVnEcCfoBfvffoyWQ0+3Ou73etFgNOtyOyVpdcS/wMb2P00X
xbHcD+mdcSiC7AX6HE4K8O2IOz5RXb73ZAgNYIAb4XffQs/5G2MjSS3ob2VcfvDPVhk/UKppWBG2
k4yccg4P/zHS4iJp/KBTWzDi87Fhd+ECoFwS9cFBhY3diSMFlF1x0Uy4ieLebkL0La9CoE85fLMV
WOA4KPJwsL75mWeyKKrTZBuH9zaJc07HketFaLIA+rmIU1Gw/YVgW4gE1iuKepoPftOWqER4Adq5
jef41ArMHn0rPAwEVzkIsyxn7id3ZYcdY7IY51gmf+w1+OmCDFdMbkTK1xExxiguAzwLC56DsXD6
87LPi5To0K2NEYpDWpM4JDSePfuFub6KXlo7BCzQUJaYjmk/wXVkMoFEuS2J8kKo6GBV+HAy4KfT
EkWhaCLVkTdIpKo3Mb9PMFkW8WZcK3up9QDxSoz+5fnfyfEkoQACrEp5BCHqmDfRpI7tIF5e60Jh
sc/r8dUlX/iz2oLuLh1o++bceSjfEZUvfgfFaejMu3ZDQtxK3GGRz6s2wYgO6HaKroEmQnsOwzQs
9pPkEF48KKBhaHUAHRe6IVL0ebThBBbo59wUfghia4VEO6KjhzGx39es6ZMPtt8Yq4bVHKzvaR37
Jpd9LJmBkRaNXeIZZrRMuezHHrJc0m9HJaOFlhZbCuh3HQyJRU76sgZ7bg2z2AzyQ8qwracCzXhL
QiW2xqSneke0kjOyGL2MZsw2hEjzxexbKYxfJyTI5h9jkocuEG1tJQBCmsqCyKFvgTQy/cI330Hm
bSj0Ny+CMydYYZ74e1WwQmVAxHtgFff2FY8Ql2zbhZACnBNLfWkofQMsWUhnK963nOAYnW7b5NBD
BYrthj3N8NFVLuQvznQx/kySvepHQjoumQqaPgtmMMrSZmv1JLG6VcNjyEHrncQh4qRYr5w8V3Da
T6qWFFdRyL4DByOtIjFldaEzRSLlpsVbvBakjWiG8fIq3HoxmMit6zZIdFk9iGzbObeTemu9abHR
SszikQWziSBDyihKdPcsW3HkTHNa/4IIeb1u6Zmx+SQSsWzpMUwTOLy9uWQcqHjZonSp/Q44HZnz
XcqCrWlO07/CTNOMtpGsb9k6caEkJCi1+wKhBSXHVz5fDVAR1HEMe4abdyHQEZcDS3wESu778Rm9
dkqKBB5LaWVG6/dZO8jI2TprIMkvtv8eRoLqT6iOQI/H4gk+efXY//iU7e0X/040reTaW1IPAZzi
tgB8YU6Vh/z8Kx1P9ZdHafkGeZxv/dNuy3yZlwuG8QwkFyLZpTebVUONZgeQZAN7RcdD/8EfZ3oG
vsi7erTzKhHo89IFXywjd6SNAXnPw9z0WjSba3G3+rb657res2nV077mwQcO+ZlUtRVNAzPNjlMP
VL9Y5Ipzf9Jwe7CFgkm7K49ZFeQvhJL56hUgtWI0/83MgPvyA1t9BhaAETMOdsJxI8L7Q/u8ORPG
lxSY4TLcyzCLPRjW0C6IYh5D/UD+3rkpoHMpH1E8kKMWyir4tD9fwfFdFcZTa4AJzM6ibSOAzN5o
47AdW5fXISR7VJScT4eJIG4cELtYRnImjyFXTmu4NEwmCxDAKGxUxF7PbTLuCjSU0ZwQn4NlqNYk
pzc1YR9THJzBhLg7xJj7xloYtgb6uvqNMVWt3XZRrXVDCIFOGBFlng8jfjSJ2n1hNiewQ5A5x7Kz
DgR0NFcWYwlpVsGJHOifiKWClen9qW5osPXZmIxWtPbcq1SLMPIMaf+iuHQL3HCtcaLo6/ab+b8x
yzVkYdOHNszU6WFpq8ZD80liIrYujLAj/6ORLSN5fAMhj3qRPP77Vv7aKl2ix16noIVBU9DLDy+4
NczvLxlkoEdTiZB/Ghv2MaCC4U848ejPPWxMZwnozYE6xUR9T1JRVsdR3jVAq7sRV0/zeq70hIR7
Z27JaisMct84ox/wa0VfEgctclfG/pbtwF8lPMUl/dPz442zvRHR/WxNFIS0vGnWJ47xXuu3h1px
jVI8IYTgy9CMVTPne/AZaMY+gOv4MfWoSm08dTXJXeZEwRsdjFgoyC4MBgCaN2N/byDEfcJOwAgm
5lFfgrNrMrZ8vBGjQC5AesmWISYdim+Y3HFWoNINJZjgt0tLz4PD+3E4LmfuV4g3osuyuWvrOwpF
kj+2IQu69xmOBkfE1sFSMqgODZJwAcyZQN7JAIzvYvtUSzogpIYQV0uUCPz3mlYaVvsPa3sMapDn
dj0INzX+RSUibVS5mATeHohhUBDCUx/2ghlFSwMPZf8lkqW8+lAqHl+NaKLfnrGuIE5zngqFd1cQ
aXxtqOimNTVnVk2bTgiw9mOhIM0EHkgOaOAzaM9nwaafqmQip9NRjsQjE+rLZET/2gNrskmcyQgo
RzKLSCEVGsI3clEOMeqt9XkeHnHxQheKUyTVjqBsJIkzpzuWys/tM1hfWKafPFs3Ubz64zjC2a9W
udmuSvoahn6ZtJn35VRRnNA+fHCaL96b3k6he94Z8WTIWrG0a4IFqUu3vgLLN0lrvH7Mrpi5fJCQ
gNOFtxKgbft1C4/9VC4XcFFeYc2O7/IyHa0DZwn4cTstVj0jzKJBz8EH7pgmCiw9f1JZW+IcLFPd
KMMSAHoZU0CjzNIBAdZBpY/efO0029N6Uce0FlxS5iCMD9u/CQSiN1jGTcY3ffXbcfaVoqwsCGQK
Gz8EXAh03rAWx0zsZ1licFhwVJU1ZeBrhQBjabNs4dk19gCWzfigCrRLMssB09XszDPF1RFT0WiJ
miv684Xj6ylXPtFZxUtBXIi+gYZ81Y6r+uvUHS8cp30AvdeRoSoTQO+pOQkfXEj+cQ4ymSwatsaM
CPpP+nSv7sXUMSQF0qaDQww92STWsOJcPOIezbppYSMlXQoniivEd01TQjo0w5fIIWFTwsNNSBD/
FSOgy0b+ytg1nLHfChoO6r2xWj0Op9WenN99ZEtiPgtfQZsirvQUeCXd4a7PHQyknX7F7ouQC6cF
yg9Bl/ei6RleW0vben8uS6LvRwz6BA/3ErITn0URQ3rkJXtqzgK5CBk+VCw53RYOL3AtkpeHXmal
d8hLAYX5JS1PVTXtP8OhQhb6gaZsTx3cL+5O9OxfikYMyi3sys7NqfOtHUVudcWPNSKbeuF2rHV7
AdtsiCUcvMxZszs9BSdzhYqGdmDUuFVONg1o/V3p75lHzV63cdPIttAKZ3MAz7R43WGIHFyIsxq1
SjvGqJoCcOyd74rQMjF6UfeDlQddE30eVpYgoH4Mro5IYKH6N5zubl5TEdkR8i+JP9/0PoH7WcgR
7ADW1mhCIkIl+WHHb1x5Sz1WWWpRpPuEy1HEjC2dTBlzDNJlDDoqwxXQnbq8jOCMQ3zBSeWhx5nZ
i+tdb9GLovAwkBUGpm8tTuK0thiDmTo8XGGAwjoonPkt4XDdDzGcXIdBMRIwYc/6ilNGZ3j75ZWM
RXInapWXWIXctSYOCljBMtiQsFerPW+Wv/UEx1b0zIowvR+LySNKsnWEmf6XVA0gFC87wkT7vryr
DNbW3N4jB8RYA7zcfk/51fBxhR4aeLTS4FcvnybI3KyF/l+VWMQUiKmAisDisVfu8hzjk0puKotf
mi3JZzf5ve2Y5Yo2Y9Ft9UqrqAYFkdzWqKZ2D41nJlHnCcwkhlIqFPVJ8yuTF6E3/GEM5Iz62NWa
p34jPvrNJff+iNn3jUvfAZdd4aaCVIcrzdubXOWlHfappIrNSk1Yff79GQ6+Cqp3K4OKQpYtTxCb
G46xqMRokT/vF+hU86D+aj2pK/YCSm9FMudtIpbVUpt8zZsocmkzDyx77Gbt80PLKwanZyRtujg2
M74bAw8kogDezGLfy2lNa82ej+5UDl3oPof6fC3kCZfroThggLs38YttbgtNzy/Rihuvw9yNwGa3
LnLAajz11yOEwdX/bqFpl4/ZetEwh4JaKGTdO0x+umCh0mqa6OvmHbXHQAb+aUWZewgw+LKPsohL
3QOz6ZIgB9gCN53ZeWjLrdXq0LeSs1Swr+9e3cGpVMn5l+zi88UX6Mfva0cNpXuh9yQJ3PRKmDtK
OsDj4olqzNtYbMft1ifzR6dU0a01ByzhBSLn5UxSNiuUMvikEiZcjr1iTkefb84gJAtyA/AjYXB/
r3d2kRTM709t8hyXG87aZ0wG+ujP/7UdgRtSW4By2uHbdfYbfR9Wfn0SFTxn8WrSfYwYdHHKW9w7
iSjMJIAddbXhcUH0pkzOCOf78niGRdfSSHVJdwR2LQjKXNcKrJWResl5N9wLDRUfh4dL1p+dKIQP
EqIz2GH4vkPRlY14esMnN4aZjn+Sqi+xcQW2vw7Uo6JijyZqFnpJVc7WcM/J5dSk1hg1eWt4YHKw
cZjJm41oHfn2AGA5EFsUgTrt4QcYoexYsnUcDgApXn8BhBWkvD1GyMtRWfy2eNBxfeDkSWl6X+g6
lt41poGVJCMe5lPpEdhxTNRVSYHwqOunnqE5UQD0WKP959tu/Mnte1b038J+ByGsYI5dSKg2QwIv
IJfcR5N5jQb9Q65uFc73Du1c+oWNm+7CJG+B060lgpmk5bCA/5t6+qUEPDaU05tvwlJQLKmNIBe+
roBEtichQnCgGQYB2FqmVWMY9keXUYIYs3hBISZfPvSEnCdgOfwSlUT0C02sE21jmHaAtfPtAJS5
wwUs49yWzV8Ck1thv5kJrl19aWhd80fIdCNt+ZOBghmQWa8XUoW4UJx5OlzOYtw+9M53alGWQjaw
A1VNgwN6is4vrxRXkfZyF1nvTRmGFh87x76s5L5jzuCrE151LvS6kcw0+t7l3xyBLEBXSiUmVEtm
uU1XEgMFk1rx1GnVYxnP4Vup7V/CHsGpXUT0KJOsxkCSBy2og4VO2/+JZXVqJ8IvhBVMgPYVMUQS
+yRnCKfN0rm8Wn9WvjzFu9gsRlEd6UVpO1qIwkS/rVBY3cUBHRCsnPLUqusxiMRlFb8h4tC0Bpcp
eZJOhiCgTPLjGjb72Qh/JwPmlW/CRfK04rNBtoZ6AXyPS0J/hG/6FVJu8xE4cac8yMQQNsZ8XpQP
vm1aAFMOye4qGdQGDLGGtVsmG5zxM1MRBrmdwjihC3xZdZhCJrzVeV8kLKhW6tJW7lUoNVAQuWEm
X6a9++Kb/rt6FSowGKRTkozmvP+kPfJ4mQb3qwxLAdKGjZ19EWgLpjx8L1GeN2Kj0as1RMZAUU46
5kwXphX64P5sR7T57bq88qGJxf9RZ4wRH6X8nGki7oqix8S+kn8NsU0s9bCP69JppygKX378C876
ItDnM8Uan4NrHjDP9ejkwRQorJsPIQTS9OdLb3Rth1Pp09M0jlcax6rt1RCM6O+KqErR4dWmQn3W
TZvWlAQub27a1ZKuBlJ+TrpdDUGAf3WI5hJhotljMu4jLkSelUNKtMs74nKBwY2jQVv09NPLK0JF
LbRp/pIeKFBYNq8cWoLlDvH0vZVt20ADz9I8onSj9DN+x+SKS3QYrwkfMPBnwj0nsOUgxwh9y4ZD
eH6Qg2+vTPGvTXK2u3zgUsllpQZ+GsmwZNDiSQqgm11bFyRaj8k/K0UB9cIwT0wD5I1B1Sa19Rbv
mkIvw2Pu6mSPH0JUu3nxXgAaizpn6Qxuh0/ZRMHOo/y/yMdzl+Vz1gxAsH0ek2+uwXvjdS7aaoHb
N+/2+p7881RiKt9QkyzkB6aNYoHP7/o+McbOnbI5FiVI+QfK6LNB0RsEHu1+R1mCWgm0IWzUTm7l
aTZiz0I2LOKBEtxHFEQyjo8YIB+JoddLu/NuWmz6f4npLvfywk1n3iHpIQX+rbw0hnFcbzzx7/Wg
hLRa8qJ9RCPaed4jidKe/H16sQJKNvEZ2ldKtbpXdH5ylO5/+/bewaA1qi+hcbir/IOt/BQdmQ0o
udkKGIay/UbeUM7IgUb+mStAxqOKTCrZX2+feNG/RuCHB9vDCJRs9XA8X4ooOuXdfBAzxp65mVs2
Rni2QKJUZPemf91rCi5cnZa/+WLFiNi3u+Tsac2SjqxyUXNz0em/Z8LJQ1lKOXKEcIX+XfgkFzZg
W16c9AWlu5nnjSFgiJktBilloXol3rIcvGU5K086IhSBHZR5HF4J3IcadpfhyNDk5kbZez5BBu5c
pnYIcftQ/4yjzw8RrgbHHen1v0i0K8+ZkEOr8Nw5jFpwYzuPF6U6Xvfp1dbIsQYbAT+XpCkcydGn
Dt0aYJIRHT5WD9d1zTuXeu4UT1EWC936Fdp/cs8UHiN2p6wdNIYQm/qGnYw2xVZZ6yBNK2XB8pq2
QUHYVz/Ig8dUwKgt0sSLH9/osnVWJmCU9llVVPauAT1aSRpWCFDHO3NDFzcn6jDkUDrbxk2t9/P6
ViCIW/+Zx+w1lB6n29tDUEfBuHIYtcSGUUJ2nHL8sEMSYdykiuZKCWw1bFPZ/d1BsLwXL3iYMQHR
zJWW0HynyXBI2NTYdctocCgt+041lC9zxlqnwRxJP938xiUfyK69YJ+y6tmObIR9icqbwsfctTlD
RqpSvQpAGyAsaYFTFgJQiP2psiPp3uoskw2XZkyad0JuzC1md909DJjtkuL8uCiQaBCt/YpbKww8
Jz5p9i/av63U13izNZdPHT7FnWzX8aKRPLw/4AxYLGiIPCxRFadjdO2e2rAqrE8Sf0S0W0Iw3s6P
A1Z17sAjxX7vvu8Vg8YRYLbNhQKpmqFQJOG3zUec2gKImF0JdnbojyorOspEW9BRUJLwI8ckEd56
fIJPGv5VFaFLDCKOClcyra1UDPWROqmKzwctsFzq46WjKIiIW9IZn4Vh2DpjDXH+4NODdcwUI3QN
UdPTZilJIqmFF02/eeMUSU0L3xK9Z37NuqmahNGpKYcK8m/aEOmV++udS6b5qnv+jDfko79fB+gN
ygKlBNTEXp/WTmrHBsMkeDy9Rt/AF7kD2hvRHDam94d6YTgs3EZTVWagf5s83cGAVa6e2QFibWUq
SL+bJAG8QFUFyUjiEDxr1g5UNeLbhVmB/Tu0QkLRDjAcSDpDGTVJ8az/xSkBW+i9xFvPm7p32Ng8
qIiWicHXvjD9pSqb3qy7kZCixjWoOzS40c9pvgh71e6v49v9Ptm3x52SLyeHMl8eufVNlCmR3VfA
itSZyu/68uzS8p9LgofAkenZTiw0XXC1atKwbZnmDsUx82W4807AKkNHxd8b75bROpqDzy5cN96y
pOUlpPcF2+c0QIw/c51dxv788++0MaZopoZsXmlk31QYs8qYHv71+RrzFhNW/TNqBLi9jeUFaa9J
C2ywxaCUFwaBepTcOtF+nbg8ZIjKTwOJEQz6pPRSvMaKYM0ITRXO0AMA/KTkLkRK9dTWkjpaN78p
WrNTeyHvBFnUaNJgzWi6beyj1elMxkHo0JtnuYRhxwhkHisC4uEVUN/VwqJIz6mlCyRvY52QQR6N
z+r+K2oZ5onHwg1C2Top8eG1M607X8Nhouw0StHVPwiBLuSrEhk1vSlUb4WavrgrsgM2J1YuHsoX
86eC5IZQvZmN2a1MiQve3jPSbKREwvH1FOd7M/6FNWHau0cpesqhA2QnP4+MmMandWGQ4Utd1/UY
qLuuJJnB8PS/OPtZicy9UStAMe8P1jHfC1gA+6xhyNMoHogRvivTo67Z8u6ahfMprn1nH8L+ZyUh
jm+PJ3U2kGcP9LZ7XT910OvFLFgh+0RXacQAleMjmr8mXog3xo/DsRvd/hgkQjyptUEnueVhSb63
NP/93Sl/bs+nfI1J1PCoR913gvl0AmaxVsxQ+ey+uEeOxb1pDIBWOvv+htnAR0YwfU+rG9f/va0K
n99yrtoUz+Ho3IbmUEQKmYxyE2Lmmm6c1VNxzyBFbUB3WKLw20xOIJfvRb4x5txrAUQ413EOyYGr
MsqbgTVXZjvGdXYJnRqXCdXvjeSjICQGWBuG+Rf9JUTEOgkSTdaXO7f7tO250BN0vZbNZTe4AT+U
7dDuXZRYA85z29ineX/QvazpgmWb18ShpTQfrHjK1RqJHWlaiqYu8fck/m7d1FWiYeJAqa/2PGul
cMeCtDJTnSxfGvrOelxEMuD3YFuuRRc7Yf5JSi6PHDlyw+4mmrk+png5HxoxcMlfoOpBV5D1MyJy
lKOvT1mt9865kEf9JfgY9QNcx1ZQC65FHXOqxBGXGPtf5Jk8+xZm48caf6wesPVPjC9GiNMEqZwD
h/fDwAe6wG75ahUCofVV39DXnh51E0JHQHqvY8xBF30FzCnTSvLvyTFtcI82FJVl15KSPh+9n3Ih
OaPykxCOamVb+pMnAk9KT6naZMS0LQ3Nxfk52xn0NYvXb44okXtG+VpGIdeZOAyBXgnF/hqm/i1k
L7oeZGpx+3UqOfTMMzqosIayTp2NlOJzbXm+/ZMDlPZJho5bVUAWFj8w341ZcYMb69MW+hDZG+my
G0vRQphaOZQhKjI3mP7vJ6+LRHsvbcYStBCKfHsQNwx9Blg0HCgDgjqEDuzkA1DxoKBUM/x9TzX3
kmE08di8/YcAS+GK9nc+lPbB2dRChnBdaeLFwesK1OyKwcxBKptGzrT1bIlzDUP2dhqDVM/MaanM
AgUQFPw9LypD0jmn22P44fZo0B1l0ICT34G0J89gCtV5R1k5bzzkPqvxvdNDIBaJGgx6Mf1Rc+YI
u4Qsn8XH956zZiC1h02dOrAOL/dD+EtmGdxDfwGUT/HfF2MfPsOt6OSCjyCfFQ+sBg3WsbdeCAai
hfebKzibWBTZ76FnduZ9ug/EYNKjKUu8toR9ViKtTa8WXf78OJ1IE61db8gPtuu6y1yUd84E1yFS
CFcAw2e0k4CWAuWGZYtf39HcrERU5zuqzzdpDPlvhxgTtKqs5r4/t11q9Afhez3WAV1NugHLu2N5
IGpXaO889OnCqt+vMWjUl/YOV03HiXFaJSZS+LxhhEOEsIVDh9keW53NwqksIj8GYKhzHCqCX0qQ
ryBtz2vNQV8Oj9pJUJrqGVoUyBbCqGx1xOWZNgdCbObrc8vF6y7S8y04ZNXWVAuABQB+wwfFkXi1
5kJq19akOCOSYpee7S9CuHisFnhtDFcODWwIGHesMYclLTMKkK/lmIEBeCEBR+33wox9SV3llT/s
eHz+0lHEogVQS3pFz1Eg87SiMd2rSmzyzMG7o2FDVdKHYg9Yu2EzppiyRl4j2945OqYo9rrypRVZ
uwp54x6TudIsakv2Lh6xel5IIa9aoevScgwqMb+batWHyC99tnk9I7/9Vp1L1LJCfue5rspy89uU
KYl8T1s3wO3F7pPBt+Zbv9xFNA8i24Qq4AejJD72+ml2ueATxq+Ei4P195N53F6Obzg5zAqh6n+J
h9wMWPsAmJaTSq+8pl917NDeHPQ2N5dOx1w7/b7R3molJ1F627wQt2N+1hC6wWDhS06Gj7Da2TbJ
yjKHwOUgIDIeSHSb6wiiMZWU8gJe/UYu/4RQh7F/7ydrg3lIwWz49yp2S5A+7VwSyf0y4NKRYiVt
oGr+NJpkTUsZa3S8mPyjB3YkB0bkxA1FCgJQR1UbMkSEYwAHDLI1CbW3UUgJTui1Y1TJcQigA+bD
fg3Bo81eSTxeVeE21Bjl+0Lj5/cyxnaUXfGbpVPll32pa9uY97HuxmAOnLsEoarL4eSxmU1wejov
YDHrWiJwwu+AybkqkBIL5QkfhEWe1jEXKxmlMd82h3baFpw3PS3Ktzt9Pjek/Dk1eQ5LdN8Z59uQ
CaJaQeNGhN2lGJ3DRHaKtoujNW4Yoj0WbmxpWCr8T0eEeUzO7AYqlnd1jJmZj6ODDgoKFujgCsrb
s9JR4267H7BLjPQai2U/x3zRj0PffXeqBQ8AI+lC863Q9x7he9P32koEKeBws95QpFZ6L9gAxxjy
RofzrNGDfQUkpAq623T3a7Ofc9Rzkh00tvn7xccDIbRLmZa0irgM1t2pU7/5I3GZxfMXx26yXBbe
t3LLatEQo2S9TiKXKLHNneey3IYrWQFrpP0u+bcb14Qj0cfXQ7O8vt4LRDy5bDKnM2EiMfMXGewh
OhiZb6orCIZsqXoUdFxaYT2VzkBHDaPM+D0Ods+NzDihidLQhlTAFYRmCxxMJRQVQ0LpwHu3W1u6
gXcGno56buBt87V0F0JhsUb1wPKwDDo7uWcBhGnehQabzo+FBXH3n1FCeTbRrku7qVrOo35/UR60
NVbx1VmFvFSSlE5eBWU1OFkHxaTQknmzeB0xyL4cgImhHkAgEDrQWvHgj6xCoQVmPlXK65bCULA+
bhY5aUEo6CIOK4aQEjx/85jrcjMfZBbLVruk8ENEGSZTh6vqb6SBDIaRrazG8Kc5I5CebJ/yZEE0
DOAD348wWkccYbYpNS0cB1FB6/r6NGAuzM3U2I0pdaxj8oqzpk24nzB9ic7faXfNvvi4frdZbBdQ
SLADQqSF2je5K5NlmQwKTVmHtAF6uY9gJZKPavjXUWJQp2Se3ZuaHMmAUjTkOQnBxT+GF68k7ym2
ozAwvJMGKZc9ZfdWXo+IMxw/tG1x4fGB7NjreX0KWWXVxbR6RHv+xHLsRaZ4hE+M/O8qfTiKQWl6
XJ/dMPh3KBqWkr7QtApcas1ovxt+G7JEA2vz6ygsV9UZjmt7Onu4Nm1bd35/Oa43IlGAdFmxk4zw
QxVBw6wZjNxn3fYI2kpW7JH5u5gwziAzT86aUwI9UMBSQvIXlLYpaHG4qIRqY3yTWRPq5Men0Yew
qdI8pjCL61viIomnJDmY5jTxii/Sucj/vzFlLgCtPRuHKKb/XvlZq2ao1xPVPLuEO8K8IxixaFCb
GsxyiN3peyynZW6cPWEaMsQ1VlZZ1tP2qsGEM2xc1UNFRXPgY8PCk6d9pa9qdmWJj5L6SVZbBbdN
XYoWO2sK7kUOiQmh/OnBmsKkhoj1HGqb+B2fN1oGM/UKGqt8k11d68I+apsG1C5QmB6fJyERYpeo
tGTKKqxmcgiDRC67Ie58uh3jDtpUoNx/OjUEdVYn4jvk4EHSdDz72UpZt5s0DFT5XvXP7sT0N/uU
IY1V5t3cPCKjmi+9f8bTMquIpxqxbldtaP/6jSL8zIdSsoLl/LD5O7dIXnnN1Xq9NYNXMzst3El+
wFN1n6oQP3ZFWK5VBYhu1y/a7KZy5XaxFfDWCrcL+E3q0V+6grBkI6DTclBE09gKgr2Jdym/nlg3
OvPpzgnrqKl98amaDdFUxuxp+0IjsJgLEHZFi1BPJjnHFQaI3fMj+VwoSDU6I7EuaU2gs6l7ZWz5
c46RmVGPPtTwzT9TUXIpmbRGepoVimvtsKopWh/9AGc27mNnih2ISpYtUIZpROR1IQu2KIiL/0ku
Th8T9GTtINTm3nk5iPyz7d0hPT06/5duqufzw+ak9XkWgaFGmBBNOgV5RD9/YjG6cmoAgvqNKukW
CBGugET7cgJBgZc9T0BYilA9Wk8UBlaH/EnbXFAtgbMQ1UVxqmp/I575Ukev9t5lqxS/gHAAEojp
c6yyqXKHiNDRfdjVB/lHRo72k/Rub+mrYuLx7Yx6dSqK3rbD7+jn7na3xUsXnqeweg+UX15cU3S3
dsaDkp87yOPPcHPPy5yRy65QSdPnbLz0qj/CZf6CezMzuhDeMm4NKbcKJwhT2bZKLekyWob8lMtA
KuknY8D6KtfVNJBHkfbtxBF1WlkW3hLY6sw8o67t/ogLf96+73B+LSUvjT1HEFLPYxtwV3P1PLJ2
FmLUdj+hPO5h8Q+F+bu6lfe73l8PGNUSY9/y4M62BUXuvkLVGETHa3j1OtrqSUvptzSOZ7k8dqZ5
w7fEQ/Bo8AvhS39Hv7hB5BG+B86Uz7Tq7UDxWMw1/Fqqa9DH8HVR3xV86NFo7BWBftbjeStc3+8s
eGirtymzh8C7snNw1RUjVmDodngqWsxiKwJCZzngGcn0EY51rHZ3IeuxFugvVkrKfRIfZGGfjTfJ
qLfz+exMjBGlg8YjCfjDcuLRmGnGBu8b+TmZ7N1kDD5Amfs5hUOuPg/sDQfcHMm8UI4iu/YZpmuc
ARRfR19bbJD/kd/MeDxVUwameoyZUX2kG8hbBndPk+hUQnW0CvcKtvZ5eC7RzeIx2X0bUQVbsQQr
WvUtOz1fD/MNZzqYNUUxu57yOexj1SGTFhzK0vuCmQD+6e0WpZ3zRuUZYUz1yL3w67Cn/3q5gt0l
6NIQWP8m/YNoUYC22sRCSP6oVgR9NZGiQdE2V01b4vkkjgcpQZI7ePoMqMTO6HVKlC6jtIenni18
xoXeIPT7/Y+MfxhW67GmfcRTE1eF0As7RwxFEvmLIkYbFDheLz6UbAijseMNJR9JBCXlUGr7DGtZ
MXY3zXq1LuPAb57r4ZQnp7z6a8FKb02WVjsjeIqBADv4TUU+qnUfOf8ADXVDcxpot1/ZD2h0Ri/0
k4kBcCgoB0z1kPfzNBQVEzAjSgEjGCfBvzwIrWyCxFGvSVOVc83zE11BajLcf3Eb90fGTc+w+9NZ
ZzaptlWMNP1pLf7fFC2GpQccRC7mDaGk9HAkflCZzQ/Kt+00FQ9Wz/ea/P9eUvzUF/Owo2Krk/Al
mWfp7fqxuIqTrq1ckmFB33hY4GdGM1P9rST1w23UkjrzaF8tN8maIn0XItN6twuq6vY6si7md4mD
5fe0blCwXUIgonIMm/E4PCOUfmXWVsJP4xL4iKPhfeJLM3vmi0lppaiAuAA1tPJ7g9buafXMDI5j
qN7xrWAk3TEU1nMFVxIyM+uhunZceoOYcz0r9oE+t4f8NfbCOY5fIf3Tbw+rOxtQL7805CPzpPBH
0keb4GSUQQ3wldInYfJnAszl4t/sMYYJCMYSA/Rhn/h/7uGW1MDgz3S1mZ5De7bQB4B6Bh2VfwWf
hsAtPgd+NtckGa13eAw/sJ3B+8xgwXRl9JHmiSNQiLfAznWc/OZLdOPiorx1hHk93W+T6xNpG3Cg
JTSL/W3JZa/dxStKvRoDuxOZkcvF2+pkLBhxtBzsX0YLRepzGQsm6KeJkRkiDtjTiC0Bw3b6WlFf
5SVj58VKbxBRCZKNc0xPHCXZXnERzNldVSjO9bYEfOKWt/y+t3nraCyFTKz5wN/+YTJzRtiytafC
X54KUt7yemw4F1UzvS9cf866bxntgG4gC3av+hbb+bt1NsUG+Gngj/NiGMH/hmCz+w2Q3sYBajww
5FpdEseaHokiipNjdcDZQIRX5Adh9JHAQcY3Rex2efgLOs27ZWqqqBmzWVLfwQPykmeKZ5p/PGr+
5TeMUg8b4+7xS/5r08vcFGqaDSf8seXViHss+pLcxFDqiaKpof5xnoaZIEj+DC1zJ+03NTV3MyQt
yOMV9f/6C7JwSZhL0p+SqgWA99UocIXabhP0EO4HbOKxpI3F9oykniL/ij0CXd7KSCffJY4nDUCF
nJyNCYPeIp2k15yQh7SlgFVnsC/aNUg2AlqG6xEMREZT6SeLB1dUzjm1TZE2TVG5uvcFWrjiZNSl
mNfwzXfJnH8Fv9Obj4OmfYwb2YAdE3T08o+ty1knIaq/wjGlYOE6nfqQhFORQfz4JqWTjqBqSwVM
SdFpxvkuUeKiaDpWLiKI/pdwbkWdUqxfn8WVwF8pJx6zrEmbPYSKouFXEzScf3CNpMTmzaAoFjRq
+yvL+znCTE08klm5oH4trEQ6rLczmIO59SPbLH6XRVQfFnM99PQ+kLBmkDvpwWuzz0NBoXZFsPbF
GZ8bYtAFer8Ck36s9cE4dcentluS5Nd2+bU7g0rIW04WWSytSdTuB9DYkJss/68FyNUK8X1siM3h
UMGeKbNNmJjCIfpPDoH3uk9TjbnACs//Y9Z+ppxScnKSKyRJ5S9GcLosmvT2dCteJmvwiQdU5L53
/nXu0pD1SKnE0s1AoYLY6oQP5X/M7+tlKbO02rHLGiPywfqa64bip6Cobo0MVfWrmBPQIMtKamHl
i1d9+hfjdQkLPdT1pVr6IcKWRfJ8znfftJaUzDNC2b6GLbXbunBN+oipyTDQ8eoremgeHrJrhe1n
iGerrT+TzP2mIUpL7R1pUjfQi4h9PsbZqDiU+X+UYeEIXXZrk13vUmTj2y48aU28BluPl9mpaTyZ
aUXMWl0/6+yNGx/JI9SgTn9sPKc45GKoseoQVDjf/e/Nce/coPjrI7wBjbwL4J19iqt/2PJIqdR7
QgiAq7K9dgWxVS25JDjiyebXTE6RO68HxhgJg24Fb8Bx2arJaS9CyZIJ1TC8byQ6rDsngXkuUdxr
+33opIsd4hHV30LxMysYg6ewY1QXeaqm99PfV3KSPMgDHUDTlZeiGafYGC6FV4uBpKwB4LFYsFC9
xcigjUAo90kzIGl4UR91YEL7KT1YHdpFNfTRpOcq1n7Dkx3yY+evTSwIhLgVOMPIJ/UhDd0Ac5M3
pz5NQZSvdWQ4WH8YHO/68GZviterQmXkf734dbTju8boCMzWe46WAaXMm8RszB21F0D5loVQRfYA
UDXsb/GDsGfdOBpG/PqVS7Fy/E26HSmmRSobrVbgcvfj+hxLiN2TseFSb5x+5ZG77jW2tWuQk+N7
P+Ck8abix4uQYK8A2MCLoZtWh9c5jGIFgcwM3DtFxwIydjF7uA+yKkvQ8orHPoS3C/UyhFv0+/q6
+CB+K6Tp1+75giZWVmVqJJ3PmWtuoO35cYzKHQgsfzv5bABTyIaCMC8Upxs13xEiLWqEBwqmuPOd
IcHhtQe7CBJTCmDQIjLUt+G2xG9y0wBbPgbKbBt3IB9lKtatcqX7f8bWv+pxpuAtEva/lpLDgKo6
3Jknlu/Rk1lsedsJqg+M/lgvjxKenKZ54L/LnV0zF3LJ0NIi08P9XYmfAmQ0TgVLtUuHq87i3VaQ
iZ2fgA+DhCFkyA4rNDQuhB0BmD2mU7UiU9AAZveLvOMDWztmPMU2Q3bfeRUdHmLIFz9W/yKUwPGt
DPYEeyXISt4XaTyUcH66uvsQmc7soQGsXccHdqSqpoONJNPIMG/JbMNecHcusjOkqEF5UK6VMQ63
c5OyY4+6HSkCroy3Ss7f1MNQTi2A476gyP6Ub3ZVCOEq/UnY1A9ANRVb84AacFfslKexnCWlruS2
0IUKKgcUnPyIDjV8Gi2giY/Gl9nNWLZYjT40eyHCcHdjjV7dYSi/Yno/9pgCnH6LLV+k1jerlkWl
oL+GYXd6CEXgMntCe6g9fOs5fCruv3fGOs4sQ1W28Af0YAMODwCmNkcxF7A1zOkL2x6vyi/6GSlq
4Fbrxos7/Sy++xrw5PtJB7btSHC3Vh1JHbicna2pXb9BBRQhTuA8JGko/ovveSKQr/WoBpdJpfDx
17gNovp9Kyba9iN1h6ZoHcikgv6q5dZWGjRHFgOXBggCREjGLEEeWX7cEqXoI7+AMIR5EynNTcQZ
aC5or4Xjk17sLgPldJ5SCTXk1iwjE1sNe5j6c8p9RO4xEluU0GN8ENvDmzbzNejwV5M9PiqFe7um
sc5NgDDe4I9eul6c0pFldFY7i5WNDXaHUFAJxV8g6qUY051exBEYWbp89C67ryvYHgyfI9rfjrRq
zMyqT0YC2yZbxEe6fVdU/4vIVbVojxNMaMffgrkTtj17lR38gu5RiWfgzH0IxDMTnFt5uBWytIn/
6PcVcb10FpQiKWSmCuwx+4EJiwI+CnLY20ASGqSggQZVG46PteEpYvjWtlqMsi//LxDPcXs8nA52
XbeS4B4zQJSrCLcQkxpZMl+ZPDPNAw0b9pe+K9zpypCKs0Xqqv5D3H2y4yWQ1y5TQ32eFkKbY4yM
V+MUWvfPsW5ASTKV782i6WMD4iQGRfBfte6JUIY5Nnw678HIwPLQZRYE0oTXlEx95Z1hBSbH1qjn
cSC2Cc0xXc6Uch6lgJlWGUfl8aefimI0XHq6yBuq1NzZZyB+jdpG6S4st4zrAExfv0gx1queTLGP
2ErYSVVIIgmRu9WXF323rEHq1JABktdhnkTiBUL8LH9wd4fHNOPq/f4CdrDd4VIM7bkZWgpETwAW
nfR5QKCHSyWqaLmyR67zVpWjFAVFaJ7yEIC79riGIFWhT6zFh3ZyCcXrwCsZJIESnHIjDiXoQuOY
8qnmemQIWiT0vzCLjL+y+W/IE89Vd0e+bLMTudR62SSkMY4CMlKlfKPIieWqJxN2BAOqtg3pu0Nm
gGUK37/ZLBoXV1Wvn1hAEw4tXyMGCBivBHTg8nMAjfOsZD7raUR2hNFnkLGUi0WmWpE11KUql7BB
lhmNLWa8ZkerRDvHlVf5aGNEElv/mK7uFnQhSgVfn6m8FzJ6dhhZzKNlpoLMtdsP17jLaxyStqvB
v5Y/KhV0xOq9ajfPT6Zz1neFnvfep8F4IpsjnRS+dCbxEWFrpryUPtGB9jCmFrCy54m2+nrx0JQ6
LPciOXHPmy9azyUpGTcbTkHZxOBR1DsbqQC83ULkj43DJMSieD1rZ6mhKy3oJZi6IHIxRaJaOavy
47as92CFdACVEdfEWiF8n+BOwqZXcXmbPKp3FQnPXdaDqPGjdQAyRttYE2HFmRQXWOhoMNX/c4UC
kwyvB3f4UQGRCqG8BEpirB+Z6eOiallKYVFmILE6Il0lz7Oz3EEFdsReAlX8ES4274H2PHBqBs+k
bPJ16Gf8zZQ2iqu75skPVLshWqNqwz57E3ey3FKGAv4lr/sbvYyZ4zGOy+IAMLKCVEcM5tTNf8X3
1qVfTPcU6w+MuVEV5NEOWcatBB1LHhSjfB0hiSdGJ56YMoqVEpXWU0l64UIYNNcQCTAsdy7/zIab
9ghOw7IO22niU6vJP1NHDMupf8yQMswMAWGcj7jP7/QKVdpZy3gi1S1OiRoY92Ia/fyDnMfYY3kj
NBKgDx7r+jgBodC1Ctfsa1nlJcxKYcE0lSr0vu0mEQxKEctiWXAI31aMlmg3W6vHVzsOFfqvinSx
Iw8rZOvPYImWWaNjN7N7CB9bZafqFuMxIVZpWKvmzVMvYW9hBNXW1R9NcQY4YpObSbESSeAOYM9o
ESgQTHifDEOCSSknoRy9EhnjrYXNwIyqZ189w+4wC/igyMGwsWJ6n4isawZHyrgAAsjM/FKkAJJV
NesQvmsPI/LjWAzl5xFyzAgPtoT36uxROA+UoRDKD48VvkZfuzqhmCYcEbXvUH8sNWOPP9DBRe+m
I946YWAf/KQKYTR9/qWIw0obVpgJfTGDajHvdY68SV7dGIfVhfTuBmkslP8Mon58bW2vJdGwLbZi
HRKBfGKWbwgmt/TgNvEwC2SNIPCtcKfJttntoyoK0fRqUuQ4n1Vtudm/UZUmdSdUpHxK0mLbE4S0
ByjkI5HkwSy9hAK5Az90iD9Y5R/j4vacigS1FBWVKJme41A/Bl7znX8vDlJ8MHbIHA5MDWWywBae
dbZBEcV1w6bVCDNAtJtRXltsbPAuuQdhqsjC2AhTa9HRnrkhnHSY56secJqYnahnH7t6RrPWQMrm
dGvSm/H5LEvDPHm7KmJXiJZligaLU28ugeL7B/VJqmSmabLE3JZxjDYdJkqgRWNcnMimWi/+FaBC
/SrK/wW/tKe2Vzw3D6X9HIfgzJ+dSK0CRYtbucOxgAA/oMtYN3Fi/MTVIXsOLQeLKZRXuSzo8+sf
kUs/jkeQHzSgN5qJ6KF9p+UFh4KVXeetFtmANqStWBq9SGn2iXLJeOwLOb4WZJ3J0jmo8w9XgBri
L9Zk2/4bdPMI2ugVmU/ZOCOTdRv3NSx5cQHMXlbI70DGsxevJ97xIWokspu6jRXItsCbz3JQdt/H
ZGw60x4Ka5VHKUzasdddJwCnzKM4ZDaC6E4Ji3Y+711X/BBX78x6E5zBMMtaWeq05QS9p9YK3UBd
1bUR8t0rssLVDOTvuqDLMvoLGjbKxEkjHqb+zu5YEb3b75FDqbnYG6ajHTMb2rOTCOKbq8Vh+Ckt
ly+02GuqVrQc+hpOWsquQqsYTkXzcE0mJEkEBEiP6VrYrpREomyNtXleMdc1IIgZYcK9hG56a8LO
2XkdwwiVD+lSxLk1dMy9Yn9aahH0jN6HAS9VuuCW1jlN84jS1rgD5OdIeRNwteFxBWeGXQ5t2l28
T/A35ZOHUomn8XFQPtcTrdM1sfx2YcD2a6Q2G/zpxvxZFHc1FkM6Ytisifb9za6LiDmi/CSB8KEG
Ok3srhHo0DPiR7+Pu87+HGPkMo6vLTty+K1swefsQV1A6yfhEjCbc82SernzzpKJPJ20FCvldMHq
W+nTsoelNbq4APRKcnEePGy1ri+C+cmT+pnPbHCevX6xoAStPZjkboMHDxJqfBp0XJ2L31JYXAxr
ripGUcHfV91PfMl7K8WGJpFPZmJ3eyJRdQTdN2JC3yIn84vax88bw1Ekor0sMfWeOpqQgaRw0lEf
3NtENO4xge1x5Plw1RvgL/R+htK5cYaF2YFHyqvPz7II12eOwg/niynMSlIclDEc3i4QqV/HezyK
C1mezHDpyxsoC6hjA3RfiocTmpnnFGOUfKB0vwY/W1NW5VAdr08WU6+CurRC5rsIksgQmGrfn9mr
GVxPkZc8lIYIcqUuvkIA5HAcEYWK9zyZCTj/E2cnZc7vjB4ZZFi8iLkAXIZcnjzzba08pJNPmNlM
hwdsTFxQKEKHUAwN4OdT0w4Zfn1Dj9+pj6ctEcD2JiomryloZglKPumj2kIUO755gll2dnqzdRwo
K6AQEg1GVcOOtu71Jnpxhjz4ASGCOjQpViOfqKxjYPWlWV4b7Hy6RNVuuCZgBEfy+s5NGHuWN7e5
lbWWW/DUqJCkTQ2pH3H/gprGIlV4eMWBS+VkwJ/9dE7/+ZoD3A8wp1O+MflcOtpvzmgbhktS5IYy
18K1Qfjzp9/vCfAfFVRGi4Nz6KdEVXTYkamhUYlwGg1C6VWradHhf3E799++zNEZUZYz1VWcueMI
hP0DbITS/yY3aVwsjUWIcbZouh4bbedBDzHfqWKJ0BYTpjTEvdccdl0ZNTEIVLfCnF8z2PKfYWe9
41ZtUIrZbTgThq8kVAql+CWZS+vdz3KtvhIzp13QHAONrB/MQ1KoeQxfGaNNyzSGjwlYtgCSMWd1
BiKrBzfA/uH0vLZfxjwDjwYooHzDhaE07y1t4g0LdPEdkAvFFZuzGZFR5WA0M3ruyTWNRy2xtLaV
ZkOrGBlqObFcnhCBLxpHIvLtQvMaOZCbNSmfd1vxAUDm8GjAHZTSoQufS3sgcue3k9WmbHEdXSwX
VwI1pMOsjVcYiOcfaFO5MWWK6pN6o5u/K+SETL0Z+dbekTi5DXMT8IHw08rc9CtTWc1CuM+S4Uut
JnMuG8n+Qy9sVxJ9NilMTDOG8UOdUr1s8QDWK7SYb4Ua/GMv0DU/HxC1QWgF9Y5sj2oBrinFw/Us
G+zn6kyqG1SfX873zYgPuvuxpsTuQrVqitpuTSoBOdndW3qoxGc0SuhTyypMuNcPuMNaNRRAnIEw
xP0Nhvt6YBXt2ZMsQX0GlUMW083VztADOlTc3JJiOf5QW0lzcPyteQazTj4z2DHYVA1nU3o3UvrS
MCmYAGPy7xThtJIyuddwNRW4rlpgn7h29NNjVaeFQxYIpDDTSY6mebm9IzI+5Y89/+b0O7nuA5Yz
/p8jpEfrwQWOQpHzJnFI7rSYSCO4472Vm1UdauOx/VKwJ9IRpBhoyFvbVLh91k/GQ0vBUBBHyQlm
ClntYlILEHZsJ+QHvsp89UOw4GhJliN+zBMGWc5x+P5naFC/8yrklmDA6th/FDLNGi6cB8fY/r3h
Vk+Q1HThvWVqNKHHEe6u56Kpj4eQjohk8s8rFMeDu+jAUG6kZ8gtp7meUCBmlS5LRBwJkSDbw3VC
CL8lJWL4ImwZ+2UsSIKzzbHeiRudeA7vomYgjpIQtWFSd8JwAWj9JP3vGsKvxjirUiwcfRx6XQT+
pANu67i1WstetYvhe+rNIhzLv6OEvcYSXkzwhG1baem/7YT394PgE77ooNOP04bD7NYiLGteUj8l
493Pwmz7Jl1s9HJ/SUxlSeie42CVZ26tPLEj2ZbSA9ilWLxZpUKvMqqzsX1rcAW3l+dy4LS7CXpN
gO4sud8DBqHmPUbFYrTB3NXH5y+tJcj4vqDSDzMDf5HULMo6QDqDqSqGG5UAJoBd/k8PYDUO152x
yVaR58pJFkQpMejEZKXN+Yd+PZxHVOVDRDkRo9As4rNwJVT5W73DDb8tTml99bczNTDJoxYznFoK
FTtrXkZmxkyiNS2egJWFldaLeZr7sLl1uRKw8WJpw4TfoiiP28PXO/Zpb7cVJyJm/RxBpnP7DPM4
PW3W7kqQA31K6hXEys4IDleTJN5BB/p4CzmQwSE+kSEOyeOvqIUTdUsACI9pi+g5NRmU7pBQDPvc
1smEh9TwmQEid4HoSdNNfr1U8bdUCNAFhOmmXsISsF1siFhFiGxne7ldBzsUM2CvaB36k/E0lqT/
PsbYOS0vbndXFBOEt7LQWSckALiNGwu7Bhuuf3ljoiUY/T1MbwSpAgeNIolSOIY/7uc5XPt7E9Un
vyFYt3cX9yU91nVUPHO1SaHQ6NnKQOVcdWz6p372y/yY7aLt8w3utmHtaI8kQvLZI9gXVvYdA7hc
fl0Ia/AzYP4ovjXb7pmqYR1C3vynRqREGi9Qa90xwNJrttVMCF3QHE+9q4uKkYFO7TTWhCLxJ+v1
0s3H8rdhLrJATJY2TyW5oSou4iXStKmZNKJvcgDLR2x2GaaPhIlRQQFSpH2EmEIn43wO/jQdGE6g
rdYnC4+o2tCf1TQlp4wgFBAt9CHZlAf+CtDDQdJrYUmWqa8DO0MLABGaFbv4wqTM2q6L72dxCNB9
pulNNf50TTC4AUdOCJZl3jDAEa+hKLjnyGRzvWb5l6Ena15dLVJHcjMm4r/X/cK1UPCOBdrgadov
wSvOmGcjNB+u1vkiCgEkSOGKEq5hCYuZ261BmuKtFeOzLHTLGyNTM5Hwin6A8TXZjKHyE16XHiKX
OIiuaKAx4ycYqJj/wJA8nKH25ZGKnOw9P6g8VmgOt1xFwKq7yaEuLPLMfiJG4elFx7VPz0kjqEqb
bD38oSSnHA4Y5dTRXDw7lcYGN99F9NGzItLV83a3EQwSVD65jZZfenc9XL2AQ7qCKbcqKs3i3SgU
YL9nU6RBaxgnAeM+Yg1OdI5FUd9F/FBOwEoiq3rUENTsGSMgeSAFBq70qD7vUiRJuc0QmxRDLf3/
Ez329O1XIV2ggD+CUVEk2zXc0Rb9jKNGsUUE8o1TA1pFa6XxUqwXxLh0Tp04Bf5DkGYCOtX+rJVv
/gmAYSSwflmvfF+hSeNJhOGRrxw9AbutyAkMq2uil1w6J2S8qcr0AJTtj283PDTgdxFSXGkZ0M0A
Mg60GWjmqnFwbM+kvYCKpGzPskT5uHjwiZGNeH+bq4zEp2yRq2okzE/9EdcFmMqPT15Twtbt7Fea
qCAICy84JyAoFasEubjYi6lE1NIOIrSxnPyWfpb5Nb2s9rVmE78c1rkhtHb/KabCxowEyyEiwhRk
O73FYc4oy+yzfI2jVm3JVOTmy+FN2BRTiC5i8trEHqcQ1GyDiUbTCHlJY8dmk0ZqvP9GcyZABhHo
33AyAQ9sES1HvKOJwkl2WKbxsCtnw60nHVyZx2xC+1DEaH+SeQfxaRYPyKmECnaHRlacRnpOfrR3
sg44aYyUwoGd6LAlSaGOshYWPw8TUzVslUFiPfKEgCItVHA9ynvB6Luqo8UpSYm6nm3Cg6nPm6V3
zmGsjH0OHApDgFhKZG9i6J3Md4Yk03Kt8FtuC+DiuBivWftHcaDnk3CZo2rGH9dZeOGbMmUNig/p
K44d/YvpUicctMEUsCWWclYjLTL8Axom7bsjd8lEcXMx0TUqrBkdAOgvbJ4nKpkZr1u9MO2Vhrux
OxIMyEM9LfkXAh1ssvZJ8VMVBot9+LvDo0dwwnzoWh0j4pn31dYVHIehR/fpCqRr/kv9vI26oeC+
ZBeikBe9gv5wyzFn8/teY/Ve4nL/d3lDYzwQCD2jBQy9HwdMEuPoWFEe4qMvvnjC64/LGfMZnEhE
XZMpvkxA2FrjjySzJlJhneqLt+m5iJdCzXgCWM+Ov4Z94xSrtFDTMK57FtL/EBh7MHd6/GmPKiOL
E2DQrqPuRjPOCpUnYdqNKUvAIMgs3Kx1+gdhvwMzIdx3xtcfRbnDCL4mXnDaSGFL16/asO3h5xSn
5beE0aaBFVa6Tqcyanv27eYxr6eHdXfdWBN39uYziJVAxDRkzw8yG6AzfWlY1YLCfSF4vxr7PSNw
J3Xiflg0BmPLHInAB1x5586cLhQ5Oatwoc4yeAisu126fUriCSDVrHGjBZpn3yGIZR0JOhs/WxGx
nQ6AOxigcr3P2S/k+Bd4cBb6bcKbP4adjoTjLkMz2EolemiO/46STKdH8eH2QksF+FzYEHw2KL0G
LBJCMoql2wCXOBY6h+Sxa1N8B6nEuZ6lr1CDlhXZfJZwTBF5J1PqcGLMHDHGvi+QngIZJh//epzG
Kjt0QqOlqeD+Yx+W15ytDtDqN+8sItzZ+VAHGxgFGB9mqBxTGTBSYr/MMrgdAg2ao5GEwrbWrhbR
LXwGF7BzEjrAD1QUVW9I1r887eAUrznHmjoVxpPmrDgpCgDluYFvX/VI+S0xajZjp3w/iTcJxw9D
XapB623Aft7oL+Uu3KHxg20GnyqeTa1bofatTraMX6I4FweqmfisG/I+704TMde4l842ML21FGwp
BIqMY9oa8+g6C6fX97H9NQQ9sLr4xzpM0eJMihaEc0wYx7/dK7tOP/YfgXl2NKtPsKnFXxksr97Y
Av7Ub9Ppel5WYiXITMhJwG8KLfKQCI4CUL0PVMBRS66iqFLQn9oNtBuCYKP0ydLH5zdcGkjhFBny
0yH5r0mdnTqdoBQWWyiPdyDIV1B4fePtDvXGbEk4eR+MEoaSDy49VKCVdoIcwqqDM2mhJ0Cn5Srl
jmzSptSKcSqsfHvqjBVC90lIT7+eprRiQbUEJJmVgpHpYvCvyJHJlD/PTbF94+fwBzFdvQuBhAdT
/pqoWY8nju29/7fs/ry0RSXutSmIGP4xeyMp39pl0WB59JqIfC64yQwoPuMsKaorS2xcXu3FLn1K
V3xxkXHz+VFUch9QNQp4kAtEg6OfaAkmLgqlRrn70Z7bNafoCyQAdm/r+jz+MGeOcAuTWbK4Oh/x
/VOROzBxKd5smZNiofH/6T9amAQ79j5oVcwSU+cvIGSpVghPtdb68cylLiTFtW1dXyGCGiJGAlly
uNXP6X7obRvJsbWA0/NhfO7UBuKW27h/IeAbm7wuhfwJ6wrhThA5++/ZsrgeMc/7f/D3ZXu9Ho42
AWwKUFtKsVWHqD+OlgM1q7Y3WJipsORXq0wuyfZwlgK7cjfwqwYb6qgFPugAXWtYE7uRetqN7Soa
YO6T4mdeTdEidF3oeMX5q0YjJTCTqZxfgL1/FOz6ZRDHSigLH9AlwUgfEkL73XWP+FXovccEPnpY
JdY/qVBInNae3Ar0tJAoqQLMZSh2xp3X18NfXi1L8Ue3M6ZHX/EyO3MSpUstEJa7wB5+EnfJ4O45
YD7yuxHN3dkMsfffzSRwc9WG/3vmCSQwcn4v1ikWV9pABgog30A3UcbL04prnsSkvvvyh4mZJC9c
V3Uv0IRiaLvPALjm9yva2C/r1acM8SBQiFVOl8Wnw9QTNt2rMt3Sc9EPTD9w0zi2UVVYFtvewIhg
w27SzjJEN0cJZcmiuu/KKyHDcwOko8YNJ9MPV3aJWqa62E7z1h0727rSAuSUWtNeWTb9O26OB8Wm
eRijj3WlFnD9JImv0+dObfiGADLp3FWkPe6Z92k+/UefJfmHoiMBGWUixfMvUQi0mqomMZulXXST
0q/50I0anXpk9jzJ5WDOSofMOi+5OHdU3kMK7H42mkgKwrf+vM/04Bd9ollJuG7Y2qUs65dkXpaF
hMv8xjWPS6X+xPoYHNFDEQ7cqCt3Rf/gqdtoYsfFfxrDCXW44RcvfHtOZMwNbcwZkkbpWS1HDUwr
K/KoTlBKLv20/cZQSq/sBFi7Y37cWjmrguCrkpybjfBqj5yyNodY25kTWAJidOd+ErnlfbL6TXZo
GlEgZRBgee/pLI9QgB1HgzX4lwWaUjJDOeHRVesNiEFUZa8gDbtucSmz1Wm8oBzTDVd4s9xuLsvt
ZJegWrCZCkSJaGqLmG1M3+tmnqx+gBK1jnWQQDdeqPf34oEhryJFTGnP0u3T3EEC2XqBaN1JJEhi
QCoiq78X3HhYVOm21Fb1HXVcdC8jmpR8o0V6t+9kQt8p6fcWJnTMuv8mTT+eujs2hhO3WkOFNKk9
77JPVkdX9f+Tl/whbq2aeOe6sKIdwP4GBM1OLJmsCRN/D97hNHIXFLGFbOnjhVd09KHWQ9lyPuQT
X54x/oIUEXw2x75h7af5AeZedkY5LLrEKwaq8gXGLZngxelRHNsvQ4NAd4ECDb/i/6Gc0aR4wJRg
x3/bzWN/v/TnlvqDq08UC184A1m/tKUr1PHKIFHIj1+InUypmJkcVn+hz2TwUhWGMnz2CBK7b7jR
khfHPKSm/TiPGACazVWnX+iru9ZbT+ZNA90/Y8v4iSDjssOm6ybZnVnBFsFL3VbuB0DFUgyo8Wzf
TxewfMyVnmZE5yWDtzWZMJV6FH8Bt9rdZ5telQqW6GMZL9vvQqxW62RQCRF738uZKJs3akerb7oq
lyI81B9BurH6XNTIUrl5xXEVi8FrJvhJ+49ptNEcHmUA2wiYLAKqLcSq0yhOsoA4RZ2TAefzNAUh
K58ateaO7Y1ibT0adWp4wVZ/i+DnzfjkoaLuDzMpfbypUow2jWwAnG3gQQzx6G5a6rxvHwF26cTo
a41fhLAP4vAiNbNfKmWAVzXRfgEIu8mY3D1dwmjWW75RNhiuzyOpDEkrSXL+O7Xp2rISRUFNgIiK
n8Ri9JKf7AXNTehLSij8kOVQ0KssZ3s7Ntztjrqv/z/bgVtTgQRnJfB6EVuo/5lmxEFdt5NWlUAY
Ai3cU5ONBrLuT7xr8YRJyZEnYxDMMiTeCKT9c5JTWeodK8dNQBACoSTWOtljz7c5iL/YrO0ri5U+
qII1qpSqCZzBFWIdSynV2G8Ff/p8Z/j9eSEtdCuK9A0T0v7w5q0BKlnpIXGnfUv85dahzLPv0fqQ
X5Px7AjZBYg8tfz0ts1VDKeDQcHAgPNT4K8AquGoJuFhkNd3jHiLhTskcU7G13bBcBdrodO71TRk
8zr4z2AAa5u0tT9wrO3OlU98BdWLtsbfcZxocrGVu3/1pOzq5RZ9Wewp4EYscAWvR79TTsZc1/sE
0mKEsPkMCir+pZmaKN00sIS+1ZKnOCPVa2D1fpaaB8zIdCXAs4zdUwc6xwcOu8DuTqlQAIF2fsop
vQn2dRCDF/ihw2RkFAejxPQy7jAA7f3vCyuzknFntqFld/oQEKiRY2a/tfbfmkTT2dFkbwS0s2k9
9hZ6aefYTk0iaGY6J2Ag0XDFfnW3XlnJgwnBZ6HvIAQynTX9NVbzjmb3R6DQhff3Ja0vwjfsBfpy
vj3edoU0wpBmpsGaCaaPNpMC58cLqRwHOpdYy7Y36Ns3R4UERsLfeoL0A0nq56EhCcIUMTqIj3tD
Una2A63MxOIXw9Kyct0yOuZ/OeIQLs4hbhcNf/lwMV3HmCejSN9A/K4S8HUiLU64rO5twC1CCFw3
0/XLzFzUaPkYu+lSWrY5UwAhG9VyD2TM6CM5teQ/Ss3XfcGEAr/BgfDBk3nHeZ5RPHtIrW51lGK6
0ITj3KK4XYobh+DIAbs3jLBq8o09nvVEEyDkkQP9i7DRseNyd9FKPxyQr+P3Wu3e1+9gp7XbC1ae
OofWNsvumEzSl+L915/5Jad47rUdt5DZacPaRkaDsNlfQ4ec2KreLgZf451Ny85V4hTk3SoCxOwK
CX+4Kcjl/mCtkFRtga7JVvAm8uhRTqpjG6lYtC9+Y/UEMBMVu11Uz0nru4BP+jl89eHa3pzPOyM5
xCn75lhnrvgNPUdsQJt/KYFgcSTxcbtHkoTZHTtBNr/yTf1+EeJ15LOuLXRCBLl9TBs9Z/HbqSQh
olNEIb71dL/35SifyJtULHG0PWpetQx0fwKedWDFiImw2qdYf2Sxh+kCNrCxch01H4H1m9VBejSx
kKEhYWpcXNgDKB6Nan6Wfdol3UA3yEQOVJdnRwNuMxcrWdpoHbBnded6aIueppS4pvaq3CnvI4Yh
ZC6ycOTuRUiT+KFEZ12V/kPVEYaC/HBofwwrwBfIu375KJBoYxm1ZoP+0N+7Bpe6+PaAjfI88uEi
TLMfC+YeXwnDa5j18uOJ2+bXEVwEYWKU/wRU+9QD3VCD1CJLsaPoT7nr3hcK2ZeMhBMjnpGHayFH
Wp2JkaIQQ2InlFKfM554TnOtBkV3kOMqWvT3eQhtqxU7IyXNk+BlF1RuEx5roukGG7lw8sJMMTab
J48iuPL+NJJ3frLaEoH7I+odb97Bx3XHkAo/uHqIC5UES/yoMj8xh5bZCLNJuAmoeFroJo+la4ol
3WbiMlCSYpxXIbZlRa2vsE7/7Gz/gYxt/wu8mzyOEC67SmTTt1uJ2BKw3TmstuEzUvNeistns1vm
vCcmNzyv8UZokq2rLx104XRgSdz/VsIa/uOROj/R4V45xlOgEwY//Tx7vl0WOBP3ef96ftcht6bD
IqkFJblvDCBKqVL/G69/aH3OVe1CxXbT0VSayRvk1nxrjnfQe0TO6JBj1wkcADR0zy/L36Qamrz6
HKSnMMNaaYmG1MLYH9WFWmfMxBYt0TPp65d/MGnbGxmHDcjsNJtyzNpRbjSQz244UIx3h4S/ZpfJ
KDD8v2iRNdAZBa7ycw4q6EWQD2qIaMpGytklm5jI/H6LqXf05aoRI6j+Vy5y46hnNC1QDEAyCkbW
LLERXcUHAUfTJLZJju5ukGgFk58gP9/2YOLk0EOhqqQ2+X/XvBKJ2APyHpi/cav6hyDQvODBjJin
2hOmiHb7Ah2xb6t+qZdBPCauwBalckVGV5nT9M7MWyum+FDYEWU8E8TLFmnWHkXc6Sm9oQKEpzkj
u+TWw/LZ3VQdP6/XAs2HtOzcrX1RyZDxhkyFdolxd1+9IYH4Aag1sF+ZNkWGTppY9RyVAoJNFcxI
Eny2Q8dbwEUuzyRLxRiDNC9qF48LHT4J6v3AKLDQtyk9Ou5VXVN2IJZ9zraHvOosVpHyAhu3jyh1
5ZwHTxjK6c1jpi0kY7SN/P1Wefoxn3wsN7r1O2dWCSntd6k/hGdyZieXhI7UDpWkvcSef/BM7Zc+
17AJgcdONDz0uDizu687sEfEegxoO6GgPOjTMaWZ0NZXRv3C83sSTrThe0GuVPztGQbV2Yd0VudP
TmSAxk6mPxkK2x5KkcqDpZ9XHKJAlBlqlQGvvw8RL4Y/93Zir2s/YP8kAUcC38glet/GIpGaAsVZ
GckTAjbiUY8hK78yVQkV6hFKKuak4ELhpPayvlEcoCYx16RciZyy6iKJ6znHcvFRFkt8fSSr6mGI
0uz/M7JWnbMLsnM2SNcvN9+zYyMF1R9nBLce5OIdweeG2qI+26as6GKL3dkHj3b28rVoezTrA0fJ
uxh4G3l0gMBbjKKybGRHJpCQ9C5uQMFLNmF8GrmB9rqk47whUM46k2fedBQ2jdXlUoZR9m39yx/A
rndYjwIltKbalPqb05LfSSZxfNhcQqZLrIMRXWWQVzY5Yf6kjtS49XnwXOQ27RSbri1LBKB3/pCg
D55dRo2CBzKKQoFcx3cfbeF3GwHZ4YfX7CPm/SzKxEikCUMpoe6RmAV+f75ShGEvRroKNCnsVW+0
hR8IJnwzzVE9ue5ZAaF+MsfM7iuTgEFti60YpTTOtdb2CjPuU+iio8Lro4Edy7G6F52FMfoh0aDL
opiyHtkY2DuIa7hP52IYuGSxPz2yXEX+HGqwGpia2BjGklNoSwOH/iOw/s8X4lf+/z9+4op96zAP
OqUk7fJzlwfqC/zF3lEZvP++0zQ7bnot1G+yk5w8ANzSOjdO+HK2/GcAfCaC1p5dhFYxCdm7JOMU
WdXR0CzD7o0dvA9ARZvrO/Ln69j278SGwlk6u5TAuRvVCcrpz+kK/YoDNNE3aRklYBDMxQ75lfvX
YXKyBhexnPTLNaE3nBANbotmU8xQCHYsAXNZrwlcB0STBiHzDoDNoe3DO+mPI8Oi7femoIpYYDXp
XzlyaEcosvELS0bLifJgdSgo6ih/67ozQaIMQ02SxrLtKmR0Q0XSnDwyoc1beF0yPguL3ZTRNpLQ
cp/SAb5vvXtJmB9Y2wxYg7b8ezzRJeRSOnmjoFW54oDPiU1NI3jrlQNAhpV2arZYEFgDpXStDWtz
Nn+4DC76nUs3QivbZ3A8XziO7dU8z57Je71dMj6Mq128mfyi/jWffvOeFLZm2DQ//Rj5GkT6r3G1
3K7mEdZacMkrTZ99eA2g/cqy4+wpTJiHNmYTGfqDAefvuHNsQwBhPxw8CjvaWCXbjnm0ejkGl2Uk
EIub5NNsyeRdbjTo0orWtbtGwNCD2n1kE2UJEwFqIq6naEgizEl8rFIyl/SEQiZtsr6bRsHM94Qk
cq54qiizLKOZjUX3WvQV9oiD9pyDHAjouHXbOYKBDrIp3tfotvlPfjWXYhzndQKxB1+lHhjSIqGC
E3E2pUIfXaec/wadxQ6Cy2syFgQ+U2MiRthBMPce5xzEDZkMr0NEskUAQzp0TJxr/H1RBbRFyr8+
+dxBOGsZWT6a6y6P27XSSWFa2qkNib0qS84PFwqfptH9C+TLJAIA+65JKt4qREXM5V/ep9QC+kPj
H4TXUdNc8YXOU3OuHOF7M8rWVAN6lcG5Xqi/EQnmmckZeXovpSF9SUH5y+Vg8UyJNTMu1AFQXiN1
4u1sjUh59+OiOxW7JgKKPjjYMO9Tly7x8OiNB9MrTwcNz9Xdk5R9vcr5KWju19ZaWQTCXo/JZ53P
b3v47i1jX66H1rhCFpdA1Snqv1XJuPWa9DvHzKcVdynqGR+3k6GcYBUlBm/2Me867h31cYTg1oJz
WkQZ1kqxsHBM+DBMAknu/9tYrG3JYiG6iLzjsm/zSvwUugrzmnaWMcmZa/hZcKHBihG1bkHeSLUA
AzVceqkvqgmsBCNsbgvKA6KI4oa9A1fXcADg5ryDWwc4X9od30vdMK+e9yW9AniVArx+fWasEd1e
qKiEY3dVoPc/lQXTfDU8zhyujEm8CZpAFKBdpugNEzWwaZYAt/SSA6VSlK5MIqmt7vPrJUpFYbpr
Va9QPt7bzc6XkjdWn72s7AMFbnRl2NM8S29i/bGwF7djj0cdCPLX2M55uubS8jIIUnjp7di729tp
dwVmeBY4aOgYrZV7oijXG+SH92P1mwTavzN7kmYtfV5HfrNk93lZXq95/sDYIL4yBQXd1rVkIKaJ
NCQyPrRQE1osjvins7UZBCHIHm4koCldIYJX/u5tKsDsgO2GJRBH0hSyssg+XdEGXcLp/OsNh29+
rMACKM1H1B/GZZLYeQUkIxkQVORsOka4hdMQRUr3woADLePIZWRpXWIhL5M07nUrp2x3byb5/8ud
FGNaAOSZCkS6kubiNWaWT3JKL272mBXyVqLyT7faZXJ4O7fMdqwRHyUBg4GrWS/2gFDZ/TIlK1WP
Dz5ny8oqTsCLd2ql1vdLqZF2X3a0delQ5WT8l2fF18qEINObJSOfzMfrbHlfPWHzAlVt6B7syNtL
pALqu2W/0lE/HqIjPg6DzAtn/nGJBTIfweCu/mM5hsuPxImIT2CLNNUC7lk87oFV7PSZEzNxcl7t
Cz/X++4G2Y61vlRwc6LjGPMEucq1SZGBjnFEY4S62sVJzbelFV2p4Gk0+NVSl+oo/iSIMmmTvxs2
rvlhJHdlNKyDeoFENk7QCHqbSspV9LTdvDgrpd2yrhGPtQ9rqVNXokY6YRV4Cm6oyuRyh0FUx9uZ
zuHVW74qFxug+cXZ9RVC7a+q4BgbpReBvZh++bsQweU5Y6sefRdq64Qjo4lpgZe1ibWr502lbmPE
0wkAXdYN9HQCNOzXH8ENCBD1lYWCBhfj/E1HqTGfN1tWEtgtie0WZdwnbg/iawZjspCxIS61LzEN
oOtxUMMqo6wYa49WuKEXWsejn5587zhXykoFkaKEl0XH4iDVW4QqI6J1nzGcvhmGfk9czYlRjeNW
qOsOs+ARopd86KYGi4cabMDDTahLreaCv//JWHMzlm7alwr4UKBjWsBjmvCaG4bseKhT0qgWadtb
VgQtkea4JPrBRUoXmw+QhHr9GDjeZealJsNyv+pe1tuVSSP1TQ4mtY7DzMvvnMEQBrm88h71QTTD
bKrs36ICg0M14HriUGqWEl+W7YUKG2rwCHK5qjc1B6/lsCIwfdIa9qKktUPNJFqTLQQi+uhHuGrI
iR4ejXjsPb9hwOYwjF0eozDNqCe7TNZN5fKFHVm3MFDSwJ9WxsH/0VS1CFl4B2V6p1r2P60VqFEy
TaiB9ukwua3ndKz8SBWWp/qE2Y650Aaq6JtPFy7utTRkmGw9LIY1w2qXe7Fhg28hj9EFF9xAmRNy
0LI8dDipOIIAmxOSHODvYx1UTbypru2BRg8bSOCginulsO6Pd0c26+1jMbSESDd7iWqdfkIOlL2D
xro5tYFyPJ1o7ve21dQ8lx7OfgBxgH4SM/1TECsh5S3RJmHazUtkujBizSY8YtBO34LXvXoQ0/uY
YB0MTNkf4nTAXmVCTMOrLpO0sW3LHkC4VCxqYkvYtRPZ0vLAKDZBB4H6SG7FmcfgVZZbAwdw0NwN
uXz9XMIsu3NPfBeKWu5pGB/hNJwwWwqT7AIjz1D2/WXEEfiTVqDAAJqzUbycKysnnbfA6LVWPKkU
y7msdJeHb4qmfgTmxMVi/hEBuqIebbTdKYvUPybcKz9SIF70p5UVjB7kfPimpr9VE95TCL4Mgude
Magn6mFbxnngDGkhg4Qz7/RoFKyUweOllV2O90U5M1slhI3LYLP2WM90EcwwCHMdAa4K5AmbDRad
99+RSHxkGoSxyR706j4AJcZp3ELKC8RYDFknvx06iN+E0x5/jnkE7bzXZ2pD4qGgBjHd+2x6Aguf
soRWGvEitA8Wz830R4uYgeNinvUO6VcnHINgRWd5EEAa4DrAfQOlDLCK/4OaZii2K37+RLzC/AzN
WUvWvyORbvOOYg6xm+/tLgOyur74h5fKTr8unLBMBPVHDWSZbDxEzANbUVQn5+JdGTF2O9Pxgr9Y
ieEeqnf6C4pywluOrCvNLAio50uV23ym9QgjjBD66OG7enYx7aCh8YxPDt8qShDat2Iqu/1f9tbS
csTPh+/vP810bDEdS1a5OB3mrhpD+hs3rjDWucPM6nXN4sdtVq5Vg9oWWreT0lAZYVzoNWgoBlJ4
+1Uf/sWj0YNgHhgZW4VCqMiCCSKrL0Wx+RgNCLfSGUUzRuqtadfMapt5aGh8Jr2ofUAYWXiZ70Td
C+SltAv7eoKgSxsSkLuADbfvVdA1ntZw/gm4LbEr/Mm/NSf0kcy/RHvhq1KkBT3MzQ6b4pAYdO0Z
KRNhdMhQCpRadDIcbzfZQ4sKbJlSegTUG0gPeRQUMvrU5R9gtp4yIhIghvOB1xkvo7Zxg9eBASmj
xe3Va/6dnlGXZFQCOqmQB1zmQl0J9D6yatUJog8hRFjDGlRoSNlNl7U3XBqpDX+Sl3l9bQPTR7/6
BRuQm57zKZqFLdqIMxfYhwwEwUYDygZIu9qhIpf3YwTt15rOXJtkCBsAg4l3Mg+tqOG2aPQk99jS
/8wFEJmC0TZfrbFKX8Zwfsd85bgLa8acBvuQW4pUj8cVWoTwAV6TEWNe3BdsTKh3W0fQHuB9VQ/n
XZpsETih5fZLnudZ1ELu4L39DLS8Mjdwm7dPxnWPcfsaylcmerKSsgF1dh/6+gI6MzoHkFngxrkn
LqQTJowanxfqvgwO3VFu/tQznvOujooWE3AuyMy9RGSSYTvgWId+GtsYRigHPuPp5yUWrgtahAYl
kQN9A22PICkW64rTMA1OvgTZHKhC00IzAPB6V8ZQccuJvPqBjXU5KmgtUdouLDkaKSqtTkNn6TMC
ykZVNbyf8Wae8GZ6+zyMdRJVGlz64xCfSac7442FuQ0hFY14DujlInmaXy6Ozyq/WLgeJHIYO+nb
tdCbhllc5uPWxFdrG6JjyM8U1O0M5onxB3cdl2VSek97V+YSs6gOW/YZkjgaTpel2zCq4/wSHnl3
0hwdj9NmSTLr6eetSaABU8kGHSYBe9pkNDy2pNIy3+D/nUuACNfZol7Kbv1Ds0MtE8VZZ9Ny/oBF
UkiFjYlMGdICie35YgXsU6E4aeDg0TuIKvte/ywr+7XVhGPmJzIBS5CBYarXFobUcggbHuSSjwwN
9J6pqVxKUFA+1KJezvq5HvjfTzBINeZJcejWG8/5oDgbWWc6fK+Pj4uPn3i+x9Kji1s8O6e80U83
2/HzS/OH8ELRl+W53wj8xXhCiVC5312Q2B+1N50OhQ8ZS1t+E4lS1R9VrsJz+rQCvILE4jC+VTI/
JuaOee4Tohe9DTWtj5b/Dv9jioOYhmzlcjP0EpGkRa1yskbna0eqQlasiZ5g4g853ewek+z44Lq0
sJxNNEIdL7TUxqge8PR7DBTD1raT8W1jTvwFco0Md9vNhIfbpj45HL352EBulsEXvCtJZEm+QZrD
mIziJu4/sRvZjQg9Ns1bwPMpjotexTO5kfk08jFen7RJE7bjM+PZ/CYqB9jyM+xFnq8jOImf4+pv
4DwpZ5Jpg1bQ6vN6kGx/GzIMkiuRa8W6P4/FLakHcPBoOWGIK91c0gXZpAZJfM3VlccHg/pXzXPs
5YxNRNZQ3bLvIdmT73H6w9GnEAHb8afPSRMHVwRSVgk1/jC+7qYvUx60QViVagE02G4KM1bIxqWj
o49LxX8iPZwVJzZ2Ur7LtcQdqs0bpQKQ4P+1FsV+bUn/xdJTUGo3MDo4u6JWCQXv2GQVSMOb323D
GJgPAYxYX5JO1eRSYT1jRzZpaCMoNdISI4hCf/V53+aRfNjdlMTMMCV6sBvF4Dh93mNVPBSPeZEz
0ong7dvUa1bYBP5wS0F14F+8PH66Ro8asVB1JAjdjWM1pEz/mOk4uR+ziHAWcL+DDacDkZaOJ7+w
GL9oBiHX+5B5v9A8KMcNase3rwcRQOJiP/8zBmxw2j/YyuP6Jhd1VcMWqayYsvX4kU3RORaWO4qM
lUqm7Ijp1ItkhV+VJgcDQT/zYUZIfBf8kDvDxEYiLYn4pylyw4vQKzRwyFR09KHXf33cNpynm/ff
0f/tgLfSjMn2Z+ZEhqh6OxgfoKe72J3pppf4718AQqG4MfOjaL7UgvAw25zb4M59IG5qQ1Wi/LlQ
uuz9Vx0oiLxNBF02y2j1i6H/SYMeyJlCDzZ6HqOmMwqzec4IitIUFkr2VsUwOe10oRUMSYiROueN
pMwBkVhZg9cmQYPeWOtSYXoBjeFxF/klvpeg1I5M4NPFF+Yfm5Ji5ORVgRRoqrR9XblWSuPgwCHN
ey3HYeTszkoRkWPfx4NSJAyI98Z0MXYw6CMIvQMb7zZlxbrK966dAb4cCJweFU3ZwV+ICDdHPewT
liy3e2QDXTzT1asvISzZsyZs7d7svFBVdPhr+2ew1XSnMDyHzIrR2AQvtR3qAUxAt+hzvSDuzAPj
AeiExz7MQGU/j7KAOQY4id4WxWUb/5DCLntInNCQdrPNjqBGmzbFBZB6BjSmL1znhRLgEO34Upt+
O0a4jvdb4pagL8qVTKwTmH7xtX9oZbSo6S9hSg1m8BYxpF6HBoRKvMfEabs0yjB9vT4u0Q8OZBjk
JL8umz4C+CuqTIhO9iVqFlkSZ0U3fG7radBFKdTeAAg309qDsSeBJXS/ATWwb+IQQC2XT7DZow/x
MGXf6s5ARP5kF9YuNQYB9c55x2PmU4/IKHNwaxfOl/Z9IAQocbrlwwPSu6xiyQwghzUKQ0aZvaVG
qP2F3qD4ibLczgoKRJmODMyox+h0w1L4TialhvWpJIm7kmbRDUhWRqrpwnjbnSgQHo6QQkWhkydp
621zTds9fpFqP6gBl7qpcS+U9SEyLahT3zo4gjr2xiDotNAr5zuvE3kmNcUc9tCMbz2Cg4PRDQIQ
Sk9+cJpF4l/tmRLioHBACcZ6nxnTckLHPDlnJRZyxVV82sVacT4A+ChSWcGEe53mKXYFePTMpqCF
SG5XBbFgLSDBHQzu4FFzuNGiKcunL1/WdbCeIMEJEdxL/QFmZksEnTBD16SOSyuZ40m/Z8fODP5r
Kz9ltOyldLKKaOf0m7H/ygoe5V9xJFlR9NNwbWB02AZRyp5J04SMTqwRD7X3CVmz5SRvLasiV52B
GLKYHxzkh/lG8murHiuarGCBq6O02+6fhGYUkMH57TkNt2vrplqvHq7msfdwtzWMsaotXYqkoOHz
K0LIfUKHamwu114SBNj/zJhy6KJOGFu5obMWnOH+5F6Un9NGZJONBJG/m56w6czDgI7jsFYV9Xc7
p/XC92vPLEd8GW9pycd4epu/qRn4lItKnOCUpS3wuNeqMVyi0OLsv/rWl0xzFlppM1ZfwKiAhv6Z
SyL4L+QBF20hdp2qmbN7znQNj4Tpo827DFugRau1vnn1iRg/xsgwdWAdYgAtR5BuQX1s3+oz3pGQ
8oW4vq6bIkvvsWjB3Xtdmh5nKbyNU2j9a5KdPaVhTG/Ov2Wx5piLJFfCWSSsm007lqYH4IyipiuM
GzzVrP8if0yCM7HjFwQLA5twb2OBYhC6fUuvDxgbHH0flY95wRwFVMuuxdz6U+psvpw8tAnCqjvP
DQqvDKdODHgM9XMtzSkbn09b3Zuu2XuZMBr3H7IFrodk0KEGrQGeC58K/YlIDSyliAefL8uH6sw9
CYdImSUoKb2qI6sEam9VzVd/61QdrMsoaN86JabHrXVavtJ7AWJj31qDnW0wjqj/Lg8LicspjQox
kWATNJb9if7W/T2prmTQF5eJE/3kRwz3KRIoC3gijKmUmbAWd/Pt+usrhH5pvVpE3o4ZCWkbsepa
QrbhrCp00Nu/bsGXj2T8B5Qv05+/mb2w5cYKrOswaCkt1HKEqlHNiP+ECLmiXbXBYzCM0QfrgdLz
Xa7noRw/sol5E7/kOB9zpc/qXaBYI6RC1MLAIhvco9JrdXK17L3uuEiRqahwu1BTBOPk4uFkXGQA
FRsth+WQCBnIpQIHyC6boQ0/MsrKaZN18QCjTtemYuXEa9hKd/KnY3C/bTxmN9BvW+P163lxGgQV
VAPn6MqpT7S0zEl8VWv7KaZxFJl6lJnr7lOJ3b0ADMG3XVc/rxGFoRMOHEb+/dHphkCc38v4Qd1K
XgtoQReYl7YvZbsbBrXAEWt46E7ZVs/3FcPLn5orV0h/28FOA5qecIaoVE0ZczhXw9K+0zqjj+tv
iTv0iN0krTl9Fys8QDvh5TTGAXg2TyAal3QMNnp0+bgm8UVPAPjhIKWqYT+ADXZVcG/RyhNY4qM+
JWpXC6MF2c7gi5HvoNaLadbANFFinSKnib24IrgPIm+tsZeiTXY05lm1XowpK95X56WV7apJ3jDn
CQNqnHEq0max+HZYsXTZVLBSuefDNaqr0W7NtqxSoTSQ/jcm0d6Cc08Ap3F065lfuCiXmlpKTbav
qvncmkAwyFL4XZVPZaQd8q3Roozji7x+uJiPLB0iRG4v3T1P2c39wMSzgPj8uPOUn7DdX70mTwyL
2Kph1AOI4ERdgjU1Z4ZxPtEn2zH/+smDYQzj201D9yQP3nTyW1+k43e6nSZuztZE1eVqswKa2ab/
H+69tAr7N3VwpOdgKYO5uNalwXGcH5GORflTZoK9UbC9Xwh1ZDokYUn5UnK7XGOh54YigkrzgSBu
99xiDRnygCSSWRE/b+m/prB2vn/kT12ibvQASHRdy1s7u9nm4EBgkQq/1otBsAL6U7cQDKmZvmfS
MWNGuutFSnukWZV2I8OLh+W1J2exS7pdc1pFdolebWwN739wxCw288suO0nO+BwxUjnM+IvuQ6eK
3g4ytehWDJAVZlTB1GoOzEI3mTIOt2x+MbE2MG3ul6MXvmoLkosdBjte5li+sJTldPlhNZjRHrmM
sbNJotg2uavtx+RyQwZQw8fXi3THI2DguBPSxkPo4Zg/eyQjd7DbJfCmQ2LKS7cdSCsKNrkZgAwn
X2Dnxz7FU0ASjMhAQ2FBZUzhL0iqDYxcCf0UxZusugXsIUiciu5AIRCflwpyGY0xTw/BX3JnIRQO
F15Mc3FVHizbdWxQmcA5gqj754Ru5xvyBkk7o6lRkkDWGKHInD686lK8zJVAGqqm89z0YZxGNYyA
GihWOsQNMh79g0LQY9zROuzxZeZ4uij/g6GIBCCfoZx4uLK+xbJYzfpZXhovf3Mfz8f/kOHkWMnf
J0eSdc2if+Y13JPYb75PqyCk+bDNXwm1Y/6fHd1Xnh6/UkRauZtclBzDSjnf/ZYEVgLLsERFw24K
VttGpmzGRtvAo5wn9nn0nF9AdFzX/XmMCgL5q56RNqV5oB7kOuVNXQUuhlvsrn21HmCJZeqWKpQT
IjMbPfcVwqVEU6voGg2/vQ/bfnzv0rd2m4qlr2qdBgqWIXuqg9Nw9dSnYTykzTCrjfM/i8a7VRNg
K4PYJa6xxonEmAXNEI38C8z8eLoEcRLXF2uu8R3pJsTUZ5+VpRCkKVka0lctK6fXOEYJydIKLuNY
QZytCwfSvpV3o5WTO5kMljJoG55Vbpi6FH5VENgrzUwXi1zn4DXi9ebHjL2ynjXPw6UOh90Vg9TB
uG4pL9W2B9FD+EaZj4Lf9V1VKiUwMEn9bXVAZXbayRF41fpi0wGeMb3lvihRA5sLuDN1GwIX4518
FJqR5FoIqVFUY8aU68Elby+9Xjja7RDNPblTFhVaWUxDj1XNAUrwt0ymKxsXmAj54GF5SMGvHWs8
Qlph915di45l87/7QdAq5thb8gcUzYIAT1twZut6uqSL4O2N90g41cD1A6HlV1UgQO5YCS8N9mIq
kwDN9xwrdAOwJfTJrzYC5rWSYJl/vPvRu4MsbSzRGrYLICW7klNMpzisOUqZweCO3P1Cgut/RqUl
AXOP8TsYWvBjfIlYxvFFc6vfu6b+gPt2W8yB+4o+aSM66ssZ1pal0GHsJ0ivNQTrgJpcIUyQ9HG3
A3l6QFZB+bkfgZv9n6EaNLkpyk1pGemepmMo/ZtJdSrcXbFBnLIMf+FYpLcKzZ/ZcEpvmTI8tyPp
UDD/gwElErSfKVnXD96Yy/1b0GNcpEOLRLqbulDeGCfNldggwE3of93tT+9cucZVRAgHT39h4lS2
I5FJH4u3UBDc4QwWGKHdG2sAXsFPoVjg5zSIOaW+yRR2YpsUptGQW58Ktj344r7TVIeZryB2KgD3
Q5uz2cl3M03emLu5VPI09KlvCFKOO0/a24RA1GnFLaOqrGX2abNSbaSceaCzWi2LuFjQYvreSN4C
kCJ8r5cRW0lw1DlktqXMzFSqsl4rXv45NUua1r3QRu3gSDdnMmt6etOjMyuE9RVQgwp8ypFAFVgS
1nhpaWhHTd4nldt/2OKmTHc/aRotYo1+ybOduB4HaM9sQh47+F1NGUcDHR77q+nRrZZ9A9QQx2Md
WV06dNxSYZvyH/qvbkx8On0FATwXG+hurKnwMZ1eAI5GATAVyAgJCFJuBPtIcL8eOivp7dEZE5uZ
dJi7mSlRtLp5H8VyW7YYEX1u0nj8+TR22MMK7oVmhhoauE0nu7Xi8aX+crlG9ZJjZhMFb+v+v+rQ
O8rhDQBDlvn1raKbA92Uoa1LZzUPdH0jxO4A+S0U7yrywfQIouij0F0rBBxy1Zbxk37SRGc+WJVm
vIiGw5sKtPplzWMH7cyQl5wjmp4qtWgpDmw2U6CE3VKL7QO/VrMR6BXvcQtOrwdhllGuTqY3wrGa
M+J73Sk3nX4UHlb1GRUSVx1HzfjqUasgwNrAxrh8Fq6JS6wnrzwgcvkahsquwGOY8zkuGPrSjq00
cAEoTVUtYAxYjt0SVXOzqK5hgh0ejVWM7y2mm1dgOrqW/4GFvCFTTETAD5YegTqrz6ukLaM2U/Ws
NtRiHfLiOO30hAQyKR+VBoWx5YY75pCuYXW68im4HXWcLckERmJxrdsK3kFqV7uQ8yWjxuf+IyHO
DBz7oUdkVvMfPNCi63kuP7UuuGONSKk/nW1SpbZvbPVX7ndE+HMNYGlI5JoN3ZXgyGaQrcPJrhPa
DYPAxmbgX9pdpKWPICEOi0DL0uUnup06ao+QVfGF92ZWbXbIkQoLWIWR38ylGAw8bjAAwnsg2Sjs
Ta0RKRzZ6vfWOELvRILm8YwKu4sfHcvCt/dL7Ny5JykhfqS/FEdOjIO4P1WMoKZWFHuCSC8CACH5
/YKngG/16EWLL5sXZtU2RXCdCqIRrPSqtWUSW/qsksqX4/iMksYEtELsKWkyaMUHQ0oH0X6e3TF0
7AvpwtAQmEwMg+0fLK7/CuqhYQxAsPRYNKZJ3Ugtbr919bihwbH3TVCXDDX2ReUb2j4g+wcZEFv6
9ANEY9ak2nxLdp7dhJYswGmbgW2GUItUyUVET+JKfL8+25BdL3sbcLVVlH2IFdaGyWh4+ChlPIta
kv6MKlSZ/g878j6G5N/6KaxjygbMpNdFGw66ASE3GDYXjY/YnrYxv+/rIPYkoIbndEmKxhBxsgjc
9+nAYAp9JwJmReeZNhdXpvjW9g3n8L/o74lmcG1Ph8FCFK3Y0uCK6ppqBQo2gjA2twViDrmrofj6
z0SSXHLnr7jcGno5dxm56FQpupCfDwoqNy9YZLuAfy+2fWMO6FqdkG6pCJdk6KcDDZ+PY/OPf4Aq
uO2AbPAlyBPQmnb9TdQWDVFYAbPhxMrcZBilx/bfqeR/8oVZdBz0J/h/RrTafteRfkgTllmhXDM8
YmEPzWvDsTefGTnqjEKRwfwWsSEWhhgchbRqYEzhU9c0Uo+9PQZ7ls8JQ17WbgJcgh84TIQVLtoN
k/k97l0tIlSDAVl58G2XswHrnQWdmITuNF15JpshNj1lj2s/dAo5qkpN9CO1kXmIL6ZeK4Ce+PZ/
MLYOwT+sODt06E7NfyJiWXrBTXGfcsXkKHx6bmO77ceNI0/W7KkXnhtlVGUvzSZ8tSGD71/IPxLz
qeLuZ6A+DVuSvdKZH2zLpGVPUXbKdOwoBAE3LvUzxGrePLuLSlb/XnlRyeu3lAmGvWaRvqT1Jv7q
agId01LfgdgeR7uvMQYI34DdK2BkXKL6Bt1lbCsmnbhdHPoBHTPMZAcwVBcUqLkjrAE0mRQguB0b
unBYrDL2iVBt1XuQ27s+HYjENnHAtAknwf2QRu6Y5Vn4C7fF9IhNzG7ne2iXk6MNzHu2lUfKoMbP
W5H11g6/Rt7AA09mxpKH9k0RENq39M7owmdaxAZOsAMyKUHvl6jvG1zKcgMUH37Zg6UM20faAqZG
aZi4emzc0jfyH0oqKKfjKx1l+YClVS0CBCsiDa4W6SuXog9p0ynqIm2wo5rzrIb/nfwsc+eNbAnN
M588yZfJztudZYQqfLN0veZeHnlMVyvOm1SjMIBl81B00UqDJg6D75imDn6XmSoRqLTI7t1jzA43
uuGETXKH2M/Tw1sIujGAF6iwGai+vkWrzqO+mO3IOux9bhSqWmbMShdykq/b9YV8XFMR1zNWO4KU
inRZvzUNC1x0QavyPRU5buZ8AvTU/tvcNSGYG+eR1CNc2SRkG+eSg/WkmR8HRD71AL2P7DlmzboE
UGObaRwllQyI5y9VywrWtiB1bDOKXwZ4kPYDRV0Wwh7bdCXRL1/UzQRpfzyf6OJB2HvClZXiAP6l
BDJMoP0FPq8jpNK8AhK+B5tSmmmFPTcqCw/X/RGFTQVvhAncyWp//i2+lnaRLuKa+BtveqJc8OpB
wqd1az/MO94FXsvHiVnveKk/efjFGSrDiVS5+so/tOxS1+InZ16wdq//b3cS3Hiox9m6EZyvndlC
3SXmvgLSk6NX9HCoaoSkREp4gEbEMmND/YX8c4qXtwZLAZkA8sIfkNfEYC2Rrm0wJah0p9pNrSfF
qdSO+GusR+h4C+IFrBfC67sQuZUzGWkFiMJnWkaoynADQ+2x3ypCkauOuP3qCt1fgAlgqvDXKJ5Y
ik91Ea4GzJeaV3nzeXSVLLkbkTXZ0xeZUY3fKe/pHx9UaCgkAYZO0rHVahNjbSDqphbY0dY8LWgo
zYOdNqLcYSD/S61FSpU6AtQ+//Ollip9oUbHfrucodIjx3e8gnWOWQz0KJzHiZmgYG46TyiZbvM0
YlwgSr79Q4WyEO/E9Zf49csH9mUF97JJVXUZLdJNxGRhvHiY3dXHfpTao/Yg0eQ2A0E1/T/RsShW
i2nZ9OdqSE58paPxfmhaMbWjiFJRUhYdH/Y33fRKxkpJaJpc/U3VKl2/Linw5za5+4Kcr8n33pg5
JxCb2B/qkQJ86pR5VrAh4obOhJpeInc93iUAVhaLPwq1rYQJYHxrPUDZdlJW/ztQVXiYQ3dp3y5E
0rPB3OqPVrx+Am3E68C0P08YIkauqOIC1M+ImT4Zy+5tAKGL+HUKZkj1FIQBqt7B/9rfxjksj+dH
fVxceqnNGLrtTui+IIZwOWePGI+6/I3ukJbFschoOYHjDCo9iOV20L9f7Aum2AEC9lxGrwAs83B5
k5G+3I0VairacDbC4zKk58Cf90pvMRQKbc1ncCTyAUZeJcbzVt86sNWDvK0VPO/NX/dCIyQPiJZA
1eO3HW/022sZf9uneG3ShJmx0Ch4mpsUkQ3YJgJ2PTdgcXyznL+h0DlRb/wqsHe6i4RJ5uHFpaHE
MNk9JGxnqXrWm8kTbwkxU++SkfC4KQH8OGq+3BI+WZUwIk2Z2Lc4IyQObdpTRpKLdlXUu32UWGL6
Iu+pFAoZxy/hjvKtJuc1uO2C/4ClOy4ydSm4IlOxd2RPrxmIpEYXQB/Lk7HmYbaXUsf+KAK1L+GJ
lvOOT/BCz7GIqUm3HAX63W/m1R0PoAoJYeTF+1KjJqoGYeP5Y78CL+P9gBnRjJWsPzlwg8np8DAR
QWKWP2KgRyxMfVJpkqUfAuJJtz6/QdrCUbURLQzy58djYTIWsqjsxzoRROHHftS0xuRx5wTYEutH
qpT0o19khUIBzxuWkpX7ckhUkkzd6m+SmF55q2cgiYybdhn1FRCS7v02ruK3UgwuZGEnQbRii+oY
8fkoHRrfRwa7mrhbD5PVuT+Wj7uhjvq23CawLnzSz7wMEjc97bUn/vRhnFDSml1IdnRRgo5K7bwU
UhKkVbdMysigykbNmoG6QWNXQt90ctTmo+OvMm3VzEjUwA0t+0RYO79qJR63yFDiwf6hrZjsuBuw
VpRBHA15/IWCKMymX9Z81Ul9UOuDxVWpzTB/WLnOe5iEMd8Rl0R3KsgqCwzWilN+mDnG+Hu0EsqQ
PrwuyyIiFyOX4J5rkBCl55xalzn7pOAssTJZ6BPCJ9M1wDsXSPhcVqONyxP4qESsBtupGjDS11HF
rP6fswwM8ciIFx49X+JUzqUu1QYz0vJtPt95mGUW3ZmRsZLZkdz1duBGtVRC9Gxch/ZpEeCMVwxX
1punJVFClmK9jDmpMIbd1BDjDJirwDQ4EmWQ7M1CwxL/FhgfuD0KzbKHm4RQtZlpdQLaaLtrHEhZ
bddlDA2ZU9pAErlccBD0sQv0xuTD3lB/0vKrX0GCVsg/Hnya7vznvLaQtgm+VtmiDAOHi3nY3Zu9
FzToZ1fnlB/5Fq1COtRDb9vY1il6wMpOom0Zwt7rj/8QeGpfbOeUZU5h8w5uUeZI7+aB4P+xV63D
lfR90PFxUxr1cFDb2+c+QykJsji68cOtfyBqywebeU7xKi8dPrPLBfc34pPcetz/3FL67FgX55O+
4oyb0KIyUBtDqlUGiwe+e8TzZt0iy9kLnh0nhR20KgXVwzHiPVWAeaLHUvZgEjtgYT5qmfVQyvzx
nqeBRIaY3phqdBiQ8yzG01edt6DZD0UgSJlvgTXyQA7lWE8gdJbwt4xzhfSuCIqa8P5W5+N4H/7Z
y/OR/3ZOFRBNUlQzNICWJn33FqwBnV03B4p6OECw5bzqMEz2pOqS+fRe10Le4PdkRceiW8GQhGtQ
i27rIe1DkBCONz0liuXrxkCVzqsUYa3D8+jKUPB7fEGY7zO0nlTPI5WTKucxLxsHdLeN7j4gZSaS
coITetFyUg6fsF6RQT6QwvcltuvyAPmfhmsY8tiZDGAy2YBAfUIfQ88I8FSheYMnecyF7eteDjZe
3Le6TE8tWO1IwB8fP37hLDd8r2/i5OPAv4gIyt0pJ/xUoI7jAl6XLFNqpM069pk8b+HlKWjmL+2v
S3NqAFLVdFMvdH1zI0t0rptm1ZwnSdXFaJiKYKj36jOlNo4vJOmlcI0xrUaRktXpCNrsA1aHrl3T
y4VHvqwShzQt9tZpimoKxM+Gyo1IwufUjJavuVz7TNbDBiEy0filiL1FNpBKHwkqmK7YOXxkEHlK
HMYTPn4vFGvMScgkNJZEt6kwkXNrnkQP548JiaekgMfeX5Mkb3OoblmFlGT/RQQ3en9+7F5aFWQA
f90vwCch4JofRh3zmuVCRBMhD3zZ2GxbzSLrN9euR1/Oooowgvn/ch/gBoHRG6D9N+d25lQXZJ/V
k8vniHtx5ljQyPuhVSOYgxZ12/9u7TMnrAdQEx2SGLUc0r5zU5yS7Rq3sLSP23sJRZtcrZ5FdpLv
luirycdNntKjV2ZpQaSEgWAtpybL+fN4Q2W4IlpTGrGveuGFW2xmV2rM9qKJCCnNH7qt0e0UJlyF
l4J9qVCqpD7XVvZWDdlS7TGi5PWAVHzcjj5Pb4keNEqsSQtge7tmwjqUbrSQZ5moscsU9ksc/oS4
nawmbNz+2GeKMmwurPj3dBUDv9PasFI0VNdtVKcOlXdpqkvGHkL7/bTXe8WfQzJB4oeduQb64f4S
tyPVVbFqUp/rTqguIPI9DAsomjZXxpxmXC9tyubiGLh6w+mRfrhw4sQyc9YhXM0ymhkXdmUfI8er
tXjBN9svEBZy7erLwl1guLQejHgxGLpiONB9tvBofTschaXEP337jSP7w5RpS9G+i+L3P1F22p/f
h7ZeiLzkYZOOwMr8NKnPmmyr9HvMcuf4BUML0f2jDQNaELLO50XLPpXUnpo/OhbINlh7olzkeOKp
YIDW5cU6pWrwcsSOLrsiNGhz+7llBv4z/PW97UEpGqq10dmEVOPAxEPnn7fEE4afTnQdCReigcdd
4jPimzWbYw4BHMK1VDTX8p9rer/dXwM0fx/oDToehWV4CnL5uRh1r9hsrIMVn3aS5iqu/ImgvHjW
yACLECjb52fT08SMRWGw57k+skjgmjLpHOUi2n/A45jI7+SiaPWS+h7PP9f/qkP0Csh44M+YvGAS
CA5kbg4h90ZrWJ9INPJE/u2jQiRD/UPrZf2t6JS6I8TKBDOlcnrNfgQRF/cgD7eBH0ZfLTSaOhJ8
VtLojuA4j9UY7Y90et8YA0y02xrXbf6Kq9aiSpfQQS/yCZ+ukXcW33Hiv8bc5a7GQfVIzBmtvQmS
GtK/56gyf+LmafwVp5XGyol1wanZxYEUh6R+jB7cJnAIOHwIBr9ZdE9/rKvcWr2kBVqshrTr+SoT
RVlP8opoDChIsbtdwrnyipsrPZNZn36Fd7ecUH3jiT881V81fktJ5SIHZQJKCZAjUCdukiSbQNi0
Yak8773CGvYtodguwBXb3WQE0pSUWS3gvShjlnIXGUa7XMFJN8gzFfIAyOkAWqolYpNrRnIE4HnM
NEn/yI+fqgRDgji8CyCt7gnmLAJoAR06Ix1gTsDlG8ctF66w3JHMgCN5yskTCalKbTlynxt7Zh40
TKcncbOHKGN5QbyJCdNRuKW9tFvDig7GzZLAJ79w3gSNsjXdG1isxoT98iOF0q9b+oEq/hX2rUo6
DxeEaBAHnjlbaPs4yKRZkYPGHAETshYSZXlEYntWHARv6S0hvZj86iQDtFIfNwvxD6v1RAWsjbTo
zPa+Ed8dTGf+4ITviW0jY1ShAv68vwUzqsmb69oFFObPR3fiDCw2inve8U2OvDag5554/IFSiRyO
0cRyWNUZTObQl3aidTuWtCAkP6aswprLnDGHHjsqvOdgeiym07oM8f8QAe5L7LXe7kebdHTbpWfi
DMsn1QZd/o0g1+WKwzPmlpggZ2nTWQPAJo2nb3Lujmt8Z/eDULHDGvRYcFFkbpf/JoEDxKJeKIL0
whVNLU/rG2lNIpek5TqQ4BvHQvRcLsPQY3SfCR6MiFFWqXbVlXiohKjPs5fhkkSZbRcF7/SxCYv3
qZ84ZKD/TucAu30QT2u2MJrotfpAF+GmnmveEy+CjLzL4smxJAIjN/hJYgFkPKnBmZ7uWmhg2bh7
P191x1/LyzgrukVLLYM2XaCuLnwt+JbXVWBjUyp+IDSz9yIeTEIvLUofhRsitFiL8+LgJQIT26CA
tnDY0rsDIj7WBSTXXHNqXNYpnPccxRmQo2051OpL3MpavLZGM6Ys2aAgpErRnXG0aO3Pz5pIQ+Rw
TIeJ5YLlFN91UNB3EuKCpk1wC1vCnoRkPmIsHkrqvEDT9CIxM99C2Nsp/F2S9G0CUjfLzDtl7scK
FfFpq8Ttl0tvfFp0k7wlGFQlG5XqfT+eHhhLizgf98DIqXuVFd3QF/iYzcGXi8v2n199f0dAlcJ+
uuZ/3bQNONwp9tkpFJj1I1ClrF9aSzVGY+hOF7muVexF7W34PiFBt4HLrZ0fcQwFSr7VHGxgpH79
ojqn1xvKLKBjl3dpi2zopUfaV6NXYgNm5FNsMZNerub+zziQCeFx2KFTxbPl3vR6saH4qpSE1AlD
Dy82S2oTS7QWdb1g7lBeMcrjlC2s/T9CZYGyhMEMj1TFd3jmF42hP646Eomijo2fsPQLMIJMBESn
bgEnVSobo3QPgeBr6+nXEwngs0BrIQcjXRKm+LWChxbBQpzHS7Lf3nmp9vkTPYiwU8Dtj5eTD8CB
qA2kIhdf+52pHN/h+hC1m6LzdQlkQhsPdTGqyxayrPXV2XRTGt0LSSWMSmzWfk+zizhZVmMggdnC
n5uYMBWTc4NA/X1J5RFe0Dq6Zl1Ebm4Fo2fmOp5+3mzbuS80gn1qdNcr2sInaZt1MnyHXDo0Zxd7
Vmstp2BTEmHNvcYRcTrZABwEQSd30UYDhRRsNqkgB2a2c4exGdux05t5nYWtdu7FM4L4ov67v2bW
knxn7Kh6t4iHyBkR4TR1uTnPbcuVDnPKvI1m4g1gAqLYnF5MYUIB1XcksJBpS7uaXYTVyFjBcVG6
KvxfBmHQ9pznBX9cEWq7ZnfWYOH3/Ko2CiQWnY9/1CieK6GjtM4ymzdVM8+RC23SiSSOZoOsa8rT
M1j9ner8O374UiwZDsqZfnA+Zt8xPvpGyF0+k6OkWF+Zrvn8M/+EEX1BorBwkL0B5VeOvgCaYB/B
7a4mq2kq+tkLruc2buct+O0IUz5eezCvEM8iyxdOWw+hbHNKoNBdJDhowB37huEbakmtey7G1yY1
VRt39Zt+BKBWE5xxuhy0nykZgb7YPArVHdVJFUcv5dVUcFoLB282ANBXBQ0xoaFRTQM7Fucb0/wL
PL4+tZjuTOqEhN1e5qrrxTp4+IAxmKwG3xunSCVuc1V+V07arbXrL/JB15P/vvNRvaDHhG2J9u7w
C4+n4zwzwSCDT7O9m6lcF4LOjaSRnuVo5hIdP3jGjbB2B5KEj3NJCD+xG5F5vh3I1NWQmGNcil9W
U0rsVYPQQUaH0MPqENbFQFFY/S0Z8OV6skp0bN8IkTmARidN3BQ8Yhsad9AzWc5+zPbPe8T/og5A
flGXGPows8MkzweXEBZEk+A3nPm7QqS5X6biHRyLx6eGZYOwjaGTsK3IXStky1Km+7EQou6s2VyU
Zoc9sTw63rbxGB6U2AplDkP0+q/hDDxpfiszYXI8zfpheYgL+/X3jGhLT2CrnFXq2G414yg6Xgta
qgRH8naZEGPJOv+5TyOLaaHibESJeQ2JOqDeLFSwj1kc+H8fAjku8/lObHah52QiE9KdnVhelXDM
wSoupFjaCNcO/DOWeAu7CAWKtJ4zBoKkmykC0MdCxjx5ZfrSJEPTGd3prFsqaHzwmdHzcdvrBq53
0J+Lyp0kupZVdAfgzfOJlSl/KyS72UDJizQzUVXyy4sOOUBz5/d9gqSIKKrjZ90o0U2bO4Q9HeWz
bVVS4dYIcsXatYU+rt4Xqg/2Pd+pheCWP4tCNnH+tvWJopTNUmxD9r032HboI+ALwoKB8l8BG5p1
SJbYH/nt6tIjFdP1mdjiSWb08/gBdeekiErav7Wef/bnJphVLggqv9BARDbRbv2vSnMJ59ANAyNk
WTXbgD32q0H8PE++/6BHkYcX/7A6D958hO93ReGgCviwMaZq3GybvJ8vtp1t/QnkcuT4Q+2dwxbA
0NDBYlYGm4YWhPuV1PMCVrDQzFO8IU2WkrD3dK44DaW1MQkZZPPPWO9Rx1Lz59/+lyzG5Om4BXTx
ne6Jp+o/WAx7NApWfcdhyq5bzuShPVYjiQrdjdGVjWRMMZGXqwdP/5/EhlE3zN0MjF5w1UfN/9Qh
Uv9FFy/fKTGH67gg9Dj95qE1QvATgzt0anW5g/qP0bw3XLkVaOezLVlDxbhHfbQrQUYJt77WQjRC
sD7tkgl6UiJt0Rkdd+cyaq9DEnytt8K7+Q5InipLsKnIQkqO4sg5xKSXC+p+LwAq1h9uSE2n57F4
wjyQo9LgA50lKIw15hyqjKj5vxKnKCNkb3+4KJkDfj4ja25/jWgrIXvcnbPVurmBDJZtfFDvSSB2
XzqGuUGgXSWyiv8GxpUVJ8FUVXRCDg8yJSPd8Sm32L9WJe/SU7yLz2g8onwp0lmkaU1DEAzofTrE
t6WbOZ+5eat3E1/ahL81QkUlXFQ30vopaXBoDWu9BadxrE+P0pEvKXzdm6biBZHa7OkVsVGYhGim
ZkTnbcYPqRhRucwsn9oCttytoem46k3HK0B1l1QoQj7YIcIzXxNHyZTNWzDfIBERgRfmoQzJEJXB
hAF7UjMmMvO9VCh7UjggAWfPW36dIJMDiay7MAaStJvBGbhfw8gtUwpZ0YCgyiS0CiMt6cUpKqRN
v2TkecxNIBg+Z7iVn+0RuIhbrL3bGBOcrqTFMHiIlbOxRh4Eqv+lf6gKRqrhBayU5oY7o10R/EQc
0BpKbXBtuPrZoTfzIkv8d7hdTkwSu1VwjgREyJziRTu+5EexqV6gQbFG6n+JlZNWhCW4jw6Wkx8I
IscgMZBWGbOyRlmC2BSkKoEzGaPqwZPjGKD2LwcmWzmMP3IAaV5RNyuVgygFJ9bPMGGC/xPSGj9/
/6pcXmMXNkkvxhAlBZs+yjjFMpwwjV6J9oqnVsnIKocYxLTkgY1qPKlzAL4VwXb88eSbFPLxmC5n
NFOXMfzrxJb+XmG+7Ik7nKbqMnPXCu0pnxiUulnsQhkj9lS8Kfm9cA5A8ii4ZhOGosbqjsEo76sG
u7M2ZATAqEHtHj4JVrE8HHotPH589uOfVYrFjQRj92ybniRvn+sW2D6+81jT+SktDevZkLRkz6vE
OTnRbrLt7MFRxf2pi1LXfRfx8ThduGJW8gmQb0GWgmhob2VSD9/Es/JMmTBbCcvfiepe6tuWUU+3
GWSGiAuqpd3vgINKW1aj3ZnkIZ+dez6ahIsmlIQJDez7n+8zFG2A3Vf9/nIJP8uKIguPh9RpUBVI
89eFOpn2X3jH0U67z30xYPXLjIPf0EdJbFsjh2KQ8qvVAj8EE+6b/qcnbK//v5FDTTkSzTD+z6Bu
1MRpIKQjkq+1o12uFvaCRy4pLJVbCUCFL5ZuwiJ2mApWoPSE3jL+wAwVayjiOFnfIQSd9Aq+qLWk
FHj+ki+k9GWfCmPRoEQ0g8le2Iuw20NBwpb4BBou/cVdEGkw8ldCotTFs6/8uWerlD3eiJBwKBhT
qb8kezuSSSIIPIiKc++fjXckxPcoJWitMpIaZnK6xNgDayNm008ewfuVj9H4Kbev0dIE0c+AjGlO
pb4KzE984uplpRoUvE5NGwFUBkpw9FKiS16dhVL3qKsPFa/90oXNUK04kUFurD2uzwqx+EFVHeHe
n9fQseSlj32/cPlugvf/bmz2OaxhDy29pl0RKbTTE6m20GdId1xrRkNkEBgH3ACOqCXyvG6C15tc
j8rVMlRWIbwU4ENkUT8cXXk+0+wxg17vhNRHorGJFDg4yzN9O3erUohtTMxlInOdM8HWCeK/Hz/m
wazLcrUUahz5Ghqukr7OQvvC6xNyE/krtHTxi1rqY3Sr6YMZO1ua78H6aSds44NrfovGWnrUndaa
iCM5rQoJMgUCMO0OFkJguElQSvGvXl/7wwYrwARkEqcNge2rS6YnW7GqbC4j4ZaqIutOZkz4QuGq
jzOKzL4T4Z78NIQTAMYrTd6LbgkjU1tMMATn0k0hkpbrjGEOSvzhV+n6duppaF1iW0rDYHFe+KSd
DmtQlrOR7KpPJQTlPKrO7Ph27vKtoD34OxhodP3zDu4eGIC+AQpQJtGMSLRD+imEnC5IezLT78C1
IZMfYdtqg4hKwUYyf/y1Ud5eRloor5ma+eLwnBtvUUpr8l1tHUMRxmFLqcG1c11e7vFNEnpxa/Y1
CkP9xundb9kfJxeNHZLlHFj3V4Y9t6FuNNHRn/9Vn2ZIM9Ps56eeRIK+eW7pDVCTvxP5m9Wiow7J
T1JPmSSTIsNPMu/W72cION2Wrmn4hz4jQDPnsMxImSSon/3BWBBgL3WJ4X2cvpsPbGDsK5GjtRpr
0NishrYvGCtWIFfIjjiajXO9Ibf0rgjot/QpJwwavrWfzCuTqtQHLhvebYiQk3Ow4CaaWIY3oXXd
WDoidqUETLh7KeghwL4mexeySVEcT6yLr21dFiOzn4Mi+SuNZlpon+N3jVSBmm9eOPwmXCxIIxWQ
Dq56l9Zb0eFIcdOct6qXRBO7y3L1ohzFkCboLaDhbi5J4+R7iHV+J/mKyjaz3xB9PkxcymsZVcvv
lYGOwssNJ4Z4x0NQ3mnWuhNFl9QDSeFgtPDJisWqiyZmDe71eIIjqb4XjQzOQjDy0CjrfRjdcUhN
9KNYt0AepCCe4TG1jwL8eMeTL1bjPEQ8E7s7O9fIdsbOMCGFm5cjO/32vCekVMvBmVPHfMaJCsEV
lPRnyJml5b7iNUXrMoB5Wd7uSzh9wf8EJoc9UJXDb6COwZ+0s0AMbY6hrON+rx062UGeMVIIH9jT
0NCIC0J5MUtvxreQfUUYqGl30CK/1OzfQWoAdFRe4Hixgok4ROfJH02JQ+NqkofN0DUFWDQTfAzH
oTOC+l7d/Dv8pRfJupPqMQZ0IlERNxqwWd+Lr5xC81JaaLEMmCct9eSSoP0CEJ7G0eaB0GdfpN7j
/5/y+moCO0I9EtD9AA/6NvOZxfBUBzoDWZUGvBFifMM/VFwKj/UcAvNLStJK1RCH+nSe0vpaplDU
cCu1D1883YbjjUZZUvP64np3l6KXPBkwOqRjpbqPtg7JHE31Ee+naiFDbbylb4HRuxwKFX7XjH5Y
KyBdSENvoktSsqUa3qVMoWsXxpUzIvSAMLfOKBb15ZP3whXXMZiDJ99Uv0F1F+O3kgJxrpFi+22w
pM030WQmh4JytafrcJp1DPok8qg3s+HW8HGLqmCwC9/XsWPF4SmLHgkqbJfpMIV1sdLLJvarVQlA
fzrcRihbrbSiAiH6Ek2YlFhStS7A2+ySiUdaOHyMgwdHD/mAF6j7nJWDXHm9g8W6sRN+gw47+gil
SCBJJx7QjbMvoGNhDJDwj1iqzDya9b1TuRrGpSY52oQGJR5sxN+WBCtjUtfZ+sGiCrHdv245Lmlv
dEZunr7pptz+KBOskdwfq/JI4tQrOfMzpHZpXK83rjO3CgVhtJoCm5i3EmqfwtrTJ3CgEJEWHvRq
F/BvYHnvktsCm+QbU/sj48qCOvFLrZ6ehySbM16oXJjPQ7UI01YzmiZttcoLgg0NHFOIrdF+Hfk8
+4yjkGK0ZCH74Sn16Tq7RqNGBuvmJM15vyouMngo53HNXrAq2twV+e97onEEaFf23sUIHnMf4RJJ
MIy1PQIPesOzWnG6AKWBRZYPqpdd6yP0hW3Xi8oGMopa+XVFlMk6mTxP/yAMuYK5xH2bWEYQeNiw
bYDxnNNtyNhfitbeHMsw3zVGXPbD4ZlMaH5v7QwqrRwh3nbniU2zNcTnN8GIm4kQKn0c0Hyyhk2V
pi1TPLfQb7xYpJ4iWcEQb8e24xpglXGup8rFWVyHQhhE1wqMy6iMZOYQ8eMFuKl4bu8vxWMs13iJ
kw6Q2gwFjnvEnFRKGsSiQ+5rJaXphe5zxWJwG0MNBXhf3WrdpYU7siOKb0wc6MhNK0hF3fn/I8nE
RZYPBG8vcjHifLyFgpW4gYKtqxa3f666X0wUilLzYjd4OFnjz7FLA3/JJjwJudCN8hTuHAcUoqs2
ZWa0crYU++TeHP1QrezvCBZe34Ofh9yiTOldJCh+YARV8/vY8NY62YXyn6KbEe9ZxZ4Z+EKGJAnY
yKReASMR8wlmeKJfuetgqVAmiHtVfjs0mpvN6Hlqm2a1W4uM3vFGjOJSsdbkpcOs4z5WgjW/gOun
uR1vVK+vbC1DYgfKZjyyaHWhsXKNGACVYRUpoo7BMxOMKR6YDgJVCKc1l8HzSlGhVrjatHxG0O6H
DYxXgYEug/sw1sBALX2tB/CjSh9btXm301aS9FLpz9WKnWQCCrAcvZ2IIgQcp30Be1a4FrHKC4q0
bLBmL65OMCzDtEAqYsuZAWTSeBQd9wuhF9L3SgrkX2itVmWM2CH9g0Y0SdJxXWfOc6WbofcqaafX
JFCzJNSdDcmSpBflbbhfah132tbG8jl03OiUs4w9EbGNmudkHPVTCUNT/OmbfCGhlqiAq7L55SpX
U1qIYu3j2FBrSQ4Q4PI/8njhlA1mi/ifELPe0pGpWdtA2Qzw/20TR/8bNObyEJPLZA03poksbj+X
xxzeYau5iBW0jzqitgDjjl2XdklPaZwGuwl0w3vlFTeRmdsjqWZNP8R+tE+8rTO5sIh4LXZLJxvR
Omxc/VMMOVQua+EH8gZmvSNhH+UHbtVo8J84kcABO2YggeOkIaNOjCc1tNBKsLdUZgUfJg4laO19
zuLU6cVN57pTyLSul/IezUx3JOcNdYxK63Cr70WXNgoxwFraSI0zUFTfFw48+ivXFhrCJAIywvTs
wlVkw7oiD9YG2Gdn7SgRIxPowpBrrfPEw0qdkpvsqpJVdr6LKW+CEKS8uF4GEk20CuMJzVu55QiD
PB9CmJk0LLBJTkFoVm4ujJnyDDxEM01DXPol+1SjmHDJbtAIOMLDTHDuFBJTLta4A+AWroZijX28
pcVfIEzvV6s/H4PrEPDgw0eXC+StXuUAEy/sB6geYgtNeFo3sADxdtSyDkzvoPzSvt5Z23yz2tmF
wMk3uv1wAsyri3vc7XPDTBNBHoK6YwiejEYduOeZVIt0MVPxECvvxEf4wfftUUfgCO9gFZWZkKSy
CB/i+cyDesb93iGLGq6iMWmV0SZqSDY9y+gzsk666lsLwEw8zT+A/AoySTuKLq959ZqNNTQRjCQk
TcZjojavl2jYZO9sP36XIcSo8Hdb9gwOEsvZWOuEw3A4rhZ6ayZyjRHaUm44Q3uL8hC1jhmdZJWR
+fFtwmedGUXlv54tHNpRJ6cXOfaHxriuO8fBajcuCVUmxYHMpK8ondT6hUyzlYoEBvrCmop2wN9O
pglv/QxjgA8fZe5HqCzYPnTKYNYSiJ2CI4B5N8JaEhfwxUB7jqcjE4hb6oSBgd+IznmXWSn3ViYo
guDDFYIeL1KNPziFbM+A/0+twfDJOhmXR5eP89/FdtzciMm8osfswmwJaKaGGJITsZvm66oIFG2c
Qo41EukbWK3QnJB/xWdJuLCLbwQ+fEUXvVLnkrm8HAvOC4ai2k+9pxeZsHWd6lpYLrFeFqV6AD9Z
ywzeosIhdshAJQWVziCMxevy2TwzFFa6EMaiRTHDf0mYf+02Pqflz93Y5OXm4/lY3gQY7/vp2tkp
LHAmDEFrRR3xFjDod2rTa3DwauAE83MXXkkDvFVo2J3tY4R3tP4SusuEYwAPm21LBIZ83C36kBoL
YCy9VyeyNXcwXh4ozaJprgAmlS47Rix/Z61CdYhyRykNp2Lw09cfNGX+9hipLseInc7xPL3YAC92
crsrqkmmoopQphQbCSVrUYApu16ED0hXmnj3Niwnqs2eJM6PZ7jjytuI6OqcH369Z45R3nL2OV2V
OTqaGqj4eedLVuoSBuC3buGit3I4598gVK6YE2YJw6QI0WxLyt3lMm2B9FTKBtngspFkGVdEx7Q2
ANlrbRc6pPqfooeS9eZiE9inF1tPnd3fi9/WsjvQxRf+/4nR+ofsBKPWUsty8zLhMwcwX1tFFHAl
HYy2BhRn566KXn1VMvBjw2bk556YZSEcF6+oEsWCJy33K4J1rUPkw8qUnZYl9to4gjgqN0REdbpD
/oWxkbpEHmkDpGLLSHu/PSO0mU1DdjetfiqQl+lwN8PHs9+VeSlSUx/mv/tQI7ir73+eDhC4rX83
d2uOM6dqOSDUtMOB7Whm0sYpFbucWG4DiQqOHqspU/9rmY/X6sAr6XYSXQkpisp6GdLgMVulhVH4
LetvWn0uXlsuAqB5XV4Pw1Tk3jzOmW3zhSjE74T+8UJFU52VwuK3j/oSH+Kyh0JYsBc9RhOS5Q6X
tHb/9omV2jmopz40eANg5R+ddP7Vr0v7p3cEXon5OdwI1yartXQs+h9SKJh0HLFbG4oXmrPRyLXw
a9mRitBXb7urUD2q4XTAVTYMh000ueOdqGQ3af41/y+CzhpGMB7w4fQAqKcxNL8xZvHd//Nni+SO
JhqMaQKOjrli28D/ToJv9QfViEPTCY6JfHm+4HjttL2l2XbXeEFbBOHB3n/dDeeR2dM339b2ImXq
cUaU3XnSAkqA8qMP3RkwaYAYm/IzuVrWe3rXjsQwaJ1SQ0tn6TmNLoPg163g+eSLHlmeMYx7CT1q
jkEIMNzErEiCqY0ARJvRWkW72tVDTzSsKy1Y8u5pe1aHQsmEGt7LigUAoHSO4eDeIr8d1xXUytgy
woty7TVAeVskhB46xF1ohWfEoCuomxIDUBRLczu0vNoROiFIIpMybMRZNUX2co8TaTt3jyS/XrOR
S+JlaLHTTk6kqRM4eNbSJl9WJNSsp7KhHdhEB1oJb1PDz9+7/BEbxcoG/JsIDa+XEmK2DGsd6Imc
iEG6x2sMPhTQcplaYULLuJWrAJmKTjzXWP+uOglGWVsNVy/Uj+RCtUhNBKe+O7PRb6xbmN5sjeUc
smTbZ0K74+93keFG+HQj3k8Nqcn6KCyJQY5TvL76cKmmzcGAHRFUpfmwFgcGUx+ZOlVhb3JPDjhg
1dED5n4EliuIP8RFEAbkwmcb5sl8GAh8XnHjZY7NvmDg7EG9XhKvlh9SBbQl8AJSoj/ILaWVU8u6
Vns5jRBF2QY8QVrVsW7jtq8ubzJRhMoEFlX3QzmqsUWP2OLQ0wEEg0ViyoAeDCKwsRHrwSP4awwp
oxeDhFrsVllGNs0pbdh/W229d0XBwX37nodlQsVMusxld8gTDydFLt82TTjKGoiCveiU7Y4cxDAr
u54jbzSJq+bZBUY+I3hGGanJ4h47rNr7PR0ljgD2xZ/EiHP+60nZp+Ky8qT+2+Xzymr7bTnv42Us
GppjwP3RdZoHRrGQxRzXLb/qgoV7SwaZh0STTNCd12FJ+0FdNem8FbZYqDkUu18fQQaUqxEg1h0x
cs/4uAjba25/V0xRi7BnlXZzzl0IWsRJw7zhHiizv67p3w/unzJ0PxqZ7sQNwViOXN/EvpLQqusn
BZLfcFn9qgGE0+J0+dDLCmrSrNz3vps7UUdNubBfnAneWWw2ayFvZ3Az13Wn8BqUu0ASbU7niCKI
pNmgeyBwImrR52mLfNXHhK2j1E3UOQNaUKdvKZ1vY6kGn2ZXUlVVS9B5IjeHGJ5KFrKxXNcA95Tq
/Kmn4sdxv+KwK+W6zkXrN/1tFEGYSndZ1BO0f65Kd2WzM8B9fMB2Wnn6LYHg5X3O5BwhvNgtjiro
HP/p9o38JfLAb8rzigTAFYtIK3USMBLgPlDL41OKu2SxegGqDNkq+xG0MXVNDym9in9bLnjliTPC
khfQp2jQhnc5lwHusbhSm4JA+QTlTSaDaBTJUW8VSaICiUiHwMq4PBwLWSJ458R7BE6Cq1xrrq3B
B6KcdEcrAu5Uu7g7ztiBwpCo9B8NzWs/uKMAPu/hcRPZlw8pVp5Rlthx8jkkP40+ogh0qQWXeZCo
9/3HSlhjwEYG3i1QNR7SxpxfGhUpbo4LpC8x2+6l5uUPcyYHBDwtKq1YagsGHYUn4VbtSaeezcER
six3oObex4Pc/wTw0ATG7CO+aBCzbxx7Ow/pyFuPCcTd2URYKkLlrmd5zELBtBq4jQGdg/mWSmTV
8OtVo51uMpZ3JMvPLDOMyuYOlntlGXO7Q4X85UBKo8UZClYb8M/4MA4TAWPBDFlHMb7ESvb+slkU
0Ku1ZJmxorUNPVtbJUPgI2ru2lmw1nyz4OJrlFa5x6poBjPv8L6fKhpk0WEheuJ3xwrG2WmkHd8E
KaRP4lM+9G35t2nr5s+sXrqQTJZ6j7u/qzr6JDf/GRwtHuT1hjOOOdzdKDg0U9CS0BodYIzq1PyZ
tyqheIIwgPmkKJso+470tyATfAB3MCSMYx16MSCPM3lFxP1aVnwzVydoIrAWBLtgd/QCu0mQvQ5d
4OcRsHU97ovfhFwnzgDUwK4imfYSWKNxw6iLP5EkRlItlCMfBMqYkoU+d99xQtYxdeF+fg3JXMz9
svTN1PGBgMaXDke0cOs+An/j4QXAsnRup9nsZ87/adlYPJxVmRQq0BZXsYvvpV1wS7C1wDlz58X3
8N0BbMa46zJSi9ZkegVAFOMuMVxA2eBc8fxRjpRnshXNy5mH+LeSHItQ19zqiy9U94ykKt/MPhQo
l2BQFTnpsjQ8TO3dXgFSDS2e77/Dskr+W1V16CtyJK7/33Fl2M1Q/qI2B+yK4JSHyWgzDx/5UDMz
3bbIjvLOC9bQS00Ds9Zl3ritkU582t/7jKgYODUn+KlZEbocxg+rLdEwXmoWa+2n6+uOwMXyfvOo
sgnAF2sSj/ER2XBwAs4zkSfrh+bgL8U8QdOxftrfoFh5L9oR8eBTRIC8PaetEkCKoI9EiO2Z92vS
ofc5n8uym/Kl/nMS/mxc7PEypwLErLrjFOsqaUtvCQ6PyFdJVjWVsvc5KMnQupOML98b00Is8lEB
OwnKiSGZL3QUwc4MKYNe9JpRXlqPteXLophuVz2Wx7Lxg9PHEmcQjfzPSBiWn9HI/9gsegC4Gwnn
q86qHxlUmiZE2OKpaLQV7ne8wk9Whob8R9jtKfNeUBULhxTrDY3ZIs0u4dyLWiXu0xp6l5Fz8sm2
mKGgL3lmC/Gpqrq8mJVshc2xPNzNXe82V4LqPKiYWAlzT0GgkbjYHJCqrPz3QWqI0u8UNU6dUwmH
bAx50UQ36XiJGDDS+T9dizK7lewtIIipu8oX8CyLZj38oyq50+7UqHaULKvqv3VRDJxnURA7OTbR
9Pw3JfM50syR7V8EgKysAHXiznarEFCab6nqr+8qdpYvwmpDZh+DV9AELG9a3hpDmhH4NyFpUhH5
PiOUkcZp0uOhz7KzRhlIyndyHtMUWSJiuEgPqFG72Uo70lzLPktm+vWOxLHrkcayzAIiMKFTeOck
v6R3hhTzRI2gN9RmmkdyHj2qhECh/bQ1SySgxyjtpxPbsRTF/GgSccRdg70kSILWD8N1Zroed9qE
e+87W+EDGolWa6AZeMJhCb0amFclPgWbv7HjWguCzumucJRO12z4kdf4+AR+fwV3NQHiLqmOpDYO
kHjf2mIihLVGIuh2bZB+qGKWixknFUEQyzLECvcF6sbF1WkOew1BuX5ABn3lGLevC0rmIcS/cz56
D3eW1UzeUAsI3UtZiGN2OhnDk09HM2hkmfLcEz07YUKnXaJ3AEUf7a5JMbBIBPHSNgiHLeLjdnBB
2mTx2sWeGHrg1T7EnzmcB11reY3n0ZKzOPA2OOYSGys2k1GWxlThNRUgeqxS6evubQ7p6KRs6ph9
Oiu8IGx+r9Fe3TKdtDamvqhHWMI1Vbnfqnnn4AyVdlO1Dqx8F3N6Vicw/l0mhtqa4ba9JI9dkzzN
0hHHYtuLLPSo6pmiSXXTVCZMp5jKmYdTQjPY+Qe0KkcUBn+jPxwViKp/BLSXJGvJrqSpIyTjfmY9
emYm7xhp6eh22S5cUL5AHSKws1LwHFUh8sdFKCZhB/hp0iTAU9ZJ2Rz3y07ThOlBkm5iP1Osehwk
sHxVeOPTl70AJrVmFgEFwms3M/5jd+SQMfivKi+Gg0hoJv24UQmh9TsTNbVfv8puaSpGFBdBNQiy
5rNLM9f+OF96Pujo8uGCSlny2l5aCDk3x42DBii437UXaVuXyCy4sdEy4sWVVSoKF2kdH3XNydg7
p1sFI92VDmwDM9GyaIGPp6mT8LAlSpyB8O6CL09UVKinVMDc0T21rAC9Z9DqjNb5zKIsQBiqliLU
RUdzHtwdVXEX+TJx+f1t3ZgFg8FhbgcOuWIjCSnsxDjXR2hsXfsDvQM93oZMdTRmxT/9Z0lQT+JI
DEZyD3wThxRkw8UymFW3UqkKZ6OJgWk4E5Mrfhi2WruUMa5W3ZFthRqkaQKZfF0pLHOIdKy2/K8q
5zY9KOepDshxf4NwrPdlzUhECNU5rcutggEMRa3kKPVwEOdbsrpQaneQOetY03wh4aDJCBjZaxrt
0htBdFu5PjqnW2yaXUvGo/RUvpy8GQpKms0YuD6UxD1xxalWdLrJiF5HrRnUdX1XRvZR4aS0mixw
xA8ozwLOXDXtgLlMKyeiuHpi7EM3v1dTGWbJkZ0p8CxIwatHzb3g942HQaQhTIwqUD5oAFEBzqYc
N7CZ9fsywnzgCcpXn8Nl+skIuzSXRTJldBhJ8kORoyoMdCLLt3RBTexYGn23xVQyvPJO+aZL9tnZ
sgRBKwcbQ53bCsgDrO3DyqQdjRlcD8e2JHcWHgUClSCojBAdojlJ0FGUix42QIbkZragNslyOtiX
333uX3orrYOEKT8vedvSCnIAm0N5ILjjqXgnxJpotq2QGJmExVKGjhAp773N9etAV/sgVoUGX4t/
iqyyFCtWiqrRQc9r50VjvwdDZTeQsOWJRfIoL31eZ2H2G7QwcWd4SCg3dUinA/15nlQ9iFqMqWbM
OgQPlLc8Y/oz3nE+uPpC+zQydF15Ex6xuvAxg0VSpZMrsnsmVkkWuu97lb9H5QDV1CIGavcKTS2d
//YdQucHc7SNfxzbdxeIUdT53BOo8QU0L/t7sBu9NSHe5Kc97wh+kiyLYj7dCeYiGS7NVFCDqxoH
DH3wgD/wbEbM9FRAZeOmGGIs3LKL4tkxXHlprTEko39lgI5xQzLuyxM4Fs0Kl88ugHa6gkpJ7QIN
clKkdklvO5FTd95vuOo7VnDw2U0bKHskRNVk3R/3ftafSkIQIvZQ8WIzussXa+NOKV+6YpvCicQ7
FtnWzKE0nHyiQY3WvB8b4DuP8IRp60QZxDPadXGIoOdTSaRtUS/o0n6ziJMFXp/yjW0nxwSrwECR
l35YNeIp2zr7Q34/141A095z7YkVLnCuVh4sB0hawSpSToUDAquEttCZzUGbZElN7wX54wcrsPrG
farkRNUB5XJlfxFd0RR2X99Dk0Wp8hxykg5vmGUJg0iInC/bcxspKfXgiPs3dHUBNHHQSqSRYZD2
OKftH//uA9bKiZdPdSCF9aS0O01eKOlbvX0yCvsaY6+YLx+kdclSB4JY8OHY8YRZQXFaaNnFldQx
IQs4ZmluZZeaLSAlcuY8nKmQbqa5QNTf9dURzKX5wS10J3rMwWWjwaoQ72RNogpE5OfQuFZBUXZy
HVR9M4E9JI3Fu2ED9sOGFutoLFRLnO/CUSOG7henGO0cX2jWnIu4Sj0gsY9aGeLB/rH8a6p04xk3
0f3zXO8FbR3hC0i8YffewDSkLg3wu1ZHjGBdfwlAjdF/AFnT+t2gB/DHUXi9uydG97PZyzcDYprP
0jvA2j/8caEu39cVjWCjlHkLEpwRLKrhXZ5aUKkkIbZOj7P8xETBwlORDvp8pgmTAS0nJriaaV3d
XGnFmp8G57fWo2wFakXbmolavSxmGgwi0ZhewPre6AH0pkdnbQgWBRLTttKm3FyrVl8adPJAKcz4
m8f7RdASEWOdgRmXfIR9IyQpQKBBACcI3HEMmsbEYzRCqCGYFWga9xLKv6WKDnSijFAOFhi76Eyj
AKK3X+N6LUqTZ3aNs0dqRwD4aPBDrvqbO10MV9Fvx33cBMqoQxVpWk7ygNgJi1AZSD8eTEEyaIrU
qiusSkhD0rHBRMIxq636OISmXf3xJcvNIGuS47JZxzLAHjaSqkY8c0yKfe7na/qQxjntkwdcDloS
Mz4SCymmWIDfuWHQ7IAckJwR+PmrQSRxHB92ysK1Dz6yP1TEIYVIlvYX6bJ0OaKAZSkdtG3k/6qb
/hG48U0sq4SRfPKO0qz/ixw35rPKtSe4nJb5Vl9zXWHxG57Q542OT/qpWRuwswQp5EMuL2YeC5Z6
MgNtZPgR6MwlpETHTP0NBxnKBdrGBT/r+G8fp963q3hChCi7eXJ1suim2z6jm001R77OrCdD57Is
oPXdJ6GRMQsgFzwDrY+d42TNdt4bcuJ5FXtk+SfsAVSyQ/y0QPB2yOUoPAjCQ6ePa8/lyuA7qRc4
fwBPMiHkqsuiwlSslqjq+bgvmcb7zkmjZH/MNGZgdQIg8mhS3B82m6qvGyLOQA2xTpPLH16XiEun
+tQ89/fp4MbuwVpapuUblw5NOsii5u0UYBtg9jWoUCx9nxeu4ABKxsHqg0qhHyn6uljnZ+HRDLFB
BGeVSLZr8NS1WT5UPxZf8AR812QOfRv0qWQ5yacPmkxBrSDHL1TZL22efUx2vteTGjuElwFATyYF
lOL8lU2UJmL89hNa6aRhXlmVl8QPDtIaKndoCu90gNlETPEOlMD/b2WB36D0EyefLNu2H73p45MM
ZGvUDpSl3puHUHBFnu374L54OJ7ODc7fJZVXvDbsHrffUfw9wvBspe01nHvIAFDKW5/LcIpMHqyc
2PlZGJWmgOTPFsyHkSGdZio8/Uv6odSMvEoOkkhYPVW1PXjl0rO+7fpS2CrsX5nUa/ausnKYqhiG
gLJerzPpRcm7+RKviETEe7WGkrHpm4koTYDDrqSLrINI3t00JnYxjwSogGGghUNtW6u9rayx5CDX
bCcxWM3IzKrBnM7QUyuKAv6ZxHHF4KZiG5V3MYKq6y2QKDDG/ni6LZPOug2bF3USUxnSxBN4aHMy
T4M6ike47FknSvkcLd4cpAMWKBL+rm/Nq4C64DC7l/oDZUqbpb2ge60GVUQAGJFt8868IHqeFm/p
StANlUoHyXx6jsY6cCuUJ28ktsp4WMP8zXgL6S9GvC/rfA2BVpfrbnJHZL/0pqLu5BDHF4uin5h1
G8Y8Tnfo7uCJ47KGANsP/64+5XRkDDx0ttobgHydLyJhdO34irlAk3aNvixS9N2vQD8JJLmrgBCA
wEPY0OmJRQNutFFbJiq5Zi+7wjfywawEuqBGMBHlyKAuLFCHX/e5nRmCbd2JNexYjfyvhwyWnA+h
3FZmvKDLzSfeb8sOoE/4w2HGNrARnp/k8PoU3mDcn4w/uAZWDMiH43s3+afKGd4o9k19v/Kd7YkP
M3O3kZ0BPvK2wWFmDqLhO1RB3Hbnjb22tl1/U3pWN58UAKLMovwTrZxdfxBbtZVr9B+2dRTnJZon
EIUMlwNGQDYKYgpeZAX2RUiPrzaGisX95Z/U6Dvx9EDD0q8yjlXeq/g090MYhistCeSzOVVOijmy
+wlaMOyOh7hEbgxLiqZt3KXS/1IUhdUjZFWZhkeREE1Xl4UGcXATQnOQs+IQ27WL5D15VGjaGo5T
rcilUzREQs5dl+2k4V5ZIpNGzG2bIpYTzaVvBwe5KJWm9bQn6Tzr2TSdGny8Xdp8jOzu9ncnr6aX
BKQjuBNOGer2PZPd1hgfhRErOzsudFxI6p4OR6GFHnUjRgEV5wbXHns6l5ifMORdDSCJlR4hvo2E
hKgXaMpbrBh44dlYMZV1eBqTb8gvZPBX7JcHIfmZxYiH2jEQVhMpSH3mWoKQhT0V3iQNYl5b4qhw
YcnFIwr6XcUIW1Q83ikBhxiZcQUtvtyMDNwtiPNtZqX6xinZaQsjYU5anSGqeA61HuHY5iOkBjoE
QBThsy/cfq4ewNSA4Jg5pWfrQZIi308MwMQ4YzwPIF1dIYTt5Kqv6oHeoycB1V1+XdtO3fzIdNND
uQEswY61+iQdRi8ov8GTxnUb2futMHtwxUdBVGfdzaS2/CzJT2kb1zqLf+2hhelTefsMBObVRify
pGga8oVfXuwoz/7yVTBqPa3mLzsNpLNx/bx14wEfe7QEGqolzT6/Uu0PVNOojI0y+e5MQkHWU+8m
4dywa5PhfitXn8kH5nF7AEM3huvjoWHAu5XiIA7ImpiVQUGy1HAN6iwsCO6+7WQN/Usoao+Rh90d
L26LL9XfqwEO5FUnXrzkhvDe/IJaLRnE9yMWYk93E6I4wWJjwaTog/hVtnSfSn4Yxrjg1XkCb2f0
64d5RvoMh+atm6jhgbSsg4JLUhPZmo32ZgB9nbTwDEyQLns01eutFMqs1LvrfHizjYj6oXRdiL81
0OLdQJ8kXa3a0LdwSjwb/wdZ4FqXsaojPM/7Em2Ew3wx0u7IAmfct71jYoOeuR2idOgSMmE/ddCL
L7FQ/aAdxjSLcaVegmQBdX9mNpvL5yCiYUl/aWz+kJDPGwcdyJioscSMIYjFKN2IoDxknyz5GT59
lt0dnjn0lqwOyCxPQ6Jd4DVkSTQoM9VRb870etgTLDk8xwIxC1k2oyucY2SQzUp1eILQgbge1/Je
LFBan2HdYJAvFYOqY6P3alGXJbaJjUKOYjw9YSpzH2TZQG2ZV68MuqXyAZn47eHD52tgbhC2MODm
OfA+Aagd1xTznod9E/eKREgodzddGyXdLrpgoQKdBhfxNel6fEDpyZ4SnevrA71FLM04zMcEUbgq
HctGD3Wc3YemskV0WviqiKvEuBy+oZheMjluXjKAcGP7fClrgZt9/nPHO5NOv781JsNp/ZvRqPvo
aYk2sHdlc5QavVFsZV1L/WU4o0Im5qMomPOoaqAlA4lTYzh3UiQYJvSR1a6kw3Dn2kDFy6Rb7BI4
tkovMDVLGwsOOEmMm+VKHeU9HGSIIk4y3Q83IsCqYkzM4+7boET/Zm11JOkPkzMlDeZckWZTP7CB
o+LQG+9UFCRnMuP5dZQbYsPIlbpO3FsIlG2QImHuDCfIQl1FwCfWeEE13/5xFhESpCTcQ3XU6fWE
QxwMX+hh759lvfEV602ibtcSJ1njIfoxIPQBjr0BkK3tjhBotDDqN0RKmjkPsb3YAFPwgfNCSxB7
Br+PXfejM+/WKsJZdBDVtDAKiW9KxhmWRvXV5K0u5R7fwZHH9jTRYwyTPOBh6n0ggfCLBFMbBXK4
4pw6I8n3PqNaKvCl9mpOFuugc8af+QwXUkFR95mSBtQ33sqWARWqdT4JkrTp39h0ofqOU+KR0dc7
Z9SUGw1vRVCzArL3+eeKNY4XE8SgmmDYnetUHdECO++HdXbTWKpQGY78M9oPTSrKqiUPBQuELuhp
baB9+X0I2KzATf3dVf8xhlMltrSAZKStxrkfidVGVAUDVIN8HHd16AAp3OScDtus+9gqAD6Lpmz0
vcS904GTfJYrxyE5V6HkQ8JWdO4kKaAcSNWz95OUM/fjkyJYlDiwV53psYRSol3sMhvjM48XaR4l
FMY1RlnKqlv9BHtUiAT8HyM2bs8sfTeMIRLyVB1km3Him+RcZtxQq5pCC1G7F1TS4RPbtlkHAy2N
/KTopUQLjXiYcXA85HHg8Pt/5ZKeks6TKJReBmVHGoAccbLuvynokIAMi7rzNR0DNK3R+JHGvVXU
00BeGrXbP6Dg85oPC3/FIPfT2FDgBlfONE6LHyFFLHHRb3WP1hs364j7YpMZlTju0jlXM54o8nIN
aaha7BOCuFu7rqaQl1qHMvYEzdVneUX7oxuaLmcCTReD+oUTRTv3MNFLGt1uCXacqFLtm/+uPYs0
XBcdBfG/TQrLVnFsYdaDYtQ5v6jIYFzVFOJ0CZQgAxWL5D2u+XOpVl5xDAnWx2RLK4QM7GBj+QN/
8oKgsW+qbYWrjSB4p75Wz/6NbIHPNLDxUe0p+mYv3URpayjG+ur1RB6qSPrruudsHvdlWIdJvdht
6Ukl7ssnCKBGM6FeXKMcOIacE3A7+6B/lM0kYY5dLO9GGkVYfVdR7066OiV04hAJlh85HGwM0Dtx
OrnPrre/3PFeVcReshucv36bIyqqDRezd5vgWaqv9ARRFDJ+HoTWcyc6IgY9RR9hHH25Rv8gK8WO
/FMW4/4afK7f+5E5ZR3p+Z5z16RFqC5SzedR9qZadw5IcMgYcRpAyomaoVsA6f8XffvXhSA3x5rD
+7dmDdaWL/L/SoVHOYMg0H11wW/KjVeK1lDF2K8yo54Mh4uuRZN8Gbr6iDohc/w8LBmpeRNt4kzo
w3/KEDEPfdSXm0Ix56/9hYLhSqtExnJxoWi9g0E8vdDOtd0gcKw1tkAUii9yq0G5v5bVkx3bNlia
FAntroxjc6A6g60EK/77m8QXoPqeayRt9aSqsD6o3XQjmD5QFFvtmZF3p+wnDuisFia8ZqEcbdIl
k+E2BgisQ/0P1oX1nd9fqG8d13qXXPpGwmsdI2S1cD0hdvWkwDtRjQUhSXNPAA+Pk76IkiJip2JB
kbJL/dI0lfJOZr8sRRv/zv5RasFf+IIwtlMseNd4ewirknpEVc4Oru5haJArLJunkJXonOBViZLe
W80QRS151kb8dRiPc9rWK3xm+B932lw0eiAwzDSxGYhc9R5cuwMVGgbk3v7ULhFqNZBCwBzZrWjo
ydCon+Z3S8GYAjHYriY9/G62vxNOmAcFOwd4QOpAUtHNNB99YaN6Wvi8MFCjrZE9lNtmlXRLy5s4
D57gWQUEUw5ME1bTi9eWmha4De1P7vWbLF7+6/uq92oYV+k7K3HNxj24HtdBXAX8epLa4XocdSOD
e487/BANbEfJvHwgck6QHNpIZOyIVsdidTm5pNC1/q5Q71ewOtCISD2GrUuk51IhCzP+j9C76HWY
LIKs2mZ5Qh8iG8xrF/dzbZwv4yTFqq8nyOOiJElPtAbfZLYwFDc2v8UV+IXxDzgr0hAh/oCes6b8
/9FqH4pJ5ZrS5KsJVp0dmuteMjChiY+/cfrGAjGQHmx2aFcFvu1OlLm3E08JldetbpC0oK+83g+I
cwHzm3ItJJ7bKGRqsdRXe57u1AlOxpNV1TW2kGbSr5WueWTUPmjOEBOpbrCur/uttYxiHD/pgL1W
km+0idoNX7osdxL2Ec/HoqOTfibRES8E9vZXfJoypFPU8Z/bZGq9ZTxuwjT8WssvITI1l9HqS+Dr
50JNOYYLW0lClo1hDA1W9q2jy2vgwqpVIQeHxM/Ozv0YtrCFwE888sO8unBcMmQ2Z6xZY7yLGWdl
XSJ5YAlzNLR6YOLykpXrMPX8ySRvHY2HAn5BckY+tjCmbAAHDMh5fw/wV4sJrA3pAiYEFfEuf2tF
xSkQH/KLqlbiER6GjksPG2VEvtUx5BPymPeOvkaEKKFwHBlcm1Cu79B7UPIGxXAK6nGS6/dWWczv
kfk8J5Cgo6Olli1xA+VlD6vKXgFogkq+SLN9uzu1+C9K8dYfKEHiIKyPInSKkHOZ9C4XYRdhXRJp
IxcXoWQjHnNHGBYHYe4/jvXlDRqwl980Kd/zSPh5gVAO9WrVrlKAU/CMpLaizu3fr5vrVN0swQBy
tcvYVa1t6KWS83r9QYfRVYSQHDvDj8Umzz9sHPYzthVFnfbiq4qD3QJrgljQYYA+owI5W/AlkZuf
QvqGntu3Fm6AHNmBbWGEFarE40rzHVRM2cX/WWvKAhQYJiu3UqVjrXD3GAeGMts30V0qNVXzFk4+
3w8/mOE8XuEt6uJ0IjgT2ArhVRbuPzI9NfEQNAIQpzLLlz8n9br+r33lt78eb49xOUF6pllbIrhS
Q4qiWt3sGzZhNjDWnjsTNQAu4TBEK7CChg3QEa348eKOTJ8YOUoRCacjVQpCQF2E9ycpAEZmNfmi
bnjzMzTTNkdAoE1UVoI/QUL0uaT3hv/4ZrAXepcRqDd6bQvT+flhAgK3wXrnXHUNJVLmPUI+eb+F
9ExIWQZZXDJ6Vp5sQDP4Cg2sb5mSfwuDVwrkzzl6c9DPcGG/ciiORcHwXa52nTHk5sInhxON/yl3
cETwE09tptqt5tb4iNaPI7ET49SxAH1ygWkokF7xcWAOO8+QOFFluGjjZ3LSveBDA9Te5FSIKhFU
G3PeR3goyJyYWQDVnzPG9OHr26J7cMCeK11jwcJ4N9+u8XYrFIT4tRNIk3wq4WYcNLstzvayFNeH
aNnKbLaq6RTN7MEc1IDtqPf1TDqhEdKAIJOwjWnFuSIvfZBPUSPWAZVL2ZxAY16vLm6H9R5whLL6
cTfr3wKdfnaAEB3Jj1ZHb6S0wbvQebb71PRAoF7JNeQOEqog6e2dfwGoRFvgnjzZnAkN06stjNys
3oeeuTdExJnQIwKNnmrBfExQEGLl4BXzjPpKLw2Eue7wIEHjcDSmo4Z+tR5XWm7Fj1ukXdNgzf0g
pAmrkIN6OC4X/saPqb1tqTlvq0q/4lGO+eyCEkompgGpHr3UdUjcYFzUIABeygO3u9Y03cdA17Oo
aD23O0nXryzUoSLKCv20lIsIYK8o644t6CqoC4Wgb+6qiFRAMGPSp78gC60STnD22O78SCyipnB+
xHBfy3y1IQQVnmCG5QFTAc22EiPyNRxAdPqKZBIilFN2EkVrx8PT+iU5BKGYnRy5r+PlODr9rqbD
OksnPT+HalSrqoRamgwqnzB3L9QL4WOYqSUEHc2es+1HLkP+vUj/exq8r/+gbHa4ovG4D+kX6HJo
0IrM4b3iBYcwJEZb+DHpJap0KWRel98LqP4fVBWuv89I/kMNv0rmCYtqMq+syseQGBPR/yAhqHNY
d4zvYJGwns8H+mAJsX7eqK1MdeW7J/f1peQ4i0pqYmqjX81UI+JVMdW2yJRZT2evRKJ/2tdUsigk
hi7HXcImqVQQusZG0QHvLukB2YETLOsJDhmCx5WVMJ4ex4SNTtPJZQtWAUGC8Wagu/uwzqAp+DbA
l0NLkDZTpPed7jsQCxNmpzPWfM4/wMTKua/ZUFOgyBXFkJ2DHi2rX+1iFCqPQ9gCuNFfbo2bxSYe
/xvQ85yHQtNmgnCsOlgOvo6976pq9jXDIFgKmLz6P/gy/8wOC6HH0gg6WvIuMGGhSXc74tEMT6Ps
gzrvfCEDUpA0/CegneytNycbTc5JCEoMtH1BxZL2gchMGIxtnajJezWsflUlWxnENncIlKrzz/cC
1sSiN6MSjuI9fMHAw0PQRfG0lALr8E7xsO/o+krmcynLE7A6qlpFtFAW3GkmsGFJ4BafrGGtqCb6
z27vBdmMI7kge7WjINPkpP6KyZZMTZWdYjpWzcLG5RAkqATJLToFMFWZ4C85gT8uOJXlRwlulhdg
zShlRhSUh4PsSjt6tlYPOF9WfUC8GjuP/Fv4xqfN0ltqKba/OhzHbECFozkLSlQKWjMkMtSCJptR
vIKfFXZIUOVpHDMGCAoIoP6Vfc51XljfOzV8Laie5UkhqF8aE2sJXFaMJPAxHA44Ph4+6EyNu0pw
lpSskvOjYjHS0vj5ggjlRONkId7Lraka3lthTdv05rNBjxNkdvEkXl8MY3tnxbvRPtR0ca1WIcS8
Jc63y6xrBl+PwdeUDavTB3LI2NDMOLqrwwUyAAtgl+yINcR04J2P/Y6ATAlsqAkwEJSyvryjlhh+
p325+fa0sACjDxSlOOI36zacGmCfiBNfvz+/u4nq05sjeEvI36sLWjzOU79ZM45OYuapb0x6Axqt
ix5U3MVFNudyiptQtCIl5Z0nadqkhfEEFCjzd2y9YDiXQMDngtbn05iSe2dVg+LCIay8JZssJx6G
8mSQXArlSqniGql3mV2ocze/otuoOs1ivKlJQUN1NLK8zfZjP8NTimXa7ecce0Bo6972mU9c8R8r
oCfnuV3z5hfdCCn8oI5mXvjR9Q0t80uM2Bc5Hb1BcDm/yh7BE+F2F8k7JRzqV0YdkOMsUfE6Bd70
jcn4y8cHE1TfQUG3F39oiRFX3vUbp/8d/5TsYWFw5PtOtxQWmyVEMJ12RxguFepAfqsUMtnLkq4Q
J8ek60j0FZSD1gdz0P+Y1Vsq93vmhhdlYflC9Iq0jkGj/Y7yoU4wxiVjJEiFE2lDD66mSs17mvvT
jumv+kBtC1tZaSFInHZ/80OQ1aF4eXDkKP4eo8mCrxK3zVKsuYIkFF9E3oQcmSF+YynJfvCCDOoa
IoVk2SbziN1aiReqIzzeXpw7p/GmbjgVGbe0Mvz6+WIPhN6i4SS4JJb9T7qfLk+oebbQi2raqC8G
SKLn93Ctiki9oNRzvLRK4Lmm8HPqmu4V8tKY277vUFOF9GRhUHftZOS3BRKFEI7Q2I7VD6xijzXJ
dMlaAs56x9HrZneHT6kuIVCL66IZOtUrWVrvLCiGuXjijCWxv96npKnXRB5nuZhY3CkBFyxhkLxX
9sG/79LXua88N+YUxgXp5Y0NvpgNgMYlVU9sk+PJTGHNfs41OmkcLiMMAYFgEUTNwVXnnCMmbDuD
s5IxG7hTvuDAL1VoXNORCW+6nxUyIolmWjvnGanN6nDTpIQ784EU8XdPVsH6W9rE6zTDSKkiziOf
l8KKUdK3Dg8Otx57QpTkkBdf0cLKYCcijXEP4zYeuIrcITEz1twevadowX26DRhWRaLhewu6PUwa
CJ09Z8U7A1I7lkShAIq4nQf9fmrrNtkjq2EjP6p5CaR7CCBI+xWLK84Q15MpMFBhB3gpIkpi/Fyh
PHjClgCavzUFXX2yqs6L4ozN7UkxEuhzkvBKg/mwbQlcSHIm+SBDt44MzU5zvvCZt8SURkdBHUP6
cpsx2PmwzyziAn8s1EuLvIrFO3Fg1y1Or3snZOCBy/HqsCP0pDPrB8Wf0v04nXu2ZnVHQRmd6eMi
2qioaDMkG93hZVnLAAjyZ6uUXNWc22NfbNvjOzQg7yDz70dQzgOUHpNcBd5FhNIpyayh1OMGGWsK
8l6mhv2Xudt+3c+YF46m6por52R7th0CrSJBmxXGGzGFZ3r10ve4jG3ciPhjjAbsA7pb24v+0aiV
2Lj6LsfvafzX6Cby/gYj1lBBSaUvS7smI/HtMl8d1FNLE1oMaPCIs1xZzTz8L8QWvGl9WVvqt9Bu
Wj0C1qPyBcUqQ1x5E3ER5r8qDEkAzcFxmHI3tV8tx9tB2isZMGWxG54gsB/ixki5wEG6FrBFHE62
NrCFHH8qt1IPtBx1tQp2BwMJW6JJ02GxqyHQCkv5IKehx/FmSuMdSi41NTWxoB54Yz8eXbmffQE1
JnjqBHV/cm3d3xF/iJt+gT/ryPqKLzkR6GCE3sZdkO5YW1D5WaxH8H7JbJDlYmLWe30Zkw7wCLhr
I0bc4xbhWZAC1uCzb8tp2HIk61MFZleqktdLOFn1fKC5UbJDfmTbikWzDn1hRU1mq8C3Gd3NE+U/
0w/HaLIAQih2iQ4pCdvZrbny/UwCkJWxqYwBRpRrN8k9ny768WiKZ3bAc8Eysp/6ZZKb8SbouShb
iVkegaZ1aEckvPMe3bmi+u8OuV2TJU4XCmayB6OSfY6zGj4V1EgriyzYvBXi6RUIhWapCYsqetqp
25lKlzhET+JGgBgy235d9NMgUq/qLzmgMIDr8jguH5ORon52VlvcDvLVgPYfHmFhoq/20nSTEUmA
ERWi82vdO2EZStW2qqygDweoNXAH1bHLbN+zV+NCpMlupJWJCfbd6IXJP6f5xEhbRteSLhHXjvu5
7PRPG4BDOjuJAaNMh6NJFet+fazlL8iUnsyK/qh8RrTRDIo6i79wJsz/HMmWxYakfjCWuejtDyIN
RUMxsJeNYfH8Mob0L3y8Qqhnq3iEhDI5GbMm5HhxqWl9slSl+Gs+/H76sMqvTY0m4RLickNeRVgO
RRLI57zE8eLuMcIBX/pvxgL4LDF/B+dnu0/oL5GZwoTpDWvlueQ4ke+ZSGyY34plSjDJ8Khm6u0t
5zyVYAs9JnlQOjaQa0Ol2Ps8ed5Jvn5rds/2azmXaBFwIrflEU+w2rXXRjibujybylgwLqIn5oMi
5Cb1vXPtqs5UY6uI+O60z9Xm0KjGs2bmJAdpfBBdFNfQkg7c6AD7GnPHRP/XXFL+G9gU/0Ztvinx
UeTNV+Xfhx0BqHTCS8nWMZ38fmLcufAFW3VCbqPUJZJ4G0LVR4cnf+K/1E3nEhgKoo0iSdlF+5K8
q+tjHo7UQs0y+d04c9TD5yN+ZYnSePjhnxLWCjntO+/bS+0obji/cBCKY9xxazjXNZ9XjZeitfkt
Mz6K0tvJb++ZS8ein83cBE6s/7bgDt5P1gY8J+FmyLMOQ9n2D9Pi6uYgUjzMa8+iZ3AkrpHWtSSe
DFV3/Av0+jWeLQeDoWw5icTA5r2p3w9A0TII7rEisWgKDjvd+PdF9vTwlXgX4s4HMwwQPiGD+MsW
M5BF1sgGHXXgfGwKpm038VGcUW3WFL+oh/WHH1UgRbUzmzIQUjQKSJG0zGEbOAcsSWuz4jy6fzh7
kwJEy5BL6sR/EK6JivEHlNSUxuMit/SLrXFs/0aX45ZcmByBghtfkD080nXu9XRMjBKUZA3UweP8
cC4lRbou5CPsCvhGX1i0Lkl3L143QJJLxacd1l04Pmh/8QHDsNO0AUgcBFVSX0pc1dmX6fblq7ao
7rjSol3MLaKTRegwC9OqPz82RCrZyRHEU04anc/+px/B+m5iGylveQCud4wEfMDi4ho9OyLxLwOA
LO4NBLdXr+N0avhdONZoiEmicsAqS3z2qxjHHhg5eZIUvAO1BN8lXmtasH7k3Atnrwo4oKZtSNR/
OUsLzOLZxQpEqYURrpoF0f4u3S5xsz1T/Fe/Hvr7s0IEhd5aDvw9jLDzirflQ4H79cgYDwQJ1J7P
vk8eeSCF/X3Ey0Q+IeovWPplBTNEr9hCiH3IvBOcTEJOs8zlbukelcCjf5IDiki1quv4rMXypJaH
tS4J+D4OaO4WDhCarESA+Vw5FKNF4ragY++cyw1L2sSsXTacD/MjP1klZTVLIPh/9UO5ZgTLxl89
l0CmJVkOX5gxNRKWX1D9rY9yn9+1BMwLSiMSNryGWrNGYBl4w5WHmRpvnqwGopIPr+WENell3CfR
sDZQ2qWHRXmyMbhBNYXAbkcjIJPOcTL9XMTG0yg1YgRA1WUB7GCbMG9KZ8TXjtw/Ud2WoJpc6Kfe
oX2i3m1UKzSZP6n+06ydkZyijfgY0thgiqllNnnV2ycpyXBorhOjgZ6rajMLSZym8nSVacfKaXdr
AmFbcwR2M8ub15nARsbw5Sp5EQSWKu4vmQH/nnq/4C5DB8bdpbIwzuvy0jWG27lrQtZ2gQd4qLDi
5ZVUQpnA1+rNGY4JZdiRxaxCjBol+SEUJzzhTYLHQzQ/d8JVSGExgzX+LazSKi9hScbjwJQKVCi9
R2t/r7OeOpEZPJD9BmDSuh3wrvkeuGStnHgRwLu4R6o7TxuIbCEJUafISGqlxx10mPZ2NFoAUM+k
vdOwarTNi7ClWFROhaJISUB4CNOIP4ZvsxbNdpkwBx8eGbi2i73XfvLnaGM98n4xslwrymPd3+c2
NfHaBKIbuc8/8zl8R18JRpRw+Fyn6gwImqtjkPFTM8rhX0Hp0QwORkGnoFigkq4F2XgL36Lm3Zmn
GSd0QqqHirs5Sv9dnAcwq+XCE5zSLwZPHp3zSqIvsLyc+n4pxVHTw3Ejid+Aqysqatox+2CQ+gxp
+EWXkHfOvu9pBcTa2epN+eAjKlDQ78c6C2Z9JYu7VOqUA02Zq6zkrzU1nBWNzUBts1yQ16KsbyKO
1H3LtAu6d9/E39GEK0xhrC7sFy6va7esdWTrHjE+FROGVWFLqqMbXZUecpABF1Bynbo+bIDFUE+L
e1yNRvTJ5E8gX1bAVUIP+YifYglqSyt9gbSBm38GqrkSXv6WWO0qTls6QWmRIs3mdOrByUJSAkrd
byZGVwu3ImnMZabrK7GXI02+oOqxhGs+kkDMXyxnhQnfKpl0liU8n3O2GgIO+Lsym3yd5G5IuquV
/kat53GJ9n+ExWOwROTr5MnCtXOwdPaZBBKRjIwSGJAdfk3zATsPsq6bLkcQptiZJ5QNxa+Lzc/O
j8Ttwq4CT1cXDD0XkI5Vd1uQY8Z95o1mOeBzbd0q8WEYRbGnIafQMueGE0zINSO65TyIzCeDfFAy
bgkVk328DsTGIuEgvEjI5VJ9+h42OSMy+QG7Q38d2qhCcYlCXHPo9A/dZvuvvy0G0ITT4POWZ3WF
KPAH/tyNVXKJXQe/np/YinJm3Y3c04tzoNZgBnEaX/XiRU11zLAeL5mmTNG6FA3ulN4eIjv0PVuB
6a/iBIwZW6ZpXabDhguenQg4cL3dB2CLpx3rGYxisZ/pc9R0wquxTt/w9hCuN7wtMuN1c6vT5mm2
hzNRhCD5/F/1KaHtnalFoY0Zg3eT6PQJ3Nsp00PgEzzCTuo655p4S33zFta2pt6fKr9Knp/DJud2
uHj34e3uOnx+3m5HOo/bBvcnSG6KKeeDbKrKr4lgXqjyMfd/l9BmC2hM3b58TgcLra/UMGQqDRZV
2yMFJJhU7JJWVs6Ltcy4Nxbho6xeAMAavFQXK3KwN/ZfHFklbZQEyg+PzqlUiRI846fJKC5p7OnV
/BbcfNN+AVs9pZzyfHK0E1hs/XSGhocqey/vZT0QiVj1FU12AYt7N7IATKo+fwMDrMk8ty2FB3lL
qJ4b7MuXfYoB+/zdPP8Nphdsct3IBilCh8sPjIv/oH/cPvJHKK88X4gBuFMnb31gWKhaFGz+nrqs
0bckazDS4R1YpH+/mitkdUvOLOHRqSwpLfL3A+mf0M1gnzPnc8mTirRXpo59ORtGickO5rJLqJVf
Y43K/sP5eY6APUrjLCamyoF7gSeDzW4w4NjrhYMnJ9xNdzmhTfe5nRo2qXQqRPBEwushwRbjptwp
ynhpjA/7ww5yktoMa3i4f1WfSljCOB9qowjhGsYj8u6qaeFMXBF31bB7W+ndqAEYns+blNjl+Fkl
Osl35fh4HzfqcToI+n+AjjYrFOdx/4iAmukOavf9gNTNecTJo1hcNBkTNoCAEfuc8dYJSGKD4zUs
DqYFbyn9Nt/+sxQ0lGelj0qvcrN7eKe83pXepX2Lvi8Jt8jtyqGlDvzxgUr2v740k7fphRg07mMS
tZ+m1mZ4wzBJcYQdTH578KApjdPfIYdVMzwt9Y+vTkV4CgwdSNDYBtyXEeqTnIGDnf+ZNhr4Dc2p
onUeYS6FS4F1E16Tg10sO57c4uz9e6mdZc5xRViIv96nxmYVDgt6hfrC2Y87gkg0WxXFFiSCjNL9
sD0GUy9MVREenkArwQXGnTrfMQrmNDgBo3D7cNnDCZobMP6I4W2htKVnYUkkwMrV+WIWHJ+AIV8p
7jLWXTjfULnzP20nmhe4auHAIcDGuHi/Qxp0MHgzFDXoZj2K8JYH/Wnn/GRd3mFFX1i1Jd0Vr5d4
kaxMlaPRnxtBCmFvzWTlUthsu1fvbTPfThGj00pmxGhmYr2PBhdYH1heaAF4+t7F5JtxLJw1T+r8
+LdEM4yDt2U6QGwZfIqs0f9y4VY7RsI7a78qJ5jn5s+YuETWIzR51vie77hwmPgmAxVUwBL8ykSk
93K1rTHbcAqSjieg2iDcTkXFmhsswS+ztBPOH5Hs/9xtmRJPNP50+cuW+2c62rf/Ij/yZOIJIeqz
k6RwZEUQ1Ug3CKlGFOBh4LGTxitjZ0uiPb8NsAbXWV+kERCYhvJ2rGmESt4C3fX9eCvaVh7Eh/5b
0CzrB7aBkX2Gge1KxKsFKv6M2iks5V19q71X3qXGbVoHMm9v7YlKiz/8E0J8q/1UzKuqmv2gzjYA
FnFGX8dyCvYOplndVptoebe3X9VE5mVrfxjZZsbdWL+c08YLG/cfq8gz62e8nT/eww/ERziTh6cp
5/1ogYc5gcPDVoTu2IaMDz78eVZM1nK3O0kkkr7K4YwCM+4nDynL/xVUVMdXJt0ucoiiwUdUhzyi
iGM8BkrIDRsQwRKy7ouRe7i5P0Av+esyo2DV2kbufaJvTcN1dt6FpBLYUGOo1FUzii6QXZ0PxaAQ
Kp1WFrjTIV0SZqNFGK77CJhFbfeX5AOUGx3PfRUBiC3+PzhxkblVdLV00iK5r+Y6N8If3n5w08Xj
e5Scr4XfahXGZ94AcAYgrN5dY1aEUCdtpl0cESFan0AkZkLmncKLL/m0db95PSFbYiXwsXMDyP52
ueRO6NjvgsMfv45Gxr4gw+KlKpUveU00kg9Mbp3LYsrIFGstpW0K8CWXDzoSpW7gaCOVXpIBhS/M
IfwUT1p7wCaCkAnKeiuUbb67zXoBmoj2jYicsBSQlEd8EjDqWTq+YGdOFGmFKJL56RVN50UnoPpO
7kIKUrFfji67xuywbO6CpJ9tzO1GupH5OranrV/lgfr+6HoUODxxJLAyWRw9VlDfwlwthwE7nEI5
S6hsT0UrfdXY4Mt+L8nNZN0VQbvpi+CaXummeevohVfO0vgm4ddtUDuKKnvxoN7wziVF1sgIXVa5
V4ZxqL+gGbC5OAhDn3RzvTIt8mVFRIi62WiA3qkCJ8HxBhxdXXHzj1tX4r9s6AKlpff6c5757XzR
85ykHSi9dAa/PZjbYzuY7ElF8BWmen/p3Hb13TIKa3D3jIxfDnV3xpZhQqsBtWEm1Zc22nynTvFY
0bFFHGrShCkudwZsvXMeiMEnMAx+AH7hwH1iJG/QoPz8d8a3/4Wtd0scYT5XH/qGH676r9L19cZ0
48KKQfYJgXeJsuVafwgBqP34QtH++b/+0Bj4PIxH5UD4zV+ZdidwhKKhgLsDqbejtCkyc76KKvXG
l+9mEnitrxjmwhf9H0wXcx/LS+w9dX75i7DbbFI9xS1exKl5ySHa87ohnB+1TRLcCAIpINVyd+t0
VGYikyj7BbZDf23vPeyDYuMKQ8yltx1GV45gzKqt5yVxeiJmXnIThbvxRhuZEVo/0aylIquqbA9f
xh+rua1j8GC4/XiyV2A/Fu427/weVwdBG5gGwdgTwuTgW82qlbrLEtpKmhHl+h8/nal/iaK1ZNkq
+xUk5dR/bWirZloPg/ZsMqZ5/JscjG/rvnRhSP3OdZBPGS4nCarEyG08+Umog3/jtPqVrRP6jl2R
xjq/64XHHFcqadxLlPQK3VDbnyrj6m0HMxSRXEUQz2TqjoZlcP8zCrwqLYU+OtXzt8MPuw+Fbrid
cOzLUS+6GiA5j2P2udX9US9p/iyEfjUfvF0znOaBXAiFg6AAVUmVZaxvXtykiJXQzpR+gSHli3L8
spU7OukI5+JpYc2M4vuhwfMjdj+vDb51gS60eb3u/aD4RUoBQBb4ghRPQ0gGo2sj8Nyx0UZkuFmw
voYrW2NEuGsaRwnEAU0t05IG422db/LMucxbMHUj8bJJ1gTNkfqbYzfaeH2GhGdUlmhwhBeNOc0o
+quupW9Ac6dCHMlids0NW9pxleGOMrjDZfeKK6sgyYrzA8tH14mFtVJakeZqBw5S9f98U58Cqcij
xY4FkmWXuGMOBca/Z++5EaYNeF8p5RtK2WYhCzrUh0GD7Zt7Eo5/91pZHIjfyyZOxhfMYNnIUmdP
n7crNkHI258ylelsJlOURVEpVZAhHLZq4W9w6bW+wOhFMzPpgbQr6qYCkKXL/vfQYQadAtEZjA1B
qIsW6mLm0E1xYOeY+3rzFTrsQg+LDNmQ+xIXoX/eSC3zb2LqK5sBjn8tkqgwangbXokG7ICG5Vrp
mu1Kz1P2pm9tPBPRaEurDt37Atx3xZ6avAd8WKAPFSpDQab+wsPIp2nLeGebaCKBJ0w7oolLuio2
bNvw3ftmGtguTcwvIg1f4OACybFQXn9YtR+WVqMcdallKbKVCDCS8HCR3KvFHdkmu0ppsg/AU7PC
nVIpokM7uI8D3JrhbNXLEsBcGsQpzI0PW6kEgmuAKk9lTg2fSQPNKj3D/8Rdjw+Rw92Bm0x6nq/k
sF00ao62ouiEpiEBL0B1fOYOfIgANgJDo088LflhoKoBdD7EIcOBac+A2qGT3EynjG5o245MYSgN
vIjBPZtUISPAxyOf0qixcJz5rLo0OgOau3Xnb98nQ9GU5sJndKh68SvBmeUPz+D+RN51QDYwT/Nv
eD3kT6MnQUtXcnAE1HlsQE3P18A6OI/O1j1MdE/591WIbe7Y6X3ukfl2+hbFSIEV57qK/fI5tvFB
XWbWe4qIsoRDVqEIuK6MjvVbzDLunSAY8PwJW1GD/xJtZkTWqBwRMxaIPvI1Osp+mX7CxZZYsYdI
EG2GBPoFBZ3+2cmwy4ug7491m61GKwFWoTmXBeL64E0g9WkjHU7QeFVvxhAKfI5A+40R9XuBMQVo
GZ0caSDya5JVUOB/ztHAZ58V3L1k5vAbUE5UW7vSJd74qw8Ph2fU4TC0P5oNKUfDId2tA82XjXCd
OH6pYQSf4XvMNE7Ei8VB2YvBGwmvH64f3VsxgZBF51ViI0X1Nh4NHJrJNl4T19hjaSxSAxh3oxU5
2au+VX4fxk2XKJN4gvhfzmoFQQw3cgeETpWQ15H9aTlivIZzJTuuqXmMtC67rBnxj3MF8cRX+EMd
FTcahUZUkLfp0SNliyqy2T5fYHao5CtFhowzoH2HTBIt7XeL8i4IW1C8boTXJBerU/XIftLWUFRy
9poGczPypLqNTQbO2i0UcGXx5kTlC0872i8T3pKcsbGALFRJd++VOjwCZWM/atIhOJ26dxwyHtZv
GL0fDL1SMCwMbkWsYrz3ZvcedLX4Eqfis2kR+XkcfTOBf5RaRrh786wnywptCmEGXeHAxzYf0GnU
DwRytSrVYxSG3BMZbKaqIxg4UjOXAlbi6fQ85wBOP9hbs4Tny5qwbSwObg/vqmNjPWXazHxaK0G+
CHe6Gfbc8bhG4G3PH5nlRFZ28sKL6rmrwkgQ6OeYsqWfuJI85VxTj1K2NkfQ2FmP0y52aw3njYW3
ppdrW3GSmgWxMeTL/z+jlIOzzHG0TnJBI0dKDhP7o1ixupVL54XlGYF7xwBw0Fl5S8yGT4BTMG9D
lxfqkwaEWCNH5cbSwY1KvzBYQn4S6lSK0Rfvl5qSJxQtM6K8RlHwTlZrdYYNv5rMppHlGTZ0YqMX
rPgh15VBC+kg/DpOU/X5KzjTouYq03ZOsQrExoc36uRxtXrukCbvRrRb9LiiTgEFJD1znlZp7xVA
8BJ9mx8pJVCcNlR01mbQmRieDbNbxi1upqV5zX4MlJgKEcljFukWWzQKA6kKQVI+GoSv4sydFCaB
vV31V8ehStGKYE0+z2IxYXBTBP142oI6Q3eGaxlfPVmpXAtkyzbpoTMBQJl6YQP1UXo+1QiaAoe0
8A4oqtrYRyQqVScgCFFWkCjEZ+Uz1eNpnfe9ZC4gSsZkFWyNIiff6/p63XtFSI+taF18u3OPujTB
lMlPapOAIjYfzCl9JbL2pUpwNvKSpPRLKmjXLMhzjrlGtOOof3UI3bUpejCHsWKvkCqkKFgZOzk9
X5GH22KSfGsIPK5VSwvEQ1Vvet1QkkPf+Z4a1/ZjTHB4MwxmY/nvpYcHfEFrxYJJt/PycFcllypV
O/GVOSeal+iU32C0HRQOu2IMm7hKN9CHu0KqrrWUqJX1L4rFxiqHwJYrPhnbM3mTZKCkWMt86CHD
Iw7DZd+b6/bMhmVQO/IwnKRuHlFfVG6VXYpIGBu2DdNyERZBMhd1fU6RzFgXBVujJMQIsoRHniyD
abm0myhjfcNs9KmJcJh+fgSTH4GrlDe78TLO6B7qUjIsvnPibBYumCkzioyyM0mqCKSEejDuMVlT
UHRToYvC5c3VQI4fK22sboGO4muKo4MSuYhOzUzAJf5NsU9bk579In0kNfcAhP25jfL9b3ycdLZI
K1ohkW8MyC+IYn15qHY0b6TKZQTkMbd+qkvwAwrskZe+Qwn4d/Zht1euoaoJzP9iqEN6aogOM7aK
lfiKUFtWSOyFwdgq+FvPSvlwpASzf4poTc17EPAjKdEpx4bDTAr/rdkv6V+E3PEhTg8U7wRnRplP
E5PnEbqZNAXVaLl4WSgzg9Ckgu8utxlqtk9sagajQBKtXHT0xVQ+Lak5DHF5Vt/yf61VHlJ0D/CO
hOOeiAEr5PpLx/7PhimUI0KES+HKq0WmFx84MqNJwjwraWlpQf/9DqbFJBUW/XD1Hiz00zawa1Bu
hsHwnpzrx4Jw5Eh0yyLCCq9H/g44ByW2SU8LqzbZ2pfNPZC3Nqf3oxVgzsRCUdcVdb+mFGhMx6jC
kWdLEvozt2KHoYJuPCfYZQ4//YWxDYKamwwuc1OH5wvGlBimBf6vgyhe72B+xNnT8MHhMtIXYUBf
n6FWymcxJJ/6XghSU1SOx3Nbyxrpol+K7dG1e5Jth0jo7d9AhMFUHo4+MNx9X1i3Iq8ZY06wJWFG
AsV7RTd8fC1yv8ty2Qh931JS5gR1qaaCvYooJwM3ZWjDFC9gGoR31oGKh0I9CKOapLKpmgOz5mRG
dM2LMQrpP4hjgSDwCx49+pBR4RDyAV/3TBi4LrPC15S4bsPD3x/GIv/Pe8MpWO0RTJ5WefN144FV
cS/BhRA+9qr7D3WhXKKBwUlhRZDoGB827V5MWZKv0EU3qR/vquiYx9bsaXbtkCbwm9dk7H49gSV5
Eh6CvcKXDLQ0zXo8EcmnJVExoQHDvIJOdno/OFVBhan/2r7bNQCZOdUXtKEHKrqw2siFK7YH/NfX
+MRxgy9N1MkLpiFyejcy0w/GuoaR7Ne6MGzVW/F/kMoV/qviheJGEWk1TpmO1/kqxnqPVD61e0Qo
RU+VaKk8i2j1mC7jFmMKW11pyvdnMgcEUvEKEreTDUCd5PHmbCSdAbv9EhV9Hj46CnTU7P0ghhv8
QPn4vnGyM8SrDxivSqYG9pkh5dzx6nqu5204TYR5XNRfw/RNlW8FDcEA+0z58SLY3A2uP4nPb7FC
a1l9l8A0Zi8Vxutp71JoZf6GnfSyXtZT1QuKaEPsXr6HSDzdLG1ZLiLt/BjcBxoCqwZwTqwiIYt4
x2MKsXGgsbBYnM7tQtSCU8357/Vg6KCJL9aQabzIM35xoJs3l3VCniAbT/oHPUU1dHFjBdbmBkCc
fHJJdLsxpamzltnBtGNWfVq5FywMDc5PR3DN0b2BwjuWB03P437dzwGNXPyToIYHLEmogNoOWLWg
RZxNcxJlMllGtAvnn66Pt46gqwo7XW1DPvApDEHcqpkjxBTmsozRTNBhwFD6/qEd/LbZpOoF/enN
wcHqs6YJ86XLPPn7oSBOkTTe5rpdGTgltFK9YSCN6WXUJygicJ5QCXvRlzR0Y8aAoCDOs3ilO6/c
6IUdj1spb8h2CeSgDKIWxZxfffm7bTfsfVkhjaCB2jQR6lOWRcKI9YaaECJ2hk7GuoFAmOqfKd/u
jwecQlHW1v0Mk+JGscACjWGjtOM/l5PhSN6o+hKjpuV/rss7hF/IRQyTMk7P/WBp1laKM7TaPB6G
TDii4+xtCsOVBjs0cDsxawRVmPj2XBa8aWVZ9v75gQIwILC/rW1YM17Lkt/vjNrKjDGozLogoVGI
BM0BwJ7dLJ7hwU1QUvQ0YjCBbH9nsT6xLyFjGaAEHPl1kd4asOFjonSvOOUadRDAdzhtyBd7Km+Q
rPcJRXqGuYwrbKhGzxNOzOTtveUTT26350cZ4gPb6P+BgByKyBtO0QtvYMNLR/7z/jwK43TKUJrD
I95W84wU3CVsJWbDo7CGEYYeUpGF5WI5DqqXDzcjjTvEmpRcZZS+dpxZnCrLOBC0oHCaPBCc1Ube
cq0h4MvgGGqbZ7NyNE/tPFnE7P+sbY7iwWwikXQMhZ3989CQPQllGweFWeWQ/t5xPCNsWK5xOkVW
4QCKfgMhsG83y2d9kXUyRSwUXmBbiVhFwrbrJitWFraxDg7hTi0EAkO6QObEP8zkX+pw/S3S0EhD
BzUNWOwNHmzdNVCkXh9i501wquNIbWrsJ3UFrSVfGXk7vc+V2xapV6oTC+kMmawVAHsbaFtKC1bB
/B5w9KzaJCfOwzw8JpZVSpSxHw06J8LF5HW69tVrno/OMGQTdbxQr6TVlpE3RTk3YoJkdAjaK23H
tm/iAikK9dAhkQ3T8roFDfRTUaUUfN36hrJklkYw9F2J7jMDoEml96f7rO2+ao1dLVLxBYcRf4ip
WxNfTs13CN4crdHR/iKeHPC3R28vx1xnxaEiiYjTa3HHVvyFc+xKNdoS5hghinsmbPRTWenFYmIg
3E1S3PT4z3y8uKYUG9VRuyPrrm6AVX60jdvgQXlXPHwgj9p53GmKpqCxJOmvIicnI3R1RvVkq1gD
m21ogVQnDM1w3Qo+vIjOVfgpzs73HiuuNDPCJqIOBMgTrXPeDYwvY8iR9EwpvKCcN4aJeJsA7b0Z
ou9n+q7ZDZ3ygGnx9xZ6X1i906a5JMAcMKR362rcF1g+Bjgo/R6NCSTpL7g00m3OruxntevAlres
zAGgwQEY4YHQ/4/zRGzZqh/N6H6sorOz2TBG4sNP0Olft7W7FUYvgDDldszyxOpadIDQ3Hlpr5Wu
Xj74d2P+6Y6DiC3EryR2JUngRSmeHSl1h1BaPAU5x3P++mh+hFtm/lbXECcHyi6zw9xS8E4uZ7eY
bX4O7oysfZ8oVXnlduwV8f7h1d5NwUxBzo1tfaz62ZcDHbn9ymYdsTx2KnOyCAnldYCqC1ra+tPG
Rxnm8FsjmB/0aGYF6LcnqCp+UZorHDMYUumYbqgKEpA0RWaVx95VD77a3Kc/rPLLfmJluuPA0LPS
CD6M2jDuXZukDJsBySHhTuFFfEpGw2F5i3JRaV/Nng3hwiB5pkQR7F4mUb/+s99PCyfiHJgCfLmP
7YVlsXGmCtTTDefnB/7zDSOsoBYO9Uj7CWgOo9MEdyx3+ttQmAcDlT2vlsOfy2/41vVToWsey87F
uEutmNzAyPOo5g+g4xyjYunfLzBmnQFB6q1modvpEBfDaWo8PDLzus7SRgT2lWv8mkIt4fZhw5Di
JVR3DRbKJKPx0nzQIUNtRCtGIOwPAdWzbDxTRrL8hUEy/BJWUvMJuaHxtTVy4+uDEozR1lzBw4y3
3fpaDtHYz1nf639TspX/YGXPWH3RdTiAz7kulG7GM4e2ccauAgSc/h4Dg+lgGCR8nCT6POxH1nEV
t5GgrAnycQ2DIZMqPOwCEyUeR+HRf4FXIsm1I6R/DisH1vSLyMhSBeOKcJ+4mpqUvqria52ELXg7
ddiMCA1T9GSjzWuaGuo3yu/1ph4P6K/KzUTeHc4N748qZdLryfFGmKwB97WQ/T8a2GuYMeFNrlf8
KjPGAIpFdXSz0y9yDG8uuEJYKXcye3XVUMhq35lXUUQDoAhLUSKFH1eUrbBvJ1L4HNcm62r5uce3
10rYHkYgitKQrhFpzbZAUKp8TCtH5J+ecUd3oq+obIglT/4a5YgYWq7OiRdKkriREv9U/d59LepY
4088xTb8Vmz4A6DBOlpqr39GpoLp/7QDQNSdytrrRVYPha3/sM8St6fbh0Fjan3D2MzAsVe1QPO4
pqzEBhK/uhMvJEsMF+qNsKXxoOIyqtWSCwK0K/wdik1Xfr9vPoWBdO8jWgT8pQeOejfL/zg9PYP6
kkVH0V/3DZpPY4gPxi7PYb7gDZ3uJ0XWntLwDjlwy1/67ja9qABW90ylSWBlKrGkS/5bNvU9WJ2K
NnKT9nwRM0C8YEZ1sW6o/GY6t0wpX3r4kaWZxSrjq9GhZ1kEG5vpw2KZYEnCpky5FmqbZeMKijDD
f+yvrfeSqtZvscUY53ews+RjZt0ChrAI1hsqIm6XW363liLybkAwtSbXM1ZRnVyAtJCZYNJIfvwB
ils1UYv+ilBjXmMLTglPcKuvAO1502PzKF/Rs4JEgZvHMEogOivM6ykn02VUFzQmZyni8tc6s+E1
0HtNjTM9DoY7SJRDNNh7/7zUXGlI9Dr4p+MHJ8LWE3WtxiodTahmKm4+o6ZmeksLNXu2FYhldAuH
v2I979iRgvK4IZZHVJNoGsWpJBzvBgYVBlVAYWeqdhtyC4vTpmyyaklZ5PhSuhY6s2tXieAkiBA/
yzLKmUBlY9Mwj4BByRMev9RrmTg4yTbf7fcrfBjBt4EYEIb/1ZNUUQNwbHAB2DjteqXwOfpzu1/W
YudpIXYXdZvsOZ69ByhDVLa+2akpz679ueNvm/0+pb8Wd/lyoV4jSbioH40TaJpnoikLEhCwl6IO
dB7U7yoEV77HcSRuc0bprkdOgJP8Cn44Xtom49taiIxEXjJhMKsejoqKzrVrmRnrj4Iv8ZZaPggr
Hn4wf9B2louaiwY2XkLroZ2f5UHKEuoYbfyxPxvqtRCGD3Sn3woHdWI1CQoEeTpqNVrZAW4QHz7X
OIxVx+2EDTBfJs3TQfjlXxLnEpPcOXG4IBHRqLZNjwpKf2GK1yu21fRrmv8lVHiqLAt72juwUvZW
QSg7tucUAbMDUeZygDHH0hYpJs6EVzoshr1NzjX/BNRbYcMRfPGJS7ACVt1O0dqV78WA+65W2+lA
WsZLj1gMX4MyQY2yMne4yAjH7xKisJYxf1ajIGCc1j2AcX4OfPGV8Fvz872tcqDG0FDvQA9y6H0y
mL1KkwOXP8MQmP3WGl9jGqtbddIx8Jz0Oy0wK3uZDV0MHCE9UaaQUZ0ZP3ix9kGZDkHDndgOz7T+
+laqfoKJbG/hS9+gLVreuOiQV3TV9jdQf2mygIJ2aP4Y6DMOv7/3SfCCou1DhaPXt026wYhbUIXB
4f4GS4asJI75N+LbBcVB/p13eYWNs+LWSbv2B6JyJzWT9zRTQFKffpF96lLXTT1Z+l3nDkt4CdUE
gNwnpKtvB5FBHuMJOBIojqyCkZh2z3cnXFCftu4CNer0lFWYadob8uXNxn9sz0imsCWcgXi+vJqQ
b2cd59nWktqNDgOMFZ5/93x1gA8nvb6faFVgdXXS/Qcpn9ZLCICtPKb3iba80stpOL3kbx+K6i51
PE1rwyAuKjzUk/hkFOI2Srz2HSJkyyQerRw/CRQWeJAg2zZbkDOw3q1Kso50oM35pmwdcZVvQinF
01pzc1W7+tY5pJkmR4rwwmifDvds2wUvDjDaBRk+1HGuWDo5+vJKVUQ1t6edD33vRBhrnaMw15Wr
Q/eBHh70Ev0Q0Oc2/YzuAz/zG0ccOUPPWUHULBfu1apZMPQ0DzaMONaHk2LqwObtnv7WQYBInNW6
z4WUmMdS306B0ziPiV1tY2EMHIUhAl8SkEbEdEkCQT9Q9b3k4IRi2nKJ1nKtEeb/hpE1ROVzYR3y
ZlA+xNrFdN65CJGtUrRDrCwy15KCxtZOsA4owTppp/Db67fI/IA7b6BYouQ7SJi46g2/a5GWdvAC
R+mzo098ib9Kw6s9A2WbXyNz4MP35sc+JapZzhJxYryEOxPGxpFosYq5Nb+Ge2h61KoNPiPMvUBY
DPDP7cYP4njtaoZFBuAb2ZLFAvIXp3jey2O3lCOK7d/16Eh+3TdTVd4Z88sNFilMld/UVuoWkEpS
i8WpMzMW3yLTPXjZ3T7qh17NiP4JPzh7U05qLKsR1U3CLuZ8BgmDi6Ub5qm5UCKoG8ZYzigoVmkF
tBzEJfyx/3VhlwExOJCjKKQ1qBehXOh5GlNDrXD/B3Qoa+v6numGbiZZDeyPcDhDzb0rH5L5eGQG
j+nZJcW1oye2r+flf22DCA308CuaPX0Zp5gEfJ/bEUzZjrpu+XxnLAcvz2ZeENyFk6BRu4i2wmHZ
XOOtui4s1jrhMYvpC2XqxiVVXabAXq/kOyEGdig8Do3OeplnKmsyr7TaDjFuX2ZBLGYK7sjxtCp1
wK/R9qO9R1f4slEgeOUuPU06EolMi/K9NSiVyk7J2K6ifE41prLQ4gWXKrbcL3Thvu2UnvY8PyvR
BVq416UnUToEXLnNRRS4ihdqK0NwBoTNnLJHUxhJrFPEDAGI2Wo4phS/KvWX2bMDxPLHKwdOjaMI
Em7E+dzvXkwpq/gemJ4aerGbidRq52QfX4hwzliYhoQpIGsEyhIfME3efj0YnI0LwJ3tOzibrzS1
USree4U9OVZFRP3KoKQk2ymUZRykObCKw3oi7vySgdqhYwf1tR2qMsRN4/ynJiMO0B9mMwbWbtN4
fH/1jeS0m457T6ujKUGxlwbmkReBlwII7+Vin5fP3batFaaP03d1+PHMZloOkqzdY+A/J0mITwAR
LPHKF6FiIB4oVGQ4e0U1Nt9dkj+cWgNp5lnzCEMzt+fu0yo7v24lQqorqKYypQLgdj5c35sG+rB0
GJTnyle2r+cx40r0jfVGSgQwgW7K0UW1qLTAcX6GRP6MHg5TCMWi59QhPh0vnD7wmpRYCC3jEjN/
ijnl3CJK7wUnoc761rU+KMAsbmniHwMpkpJ1WKIgA8Ki70gKVEV8GknM3weLVx3lUjbiKPgV0fxh
d/mTps+y6aOamzDgzwaL3/DR/i466KX1RCsVXE+GykvueWMRCiKvEiGxtrnQG8EzaJN7SoIM5MZq
i3uR7lTYOe5UGlWsE/tAVf7O7PZYPh0UrPqqq+JDEtlIkThe1qsE5ckg4fYZEh8ssLL2hOdVbaXK
vhfX0d7flY89HfnmDa4xbu/hk1DcgVk44zd/KVyrQFo5+vuhu5a2E+9Jg09UPh0OBrrdpKBD98kK
4ppa6YA7PVQlOkACcblMQUzPw6GRQ+pPjrmpggjSQmlxMWqO009opt2G7C5VeawCsGZ1GD9KvVP2
5cLxdORz+7VHuAPYL6mYI9bf/z+Z62Fy3uM6Q7YQcr+Lhe65WMrjwFOm0xor5ZPx1JsI2h0eyITD
VupdLgd/jBBYzJ6RxZ2OTm87ZjxTbxCViv97f72sW9p6CkdRyidfw2J0EtEVFfFYlWG8xJwuNjlf
YUbaBRPXjGza/TStDch1h7j3EdOZA+FJ8E+8k1rBZFFzr3v9R20jrS2k56iUxZ4XRdYiYLerUfJx
0/MR2RFsDc7m8lNvw5nujFp4VvcPKOa8eIN4GniGqiBiOofgtRaGzsgwG8mz5whkiCKY+Al8q7Xu
IrBrkCRvDEYU3bxoqf1RZjSP23rXr8fKuI5zdA6eun0MoXghcjGZDwgvBG0iCn57k2IhJe48KAE9
kNYhKtKTJ5XWmZVQI/iKl2n+OM399vnFXYvJdJE2DXHmZleAXimzuGazKbTLLQRHad07ESMTIDRQ
V3anpNWuLZTZ/RkxCXHHkbZTcCha5pdzhmnGcq+7QdXfO0+LKk+sz6jNE+71Q7HsFpodXXpibpIX
RTMK11DS4yvXKkKGkjQNG4JsMkReoRwK4fRtqFfSaIPTBMNcz+etGOGEyz5zYzBuzsJwySyxIBv4
EsB2GNKeZv87JQRTGF+P5ZTYjCLp/bdaTUJDIwE/VTIzJvglDPQmIyngq2JhGwdLZboBtTAC9RB0
vy4aeBkttkY4FuJNu8b2axD0N0LHv9q7uS9Azu5NIrfXObXOSjYbjJnO0lZ9z9HGwP8QCfsZKAn6
e6+GuVqyhCGluKOEMQxzZqKkKeeTgukvXbIs7EphHirihWvTCyNCBdkviw536eMAOBDWXwF+cmZC
qKncETREjqYu95SpGhW4OAeY0I70WMpPx1kZX+Nmc0G+l6ve4b5sZb8UGsNuRbN27JdRNUjtCEdP
vdqduYvIpEXfFEtsB0ctai4FUq+kbZqkPfbh/ADDnR5eVFILB4ilncoNlFPrIr+dhWGZ+D8p5Z9z
6ZrAJsz/yN7KgF4ylh+ZajrL3baNGP7s93wFVkvl7Axt7hvkEFd1knyGqH8VBRYycLKFtTq4HEtX
/V0VKdsuTAlSTOTRec00knnw41PUjm64vRV4s7aiOlVWHrGe9m0HwIC4/2Kzl3dcEEFhQWKCeX/o
2IBpB3k1N5zxJbNG5/b7rPobnOzYHvXTvWs9hnKJ6g/pxcc7urngHz4hx8nFPTfYjnBRxuo5aYp5
ow7rfnYm3M190MH2JdlIxQ3XZYR4ilMa1gzA40z1H+1L3If5mYiBUr7gWWCUGpkOQ/ZAJShdc54A
7m8Aa3RvLeMuoPpN217lSrWhAYY0oVFHRAB38vxPrJ1hvCv0fOeyBd8uEZdBCPDpeo+rKmyia7RN
uJMMGyQnRcbG8AkL4D4X/i2wC1ZInCtqIQZo5vxQjEZCCL678WfoziHwj5zphXSSduVHELUn4//6
NhvKl47Arc5l9aRQKCCHUIaEfkaQ4dX3jERQGt4Vyq09qlIUmEEmszP9Dh0o9BIzhSOsr7ryigYf
zLqgCua9QYypXrUUvGyoF3MiZkTbvx3gsdfs111aQEH+yEcr23jg7Ay0TQn/r05IamB/BfC1aRzz
MOp0o9bDcHZWSKC0nbzwK02hOqF0WJrykdkIZbnXM0E3UkQ0KiLME3xKHXNzaH2i6Bocmm9/KTgO
OW/PvTWUKAtFXDJxAhFYzHTCT520C9G5U16GM4hHLOxg6gH1dUYYTVUuOshv6qLRNjAT+FHUoNYW
J7HqPOGMLEiaTFnEl9Dgnwi6m881H+NPi8vvKdB6ZMYDpUltgEVh4WQET3MOsN+V6uEK8uowN7wC
zV46bbQMKHDcE0z1OY2ge/enjILvbFhR4vmjukspTY1gammuNsF1UOOOiuhGi89lBdzX5sPPXIYr
3v/97TLjNeiRCfLmafihV8yqH4zVuz/isk1jT6+IwvKNDb6R0b020r+nh4ak8hKvz4T3Xjgztp3l
WzK5ybkMHMGiA/tmu/KOjH+tngQZW1f9Dd/d0CCydIrL8E8icz9qdCkRLAMPZqANDYdCcfQJdVow
Af8CCu9T741SH4iBPVTLuiLlsgEZT2sBiTPEmzH+shR3x3Doxzd+OlmK06uVAgGoIZ7qKmPbvCyx
tfEJ8fD0C9Ic4AKewAKo+ci8ZeL/KtAeGUq5NVwV60PDLB/ovL0rns2kAp7RZPAWtMO9Nes49zyq
ox3dNS+OakVbnBx20sl+tbstpwgGzPK/23J0vVqPUEJe2uWcyK58/UtDQqQVST1te2Xvvp2Yd1dg
vIqcvnVT1WGcnW+GY2UXgxO1Hd8sAUUwN2FTE03CBO+4m8C6bkNcLz6fZGli8AuYNM2LUs/KXK9l
Mzp0Tqoz7lYG2A3S6kcFccbicCgZ789LCaw2W59jBdnG7B1gjMnK60jeyOWMczUsTk95H/056mLL
hl+FpvqCvpYbS+e8fhUuHgg9cK4qJyJl1i16WYvpVdyzwjnhCm+m7uVR0Kf8VLVZwdMZ5zFLS+xb
OhTQ06Vg7AKQJ4muoQPqBu3g594ORcd+cZLk/e275d/XHrJKmHeceF+RlOT1U1QZz8KuszhGTcDv
5sZ4FGmitoozhBSTANL33iMYD9hD9IoJBfLQpDUCuMK8mhw6KZZIOMCmgxvIWVBih87ELU3ZpNHO
RVD0Z7MlzUZSk6xxfhX51eWPPFdavI9NrJ1FT/WZdJPgD/p5y7yMDb1PK9gTxM+Q708Euvxyqjvg
hRZ2mg/me/3H0u9lh69RW3m3WrhKLee94y76lfBW4Yp7vbdDJh/RHC9ObogFdn/QCod2KXpltvxe
UyPL0deGrPLK5MHalmENfsTGlnsySvgjHP04Zubr8D/V8Rz/hjgAU5AxyaZyXh33hHRJiDbuLbgW
3a3P3nTiftvTyNCpxQbI4huyHfKlFWXWhqf6MjQ0ZnHmf/Xm62yzasmMsWiQ4mSIMu1FjBBteVr9
tJkSzjsl+YfneQ63E07nV69QSwjf6N+PYbrVbRbOgTjT+3+Va21AhgaRAhErLce4tqlJ/YdQ2kkb
cfG36tlLet8k9QYBKhxFYQaadMBWC/MbH4RwsQFb1CWQO7ZlyYed9+wEdCxJIhBAGIQrvQXT8fOB
BXXoR6+i1fp5ZFuNpBRMmwr2bnCvp60V3E2rO/poVuUtmTYjnM/6nmYshPjXtJY6/RbPdGNypek4
LAQqZI1vm09f+PPArGl6zFQs+i8sUoaX29M+wFi3KUIrbCei3Q9rEWv3miqwA08uxynSrBKBzvph
5Hop/M9+QXIzCNDMcpvJSMmUnixtu1XpcvATGmXTB+7aw9uBsARWdN5q2leyAInM/1aLT76oAtG5
eR5RDCVp0MxoFZKbPRRQgDK6Gaz3H1TJBmcQgzF4vWvMmY3JVj0h9+O+pQ7PwyQ1d7LWrQGaELxw
EUJVDI5f8DHo169SZhlIKJgU9eEUm1ZPIHXPgS1EBEcz26V227b2HNDYmNu4MbBXT0WXG4OgEXGq
NJnx0po39cv18FF6FPW8VG+ADn2aaqZLhsKxzXYKjFn6LOuAgo7+ESNV0YpxwTiVDZXdM6ebBDmO
H/mxxGZYhKDNfuwwTjXsbTlZ6370cE6w7YhIrdV1TmQ5Wk0SQD6RU9MqV2Fis3M3c2Mpa/aosHuw
q81AzEvFCTmRmcZbX88dCOfJFMy0gxXD/64hDleVeuZwz0FRSnCtCgkORnp16GOyWuQaPj1JiieY
JvYUZn9efPdDWEUgxwMtGmYNwa1Mf2dPX/K+zrqfKE7ZXcOuusiekYBxx+1kwA29VIuj6gTTnKkx
iORkVutRGSlKiA65q5FrKF1z/9vMYWTqIo3Zm+BTbTSbHzKoIdDwaTsCEislUVxAausZSwNPxmcP
hyoVaQkFZiRHM3wXKPXgbmKdZ/h/eb9cR3wHN4x0jALIWeVxbyRK9BatwCsTuJOl0onsJ1zsIFPh
j0rdloUWe48tV4tdTBK5uckRNZ8UkVeQmg00GsUrBVye4KFMOlbkUm7w3jrgmih/TWKJCKKvmqnh
8rmL4wu1G7YyW5ZYNq43j7IP5UU9s0mcDoPKUUaOZIfmMy8bSlhyRHgcQCC7+bo4hTfbms1NxAEh
uWtrtcj7NtBAzPmavYUMnruenwR1jhLVgFxNpsMqWtWNfAELm9eUW8y2v1OHkSQS/uy+pFKx0WZe
4AycSVIQPziE5YRyvDUlwtit/YS+nqmytrwD3TnwsQYxOW1TGD6QpoObyTu5Z07mfD56AGmmQZIX
olwc8WnjLIU8qPDEH6mh/vS29lX8y0/6OTbLzJI20BwqaDsPYePjFhraYi3RqFYs478BsKeOmQDm
4lAVkHD/1+57hVkqE5CVbXtdetGpvEyEh0+yvwVI4tst4faNuULL5NSSkO3Zgaox2vKeFTNIN6RP
9QoB606ejwpTaALbsw6iGnwuidXfkCWtVtqspz2jdzFHSQrdRccnAq3gDGauOmAJYN3XZVLkU7n2
yHyvvdOjAgv4QoJ2p9X44IVPy7p2yx4m96Q/2xChd7Xr3CMU4zmxG4bF0t9iZtRmI3mH/RT1qdbm
Ewyv6HAH/hB6m6ElcSM7XKR41OkFV9ufJ6y3uEViDpcyOEQk5cQt4zMYLJFLqN7hLksbQyuzflnZ
LIfaz4xowilnLJQVQFg+t/OCgf8sInsOjNRPZwOWgE1NyqKAnanS2m3gSczlAbCsXdvqgqwYlaTv
0X3PoMfGyEBflRsAB+dHOQhE1LqnqEeL/6JWBsfXO8YZgR7iuCJRzcZxKeQM6nOT80WKVUWIwN4c
ETymSgUm1HS+tLdVgh4kq84SOQ6ibUqFdOyxVWm9EQT1i9snafe0Hi4ADGTwEb/3sOGIQ12aRL7o
zbUfXKgh1si6fUS/Yxkplzz46WT15tJ9vX11hj//5lh9i4XAHOLchGgbFZaNfPZHYMWQjBTAkYbJ
Ax1BiNGrR/ialqJAs8Dk5ZGtW1328kgUM6TOd8FJQy8wkCmxYB1zHCyPL6IPm314Y0/5ytUkVyyP
McJizJfHOTx+YBCE/9jN0J+styieNGoxamyJli37KZIASJcqE6gSAfsVBaVeAFVop1HzDDehybIV
1teAXp5l5RLbytZFQApuVwYdfW1yJtTCX2lb0VQ2EViGhwc/2I89jbz7GR++q9dXRAAtZaQaML07
brZY45C9pj0kxcepqT37raZMwMKAn+/4xVmDseuQOtdXdiz+S9D0EsStBxMPfo0a0fldMLZqdkPH
1k9JyFpbmtlwsDZE99/tOVhvqOXf1wIno/wlBq86IGeppztp+hH7gxdoaLhjOb9F7U/PgJZto7lo
m1Sj9eW1suJBeMT7qrTJ9FgncmI9EX61vmsLj1Iej1PxMOVD8OnAccmjoXHmdZFs8uEbL8EfZJHg
BwpgOztKu5xE4mE8xGuiO8conWMrKZckJRIpuG6p8vpJLHSiQLNAWRD1sNbhWoEiSgMh1sGUldag
i9Avf3gwA/l5eXsK4UcEpnhk3wpPcFLIWjB3rO+iApa84au236GXYeJxI8XWbCpUmbedTIFnmXZz
9c7ZQdot3ZaNeaoAiyaKhlGfC4L9XGHF0gcIzAuc2rib8QXFfwEJ6GQto+JYcA30AlHCArZTwjqc
2/wJ9yu9N74RhTMsajzkH9H327ea6ludg+q9Xr3fxhHvWNf2ZSPLVvp4z6egKZqQacbnyDLblg7x
zMv35jCJSDWbQzzb3MG48UHeqzqxSEc4uLxp+LybDMTPVh86DVagp9crxSJGem2ygpU9jrIdr5YS
nYOYrFHQI460TInSHhpFULrh1DrSc1n3pUiUqmKg9o2Z6Nbl4+QlK+NA3E495ImEt73559P6VBhC
lZpNU9axRGxpbFtEpnr5aF3DtzXHnlgh9Ej7HpIDSeLhHtb7kJ0adRPYvcrF68mOQ+7E/8NsC58e
3qVketkar4B5k91Hu+cKcT/z1nfcq4RtFiwU4t1xlu/Aj0fiDgG9qPF7xm/Xi3WhzNrGLM7jEeaW
EOV1DhH7TVsEKpnC+9wm/7TXSrGuypC+YpOooT7JVOKJrbMib/SxB13sk0aoTrjI4bc6v67E1d8u
nVoZKcz8eDpVqt7DFnJ2de1YdWrBNRYUXLXtd1CIWCShjJWM3+6qFhYq9MF5Ff1VCN3FOCsIdMmO
4i4vlbO0j3vaQKRpvgtVRIYALnDeSXrTY61kI/+qdj2zTjZMj3Cxi7PpO2GSln01p5dIA+qhMXe7
KzOWoC+CEla9sgCWkYB/KxS16k+la+KXIWHRd7m+oFzWNqFQcdA5Sh3gzOZB44uQReRo2zYcV2C3
iHxEdkELpZOWQ+D6DAwIEdpq3xDr+MzyX15VC7lkNM6oGwsNQbfBIIYIuoVWzyJwV1NfPcNmLVMd
YlJ454ASXxiFJj5S5WRHnYmt7N9h0/5IVVZf65Uh4TAWT2LkDaC8c/kL5dNvM4YtTke0Rapk7gNn
+hfBFeThZ/NtgA/4E23xQcNnOGd3YQZ4lFyu6bKGZcEHqO4VkA8MCL+BekVnHkN1JxOCTMa/VZ/3
E9rFbIdMKv5qr/gMngAtmvf5yVqXK0X/bRPGf4+7xkZ03Tv5DpvMmS9irBT/23QlfpQYbbeImwvY
NZtdfl6fpqAs82yxl2IST4Rj6hqDGwkSGLCm6TtQwFnE6kuu8aSvxuqB26RcGV1IuE8c0lLCrhLW
dAenE0AdvxLLHFUVsJ55SFekLewuqmqkLzdEQn5khmD2WvEUfGrs6M3LSaXYk4u7RoP6nDGZZ6Iu
J/rqvT1xEfD5lc9OKDKVMPFEY7Iwt7cbufmEy/xy02UY0AqAAFMiDcHoj/UMafbq/7mKQuwXewGs
47fAbBqM2s4IdreV0LYP4hq9WMv28ytqIkFEqwKiKt5zk8onkEC3wxlCbd5p9ipp49SpBE/KoUfd
NBnRXUKAVqyf8BYqcVME0AHLdh200WHFCSm0rN4c0067Y0DgZEVG+tcruNiNCVHy/+nTlETepuUH
Vy8SYjS8bnZQ7veuUxRQiJhYWlAF8iDVgyPqUyZF1lbQk6qD1TVVHNRPasDCGu56flANCk4Io05N
9kvmulptaiY5iHwakpE3FS0jo0xCRB3NxzhPWrt4KFzoQUUpgsUhPRbt26XNM1s8RqlJs8v6WCFC
QDvJXV25uBce4ExhutlwrGurws8Jig/gaa/t7oubpsbN+9EHBUR1GpHmnJudQWwQnAr0H504N6Qe
uq+aKe89xDg9TFa8T9i8ho+mBeRmMzosMQTOPUD8LSrKhhdGjksO3xdU1BrfbmupXjY5QH+J4+y2
bh+YRC25o6q+xaTqOzfgI9YtpK3G3MQd78c9Ns3c2jIPl/PJsZluZMdvAHLXXgQuy2jO7usB/hZ0
hA2NtkWuYP0Kj49McisYaNE3Lehvz9rTDU8A+zRcPZ8TgS3RjQe14g720YAMrLLaUeI5AUAIBBjs
2mamRgaJQcKtBbOOntCq3VejDDMWJge1C8Q8w3Fuo3U4kNvVCOLoFVcpcZSmipIU963ljGSTARNp
7GBBKSxqR+LnUFZG+jJcBq+/jCXFCFlZjiRkL9RQe0nXIajl6wN7RxeJZuYaPrES6FsNEiehAkeX
UcXH85FnCfzoaMW8F+y2QB+OJ8MCQNRTd2fWiO4bj1NiZVsXxKvC+mb8MyBGkWBjjLBGwORRhcgI
4IP7J9i1GtwX4AunrsfpVe1k0F7iWCGywMgToZapdAEPg+nsqCVvIWd1aaUzlyefyZgG9CwR7R21
j6xKXJUfRcVsOaN9FgJOPZSbB0ddLNRubLIv1Zy1XqNTQboxKkghjFRuVs3AkflbMCGm6qy8ZC0U
RVeNQEhFOHg94j0Q0l0Hie2Yh1k36CHyKkICGGtXQBkEEghHNn6gT1pAkTI6q+Ly3pZaVjq4CNOh
db2vLP/2lXhjME0fSq0bWym+x1LygXC9Tkc9wI3Y7cbxBvXFUeFOOev/tGeSInVRG/Xfy2KXqkZc
1q4cNlfdrQ0EV6khM8ER32amZ98+FYqwH99IYb3+hAECxTtzwjUf6RV2FAM0th3cg/B1RuLgVrdF
bkowhUMDFws+PpneoY0upI0VQTDyn//EZhbOPv4FlNaDkFkciVOxOCdaPz8tIRg7bHKegy46uSVn
8eq5BNLzW0fszT6L5FvHvcbFigFGGhN/ewEw2sq4NTaPExW6+XiB1iOvAAJMoe8d6j0xGoxhQ0E1
lZBpPgJ4EcCTnCJk0Rn5OvsphY3n33DKRr1sjNc5GqQI6Ij2syqaVHb00lhaGzC2BGKPeeTtjOiN
j/wz+qGYmzdhk3ECHciaAIqNKoBoSMdGuTQUJJfkRzV5ctkq67rxNEPORgBZ84JP/0Wu86scOPEU
F12RaAfr7xVGoYt1skClXj0SlCg7rZm8IWFMpGbINrzgI/fpULwNTAKDxyDH07BmUSZle9ulQjaL
ShisElPSBpn3aM71aY9bh/6YJTHwvrEcPiEfTtGnk5f+ocrbF/CNSmdWvDI2CDAqLhmC/wq2EJAl
Eu7XGAl1t5CsEf6GdJ/x22RB5o2rkA0GKaGMZnK0xlyQwqZuoIFnZr5wYvGlZzGCD0fBkQtruEkj
SmP2GT7bpSdVJcsAn7lPUJz4boxf2GkNJ+MeHga1a0+sD4XFObnMzmdSHifSYRAkxZSom+2PFFgt
0ZSR3aBtXDS4bnrAT4DVo0XWk9aVwxrK8nUy4J3X3wpgBb0LvKt9fvlrlZVhpggkU5OlhYVfGYyG
EWp0U7/Qt/dvEdhOYnCkDZFd3oAplOY0xQkJ/nZs3/fWzf9lFmEJ7hzUuyygq7AlbDLowYxD9c1a
3e09f05l++R6Ut2gs4JE/W9/JmFLzwP3DJ+xTZ4iXq5sxAY+JoBw3Yow/8Z/B8Z7WGc0NFbQ4ov+
zHmE3V/sZ84tzztIWT6wE+8tGCB/mt/7BIhds/FLdI0lY6+BhZEpaSaPEN9yrzUey5k9du/wiOBf
is8E6Aj1uEHV3SEYAr2uKsWlX97B4GE/MemOe0fukMjHdz24QW6cPBD52Z9E5ALoOglMPwVNIMwv
WTXN3rx9iy2D4fXN7dE6PP2m4frcvTsejjYvyU2vClimBCOYiCibNlMqnV/mAya7TzHjZEEbr4nj
1QwxvWnEWsRTwvZZmsapib0Con0iKutysfqDijchsyRlgfRPMcSq7ag8TvOh9N/EmoWpvI52o6Sc
i/IlEXwxQgHhwgLUoaP2k5qY+AmpzSNAfoKzBRCb5rxlUXJN5D5P3o6Et0CW3fWH59sOBXeUDriE
SemN340z0ZlHuTrfAsvS4ceMSiWCCfBARNQKHr61wB6W5LVLNZFxO31zFRuKDiX899bhBJRRArl1
GqFTvqxi5FUfhNj9rAaMh69K8U+Eh/fDbrvJvDoOAyOx5AQF6wUviyRDWZgp9Xb2xw+s6oFcmmWT
keZyu/o5M7MrH9oDItQJ6aoibGfl/OxQuSAs8OUmZ2d5cK+hbpvH96mItgNIOMAUYxUvmkfHPef1
A/WchpcgIJKK8sT8R7QAAIEKZ2x7UTyNcSsQikF6FpMficvU/JiODvqm/BEXvauvbfoxUj92Cs5U
DN0GZBHpEOeW+oVILdzE852KwJ801PQ0Gv/HD8QePifNQKVwgnFAm40o52DFG/GXMjkVAbpiKmk9
kfFWHhN2zIJQaSTrEXsuEusfKhT6Lo1+3rf91Cpldw1UPUb775afCdWFF8tJ2hiOWwBWCdbk8Iz1
wU6GsIRZR5yB8daJuDFY8MjPUUxUWsj0OT0y75N4Kh8j7o5DIKTHGefzk9ixJiq6QrxZI1sAGgbT
XpUrQumoAo04fH3IifmTPIhUNIxcS9oTXg0bQANgmBMwkyXqzOt+9cDIsRP0tYLL4bQBxRY09I6Q
WrZXt8pPONs+h/lY9/eUTRLVH46FdYeQEdMMPLb91wPbEXhVdQhGDaV0qH3oOiz6aSjyPkQsXkTU
EF0rAGrimb5AwnwWAXEIIoZvnNrTcE36/Mlgvi7ihjYI3oSN/fpB09Yd78nnnw21G/VCmpurgCGl
MDea50o6NCHLHFOcMqdodka1m1vGvOC9ZWGwJ1R2oK3MnWBAAoZQQGzSSlPXjv1iniIYJRU8n4ID
BF0NkCHQdK7CwR7aR6Rc/X4pW+KlXlwILNS3+33/ZUy5jhy0VfikicbB70/uDJiWN1WEpM8kWR85
s2zP20L5GoATUaFYlZO7IgRq3j+aU2dTu6/S0ttDGStqJ8QH0y94KhqY4WtHsiHszBG6VQdPYL5q
ECk8DvFVFcvSGIxUk/ejhvskpjWM4B6+JLvDEHxCxggvE52phFoEZVKsdKT9a83uf8V8ZKSt6Pi+
Bqxl/E4m/SLB+cgBjxL9HdYbSzstpIkyZhl+DP9UZVU0TBafsGgVvtF+HfocQRVanTg52bCa5Pk7
4vztOFlg+YQO18VPzlg5Ml7z1ltYGNF80qXGrAITVwp3OooPYayMocqGGLZo6hXpGSru9P3lp9hM
1TsdCwGWKvOxMVZrR9SW7WdIhiRC/uHGPyyMN/SbOblW24qHrY2Lv3qlcoQh8FxKkb9Th1noSNrb
5yJH1bvMo1RStf4kAp+mREoSuLBmzYHVMIcVblP1oj4rcmj//Oxpi9JAcl9jD6r2eKJlZdGJ7C9i
Yu+gOiWhs7wIQWbzzF9kCJkLHKh9w+/n6t7bKuwyA+nkHA2xbelarIByOj1V8Ufr2WLTEIYxjXo/
4yJr059FGOQs9d387jsfqZYobK7Pku9s8uMz8/cgoSEW4UIxUuibWchzi7bCJqPvFSb0qdRlt7+K
LOkvFgjQ3xEcZu8mM6fW++7DvEelMNnnK6vnXq6EgO9xjahcWaEp+M+vLb61XDG1g485NtT8TXbq
z0qipmlU80oBfiHUAofs6J7zkTxsxu60nr+dBFrMv0ry/On5yyu9Lw3qB5dDxZd8NMiAcYghboJI
nvouWNr+sw9wuIYR4F4eWi/GsSVA+fiwPvEGGiM5+stSvlF1odiL0cbzBr4Jzwjf1Hcq7m28mSam
KAekthDouRtcZmY/Hz+NZAlGY3W9SL9ArO8s6YEIT0f3t4U8RrpkpFrNXnIM4X1ShtS038LLqlUp
M6XcTNM91+7XBHiD++qoKJ2gKuWX7hxbQ2PFwkZV96KWJwmjd4FoDHn0Bl9s2Ighh8jGiJ1C+b1H
O1STDSbDJREgdzKXoJu+1cvIG9rYaQS+zCjzmDYj5lHNQxy7T4T1yvKWobetnZjPBrd6A7b6xiNa
GKRUrOeBGuvAr3+CTS2IyZQ5cGy2Ig3gz4jGq2aiXH6K/mZiOISWsOctDjlu2Sd3IKlBT9AlyVT8
9NyYt0HuBKvfBj18HhWKuFEFVm34Iz+IfhVejC2m9kvjaEmUTJ2Ll2QAw/52wLgKYt6o38h79onk
opuzvO0DRY0RKxnHCQW0YeE7v0oXysPd597BM/3ksRM7jtbAi1PVNnzwrkWyNixcPOMt4n7CykVJ
A4M2ypjA3uYxeJFzdDrDpBXphqR6+DJhUu28nKMf6KSqrP8hnEmauxvWQaKrkOKOoEosRD/CKxO7
fr5ZiOmnqr6kIrlXyOcVlC7O5TsFoH+H5uWHwfl37MwHQyEuafEooqeNbO3tF08Z/wMmiU+nmRjQ
37vC/YDsJra9vmSdqq7kLAjwovmF7GI5hnNzISP7MNMLG5VXGu/UVDiVZCa/HDQHxlMZ8oj5aBq6
3UQpB8NpUVdaRMWZVJAdy+31OOHH/01KYqugUcTb6onElgbcRpTzhn950rbTmUrmwBiFuUKuvtJ6
wsRStoFO4JwY7Lh5Bb/wj0jFkBbTji1P6r8TnsF9CiECZih48sFMtUZ5xOwARrDMnsvRlDez0sp/
dlgjnH2lIMxDrCPHXGaRUZnBA+wDrvwPiefuaWM64xLEzsI1mkNzAJwjWWp5TFmGAz/bE6Hr0lws
GGnA67hBNhwTAhtJ9bpC0IN9nYoOqtaz1R/P7n5Vxaq+WQGfJ0JHSRZhv3Na5jG0uwKeT/XTdWvY
RaBTcuMR+mxMHbWv3cMUIiafWI9ywu3fURI65MJh1fHjRKRmD3Ex64iPJqmWo3OhHTFbv2Sc9gzq
j2BkaK4LUYbw+mgf7nPUrq16rNgyMarpe0KCEk21GHZinT93ee/7DdG++nsO0gjyZfEBqMdgoxM9
M/ZGvRnmfGtTG3nvO4VHvS5T3OxDcVN14WZOdOs/y+WUUC+UM+6XfnjIVevB6xBhYeU9j+RXE0vp
QuEBB6gdrZpNUC8fjLOTWSLAgoGRVqy7P/xUpm3MUyMHxagNswDJcWPYSJjKHD47oYjwA40pErA+
WwFA0y/11v5bwFXpBAKcRqG5P3in/FZ4utkQLbJ2kv0aIw+pAZsZTm3ev7/hYp1y+d78VWPq7fGR
SMiKnzFwGeVZG/JIDYHOBWV2WCLiQBTkko7S/pN7ybtMaIjdgVSgY0Z2I7Iq5AiBM/BMflue2O5A
58emhROou40HysgbdjB31aW6xvLUj2b3TblfgFjNAfOtKROXok7yYPU+s8txU0RogEg6CdGjoHzO
DSPjA15EKUzJ0ptQIXNV0jwTdhk/HokUhtoc3gq+oyUrWqYfvHf5qA/Q9X1DG+FL5RHBfYBLOYfb
SYaN79obRTL7TBJ4O964pHPfYE8zY/l053B+tRFvSMyesTWpgrVxyyrfJxysDG6dxN2FFQW7GQmF
L8Ubj2UEb9blCSed1wkn35sduYNdLvz4naEFQdJLjjL2rkToCIbe/e6Z0kO3oZCumEDuHjzNwncq
f/ON3Afo/wafBUisY2X8JZSXMZTjPbWaQZgsEW9KfORCfV7boQxyJh3a8SB/zmNgn5q/KNTXGVse
rruFn2qtqQvslo/lWh8fUALiBQzSOeGta6Af6fp3KBGSS5LVqR1d5UvmwO/fIU8WE8DQLpla02H2
G6FQnEkd3MAhOadJXwgdX8qBiU4RT4GKbZCiDzDbqBnyPQ9ZY4qJk76nv6/sfmqLBe4tOE5K4yPg
o4Cw+KZHgSbsSlZitj6Y3PJj67ySdJNj+MeAnamDedBumrJ8DbSA8uC+B+qzJiyRvm87jXabiHkM
tUw83xsYytcGwJX/DI9uldxNO05oQhkjQk4ARWA8VpfUeKLOTdLXdMHI13NWzN3ruMGj4tbyh9cN
CBwbF3sjsEKg3BXklZ1HFESjXLSvpKtVAHAeKly8a7UIw79FM6ZWiq4LrkonYtqYVxPUwVrVkP8W
xi4U3oTu+FOzsYkeaJSlUPJO4ie4yTFxhV9BiV1phAs2/riphEgeYDgnINmJZANmuNwclcb6/Vfx
P5CLBntzlnDP3oBOA59ozePdFCaDTQETuOwyc8ct+gC5QlT1cZUfMT3SfjPek5CNfJbkVCCUsd9l
q4CR/QvA7EnnTUctpP10BR7n8mA8bcgYNQFNm7PNewUgSIBtijIAFwK/Til2Re4TjBpkfLbA+pMN
K4iP22BjiW/pfXkSHdc/vvfvEJCh1FCTXoW+6EKdm8whS3iM1rgMqwJN+bLmIH+mPGik4tnG9u0f
1yloE38igienTa3UoXNUrVfOCnd/uWgktsftrt8d5ELCOj6hj2e5sbAEOkY8s3MOvXseV09p25kB
vq+0yksIWqeqPNRFsNjmwsKZGuiTzMPyRpCtmS7yNmhGeB79BH93QqFZJtmLqQkFaXedLQOc+KvT
s8COKW4GOUKYrdjjUxlawPcRFLa9AgyTQ8esOHrYQOObACC8RM6edDzpdTr/jHPyoppiutmgrkCj
tVpHErYCr58V8M+sj8HFxKgrLt7yNY47obZxMOuBH+4765bZEFOLiBnu3UWDJgF3scYawGnVfjbu
Zas4UK4R6FnjL5jmjod8powzYnO+J86dUkPf+REPAm7qxY6CL3VAb4evSrTLcSkNevcx1SIIpLZu
obZVLpR7AYJRsCszhgH7WTLD3yAvqbvjK9OMUk9xP3tqaOqGbfRXqa18AAYXPE8Ux6JHdwJfvlIp
JUDHv/OLirdlatMiV5pvH9xPaPpb0jHI/iIfX8RcG4cKa4ssOhM95qZakCcDrCk9YG2iHR9tAQXu
bcqko+lRkkwPkUp8T5uQDHQ47+UOVD2JVXLNL4HsVzd7I3oSmML3Y6T8OOgZQ7aMOk+3ONvyuFjo
xSzKArJGoaDuOPYrHkyBDMo0EmC/iEHKklssTtaxRM4qNDaIs6f4Qym7PCfkkygwzJdyorTDVJAJ
Y8BOuwG06Wd2BYuQ+Jp1kk+qDWoColXH8d/jBdslTRrjndTNgcAlTwMc01v+bCPxF/YH9HRS7jlQ
IJf/xSESQj2l2J/SYGJffKcypBY7iQ3KcGudz6haftEImI7Blb2z318vRV2r3WIGhA/qotBY20Np
SkYUUNes/IragJZ9KADRxjEygxN0yQyiXHd7WZHuB59fHRxDEbBz0cWUvJbVpELMXyHM9ssNiO4q
XPSdGTQF5FZT6cqT8BJVskdv7CS4dvsrn3i4TA0+b85G1OmFNPi4MYC7gsRT4kxIQL08j/gtynC/
CRLcngOUG0AP9Q/0Xcrmkc6dKzm6u0oyByIO8MTJGp9tgyUvYx/yd2hF0jRDnJqIR97iM2OLlec/
o+8NU49tmc+u9SxEpjJmtutTj11tbVbfD43C/gICZwMBQG+R3ljYGCepXB/RwbgVDDYuFnmyclNq
U2jJQKMk9p+eegQbfFFnWBlgRl32eoxjH/WNtE7YP0dkoXMJc8j8uSk8/uMtqOaI05eBDgbW9U+0
hW3x0b1FTo9fHoxJBfCkSKgM/39fACty6aHa7lY7iEjQrsMwjboHnQtvC63j246PeA2MBmS3+oPp
r9TaPLW9cvHgQa18QUCz+z60WDNX78a7KlPP/tzyHAVG2NwFkdDatcWNwjsSb/dZ1pwDT/IZ7h5r
A/RiTDo8vv4KWKQTQUh2HeyB7MNs5P9yFl4fO8p7K2xYQr8Eyqo3QUhh9X9Gsz9admFd56QH+pxj
upCs3hKULmO0GV32KipVVwYH8wnIPrz4Y/ECKTIK9MLw+PP2fEhfLezvASzaczFK+7ZXJN53zppo
4+ZvgG+o02945tVSwxStk/+fkmXsP+btjuI70m/6572Yxio4a+nlvT4WPo+8ZH69+IfqFYkCEytM
kAN7nuUj09pdvCRdkXTazjRtW4x1rJFxhM5A9fkI4uT/Xztw+Y3OYZLD1/SXcP7LWJQcF/D2usqb
O4FgQ6ZGl8O55l0pJIsbLAXKqX5mrq90eCDRjtiYLRsyJjY8X6Bd6SgoWhwYsJU99PQHZkL72aPX
kKTt1tCgUKXZeM8lNQX0CIa3nvN9tfsLZMgqB8RT7t0NuRd6r+JdT66T8vhlGi9o40SbXAItAcN3
EZKSO6552SQAVw2rEAuxlQeRbdf6t+Kz0rJTS7ysw5KbXlrs7KZeYoUbJWecAkFkyY3WZpfG+KIQ
X8Wf+BhixXOfoIBxAoPVvehYz+etRcXCOM2MLs0ZcSlReXc2C5sfUvjNGQZjwkSDanecCEF/tZ8r
GlLKQ80jMTwh+PdQwphfoDdhbhtGYR2g+Q6nnlrEsJ55iiuNFlJivQVOQA5Jk1aSeLOWpOg1w0N0
TbJsf+6cfI9dwnGxpZJqFdhSZQ/Je7RXPZaoPdZotPgKTehm3RqNMQg5YWVHUoY0yJX/77PN2LDo
VoxuU/5ircL0MK+ZhuiW2Q0vBwcWDsZaQqFEyHBsP349zp/HO9awepagvYqM0AVzqEE3OFIQcdC+
8Mm6YPEvMfooOlWpbmWfLXJqPkVYk3Xa2lnaRmRXAtK6kjNUD0tl07jN1SizIeFjWN3Lu3FflrEM
YPJnFHOokCmi/qxx1kftP1zXAazR2Vl6jpWKUJQW1Hkn1S9GXAE4r6o5a76rw0a8cT8kpzKUOr3e
GL06QekbO81vNxfYWQwivFJGiXpldJh1/j8i6iZyZCzkVGFLU9hR1wUw3Rp5uPx1xJysqTM2R/mX
8LnhMzIxo9tY08R21KRiv5mjry/rqw7uRroOGqJn7O97DV+gH6PN//1rSHe+PtICFGDRK6ORQCJe
0k7mvDezS7mJt6ql44PfI2pThMcJDDrG4XblYX7s5IjQ/HsNUOGEl/WtHo6hVzZ49rvP/cHg2YM6
y/3p15T5vpzfONjSElTMS7Ij6zJjXikeV6r2f7Du4mbGPWuAQaTUZSv+tugq8bfu+ABJZ9YsnUzi
fIZAKWzXPTwdbJlUT6MYBYFC4IbUzpYgRcBuAmhXKBwb64PF+L1B4ng708Fdfe+UmVPvWA1GQ1ES
UPjmnChHETY6Pqe+ArzEBMklPrb87/iwOc2JgWExynVxGV/cIrI8sqE5SpMHVCKQIOvSi0aNsAPQ
ktUIAgDa748vML/Rn1Mjsu28Gxmd5EBQTRhGmAirB3csRpPlfIyliGq+X8sYKs3UCHmcVynsrHaZ
9apDLllVMe9YeMMLLdPS5fC7tjzdCEywy2DFaKLuVaATkuzg7sA7dJhliEFcB3UWD4E4bsFI/Ypk
oNtmpMT6/yRe6K0F01TWTIIHuH8ZctVC6vqJGC2vQS94ORcu7Hy9Gc7P6fnVT++FAdjNcMxVWo+T
leIW3xS0s/Qxt8IPCWO/ZmEHEWFB0ckK2r1GiwJ8AjD1cnOi6coFbTpt5E1Bk8DgkbzpGY0DDorQ
MYPgvph8lZ5j9L0tkH7OL1cNEo+1rMUpWyKsmwa3GV7tu3qkkn9js09ByqJJ7JMl9iswyyrkNyZJ
xNglQPG1oSM2f37c79J834XE+BgMf8YL6lEGFGYvp2pjJgey2ZhPaasMda0mhwuA31w4h2vHbLjZ
ds7DkSjskwezHlKdtXwoUK4PSDm3ZCg0jSaUGZwGvDvPBWYHH/U0KJrARDV34yFiTG+mK5FT1PKT
09AKR0udzxVDR3yvNwQFLk31RWJOU6onIcCx6O+NwOogB/HGDCG0EAnBiWfhwC2NmM7r/JDlbF+O
s4IH0voUTTgWk6FbxLeo9lertcvfrD5W4OboyIXzb7VN39lSQe52nz41mCCzV9AiYNvJfwQT8SN8
LwQQA0jhxm0uSmQNHnlZnSugejizg4bQFD1pqQDpdoqs+LUgrW/qjbScrgXP2RbCSpZVYHmFFI8E
tLzJ2xUaRLbzV8lLcmUnV0PsyFRMV0IE06dEskAFtPUtsILwoq3P4sIhieM9XRXpsjq57PDyDXUE
/js1g2VjWaPOUQukeeN3/31BK/gtZcraaofXmKZr9N3c4BHSBqhjcKyR1rr8H5Gr9iU86A4YTGKj
zk0UzjzRU0qqytXHYv7rNSuX9Xpb3Czr3LEA+r1vn6eX7ekOkJAisx5zsxY5BMRAoziP+PeWQW09
izdVx9RFX4yqbkBOQ/1mAGFIvZFpq4r2J+wMkFf831NxPkhs+Qf+Tx+LVL4MixDT4CMySUm0/s6G
p68xsOwJrsG1PDvUdPplVsx6QhmW/NLz4qMMR3wSCp5wM0+lzG6Qq9FXHETzqhpLeekR4/zEeZg1
iuK8NQwEw8DFqniQLy3aUWYCxx/9PSfJy3gyN6CJ5dYQ5jF1Ym2w/analAtUQSADZLQKsxdGomhp
PePYkshso6TjapLrxoS9n7P+lZME0jLggvxppS4lTup1s/ouiZ6gXbYXEmlnQj9Sc0Wu2Wo4JRzy
PNDEu6xw59ApV3gLHuAJbRQ5fTYpd99t/1j8B8gqVGeTTEIGHqYygBcr7yZjZoOPTfeqbY/dMf3k
N/wvaFLblyv4DWz5dQNiA6uNchPFH4Wo9zwbV4f6XWaRtofN1jVES2D023A/aKACvHBn7lYYqk6u
i5jutRZpMCS8+L72L2KXy0bdxtClodq3uF4Ax5rx2qzjnIp/3qciMD3tr3J9W0EAd/MWUe+CSMcK
/wmVcU5+h02XxWbFCRR9t/MHNgZBc539uKy13A6UCcYVaM9xGYOEvhQP/ZJW3HrJ1iAhgahkPYyR
tyfKyKs9p/pmBDkng93tLTlCaJAsBBRohqWd4XduzYtsZJXiLxa/1ucAISRHiHVV3uoPoffWqAZ8
+sh2qtloD7a3TFQ70sux6Hfn1i29HF3VIDdc8pjcT8/RtqyiYsM0S6XpBaAOHZ1hUhMKrtAqnqrL
ZZgMndP2wzoRoZViUUi1by6xdRmm9tvBb0zYuSdnuWhZqgI444RqWOidR0sVNqmcK/wC9yb6xvVX
uSGAvpxMJZfpOLMmyEjwhjYGViyuLXqWICDza/O6BSEYgDzP3/PHCYPiIILYzBD3gzO3s2VGpD2H
rss2IWxTaF2nS2gRuGWnDVj2C+sw84Nl562HQtOhAMeeZshbuaBhYIdbdaWuIIARS3/vshtoYgCD
AZmhKv0GWF9i3kWkY76tSLkpss9poTmV1quN2Pp2u2fsNVYoiUGAX2Ciitafpf6zCOOAVmMPn1ZD
nR6QITQGlB8CB+t3klzMKP4/Ydd9E0RP5MgwX/sxftmn5MxgX1A6NjlE3tnVMj87QvbMJyd24L2e
1sPmdB967zgYFKTF7ypLt5wwKiNSeyobuS+frLCRpWO+aIMf1nyhntZazjK0Qw36cUzlorBcmW/E
NPCjC+DGXIe/bu2gT1w6JroyWfcV+oz7fS2XNRBGH/mO0q4a7oT892hAwX3/uthKx9oecR/s8b0m
4hxwaUT696zvPoyLOCiVz+IB4X2zLQmqYCsX3PgB5t/HspSR8i/8zb/rG/Swyvu9oZKc3rl6Jdeu
RJ8KBwd2VpxTAm45M7F/1BirPAUn71WHpatS72vLzn4q9WOZXKmw3h45/s81uzxZUXKwiz8ZjnUr
XsOiTwedNRaSl7agV5h2eQBnSfC88bATEaeZZCqxse5Ut7no7vvPcelagq3QHcSAIzOtzPCAcNXl
kF3Wv212hcIDNbSPn/acTZLX/HL5QkKaftetwRMWkEDMKn2etBd36TpZEVhHaY9QO2lJMqTFsVtb
RirJYE5yfFi9VtlBnlLbk6VGukH55nJ6QUqeoFJ8eZSJa6LvemQ7vQ1KNaOGFofjT8XNVtJf8ZvI
+8Jd76JrC/5zO74HPdADerokIFT4EcMQC42G9/CXK/O4775ArhjSNVVy5NxivCBOC1FLnaaNDmHh
E8eLTAB+S+v35d9Xpri1kOvagVey+rNvJ+AgOEc3wRI2AiwrZClkWRKzzI7p6EKz+sDzXuqUF5Fm
TvthNAgRpnIK/s4Gd2AOTIqzGsuSFVsMViZdEOa7l7bGhAnrziztHEgjpd7raZGJQvQNf7+ALpje
Y9TO+1oCfhWcwE8+g24n6t+LO/Eff5dJYxzDRkvuQ3RElJqpJxL04gIKi61um1lK60vdF4CsVsQF
lALyi9spfC+8PPpU4TV54pl9oeVprmBqfU+pdAZWP9O6ElqOl7ZSMAkVB1aJr4AdJTnFGMS2CGyx
+Fnh+A770nizOTTZuLg6SnIsGXIxSyKBdyrnFp5ccSQprajMYAhDmXvKj2WItKGKSuYceywS1tyk
J01Vs93+GvzekaN3mqTYMqdmaKcxs4aDiU9cwcq58hE0sb9EjjIqblak/k9AsfONIfD8STBWlLOp
axeC68CIyeAxE445ygsvu2gKCUh0wgliZx6vzP0zgUpCsI/Y+xNs96Zv9t5/cPr2RuKglQ2ZsvsN
v+dF6rbBeNNdyM/X1G7PHmaRebu1u5HdhKCq+xVHizf6NoXurSMfttH3gKZU17VYgUThnbzlUSlO
Yo2IjajbIcB3bkESfEPoL4a9FmX9KepX4mKNdiU+XZW8rq648UgVXtx8mbL+6Nnwi+Rpc4S4Mtiw
vfyHsjvyfvDck4LgwvGaqOeX2Yfr51ZGgac2m4Xlekd3fQZ9qB3vePdsl7Rp1HCTOnm6FSQWEIv+
q3aODqs6CE/3n4nW45Rzh3/gcImmaNmiSykYRkRIm1Apg6QNMg6YQ/iSenzjLkef4Uem3HOmvGet
yzvXQLeuTyTZRP5GNb21CCurchDgWLtxoJnOyZda4QgXo60RCVpNwcSYBtAbHgXltB8A+ZGpmxm8
Bo4jH1ImOSHl1ksaHTeCFHP0YH5KNSf5G284Z+sGTP1Q4alYccO8ENdc02c4RhhdaqqW/nDLzj0P
sBWiiPuBlZwfAVYMdEr1OqqULJiA5KqW4aG4C9xdVFvRrjMHqtb41uWy8i2sugjF7kck2v8+q1+F
N9Svm+JLK/TMeB1cKVFIvq8ZsGBrrmouuhxNil0LQVfmUJpHKPkoaqVvtb+m9os7i2S8mc5vB4D5
orWeUekiPDFJhOblOi/QR+x0eYu6ZNv2xODitCPlIQ+1RyLEFTuUAokOEOG8DsgSddY2w2k/AFdd
6ehWQWI2TUUM+pX0yqCNZsmesIMy3xRIFLot32JnoQoBPnGJcxGCKdxl9jhIROIaEY/gwn15qXFN
EdRgq4fwksFJYRUhh+N+s8UooaVoR/4R14TGQBLGkmE+a2fqU3oC89WTLaA/Ebcaw5ToXQOFFe7d
CxZNo9QDeVkxF6YJJlk+SwdukWA1vAE9s9cTiTq35cDNc7CR03iHSFEMK1k7JY0uPKvgnpx0u4ZK
Hrhkmc16R7sRIhHnO4VMnWHCOXsXmyCNugtNhqPE3gSlBlsq0e28OJQVezxPsEsOIH8dY+222Kzr
W05xoB0eeY8/avrg24FnhdjZk9DN0BVzoIPVX08VK+Had6FePMypsTIsjrMSrko7Z9bqQKNloVdQ
MAZWO8faMXiZCvY3BbOzAlUQ1fwDcONqWB/HWByKodcLVeuEy2j2L/W596fnyO5AqdaJDY2sOsQ4
TdZx0sUFHe8nWnOW5N57JtpaLEyx1U4zXX2x/2xkKA3/cxhOW6nyJKcm+VnXb4sOMpReDsG2B3qa
2mgwvroCDWaR7I4Pa+w6F8cT9l1zuOFPA1UCc6AMP9UPiKtgt171vA66PqYb+6fLq9FH8xrVpfym
l8zKtUUTkEC8pCatrWOHM8lx9PuGnfBWpXsneJ+/4axXMOylZeAUa5ilPGOJho++tkHo+FlFG5Xq
4ZxqxAu9zWC61N4rmUKWSXNL3Xf1krOeGoyITlMH0S6t2AAkx/26IyKo1Fcil07c2cDyjwCkuIkP
V6Etxu+YuCQUF1EuBIvaU1AELKumtzE9uFcuw7BW+47A8m5mSO8JCDt2/ZFfiJ+OcjwvK9IdfF/m
BbCmKT4PJWyNmYVTkaGw2Dpvg1bOs3cirzvjWu4OAIgiqVV6PzOYNdZMJYeFpFFy6TUtpH89tHeB
4wiFO34+LfHPyrDP9cuWLJ5JBm0TcjnGmTwJyv1QKxGzcaMivui2JlzWslvnP7+guksgJ90XD+iy
maUpWX7ntgiZ4xgz+jdkilNgcn/VtZ+C+myWcx8EO3j/5ua95F6Ohq00LGjkLEWcr5thvuLCc5pf
B8ulN9xHx5izbSnsKiPV9Lr3IXqcvb9y4rg5Z/bj9d8wf4PXShFp1pIf5Gv1dU5fHRYcI7tC5Eq6
Z0/Deyg6vGWW7oMEEzG2qPxq5PN4zYWuxKKVtAH6b55KjmmS3q7Mr7IvACLbvhwU0ipAH9ToR9IJ
eQCTIRz61IIjO5qH/jMjhwEyhPTJha9wiSGTEmFlPfkd8284aEOV8vdjf69DoutXGD5qWIgx9HUx
qg4hDqIAtcq633IycYhGP2iTDTjoXMG/P2w8NdR30MIFh3G/88Du9MIHzdGlRgDERapNwCwYqX7X
pPqAf5qMa5TzEgcMCG5zzuae08b049lXqi3CAUZh2XCuMlPN/Q+9SAc4aXjuK5zXDsMbhbuHm0uk
Hir6ywXPjPjVo2RIl5K9LQe0XA4DKori/h6qIj6TJ/7ZdYafDcFqxQWBZWcncz6sRPvGoxiP4Nyc
2d6c9Gx/QFOSZ/KPYzoQxAck7x5aA7L+apWONGxwQJtp6tHV2xcAmhNV/2UAPiT9Z2OlCtFRI+ie
BH2xvGqCRV6lSw/5LCjEUfv4nS5J+CYgD+vr6cGcW1VzGG3r72S9pd0lkbWwHamqR5i1yMawCJIe
x4L8FdvEKiG4/ODvteoGW7uSI+olSH8jZkRiazisefFzAeuBZxOc75P8t1sXd3G0HQGfzO0BWJDE
an5eqm1TlbCG8F6uqNj1FjthdedgdR1W+bW7yUcgj2sRy59WhuO/1LQ1WEgInCdsDuqC2d2WRBWc
Oyc7aVvtSB3CUEl8gqFqy2OwO9n+Kp97/n2NfaNDsuP+T9cDS7gdBLT7U0UJa2SSxPtN2KtmnkwQ
cNZ68HUYFQYPTzxPBNBDhA6NPzgSb2aYOixMRpTadgIsQ5k6KsUHca3jITbmJbFr+635oQP6Ttns
x1L3sfl5G4jjRGeC1WC9URPdcs83SCpm3DvtZzxvwu4F4IWRxRc1l4ktLab1ehxnEhJ+G4LO75yF
p2s52v7Ibb4YrTcpDYEcOsceoBI6YAuol4VMtnW1LsjfXw7uTDuIfViGQNCrlYD5Aj7liLD1YlhJ
rgJyGMAODA448pOEKVegG2o0wYdT510HvfkE25HXf65uzO4GC0fJCYF7K3m84zhW/11RPeRyF+go
tO4J0Jg7pJVfWDnTsQff5SqbH0Mq/spjWfeNY7d9GupSMRILdt0UUG8HbBlfD5utP/GCSYtbWeFE
4wJTcle8rsm1lFhwTlHmh5LTEpH4AvRGX7vWGuKA65d5reOWp4tyTahJXDZSx4mpHc8lFk7L2O0b
LF0jBUUq+WQnG7HS8V9+wkJLXeBe9WVJCbMGiuLeF9UkAh7Qm3irIKbfAi/loafRS1l0fBDVN5Py
JPl/zDb9fJM5x9F7srOhUKyy60ooFpY2pOKyjf0WvUmtKqwpZj8Cjwl3euHXZLBvtwoUAs0CKhPC
9tKwgIisVfGvjG/F4si1NmBhyKr5Mq+EfDV+yfgdqxHdQ3OzY/JyVmhwP1FFnYk7OfgYMK9BPLPh
FeMMbMuaHOeqCwX9v4zEArAsPUhM+TlKMtZxpK/wc7nwoBhcrw371lS0aN2B2phOMHaXBXhXpXxi
AdPv06LR//rghV50mX93JHUN0jKa2yo4H1qgqj5ym8tmxutucqVRdArMypJP/cCg5VKZFjWu8P2u
m+dqGeyg75pOZPvwJijq89RMZm3ESJ22cRrxoDgHFSEqEr6C5DI9uyYvzRsvkgFI3q/Yq+50bvCM
U17YxdgPY0bFlqJmGINEfn2mj4fMBgvqFsuRLuZhbUGzZUb9SQGb65ICNIRYsXiw2/RfS3i2+7Te
LjZDT57qEn1lUyTWk0oM4C4hlhEcJjIlWwCr80ZJepHLqd1dsRkTMjwKRvGz4JbLtAl17oRBOiIT
03FObsexMLHL++PukUaBZzUDljuKXufDfRW9oKVnDOlkQauL7UZyp2j/2yD3NTBf+nLmSLYyKANp
cMCsLEK2mjnzIzxj06T6fDjX4bjBNkTK5yZP5CCw8L3dsAVH7NjXx/0DAdSWlmSH09s4C6uAwAYD
f2UekuH1cvv3jDjgsp6TL/22uMdf2iA6RFChObulOxbn/4emq0nIZ0ZVkMzWz04CNEEjKq1hy6XJ
fENHi+teXLORZDW2jETKB0RYoYkzWBbZnoVomsFAMvBLn8g5lndbTKRyruSQUknI6Nj9TuQPW21N
J204mxlLkyEd5pN87PJdo1O77Lxo/dccRko0kNiKQ1iiqwOZdz22tl2MxAeV2brrmmuDZ0oc2F/L
usHgj3+jeZncSKRCZ19x0F5wmP9i87/NFao7XRrUfmTIPX0IaX+0VoICgofa+xfetlrrz5Ma1PCH
zBUNyjkngUA9Btb8+983GoPqoaWZwPuy1oqYtDvLWGhDi+ThSc3aSoWS2n0I8xTte9v2vV6J7obk
sQoQRg/6wF0qyR+JL33PFFX67SmL/QWN8EzSGEN/vJxPH+7TpQFUIn/iAGMn89nlNysZJ3ms2ZNY
1cWQhvrpdPIbveB8+MY4dp+avXNODYIHSmy5Ca2bIQTyPy2Frj1t6Me7ovFkGQFesAalkC42prwQ
RwJvnlddpnWfEoaW7GdSb0hX+CUThWQ+ZtFitVgwFLqPonJIJpleD+t92nzigb0cXDsOlAjpX3hh
YqtrGMhMEl5JCu1a3UKLS2qYUr9r+PXcMLa8ATL4XmeZQZ/d2IGcPge6F9Xfk/ogOHfpIcPtKr/s
oIDQs9yE5lcT3bFIscrBfjejij+xJ97q29OyexVi3vO5VDBRatrywspx9F+fJEGaNre1co53OA5f
CtnaNgKTlsO9Q9MlQ6ypt9cvLNimu6WhUAq5xN3Z4epO/2QfEDXsDj3mL7MNlPDzPy+NHSEB6P3O
J/vbKPn8xLEmYvnmyJyRAB8JCSFIqlvSAi8bae0R4VTV+APmxg3f2oQ3suSzu/IDsh3isvzDxxqn
F/Wc28T+UgP1sX537IJFQfEIAUvZu8rsc5rJpCA7/76nUn/HGeUbw3HgHM7HkHvsqDXfU1XjvP22
Sg7vlVuyInJ9rPOk9ENDBuBGohUJe3heIbrpOQgu0CwHSdybi/fwml3iSCYPzq8xW7GimxESReca
KaWEQBZjdLhU8DD2urr+wo4a0mfWN4zmxrDWsO10BixfmhmesTvLj0EISoCbXUhCVRDrvAAFw8yY
aggthbeQxYudAZxqAr9vlcWoKrDRbW0QkGb/CqYYrJgIjiFMRbxXKfhS157kIdCqjXmkBVsHXjbY
YfZZtaYphxXHCu4FK3/bqp974H1L4S7MF9LNOORxNgO4szZrFpGfbIPt3Xt9OplMK4QRrRgxYAwz
O2bXg9siT/Ja10T68lleOKHxyxE3VPyU+4Oup/nafXq8yt3v9ZQugrd7a9jdLnREdTScpXWpq1G3
tJ8lkfK9CI8E74VHrbs+lNTSxLHXNTvCV0yt6ufG3H9mSkNnd7CISFxAoTeXPxIntckUHXbt29yH
g9UCiDDtUQT63R7XZ0xqjys2WF7s6gLK6ojakXwOlLODcO43Erml6ljxzBgxeu6dYsIy2DrU9Acr
I1jehA8w/+84mqg/RlAOEEXfb1ttW/516UjONwkFg22668eSvOV/KQ7JIhZHSD8ST015NrCsp3Rm
FhBjX9arcMCR+o8gyaNF9SWfbcLue/mTrQKP8vadXkR1lybZ+4HLVK1l0UTsmgWBu6zBEX9dS/kY
lffXGMO9SR+p7jQ2Ov+0p4vbVQGuT+g0QnkS+LQFhDbUmUWGWlZeoe+e96WgnCNGglv6kHwb9kEP
Tmq07igcZi71O2NcyZ+boTzoEaKNO1xnK9KdInoX8J0DcpY2coJzd8sARtKvS2nYWbUH4acLl3c3
PMAl+Rd383QA9PE5mWuVRqnYJzxzPEeZKqQ3dUTzpdnpVtNCgWvqNsN3AgFJeKai50W8Pg1qxwDK
vUV0h/NeGXjwxR5RGdWjxCDtJBnYu5nim6V9g/w7jgf30+1pIeIyq9hvkDgakWk+y04VY/hCn1F2
+a3ZnNMAN9dKGcDEeyZ84EoF2d6nFKO/2KmeogVmOtTc1MUk2xjb0Z4pmZWhlj1qiDVh+cyVUXTZ
O8vjtTOcf/MN00HCOf8mYuadHtxH8nuGotI3bODk6QgoHVwu80hY/GfoRnnivDwF6bM/rfoOjUeL
pY6AO8MQO5SaSJs1Bkq9JFzbBCXjom1CZHC3Ajo/03FFALcLZjxYb7+4Q9ZMAHqM0aEgsAx68NLp
nPgKyJ/hAywT5L+/Zlpq5zUw9ANtp+aUvxenrXjbtNpXeLFjcKPC9dnY4D/8OPkbM0E2+SKyF78l
b6JfGiPGd6bipdasBMHkYNT5HWEKQkhUCq6WabSvI7YDwjC4bx3BHE49npqyoPqkBNfE2OXk9Qvx
N2rIByOMPdZm7wgr5Z6QLiplbE65XzJxxJi6/W3jGar5AzO6BC/JTZpq/YrPKLGxb6O5PnKpQmsi
EPN28CgarNhflczJnD+f2TyQgLB3piqMPxv51siUdoFqpyiedGxJXofCFvS1f6t97tAepplPldc5
wTAyPWLeSKv6tvyQ4eBcDY6fHnc2H7+DDaPrJdiTzIb7mwFzdvjgpworzjK9/k72Z1nOWQNOG/BN
+17CA5CZsrLku473Bk2Ndifx8SVCC3slCLp7VFS295p94MqnBit0xQfSHWU/IJlVIgGn7nz+DoyY
dlcdEn1awdUzIPRreozW3YhWuGZtVKaTGjYVMuXbyVOk+nTWkH2kXtyAgyJnthg9Wf5/FoNulACs
QWzbwL16SbdBjkqDcb8OVOso+S9478yN12c2y90BpqQ38T3UYyr4jU8dIeRXki9yaIxfbxycUzP1
9M3KlFdP1wOTb6tjilNqByIFgEL2lyOPyr5pCjjo1iE0dk/MLxWE2fvcrWECW1jGX9M4AyjKJO3e
5GG7VQ9aDvk1iZQMHnBnrX9QaLLOw9s/FCn3/Yjypa4u94bmscDdBv5rr47lzmAHba7ls+D/B5po
bs5TT/vgx2XsBII8kUR9dB389IlorXHp3oaLOaQ80u1qltvvrOPsT6MPGtqnSju3mdnJhRwD1EzS
p59vJsqmnqp6jXksWi3EyUewyu3P29YG1ws0yobMqkoFEkdh6aeuD4re0/DR8uRKeG4P+sQUzxbv
rLAnfE4gZk+vdu3ovjYZjT8gTU2CO0YwTrMc0hXd01ZG1inhahLS1ShBuUvnjt3UG6w8DITUpS5d
I8z42Q14+hSsCGvCYXNtGeg47J4zupEW8o+2yOvEk2IQ5H8KkdYge3vng7uEFPvXGQP4srGXSYkS
YNiUUaaUr8WPg36X9TJcZ3HqE5KPDpSj+qo6OUiWFNcIuuxqY+8rp/mgrzh7pKkp8r/84Jq4HNkT
HuCteDQ7r5kPtOKToXfd5pEN0FwpHIasPB4xCvhteTxbPJWyeHwTTxy7e3kpbKAzwJ2xllrUMdhG
x937/tyoTTA6uzOnlLvhqhp/UVrX30nQUHcdh8tKE68xOrvhAuqLTzywvgDU5Hi7il0AS1AasWYy
I4sqOBn93xOh0xqdt/t15f2zcFi/RGU7iG4QyL6MxaKU6uOlH4IZxSahS+1G5DIpSOTip06ZWlu4
eiGeRxQ2uT/MeaJN4ggif303TEqpMMCtAFyJMEEdgpaq8IW1e1Ro3irgq53YqtqYPdfApucxTY+c
jvlOYQK4c2ufeZsftyn/pHCM39klplWlxeFk4DBGNeEUrSXl8GMbggEGVy5xldy0f5Rk/9L7Y5NI
IUv1u3F6vimWitcDRrWLXw2gSxEDELJn5075sN3GKc2GlajAXp1cbcyFD9dAcanJFWxIhSi0YVRw
1XGYgxBnS2tqLHhWIzbZvUfz1QRrlTORgbDO4z4/vE3tCHqPqzUI41b41qqfxEZFkaK7ISq1QFG+
b45W+3Q82uRCgqxg/7Mdao9hob2Z+KyjMOJzyY5etNExDH4c39XoizUHHKLGcKOqXcP1/cKqEZgK
c+n4/pth4MLJLGsxLBl9DRjIj4wqlK136pMoCC2IyMGvEyCmq/AM0IwRFEReBlMN3eG8aTBCLN3S
fQ0F8Yd9tMK7OsWXC/sO/QL/o62bCPnNyiPXRd5TtcCwY5J6AYC0GItRYQYjU1GG42LfZhlYAFao
67viyPXsQ0BsGfJIvqZhJq0mAb54Zjws2434zJ6MdKtBqwZtXBzEy2IA2Gp5Yj9Zb6Vv01pdNciE
hZJ2vYzdeZ6mLCt55K7L3OSyPzJQ3ZQ5m1XdJHTFh3KM0ZTUvRdRbtcDK7N+5l4Aee/OM0GazJBa
DKA3npctlod3E74UHGMce07knMTf4lNfCOyzCDdN4vKztOHtuiVzcZn+M5C+Gx/21jMMzjXOu5kz
E2w2I8JLVb8nUNOGoKf3YS35GfIP7xInch6XGogEIIoAL0afLSE97zmQbT6TNS8SuhbOAU41VVH0
uZZRzZ1/7fcHYIeTi6rEmafMIRKfcBvDJrGzJCMGJTL2lXgGz3FYivVenLmaRSvoefwihlVF2ZzZ
mZZ+Bcjx5bEawcyDIhdk2NCCDPz5ghocha8tZ8bm/iaRPVYvmhc4O2OqDEsIAgLh0CC0ZeDeEdzx
Qs2pd+ymy5zv+MLPS3IJd1GV6dJYEJqEGnNrlFhDP1rfpNEpATUnlS0uE08nfEuNcb/7oqr23gTL
BI8lGx6HexBRCqd6B1CYCFW9chOWFgov7Yv0C51gotp2Y0Oa2pAzQDcNRhEtJmbwX8de4cU+qZ3w
iIwA2TO8J3/umCW51bq6u6aNjFN9oT1qXI8KESDgu2F4TnZHZmHkRyaVMa1a3d+Qjj+gy2ZP6f8D
u5UuBl30L1rdjyf2W9Q8mRpqt1AeP7hQKR/nWLh53HrEH+hz2JOrE1KZ0G2JoXA6xmTExfhGP4aN
a4MMHlpy0Fmevo9lOGXcMNxF+vjIZyIeoOqOrKAbRcJTLK6bNMGIAz6HFREXo/IEIJxQDgVkDgYJ
9AZEz6+9SMpnSRt0Um1aKCk5uFhgCDkVv5ne07Ds88xHNaaTcAZG0yM9BiMjTTckClWb61UBzR+J
HdEQ4+C9+TRdObtr1cTP/zpWzbqvggjJ8eUjh5phr6ZArbhr25jnhjIiz8Z3LYkVrye3qZe8O2yo
dbVSAK2wNEMky72uMxz2+7GhGanRa9AUTewf1gRyC+n+hWhsm/SOxHKDP/Ja+9gJvveMDnS5jOLM
2wkLsB0IetNBUHjXjc4qH5xRAAKKglNsP3kEJS1fUCFTMas1wze+7qsVU1rSZMKsAmFpYrt6IcXg
nMxzEGct2204RxfkAtV00c33nJ/RzQ5Ipo6JzepnsqfH6h81BZpGrNuwFfEmrzrEGmLnzzdSROfo
45uKnzOS4ZKcoZxRz8oMsY+/n6s9AFnmQT9RzQIIVqw/QzUQPicqysKamzqyqKWXusX6fcfc/++v
cPpPose97gZiu6u86lVrWI5MtWmrHbZZt0bCNbLvc0HEHTxIWzOZEN6wHGhWA7bJqVsz3a+Bzdv3
Zy9qjEs3JPYPrKZ6oqgQ+qwgnGlFanKzOGMgRJjdp2pMqsLYFPOI9jiPKSUAHFyMZSGSO6g1HTxU
hzxVuNiWZ1dZBzJbiWqD1XeLi7n5wjfpSwRuSZBunZ/Q28cI7xaDfkBn2+1+EFXgVlFCGV3wcYxf
JWQMPUzuFODHUI3AUsLsRH9rY6FwtkcijnPjxyrR0A3C12Ux1ETRO9Ic3CGy0PcNfkWwPkq4yona
+t+A8HqbkTe9CcwY+hkmnSPs5rb8HZ43axypIeY8IgcDOdeDr8rF+MyMrKaXIKXs+Ki/KVcv30n5
5qtQwyTHqL0hMEtGSreFxDrLz4szNv6I2OEbzPqrs8U0dCsuYzR/RitdouJZKVXASSQcUvpAuz5q
VQAjywEPtdTpGkVcYnRc7RKduTgonY8fhA3IS6JEBO1bwiWgMuuY92Ps6GvGWcVSJ9teYCqFzkfj
4vBxLWoHuG18gSx69rhrmplurpXoM/YiR5tycv4XRZeacNJaxBX3RhEaAdBCtfy9GCPzxlUhe0OY
8Wqw2y0FXgjB1WaSbHPFQMKrWLr/WIDgku6cijwnb9z9s/OnTkNdOipEdws69NCOJbpvAHc6bD9L
S9V7FTKg9HpO1xoZTgpIDmKo/aG2hWwkPaRdcIwpD5YHOaYLjJLSnyFlyYvo6lgi7Kw4Zmf9J27K
dz44lAPFxivXzqnRFiCLe+8RQOW/uuL1X8q6nezKic1vDFCuOzWKmDVaCI++2Ap8OBwXWvRBKcqG
0c2L/tYgjYhORPYOscuFaCnUJhRygPG9DT3R3q08AJAYUd4MaSBo3JseOgIHnziE4d7uLj8W50O1
rBm1Y3j3mEaNciLBP8JgaAsvwsi1Xz5ZSpg4ZdImIUrfBRGZCwfJ4S3UhN5rH4BU+KAPCRuTuIJ1
xwtih7LK5vykFnl3kDFzAI0PZ8OfnZEteEwYVv70LYj79lV9DOk5Dkgeca5QgapHV/BBwAJ38dWt
I5n38AXgpiuT+sQQzB5/Me8MUBzNyYpx4pbYR6bSmQ8TXlOnhyo01Qqu0pHsxO2farn0GC8nqFk8
4FTEmYDtsdZFw3CrNSfjY1+l1r/Q0I4RwJE2Ue/yLoFOIImEMeeoIviTdHhi4MGgj6wq+RIfbL2n
C2xD2Pqn4JVqMFJIA0rSWuAmaWWKDlCkmEa56cJln7SAfnxO3+O/Olv4qVa/JEdCJDHtMrlOYKRm
OSOpWZp+ucEhHjWedTvZWBCUhdPqHb3QNio5FiTVTx9czN2MWHt/tBNVs422mIrSHX9yOvxX86K/
V+XBk7zyKILyM6vy204v8vUR3ogfTpkDoBxKrcvqiv0yPysm1Q8pcZP4nhkeviURKkvf8MCMxt2T
EPeMA4OXtYpS0LSR5YozqZQfajjJsHMgsVV2VSDuS0BRAKyTI5SXHVJ9BCMIg6USrmXhDs0FwAEV
kvMaRs7W513aycL2q7D4fevx/Ik4S8KqRH+PUs3holdSLMw2/ejZ9bYZ6sh+p0OUXie5uplEKUaF
fH+PoSY5k+Tk26YHPC3gy+fmlrj8/kq3hZ7IV/hDvi9Yr+aisTQpqf3H3AbI3TLxy1+woOSzD9Pb
ihra90b3Kt1VbkrdD4qRf+Ay602rqEdoJ+AFI/5xagtLfkr79L5Ptixssxnm18A8grRvFj/op5LF
MbKL+hxrFCEHWIZ4ZlSigpqtad6G1JwqUIvfvysc6gRoYJEHY2gLrTdgVxewdZ2pv/8pOlNjx/J7
jK0F3o2SYCO35NlMJf6nJov4IHHuDFBmvqulumdQm6rydmpLsDBl0TrJ2DD78FIIR3ju9SB++mrZ
fFr27lEj3F8tvSqvXSFZdrzpjBkg9y4kTLPLHOIzhcXRC1nXJiQ8bdrLvo7pLCyC4UIKPygrumSQ
MEdlGi6cQN7z+zqlLO5OKwUUmWAlGiX9/LSWJDil6hez3TNt6X9bEr3lsgXJDxXc2uBP9MnlfBE2
tzGoSQgdk3ArYijodKqJsMf0ktoB+dMjBORP2wWQ1JJeJOx7veOsdPU9FXVgnLR1k156RkCFDiSo
i0sjC95sTfr5xouUIObVcSoc/DafvCwjgphf9v83kyLp9UsdRmFYMkGs5KvMfVKUI6qzuBjS/7fO
hQcoM3Lu9MvvnhDMx0r1ozCFuXKDhHxCAG+Gnb7oex45cGV+UB97xO6jKVRqzmDOFEg2pdehduEP
5ua4KFkVu1z1bDzhLiJ3NGY6k9AKnGghkDVe3SGqPOfjZiOF8icsjfyYfCndJB5CuKhN7OjbIPeH
+p04MkbZ4L5exLkrFW6lJhSKRCdL5BI7gndCJz3STjGz9vimo2MoBsED39IjetrIGM5HyE+i/ZRZ
ig2QaTkMZu+ajkYtYZJn5b0J/wtu2vD6nJHrO2G9Wzx2+F10PM5MXSHD2IbrPvyVYhlTChhSabeM
EdvnRSC0A4XQXk9VVY7uLg/W33JJS/M7xcj2hJzmJ0mn8UgUptLiQkuywat8f0PpH+iElrs1/wqn
ITtjG6Zt0UZr6uaxJAu35SIsuqe/Txfn2H6cTRA5z4b1MeFb5IlAmCOtKbEePnj1GdniIIYaizUU
KlMS5WqHNHkVLdUZQEkYGiV2YYSE74b2eyajYJ7c4UjAtnd21JNvZpXbNwk1ZFMEB6UFsy385/oI
i0AT10FEktKEaC3LIk6cXgOUlCudJ/YGdIVhfPiMpLsLmVLHjoArV8XquCNtdd0WKssq09Q9kupv
ZNnZN0xq9ZCapq2k7CsdFwq/zCCl+s1HAzXCmpzmPGJjETjlOeeqVAFF9u3Qf9CoUYn3rF94mZh4
ojuOHrjBo9yXYlehKhNKyVLFCRXe2uHujMlB9q6i/x20jvY5vqOCeLVWF2UtuCHiGJLOUE4OVlnk
TOut9LaKoWujqHdEvRTjt3X+gBxLQmLlA1KvzYCCaqiBrWRHMqHtKiLh3eKo/jsIzdXX57MCn5oQ
qrkH4JMni7cqXX0eC3CLsbVqFoy0kkyZJvanx676qcrJqx3aw0U2TCn0HLmf8Oeg3/8WCRz+uRTv
Ou+tpx7b8Ss52q/OIh95g8a5v11U/81TUP/BPz/H6kMcW/q2ic0mIjReLvruWEhWYTEy+28BzTSF
r4E1yadNGh+avJnRcEiSlPJwax5QDBCwOFO5jEjNzP0e5vaSBvn4iJTPp2ZDmQkr0q73V2G3fDyH
D1Ki6EaKDiXu3quZ3mGkjSUJioaLpUJ0NLL5VWvnXFcvKugHGT0qx1B9yKDzXR5Or0w+5gzg5rw8
f6P0E/TrumonWWUvsX5E04XlLTtUGwO+mutAUhOKHmK393hW8Ed6MgjMnx0TQMrzENOewXQdVWbY
f5PQKjFGyCeFIhHEdUJawErVj8P7NAmSjy9gDY7h5kRkX4IT59iZOzaxPy9YKFMeOy+tYdUvb61T
zOJpwzdkKn3L/c5Z3dRTkn/F8WOfzb++s4MhiyupurDevYug+jNIi1ke43m4/nZRE+sjlFujUkkY
XblxpEvSDYUL7kKK5E0p8G05L0ol3dnvAeLIpHd+/FUKKezfPuNqR8Y0dMADkhG5uLOz2YrQ9+mX
mVrcVSnwlJB3rlwvo4fHpa07VRXmRpW2h47Ikz5Z9H3jGHmUUaDJDxxejJEp1EQk08oHa/+pZ9M8
1qQNrQAqJ8cmrp1k/QH0hKNkcDD5umTSrEIhk4TtgILN4BITIF0C34z0kNSoTSIf9rFpsl5JSwtm
yQ7/wB483bGnZpmEcwR2gMY6KwFmyZPEJ7+QNIEcEcJ9P924cHwjt4v5ncuHoLQqqb+9v/AF2Mbq
dAd5v29myTdivdD2Wadcxx7GfIeuHRoHIFmfrYeKdJHwK1PvswSCEd+RNoJU4fEq0UT8BJ3upPhJ
6iNLLCljbe+qW/wixvI68klhdrVJxpo8K0W5hZKWfIJyoCb3Hg4YxSiyh1hkqDpOJDAnxsFt3+NB
XJfeSrtwvY5KElq4YuxBZlAuQ30TxVWYCqngXinj/51OuyGAQ1nIekAeoNvgi1bKLYQeNWxyr+E/
sTsxYgPwkp1SNI1pAqudgDK83NJpJ/CPagNbBS1mN/BtdKYx4YaReMWpPbQA5d8jXJpHUR4nQmCN
xXmtLMP8VkVKZxmaGfo1rDcIanN5/tf4+wlX429rR3mmu+ZUdwcOzcAhiHjS7aNpsClZQm4P/LRc
hZXFzXP7YWhDbRwdffyF6DYwXTW/wY72u+WdvMGmuGxnYfIHj/rpi8xvvBVxj/EOqaJEX+8edkYe
6H802lm2q5anK3wfR9fhcGtpM0D1jeObiYiL0S7W+Ua14s0f0Zizl4bsQQymvf+jn54kt3dqr/vN
VaU9ZB9zPfK28H0x6iKTzFnNmQSeGuHaQe5wwSnWUAPmbVFiwTPuLgw7sZF3hhXYUpKwy6TDHBqX
oAhXD6KkmA41Of98dq45y8HFqG3wf7SvSIKjxN3LOkElgpdptwDkXEytR8NwghLLAGGmxNC1aI0p
ZKD0cDBJLfY9eRyRC9yppWjGvyDMbCrz/noHa8jux8KzALJE9gUwViOBrUDYuxjABlbNfSUti+MN
lh6MEHXvVmldBhRKUbp6V26cacpjSGjnYs5EfIK1IppzuA1ZuSj9jeFxZ61L5gzl81OrwMhGNuka
RrfBEL+o1jD6XvjS2fMBO6xMOeY7XWkvt6Uh95LH5gVFV2kF93+vdIP+ZWrAbWnjfk+b74wuUZid
HNtzx5bWOysLAwnjjyoNylvfQyWhETnjv/+scgTUefihYEKi00cccrpbburjGVzM0i8fZPfzO8YO
tqjHwU2mnELSlgmx3e+QdoAa3sfQLavOVNqP/wOcLE8wmVJpitPuoP138kKj5gtQ6Pzq+91vQazG
M23e7cdnnH5qBNy/I/kJY8DP8nuS9hKq+eSmud8nOXPX7UhRJcWIafSe6+et0IOXeKTNNdI2e3e2
z2WfGKxCfEBIAWPdxHtwYnM6F+YP47NjcGSafY0a3qimXH2MavEQxne3UHSl9kOtWiR7vw2GECy1
gJx8VY3D5VpBnphA5BrvDRJAjOxKswhatSkYZT6ToLCPpwd32V+kye4pdUuqo69sUn3DH8E1KwZU
jpNZS8m8ajiSl4VuYTQm9Zg6EqiliCsskj90UxWgGwHt/yNo31l6BUso9zPexMUeH03dZBiahzNV
hHR54A0ISzo4gw7Lmq8gw7rZs6ahHogifacGQjEGBS82LVjXZWC9nOFMFIlnmAO2msrytUzZP0ob
GFueYkH9b4sx9ra++fPog4TatlKjq15vuBKXfMROCBgShAyQfDQhZGaSerAfcpUZ/F7xqeK5LHLF
gl712TJxtyx1JVjtbmg35iLIfBLGZmxxo/zJnkPwK50NvLoUpmpsUNhI5lGysjjQ+9fVphmaj6a2
bptrmgiocFdOpHqTPxvsuBR4LWFYR8NPqbp4ZcT54q5/bJBUYXrwLoVKg/zb5d6JYBzcSCzDFx/S
Qf4MGePNekkvuTBlWYbyGh38hN8awvC2cFyIYuLbMDMQzcBcvjxTy9FWLusEu/KsFOQ1nMrqR16Y
/x5yZvENuhfspGG9ROWBGwdb1yA18iaPXGIwBt7TZ2jozeU0/B0KdLVk60B+nicXgZtxPKzYVKfT
YfXwQ912CqKHaTgtIIQhwkPAkeWsbO5uNl9uoH2KZwYfmdykyVf+SKA4GQd21YWTNmhvzWbsPE6j
WZ8kJEixX9kleMjp7MWYduko4x7/QsRIF7SCac6iGsMyWKjAl1gYYeRfNe1Y+YHbNgtIhlBtTP/H
ts93Qo+NRbEetHjVXeGobg6QISaffDBr4HCAAVZjTyjjkqWvXppYudUtfLfyUEuw+IwneD4FOUW3
UCtTlJjk0NyMbZDvACVXOYA7ItxlMH+8ORl2cF6vAjU8g6vZp2Fq46teb5NsuHMqfq/2a/tM2lSe
UEyFIejQZdrPPQs5X2rzZoAGSKPKVkE+O0moR2obZEPMlTpSVuiULw3zJwv8HF0Ypdl+XeHErmoA
QY+lhHps5YgdxzwFI9Kiwd+4zhe2vBArUOpw8FxFECXiD8uhFn0VP8R7F8WWK8QZkojp2M4hkzue
S9ZRQig3fkR1PeQqrQuTSoVPImm+GDZL9kxQCR2pMN5Gj3S1sdk3q9gTuEwcP9AYj3RJIUmC0b1Q
Sd/C3MbbiKbz0zXB7eWrAZyhKLk9cXLeYBp8ZEYZeWIASh9aEFg73QPV13GPsEqFCIeArYfagg6V
83Kz36bVK3F2vZh+gAXhTrHsDkoefu1PA7vRVdrIsOapvsyTXVXL+9BGQfz23I6kJ+VZYz5Q3FU+
Ix1BaauTApXev7oPPqgMtuhjN9vURGqnWjRVOng/bjR5n/UjRf9r4tWLNAH+xOMvMSytvkkxQwwd
erkT1IyQInX/jR0J79tLIOOMhPnT+UnR822oxUnqNtzz7oatqMO2mU5IKpPoXq8WBUgN09SWYejC
8IM5AQw6L+BzK7bqPEj+SQRna4AUtHHtp2cWdNmt6JRZwIzXHE2w7RnSaoX51wmBDpwWzkETtpLs
JROua/gNm/DP4FENr5A5E/l2VBPnFmQSJQh6cd6aTtjsK8r53YWYlLKS2pNWHw/+1OoNCa+A+23F
mgatZRwix0h6oeZf+VdnMtsov5rdNep4FHAz00fyjqazp+McuPSlUilOqjMfbgIHrKMqndSL4df4
Oc/mGdmDmvSHZT8C2sdb0ZOTwxXWzgvSNGM36vACl0j2o9mY0qSmhDSDOl6Y6IrEtuUOAqEioARM
2ldRmJhat4tkocsRNUs6Qz3SFR/JVBTZ2ZPAF8t2DrxMZIP3jMpv7cXq7erDHU1gPXn1NIHqj5DE
oqOAcnFKXB5v/G0I7cNKoVce81gzfJ818siucJPDLzD/L9VafLTZpPxTNw3vyyyvznzu6Nrt2/te
rqAd4IlUZtbwUNhBDofe8PwU642fr7OAMxaaGEyMTdbNdHkBGcIevRHAraxGJQXu2yeEb0KIVTVx
4iRyHB+TGTxAcPYkjho6JEXvF6/annPmxn6aTD5wLwkTcp9roskgb5Uj1Bn+HPz+4KzO3KAGR49b
s9QJBn7Py6n28KOLXGW8UypnohY2VLjeCaw7rK5SP+PvTc624oQffWCkvGj/mWx4UGTGxTzMQ1Ke
+T8OHfao05ZkSG7CEasF1ZT1NKs7tTdblct5mKW2nMG+ZTMAHP3Fe1WoBsxai1G5EVwOd8UTo1MZ
a5217LggjuPGWLaUmeY8+++EdUN9fpVieyvDk8sq/B6+wsCCD7B2iToY+UoRAoTYpVNxpOWxL5r3
nmi3tv5MQNeoEdSsi7haQ9jUh6dCjdRCefrrTCcRnb54vFYhSbfyon4GjbHj6d4ii3Ka5OkPoXzw
L0ea7sAbcu9LDqIAbXlNRITvUy8JPmW98e4hRhhVKZRrlJJ5TDHNuaoHwelxea3OqH0M5ypbs2c7
ZUB3fnQoTLI+vdB+A0oAb56r8y+z9ccc+sqQyT1GVjh3QCo3MxJX7ewDc++I+YBwGpeLu7faiqlq
4uvV6EEdgdMqL3iAGShT1bPCgMw++YR8ACThLGIyZ6BPCCGD7rNCWcjgzPp4QgDdJ8qTA0AAv6Si
zhyQr3tMXhXgzf9SJZB/mBCqPKEB2go5zZIzoxVTooxcLVHGZtppmfAnHU6D6vcv5rmlMMCUmBNf
2MqmtfX8wN9g07QW4kBi+ZUJmSLDAI0pDuPo2G1qfk6PlVFjj0cRj2EiTOrrUdzV92B1sN7/GOkz
/JXa3s87/Qf9/VINW2CaRZXWR9sNrHn9qQiP5d1t99AZC3CWH1sB4bc9Ik4A6547ecVz7Q0H3Yfl
uUmTlFqOpl9SfXON/AZDXnhbbGSARtFpdgouRD4c8PNAYX/iFcWaoyP5TmrwYXYHz0h7XGDBDDYU
yCD7cUZZ8Hfs344xWRbuMQcij972mlkgOan4fjiMO2gxkwkhu2pOHK4QZvEglhCSVgrySgYWwWit
12rewisH3/kD6vQ36Vwc4xVRtBJN6QEaA9QpEmI7uZ2gD29+z17NdyJruYNjMFKwi+b1Ss/J1LKF
PCygjiQZ+XHHmV1gg56udTqSYJO4T0N0lmhleSmrwE9xe2Agrj1VzsymNB7hlkptBNQpB2GnAkYk
YjiSSLhIEI4OWEgS7zj59yHQMakN65N/noes2kZVojolTK+PKun4BUq5LdqxPbaPrfCdwyZNsjku
yk6gi6uOGNe5MD1as67N78uackY3fpFQH26JjIpUEvC6BgnfF6n3b57jaQ9kskHsd11OxgKdAtBV
wC1xRtLtPQAid1nyhipT48F6lhButuNkxQHgMSwrcKjSAe381SYeieyNC9/p+b2YzsMx9rtBy8zx
yL66eh9TqK/2jeeAJpGVvHUdgX5KNpFss2UWY7QXfmr2CRecdSLKOK/onGNWcIwBoqtYD19RcfG7
Pxry6J5X2EUzYpz1mRYfUauwvfOooHbqrc4xUUMNygJmFFimRsPfAoE5mUUOIrBjFijqHr1+es7Y
m8bR0B9qgRFJcKvOzxQiFlaCWtM6Y4yVTV+HAeuAIsppBsc2hu3DJuClmr9WbKkMZ3JgGjfdwGqz
Czh7c6nDAkBHDHG6/srGGDN40H6Gq+ujKO+V5BFD53PkRu1AAVZAstjg/17/3GnJyHauM7PplAaT
HqeMhFMuQfoWOiIqFRR6GVVXVbKU9l85aOYT36o15wEXlNt8inVnARYPm2VmyDT04zjAJDdbhMh9
vbadjHJB7/U3dGz/bceONIyKXzZTpKjTFJedg9N9QWuLVV08of4KZEl4y1EMsLtWI++lVODJ8kuL
iLKcuha7TBWWN1f54PXQdobqm1te4tn90jqvWAx2i+Rvxne7wStZBX8DZZXv59c2l9WIX9qLCkBY
/ClElrJ9KqYCxjzxpBhBdQZylTQ1J2C+/pgfaOV8yWgMkA1ByXjvly7k3MWfKFFOKpLU9U3bhfSw
WVDgrXpdAat1CtB/wvu0SlGkZJQM0f/JUwtfqZLGmmVC4peULse64gs7PsRCEvtlMe8xjDjdC+h8
E7iWmvDKKj6zsXHV26EaCaRMQNHobd18jqaibAeZFX4ZXud9A3U1sef47nRM/U+CNLBL9xu09183
tDD+5UXpUaoqcR9x7C7mhBICEs2oKVtABlC1KBdAul3Vrued6ckVjiKZbihGCnTEYEtxdOZU23n7
C1bfh+1bQPMpoJsY5Ybbbn5oVCcdUJ2pyRo9LoahBFJhbZA+Aoaq95sZnGjFoPkHwds/F0sJath7
ezHa77Y8wcQKinOT9c4jKuD6COsRPETyeCWzoGKqlaEmS1+q79okwboChAnoc5fv+L2ID6enLmhT
BCVPqQ8URPNzYlD1982IxzwJuHw4d18yUYyAkiIG9XS15qB9ldYd+RrjmIk28e/g51c7mwGxf5OR
gB4K0rTmD9SKFnGuwzVbyb5n5EdsZQyFdOPbutcfMd2LJmtebN6u7k4Jv3/SxPzjq0CFp782Kody
HYBiLihOQSNDUUghZpB9GejcpnrTrLo4Sv67EtNDEeC272FIo3uhItpFPNaOd0TxEG1cKg3izUd0
0jswxzXHTqUjhdKQG28OBJMETYgnPK95WnK5QV1r3HUTJfT6CV4ST4y8qKGdR53PMbG4XE6i33ri
C9TN2Xfe8bIrdEA3lGdcwiJQKf+4xc3VI2A21rD/VdFpOEB1WPkNXp4SW5911RhzF4//USY6zfLN
QP9K6YdobMuxgh+KJXwHddyK5TfdRareEoDLOktBRW+cy1kk7KJ8ixiS8VilJWMW5tngih7llO7H
wTlNTFMsZXfJBRF+bOzejYjl4Wo8SEceHvUsBm7D5QcLQkvXUlE2tqXPucFOfIzHcapBu3+hUi2g
9K/PGN4q1mLXbmn1FOp3G+/aS2rPTuTUExbdFb7PbXYQE/GaCDtwowjS5TLKOyLbYrk74MpscLtr
01pn7lyK4n4ZjgAWNv1h7tjad6tH78lyH810/vsdG6NWYrXyyVnJ9QRIFWx1F0sQrfFI9jpZb4a2
mc0Z6UkseN3PwqZ7Dd1W1EkP1699Ujh6ylcYNIS2IDvI2waaCppZJ7xFjrqFqay9kiedmOyURJrP
CpALGviDpuAhqledb2Y1G8MRo3K774N7jmtxFfBk+uyO+CAYgGpL+zuussLBHGC37aCB6W68UD1b
1IWHfPU3KXtDXGTVjeEL673Z7BeGpye29XmMlR0jScN/ihM7I61Sm6MsjsJi3yqe0Qe9w6nEqfYh
7zbP2FAehllqPzE1T5PHZX0PhDfqPOaVwkYQf9eUw0RdQcA0X9Ick7cTSjRf2qirW/G7w8RNapAR
ZXeNdAcEsMAJ9TD+fBHlTCm6IOJ1LPP5KKBI/sanvdjbLLgY60NognlTzI+eX4F39nkKdG4EQ63e
pNROugwOi1d3e852UpRJATATpMdQnOVc/FBzgfLWDqt6jFKPevqhPu+toYCHjQ5/kIpYypIv60f5
FdimshVWQZdth5R8KqTHg5xdypz4ba2jIq2ixhosZvakYLc5AaXRpp3Xh8Y4b/rf0ch61THp+GnH
RoUHpjvpbRtRJx2LtoHjwPOvxY+JX/mrVdH8JxefgsOa+UzDS3o7rVDP+Fy+5+37Zq6AzRGaDwTX
Hen0mMy1eHFW7s/y+GP8gipe2t6rVskn9VDAYFjsDhbzoDRi73bEi0Z0zvWsPWQTZv+KBU55wwcm
NlkY9Ek/7tnLB/KCy1k1sPgInndGyhJPs3LYEa1jYfLiZHfJQQ+IZNCyrbh9zvGwfkd+gNDWOHDx
RIw2Kh8CtynFZzNRV2hNGS7vW3fCxQUst1Xn5vnh1d1Y9MXEaY0IU4Ybblack/OOxJmOPYG/nS/h
CrS6sjdBfVUrVBrb2aS/VKcNv9elfXhgJBh86jxW8Wl4t7z+tbdbEIdHjwCbL8zJ5/7eR65Gp4rN
pGdO4CRbFL8akV+HrUiYBaQs6Vs6Bg69OPpAq6/HqwnLGsrnHNI3bSR3RqiVS0u/ssS8PYokq69N
6TuEJNp379sPOgKJI4dEBT+kuSdjI6be3sXZnJgVZ99dPC7X051a4ltd9raKKKDj8TdNVGLQJoh+
y2h4WFQVPJBF5psYoGkyo2QF7Cglh2hvVP0O3bzwlxm637VKuUKB/wtkTVlWaxpkbmR/UL0sibX8
NBA7IK/wkBho2OMyxJzY5GPE+03XM6SOgNUxBhAAYyqS7cZ0H3AnpEXrDmOi2xwvEFtr2y8LGum5
f0J3mlV6DcEKInTRyhvFyQzKW+QgJK2WvCI2CcU4oz99AfwzY92X+uYfzbXRlXoiZxVw/R0nt1S4
ZzORA85ibo9CjiQWgPj2cuJt+8USf+mq4K9S64QRchLQfAq3HgB/vtFxzpcyPnhpOOfUkK2H4ELy
iTyGJQ2lNxehYri0/qTJgVZoD4HRBV+fjOI2WG9kC2TQJ+XouZHGZ18hX3ThuAt274budaMltRHJ
dSi/cnBNgZd3u4uceZr3oz9tjhKo+QeIn+GHVtiXgv0NyGcWTIXYQzcyEKz0e5H2zH9WUioLXztc
CQCAbNsLs89lC/zeEbif0JwbzV8Mfuoy+g86J08Q6REnhGY6rh+RMcvx811LKB2j57IVPNYhIBR0
LGuVHmt+8zPhQR9qRGmHdgmruP4ClUBk79H6NZiaUzLKnZpmolkAvvyH/+tIM2nacQtXvh1FLrjI
/LIonxAmZH3uzotAKbTKQrh8FInfQwgrrwa9vjsRwLW3CwJo9ZUDC7DkxOs+S0JJK9WNzPxItYuH
5LIbAtTVvARs62wNBj6X4Ba/0CAcF2fo3/7JqGWFTMFMcz9RQX+lZKFZr7WgzHB+gPiwkhBTGvTJ
hfJbqF0xYr4cdQr8+WXVRpJdoTxNccHo3fOVETgqDrFXnhE0qxFubtSAcXcdcF0oFKzaZj9AiohN
mGYApI28XhsUH8B26bwH5c+utWyBwEuUnBR/0dIussbFAXh4AA1VBFCP0O9ajvOsznSs1VIPkjdR
8cfVhCdPdB/uo4GF6v2wXUzhPdxhun/8izefxb6eg/g58Yzk40Its8dCekZkz1Baw/0kPpLomsyc
ug7cOhUUwcAiCm0+tSJIw60JykDkts+DE7aHx5bCaFWqK/7gn0Ti3gsgKQACgmTUdSqrsf1o4N7+
nsmyreVHiUq1yeMP6nZi5Dvoaie3I0sri8v1fy12O6LFlRXYX6qV/gkvhdhdrC15NKd1sZI/Jx2b
TKYZxcV3K9XQAfpkP4v48CYF9XcJPOC5+0rGELMf7x5S5fHWgXKwNpab+iZqPudkTj6Ber3j6f38
KBzqAP2c/hA6IgSi8UlUlAY0i1OhwdfAAQ1r0msAcGOlCOK3nV284SzQe/yILGUwJZ3EpfTMBZXY
2vEnvGULyZyPa09eGHS5STfi5CYcaqO+ygUhRlPxt0GEfDMajD4jhQT2q8ImKx/aP90GpUcDoowZ
90jBe1AJqTHtgq7cbZ9m8ISh6SNrmwr7WIvTgmWUYAkfL/0oTZmjcXlvKinvKgTm8mEzxrcK9Z2h
nhPlppi6SHd3E0+0kLnSHK+vEdu00jmqMu8NvjtwsJhEM2kevucYnyivHnHKW9+rXLSZRs6NyGCH
MifHWumnQrAF+JP0S3K8zYExFuqWtSkqd19XhfBTA9YpHz5i1gpsERcTInRdcGXYnvWOdxHVBsj9
KXa98OZ/PhwmD7FZJqoxp6F0tG+UuerLNRWhls+0i3XNDv2zBgP3MLuuDtMepAG0rDtqFJ7LyDMF
v7o3BrD3xjyJ2oNTNuT+rLhm35btjKF4KFEb+18ZSepW9JodV/gPbMXiulMl7SLQ6wI5iCE7nIMr
QX1c9Iub4wT4f2kaU4SuKiWFs1TTMo+x1ariTdz1KUCB/2hmqTmNEQhcze6LyQlpwvAwY63sTxhK
t/tYf2E2QnBmHUt4edWHSJ2qzJ4I7Rh0LvWp3pAyloQ+CFalfqRUQWIHTriojKHsAtv2nsW+3FuJ
F6A9SNizV++5aJKwKk95hMjEf1P9qLyA2/RqzXxRtX5OtouoyBopbWK+7U2k46POkhLaEjHjj3lM
X8HfQPzjVZFWJUqJRSZdrz8V6HAsk7U2/kB6H//asN4LNl2WrmSLlfmmlGHk4LA1mm7AR0WIwqeW
AIyjV6aNWVwIAAPK0hLq1peWw7KIlFn8Ps18Xymi8oUrBYjE1IqIvQlaaP8f4EGEpC6wwhFiPGty
c8E07NooOFSGEWsjP3uys9srmZrl0kmzKv52KLbQPv9npOETdu4KHdwm8ltMh6ek6yYTC/2k+898
wkU1Py4kuubMRz+19+b5m357OoSOrinlCT5EUcrm8/+WCISVh7UtiwiNi1K+lG1hlu7tjzZf3QqH
yyK6TeudU/3uv7WGf5WycBJfBGijmty9GljyuxdBqi+gKBto+KPv49vvYk8vyuoJGjaxHA/Zsqo5
itHZDn9AN/yAHO6DCha9zKq7bVEIywYKFOm4IRglmrIvDc2+7EMCsnQtwjqcXFMG7tIwru4q8aem
A0qVSNpAv1hIr6dq4QFGUvED2HAp6TYsxs9HpynuEzZiEHyy67ViVHU1WVrhVf+IOsZze/YJ1pLD
v2uluXcOkELGsG9la+zOhM1BuvH27EawW7x4yW/BVYpb3FwjtCTuDWSb+NB6MzPG5ZoEVRCpw3tM
QVg3c3WZU4e49ptlCRerl8+SPEAf90/2vFY8FR0cIucs/TT66taTbhl2REPjroYflSTAy5Mudtm/
H2wBDKSIUVRhFcbdpOc8SQ+E66WiJMXrOCUKVGYXYY3cr6idoV8hAMy75t2tJzCc2+vbfBdrNyoR
hCpO83rh5F/IDWKbvBngT1uZwsaq5BF6+9aBGoqEeUeYmnEh7D8e65aA197+3x+tIUxT8xmr+BJ/
WhmYfYArHuhwgb7DEBVD4hNRLQYAxf8EW73HNK/MHF+anchrtvmStag3s4lSfjanwzPBvQmo7Qve
tggBIrrj7vVQ6ZvwMOp1Ky0FNe7EmqURSSjDdlU6PvFPReBrX32JoKh9Q3mxxvKZDnyQzfpBSl6N
CrVYX7NI6cRlO/XT7BTUpHGobYtB/QnV2lP/T/fRRypLReiNlRbAkP3LWg9ovNby38AOXgDujLaE
PZX1IrNK7KPC8iN1MIGHHzlf6+PhYwaS0FqlEA68Bn09GbTHCCH/zQiIglbB+5qMh7Cagwcxvina
pdy+8JX08pfsXRlhZtENt5DkPSxboWl7dmaAx72kMeoh2p06JOV3FHdoc4HltMnUNPXnyHyowfH9
nhyYVZAc1kmAmVLeq/9L/INAph9l7UUNR80BvCTur9ZntpBUBOz/u/uJFkvs2cqU33iqn41kPRun
Ay0l1ZSm2BO5VyDtDP2dPYQO8BO0TiZmlhVP2TZ/6OMO/aG7OdHB+H1EowJxI3jStv7U0xAbaQLG
+Xn3WUumz8aQNv4nSToDyvgMnlPZ98yLZb06CO5adO+8H7ZbeUFyOzghB2hxyIkKC3zrsfoh2hLa
94zCJDaS+an5P2RBf0uJNb46MDcyOTj8eQ17R/qDYIIOBHKGIp+eMgia7KGIsMlY7VWWnEfHNq6K
cCKfSThXrbZja44OBcGAPa4S0dmlO1yDXub9NI0bjVw0UXIKdAXIk05hlZJ0W5sMli+x2YtDSpj5
Ni5NUzDfXC54sq52eJ9WjG0cos4Zzmay20aWxijqFqB/Fre/ZIiB9EmrCxyGiufYsRocIkhHZW5K
7Q8wFjZuuBFuc2ruaNUs23ZFd2sAGlO31x6FzNaLMr+esA72+qv9gMEEsvyf2onBcok8XiFfUeJH
iROLgXBR7ce57uch/xEpu5Ho4H4K+iKyB3gYQ0WIzThJZGZf3yKFnavJIkJG7Rc5+p3nWTiw1j+Q
anj9+SSOK2GwB1eRboKkHq/3YifYv+m49kZuFH63OxzRuMXYM3TXM9bt9sOLtyD1V/oYkFLzwCto
fC19akvm7dFDjug3KwvG0SyoCJlsUKHUJglffp1ppqm5cv1Uqj8S7cvyz5Ec22xcDn51Kess2yPK
r0Wxsgxm4sAOvS0anxyARdmvNo6BbREhFpxBetAndxwjVFhIuDeESVhaF0sIQd1MN7NcGGs0zd2d
4POzeANEgpnXEepUbm2ldZimMT/Rcry0KPiAmEY5uNjGupS7gPcglCpefRSi7ceX1ApyHQcXuPso
H/R9IuqwCJEZc4bz090oTt9CdABVxPlyKxKi/Lp1Ly9y2X/IYm+SWMCfLE3ZoUyPON81xWZnvc3s
8W1mMQNUYA+7nnqBuBCUBIutSH/32LMRrawoGZKEsYi99Ht2ruQ6c1efJoiZB22Zs4HoTaCJyKBD
9HMNIyy1U2/uwcRP9EXDjLDleUrBIQnrQX2gyP/lEnVA32JoDZu1D9pUf0ZulWZ0zApWBJsVDvXX
LWRcoGhTiNGx8TpGETtBvMr2xjt1AWV4e0nhc4jcGDtwztORsS4H4oRmXWhu50IK5Ih+hbulnPZc
5OLg/Z6maJo0e/1hXBdU2Sq0ZhzWWgCanJYGmmoQmHXbq3tsAnXe1u7lZPxB1HFw14g8qz5nlH7Q
Mm91e97o/T5tk0Nqcja2IEk3ZCLc1K21W6NnEhxkQYCuTPQvLpKx0EISsAKZufzCtgq2BFCxzQZw
7iRO0FDqMoDch1XXfXAtQEFaOW/YdnNOJ7AvzGqGK1iam8ntnZYA2pTWGzcF0nFgfPLQoweYRNdq
wlHxwocQu/yxeNHS+Oy1DkT7F1V018y6XO0aPpqZA+/L/6m8qxidEJg0L3uhVSreK5t98q40re2B
vjDGoxjqjzO/FmEUqOFa2dEKDkylvF5bCcotMgC/9H0RgYBc20CXNlvqbRLeiLE9EPyjot0ZDDLy
VZz5zK5zOwU6+8bfsQRod8JiIMk3NitJ//84/+6gqKprjTSNFxk+frL7bPjsxMjlGsmzshp4Tj/y
OZZQ15mqRnDi5X3hsyH0fltAXg3PswrGj9eEzwRAG1K1VqJIT2luXdH7nABi7GEJW+3tRExGL+QG
UyNRLq7+NzZ/YOCnf8Sgs1clu5obaS3OAGwjN4ROo65Uqsol6x3i5OIFfFzy3MaZoswwKVtAAiNt
TLDH2hiyl8y4LwNEgwPtNqd5IgTrHaLEGyaXhOyBeDFow7YmDugqCja1bhEvdmJEKIDGVdI9gvxz
f0h1XqYizniwXX349EOKRF7NK6ixqyAxZHS80J0oQdYOPyEqVKnvYRV/tRgWWibOG7mE++rBsJNf
WK3nBOuUT7hEyzuX1vcNX5FJA0G2W/dewcfnWWowsBMdVUUoJ0mPC+8fq9yUFFYW6A+OK+3wESuG
6q4eL7Uq97k22h76VmA3rnI6e127EC+LWq6qWCRNDx0PzZ8kVgs41kTkVHxF1BzAGoLbCNElfxdm
zpCtHKAgj9/rFF+f0c+NctaErVzFSNPVrE4OUtcM80iYA1AMAHu+lUFJngjiP3gkSuZlIDWJGmXd
vCufOU2NMSlDijuqeYwCaq7TCq/FcaIlFQ+DM7Fe4tqM/R2Byh4xeGuSrlBDsDPwxZ+PoXRTbjLt
U6tm2rBopipV34asvDtE2Bat+DcYN21IZYGJJtS3xRpJoiRuTSUByOBGY+dRKNOstZt35gp1+nD1
Fe5tzT5bXQhq9m70oufZFsAEHFI364itMyiJ4b7c8hbPzd/qVWUEz9qZe4ll1CZyLhdlvf+ZG8qb
vFmE39BN12+VD3yC/9ud7ChbcL9QJ/4lSnmIC7BvCrfNFw4DDxJvt7LDfWJSSMfXIMTBA9kT0M4K
mV0Ye5fLW1PPQZXo47XD1GZ8h2BNkIWaNhG/Bb3/bUIsJ+pgGp0lPBW5ApGYNMWtbAtA2Zn60O5b
QwsyXoE2yX6Vp3rCz4D3e9ASHXk/q+ofAx3tzA7zSoXREPqbNh5BeJKDTH8Was2NTqXSLwGwVlsJ
yUjeBfGIQiK6erj+Gnh4E0s/F878KV0fh7nH0SIJKRKjZ5wfWidHRafqkhy2vfymSpksdUpfRV9E
1BE4fTTNe4Ae/B6cjyqLKC8xOEtdib9KkU7FoQkTc4/oOziv5ECMOG2fG3+HXasnDGMBq+ZdbasG
BfJpMw+u267A6nnzVTlT/s0FxxkAJehNOQQ571sbDkoaHszPa+4y5hk6+mpIE2VoJFNt/oyPgzgH
v/NyaHbd32jXygbUFJRXJjbxALrUksCINrmbxaUV7NHMFDoiHkmDFsnFVFZtprJwf2k5/TdJYjw3
DxxQCjlvGmfp/lRy14mp41+hBDjp80vXsX3xEfOG1mCzSkLTjuishBkBktMKcOhn9LSvYehpzqgG
f64a8xctBXzMLfYJzgAC7LzeKiEhevsM0tKuRl19EDhBnUSVKChFewI9+jcOi1T/6bXA3jKMzy14
ayrZPJzQGhTjWsLPhS4fYbUuTjXUv/kfAuE9t+Y37njFqxkRlqSJuTIJcRoZSQz1sKkCR9/nlKES
6tEU+n6qXpnLEo+xJsCtB8dPPU/waddFxYMfehmRRGXaDtOPO8+6M6TRQwMOz6ChFqGDSbBz2Xu+
1PsT3KeHKQ5GZKwRyUoMM5EZCb301vbCDcx/5ZBwTKPm7wTTQHY4gfZBzK1lzKFrbfmQyRl0k86B
LtUofTp8lNFF8wbd61rcgNSBfOywNi5VLgvoSxmv82atnDbW3R46G8AtXS0A/+hn05BeIhDN/pds
LIc4F2KrP5kyeaNHjzN75XWacMXULW3vB5SXVP0+LJja3oknlnRw5WLkCHMakihve1f4tdQRClhU
JA7N3j85zdfyvaPSKmT8hI0SbOSXSUpEk7rgo6WY5GTeajjjJHUaVzp4sdvdHdRd+NZSIdFjsHcN
VMrfMpJPuOTgM4qlKy1GTda6WXVX25OBPE7/BA3eNlkoQKXvboOHkspHHMx7XyOZIGN097h5Iusy
Yn7ypRq2VErs7qRDO7DHBe2pT7sKeDjrDfhodDCzuaYySmShOdOlVa1sHBOQIxaSu9FKVvgM+NJO
MH0SzbvnAPt2f+FNf2VjiCMXdp/m+mkSzNCxhq0ozePAeodAEJdGYEf0y1ZVSa1VNYbdilXyhAD+
BCTHO5Lu5Swi8nxXyyxpyZGIjbwjnjF1JbLlSurGpvImVA5OBzF+yvk74hw3Fhg+SnCdzrx2pcIB
yKhPt8Ey+oUKU/OP0FUN5pRvA1Y548wlA9eDEZI/EEho9bMBzWstEIkGOs7fTffvkVO+8sJYoOrP
TJvqDR9kvGuA7OFlvVDbsNlBRljdMNRAwDlj989vg7NYZKtZdZHegyiIJrqMCHBjN2GRPHgpoDaw
vmLSQMgzV2d2xkQ52qnRwW7NA9XHzNHCFzzv283lkNRe6RIqGJH2VHmSmrqD76B+bAGr35hsL//o
htP520rnlFDUyoV916Y33EUoaXjFZ4Ot96gSZ6BDdBeniKHsaAnZJzRE2KEfHArr9piCySOFMquM
WJpH6hXEHN6gvCWZ7F6L5Wwqc3UHU4Vum1Zcoa7MTX5NgUHZZvUdDSkBwt5WHarpfyO1H1LPETM9
kSzDprkn7zlrLSEFbGfjnPy4cgAGB7jA7SXrk1aR7BAX86oNNBkGmMly66y93D5bz1qjqGK0auG5
8V0v43HufxMgmZWRGbyvXUkj1xhGuOU5YEoKGs28LKg2tAqIVWWyNcKBpTui2NfO5BnQfQsrG5Fr
xmtcPgaYBLhAekq1/ySy7qQiWkS+eSPmfUOoTFsEOfC0kJ5GRsQfwKhmO0/YoNynwGboH+8qHlbH
906YVchXneqHJVwM1lShMubmZuUdnEevo3kbvtD5rFGvHcdj/OMQTamNPXYe3uSn0MogB2VTyG07
HHp61JdXmbAeaRsB2AVwoc2flInfEX1UBiTdyZ9IgH5tTkVnoqcCpZVawSfw2KITTIAZzkwqU5kV
oWrjSpwYXLAHk2T1gZdsIQol08x2+ZmuKUMFVQpziTrXzhypA5eJhvPtEW/W5w7O8Zrc0miN2NOV
YvEu7JMdrfjWwC5N6Uf8d1vqidYP6TjapF9CuJeERoE1CrrIzJJwQO7qijFMKpUlLCvcrlwxkoR+
bDpcNmkeTQe6wEl/c6MyltdZKFHQYGVU1AVdiZYo/qWltQ7u1uwpI1C+8arwSa/vRo2JcTsm+oeT
PQsoPp1+B2kCJ3NaoIapuODX3O3U49xCmWV3Ebc9fnzcn0EMtAeAvQd56OMHcM9cw1rSEAfT5edu
y/5R27nmXOv2EWcvBhJFEvJ5hkbUoOUxeoYs97y9qA9LMUrtBf2Kxxs+EwpXfEe2sQsRhVuYtQdx
6wYkmgKlHFESiCT2DH5RSG45TzA9Pq9I+n4B2m0IdNvFjili+lotqH36fZLKjBa2pCBZsVZgH67G
v2xXBM4YbK30SjAYO/lO6IaNEC2SbG9hE0jqfTWhqL6y7xbpmF9nz0XMNC3fDvXOXob3D6L6kpLx
jgx5Nt9wYl0V4OZn+7G2up9u1EUbrJTaUgAOhBBhSAg1N1lvG+VvOPa4HkfZBREmSR2yrvggnSb8
t0xdUwlWT36vkopOCrndAV3s33eGaVvlanQel0Xuvv1cuR8jvZN6Cq1EPAUWYD9C7mHATUgf7yMG
Q2WUxpi1zYNDmzQRxu/BTOEu9+zCBXFhWz0W+QRZJai2axVaTBAXAcnxAzYNgD6GpoP2XCuVEnpl
KjqRZKacsjV1rfdYLL0Rbd3tr/UvV3uTmT5rse6MIb1MHp54Y1YeV58o9bJ3f8H1j/c9/LGd8EpC
aG5mi0OESQ2QtOd/d3rcfDvggSTY0SmZLXuu4jxnHQa0v6s0oGiNsxtJZykd112atLdH6T4+FMJV
RjVHBMS3B8wg6onVMvCdg5A8u/1WUP2ocy46/H2yi8jUr/PPF3NFCjohhg4C9idsXdwDphDPIFG0
lntn+8ErP6ml7r4mFW3R83tV7TcMp47mub43OW/OrecEasIjDXIhdi9TVwP86w5ntYs3Xgp8WYQI
bM/Zw7whsKuszKoGvgiQHSQmXgxPUOpeJbj+EdW5IbwAe/figgzgYQAoPJ0AycghuqOa1pktd8Rt
amlawP51ljl8pboO1NBG9gJ7Y+bWUnzKJy0pbZ2qX5r4HEITSrYZwrFyClJSuWlM8q5pJdEamBLE
PqfZmi88i55d6y4Tt3BaSQGyAjaEqUw0LCCZxTYsEpjL7ieOIwyB0MQ91d/uE3CbFNzAY0gkosih
heHKden1MPZjZLSuiIN7o4WG7YN5VedRfkg8TM2IYbGBS2y+YJArUkniw/SydZOSFYg08OjBSrDR
FZKYFefSH4hB6fstOjPO1MnXkMifw/MXB1RxrMcmVOjPSbHO0p+TMGCSItQLo7MTu9pmdUStU9Fm
NEJkY+fsRDhT4/2IJyZCtYBeo3D8nJs4yvgk7HoElPTNc+ds997lRMu6+uMaOiQAOmMzqkDVcDEn
J92f/X0j98ufBRomKkH5zED7xeOFiGCYmH/C8G5pH/4aawG3ry4vC55JAZu7edqaGBhzvywBA64f
O6j79jrRaiQExL3j3jFpiodjnXpmi2Wyrcb0rRRvHj2/nSLlalyWl7DX8bZhJOnpL4nIGKpz4eOa
7U5MPU1f7g8MsCswR4hOb6LPbANa4B0LYguMhbJeTNlQmSELOg65w/NfeIWyrqjMF4rGi4GPC+BJ
WlwnkRL+7e7EYaosDq/c8IScNZjY6M5bgY4PRMPFRkcFrTTE42rellnOqgvcXfULrmnLOQRz0UPc
prp1S02TEZ514UgsptjbyinMvq2BuDBnNv3KYrQIKY16cURjer7bVs4y7odvzmokTE/U/X0XpSfw
uChnGLldiFfRrRISpf5W98yCk8XUX0+ATzjTSWVq6CqO7+FE8xV1Eq2CHmcbdkCBKEcwjcyMESsF
x7n2WOH0dhXvDgztPdLjjVpQPE4j1xUVRbMalSEbWRScGmB02/Yv0N/TMSh/MM1D3aVpPy6GV6NL
Txh1yvurGb2ka6RihqJlUITbXpI9rc0GExYRt6JAVticPBiFRGY0Kk4smGSW+EqmwXaGuvR4c6ty
JiOdEPBnlWkv8zU0R5zK1m2i9wBMHOzED/N2CcdhHtk2vGaI41W9WTWzYGcUINH4udTjvInYOJxK
+Qm0LtEuxywFF+GbiDsH6ry5CQ1IZbjphDQR7NGMLO4pqaYvCEyN7TpKV7h/1dhoV2nzcdLz+o4h
o9Hvm3v+UUArnFOvr5/EMkUIjCtBGTiJNU0O6y8AFMQsHc9xcI+p37mNjp9IMFIjHPeK7amOsrFb
37Wp2YMnNLww4725OVN4ywxxaoGk0ZyBS2OgPyh9TsdU7O5oJhBqePiamLdAknXp9XXtOwLumbaM
sgnPrP36jZBJN1c97dp0hK7/XLVsokVCNeryAEmPETx+dnhlqQ5MXgvddQ4V5m+gmt3FJ4XLLgXd
MBxibL7Urk4npm9+R/rUsn1sA8rq3RV+Au24tf4bdjxUtqETgw+NPJJ7qc6zxUFfDsypPiNbe9/X
oO9l2kQwY+gZorl4+CuIVtnaGZBgPr9bFNvuTQeV07dE8FofsUC4IY3RjL1jxgyizKjyLF7XV+dj
1I8WW27f6iNJ5L7s/jNzRGpYUhIi7Oe/4xmrcejC7HgMblan+U9uP5BEjIKHEe1bPpVqfQYHn4Ix
of9hbCImNbByGdyg5S9J8QAUjX+/UzXvZeabZZ0Ew7NjnM/7q5oIcnYlEWIBaOMpBgIucagMY/U7
unqqKRg8svd1LUNj6zyOC2/J+P6dUtGdXrW5PXR1/lgJMgbG45zD0oo8vuHgBE2ZX7Kzi6ahpeeM
ph+DJZ9rcbprDs7rteiXIq1BEABqn9MCEDVOA9a8zy9FY05LpayEglxHI+Mj6e5LKndB6yJDXDS7
NamX5plfnJuDKAVmgzLRyHjiAf/dutSdy6TzMtIWs7nH0rQq5Y3cM62qaGe5L7RmEzJxsBje0Qm6
lhzlf+Yc8VtHQpSNX+Y+wLy9BKf1lK5cWrrqthNrKmMVRqcLtfHV036As86589k8GEMlLBPv7DKi
pranyruagm+dVp3p9eUam0zvzNFxetcrLIzyk1Izt99Bsne4xq9g6Pxj4pXMDVa4iaroApx3NqdR
IR/NlI+NyNJOieSG7Ww1+lkWP48Kwv1yHtFlAMAyE2ar6Vr09bmc6Io2W7T1isBkKuukV2TLfu8L
Kl2ZKTipznvVvQcSG1n/h2xryRmCVojwLiePnVqMB5sfeCvtQPvmsm11O5SBqSk89FHHYdYGqEIa
MHDHe6+H9SSnv9X+iHT4TYbE5eSWPqQqt1g4oIJQ2AOmSY8QfLD0qzWtjFmF+R97BZqcylzgzeMe
7JJI+KhzQ4skWHQ2TIIlsonW7mRg6u3bMKiwQPDz9YONpsi8cjOQXStsuGmMbcbNkYW5DhT4PPLC
mVKsgTxZIu/KVmAM/uBXAOfxf9GJgzLe50dljaMXDeOBbqkI4Sa8qUPNhKS0nfjnNazwpeKEnBoX
uuunoyKNy5JSZT+NERF7NnVCF5TBG99tDwa7zWJKE1Ec9pQYC3VhjLZ6dXmvUtO8uhgVmCFGFnJQ
nCwYJgPcKsYyfEV1GsTYqG/alh8H+PbqPTaeHgF4hYI2DI0jixatMwlsNIwYPNxxAKnbPXJ6Ekxw
VqzYnCMAzUjfBAWWMTvMVmwKcw1E4aht9m1CeISXAzNi5AW14YmYKkkk3osPIa+D0IgmpIyYeMmk
QXQOtawlCa8d/SXYz1TLDcoq49dFd5didafqL9n9mB2JNmASqzcQKl+UzNH9bWEboXkMWD1d0hLu
TkWQ3aykyo2eEaCizoXtSO2X0uDWtVTy9SMdNsLbZXXoHtFuTaC8AQJiutsSAlRVMyPgrtbcD+fp
fGjrkXFjGpQfm49ObTEn00wqnITBP4/yjVI+FzIV/prQN+LFalCQjCo5b8LLjpzBsLUIIvDKvo7s
KKYedGq+9U/vOeQDb9bm9mzMHBlwqkEXgGTpnnJ4cmT/PRoKcG5FAZjXtBy/XyWMaOL04WlxkCo0
3+Wq3702trJF8AYwqoXyUJ6BIEHBqFd9WpBkbRyP3kmAtEH2n90vbsG4sJAXkaUzSA7BT8GFHo9S
9tlCD21h6fc0QYMMKXUq7y/z12MOm2Wf8tBTm/uCSMzGcR0cynSkOJ97y1Cvdbgi3eIWXpwMsxIb
XiNqmaKUVJOurXcR0g4IC1KToerP4c2obLXL86Si+dfYkP5B5OoA66ofI4BldXG+In9HPR2mTkzG
LqmXLs9ayjvARz1EWKPoZTQBCB/e9CkbgwT7xQ12sTVCI/ToVsGB2WngPRxUwgndfB8SMXbuAD39
vgiAmZpsk8w1XuGxKI69O9q+Mds+kVLgv18l5hn6QHWGbdWQDB3cUIoSHoxMAmvfl247gdk+ZdtQ
w2dSAPulUHBAn8Lds2PFgFQ7pFarVDqx2cpKvmLvkMYUSbnxudilfglD95VydiOiffbSSpIELTLx
YAiESIXg+nRrQPLNeyloi1LzSyN+jOaiSNnEY1bZktZzISltn1Osy0nPI3L+cvw2agyA/iAAAuX0
3dAaExhEAyBHsPd5ZIZroza92IYJX48xD9PKWP/9uIVU5tq8XbQMC2GIz2HiiuWZSlFnmIPhCM1Z
jyG1qe/I/ImcGOTK3JWuKsVjbidYGi8b8GQw9usynsOzxx293g+0a/Nnma+XLWeBG1Oegs0PCxf4
IUpfavCAkGGonBzHaWkqk2fNJ5YoJWOQIOsoFDHnoyOAtbsOJoWzTx17Xm18KWbw7zOMtPjJE6my
LEXNjV794ZiNfjyhCnx6ZsSWkKQLH6kXs1miwUEVEekTU8HcmxQrVLpdsgy6dY13WJcmDtq3crkl
THrN2/w71nAveLE738mDJxwF7v5vipRfS9/JYTKkvviyTDuTW18iH46Wo1+l0+pNOkxqnVguVS4v
ayLrwMGN4jn0oSgmJNPCIaNxXhM23PFOuJ7ACwZS7AqrBgZgeGzYv3OIseDxZy8ppGmrDwAVqKYK
cXAE7dugzOT/a1EnFY0HU9tIkk8tIKrLRqb2MgoN6hQ28wWY5erWXqaveUvXwWQWmwoGCnvRFxQ5
Q9yWm51tCt2iSJG2CAWo3uR4fK9tXx4DwEU/5MDJfehhg12JlUfKYGeB8SizQKedBFjzmeo5b6wG
LQQ3XPMjzwG7EhSG0ZGDaS/LGwalfsP5AjEr/umezCWBcHorzYCdkIw/L7zjzFdEdx3hP8mX5AVm
k7ESgB7527Av6tNEU4xZmq5RcxVckdWgu/V23hQPlPVmTpJ9QkEcKCHnualZaRidXAIalQce6ZvH
mOTWpes3z7JSfpVyPtA/8DyOB00fncZbcw+Gqry2uy/QuUTRKgOv6TIDo2Jzrdk6/cUMm5kH9ZYL
MmyXou19pUXBFHaYxMa1VtHHN2Y0s492ZdxFrXDVj7xNTzaac3adtk690dMto1EOhuJMjTWnb8WS
XMCSZ+4SHE2WZp0cGucx75i/buRZBsyQ0dAYEZ3J9/PUdY0k+igX84KGRIdSqAoI33Pijqp76R06
hkNv8a9donk2lYtSUfdNqapNEPrH942NOzOV5M3HRz4JUwmnkys7ML3k04/0IhYT6226xobcSgg3
tFbae1RD1PM57NqRVWaFRJCy3/GZIQhoCv93Y3NBeLjgF2hOaWvTomHVgkVq35K18lNxbxirVluk
GI7q/C0r+a+wP1lyG5+yUuZZNP47HRX2wIaScyD8raSCz2v3F9bp1d++YOtG6xfqK55YzgXpD+AH
preU0fpDqTup/6+UVmykcDEGKDKvskX26hD4hBkc47sOFo0takzHyFB9Q84uEosoUhoDZIwFD50f
B2G13NhBgheR6mnsPKpUQZX+Lq31HYNqx9dPJuZ5VsSFmVux6lL1LLccd2OEb1+tzCus4USxGnL2
D5YKtwZt1DpiGgEqIb5T1aDuEk3ddAm5aNg+g13C5qx3BhjpbSxI9BDiwsP2BMrNs6Py3XFNR3sj
6d9LednABEcw3Lr9dWUiTqAOJdAlTeCnsHyS+XW19kg6lNTK37GbPwFxgQxxktFtqItX0OJVDw9r
13yi4/dvpeWfC7lPexmzfMwHjKZZtdq6DBaDpzjMw/UIemU+QseqlKWA1TgXf636R3yvjwWFmxtR
jUULRzlhgam39QiEb1BOrbTKURO3a9OmR3g+TVhRbgV3+WBZ9y6LVXQkNjypqyJTarFn9nlHVVF+
9abozSIFvsZXnJd2IeZAXRZBlkuZzovclI75AcdOw0hDkzrQpYdWVfuCzVq5GlAdTWeirVdJ/DBZ
jQI7XWKlW+xzRTct9BpZbKsTwI/kWO2hm+ctZlqHrKCP59BhspCH8XtvR2UDMjGUHzrapCd7hkko
h4PmzH9nDoQpHgf4kMZvX5pnT1JCf1KiJYSGPGNUG50pNWon1R1VOAtVn/um0l9fZ1J+TkeiI7rv
8IP0NvYEMAJkxtkTlTVg/jZiuCZp15+DFtnaQDlVfCC58GcHVJg/9oQCL8UwGn+BdmUDB8+t8qQO
hOtWnHFVoLWkv3+nIF26JHE5HnTGo7cU0K4To1TAOlJuJxWlB2URJjAs85t3hLOzgDzM/j9pK8la
aZmIN5xgmxvq3wVQVK9bSft+wrIW9Oi+4clSJRegdabOKpXqyKDesgwhxu5LVm1Yo8NEpLxIKSof
LmUYdzg2nLd/XL/5cWV4J5KI5cbUPRfrmfNg+AhX/6X4SGzYzhFu9yuvnCWKT9oSyBj+j0/W79eH
i8eqDNJBLqHZeXxqs9teQ/SsEGZMOv/y+qOASI9Lz0pPKmzeeaje8SXZruMLPmPzQPf9ZHexiq9a
ELn+w+opK9zXsN+ogOhC1uvXXYJBJKSKHrx9RkW5CTDgo0ZPJ8Ks7ByttkPPjeSzAh46v+L5KP/f
xk38E7pGknbbcQo2WKN42MU016BgcuNNOmDsdSYf++1WFXDKDwnA6gPeV+sMVJGwU/KNb07m6Two
mpi439XO5vm13gIySrBxtvrEZVd9B8w3BUEGkD3aPIlOpX/Jfc44QPA2/07V8VYup47XHasd//fR
PgF+tvOQNgO6csVPjntJ+jH9eP5CDph/VuyNBCrKzn4vRu090vBe/r9HSaicpOvW1bb3Qq+Bv8K4
iv4xphWVuJM9TBI8RRmIMazZPp3187ZFfR1hms8Ay9ff+B4W6Gvx4INdsDsNC00KUadpJXF+m/5t
fi2b5XrP0S5HKb0eyGUka1uPQRdcTXyfdHf+JYYUBTPPDgP7jBjVwMQ+0AhNAOxpwvv8Wy7mqUTJ
ijwnQcXI+ke03jTcGkpUvyL1C4KYJFVQ9Je9MXDx+wLhYSiMMd3hgRG1ebhDvn6iRYu2tYwCquNf
1/TOxwpsC0kzbE6f+50zG7LLkK5vCl+9qFPF30il7puAlIeUUJy11UdVn41mpNsUraKdY1IXmHdU
m3I6WRPgTpAHe/bmNl6OPmjauRDvGD6q/bdm1nEyEf0eMrOVdcEkKS+OvqSCgeeQxyy/idqO1sVx
7uinhF2dErA7xV3bEs1hr21NQKGpymMeclG7jFJokUaWIpepRBqR72O+UljBMoUnKzzvKodHRu9d
FPYj60fOf0+TpoR0p5N5mNGFv/BXcbzN4nGhwu4EtJjZsCMgyRGwnKWRvGNvi6c0zWXpJw6UF9YG
k5RKFC8k8awkFVSdUepmyeZIPG40hsx6dS+3wSuOjHINchIYOCnqo3BauLMh73LS6eC1yfLC8LNL
ADHHtnmCGpSUtkNB9ekoZ7xeS/PkDfFhVCz/4D2rNLYFN/CvbUj11ZzRLtMkfGctfkjpYxyulIPr
AJZqYwBYxHWtPnsjtPL0XRUCaKE4tblpJeZlWKMseACz7pPDD1yrXO3I6SwT9o9iw6B28eagk0f2
y+YoR6XaG7LVXZD4NVkd/TjI/6M22HUJpZ0oomlkWkAn++J0ZWEpHTEOB1dKLTOn8l5eqq0I2QVa
L9KjIuM7Vd+I/b2U7y7K9qvUNV3HxNSGYHNsufLcE+PRY7pPEy42btSNaeMoZjo1hgkWVUMHVgxz
jEpJcFIp9iyGlUAqeN44h0B3UIdAd4Y4mwCU1awAaY9NVeFxRVaDHb+98TM6Xsc8GgZpMXFGEveO
n/XTCQ3WLG4EBICmb2p9YB5RxsfI5LfetmMXZwg7vD5FeX3BGhWZe4qGCjlAarI8umR4ETDlFxNw
fllfm+g5nhhTvcZp1rWneXY5E9fSX36wVmNcQcaz0+JLO2CNM7UA/zV+xGJs3csd/1G/3CudLxw3
IS/Gsp07F+2sqy0UrvBmr2GC2GRLDotWb1X/dhkRE65tmzqFxbQRcHxmRkJB98q5MUQOexVOiUyM
52hqvKajYtG0/QXknZqqnwhoMl72fbXmbqDP/YNOaT9dv3q3N/5660ARr8zG3gDTv7+maJL3w+NT
JOTR1Po+cuCHrw8JqxDla8QrqcuslSiB8uvCKaalUtmgcOKKmWsDDUXNQKowh61HKPpklyjkKTG5
nuNQT0l8qTGe1J7+Wv2lFbDNr/7xbuaW+9OcMSqFYxO+2+pcS1phADYp37ZEwa7ecXaTsJMnT30c
e73aZ0FqpToPvi1TsHvnmodRbqoUB+h2kCAi4Uk8S1ht1FdKSbvGNZv1aU9wg1m2SrRLAenwegRN
E/rrQl8tmjF1WUqMXz9rj3bJ6zFETjRNMVMyuyR/ScmCw+2VTUfWpi8Rs7K2WiMlnQm9u2a4alHS
S6KW+JX133/DzHGtThO8zzqi1ywJHJH9kLvsMzcRhtB9jssqV13laOrXf8QJ4Nmkze4jXl/rJAY9
/psLv2dJYfSe4+3duN5uZlatprIWN8MipHQ9TQw1OBk+wB6fPfhCGsCJJbwzHlixBwGE+Ze+Rcau
ruzee1p/HsoN0RNBay7+p6ZMcHOaUrg7hJwMWYMVbHxhMro/6SUUGr9iyXZ+qzyx6EbiGfYzv0Ih
1IQxOFI+hMG4UNDF3A5vSkt8AbQI3mo1i23+NRxtTeTV59YsWEh4rbZrKQBDQAV+jM3ma/pPm4bB
qlzoC/qVSBgu1x/qMwPwZaWg9bkl+5AAKyEPThQNkgX/9sUa3677OkjB/GJka5MI6KZRD2Yt+93r
QeK1yh8c0ykDyBlbSOt2yPNKiBrbk9wpSHhcQP2LDDAQQUd2+/q+yFh7fSN7un7tmVsxj1y/ueTF
ekQQOaAqTms2VcpWRlWnU/An3J/dmcFhEkC9CvPvfYQ/I89Cdm2Votn+B8m+xsTsjD66uJiDhc88
fMcFltZoNp9xbB7RA2VWx9/oo5Dg7cgq5VPuKvbFJu/HC8/syURX3rYDMANtzmNH1H4p+MJ+LKEU
6Vs346oCqzAPbnFUcFe0DuwQI2l/4DVIfvpEoIrVrs34Y0cSC0loY6bqJX0Yr77J0O5umyhLYqjN
9C0j81La/+ueb8S9L7VZBineqMLk9A+EwKVr0UrsXW3oAJn9OuXl+jr1IRaegMC/OZgGZRXHP16y
3fShEnE+96jarM/4SPxuBxQ2uaCT4JiXm2scVMryxRh/qQuBsKXGGIlfO3tKaMMKP+88aseUEhLm
sQfERzwTAp7T1vHVQ2SGpNr9rsiR2AwYJcqJeX+wGrmFgWGbrq12Zl2xndm3jJULUCct3U5Vrjm3
48AeQGLAbdIXINtoY/TM6yjxMidNwMeEsGD4l3J6ECWXSaMLRqhxRkRpdkFKlPfpoaKP99nQwadh
wyiHKJ0WBqHRVpT3UIalbmTeqHC4ywgR32k5QPvk4RIuiIW/qfZJTShdsi/JsfwylEFNF9yVs43G
v7VTIZ/w0UlXA79dvbsVjobco3RNDfH01Q6XL1WDBwXdNviIyygM4F0rrZ3wKaUuuRwkTh+I9CpF
mF43MWf7XO5uYb8f5gjX5wFRFHMB1H6kYFb7a91kJo7+PbOit5Hnp/j/V2TBkEmJEtzw2goYJtlT
8yMJQWmu7aOTKX0rOJoj1Fnv+bV3MyOhhNGbBSEghj04F4AWOJSN1YHny7zcypwPEorVU6kWGErl
fHtYSYRgg99++k2KciBNGyaislRXRelW3G82WaMkMYRBFLPnOfrHeFx/6yK4fXyvQ06G3rXyaQ2a
7Z6/xW7PIeaf7yr0KpYdR4rbgfj01L65Ed29nHa/nF2ZXSLfBXZJAiOUK2m4WysAEwne+ov5n9Wm
OreA/sEWfMhn+v+QeP5JakcsGhu+jyu49zG7SIkqdcnguRjgyZgqcnMUBAVdCDGaZo2PTtyFM04V
zcmttTp34IHm9rnVkDBtN7dkx7h6xt/II4afzL0+cY7W7kuDn97nwapf4ipka8lbI6Hin7vbyM20
8rZMEv5DeY1/HwXSaHsY8qPeWEZsxD7Pfb0+TMkvuXGrOxFlQ4uzp7vcyeANN++vaf9GtQfBvU36
RBJNtP6iO+YwYpv6+qvRAST3IHcKH2PzcatdtvRbMI+7m2qdrU/CrJpLdK9vdRUZ8VUovsPEe0Uj
wJvFsZMuF6ZBNr3CM/v2LmQ5DgITJSdsPWOlMoRdTHCrX2g87DiUHkHg+YQNnLSRSFJeplPxjLoM
b2iIAD6lBdDOqOipNJPJy1UTl3Pf4+c1TzBARKU2oL9ZEbAd++4N/hcQwbfO5F98I25A+0rPz1VE
m5tCR6nT0HYM/RSb6le8OIc7zow7leqNix4LfOqiI1nwA4zwsJJZYkbBbQ/SKyw6MpuFlh8y658i
zjYtaWgt+WcskJfnB0LUytGENevjkqWL8s4MQiDe37qcMTmEdi0re38DgFdGD1GM8R9u9TIzGduJ
WjLbFjIJaBS4tZMRW2Ohm2vhtOt5v7vpx9/EiASWk5ikLHk85ctBF7s1Nx172FLpfS1M5ykmTAc+
X6V02sRF4n2d3mQ8+WGmKmOpm/1oaELnlMytJn0oM3If5nXhYHNqJ9xiHfyOyUJDvUvEwl4aUPVp
L6lPVhYkZ27BHRLD/qxWdfeCel8JXvUt2TgM8pTo1xvpUHC2y4uuN3FP42WJQPqGK5BMRbL07Y+e
LFZj4jYmnxRRj56b+LPj3GSTmAQPM5ogC98qMgu9fLG9ro4s0y97EvsGPOk47nG+Ls9Q5Pe9WWTt
2lIlksZXiF9qEKDOvHvJf6es/CrWzp8BZ3tO2vFpd3f57AaTncV2mV0kw0OptWvERxCzH7fFLciB
MS/QxYqa/UODsNdiCAXUV11PdSkOs1PK1J8eaZq9XMGdd8f4reZJMwZPsbWX7G7M1wWc1iPeXWUA
nHVJehlYy1YwsYq0jsbBUbT/GI/I8Bg0e9+SIACapyZ/Y/sV27eC4wux9p3YujNu8xi5dFnFThPv
mgfIqMfkeR75JJpLJEju7byckUuCGKACW8dU7FUZ390YoAKC1cAllTYwPjQHNEmMq4KN/Gl+mvDb
i0yy38Cu1C9xeTbNbYSj1z3fu0Z0DwUST/QNRky7m3+I3R9Vdzaa3Z1nbHeodlSIgsSFIFu9UlC2
WRrNaWY+Gb7JLtK/P5GQrk9KVUo1qDQzkOg6uYXZlgnHi0tZafwUm4e9vEQcBqu7nRlerD22wnVB
q5Rgd/OzMbmS3o1d3E6aU4zsWp+mHqKV7fSf7wQz20693JEiYabsiNlc6/tAHmSia2OXHYbtp17B
9oYkbppPYYIU9G2zKyWbl8UQisd71/yN1RUaXWrMzTbf7YrYnBCP1e+mx3L3LilmAMRzc+iDxIjp
r4Goqaev4sT98TSrauzXiQN+oroLQlLXTfBYbfzLHqAc1igtm/M2Zo//nRU8aIml2+LHYg1W+gFb
yyK1t50L9D14LQnUSqpfe21mz45ltqz/rextRPUFtMV8dbGsD5iD8yHkmf4g1aYk7zt9tCDR1UrQ
r14rkf025F5NQBwypgUCfZDWxQcj1QpSVVUVbxYSyOVHS0Kq2xn+NEfVHMyg3WgagX1k7CoHrxY2
gPDj2MDaYUYGJRtyiIy40eyBDOx2rvVybupYFdX50mTZBifrZ2kcOKUrgsxFr7yhNU4QaXH2xCHX
ysqaMQHR85Y4t65Cwtx6N3+68wa3DEtdBm5ZB+QyidfN0DuCWLt5FbwQnjUU3mSNefCY7IG+9p7I
yCgaoLuYlPKH5lj3NME67DlZOO1n35AcfOTMPCWfrrAOg0tngEyNCcVygW5IwhrKl8IMFhW0HsPk
VzR4L3NfhL5cns4QveF69EAF1TfWv+7sjAF7jZ2OrxHlEcYeccFf5DhI5F4yPJgNCSL3zce9Hn98
u6nYw8zHeetSBLXb+eT0nVCk43oZBxAo3S7oy6YuBr7bl5jAYpbzuJm7NEuO5lxfB1tLYnAJFZCe
QFpjLcBGhYW8m5r3tSJMBzezgCxGSJGi6WOUBZWPo6pBFIlnIFpc4xstPcJ4u92BbNqP3yg7yUr9
ZSEyDGP6FEhZ6uVareaLr9EWuEIlD43vtdrlurioqz8IJxmMIBKW+hpWYficzjGPVW5TOoV0wnaI
WrXrHoZw5tN1dx2mMvkTfOC3NW4aO5i298ypEzMzIi4t3Nif7IDPQhufBZAIaEnQ+Ovi91QaHNzj
2X0cjmnlQED6vUh0JEs6Ex+VHSU/MWTlOO2MjeXzNiBODHscDCHTm+pLX0qawzz9ql24u5w4oHw2
OncTirD4Fxu55K586pGjeB/HZH/p3ACD83aFD8S6zxhJvw0ta4qv1ZpKh74+S+FmItEtscdY01aN
4N71eYB69F9nGVfXiWIPEXI06xzSHRRz7Olh+5erxx2OFnew7o0ytTWcgb3kPHO5pAuPGlqS2kYs
zkeX3B1EaUDMTUxXLqX+F4j73bKHM4YYDlTt4OP8jwycKAebZ1p65GOgk+c+MijHmpDVLf0cEONK
0SngeT+JxbJNr813ktfYNXG1fj8iJzGP3fT7hx+eglb25qUpL9qyZw6msYh28uEl8aB5M5tA3+qh
lmV9Xmikernwxwmj0MBsGln+bwzgMbjBTlRziUZ3wudKeSUM0Dz9Bc+6jGTk2Uf+mb38arprzIk2
bzJ7qvBFQJ+6C7CtSwJibaLi9EfH6hY0hwk7EkMbZKLuTE32BbRveNR3HLv4FbwHt/sY3h45sChI
Wy6P1Xj72AuN+62dxm+eGN6fIVq6mQFnyl4wDRwGBF4XndFW3HL1QBvPhyj2GbCm7ehZM5/7giYB
YQAm2LXEiG8NTvJMNjf9sKZy+KY2pIUNb5+bMMk1BfUq40e1aXIMtwmf3bgPCQxfdby6NyJC+QgT
OVrEfU4BVgykOaTt0iQ4Iu/mCHbjEWEpIHl8oCE1gr/buFYkpApAK94UK3RdWV3CxgBCTpmDK0/O
B0Vql6hAiWgmDZGAmJNRuLf62sMirL2/yNI1tLHxNM3uSbfrYxy2wtyCMfQqeC6ci2j5LHXdLBqL
T0+7DdeAJi0WxnEBQyGNtCdTKRoLE39qOZGlsn2uiQYBfrqCZgsXcdidNVB1Fxf9fqUANjoDZkAG
4eQhvlPWXRRCxJUq4DWI3Gigkhp4pKAy56ttkT6CYqPmLrl5W0lLvjk7kEwvsOpN3+F95AwMOCEf
wY43Ltr5vrP5mBk6VMm2S8xzLZjjn51ZUIxKwFnEvhl9bK7SJxpL7Zwuv9DzvoxEEMn7cX2RhGEX
W2SOigdSIje5MCk3LEYHU3d0C50MrKsee1MmksQiaZHKAPZfiQIB6RAYmmgCgFIdRPzvoxp60mA9
kSo6NR28lxhql3Eds2H7oz22DF07tnzMrCp4+WjmrkK+7jWwupvnH03W9VE9OcVJ6T0sX+3py9dD
bFAQ62ZIgf6+DSwZUmkDLcOlsV5mVUx2Y+ZtXJKr4Wvx5+BIbFK0MdDQhZu2g0ewWjcDO/Q0c/+o
Hv2SJfdB+RjDWVRMZcq/c4l2mtkeyqXxNUuXdc8qTV6ZzufdhRNRdLsRnEAHLAWbXTuI5EuebwSa
18LmDS1qR5K85/oVnAULqA1fLcoytBtDx9nQUEyJS7+qJCutIxjYALyzbVHNavQJm45T3phgh/ox
8fqVXFkROnvxM6MLegcIUg7yWLwOKn+YbpIceY82nT/0kdvo9MG6hAqhA7agUssQAgxGvPSv2RQV
Ivkg1C50c001swlYRTg3MkJd+ajPUnE3hLqjFvDm4Kw2gwsFB8YfdKSR2yyelZ+ao5f9MzSIK6bH
Htia6INPAFw8b0eYQOVLQKuR4g7FsHUBKS/sIlA6QwpC7zaBEITPsEHHWLFcuiBK8iA3e4BzBqyS
du0YpQHapaF0g0r6dtq1Yoc72DFDzDTC0znTwW4quSsfcfniASdGoyhlw2zfu27NMTS8terHdFSp
V1L/BZR14dMf8zINAD5jOmupXTFpedQj6iksUpp/XFTRfiLJANXmZgffx2zxIm8pV6B253DEaJB5
tSFMYw8S/q7XpugRZHBl1eP+megI+6Z3kjAqFFNMRt7b9NTtv0xU//8GoFeeqEwd/DsXKQPseM4x
KdoLLQ7ynpvq9htFcl/ERrDq2HKBOTlacl3L+GPlBASrZLwqHJ6RNFXVXtMUlldSPyt0hztgUPBE
0O4Je088ObwTKY1JD6Lv19sW6DJeM6AHr3uoFLmYYnGvZiGIK7VAzIJxUc9tpbQTz2ygBRF78oyA
kbVy5sj+02qZEia3WK7WRWOYvUsuLwkLHb2Ib67UmimCjlh2BhpsSGSLyKtNRXCLfp92+XqnoBl2
ig/bVtXqyFwXFhu0VjDDATU4rum0Hf1x8kOi8JvWFPbny3rJemzyMqp9K8ecZ9moetyAVZ/BNlYl
nQPg9wpdAji7CfNgl3HiN3RnqZS9fFkVm7OXN1DXnuucY9ZiL1M6NGB0Mva5XR/4oRvJWULh9Vsj
OoziaRrnzObcW3TNT4RWEyrmFWPIJ1xea3XQLNJ4vPYtitv/cOeCkomtBl+yQTWUTuWPIXbEKrAJ
dJd+ECQ48Rv/HJD7e4Ttkn2h3SkqSmZe3DLRIQLKCcYD0h5R5CFd4jhYhcW8hVXL56kUezzVr7Uc
u4raA0TfMprbhsFKRCCzqlk75F73t3+Ckspk0apU1SL3MY8IrYvW/8dM3yDy9xMn3j09YMQbh102
Kr33+pnsTt5puj3cgxlyogMsOIF7inAI9hHYRsNBE1JSqtDGUOXuDjNz6xgJxZwAe03YpKEcb/k6
ttzpVWlfX+PMQsODcWd0fI7e+uS6boQbmIj7yyTgdmMehu+BwVNsbcCVNYLeIppempmoRrh0uFWi
Bgtqnmr4WeOan3UPelP38rzyVV6sHvF4GqW47mf5OIyZ2B0uzVb5Yjz0EKQ6vAqv+h5HRRxYHTRu
Pda7ZwDwTg18FkMG6UkztBpxy9wtE1yH7f13FJhBcDWpmKX1fwGQLEiPUwvuhB5nGce7tcfx8TH/
RlrojZI2PHxejCDEbsXoGeVvo1XiK7NHI2FlEhjUOZ/p0VyGOfjFgBnmfKEQXFdDVqGUtPrX6b+w
6Nry54BWHUhPHm5hTLHLP0UdO9xwYClnNZvqhLNsS0+3xg7ZC2pOBMmPLbrngvfIQpJUZY/HyOlg
l+GcH6+rSDyLcZwlRf2SX6Mix+nA4iIT3wFnYa4VhLabsSOxGrJ1+TaVyOJSs7MybaUQSdoG9+QE
kXQaE8eGQ7cfnL0kMfStWlpJKKnKUuC5Kju6LR/DcsyenF5KDxcfz4ImEwS0n0snnPhX5fyZAhnV
eFvcqpMZQ7ufAFLuiy9262zYAA4B8EVYoJ40kVJS4i22Xm/ORoGLB7fG4r7WU/Twxp09IAkfRmgG
I0ngU+taD9Nb0lwDNe72/jVCRmqOs+qEn0jI+cqVT2j0PJslEcX8/pZl7MF+aDHYcspekXHc1UL7
2DkqdLiNyr1Gp77Gp/PXVgNiuFZS+AECKu37QgmzRPuJ6NAlx3m10o6Sk+NlsO3ijQxYP/fGNSfv
pMzZuI7oieEk2XpOzHCsj0Rz7KRvhOAWPR5RYGBKXRHsS9QV935zXn1/1ULIY3K37VpDwiS7pib8
TmUMyB19JAx0VLEC6/k1LrIo/whR6fLAwSU3fUfUzg8mU3iNBql/nogUuAOXZljQib039n+Plr6H
v3V3I3LT0iHMJ3CZI+O6jzSLwnKZcylmsPYi/TUBH2cuK88fdC8YJUhhPrcsQXu/G3Vi2O9sajmZ
lBbHDIJn8pkRXpk6lM3wcl+kY588J84/UZe0sfJL78rw4riAHCDZyBeNXP96lGcVb4lixVoskvFh
bDx4tVnUPy7xpGUA2FPmbUBmBuJ3AQ6C3YzQORind7sEomMBfiSQoyK6dABOQd15Ra/pSh6vMmPo
DyMYW9pX5oNz+lija/La8vNmtWnyjCR1iF+OJfSsJFHKmhH14D4cKdpR5mEHna0wtDcfs+t4//4w
RaTwLIMttf/fm3OwYU+RHGnLBzLmWe7V74Y5xCMtdQuGvyY3C+5Ha+Q/OMmddFOU3VYMCyep3HLT
G8w5vbaI7zrwevf2A9k51PqCUwyaDE2TvD99t9C4JLNPQ2yowRAa/yLD0IOYq9aAGC+bItDBgOUz
9vCrLw3pzdrPhqAisSInDLu9qgU84oO5+92nA8td6y54qTzBhBKHoFseTk9GIM13plNnOYswdd6Z
s606dt9l6rhLAFjI2HXWsNPK11ZUlndYIVLCBXhpLN8EafPmgIcVWNJDUrAwVxEbltkAm3UxOPSr
6utZG8WkcZeF5LnYeqRNJiUf/qtL1us1hr7KF0OGM1SNiC3rCqkbwV57Jv+yZwThZ5r9pBe9PMYf
nL+fOkHv8AMg0STNDQlTA7cO6dnr2rbSnixRDIguQSC7QkM9fB7DdKUwRttQgeahqrm+ADYoA/yl
DEsJ4zcBcguPhXJz/mHt+ICJc+t4GmZaEizREo3jKB1l6ky71tXFo0thTidbjG4mpeDMDEcrXT5Y
LJhxpRWVm+PsDkhChCp1MXi5aIKEHAMlwRjnyAjgG1cV812PBQrLD210IkV9WMevsoAq+D+pAD3G
TNuF/WvtpQi7tfzj4KmrB4dKV1fleSqos0w0pQkr4QCF79Fv33uSMEMreF8mfxMFI4sV1dmdj6qO
/UXWVUFbIGrbhBqkG2wCMLXMAo5Qk/tVnfpMf1vyyLAVCor7+FZkcV6wmPvbzzACtmvO5xzdU5oy
HqFLHNFtNwn1gmocXxHTywscyQoyr8zI+uPzIXXD9gJZIfBXav2C0PdF7qNw4SE+kt9PeGrM6/zL
dp3h0KFveS3IEk1D01Uo9O4quoZROev4waHDpPIB7uez5TfXCc0nBVB24btXk/cggsX9VWmYDCzn
s96qVKid9Z1A7++xmkIlM8XiLUT9USVTG2X2jT8ZjntndWKI+r7vnSKq8wA/vieaF8L25zmDFRNw
64ueBpWkVQ8JsFT61mUhvSBPeo2REeKHD9Y1flA+IzHXkoNmmgyeF0dJuCBLUiYv3S38feE7M167
KgAZW5q6q9chb4U6Nnbji3wMVx/wMRE9rdiC4aCyzHCO8s3DeQjRuF8tcIh3vKRMtsNPsDo6Kd5y
O+eVAY5Ehr8StSGGYTIaF4A/UI933wMQeU4Dc8fQguOY73caFWRtiTt2HU0Lt2ozrZ4hVrdwTq3K
B8a1ZQ9Tj9ap5KI3uAQ7G6kfGdyo+L//A2OrKzZzkJf1L40QpVOl5LR5LZ+gkMlwnPQqDZ5s79/Y
xzntcuWExULwUK2gkWpPxvC9OYMFGXGZMn7MElV3kRhdXOM8GcpcrTbWUwqfClV08cxSPmU5u0Cx
mJ6r7KDa8hqwM/ByABLW7YpZ9LKcuwholkLO4DdL8FiS+pEff6iPppuQjwKzcQJep0sH7OsJ96Az
6NN44i2FniKoN4yBhxelca88pENbL3jasGGQcHAjipom1ywOWiEYqBOYbmsdlwAfBI6aRCnlsE4E
Pna7vJJbXT2rwFIodvMzazqRF/YES6bK8/JfOJaJ3u1YAdrZQA32hjeawRFyUGt5TON5tYClX36A
FSkOWSWr0tFmwRGZ874L8WR22nmxFfuKbiUV+9KpMrYm9JglXFGjE1uMIUxlTOw2P2/qFVazGLQv
5mQFVG+F6KMXjmzxbvRKcSpML3L7csT93hIwET7zOXCX9lDrum8USaNm3mE3xTE2Jy7yO9rxB7Ji
Gk9Es5L4dViSXLxGPMbsPuKYUsUW2z41gKgi/aU12ZMwiYk3Lti050U0VLEX+WT8K8K1xH3fHIof
wXPgRYeNG0KdTFfIKHjRS9mIJXHdl5Z/Kl70Z2lyKYygsuHsCHA5gIdieLg/NjZ2nmwa9sTM/qFy
FTqLr2otI5fVJiTon/lqhjhgfNPRy3zdXyVNdliDyAMUnZLWlGfj1ffKE01gLVJtezB50HjA2aGe
XAYCJRd+3tdYw4Dfs4feimJzAznAZax4ArEcKQtRDcj6iCajXvv49fhmW5c5im0lTfUDoSCHdZgZ
GwXj5QU9PseFpab89SRZAO9/DUmkkS/CSGbppARwSWM3M8GZPhBZ2mxpRi6q1kWX9u5Sd02WipHh
rUtzZuEIy6ELZ0Z+PhmvELeRUzT1rVOIsK3qIy9NhsN+0aQ38gsNvAV1pexdMSuTRvMNanWbZ3FR
78xgaDS+UgIeNSqJhUsQvf8oazWy+E49TNMvXJAUzyCrcLSnkJkOUmN36pX04hiYBsZkECjoLZ8l
JCGOYxl4W/9N1sWxla3to4sIvxJGnxLk/uI/iUFRC8fuiaN6ag1CnwO7JT9FABcFNXFyxgFQcYDi
5I7qcbvxr57nuAVhlrva+l/TOwdTIfEq8q4fDl+Np+MPuqFOsXVD+Mx423+mHd7CPnxDMGDs3jT/
yKc/eFJR+rFOnblp5UL/xmb2ZwT5OWUhPZK5bHJDu+ht9+YcU45wZNIayoJukukl04UqZ4vSGtxj
zSzcYxcEIvCHNLKm+CimGIPuuG/ywJBdLhW7k6CcXvm9UeJkE+7a9oFgI/jQk8uikc/5O3BtQiTU
F5zWSDVKGiHMYwEDrDNUBTWKYbKjsXqih2M1aeko5RmWoqaEJQYGxbJjHL1AcJJNRk+eDj+64gis
UQCGZZucFUMQ7JZD9muqnAkL1JigdhLowSrK9KeLAzzIB01k8mLHnfL1FAHmb8Hdnkv05UdVoN6M
gSTKBcaWcS11l+WrizKsysEFsXq67WOhvMZ8fVY9g6SEuaj2gr/CAFv1WwhpECutJUVj8YoL5xl5
7MGFUS8xez3SgFfOpag8Oh5ytLL4VaFVTstzeXW+T3rtOs0XIDUmzYomG8aUmseKH2LZJbzZBy0D
hAEQb07w4EPBWSIKlI3C33wim7oZoKHWnkTri9LkpbZELi83qh+l+LIifDzJ8SPF2GWyvwB7H7xK
b3DI2c2gvfBkMOLBI+e0rKB3xvddleWB8TSOvuQX3YpX5ql9WyVP08OKTfvFUVaSVYNV3qAUaR3X
8Tnm+dnEbhCGAeJj80uBVLXZLvmTE1+z9LpAUaZ4kg/+l14ve7eRjAjTCWsu2DTzeT8Bms5Cb5z0
ItgLHuMFfk2Iow3e3KheUsRt+X/pgxgCpPFXLf/OzPbCPaeSG2zc7HzTRflMvHZQE4OItkN1hqzJ
97EgkfIy1/FiDwXf/+WkBRIkLAGMBI5rcJomqqcumQB6/j4JAzFCF4Y2k0TejhquRLSZqt+bXTr1
c+VBQ6Rf4hEwl0oZsX72MG+l59iRQohNXDpjH6GIxfe+OetX7+mA0OQMlsWa14RuF0Rm8+3SnvbC
yCQkXLwFUnfWAAtwDJpwEELiJXyAkjd0GyYkoiJxr5R+o5/PsWH7rNbSDOIKYoQF8kJBGaGddeS6
+amoELiVQ6s0ZuRYiInHAQlgUwJv2GTFvXLGiJf6gNEDCqDJEUOxZkTLNCWpl5AnvsWsKgCzPNDa
Dld/Dmg/UI3kbkelh5Yie1YGlmnMeJp0gR9yETMkLb8iVXUNMtmCjLYFkWQ46HwpaFc1MwQuFhOJ
t9HtjHOIgnRrN/ohIRiDBMcnT8iuc9/bgGmM3Y2fvSJDzYus1OAZ/I/ubTdLgB6wjW1rjfwhc/p6
n9cUoObwPsgYmS1teNpLgUBt5TTnIV6jHOSAiN0+tmCzIDGMRPrIMqUMuaWMAYA3kXhFy+xrRZ91
nFPpqalTFvGtBzjfTOJLlR3QO7Lc6IDZKJN8VdAM9jS5cy5jJ3+It1meEOIaI0TChDfpIU03Sl90
Qgjrl6fPsKRLUmSiiIwgf+gWVTzRuzTnXrfyA5nte7Z8xo5PP5s/bdTJMqDxFx/tmflS0kl3ngzL
OG9VXQGoBHQN6TrtyK5C7/Wpn0obhLX1yO9UzVzzislhkL+Ewo2UBXG16KwVhLsiCsF1v8lKQp+N
70jizKJ3DWZFoECBUALpGWD889QC0EpmsbE9iaH7MIftpNjkTKFK3EYwhvH9mWydwhPeBGCyAD86
kUGILkkA1L7JiccU5yS9z4VtYMnFSg3MbkbU8N8QlTqOc5l+I0qT1DSo8QJu85BXuxRFA7WUhNzT
LJO8QYJcAH+0KvblyOYFDCLXH0OXfCuG4HcptTNdKjXEZhV6BHdudTwIJqavBStU2tT/xtnvUdFZ
Nun7JbYJ8rXAwzLrGg4pvmOg1fTWplUxoTefqfYv9i6XpUZvn+jbrDbpMZAetVE6+uoyFW/He2S4
EgVwW0Tqu7zA6Xy9/prINdBL+K/HntE50HAC3lXGKwHRqNIFXwRH9BWvHLUqmmo8utW0yhJihv3d
SxsHcoZzs/k7y67/iBEAfycw5b7BXtp5/R5QRW88egKpdw1k0jVB21giNS+/vtTkDTaeg12n0bGe
+9SRm+e3SZQFaaV08aJytzc93Scs5VettkFChNXkOLMN+Im8K1rzoeN57K7GDqJ9aKTof56qWr0A
lgR3ig0CxrYlBI0laBQDnYfDFMiDK8xjjSKI3iBZ6BsWCCsiMwOBeX4TQq/FTsr8DWkhiU98b8OQ
MHjL0678R+yIp4yOC5qePTj/0peIvDwp4sXOWy/muzZxyMTjxnmK2McGJ63Tm04wK2Os+rQPJxd5
xnxHIwp/2StMixuBH132NcJAZOQUKK70o/hGGfLHEntCKCP0LAgWZfCe6aBPtxU/rbug1El2FTho
CLER/Plc5tz8Tj/p2FsyK5cnLeOT82WGqK1Ysg+VuCjCXtt6zFBNYgUTeRayiiYXqR4LiuryUbzd
FRcIMPgPjRlG0pt6a3JVuTrVYU31NtyOb+I2ylZZMjSCcD15AwE1fHMtbXzk9OyPjyGdU1k9inLb
Ej9Nph6U/ZNsuLsYpD+8AMdzY3IVCT+IbvTSriNPewCsphWXP49KQVO+zxio/3nUfffpiyC0s9/P
d6D3jWKy2BGPirdz+ZjKTsoujt0lFlLbxeMTDVHuRWfOvGXcsSwKiVBVD6f8EfkSDDsJgl2nOEIC
n47XWWb6xfSAciytH/IARZbqDYbkYQFw/OM357DOynBVp9ZumO7tDsPdMq4TrwvXHvgpsOMscDMx
AB+NHpOqLHWGjCzJ5VTDGjuxytPo0PaivubdK34bibXYWRHLlBXPhxowij5y6955iXktFeYqhufR
9Ga+t4QY5YYwgvgYYTe4XE44AEHs8q/MfSP4Lrrmrf32Gm3BRg49wTLZRHQW7Goq+ogrMk8Te5wc
9IKNxewZvi156rDUlLr7LkGzlmMoQFMNXiqzYXdomZI95ELXM50NPCL4m6WEEI0mG41jyGdoQcul
SDxXeVnxoPMZw4S21Nq4ASlhnra1jCWX1KtZqWfnsRtiUaGJNSwGXfu+BG7AIZDETUVIsrGD+nQn
qZvYm4FEiMYSq4uHJBSyIWRD1OWc4Vh6K4BORsubCGWr2JKxFAyets2KqJ1OrF+EktX2Z2d58Stn
upFHZJ+3TFy8XSalWsxHi9RIjTpEM67w1bRX7Oc6GJct9ITik+Kl0afdYwWIRLHXeFECCZ/4KyT8
4NdY1NXf717eo6i87i3lV0Wc3Z3WCNyNGz96o+CQBPby+/ILmVJEN3xdfRzs5FRGDKE71AOGjGNs
hlcYAc8nm0y48ILedoe8Oj428yO7Dz9QrXgE6OsULgwsB8UeAVLLIzjTDNFuklqQK7lqV3Tu2+So
jxxZG9A/0ihAnGUzuhqBCgb8kqj7iwE7R0wz0yraf6gqnY1Eyp5FcD5kBFsaaSaMADukTuBEGT2S
XltLMW4FniGHuGlq6k1wydW+rUs78tjjbg/KSlOJ3nynW2dB1ILKRZ91Z73f19n9nTBGuMgnj/QD
jgPs4YaW+xU0XNCwLUaVNHb62IqE0tb96nwWJI0fq0GKBna1wfiQiA6l7EkGC3axQYMsuTRVwj5y
uI8vW6UfaOmccps+TzhSLdCGEbwDhcIx8pxVHgbRwIdEPNIUzQhaBGcXzMFKFJZMGarBo34qv+e4
FglNWXQmftlProLdjxBx7kSE9b2dCPXnDtwJj4b/uUwbrmzHBSapiy5z0JdeCFPADJs5y6T30Mpg
/eTWU2s/4d3Kzs01JYSz7/NeyMZJmjIQ+Yg1gh1ujlgnRLysE8Y1uzzZIdGzOiW/6kcfsFItn3+3
foeWb/qYzce/3gonzwFv+evU0LgjcQbqNWJUI+c0qy1P8tGMu6R7btJBBnBtENawc0+RLYkpzu15
NyPHCLGDSZC+3NSMD1T5I4v9D5U75cJgSKmV3wcQzwClatf5rBU6Tibjmu+r4W6mLk/O0zd7ozqg
lQQ+qbiS6dbCGGxJzpF8eVF571wRuwJ+cGcOCxJ9b4F8HBnjyIwpLR1maunsvkP5+2HpIZSgPfhp
a+o3olc2LZRduL/pA6AuHDGj4bDA53N3E0l/E524brOjsAfZEaRrhsltlEST3FbXdS8d/ND+tlDU
2PL3kelMmVS1Ex5JVCJROQVXGQE4SuRJ/sTjaiwxjtW757ScxjTqpXPK5pf4j6wS0t7MFSfmUHh1
1CijRHLYAivBIXIPEdoCJlkEpAk4GEDF5lggV4XXiB1cUcn7HbqmoRsFcoJWIoqXPDNsQCeAePrA
OPAG0iM4PhCgYNfLHt7/BZMvjNiuvhW6e3uM8CN/z4XWA+PNsF81hG6FyEnss8nngWyvXT5Di9kP
JUCW9nJ/P6Wkb4ayeMlu8blXkVh4a7gHfaCSLaUtKhsWMMnyGZBAr11eV9weAuMaI/b0tqq0YX+m
g3lPfXEXV/vA10EJdTOKlo1kmSUJtqQCs6RGHNS5nsCX4hHIVXhnijxsywegT2dSupHv5pQiiRxc
qEJguruKpdsbf0M5Vw4PkK+bIKwOTZRzvBTzNndJZCwOk7qlNsZQtv/6Pwxhp57eZeIuHE4oWMzt
X1C5m1lVXneGPn8mwu4x6jAxNGEYAHPTLK4bQLhgEzKFHo0Do3Bs1+OgBFD0JWsUptPJeflD4Sak
kExdcdQVRW0F4mrFmsOI0+wpOb+l7B/U0eU58w8beZtsZAupLooI3lxydtEEzLjyZxtTBDGI9YpE
XcdrHBzaWkghiscqdnPXWvRD2h6dGtCjAxnuoPH4HOfe/3BewUwMBBQyArcvYEqYNBrzRs7SsxYn
ekhQ9uDiV9kO0BU6mBYIjWigtxoV31WPayOz0XqxMsdPqUsIOSBXTInelazRJQV/AJ7wU20ROiT0
PR5MvV5bZLgPQOnENK0gqNM6MG9xSnYQULMG2iFPxY/sdv26RCM1/0zjnr1JBVznHYGpVo76iDPI
8OYNDpdW0N8aBEUW2g5QJykllTmQLaaN+yYhJl+rUr1GgSgC779rtH+ErG5A0/swo7hMiY6HfYPf
sPl/ewi4HlrIE0Hk3/mSztVeKEDCcjnwp7/WQXMl3XLefHBljRAOllBKJSqmPB/eABzkovoMawsS
p+f5Z6+BB6M1cB2I7s0jKF8ppJzL+s8jtALc6RGdO0yCq9MZtjBJgGSG4m47DG3hG6pIbGfS8oPm
accDXhIgWCAjacfiop3o3CiLBPEVg8gX50iEcaJL6feThLeyx56n3g2Ow7+VRbSNw+0VcWW4mDe1
mP7aOqH4SNkZeC5vYkV3YYUB7SiioxARItY+67F5096cma2g8XLllZzszHuqBxLADghtD5AdvCuO
9flPkGLZkhB07QzYF1hKdVZhy20Gg2xNoPFfFtq5mZPUBFyZsjHUQqUbPKcNt/fHLWUidi7vunGV
uh1mqgRRzNSsFGY31hRVDx92gWzVWYntwBbOzCj0osdezE//4llJ1tK3omTN3zh9bCJsLZ1R05PN
XfhN7Nb10Qvdh7oqdDanpgVN3yZXef/YnOBrgZcWV0XWpFWtEAKfa6EegpCb7IcALr1Ruu8T7ETA
gyh+qwLRG8MclqdYzerycFbLH4UWdzv26Rnpmdu8Z7E6uF5b5NByAGL6YD/vc56XEn2rru6wAJDz
ulCfoAAZ07Q4TsntYoCBNiU6bTq6YCV1cKIxyY48lBcInDvVb5yIzUuKDURJBmEBibJnq2Vmx5jx
D30zLQDz47wA0GlFKnQqczhAqKM+dfrcsIaJcujKBVSCnnXEug86ja7YZFAgGmBc1ThRd5Qg+0bE
axVJjuLoa6Z57dG82qfd37xWCqzuAi5uwAPqRhMNFqO/6cLvoRf+2Bo0d1iYjvgKrD4wAv5Fif+o
Yjs8cg5nZRFoOlYWuDOec7Eo7SlelT7q6uanAesgyKcRGf0cYZvEg6hGcqFR809s31VNNCEFLRWz
5SaGVXDndyFHupDp6miJuGf7mPzLika44G1edzUcFnCy4XxGsaA3tGYLrk5KpRk3mv44zK1g9d7V
IBQ+snde8dlYoLCQsbcPWJ/bX0WLN0fNdDSlJ1cb60YR2yYNPUtCGd5XBvbc/FqmWkYS4tPA/Fky
VLHo4+cDcrSaX3QFWSWMm0SIurzTG2t8+RhgPB921ddQ43AvbndW0I39SYDxACStEUxQlMGJHvks
uSrOOHIwS1Fma8cIgNNhmmfYs4dHioHrRxLDcJUnqAtlqjDgYrxxq3pAI+GXlcZ6krWdtMKTHZap
2BHbfka0+5/FkNxqJcBhUAFgxovbspqNPBVnBoNRL8i7HCBJvjRHa2F304ceA3urETFLPZ6X1WS2
U53UdeHO5Ih8ZM8NZqvvlDdhphXAMgYB0wQ+1PoHVqs870Qqozh9aScZ8fyzxrpoM1wUyYYAXCpu
/6xEW9NbepTD15Ka1yNT1ubDc1PEtKiQtdDTs3tMmblDYvkmt0+KVYfDE/RAQQxkotKbCxxEPpNx
YZJ1O10V3TI3E01U74uYMo6W0ojIhSWHvTKm4mbLy+HA/v+xBl5N4HSHatK0B2rNCvY9vQpP+Ozg
XdRTTnyJkDQ/vyJLaTy+H+9jN1B0JeoGp5+7wt0R0P27OPfgoUwXjLgYqEJjKHLApg5jfwJ5D+9G
rHxpked3cx2JKIixHKsEwNWHSSQsyzRL5jSXayqraktMPSradbd80pwsC9qHk4Psv920XsbnUBqg
4v6JNZ7pCcb6SS0q9N+JbxZA+J3UjEeQh8JBZ+p26FM/ZbLNQY4ZeFc1rrakv6Bvqw/kZmWv4KaE
OVsJMMeKPZliV+4T7XBQsIeSjMOtzenHjSKS5pNy4dJYMWihMam3uvMhU606Lp93CXY0ZlN6EZ5a
64WNccHZZSoTjcGMTECzY3z8n3M6z1bhSBovCYzeZ1ptW45V+xaeX+tfYbo8w+S+dKDARIjjhgei
FHSARVmBiHr94WCNgaT1eU80qucMWPcuuL89/aV2L5Wlan7JizF0jlvZBnZVsdtdySPgCLP9bEYo
DeGksQuSdSefOUbJoQ4/cUnlXxDLXWeLF44S5it5DUOQvinMkt86BgjFM8HV+fT3c3/OEvMq1ysK
FkMap3VaM1H/Y5eGyb5dL5l+EpmNrPNQmI5ZgwW5ISXL8mvlOwJxLOVS3JVzOKjj1UjI1PqUj9/w
I1ymvCyn9e2K7NEPlWlN+5WXz7LwtAB/eWOXE27Zh2Jk6PoqPX8lFYcbglGH9wAr8oNFPiNdMsrY
avWRYbLGwzvoQCAHS/AGLheSUHP15cOIej+o8xWvFtWFgr/RIvfKfbEZFoIoeKMLoswnlsUu+Vvm
SJDqqn2Ej9+GJafSF8xJ5XlYlTp8Qf1QDXLc6nNi+yBsh6sC89on0ulGgwq2jB6zA/wCFA5SjILT
fBATQS2tWCVNyI2/YcZlqjQ8/g9LclvWAEL4EVCicxRychP49Y1Vddbvj02Fl2+5fLOHUoXWW10w
Pcc6cIE9A1VQNCjXYEXtFKTKmgsFS33qdv1AURHGANIwKCVJ9H6/np4PGZEyyIxRCv/Xge+kOotR
Dgaj1aRIXze/qv/hdPmcWmY/LCb83N9zZv0UKHmQIWPUeyc2OLx7MVOOL7x9grf/WVr2K4ORFElF
jxOqGAP4k2J36Ow0ZlFZldBiXjvgCek72RX4DX2VFvnOMLQQ8YTbnq2p6+4etnVM482K4eYGP5P9
blW3nOnE8uSMu+NR1t/iKRCMGjLNdeweuB+5CqrfZxrbngkNB1B+O49oOQx0do6qCkHfbjEjLiSX
U99vxJm2vU6KXLfoRO3C6fdFPfTjYZia4xMnCQhHMZRCGXxxwqBJLRR9mMZMFb0pGsUjKAzBJb0u
+00E5morsE66b0m69sMvRVAx4VzraYpWK+Cngm5a+HtM5HTt8CXy0400FWelxloIODe0YJ0s+I4A
X7//YPWABqSwb0euf0A0Ssf26h2OuKyMcdMn3mimiFTkMhYURPRUaUqbbliVx0Tj1E5pbyWffm7A
ILxZ1RMUagMA3e/paO/FYkDrzha3bRJ4aT05cCKsVl7c0WnalXixnGASh0QzmDrSrVEqxG61ABen
Xsa1PAUO31TeSZ7nqJ55UoZZA1SSViUf898Ag3PiKmL3LtGLoQN7LKOg+6xA7X4fOR3jJ9BPVODN
MVNS4PKxWWxqLYmx5KgrBYK6Rxdj3zzwqfQCyzIXQ31AN+GbjxnTmA+/cGA07UGG4RVIPelSlis6
4A/hN+Hy/zurCb50McSY0vgSXu+aF91CD86K8mNtsUpyDpSVUX3W5V3gZasw4kSluB7gYm2HkHIU
C84qnSmaK5eeZwLfrXkjZBGFPmPcCLBK0eHlH1LzRjKzMq1FUqWEqvWhtt+PLkI/vooMZuhq66PY
OiZbwbIDFNH5StZgLfOJ8aS7e/cqE0wAm2XdYotdhoiejyQTmPMM1aUvdZfoTznIJtyoA82VeCxJ
zTaZvZLbE1X4GuoWKPsRTiNIVNeqsfJnVOO6SjL3ctiJdiHWuM3aZ43xR1//4H31e6y9WvOXtZJo
XzZjE3BRdBXjPw4Ct9rBOgG0jdQHaJy210AbSgg3bTF3tf0nO2vxaHLa4d4FakSKyYZ27LnkimY/
hs1szmv84eWr4/DJNiWNsetKzbFQwublU8rGEEONtMhyIoIt08fCtPx/59BE3eVRrHXkn40ya1/a
WGYqGZ2jhXeOO36EyiJy6LyS+A/a1SUgvDXwJql+nZak/v4tTTJ4L4VvRo1RmUsnnpeR+2NTc8Cq
qEFlXqJz6vbK11d0DjI/lHV0+VGb+ms/2eNFQ8CjyiezaoySm/rVGEUnqbXv+F8CjS8gJItSZUkx
jqBeuA/RAweHEav7qOlAPUV34jQaOis8ILpFzIRRl/6OxFMYRKwdaJuUK+f1fCHwvgyBa8m8WiSn
OEIOiomPYp9wODIs651SJT9iasYuDnUJ7dsUljekptif/+5/dO3i5DoCVaWOcT+LArB66hVBHVZ0
WERXi/Yqz9LSyS/jBeur0uhqpef06Yv1LnaagTS9y0bbvtbDUETjAkaAsLJTkl+ILqMbS0Pu9/A8
RiGWAlQJ/JTM9P8QAyTBfhjvJn+wvWsN0T8OcP43fTk/NMZSFOG9baovAiQRRnnKe2fOTl6bpFpA
tNvChkMBkAGNMTVfsyK8CboDXg6xqtp1UwHRgVAjmelHghp4Byf4X153b6YE9JS5P/6OwdhlY20C
GcRQdma1e/7ssmB1CL+Gj/RYFofng0F/ssbGuNgn+qsR++mq4wsFf5z+yUqmdRh1keSy6AdI/B4b
iX0HdqTRl+viFNOTZQ4FN0J9IaRtfTVn/r7OfVaLKmxwtjJ+OJAzv7UEgOopvrcDQws/GnAb0OnJ
BjphnEYC/Z7HJexHLhx35De/1NxE8qfgz46SMF/2oNy7OgUHOZD8zKI9YVyhMXBYbwPZvSO5AhCk
UP6aqNnHJXRthng5ywaOdmeQpcPnD2rYhCP/XHpJfUc4xXxjMO+vq4520+1KtqUBqtHGl10sa7ZC
hxSi3F9lItOS1DZUoozz9FFmUSOjSeBYp+qblLzfsryEMlmrL3sz9kwiyM/MfAM1FJZhNBAD0cGZ
dcDz1EHqqGhRzb3e2E2NwPnTesTCZtc5zI+oaknsPl3BBAkd8a29HpkSyZxK+Qu40NfoLJSWm+ap
j9vIkOz9H4L1DOA/GPGmp5ILqF2YZo/F6Fezsh4t/hbx5wCzD7htrAkOjROzexI69CO+07wNB7hp
XzdVoU86NgbK8RVdZocwF6BzqNDEiFEnMiAaSPEC+puS8WRSAjE/IpzBWDe1IvTM8/X5CXPp7Zo3
nr111M9/OIi8LNGYnppT5qhWXSZZboh1UIHE7/TY/0gH8BIjndhSx502Sd34tpXbNcr9z2QFCacY
Tu++iHMYFw9airsUWxo+fRjZ/Euz/CN3rOYSaNbsXKIMorVZbvwnCEbvQIPw45b7h00WfBII1FB2
60PSp1FLnvXCII/mZEDsKvkqRPJZdPD+lfP4xSXHsfQodtxE43UjSTBRXpMRqnxoKw+98u7V+O8i
lnZ/Yp650FGMDvDigHeFJsYjJlAMyA5QDuzYsZw9jVcgDuufK4BRSWYWdxgBfgSi8JezXNCdv+72
4nE++Cl2Jryaeh2G0cZW7MRkIJ/oye4piPrPbWmNccc7AjDp7CkMr5ghDrP3b0QQMu5sJFgARy8f
gOZkqS4xQQUTfx8wcitLXoGLtsJ+W6EAA+yycVXyWdjw8IFLJrEBTYUwU4XpC7rg5O1vOIZM2Vu+
2CQx1DSXAmZgnRuxloZjUvbk0xaa3Ad1jn9QO/qKNlwztVrHOtKiowPIHjlds3nEu+odM9FOETmx
icweAwouhIIe+x2rOqLOSJ2Uv242YUZAJ+uObXaDBDLFsJuXU7RzIBXJPdD2et7bSsEYOFLzGTkF
Ze0qHeGfvKok0Hh6qO4E5GR+gV6w53Yj4/b3Hmy9cn7SacgZoWgiH0m1AuC5LlpKrySMuiNvqxKt
ToAtex6jMLBIAkxkRkNYm3ZfR+sopHIhmxnWoG2kYXv8KVy1uWxXE3nMDPZMXtJdyunFNqyHrgX9
eLAGeeGBxIFmaklbxUvUfPIzRneKxrIgMUzBZrnMldR1slpZTBD+zbzkbYS3sNnDTVP70v3cnGdc
mYedYxFnWsyAeR9V8ts25NUffN+ZKqLU6M+w8JB74RYIJ9vZ6gG+Vxe2TO2wXefNXtMY4HWQh4n4
w+dytRL82yB2jC8YnWLjoRSzIok7kR9r37TZcUxLoHu2+FHRkBqAzftTf2zoORL45mMXcvGeO9Gb
R+mNctisH83okPQ1eukAf9h2We4UWC/b1wraPqZ7b+3jmbmCjRHheg2GwSI7+pEl3nWMAqiZ/ShJ
PKEMz5UdhWF1cj6eGT6OdsotHYF/5GIFFVO/xhzvm2epCeKyqj9D/dYWziXqR2pG4oOQLUA21FEt
ks2+1xJgQZt18DzM6bsbIN5dvBi9nth5tUSQXS0S1VHgN+x0qBLKpsuWaA2ok1HB6519mnspVIN8
7jW+IuXAVlY5Ww4WgRyWPhT2e8+8XTtn0USD0MweSNQ0dy0SrGAupzeXbunE2c1T6GgVB9THSLWg
uySfZTYiP+VtXYnmrTiNNhKe6adBxRFadileqns61T7SVckaeo1jQkkqCO0U4zT7q/8H5U7sJTmr
FTkX0usAz0cPJuu/mL2vlPBfbBZ2Pw2IuaHM/5MgrhQNy5Wv7Cfbao5pbJFl4Wjm90hh44PysKjT
80HNVL1PHm+OKyJAL840nHaNFUW0QXMi/Z8lxWII3mtu7YWz9XTFmRsf5bedJxg4Pepew0Ot4KlH
Sg7wJx7obpDa0W0A3qJ6BoI8JLGPhPfWs+uZjmT3w0dTAmGVUzC9DGPRQj1uswTcx0isLk4xhTXe
BX6YQyGK+aS7yXo00DK19kQrp713KePOErERISdbAVyh95uS46TE0jq1dGXqiWBQFsW8l2O6z2Ml
77UPombBK8hXGMGPIRJeuFUHzvCLuJKI+PiTZvvoKSINSt/JH635cm2NFYoq6DoSyhM938tTTYK5
t7CuO9br46JYRUIbv4d4JGh9i5iKbpwc8kbwHYL9/nTd/Jr0dRpoEv5IjBoknMnIObkhTxkTPUJc
p3e3w+HHMToeNAMSstzbYMey2lEjxmtoRQQZp6aA2GXMXUfnerDZ84fv6fBwN5ALw7h3rVM74IJ9
87CptLdUixX0LrQaO2KqV1mhATBVaDPPLnxf7Gec6lcNbmr0wJ2800DpSRScLD7UK3bJYTnJ6NVZ
ymrRfXSzs519GQNenFMlpkMm8XOrw4ea57OieKC0hKNVv4aoefWJn0tU5qUiOupVM1WiHwpCW7Qg
n8l8Q0IS/w2Dydlai55ofM+7qxVw352g35/mKeIFcvsx30APCB75chA7PPHrdUF3OM4cTl36DCRS
bJkWhwXSBebIM1cRrD4I50IosJGZEtcP90YxcFO5F6anckmzoBla9C8i8uocJJVLFiQ4zsVS/6OM
3cZkNM6TBnjJg0SsEmnjIOS1yn6NRQkjRjqmGoO3lmQBtZk+0T8gy11yzvHCi21UYQg/G0rJLkUB
YVb1rmAU0QTeyy/3GiKvoJ/Dh+5GJ97M4GbnKgx6REEvHOgOTomKw3DTCu482Ol2aN5447h+kWEH
ryG7dlgvSG8jmO8+x5lVY7Gu6QTyyFiFHphWm26Ho4G3Ej5DTTgho3XIavW+1ZSiLECzOPwIInT2
Jo8UbuW+MwEqBRzACrwC99jCPs5GPkqAVlkflR8NwBibu9H6mDd1Mm2KPCcFB9rjQIO4NTDSmcQQ
06vvV/UP41PDJDi+ythOzIGBzN6BmUEDTLjjjPSTZbkNMYpmqNUD548hXW4s1w19azwf2ms5QoUu
ej7N8CE2xR4QqZv9k1NUuKZSAEcGhqq5g5Wpu0dZUoOM/OAqdqcEJ5jkl7pY3xRTjjUm1AD2fxqB
8HeW+WAXI//67gPBxwz1V0poVaRIE8o9qzO8F5xuMEZob/C6+Cac1nmXy7+XzUsclTTqXgJXcJy5
6PNq9TYUWjSQNv+m4JnjBVp91O0T5LXDNprkR7Fe1LsbJv0tz+OPSGdC1hvych5f7+7d2Hw7CJq5
QPNI09EWUf2vJD6+Q/tTSa7OXrSCiIgmuacojtsGH0uwSQWEJa8/i78A15CFx3cOpVAS+wIRmGwh
qpkjAZBJk6/taIxhXOV1GiQjVVmhLZOjlzA3whYIC5MGQDEBrMX6s01NZsr9MDPtgWjKlVveGw9g
Xxt0yY2aV7Kztd9gbhCyCa2cpXA4+Bo5J6GGcJLHuBOeSa3iSxL/l7Vu4ZtJAyKC8thxzwxbet/F
qAL39NRtgqubBRRR5yhY8axuF+9K0W/iNfNEiFiL7cga0dJWMSab+OgDTwMCfnk179Ssa2WZlUSv
5MwLPvcaNR4THvvbESPxceydFMmfpGlAm+pC5szjiVMo0Bw+8nJQ5r8B6fjeb6+cMUtbnZr+BeS3
Ao2XQjDBORjWAGDuITI8sftyrcf7zfT9nGQAjptENF3QnITMIsNZwKgTbut5+CBmltOwZ7GO409+
sDLlFdfPdXxl2e/qA4bimSvsFUYT3d+qFircvp2aebgoR6jKul1TU8iOW74e2X+SAgLO7eraqMMM
4JMZ8q6Y2u0ADZAxMwntpdSWCBHkKl3S2AfHFqwO2J/ui9IXO0AUgjGNcECNyH93vd+38ROVtBKX
pv0JyAvZ+Qs02EWTlOxOHdR8qfZaZhu01PDb5+1yVpHweD2EK2pvZ0R0/osEsAG1N3UYbTvj9CVr
TFIUjd2FwRx+rCLlEMyvnljo8sqqRfG92m1PgDoOwjEmXq1X0BSq8ZkG5D4YkLLToRL7tzBPGOgS
7b+j7VwtmlRFKCxciDV1wi6jiCyEoT6gYxHsAj38oH5wsLbtr6bQcRX+AJKQMggOr6G9PW5cqJdg
tw8DxpIiLmvoY87hi436i7+S5yzIuDC0FhLIVqf36REDV9W8CikTX6ORRNnr1P/tJWZDTPvV7Phc
dYvy24dGQo6b3SNqF5mOEtRo1AHWBs7LLbXr95rGLoxHD9QAhDkWGB2VK3IUFZDi3kDL2m7b2Nue
tREWt9IaRUIqU8djO1FXtoIIm6tnsoQdj4jiepUgbbp5Nu037Rh91Lw9gUs1kJFw8vKxYWp9NsPj
j+sYL7bBUANuZghuLFm/Zo34zjhClQd7FfOtfxh81dagonlBytauDtRyk1wK5hhaGoL0otFyV9P8
uHp14VWUQ6hQuwgl5pE96JBIaa7KRJg+hZq/6nSHH9ozK3F8cQy8YfblEhErtCXX1XSCbznWT39N
w7P8AlluB1+cYgVvAdeor6FCCDOf6AbFtiL6iVOjQRJl4Uv1AzLwDKoVAV0EPGfdYI7yl9rb7YV2
DIs9XcVkvZkFwCv82Y1eKL5M+IgcqZXE/6qugVqHO21nL5lQTvvuz//MDp7KyXPyqNmD+UDVHnJ7
iq5bppFzCQh/GX/fojo+Ham6Y1sUbdo+ClIoLD3l9x8LdR7ngyMq/UXjCkvGqU1C/1r4fSpQMI1e
2CdAl2RcmDChtwb1AdmmlSmDNCuhcTXo1D3A0c2qR7KxrjONj6LgZXumSXnp0ut+yFz95Rbl8Vsu
kfOrxuavqwNvJkdfU24T6H7uHNbRvnV5D/wGZFuCWZPxWhOYYBnofy8LPPHdSikXHYhJ+iFXqfp0
bir3K1PU1gv2+cSpebu6VlsmAvG4JThuL9H1oYSeM4zAOh+EWzE6BkQSbgvdQVIZGUsqyFU1D7fQ
p0cE8Ikd6L1OCU4R/ERlh3Q1QURY6jj2Wi7P6GGwQrx0vmzn3X8kX8J1aQNxOTbAX71Hva+FvksZ
jrdo9VAPH/QxrQy/TpatvCNhNeO1fQA60CtB+xRKAfm9iGSpfyqH/nRdaW01M1tCdTWGOaflamZT
YBHNFogksV60v6vzM7u2zqoLBJfrzfvXpvrJwiWUdl63LEksC1Urz2qpBjukNw4/8GRySsBIanwb
+CUevb0mGeCAafqXh7SwKGPsunQl8WruNSbW86kHP8BmtxFHeMvOw31HOu4TZf8tOEjj006TU9BN
FtvKBzSGtkKobgZ5a8dnnv5smkdk9IZ82BGX2dLHrF8Fy+o/E5hj56Uy3GOq/RDjSFhnaRmmprAX
aoDU/qEQzYBEc3MS5gxOm0bIix+Mm5CpgvYq9F6jqa3WeyGhWPK9LKhKd3nW5VvL89UBbTSjD+rd
hzuOa1CocuhKq+ddNjrqGPc9f2sVdvEmHRFqq+tW9LJq9Zz2ll2IIfdiP4gskSPOkjayqGWdpa0M
bRtTk3S2nOVx2CZPhdzHFmuiiKQBaL3ytyxnaMvmy1uRthWkfEblrCjeb35/OXZ/odHIq+AYnYRp
DQ9h/nR/uidlH30OfkEClIaWJlgZRULsjIv/Aa/7YkJlWkv8NsD9m8wN+zm4GaxcqMrFa9TClwCV
h3TNM+2kKrralEups5PIoJ9l0Pv+HZp76BjOvZ1EG1nhp6Q3EW7a7Kkp1MhBZbBE7WE+9tPj+Ouy
1Nkaqf2O3OhgXH6E2lhPeW+K9kaUgqV1ZOmY/Z8V7ylS46l46/s9FRBKU6bCO4sRl6fYmyNGKqgh
a0/PXusPtbtar/4vmMM3EvXvrNNkef+k8wRsOqP5YUJ7HRSksIv3kQJ7RQBB6zXpi00vLGa6tSmw
GrL4a22iZZ7zD3esv5vdPdu1eqMNq8/fX8ezo9SRUt7Yqdz4cTDqVWtd3GeH4VfLsUDt43Wl8a5L
zrsBlX1Jy1HfN3pEtnTVoAOOD4js0iz5O1J7+XmSjR+PiB0QK65UOsbM4/tYWrL/VZ+Kx08f2M3a
XzcSVTyMVMEleVE7QvPjvplxhSiyKZIf2fH3EQ4kAY62jbO0AP4Y8I0C1DgJcB6efUWckR9ACE/M
0fzwF8aeo+As/VTqZGeJp9M8A0CbuIcxPcedPJTEwbSZHLr2roIhu+/Y0vKugK+9fIZZC6TrJrU1
7/D7AmDS+/SrpAxk5xDVfkqWj4BDfz8TlDtId9ZhYdlCUhyp2aG9ToUA+xfMyXFlKf4I1idZTiwc
BxXmH4NchQ3NHJYELKLXaXq7mwB6a00P+dBXy9rNvKV1TcRsWDiG3pWfn0DzaZoYestA+QBR/VwV
xFatswqqwkwD362gQ6bOhemS1xvRqg8UC87zonj4No3SRQeBnjkJzVgvyttfrPcUqnpHMYj33dZy
74J6Eh0dmOJpui1ja2GFd3R1V7gQeTHUmephzh827BbSVJAftXCD7yPC7m0IvE7Lr1BoON7M+wgJ
BJK6efTZ7CKfLlrubUwRRwqsxY5ANqmpz2CfCDXsarfVcU5Dytz1MM/YdGyMWfifQv3fo31mUQIe
q6bqKM0by70qap8kBa1EQNVlLLrghHOv2XxglwTq5g6cAq/a6wSu3OvKinYNgsaXlSZPOTKFHn+g
n1m+O/NqfaVIblnbtoyjCaMYGDc9H6PHCAigDwi410bh4V4xDZp6uz8DJEfKEsFWcc/kDf0ES0aT
Ni2bO/EOPPCjWUTqV1FSE4QxsflK/I4aiWAJHae9//HcQ0Mg0szEJi5SgUhn0FnjEfnHY6/C7C9j
KfR5JjkkCi499FYJ4HRXJPy6vNx/j2+TCXHYuFxuu07RuINuO+EX3ZswV7Do2FjMx2Ekoqo8JOUW
EPaDTXuErnE9QK1QpclBE75w5URHFMSLJ1yyZIb8TgKYZyZ5Xtatp51mpCpiWeFDQiASepfGjZjO
jlrvs236a+Oq8E0s6CnfSlLxHjfjwT2IiU8K32YnynaU7w3GXhpVhpR+o1dxdTkhwjxxcQKQfTin
v7AjKKoakkRrfIIVJLiPeI3cFsFd4P+bDJ2nkRJl/F3xU0hjtUL20lhz5owKAOSrt2hu4zVn6oUy
udikFdlYXt9tWuRa3A3X7hkZIk70VqUfufM+2aIJyhQFGzdGCzD/VlqoS5Vggntdl2Erqn/pg2Qf
irWjWYF4IejQhW+nLdrCJO4SngpulH5wZ2/mWlDjUVTFUZ+3fL/MYdQUbmexivbpYVRFHeV3+SuP
Qk7MfYedUKVNg04Sng+tVnSaoDyyo7/u6PBZU9xHPd07Eq0xCjS/gzIpfXX064Ce8R1YIP52khOB
OKqkauyXia0tqhDfxJId64dmn8rNvw5cE4cz2/MiCP3WuCyRoLPlfEbb0uOg8CopBwjT1ICzLedj
IIYFxIcqTWGmOMDn9V8u2aY8ZCcU9OThE7QVR1loYZsH/xmtiXfanZljLXM6xLa8c2uSIgTDnWAA
rM8PZ0q1iRG9dC2DH4WUvRW2U1DX2gDh/45PvZrm45HX2JIDnnEFHcslkJcdcWZcA7prOQZhUDJ9
mPrD/MC22qAEJLsLwio5jtmnWICRklRBRMSzSdJAhcwnaCLlGtAV3+x5vv7RHg9GqO/PgMuagdUR
apLeTH+xSftPezmptj2/gE4AyUedU7puSS0OSjVsebS+I6SNQeB//QnLo00/ZkdWJ55d2AtYh1Bf
JzrMbrBNciP52V+2lCMTBMqEDLMf8wlUwQ4/tKycKs+Zyz7FdNSDFt9DniugTT+24uUYu4PtLbUU
fpUda71okItb/4PqSHd44fDs/e27NrAQBy/n3s/RXEadHtN5tjLHup9F7faUIZE17LuxUVl4wwtB
/Ja7y1VfzAwE+3Ip/M0l0wPJr0HcLHTQDkUywSL5YBUKTRzOxkWH/6M2D1lPqmumgw8SXPsl5Its
+uTZfskHIVMOQhglCyCLZALp9DjRml38MtqKuoZFTeEj3es2lAS2NtsFAuENFCsz9M/AstSfMSWs
zvkXM+QrIXKRBsD1T/mkHIn7Pnj9nEzlwenUXQXf27XWV81mY9E58r2gvLr6tttacfAl/KpgKxD1
0QyoQz7oWjkAXC+DUGmR1LZRitNF9r2+tsUwbz/KWugSG6VWMiEft20okWJd9plGgnU/9MTIBaaV
fxNdh3soKBKYBlbOmXXOlVgZGy5YRB2xHdahrRmg7px3mBgKLJX4jJB6hvcYJguttuUKZo043ibH
3ZifJzp0RLxQD+DXZtWHJ1xBTK7HPcienLOdN/y16znPDAwLf+DaH0NjdqlqGv8zAc/dyFSTFPEh
KPpcbbCuENbU+vaV4sBOh93dgdf7QvFi9m+4XTziDwoPwB0yW2gJ8lEWZ105f4RgaPe9dcbKsWT/
wufoy1+sr2zritaTOuVmUxZ8iDdXrBKoeNr12nko3F18OeJ0skGGp1Ig/kz295ISDxymxLqjex4v
01pIFgoI7bKjSBilDjpSH0Tha6KcZNt46S01oxd0DtL3Ll2JkhB2dfSkMEn+TYTUc07pl1QL4CKL
6yOrS4Ikz/Av7rM8Hjcx8eiTPKUgMk+REedOCp6LcHnPNQiDX+ymYR8IDMyAjhKgD5Zib0zuzu8s
TKXkk0PldmpjZmX35r9PJiqYscujmPeasT8G9iSLPpTGjIVL4DADg/TcT5ykydCN7O0F8QFIa7Tg
jORuikW/ut28qgSmEpodyDynrkar96ow0fJ6+oB5+XYo5dcQtPuSO4wr/bsZPWehjoE4yhjWJKex
fYRvxzX0+DDYpXEBAexBwY+m0LmwX6ndp8DCxS1n1gfZBLaCyUYj4JtVdqB2Z3xG61V5VHWBxleE
KonmivdGnAPSVfWg1iM4bEE6UVMVWCmTIAquAUW1Qisw9UG9HHKxDv4dd6nsZ2Vap43s9Ekvy8Bt
TllXs+tML6icd66ladfm+mrhUwhmi220uGfdgXT1JfFkyrd+umZNPrWnn5/AxW1sYcMSY3CUXHwJ
jOc5wKHuoiC50sLKpDVeEiElQn3nhbtXZNSIAbcBrDa3QQAlDbmOIqbB8ueCDj12sz3uT6I/9SPq
+WHiLZAOzqzyfT1eK0c/RDS7NnvH/s5Fs3ONrgrTli0T5pvktBpZI8nJZxJpGOKj3bvRI/yTQ6jj
CHlbh1ByDIom1qbht8C7u6/W4ivbQmYtfW+A3OK+0S0V1pLoNhdwPKJ+qNVq+hUgPqa+Rs1TXsx4
eUhaugZmeyyRrtgBrsw4Rr9Rh1UuuEEz7snsJnI3hSkkALCG5twkFyK/mQKx0JQgoZwlE3ZBBrjS
n2Oz+NjrxHik633KCZB+9ujdMJrw7cnCvoH2a7tVgXfJhprt/X+0pTmQ/NhdwHeN3iejOUpgjsE0
HLBEmnJynECmQvIKdbWBPpLvyFpKj4Zr9dEGIspm+6PkEo5Cm285tOkWj5PgkgFv0GTLWJQIGI20
yDlf/PVJ5EFNnLA+6LQF1yWOkIxIoCxO7Q1EAshAUirIVOy1k9M3m2wzn6HCarq4ZwkxzQIpPfhR
eZoIpe4wzYB81OwGGVxZXpqIBc3d91AX/O1kMOSr4PDhSYv84X1ipMyYS/ydcszVWVMyN4uUX+7+
kjL3PjlP/3HpawtvjMdySd+O+yyVoVOB73H2WilSlBPYaIM0sYKaN6UzeXwzoLl7AfuIphLUGGdY
J18lpdvn4JMAWRzYfH/e6v0+0yXWBYZGpJlVeNVpExenO2GuAPh3AoI9fAIoGUWTRg3fsaDy2D08
T0MKlv8J45SxUTgms3W60ny+Z0bpEeslrAJEQOoXhfJVGF8bkXipz61PlMalfXIriugnfIgT1xLF
68TwFfcn+7LaAyy69YW1sISDpEOqIlU2N2YmbRkWM+SN3kxXjyqRe8/hPsaTHqX1PB3j7n8lqS6W
tPxz1RUTd9Rz9fIeq93ivC1bvhz+uLtU8loaDgPkM9kTasTenxRbsnGf6OY36O5NXZCmAxhLx7LR
TENOYBstZ39KM23NkHA+LH6Ju/h+phAWct1bmjRXPMs/U67uECWHluYE4jW/NEErKFOSO/O16cMn
38AHcrQM/k60un/i0k08hDNPyRUPxfFESDpMplK0hVJSj9AEdG/2YiJgxd72yZayII+FeQYhg2PG
14K21QsJd5ltX/kMjBFv0euGy8aeoxDbmYQGDTlW1yUMPhmEvtVaDyDnZZ6GUh+MyH5/VDTzyOFs
LMXndGKnJqYetrMfX5lLaE7PZ1M+MVDtSd2SybPzccqnoEKxPEQZ8R94fjZive7bJUG7KNLIf840
isU8xeS9/k0eE9jBXSEGRnc9NuMtfi78pLHadpXeZRDxSKDKAA2y/bwGMvNfHUnL3MbeHq1ws4nu
sdB0T5WVaeguMEyzofqJdI/gB9pJgfiTaL7tg/KbkQdkOQt7izROuMqiFmafIi9Q/lOwDVxZHmwM
eMBATgQDCafeTmM76bEAlyXFIBbVn5uSDNBzHoaHxtY2lj+icT5Lmz6p/PzoTt4AyLXqkCTF8q8X
ZhC7eCAlLMhRks+zafr0QjeE0OG4FQiuOC2owrwYFlApKzZRYPYlj8Q6zHxWZFDm0lnPRdZdTrhw
XhD+7eX2bbYvhQYZFf29GJnYKHVoTpUqrRqWiyt/hjX5UU2Rv+Qg3SQ3Mvj9I6ms9N9ndVY55t2n
EP8vw3eRb8ibwTuT7l3j6Yw3jTwTQu+QpOFEH3/Dj5pAIuo9EnBOOUfodAo7AEllNkGTybjCLj22
O2Tc/3Qfa1o7GFlLQPyQG4cfqtwBk6IzEUap4kixkfrlrl34ptvTxHzH4TGWi2mTVikPMm/3PGW9
ECwlkUg/MaZFP4BCumiE7RTVs+PTuKRuhochbk41gZThSZ37cvg4qGNrXzoM5xJjrILVJ0N1eE5Z
LcvMIOY1WLrxWMj3gEqAeLVnBhhy1G8KKKKfd+BHT3dlGXuzmW50mCbPBkkL8EFuww3qmi5SIIyO
aqAHvRDFzzuIyJFP8VczNpDnkbm0XIzVPMCqk9vB1BVgJFN9YrxIqXT+kfNpwf27a6PolWdle54z
NLxCPYcMmCUAkUiB7Z7SEJzIP7ncVthaVLaf/yeUQKsnYdOJbPc1n+9TQyUA1ljKdCd73+ZXnkmM
ZGtW9NirQA7nNcEQGv6NcuzHG0JQftwoqhldV0FGDm8Exxc4ypAzB+aVZmwkHkFrzCHtk7aQDVIB
CulQOqtUcoPAUANZD/urM9yFNQqqONE1vPJF0mMpv+BJEreXvpa/iS+U4+/xLvtUOPiPzjkURFaY
NlXsglvUIpV1R2kCA8D3VuqLMvOu/v+NjowHym2iTif0Hm0V2ofMP5mpzqKe7VOmwIhOeObc6g76
8yd0nJ18dwdqftQD/ywkiZyMKsVfV+EArnxG1heKTVNaFnwvWCJ0NzUJVhQaetc1Ij67x/TVw+i3
mSkAd1VsTZZxaQSdCjFDjbpSfpjCw0bb00k9SCkVFYCj13ykjKKwpv9VsSKOwJYAmx4cyJNtGWdP
22MAzCkwj448iHxH7/dBRNgRLJ8sab8OZUVNGTaHhQaq7t0XxJHsJUFxgG7jwBp7WPOczgzq5nXU
idL0ZSKT7SJYV1/Wm8SCXNt6Pihe6hSFO+ZssUBZkMjOgAtQAbB1DZtVPhnfBbytIyS0eqZ0fixC
9WHx78frMbpXv6iyTAhONT8xTrnEkBdKkIt+GNgQHq1+6EuUeAE8lzzd7asYPzAr27dUpAlHeN9M
nAeGb53+4/OUhwtlbFkdaWeumFkz6FkS5/opBC48n3LyZa+poeMTfmwcwvXBNuSVjw4TFjfxtuNG
O/2s3Ps5WROnmsxdz23I1CclvjQ2sNUp2u2DbzpFVvd7VILIdG1SyyHQVKqaiHNk3D7+9frPh+So
BeXf6vqO7UEs2vsYArZva8OKP4Lpi9zrHd66X+GIBZ//6VYC2VS8xrClYhlaFS/FqU/lJDxH3Y98
FshyR9jZkCrc7/bpG8e+erRRGDlf04B80HCP5u/1eag4V1Yimz5dwrHJdULDlUh0G9/GWTlW5C6Z
oGWfIh/AeeCiV7mTARxr0bq9Zz0dc5m5VcyUP5Ts1D6WApaaT1qhemW5gHs1LGel41G9lT0xz3On
/UUcoctI/JG9tW2yOm7yDf63lza/PJAXZJxdH06s5Y0W/zbAipPfkLAVhJeu2HZKrPZTplqo5yS8
HurS8XK6n6vfvV+JClzicbgGfWN6srnd+Gzycl1HC5LIvw7AsGJ1w2mfNrBGhJiGQYwanQPdllEL
x5jPBugCECVLvNgCqnsKg6VR/fE/AcU2BKaZk9EadgFAVqsXNC0oSsHl4XYu+J1ehAnbG215JVrl
+PHTCVi7tRp8y3Cy/xVTVcEAsNz/NR1EbcPf8QkGW1EhELFc8KXSF5kI3kSA26bKWPA49YQfnXZQ
UBcm513p6N8Y4uQOyghBZQVeFHKmnQyl9wNn0Y6BlbZHlug22H+W3rPIW6N5ZnlkGL2J2Q4DvGFe
ov4Fja12Lx1aBzLq2XFw5pRF+TfinoBpuyGUl63VnkHf8TvCVECqLhOFLHOcAueOL04kxG3yzjVz
mkAbKkn+1XyYHH5TptzbehecuUc5tcsjiFd/sQ666ZRs5R4M+r1GlOmZNHoeJK/Eb7h/FV9uCyW0
a0wK9lchsEXMMIhW8XRIhc936oLfoJP/u6pzxNxg8/CiWVru5qXNoogkwKt4FlbEZpeQc6edg4ag
/eLYtJeoxZOJWKtexRQ9NG+S4N2n0mBuE6+Tyqx2ezzP12n3Qd7gDnqsPkDGdAGW+HbZp0UrcSlL
7e/IUlYt9xvo4hKwLDT7A/5+DPSCL2od+shQB9rCyLv+s5eMUCH+Nt2pRBQO8NX737jrJXwMf2U6
QrXwz9Sw7JmoNa5qQIFaP3Kx8oyU16p6dk4PJi8Midvv/2UwsbPLVpVZCZmKnz8mBc9YCPAcp945
ovQnURA2HtaVtr0oH72RPBvjwjdb8EciXt3WF8XIGVn4hYBq33m/4PuyE+SZFqtn00gstuVPdi6m
BrQIjuVNMdf3bLwEdmuSDImZoZ1w5NOHyngNk/Gr9PLTv9StWsSSa9bGRmmQdW3KifSQ9dmD6m+h
ExTJYfRvEwB4YdGtVCSRfUW+5evjxNBdpQE80Aadnj/Ze04rvCZRDhW9ursHzwxVm86PiWOP18Kz
trKk0lsuKEzInALvjonGibSvXw/lG1CW1eUk/rN7k4XryIqJ3eSoAR0odzF2EKWz3AdRXEtpUoXt
M5X4E5uDFr0/KYG4aI8f7S+eQVupGmFtJllWPRRw1NgnBnC9MQ3hhFyNt8fDWWJU63IDypwgwGUv
pdqgu3kmAfsDOPb756woGdpu6NWuSL2tWMSedA1I9igTVutOyDs7k9wGrCs8ebllpaapZ9A6yXzK
EGPjjXdJonPwoLYkszvfaE+As6rM5K14TftbN55TyRUhJwhgZXWqQWzTR9TzD7q9wduFF3wC53bi
2qP0mBDjuhfg0DlwFFN+HCP8nHgCAAu6J1WTECSe3YR77ozKWR73i9l8e7D/m+Y4YXcLhWfLOX5B
mnwb+T1nenNGvg0NtpI5Xi5NfwFRdoo3pcPn1EleqWCF3jP4kal9GAywjxx8gwCDaPI5KWP1tN/6
BW5me5NnhypQOaW0O+lhyuahuSYnHdtFn5qtUex1gwOmlsS24yLRXtA2jxn9pk7SKf7O2zFy1l9h
B3aEdkSsHNW6Y3LLQZSWo8NMWitwKP0dWgHXIxqNgC1QqAAbg8+oAz0332/5snwaH7DkJ1+ssLWV
k3Wxfth1/+95ICoJXdbpRGMZZ3IT3Igs5bJh2dJYUnwuTINZDIMrHRZ/6cz0kjN24HkXHjZ8xz8u
h4zlh/+a8U3MU3tVCzBkoIh4SCZJWUaMy6GJrNj+/JKoqmu9KewJvo7nsOqyca3hsSrGqO07MCgv
nDHAFrbKc2Ne+kBDBmfJyHUOzypSpm1micM2DTN96xmAt+Y1iNLNeCpvV/8mMWHex8pWItNLAet9
NVmsMYyBXv8g8M0EbtMUtg3Dt8FwHOJ2B6yf8PK6Y6kBVmwjTxNNDkxjey+bZ9siy+jxhDxXCnB4
TMd3PortyaMRpKJTYNIvfB29F4ldCoFcj63b/ejidCWBgeJNikSKn3cvaGVzX0N3ruBrzkIt+b/y
O00dkTBHbAcS9HiIHTEUifJLb/uRMxRqHwSrfqdKXtmmleanfKT4xLruqnW/5ncjl/zFtJYivHH0
fiEYS9Kh+Ae47oN+iyvbZL/J+3wuwDMSe2lpVkrOv7OycuKjx1L7F6P8Usk7FDQv5pvLhjYjrBAI
o4aLJ9NfnelEFeV/wSLuVNAMiqpHZPmZ2W0fIdNXZxFuan0qixMCo3nkK4K+il2EBfUovTnj5Tcr
1u9E6r3QL0D44zUDxVvhs0BbQ3tgwAbufeuRGqaVcwpz81y6VAAujwkaf1FiVX6r8OZAt0YBpYDh
12gXZLKW1Ej2f7SGeksN/P3XxETTR82xSTfmU0aRPKNjAU/KQBn5l8izU7eR/7wrKdvh/HtaK/dP
zg+2+08ZxKxfyQfipFyP6gbWLT9PDmZLeZ7UCGRcPm+oMoec1zTwYECSE520CUS0Bl7T2vbg/RKs
RokYWrYpT12GBh7Dpw0mIl7pGpLJt1VEihtotWlwTVNTATzNKYVigXpZJJ1B7gFzxuRw1h53iE0O
LgcjVjcHdIJNW8ueHFiYcltOlC2YQ5CV/6wkSay8l2/TjsghqjI6i2EKbvoEqxGtbWk1DytWPj3F
Vim/3oIKzhiPVLzg6h3EdDo5iTsq2Oq3M0xjcZ092LpoCii8SYazHkp8vLhR0jl2MCekN5nFOKDY
nK52gM7mcUzA8kjL0HJgvVbpMOJPzFv/PRNYHFizSdRFLOSLzJ1Sp4foRwyR2X2PbYj8YvWVyrnR
zyQh9hOecWLLhTLGkgwb6hGigsBWdEkhbDCwc8OEs6UaSjl9+mZUB0OlZiMBjBC2MkYGOaWgES4Z
h6MhywAmcuXo8Qt+XgTlihM1UOD2HzP8lzWoked7+HP6NZWAYGaDjIoAxuQ2sa8Tlshkwxcmkn6p
eIuYSYsXn9CfJ4hHs7w8743bAbR5+dDV9Kgo+3JNIXWHzUElX4sDpj3zNI0QpQwV0T/BWzR2zS8m
n1SOcwJ2hXAWt06oaeHeI1tQcgFq6ezDWaFcPoDYfLummKCYvEZ4KzIrTkDxBXYER0ZDDDCGT1O9
7uIfFr+ePYY/CrM8d9lkdb8vSEZ+QxZjLChf0O8Rzdh+8jF7pUmR0hnso1klxvGN/ZRzZRke/b7n
QBpi1BQD7v+cmVSW3d/mq0Wgt2n4AStULbtTg3at2Q+64EeVgYYYB56Nn/Fw1GQawGOmKWPcWQtP
YPvCqE8HlslINTA/FhYJncFSri0+C7nG11KniQVLt61aLU27YwOn7yjix9BOXAleCAUjHVuIdK0B
bGPDGGfmzToEJlyWyzrSroAxin0LQdui/Gnz6cuI9WsG89ubHt3OkQiN+nE3C1qqmV/U/D9bM1Sl
/xPi6HbVGMUhUIkZp9bjE8LizyT38O9RtJsgcg9J5ZB2Z6JcdPQR5XTMG68k40WdEXe409xFOIuk
wfvl8bdkMI4PGbgEXz7j5c3ia08gqVwvd5mQ7FyXRu8ulL4jK+YX3HgcZBu+IONUXomNWtCPYWLP
CJqrYKwxw5/tzzNGswE1bZC3Nx6uHreCwce6p1S7N8nSJ6ZlpBdaweTr6BuudKaEG57H31Q5rR4f
MkEuEDJyMhHcB3j4Y6jh0cpXwrtRUzEBH+b0iy9TVzuP+CODFbwXp9D/OuMIwwzI7GQxhqulryxs
bidMZicZrOJiAoucCiz9cOCkQOAglIAz2mivzJVFna/xH2Z7BxUsFzYGC2TG/u50KQ//ou/0L9/f
d6bElJCZgglXETJKeE4HO7IdFhSdFmtKBP+K+kYPgY55TrFGkCNc8QbClTQUyLyAp5kOx2kqgetf
nUhyQDt2QcsLBSHhVsVPpzBfIibIjQA93DdCzshcJiHXugBCnmtc3+cOZc2QodYkP/mRZG06DLTo
QeRRslJe5SHQHNwrFOUki2rIkp1Om2e5+5/e0AzhrlNZeC0ssSrFR60VRlYJmm7yCY+Sb4B5+OpS
5Z+mlK9rsXueXYli4K2EezYnO0zFCwplro2fSwqmPtOJTGzMJDKWL0UQZpX4tT+Fxax4oXIQSRMj
mfPcOCPpWINuu+Oyj5NJ2ZBjTPZ/aML3SNHKlCX14qECjKOde9cW81EGqaBLd3gBEc+c7PVJnw6o
guycDEdoFFaJGrXxBQIPMuCqk3ZRjokvOGXqkdyiyOctmARKsRHiC5cPmJ5KOyzPmSX0G2vTGz0K
0w1408Y6D/naJPtjj5Pr/1pgDNcqFq1HA8xqN4oWJUfoX+aBuo5xkuubf9LB2kG/rlt9JQlvBZ01
C9rEcI7BtHT8Teq1TnGzYDTBpYVBu66wo8ILyKtsQRVuWJ+fgeJ3piUsVcuPZb+hxy06OsXY93S2
6RU2bs6fqaex7dIdpyGHz7NjT5WMGeqE1DW4G5wOEivVcHNiPYkCBFjmjYHcO9L8T4BHdsIKgnbW
eCOKj1ms9Ggo+mzWufXBNOPK1Y9YowE1lzjJ3mzBuRHwkcn+j8kmVecSGohIwP8GX62FVbCsCNpZ
L7/1LbLJeor2qm8Bi4H4dM77dI8ge7ypKY+2uWuHlJAqNjsBb+4ptRxlecxTV19u2zILUmIWS+QJ
ydgi3nBji3+xALg3jbWlj+m4Yk5JRP7eofpVoPEC9rTLOnwlGGRfVFEIJejty4A4ueoiKyNlK3Gy
Kriq3AkiefQhATMrM06gQpB+bhkWIoC+3a145FexklNE7PdWDkSLHt5MV1ENYIXEC2IKAv54ys/Q
1ZfWpC8MK7y09NSrW5I6INJHv+mJz0oPoiyO5AYWSRjne3rbm3UD6x0Hu9ylgajwJIDgMbg68yMm
M27QKB8biJFC02osa8iw8RsXdR6RnhrrtHifC4Q7SZZj51Fo01yYAGD+Ku/feYeSlpGCpxWCMWHA
I47ghsZ7FNXhv/1jSwWkDhYA7tNURjGxMKPryHNlBOAOuT6dJq/UIP5M48mE8GZCDRp06KW5bieN
BSrdqDN+mbieQ9Zyl/g+CNqLpUMlg1wtDho3+0Ji7hbe0kCrTaMcApDxm4fezbXYLa+iKH1zIi39
h13DyeXW7zqd8UcjAxjjU/k6wv5qvK6CIcRoMtwZqZswMK1ShVKqpCdRJTWn69xqXpNoJt0tV2Ed
YcpfHnpT0W9xPEuScZ1He7whMCYR9rq5CVHq5Iep0hDz7xpwpTg0tVMS4gbl3dr0T+CqZJgl90ii
jSgn+vXQscjf5bkCFsc6XQ+4DuZcO3LHuyTTjagO1X8NA4alZL/WQgwt/hBkGzWsGvlEIf6Yx2wt
vOHcWplA90n8fn+f6F0zIktWE2n85aMliiCdpsqAlONvYGfrlxWeq62m9pbz+OqsSS+XdENL73U/
yMcMKVASYytBAjXkch/eJEJMLsFed3NWI49CDyafy6KEpeky7Dc9nw56pJ6amWmkFZcrod+Rgbuv
NO/GibZUZccFNUbJqPKPQ40Wqv1VAwrzmjLfpEUegp45FC5jE7C/+FDsj1Iy6Jta42JqsURfBOfE
mgUiNHLiDQtUVGlU2JiBDr8ynVWmo8BQtwiw54F8N1t5WCVoe3x8C4G+QCRzAWB+ZYhdbh0EKkd1
iWrWfMM6GdAuwNtuNuX1kgbu6KSPiME+M2Qb0jFqUeJGewk3KtpP0fKFt3SBS9FJh294dbg4YRvS
DBMqAwblmmNQ7ILXzRFo53AOmz2v7eUY6np7cj6jWeI2aEyrl41uYnQTY/IWpXfJDkgT9jewj1GI
D3xYMugsvttDC2sbHZ111VD24B04ZJ5T0lCZ3m0GmZ+1KB2QxP4Q0ZweGrJSYNOw1iuXdsG74BI8
agzy0XlaFYrz/vxyu5hwGHXGY/xmMxBDnUfNErbA1NuChyWjzwqFKo6pkKmz16zR0FRMadkOHprO
gNPd5ztnX9GcX5APdyrRT4G7zzkKZc9ElTfn5K0pmxYc+LWQrf9i11WaVVFGE7Bp7SNVQY5gsSYS
jfJ/7kNnPON9NXaACuUrL/OCQ+90+d5WNqqjciKEpMODigfGCUgSl3xGaTQ1k3vFi4cSvI3hm+17
VjX5Xl0ARUFCAcL97PyD+U6op4epFLdVG2gMMpIl+FiU8Ux9OM12/y/KEW+kjD3RBGLG2yruLwbz
aJRyS0F/BKNYmJ/7m1KXCPiiE0pIpd+8IfrPYbKj8qjAn6Grsfwy6JOTpHmxVwMj6qmunhg56suC
El3sGuB3REEGctMNzSl77lqtfXImnCwndla9wL73SyKgqg4QS78Rv693Hl8z6zDAucBB61zfCgk5
416qafBEMFbs/5BPaqY3ButLbZ8hMVV7X+rXmt7T9Hln000IpwtXjAMYOs7n9v/sI0I/Nl8+HTCj
3evo49Zqk+HX7mdZKA9zKB9v2orcb2BxMbUC1pPMM8v49zjWmK1AgdSQL5L5YtMtsHmyECXZaGCZ
WIdMhtOrJeG/6up8yz8BniEDqu4tHQch9NOtB/bGF1g+3dsyUDPwDnEZf4K1TURG5YZJktC5xlAI
tSyRgHwaUzXsnWzPDwaougKeULNNv51Wyae+MWVQM70O9LN5HYlb5p49IwWbt21hZUn/hKdOqye5
m3hUtOLGaBRfXIMJSuHM5/MJWIFb3hj8B20tfhucL9mDaOB1F3u5ROSvx9CIfK9smkIoWKop2Dy+
w1cSjOzdCop5U/4nMavQ6oXGlLgxtiD0Fhg6IpkobX5C23jPQq3IcgbhMeHTFAxk57LfOEzj2DrZ
q8bdFsMMm8nft56GJ29iwObiXmmxth4v0LZeAD69KUpyGeN/a2y1sdUHk1X+9iukPQ3ATsk2r5+v
1HZdNj7bdyOQY4gdUJQJOoncLOwxngXRgXxaTauwvXBzf2S7XeFXr/k37LqN+ezll7OUDUKb9hJ3
5Coh3rkmKuPumxzHqfQu+JwGywsy3SRtNrjO25CDyZvo/EeAnFoK7RjKschNyXOfAk3bzwmWZNrt
Rwp8yEcaT2F0kRDB6/JC4gkyTBOmsBeAc+cNSZuHbikZF9nfxpWQloNv05SHow6v2tZunKUcNDKp
Zi/xCId+glVe8DhO3+jxNLHczdm3KKQ5KJDqyudYlQRB5sPxxAwWij1M13ycttoSLM1lk+9o1i2g
7qH4hyih3a7q9N0VjJGeDXphx0yXvpPscwBGDT3Gw4IeHibjTI9FIXUUtLX8u+BWXed2DVOo4Bub
4g+WsjCnKjc1smEJgOEot007u5CYhDZmbRBx9WgEAGFa88KFR64rjd9MdkOAMPwsHjNtGMDASZGI
O1xUDhmuDoH7ShrcWHRZJ/2PVK2gJeO0A+yqG2Hsfc3HiAYi78kcPGL9EMBFVJEys6G+ZhxksYZz
OqQCcUBbNQRzU1HZ+u2B6YgaUvAKpgStRmnwmvfg2hQmqqugBPb15bUR132J52lveytKbqrLCepn
TfLs2CKmj1wPy7viMzuRAvykQ2g2zWbbVokFJ36SmLylDStdWToTMv0z2tTKwKIJQ7DyWMxX8k3t
0JWpSE8leJ5s6rpI5P1uim4iGG7QMjwBYcqHcvNA4zz2kmt8ZuRYiA/k3NQK00a16DspdoO6/WkK
xmyPvqYQ6hjRvu2spyI9CYd12sAovvRw2nUhfe/hVpRgKP0xjcPxgyWwRy/Qxc2/k52u7gdUK6bn
o9PbbuuqqOQ/XgYihfVQu0KlGotKE/Z1gqdR5OZxAqBrfCIGJkGjbNllVgc8T8sUdV/FcvRHsdAW
/aQIrdaN0E+1UGvwfYhk5B7SOgW7YssqNUP5H6Nv7/VbElD5MB99mrXD3KvcUa6ytvsAaEHH40Az
E7zfYqN8HFSLJ6CdYo0x+xWipGU1eDntrk2O55P6CXlNSIjR+VuC+VLUYOJkD2nVYFDTMmdlzsqQ
FhTC+U1VAhC0NZySplqx9MU+IOM86rxwurvUpiTSvSVrAgDtARxrGWOUhNWTWR/bahaLTqrja7Tp
pfTshsLGFr4h8qS2FkmcygMX5di4xnUAHBMZ4/mxkn370TnhavWsmn1+5ddELsE+o3wgiOYbOx5P
VbU6hOdb/DADAeLXEFozgGl3Dd6yD+KQMTgkKsSxb+JBMVypIQBDajb+H8+qBBMc/i3N1tzEX1Iq
3h2LtrUE0DSqWsXeQ8ghRTOw9g31pN2jw+SRheDMFRqc1VVEK0A7S4wnIPBWGedZU8Es3QGSEcH/
+eHjb9sLS6hynt7USMB0HTQAhYDBh7+/tDExvtSVxby0gbFwPwoS8ugLsdLVz/bwig29YOaacghn
fpCF2G9Pw70viGZ/E46dMfur4mo3M/8KD/6cqd8t6G8M+IZilGfy9fCwe8RB4OGmmsDqtEf7VaZd
IWzj+Fk2zDtRy7aeyH+6NRnepQMRSNGW0TKMxkklxwp3YAc4nKUkmynN3FKqaJm+RY2U3MfNVYSQ
M00QsOGg8pIvrJCWiwJGqY7yRb5Nu4KJuBCkReuk8CxJpU3nMlX/f45L0wK46ac7UUWc7KWUwxUb
hh/oX/yjvY7s8nlkDjTmTirMZqkiwGOe6QmCI6qcVJGrrG5ffKOtK7BzjGNHte7O7fes6mjs1n0p
29FeP0ItTxJyHP9TjRcZgGdGLPskaoKqSyMIJcTXorcKIfbO0oJ2YMwDxP3rBzPhHOAXZvr6bkAU
WUzTbF4JyapK9sWkr1Sbwlt56ZJyDJJvdPgNcVb2C7w4gR4zt0Y+PoI1D9ClwexghC2IEGoKT+lc
64VUd89cIx2cC7VISeeoOeOetYRMKEhpCq+P9odhu3CgrXdZCRzEQc7QeSfAYBjmTcXXFZFJn4eX
x5QyOHAclYebbNpVQIBzfDiQTo77VZIHvwcqXU4AHTFlUuxbzuaxi4ecRPb7GvYkHoCrJ/Olaj9a
htDKX8noA6w938QPAlSNUyNRuqVl36S5ACK3hFh95XlPMYJQiDM7JHfmmD/k4JzLPzwU4DKE31OC
uiv82LtOdfiSDVUF5M/KipDsWfO0IDtAnHoQZwgWw8Tjs5Lu3gOGOs0NQ5j90VFcH/BHC1B8PU+H
GatbnSYlMRWOPHxssJfFfE6FWrblN3RQOJukm8JWXgQ8Ibuvim1RhPL97GC7n/mbnZ4YZVBihRHp
jTgT0L59iMptDFdnygT+vKGahdtSN4ZLI0eSvxTyOeV1jbjZfZKDdvD6aZ9Iv8nS96ySakxi8pDk
XEFHMNHm+7jvDb8M10yJBJeu1WTk6ozVRhPFzoHs743f6bdf1bgAxxvY/ELbNai4pw+q6pBB/Ew3
aJqDlF/YFbjNFSsRvR2VdT+wMQTgHV9kD9EztWio2JJxRKXHul0NZ9//5IL/6fHyUqaoRGMlNuLg
WRpguISp1C3Z16/GZ+2QrETR0L6QppVmrNtOoBAyWIMtFlrWmlaQhziYWlmkb83uOo48Gbijs5aO
xMTjHgkvOLysAfXSKbmqzwqyRQeLiRn1FKeBw/fPQ9YB5c4EkaF93W9Y9VWm2curZISiVLgdE9tL
X0n+3L0Au9wItGiP5h7LxGBS2Yik6UuvVo6tsyiYodJNTy/kBjBWHjnKgxj40FZx7F7uRKE/yj+x
bKF+y6xWSIN5nZe2oNueyY9niSJO4wjpZCa5w7DC8SEhXKPEfbd26teaz+iMwlP1VkpIMPfEBZXL
LJG1lUA6hRoYjsyMb3z4aYfyk9gD05oXOMNjf6rXXawT6x1odkcaFIissQqaJaifAAukGHKChLV3
SwKdBzZpzSn/uPJXbVK0T5NHJucpKN7qnfqTJhz5hxTCOUFZGg+W9TrZm/ERDohtOdBkJPrY++qU
iVYT8dh8s332ABqIJWppQhWF4LWNz7LEJeZp3rbRnU8HV0aNhmQyd2rHYybaRLIQVsyL4yld1utm
jGoM0Cg1E871qb670+LCCQMjCY6qzN5AyISmQVf8Ew0XEx5LCsnzhb1oLmZxr3Eo28/QNRE/gkjW
tA0K5yNE04m4CMXyroAJjXeRFKYarPOAt6t22TghV2UZ7RZ7usALqGj/EDZBDpojBLxYeKF/wLSa
zcjzV3nQfevBZSfHzs6w78PAmkb/Bei4qRUXHEWi7YRQR62nD6e2Ejb+kVIL56fJpFdlmH9ujND/
P8Iqlmj2TYQtbLBDJm97JRYPVPGRq0tiKFk9lJhewOpIscmKhgm1yXvewZ82fHjtkQV7mVU+t29D
7DuWDYecmQysHU1peUiKp0NdsFp9xlBZvk0RRe7yStlr/25e8vOIEDQKlr9Pttd8cuRlj6YLXzFa
PaazzOmwMT+LJBqyW5uN4iW55YBqzLMZElKOxVxKLgUId4Ow2esfB/wHz4k0iksdifurgWqp/GCD
1zguT5WPrrgvBzJqTPaJJi31cs/xKDQH9GLSbJqU7lKH2NVyfm/vRUwEA6wGn+h3CFU7Oi7Xe5/m
iyFHSlv1YTzlwG4BfWPeMod2RN7KlhsJoe34j0WxNEkqvvwvhBHkTXtf3Gjh24Cx7tbk+AtOqR3Y
JmXOwrswsLHkzR+QIF2dGeoYg0wAZ5iWnlGg+G6wg/ethghZO372w4HUYrJKmX13ChC+1ljV4VFD
o+Xd37smEi4NZOMTQZONHl6V8URBPAzXb5qgXNDuGB/ac8KtnwCEUSwj2MUZYIvqDRkrddRWgi7e
go/8GsL4CG80rBIFpJuOYxHnEmPnu4+nkqAwJABAP6cGhpxLJB/lIqOrSTq1aToLfwztEUw7Ygbi
tleTVJUXuzIO37YWE9FOtDhfvjM+JKiuvZ1Zfbun1QniYrK8mk5E/5gZMYlAT5PwpR6zLyvDOGJP
+aM/HSy6yYFEcj7+hsb5m5JqK4T0pK+7LA/IitCjsT6/PsGeCMRXoTlkaxPUAwEKH4G5UY4yiamg
hr9n17M9hBfiuo7mfRnnlyVHosF4mkdvYSEHNjoPgnJtcuJ5jR1kSp7HJa7X52a7B42XXUuBoQ3N
oy7NJW5Loll0OuzcwqsTawP/K1AVxqy+sOo16b7dGKBCIz4ta8dBiws7xdVnYZg6LIR75Cu248Ox
08xpGNwg5HufCG7geVIVX2AzlvIJHVY5SYtamORc2BJAWE3//pgJcOtvJOt1SEnA1qWVAC13O80J
kt1SC5982QKvgqHCEZTXf2xNoGtJYSD05LULYYCeh8yL4RM0AhAgACYExTaASsx+bthDv9V7sD1/
XudAtAph3q5EixStmCFTmt1/7/+cJMbcUyBjy6DwdxahZiDdH+sUfLLSEOAwm8dLMIdsYxnzeKjn
zL5m98F2eF8xCjM1WWdqTpxgK6rcCyoi3TaPOBiCo//ssLwVFNePfcfAl/El+gVp9bWY1SIcKxkS
Buuoa7Hhk70GObEUWB5U2UMDj8tcoWYPHOz+PCdPMAh9aMbuqCCJGvR/msbm+cTMNjZ7lvdPfwdI
Mp1aiJyPmE0/K3mhnbibzo9EV6mQy+43a+1/iGxfM3OoV4WiKrureodBQwzyrouVpIH7VXNdxALo
fLRqoC9DOV6NXgcRYa/7+jJWz5aK9eBGB5Y/5oaQURfhxzfEFzGrGnJC1qBOtpzDx9Pt4AdyWTUG
Djdk9i4o1F0FRXJo/LWd6lphI69NaAxnJWXk08hYejtIHWAv2mRKrJhoB+021x++cu/YcbtP0EbX
Nde1llkGWFodNVIXG4975tMUwznsk4ztvzt0SxxWUj7bbPySzLITLpB6u9mIfCsV6D2bD9oe8a+B
ikoJnbgUyWVdgZXMNQxJX9DGsXmy/strAx4Tk0F2nAPzHzZXobNlLOYYbqgCZEwo0b2UUPpp48Sl
l1gHYIL87Yhmd7IAQCYfekdYHARFDyif7XQEhYQnQ2coGQ8jR2M/efStzE5N3KBHatjz0UrzVu9z
DZOuEITpFrAka4+LBJi5BkffRnAPPWAjRM3zvWqRUck+IaZyoQZRWzg6QlUTikzB2SrAFP/bv+yy
Rhf+RjnaDSwmtnsb8wUG6e/jNa4j/6Cf+m7PVUYOoOXVpEImXtun7ZxUP+ZL6SoKrjpwkmJyX1wk
UFINE3eo6NtSLFdy2opNJA48bapJIs2aoGI3ytk0fy9j8jl+kTWj4gWJU8m5kW+ZQfobIyQkPfae
GlHAQFci63fS78YrfqfEKobtFQz2yo7X4ya4zX4Sl0/y7vqq1RKPQCdXBJOOKFYqP99ZOEGsnXUE
/PVp0jhMHeUNu2P1GwqnNBJiYO4nA2R7Af7rCG+h8SYdhqT0qLuQ4QC0LrIl4HksYiDToK2NRM1X
TJZLXK12BZUNaNR0FrD34XvH+X57ATZbliba6qNe8xJVTj8if4pOzUUNsFlSr8dHz6cP/4fG7CBk
kYR694cnWzYIyXLmBhFKHjqNmGvh0GTK40frNQiGstAAggcClCr+lDGcVDBqUFvQU6luWrYzrn3C
RuY6zrc+ehARrwRCEq1B0jVxt87DR/DYjaVyxSGJNxkEAu1yYACGG+0Ln3GALcEtqBuw3cXXAFX0
tVU+chPYbKoG799z6O4r3Ep/pVofzbiDHZCGFFp/3Btw3SLe8YB0d/uRR+xZrtv6m6pw0qNyGgmi
cbbi92VblPXJrfCuWOlZg4v8cfWikECP46mRSWOUfssnHBzKvghNRVzY35OSDHD1G7JH9fnyxhnb
2fi7dS+3w5VlJu7vWEOwv94WUy2ChXCGvdQtmMx+3pcjsVG390rkEZe6X3qPhDCi/84kO87sHXd7
TFTTMV372dEH0SbqxaqHorGin4y/XcE5zadAEnx5JMK9RPJPstuzUQ1q8TiEohR17EyBC1wgTxYR
QKyF3gRe5A3rdpv1WtWvFxFgoZYSZH9dnNraOkmpLAEOoZorUsaNCQIsRtIVkW82apUX3kPbzimi
nsZG2HHJqJERpB9puTkaOeJxTKO4lU12Y9/o6w3Y8cXgXhMiQhZ+WONriB420zvcDswH/x17Qtd8
m+JDEyOGu4WDHpOOfATwgqkgjmlUmIaAJgsLM+zrgq6ZUuqB2FNBpPxZ1S+s+I+bagDdFsVEhpKj
ynH1LBVP8laOK2nILr1fGuImyx4PYdJClyGqq8yHbTW8k3Vj8jKLFISaAfQ4kSPHY1u4qKEFQl+3
gkJlueTNC++FHNMY6XCX8D1FRZ/lHCXo7UYg4DQCDAmF+jLhNGpgwGCWsrvo5GAlE65qc7d7fqkt
iXbjqOgm6mvZuTcYHluoPrHdVn6FmXhmM9WvPhUipZoB1aP6Zkh7qJx00YImrxRWSsbhMTMmYnE/
XhCoZSy/Vtmi42l81bjXGF5bA0cxGRUb+dDuPAzAP57NVr4mlVVaCFDKwCTyOKuRWh2x9J4RJJgo
LzRjntMsgMHJ6J6XYDsN6wWi01LDsu02JoSxjblaenIw6cxQnhtPXnUpf3Aufu8TiH0Pt092c+dG
iT6NnBRY3ywtAnyQnH8CAri+i8FijNrWtZGe0ZlO4zT39eQkvY8X6Y6cPbYkzDSXdfMZr7omsph0
eFsgVlLXJiEL3GZJp3X0SbANIt/Svb4jHzaN4RU2a5NUF1p4aDZ2lNIDn19SXYy2Tc80VHPmEaYp
6igJA7JP5aP3hsgGUYf4y1eQ/GDCUWvboH6hYF5mr2MahP6vJ/qGWwxk4Vrjetr/ybX0cWUH+Xdu
QQrIaELS7eAQspshpcy3dk2mWjKpW7pvUwwcfsVLn4kAqnwwp1wzy5jRbL+jq8SLc/90h8NhZM3H
cp84fmdtlrjvoQZlovNftejDnLMBhMTNRuCAs6p62HF+dumh3NJW95nIJG3z8QCeGk68fIxzPBUk
qaHXFdEebWtwb2TQhHOF1F3G4Uj3oEIyXO7GSf1IIh2d+T6WHDcLTOsOnbZOsReocUfLAHN3YnF+
RLa996kAilz1SnOD+sQE1cU6T68t/D7GK5R6OtdqJzvl5VPLZqzqPaTBbDOb4qqQzZM1BQqQapeB
UDVJKCVTNYbacqjALbfb/gAsMRTa29YFxsSg9xJ61nd9s7vhBi/NghrHnrJKS6wXNcX6W44unAHp
5lfeyZr5xW+EFGlXMMG9TJfZoUxeK8xConL3DMxTrd4pXA4ICc7HGU4DNNroda+7C+3g45ssRlI3
hmb80lo9zP+Ll85dcSLCBcTLBiQSbUjKFbqFSEfQX5puS7h41IBzpugBBIf3Z5wjM1vAKiT65KbA
j6oGJTQSwi0DL92UG9u0BA6QsqWWBsbKAIN5EC2URzEpQuyxqQHiaZeRkSF8DmdmjUlNVR1sUbpi
zAd3b3YpuoQURhiCseZAmBjb3SQ2/g1x7dqdjwfES2Ph6aw57vkxMT3u88FjH5d+mvSuy/Q+mQFN
yufJy/WEYDnECCZumPnRWjKL+BBW4lUdRyxNhrBP50vnMguqlBSkzpp2SajDx4EN+3Pc8HxzS5ED
03sOCn58UiSu7sikBjai8vzDyTnwIMrAUqnPnMhosw+aMTUXWK5/b7JYqnmoqeSHR9mjb17BdJkZ
qwqTcJrrWh2dfMpGUwcefVg/zb0dDsFrFRFqraSfpz2DhfcNeA/HzZ8L8axfGPlFyluLRbrtRtVO
xCfdm6GIr2YRbTacJ3I7zyUOMJ24z4BYNR8XHzEiWokUdKHKuAgDWdsppEAW1lyXKIDZGJqIRgOB
TgB7GyBYJbgVXim8yPoxsI+UHv1F5zompGoyDUOBbxTyWDdpccjE7zmwbGzS5ZF+VBunm2spT8Gd
FiY7x2T2ygYtWfc+HiXYanBozV4RrM2ZW3sCWUeDyq9IEnubVuCDcdtbIGP+0V2imQ+O4aN42JKY
kAAL5YdwJtlO6cnw8P2yK0KK5vK0SMekEXVDbMPOnZpui7W7JxrH7PF7KyFtKAhUbB2y/DCCEE4l
PQrYhWTKGyoE5y9R+73Qsng0daSxY8ZESWVmwaAQgcRJV07XEVp0uVfjtPlBap+jmaHq+iXdfKO8
IUv0QwTjJZSXSrRymYUIcxCC8HDsGwZuiQB+wdAoexqrguJajUHZZOs4cqln7fi7tzE149hJbW5v
Uw+Awczn9JBayBsT43mWBXqzl5uxat0uM/EqL+Ta88WfTRoGGHO3NkT0ESi02FewwQ7qyGv0jigc
B7dpAMgJ52h5rmbD21Rh0DCOaYUoTZvzVGYZ4IGhO+DnffHZnj4ERZnO/xm/c3VsypHhcDwhbAzI
uBk0MkYm4Au38WjsEEhOqsSXtdBXZVn6fcgruZOCIRhfEnwSWQfMTBaSp7NT0uSAV8OEp7qTDmad
gxKWgAF7YORwK87dQFzCMrwVD+g0DbGuxtzq2Xbe+GneD+LDGNMu/yeckO6godtbKHho+bhQmWQJ
CBuyzQuQ7aHKt0iAgiuPlixhyL82/HVhoXYfEKiGTgdakmIulidmKMtEsID5walb4b2SfuBIDh11
3f95U4XzCkpfVuv2mVdc6PRf74L1JuwFi64+x8WppVZRVc9meqUvbVj5htuX9q+R4yp6tlgJH6ln
l/mikfXQPgV3FsMLuQqODfyY14CdGRDg2UDex0A8mGAYEXs7fvmGvSeFz5XdukYwLmkR+v4aa0Iy
KNZVm+ygBxPzLFv++E6qvqfYQZnnDdXXrcHIEaoBenc1yH0rVzra3iD9W7udftxeaG+a+l//6/rk
SaaXMiIlCY81GdygH/aSO2564wZHVzk2dUY33tsxoV6SbFKwqZuFl1sYh+oOejwU5w0slO5KKNE6
NaxqfQlacyaKKLgjVSrf4NSl7igxqazBVWZvpVLAHtbyTcrxZ47rNQrK8OLRM63NR3sw2x/Ku7ZO
m7NjNn81hS+NtXAtumc3pWwjz4ytZTqtm1+7tnglVfCPavrGSLs7ppK1Spwsgf2v+wPi8gVJMVZc
uhL3j0+gZepWmlqNCsXFjeuWvjrAFjnMKjnHt+Em73Wasnl41OMvsBVvsBPm5G7Ye/E7zT3uVkst
K0OkF2m3UVe7vun9n1Qp6zcuumbN5itEE5CrFMjDgeRnuF0og9/u3VJhfUydRb22zVKB5LE4hYmG
6IMthg7yy5VJMRiAxVKdtToXlmPXdFrEF4rgsZWnna//1CxUsXsPTxVmoTmVVsH+jDboL8uc5clJ
fQZ5y+vyS7aPkwwf/NoDMM1uJjiudocSA1+5m76puibeRY7z7QHu5zvBqqB4Jd1wsvU5mpso6fUu
+xKaHoOCZ5UQjOwVJKwhOOpKeDsDG9JSCqRBy/fNqbydQA+beNnTeSG0U+NsojJOJQrQaAKRUwlO
nmb7JyeoVQ2H8RuY3KRzOS8Lv5SY5Hsh64+E7rVicEgOXtYeN5Ydfp7ScAdeQe03jQlS+byEH/d+
qk7PBeyp59Z5avPfY30YGfioNBB890LzbrZ+k3VhFSl5RJH9A5DaRH0rl4nPFpQjetKRYFbleKgi
SrujltnTUkW7cDFk6QPrny46UIDGwZ/iw7nDAHc5FtIDb/OH67V2hz3htgbXVvCRGcBBPnExkZ2B
LFKS/NXirxoxx0YMm0+omLPNYxx7CZPPv+C4kt3Zd3oAFZZszrkTe4qaCBCjZP3KDul9ACDh6DU8
GsbLtT+qH2wUvd2nTTD4wTaoOHY8bGbI7Q3FuKc6vB2kfJyAC69Vu2tcvB2CcdIbhFaYPtaOo1fH
fD3PMyKmr9/2r1zFqOHrW0YX1ML+b9vPFf+FNJ7RTKCV298Fa8VZMw6xrHzQnnc4pum4Dx1oRcN0
g8Rs/ow/1xP/FuRqt6ptncLnA/ZN+AT7Buk8AIBhpJQhZSRsIMgTLhQapVHpxFIDIB8wf7E27aMH
Nk7D84SWLN80IIItlDYdN89F33DVHB1D6SNOh+UD+IIBg5dLr/pxxRc7X+82lm3GyJYByZdKwpDs
mXrsEIBWW5NPpvkEpGVsQtFXLS3v9IPvWQ7H/gH5oPFgPY//MpejxxFRXeArEXk9Tn7bn/JQvckG
AoT1BGG7Jmq6KLfbAyVXagNUhTfIDEyBGmtmp+rW1cI3C2nLtYY/5hDIK6LWLWUWT2A+5Fu/f89h
zdfLX203ctM5bBIMvIbCPkkvMEcM7cc4BB+pjsCxN6XgpUILZf0S/IjclpkoBoWS4Yvx2u6sVy9h
hht/S2bxxfLf8TXt1jnb78JbSrOkUL7RpNH9w94wfwjKe/yL3Z/nXl+t6zdzkG6p33sWs6tVr4WP
2nS6e4jSI95spd0tWPN6m8ZaXSvxHcz9rP9kOcb3nERLBbSkua7HZTsSjbzO7y10l3cGAlSKXQdw
j8WZwoqb6TxFPocoYT+DV6quGaFkDQJ104IgC3Zfm+ulgpFLAuu8Nua0AHiMjemkQAc7MMBjS4G9
jfd0/klfZW/vRouTAO4kVzMgD+86ylhSOwhmy8C2cu1PIx3TELDfzo84XClpTGfbERy/igyWflCx
H+/UELargpT+IbDFe+jDCvg4dkF/UUVaSgbMDftN45hGkNCGDGuTwwz8surteQvvqDW/NNxyzs0U
fZiSinmEwTmhm17HPX3Oy9HoUYQv9ZBj83LpDevV/zKyFBjD5lp6D81RBc4QymhXhI9sBh8h/qQu
6YRuF6ROM+XowHL7XAcThepOdBpNISnWYd1XF0knJmpcxNifniyaF+/vMIf1fNY+Zt9kSSxf2qcO
1c/iCjpl7216HM3UuYS0lz8uynvx+2K+n+h68vt164b6HyfLpzckcBis5oZgMeZl224gSdyTmQ7b
i8FPn0DcLayiOs77UA8+Ekifhow5U9YMu/XktSa/dZCsVnMkzVNMzeGcUrN6yk2vyggOrTo2iZih
i0Ysot5l5O/malTdlSSwBUGqOg66jUgTvPyx23nIS803P8kCmHyQ/ljRc6052mXuivpJdJD4xlV1
vjskN1AhS4/Hc2MiqMWc3QzeBZAsTrEuF249TwYmFy4bifI1Mg+/jy9JrBf1kKtL6MFh2QDUSW0f
zHUDMfQdS1j55EZV8Ifw8tXU7Vmnqq7zlNyfn2KEmr8HcH9ufWK6xyv8EVxGfp7U9zCi0KC28lJE
1X3kARBJO1FTPNtJ0xY+StSzAaVJT7OVdQDE31T4wP8tRuIdE0XqFNDUNPG5tdg81UCgBYaDgGQE
yV/cZpE/H04UgomtxWM8deuzo07N9UhakX7ktcI0czXoOeRT9NBxs85DD/EhE2tkrpG32ewJx2bO
Z1Ura/oaK8iPmENQQzH86b0a8epTKzFvUD53BY9tFJQRWregxHYzk8gBWwT1+Hfh36z0fSn92i/W
L8nRRfnSfv8Tc+fg4xGiOYQ5C7b1guxQynndUix44xFhKmNMDtXeSQoVjNJkAgDa35kt5cmMnB9q
Njyan/KA+QPjNzqZI7QtIEkSYKHsRpCZ9YJt1PyRqIw9dsZX1hyJgGz8rYatXEqlKpULm/dNwNL9
bE8s1M5SQt8XdwBL+224idyX56IrnI82DZGdMx48rSxXx5b7YgiB1XH1EpqmMePHDKknQlI5njxR
36VQy1NqfClTsfmasJcI69EoJDfj0+VWliyTBWW3dBS8y/URBER0EIzPol0XBU6xlByRC/tVeUfL
VySKpKGL9KHyIM7/XV28UWzMTNYgxZ4AEY0fOpfT9uivA9Z73J5ujEnTQlCngvwo/30uBPN/b2Ed
YeCrGIP9GGbXn0qmU6izy5iTIy1hRo0dxIhIG404/Kbd1BZskxdSj03hp79uhp1t8swH0SoAOsQ2
NiB+H5H2cKnY2zdmc0DS7T7nlv6NXdNF30ZSIxoyGTwUC9BnC2JAGD51QHMNWbkVa2s2rvpCdoi1
5BgaDYhjpYxz5cI4UzAF+pHek9KvcdkoKxpWqeEyJ+bzlxJSkQ6LlWg+tXdbXOXAVZ7BN3lfmt7d
NivVbxJ9V3EWrdvM8T7Hk16MzJL+McA7lUWs0ziwpEoWoEhB3gFg7S0dgA96lCScGgPOBkBlLuTV
sKX0nfzOUuGEKe+SePd489pDJwIS+lV876se3Oal34esthESWzuZNMxwmhGxeQkVN/h7N9XpmRwv
vqJhZZxozbNdQ3EZBxd+NeH9nwQxaCjaoJfVl21aoDQ0Os6COvj6hCNy8X5L58l8NayK9d1O8+SU
XExSwLw6kPv7mjk64rfA1oKWRc4l3u6qizgAn/4Y99gxt0+ASoVizvfnbh49Th4wkjoTwmyQ/Z+G
30svheON5oZeI8CflphUNllNdY179KptiYfMqwq4UzRqX44ZlhZ50+7LkaUlLBJ0IV3b5hSPSqlM
fJy1yITBl/9+h2G+9J0beZM6/QdB0uvvXte/cdB7xA8BNKawOkAaH3gI/xWZgqro87t2A+hukXi1
qxVJHIREJb+GVSsCUFP+e7zqyuglEaYK/tx4jJt0n2xWuUIl6NYcwLXZXjyG1hUrzjbxr6ZAHsYk
pLu2Cvxqk+C2f3S4hhhsqV7uKuGyHUfixhm+D2GN+UxZEeRRAsEUUiu1SIg4yGh5TuX+OTwJKh7H
8+f97+yMuMwtoOQGUS4y7SxlaveJEWmWHSxh7DLVbk50ER0k0mUJ+rpP9HFcD1EBWoG0eDiPmLSF
vhXx8F3CBBRDWcs6X37pqKEnLP6vo2lwe+s/3mBVmUpsBt6zNOzzzibhZPcO7u0Na+l2ay3m8xzc
WgjFs21YUxX2hn0nd6DGuRCgo8wumavZC+jIMAy27pXTXyvwAVtL5NVAX40aa/ukUcqbnadaTZl5
ninQwWA9l/HEluO4trd47JgO1tvfAa0Bb6sSQVuoVFlHoiaq3nZl20tWT/7zckJMLy5qqxFMP3d3
TTmMiafvTORW41W3Y2LD9uWdwAk4kVi7b+tujdklFVJCfyl/928P//SDpx3YPafnGGRN/jeMfmZ4
qsH1RWSGYRMX0+8Mb/F6U2F2DiRjx51CYPKBX562VDTeOpR3/b5M6Ih+UpPWo4R1QlzBnJPd5MhB
QxHjzZVja8/PRAasOH/WpCHofdBkVdtkhDGSI2wihIEXi70AXAi+wTakDMGznhm/ebqtDnGv2+Wj
oxyFuPgdm0nBd+jGFe2EOacV1oCld+0zMb4QWzDyMJDNmOBFbModiIIgzZPgNr2CdRpJrs7MPcnH
2hgox46+u+fXJxmMhSvyIz4HAqJ/sgSjmtata6f+AFstMieWI4wBQOswvPzFlKyEZCcIbMdgrGmW
uGBThENZqAXKFfW+Qg7TaoEtSuHPQqCYOojdOYJXTNyC6y0qzMX1e+MDD1VC3NFVVpNmXkqKg0i8
f4fn09B0Eaq2gSXSTJraF8jjvidPsZNhdagaOcUTCUAeHUYfI0x+sjVUn3iDo7N5dONSJs6axj88
RifjdA5fUZyEYCp4ZltPRDhirlWda4tPZrArN340+e79vnXkBp0c6Y6kyGurGYX3n2IieXRk3GrE
vmZB31q9yZecwRVaRoRq4DgUhS/Ja0fKRGvbpmq/RKhvO8yaYbxNOgHW0rta4jk6B2noPb1frsrj
XI8ULKuqbuaCNa96rp5Xggfkb+q6bbVM7usOjagvW2DmqbLMgwonwt9JCp7C/sAuaX/caTukEopm
n6uxVz0HAtVPjhuo4GgJcaIDlHeisRczkR2afdZqzuw9DVtMDz8MmjvdGARFoEnhWBd0y2dSRmyH
2+dWP116O+mFwiLcfK6dHgK1b4/41F8N2lgvHOjPOGEpLK6gwvfiLbOK5XXB3CZcWbxmlm5R98Bs
ABNoJE467Wd+wPvSkRbrG6nccUChFC81CbPC+0vRMVI6gLJtNuMeEu5PcRBL1MgC9PsvvNVLrgri
S4uRiPUpPEdU7Of/gPZomdX17YpAs0kJSb4cB7TdFHLaWmfau44VI9D7vDgGL3L4sVq8LhGj+GEJ
ekpbwtNUKaeMTwJs5sUgz6h2lvrW7X09wtuwxCCHEAqP9nbrKGqFRRNF7ClyvWHciQ2o8eddyUxW
g/FMe6Ne731/uFCyexo1197YVAmUNIeMv3P/TMHeOv7o/i7AQKKNB+Roe2unWQuE1wy30YzmzvCb
FvkF5ckLVzWmHKCeMhc/jI6fNkcFNxOrkX6JjaF0FPym+9jp9f0xdyPh6lRgfHhi4eFijMQsd6ZF
AYW55ZK9+iZwn4aBEW4h5Lh9ga3eM1OBbchdxq4Wspt/bplO4s4UnrdVzm5JQ74PU0012I4V74Y7
wOfCKHhKVDG+zvaJ+GUZF2UYnr6DNmgBpOrWWqOgx8/hC+JlFF/hR8um5J6Z2paUU85RGbMQj/aG
52qzPGqJ2DUHRRq6x74cPHM0y2pzdFHcYKhmVkDQMhFMiayRLmydyty//HDQT6tyZxpzNpNbgnPM
5u6AqY53dYx8nI5TAVZ854x7+udl5tuu6kEDF+xbiqDiWkAXFsNfqJ9pVsu5bZthDf/TEO9AD1Gw
b38T0qA+5TLimoAyGkD7Y6JPQnzURpqxDrgKkrgQCLw2BczOPXj2Hsswexr6JHMVwZsOXZnss60q
1QfEpRq7VK1gBfIDshTARgycQ+0A1BakiUqP9fhgzBCErg+fVwrc909QN4VaZNKnLGOLGnKbDgXN
TCC3gxAyMyIuPGY/d4ztVFFvVJ489j7BDONNI0uV/g9LCymm/6qBw+QyjiHmvUL+v06mpWpKzkQU
uqhbS8beP5bBafg7cFOgZpI2n0BuboMCA7oXdxwtsJBTc2BESNxuTwkNZSBX4itdbqKQ/kNr57hA
FWe5NfzglgvHVj6PEoifMo1A5lAfH7UzkOdgOVgt6OY/8mRLLMPPUQmHjXKMkQQiUNDIOT7Vvhsr
hsvq4vKwtlyrkRAQ81W414PtvVlhE5w15SqC7eBA7a09yXgEbG+1nw8moww+iAeZaZrEgs0z6XEq
QQ2Ct2XTmOpLb8nEcK11Vp7LheM44xW36tq88FJ0n+68XqmyStQYcWLuIOhFqp5ggctw2EWzL0sa
i1S2FP1eFuZvAiNzVS0yOPKZeK3QEQr6+Fgnk+12Y3eK8w8IBfBIoz4ghEEjFmIEuXFxSq4u+RhN
OWcHmQrSZNl/TT6mDpcPrsxC/yAgu87Lz3r03kXhU6nzkdijh6ccPY/TThfB1/+Me6bOHC3hDWZ+
qK5SsDa+PGqrw0rKMzDFBy9Wf+v+sZPSj2wfM1kflDbbd79/LJmsmZvxZ96kF56P8VWv4c3vkvBl
53RCROg0V5H1S1fHWcwJi39KeotqqNlpLgoIYq1+l9j1XGi0xvsBUhNUgfC41/LN7hc85x5UZ1LE
2fxTQCFDLiAbN/5y0oF1X8aJBGxu/el/cBSvuYYVhP8JopCQR2BC2fcZNDYoeGla5y5dI8sD62V/
7+9L14d6V41We1PBOpl+LgX4LpBZq7HGNuMitH1or2Q8QupK+Ezt1K6EzvRH/nfEq19VJmuCrpZ7
JRYRBZXSmz+9off9l8++BIvCKWhRWJUcHkxeVCVKslvJ38AecMg5j23q1czwHCbAtT8a+9UXGhez
qVkT6eUndsg+AlaDQ10GESlrpXFRBFAvsdPVaBpXDisX0F6t96TLgRYgTnAo7eHlFc9n+HvERHdh
wqrpdPigqEslUionAG8LPEcXT/4ZTVXWqGsyNHCoCcqI/aitMEQqmNb8O5wPJg/tCRcPy8iYHaLQ
zJrCIvTSMr3UXtHp2na5Mav+N070FeQiISf0CiyHrSsbc8JjOMfw/I/FwD+lFu7w540JXS6BnrhW
gGNnp1jrMjLr8DAVPzASvu5t6uxwXr6GGxKZYZy2tBREJJXgbds1IOwT0W/TBzp69edX76BcLxWe
q7noTkQiB9DZV680iABIkt7uyLoQvZELpovVe51jbeaWyE5UL8/nk1DiFrmRLhYTDxD6jeHTyVur
kBrOcuvq97V4GSXz7O2i/EkoYQfIcUciZj9kIcheAFaiuS8DV18QAkbbhz1sXmed7dnilaWAyhS1
uBO9uN+S65izi1sB2/dj+ZYyOvxZC+eQmpyOHVpTtikXjhIpiLW9jDMqpZPrEkma6QVkZu3dqFki
rPq6BikIjZpVBsU83bPU16o6TPDP7Pva07BleqaQRsPs6YjWGfrjU0N5Utg+Dh0DVeYs8NQ0vlQq
Wa8M7g5V8BsBeXCOyZ44Ua0uDTMeuwdL3iQFYH5K2D2DnjeVniyMOlGzPYARItSTZxvwCJr0x29j
NR04MBOafIAY7GVdzB4bldEZ28qkNmozavUcDX4R2mMdwU0ZqnwzJASPsDlCgI1m4m61mf5Iq2v4
F+2Htq8mQPU0homyJCujdADbko4TuyX9/yq/bh49B/9SUuR0BhFhGZCQ1yQYVI9Eo3IwaXk0je1z
eBJSNCf84ccpiCntDaPQkTiJnxDGMXxmhh0VMIZrXgTbLetaD0wao05qH1iXkJBD+gjxUEjLFXlB
nc3t2Z8tZs9ZhaGYAVB820swSqZhbnRF8Betu0BkjFeX2mOmpb9Mb/jMB4tFmqVicCMXgfe5vPLf
8XZMeO8bNGojz0DP2toqqMO1H3sdaQjQXzQAdhBP1H5d6CeQFLPYoMdlittwW5QnobXKuklkZ+wV
8An6VEMFMZbE32dOGbgfjubEqt2DvLZ8KikFsXkjX7Yo/ZJS16dPQ+6Vekhg3o7VNyXflAzjQ0Jz
gFq/+JW5fSZPYcFsbHjkx1YV6dHyq+f7Bwdr5XJEVFLtDhII8cKPlUeRJCfURNilPZ0iOM/ptl4r
wL/NvpBuI6AxjE+rBXWxf756aB+GnyqJDijondeLhMPO7EyrdtxUcKGy6TJBzWbZG5n7jwy6qWAS
FJSqvm/XXez0zENCiNehnS0Dd9aAwhBcMXOFwEpCbfgwXilN5ALgOqfNBfpenDa4Ej15l26hYfZk
9VmKSRtxfN5B0Jj7WsUl+UQcx24rJyQY5+7Jsb6SwKCSiVuGDeksj6oWpfldaUOheUnfE0CXHgoH
hjYTli7jma1ouMSbMLRa7Qy6q7snkBZqPG5PHU9onQI09JWWkKrdf4ZedwnkxDIYjmX+w93h2J8M
xnbXej2TpqXASXPF5+FWwBw8yHSP1mSRdAvRZBJlipIsciqiANsKC5QxEuVTrbRHcBlqq/OyIyM3
qyMCGQz4vLdr1Y5/e1D/DOSCH+LJU3Q4ABkhl9GHSu2sQ8+MQnCFng8mTwFq06qdBkD+GK6jhQs+
SMNh7gmkJlkHc23eysd2R5iCx8r+DAaI7YaJyAWggFG4ousSaDJwLPmGI1bnyjXrkTCCOVVjN8a8
akPD3zsn0qDBaTYlNwBCJsW5VIV5mvE7QWj6lP0vl9VT/whiJsLbUyd+LxzMcpYTBSxR/hW74eq4
JeTgA2lwnZuMQt72IPGnEwYGt26IraCtuw3eLQVdIF3FS6k5rzYUEt18vnpaa3qN8aohSLwzWo0n
vu1VERJKITyoMMPWXPhnrBvtEoRt4x2hT8lbzkrhYDgCqlJ1qqSrEMyIlhQTZdowntnaly0/pkDg
uwwi/C/PMzGvXF6p3lLiwUq+OMoQBG3edTuXEaCESEm49zbLhvEWGJTh4N5oON3LWaf+HZVUYoE0
wzaxHX/0/Iob79iawZc77JEXZuSgP/0dvQQTC6XV3yUlcukEAOwCwULPSh3qGGvQkWYXeFpfxPZY
gZ35OlI5pbVeKqmQ9LWkv4tnLiCDWPWdTjCUBkti2AcIg/JZg43dGzenh2K4q/YuQlarA0t3A2ZK
9zoVJ91w2hWdbmhit66cbk3kjnwiJluTrJGSs/hDYoFso/zLjQ+ggpGYn6526Bvk8J7w9sQcubAH
kkshU0KqdqQCvLrOhdxu6ZaEGTXD/sx796nrTA52EtUpPSqQ2pmsohQYH2NPZeUfKepL4l7LUSR1
WUteUKOir1sw8yNwP2IhSsSzDBzVC9oToMu0B3OQpMZt8995hyH2bB5j+5ux10gvizVqKxtCBa4P
lRT+LCbQ2Z0VuH7pDD/59kRP1iKvS3D6S2QD5HrCNbPkpacd5PlCDaBp9QYuz9+ptNA1dCScP/jn
co87JhS9qpYUzxZSKOX9PUyfcpuxKe/hRY3aQCyu/DlmkcHkqqiAOWP8EhgkzxD6Ub3/+Qe0YTSs
9wCK/KMbh31eaEVcOF7tsnfOBo6BkvxkMjGFvbn5iH6/V1bzpzOOPmuLXCNPgbS8HtZ7RdRUaZl0
XmycVv6VYVZ/bz+zaNglYKrgtBz0GCXrg4mO6KcZmx9q2VXyzXfo/a0BtNyYW4sGLnUT2ozlFMAZ
iSa7NPruqXgIkdr7IWzRL21hx+X93eeOmhZ3vxOa7exXXZWuaXtup9s7NdWLnA3lnx99W+GEFaQS
kt6cwQY8AzD24rInAzWu6jUEgkBJNy9cFHb6AmjCniTMzD9SR/RnMNWaJoIq7RkRfwPhTyhz/svj
vbblVu2K9kiG2YYWu/YAjsCkw+x4K+1t7KJqMd3+S2rh/04n98MSDfgpPMmBCtZoSrVpkajFdZZc
ksw5z/VTb9q9l7BnM3ae513EktAk/i0nSuL/V9rHfQgTl2BVCLg7XKQSifM1Lc5XSK0e+DlJTdsb
RZCPZqoEY/iQ2v0Dsp1S0gZprceUy2zBasenZQZuF2wormFzk5LSw7K8/XUACwcS0WVA1cXSsiz4
YhutuCHUZiPInZsrfq7iNwqkN4aUgr4Delyd8+FSf72JGyqriUbzGETSp/XcYe+m61GxqqTexJDs
fWYn3ZTYLgBoSHsPktaTetJzAB9bFv526FZ3rt1fQFOIJwsk2X7l7xhKH4AH3I+PX4AZ3w973gds
GgT8p8mOcc+w7riANC6bojjuFizJAI41laMoKTzNSkWa/ohoMcVdyTlxEmjMaOx/a5q6XiQ9iC/B
2hbhUxK8BvsG2KpzoDRCGrJwMrNgE/m74ZGdFzWTzqPyE7QMyBt1fGcbqqk0XL25c0BaJIx51A72
MU66whNeaA5ccD/mi4JZEpRp3w1bQwvUu7P59wckniZfBwufkXIXgqV3g95yqPXwUU+pl13g3q4M
DfJ48tTVT2KdsJJtoGT39RMfF5dtvAUpeixqgc4FW04d2o1l7tBo2fJ6wrxs7tpHz31sS5GZmjye
S4bwNS8izTP1ZmTPFWh+Ei7HC6yi1/g+6nK3tanvrRruWeA1FgVhmS3TGlwpRwDiKZXKa3MtdwzS
vsRe2FU7OCCBwVCDsbRVSeI/XIbPVICazYSjIS2apN5u7Wj6JoyoLfETMDmY75SLXl/ZKAuzGREU
ZquX1BgKHrPdUF/0e+AYTzHICeqWnverFnwvPMuATuy6FlNzOSWxZwCd3vwzsqojvlGe8qAgUfQ1
WMzXeadkaTrXSw6qu60XIiXoLxKH0pmA5kwyIom0xE7QrkL99R9J9sVCbNxHiVaB/G5JPgGygOBr
ZM35oesbkqLbskeREfGbR5OZqv1eWTc5SSG8EKABroCHaUWAH486aqQEqirwARX5usITTVrdNzz2
m74bQvai/Lkv8XE7fgFUntUjexlOa5PrEUb4eqEvilX3pTK0bjLmH5jgQ/gd5STRxkYipzY6bj9F
AEjScu1ZW0xTWoTYxKob+leQ0TnFDThsFvHxmvUHYWGek61s9uRYpFLMyYWOMPDutRX1jZEPTL4Z
Hs7hfVyPI8yHIeYYlO529hDfaclIqmWtT09P/exlg9S264codGLr8Q2mpjogawXhdUD2OJBJIfcP
bN9w1pdUIc3//o4GmOXHKD9spWb0d2Nd76jCHn1dmUJLJ/TVhBaGxWZl9EV16RJzOYCiuv0MI7c9
N2HCTOj5ItJI73SHvHB5p9rprvKirLuZhFBLoXzG5GVSmkchRoow9DCqwqpdbJIWAnuBx2UItqZJ
ejMV98LWs10DS3RUptGRpwVfMnTbAiUvGG1LGMKzjbAiYhOGZtlMua6/lYGXprKO7cj2+1TR0UxX
ahxW2gtbaOUU7GjOMBz+mWnWs9EGYn505s/UI1ANYtaZE0zc0PkV1x0C3CxD31S3R8jHZCFZQT1L
dH/V22gQ0TPf+0O46J19XnSBGT5zzeYqffTaCnERqVtWQAw4v8LmLdMKGXVyS5rWsXxn7G0F3GJX
BBDRIZlVSc8aRmnYfNMfUfBgreHyVREk9m+uGj2tuxiP0BlIarnKtX0ji4NzhdxqlOfKt/ZQ9ObY
axISZPkt0Zo1fZD0L3hnGI2pJbQEjU4xWBFIwtXYnnf789Z64XuTcFzq+Up9ePmLBebXSxbNIczn
6PYOcqN5O/aOPpimRIuzLk8cDF77aq0yNO9C8H1ZvjjI4DGFckGcQvU8J6IW+fpRaEeVX2+OggvR
zMlGKDN4IOK0l/o6lixkAiTMu7V6yVOAJ717MVAxdVxLYOR0lVbU2IKjtQNQtIY/PZlGb3GKsVae
dAoKy2eJuK5/fXHdGjzTVe35MJsPFY89yZ7RARMadT4ohuNt9K9v5JqbAHFaK+ScBarRQxrcYti5
XN9H0cJqpwzVL4u8a0yKPl27C+YuCUt68cNH8fZQm7HCyIPlUH8Z5utnBGiCvqygu93Xk9j9HXUe
z4LG/0zuzK0T7Hx7rF0DXiJZtn8rX5zt7JFVdQMnTvqFy4eQXqb0JFh3H218Zk7H9zei1CsRlU8H
Pa3Zt1mlXaOQT1pbJ//Fy1HqNMTziNTmppC4lxX88PrZqrfzdqEOrrq3bPenXPLUMqYm9kCvU8k1
F3GOQtOytmieAbIv9CYpgNcQaToyd3NGVSnR5QZfiplqzwwaC50+akGwcss8O6iJ5uGlgvho3RCA
n+dxPEZ4HgnOdPLwHCtPAngJGbv8to/Pm0G/n+YYTi2jcHroHOqYWBkjMhv1ntdHm44KN45gnrJb
hlGis1oXoIA858dA1FgS1s01SqV64RNwZ2mbKmhP+xFd4KmjNJaUlasc8ckBFqrsI+rLjqFq/L4B
XWBFI8RJadQUsqRZ7oh2O7tPwwzy3Uav6MoTt1yea2bebj/bzvAqfSoGSZOdkbVyPTtI23up0RiJ
PojFOgj02E8ah5ZzFkG+GE9JPBSLYf1VDe/6QZrW3CuZYRaxRlJJVLqAunxftiAH43InymFVWnfm
sSHHDVnZaFty65YLWigW+KCv/D816jBQu7nzqU1h1IwlrOqs3kkuofIQsDmyPVB0SYA2Rq9Kj353
OQYFikoVrZUNqsaWUn6ZZHnw4mKspOmufaOG936BuKdUTVKqs7GNuCR2MyjF86qzR0bBmgad/Bcz
+JlV4m+nC3QTaLgpu76cR93ZtP0VhT7zZ3EIjbSO9NLcPiVMbQCnmEkg+aXfOX3viZXBuzQeL56W
n6iFB38M86elNsevTGG/u4Wto7tjyL5RZLirg4onOnBitN3GyFIGpS4vtc53+hGmTEnwYyuDCf7O
9Rhdf1mmm3WqD8QqKEGB9ycP2gT1Lu9rBjAvzuwm3oyuToQa4pVqTHJAkksu1wr+TYEfevKdUlIo
p3eXWTbEU2KpFxa6pm+a4+EFnXVlnkSYajEZ7lE8ATVkYjjOIASo23+Gr1wJ+4b9vhXjmvOZykBn
etlUhFGKyVdM/HHBqumO16kuX/fE/KgeT+ZSDdjdLqMhemy+DYf8+KZf+Qt0HKqrQG/bKygQ6LYh
X77g+fdGvlInJY/Y11z5WCflpfzAKugL/tu6sP1+I08d4ny9AzQcXToG5jJHyOmHv9aqaz1HyQnY
fhkUdWNx0c0bKayjNDgrTSsZ6G0yraRlunIugNACdbZKVX7zrTevBCuxJcL9N0FQFnEqribPNL2S
XSi9X0EN4MX82pzeheH5wNdiZscmWDkJvhcno52J/US4qtWyeKtSvaWUapzOle8pb45siXLirtxg
YpQrezpdg5lO/In/8f4baHuXb+1NYFzYJ3uItrl9/t5dYSqCrY5cpzx5iGFwpsxf4Ug5zOyyl0uf
SazhhuA4JQquHMhQfhvq5W3EmwcDRnV95sX02q1zcvB61lrTn53c2RhQ3NIA4+FO3Ss4gw/FlArb
JIh2TkQSHGBoq7QdL+OJHqKMFTODW59KOkAsbFWcN3exvsE250GEtkSugfkQcxhiQc6g1L8X7Y3U
EoqZjwP7YrQ5plqCMzdIQm1EE4M6yRhQ82gSXZsTDnpfYKPEctVBH1JZ69l3swyI6adUm964wmtU
BgKTMIWwLwE9v3JVUBmy+mmY5y4uDBGOpbi+fSfDNju6MX3ju4Jw3NXZ5fgoWFAaEtOrCM+rHJTA
tmqeo1UVIc+GovQLX2pT2fkDaf9gZvz0U6BOyF75BRDES9Mpm/32Y2Yd4QI6yHQ7IG9iVvYjgX10
Y46wNfb6QJ9mSR0J4o70c/eOpGRdPD27np7oc4wL4dj+G8wOWnouzkwz4sAheyrx5bMJ11QFqvph
ZdQTPwNQO9qSHLg0s95D9XB42rof/mbCWvKcQzGmh0nsgDUUupVxJV6oqAl2uLlxtXtsTuG8zK/o
Gm4pBA7pVdv36lQaH6mCVoBWx6vED+m6orIxkQTH/yNgQzm33um3uvOXntjwnDecynkaKAfqQ9X9
v2XP/32oJgf8yVnW6HUFVPAt2fB9LSrHmqYzdWAZ4s9ZARAQNuiAki1PJl0+2vqnc+54ZVPCeVrd
2Sx5HhOU/R+w+3nZcOl/YqKVxFC2iS7GdioC+aHJgLwwciJmBCcd+ZibVNpIowJXXQ+PGDx8srZM
WyoBdqQ9GcCMCRPQ9cPqhg7DeAGopVLzkE/dY7vpXwFAGI85n3vuoKyUufG6v3HA17iczgzZP8W/
GtiS2jm7AFTN1Ja3UuY5Vf+7GC0UWNNDfLrsCPK49IG3q920zNu+qTNjZuXb/d2wD8VBCG7PCDTV
9vGK2WFxHWo8a+WVEgdTYhvOSdg9EzjaZzjzexdJWD2LP0f2wEOHNbI498iE/88uWGBncqpwNSBj
7m8F9wkO2O7uSunlKT4fcNYB1CbVPWC5EZRMYmPt+1tEbt5LxgPcYlg/tvVyvWE0j1e7rngqHpG8
ttO1w03cJM4wspNicCAn5+L9GL9Wuh1d2428t5HxrLBKvbVnvgaGmEN1TVK+mi2FZDohB+ShqxtI
FUydQ87o+zX7Ci9C4CQBudEqYMuGvfTAPkSidEIl6EIcpw73OCq/ZJwrQzmKwm6HCu88EXjWlFje
XxvfOX6w44uZ1yA59vTSiWYKljLqEdEVP8lGJZ30OyiZ2SFs540rh17yS6/1A5k34SgqHfr5MyHx
IROTchmMyvpWnTF7Jcdiu7Ffcw0J23Q2Cg9JVdRUBxs311WKwIuU+i3SrKlyHPCVvrKhX9mHk49+
u5M2uYCTFWB68JTTUSy5MuTiMT899pcdvAkCaN5e3SARgkI4YXSCv6byaDo5JkGDX4QfI0lAoY4X
DdUlqG/pWEj6Tq/zJLzTbLD3xD7tSeYchc0bPI5NNUIdoUTZmHZlTeorknZrwnM0c3FDJQqQtuwy
t5/kT6rWojyQmYhbqCXhOxFb1YiDa+2I5YSnhoLcDkf0+bEos1pWrIrNCW6uDbjcXYm8/JkGloom
Rg7eaAoSrsxPRWczP6nBg/9lFG4munP9bciC3FQyHe4FxAZQ/vzKuBRrHyOzC80oTwG8u2TkT3/d
mdTOKDBygZ8wnS1CWaRCeWprw2YnINjNfCpxFq26wxx+GuMznQwhlKNfwdqHE57pjJgJqgETBhl8
wIB1maYwOvvVyMvzEnwUF8kxn1kz825V+mXZpiLeB/2zAmbBsyI2LV5wxQqyQFXw4G8pLkRLHwIc
MlVuVkDq92d+hwbTYw4LuR5X1boiAUamhMaiwEagGNwSKQGNEZBkiW6gfcsbdwG/jgsY7sfVSwvO
7BO3KeooegghIb8rvrHJvampus0L3mzx2ggWumojOtqGaUjuPvx65nAnsudjrMEby+EV6hJDODqP
BWNsqvPEcOUV4CUfjdhTadFFps5vpwKHgYNcSiM8vo2JKBywwXly0U0aah/Clcj2tHZUQGRagHNR
K15a8XzPrEzFtx6FkhOdBrG9qFGpGNe5q5iEiqV00CbTSmLpdqCkh0mXIkRKUpEdnwaMWDcjI6xA
a9sC9iiM7nMcpa8NTlacNmIojvUxhO5iHGxA/hxXv4xnXfTH1PcHfjVI0H/Q04kH94c75W6doWPg
LLBKA7dMOvWpQls4LLI6XbN9NrLkcyxONywDpXjJqCPcWacQ/jZ3HUzs4Vrxxm+LIjbMU9xS55Rg
k+fwvfG2uy0XBHhQoixNXbAfQ4qnLYw/iVeeIKZvMqIBz8ZmpxXGsVVrai1mgC6al2/aWE4mAqVr
WXOsst+ulKe4xsQNrIcdVuSE3JdZTm8Q2zpjQbU8hAqpDo6N2Ob8Dx1p4ba4nu7I6iXKrWwb6M2H
gRNpbH/KxWQmD7fDwMlNNQEiaztG0hct/tdTp5+zSYE4Nj8Ua6VTbDdEEpBBg58dCutS+iel6qGh
CxH+wKemodjyhWTUk9Nk7TNcL5ft0/K8FRb6bCCYmyRP8rXtxOSFsUMx6iQ/7VD6cJcM2C+JbqMv
k8HsP4OV22KtNDBaEZR179PxNt++XdKQhFAJeTfOudxM/2R8SwEPZDkqbavvMJ+GO5/xD+nlDxSn
6wBTkjgMb+jTokMkJaZB/47V1N/aSTJ8OOJgrInYjPjv4z09koVawshhFX9pTmpOCxE/t/HPDjdZ
XijGo+vcym8g7TQOWNuwcEqMpK9mtilbO/9K5hvvz64XR3l9eVACZi8mocNe3mapETTS5adj+pZL
LkjIeJrqxbutJdDKxXzxSNgzLUEmS1h0pTT1Xu5xLF6t2W8bQrkPFGDYIy8s9J+XjAwDhJnTZtyw
yxFTUPz2zOZlosdOFPz5L2/wANl7pRJqK/BFmEDd9APoOXyjgXnRKK5k1yb+1MAXPlUkTL+VS93u
Twzkd/L80bODN2vbhOjOqjvllmKuBKfSlZDW2jvkfUf2b97yd+D7UIeq64//O0kEO4dbF7Yu75V/
cUAzXSkzZ4U6HhxMjNpt0DZTptEppz0ARmFA5YhcN/f4iZkFt2PZ2Omg5AowGW7fMgDfYsP71l/v
150BDjIT2SXkDEcGN7DBlzXcvxyIfeO0U7ZDY6xgDwlRciumJVAT5uRD/2JYSxc79oaREXXDGejE
v0kUx7uBRKJfRuOId5luysevA8TxtTCTF34tJyjUWS/LI3S5JJKgTwYAsRfwF3xySZFi5UIKLPl5
Gu7q6KoY73g19pFP2YIpqLZ9Mwkk5+OTuyJLRbr+6UO8W7RY+jDpSIFpe7xCxthRgM3obLzhGCoo
QazGnSoSLg6TdW7bTwVGyCgOP95BNiJKZDr8BBjKtQTicNJ/rrZq2+1LI80mYidl5e5PbnGL2B4B
tdxmse3j2OKKgQHuUN4zWj84Ea16IWtxj3H30QJh1+tfpXBSrVtDBxLwsfXfnI2kLkNOnZg6LeBO
f9x9JDTzNUeZTP4EcJkT4N4nD9ZZ0kDsALNK/R96VItfD806abWVCoZ5HY4wsRLR3yflN5dBncnH
hfiaVsehAdSQNDJZ5UemU2PMx0Dt8miIIjPucUlgtwZixgHBaMEwvR31n71e4JglDnd3pPzzksyP
euqS70I8uAVFeKv9jIglrTcX4hnW7QZB+i/NHdHWHk1JMWEVPI7adadZwzR1WR01HTBC2+ByZl7O
kGUW1JeplQFnjMAL/UXtqrRkmFboLJAWau+sSKFN8qj0MpWaFpO/mYvTKQwy3EMF8ktiQgqzPLLg
Tn4Uh1eUe8mT8M7VSbazkmF1AgPvVHX+SGoX6DrHWMm9y6maFg+IeBQ9wOM7UZ+R/OkVlA+b589W
pmDBLmiHlaXwSBKshFWkh7lKrjkI6SsZDeXWmITkoEXOQrHGk+IsT0tR51xP7KN9lcrHlTFQPqFw
Syv+g1ig9O3+yCJ2yRYMF9jeTjWbjx8i5ElUBU07SpX19sRvPF6a1lwAzLQ/OpWdJTZ4uotDeUzN
osfnZ8c5lIwt2zzGpHv60LUvDd1IXIaJNfh5SnTAVZYN+s1cFS+2KLHac6i0ycGuNXEPgxFVZ7YZ
+zf1cqF0zsT0kbAHQcxEt58T8mhlR8tN6lSVfsLjJYRbvop7hvdJ/6qtonfKYrf2iJgVrB5tp+V7
uPOufAEDW5AsVyoiKqKoF3HxIh1+drm95eQRloHxITUIgDrjRBVP1FCp1xevGBYAOVGkgDw8Pj4n
S3xDaNYgN4nXwk50b+waIUATMGGs2Fh+dCCPjdlFgfQSC+/ATqq5sK2nc2hRpOQRM7WjOjh69Q2A
vj68vrPNEXbx+vg8b17jjB8ktrB+/L6/qx2N5GEWowTburkYdYZfhi49NlAqgxgFVpt/4Y6QlIzA
hdTbW/QYGx2AmGUQa6DIZhWuhoTk5rKbh4nggoqksUEsUm405G5h+Flnpc37P3WamoukNpIbfRXF
OfTw1XwqpHvjVHkssq3qCTzUNazboWK+p5rIBo6ukE5HHJm3pGJu+IWVIwWzrfsV+wZwVS2amWEr
eU0n6Rjff43DMpfdyfzBqQK3uRO53EWx3tPzlh4WgPnJAFvzxmt6iO86bCDXnd1fxeUy/WA/lcWF
VYt8tVvfVG9DADf0K5QneQM2cEzXCtIbbVnRhjhUA4gULDF42lVHB6KoubYbKB6JnmVJQMVcaflm
aqrF6DXBYyOE0zS+8Ps1XTRgsQAZXzZ25+Lv+Te1xAf0pqwglSwhefkYOOi4+0R2kUaqc/ebDgHW
uszZGX4glt3i+be0ajkOl/hR2+sY+uXnQoimUvfD4+Nxxg/FK1xXk+ITfHRCNtZKadK/K+xFpGTK
toj6kOs3PBPD5/M7urUdTbTQ9TUBUF/gzI9I8BPlXUnm2vQw0z53dPm6vcHyntc7CVQyysuBd+Eh
YVvzD7lhPxE59ehGmoPmaFKL0dzcrjleVwNpRwYDVQBum97KKdVMXPmXeo99TV5M8VINmIS7ZLwS
Vck8Vo6m//biE9yeMEOPOxX7wt5lHnS5JToksuqTp9Q91aN+CPpJojcEe2o6iuoBNTieP+KWDPuS
cQ5z+4eL5UdKkkQg6pYaNJb3ey0N9gEZCTeQM4iDkxPGQfxUs8eIy1PR6C9nr/dNXFTX3NsUhiwz
HLTwhE3XVjUdF4dg/E0qXni3hAtj+RPzYQXHcE+nkFY9xffXAizVWkNx5ailT3cas8aDsL31Wa1f
rKza16l4UFBEOR8UKbvD8s6qVkuWtuw8HgtXCX1T4ukUbCWnD32JmKsqHTj1gN0XIPdD7CfY1bM4
intRqwFzNnk86JNwgPIrB/P8o57/cbI92amke5c/dxklpupvuYWgWt5dSPhG7/8Rdi6j7qhSfIH/
OgAmWv2/6M+xlldPQtwdRw2oW6ZE0e2RMeNd+CIRJmIZ+9rCJJpVoZyWlHMhCqkhdLL0LOsGF8Jr
Jt3vM6hkftIyalwZ2k3MMsSZQWuBv7tJjKtOvM6nOqTsDnzQka84S+6VIZxy47w/4QNMvHgbUNy6
TvBQU051xwbx6vQfZ3XP7uoaBkZ+/UKGuid7sZeUh8g6M1rFP4RhggAL617auylZyw9gaQYcrCRm
/kGp4HZxkOdYCxExtqmvUb15o2WRNBBNuAoonmC2zijrPHqPAKDYR/7gNn0A6Nxi4zH1JkxfwQNp
QjIvL/6EH/0HOke21Jn5wY1NXYbU4uSUfxq5/40elW2rEalodZd8J6AO9AJM11C8bA1iisiN/MYU
k5Z8aAc1oKv7ukg8mV3vg4yhqvvaHRDfHpgTdakePN/bC6B0LUn+N4lC0qJky/OllwtZxvYc4dAe
LARmUz6s9G8SFmAj8QOfWO33iXy+npkNzTob1YNehEp61V0tMu4e0VPEVcqkhD2BYFrSd2MZIDap
cjrtNUD6bQHLF2A4pHQU/fqhXaV2drpnCV84NJmq1CJOi16VpBpfUvhavYI9l16Za6VIaCRmJCso
nuvBB0C9I6/4Jnox8W2W96NBQkXj3xBtyyS4o3vKQqMDJEYrIRm+uwaZVmoxwKviAR1g9YOGJ1ha
Ub+DCr5MiG1rMLBOkF2iSpZoxImGxW81nHFlAE4or+2v99eZJSInWFgtD1rszn+ZrUtZKSHnYRG7
tPvi2s4/T94Cux+guY5vBpZuQ6qV/98dt7FfudV9qJm2g5NrZ05JPj3U79Uq0DoVASyStIoUqg9g
obnBh8u74nlIc8BvQXRP2MB4RnTowEj4NZhXazPn9KrTKQpRQCaWZyjXqsbPYfuj2RolD5TLk0c+
KIqflwtfq2DVhIYqfhQ2cVLyIp4OEBGONnBvlTBmgP+ZKzjazDnDeHQW8j2qU+dogndiz5IsDdtx
nu1Oy6c6U5FDxnK1OaUvNyyGw/DBaXhxYWqp2EsCJXPCv8Q/AIjURVHZWSqeiWUjIR0MUHwLXa2i
tNcMM24FInWL5hpZmS1BrpjDgfpjOjXnSTkVnabnQrEwPi4aH9cACOAcdIonuSwvpqyAZlmsFo5K
yiu6q7yiMhNTz1ecX/m5m7vhotxIMzFA+FbN9tBSLXrclXGds47OdN685TmvtYmHja/SMZkL29vS
4RIF559zNbgBXqV+hcuhLQwpC9/U4nfDc+vGdlEXfm4D1wlt66aiORIu3C3JpjbObc9scODELaYr
+IQZWjocz/Qr06NyfTYAEYEh5fa/inkH9tHxADzoiifvCvgTwS7fWD/hNusM/9gKGoMqkrv+l9+K
Co0TATZeWufp1s037cFTTyOGCdnxQvmn/tMHeO1f2zCBiC+QMrPL8SSXYmXIOnGS1CCgmNaOqMqj
jGpBMcycGEQewv7iVOUAG8wnLJ7bgagcVy9WLZB4x/zQkbDE15AX0W734+vnFi/niTbi0QMXQrpZ
QgXdb56PCyuBDkgLmXzOYYzUv1DPa2+8smsO9yNSX3YEtbyx3Qw5YgfHfHW4T2JyFh/7YUc3xeJp
ir7vY3Et5NMCdsP7jj2KbHdRgZqKI6ujdnZ9ZglNrNbo6qHLD1IqBcdbCmk9VpTqHoIgFkYYeWS/
6NYUVFvGWG4wFSXYnQPJTk+xjPNlM2+UqsGw2iDCaRRPN4xBlQuvCEP/Nyc7Ja0Vd5oQw6C7OoqG
WIg4z6DkWgJMlvZOAdqNynZfS0QM8fKb/gGrRbbyyd4G8URqtQbHepjgzHFFGpuuMHsNwIQDA5YJ
GLfEu2UBY9Lb0L/f5TcHAAKImicrhsiqh4w36OHyZPcAAJLzC4OlRsabUkkW/5S9m+krbsZyPAQ2
7IOfA8+Ad1sxeyHD9awV9Npjhwk1Cq9EriQQbO0kls2dtaE1mpmt9/uQe4DtXW7PpeeB0mSUGM64
XEObDTgSJOE8Ge7EvJmCVDqzxzPY4EpKfTAliZPdDNgSr0wh7Aw6ThXP+rJX2QZ4z6z25PIExC1N
vYaVpKJCBvOxF6dqTYIndc7bobvCs6bPf4ZEklESQ/MiQrBvQVmVHIFW5NP7L6CwWJI1r2s5H6V4
dcrF1Gn3MTUrfhUpkIAyjiAKt4iMVdgVV2nUtoPq3sGyQT6HNTygQCf8glhmWmrTthzoepao8zNd
eA+YIjZDyJoE5fg0aoxxgG39HpmAw0hw7ewcoK7E2GX2esLpELNb2hd9vmA6ruPiNaL/EJ7/CPKY
dEwF7q5j9Z4VQ9N2jKeH2cUG11qGpjc+53bJZdG9UGk5fqqzhJ1TxzpyeEYiV/jRCoedvg8rEQ9T
X09qWh/3pRgShqmgQM9+/B6EcWwWFDsGC1ZAP/mQIAVd3FITiKCYv05fnvfcnhEy05zIfvnvRatp
LWdcoKvWiBL2ZRG2IymqX7n3kseK82lhI1/LanjG3qxVqimNEkkAIfsvTTaTMZFZ83KKTgPIjTAT
HGVKt+QUp4CmC7CoVCp+txJLxFtZ7CeHgImxJ3EqnWicsB8jFcMI3o7uKyJLPEOey31vmefd3apQ
Lk5Dz7nFwt5VwbH/dHJ++26xnPVDNAA0fLUO4MdGOUP/eZj+QiKl+Z8NNEfASjJrSvkN/fMR8Dhl
ksa1aqUrLrOqNBTpE0vrLLK0V85OerTPjyqYvAJy/0QNY1oCPoOuk3uQq8epVl+Dd69IjQ19B7o6
fTFwI2VEHwPlxHe1WGxDizwS6sjAgQZgKHv2oPed24exGoq8DarFvupc0RA4IMTKYtv/LPI0pUT5
upn+sVQCHi5sD2OUyyttM8usc1Bb6KGf+NR9ljKDYXyIm4ttIccUeNgakYcJSk5NhSzZfal1LdCx
2T33DKG/4cey9zWdnegFIMJAuGmydDD00xNpeHolgxjWfgDZclEDtH9m7Od0l7REqZaFH60bVI/S
38b9seQ8grllrfUcWo8WJHlJuS6cosmY6wV18aUVzIqQ2QTxrG2h287zbnhRSG1w14OeuwiKfGuY
RYSLlpKlOmwwX1Gqwiv5seYGIhoTBDmf2IMbayxmklqmr2xiWmel8OXex4DRXbmk7CC0+Jc27ziB
Tl3RQyc31mIacC04jKWk4qQ0mUn8IQGHWzEFALCY35yqMueFbK2oKATdliUjRS095POUiNv+q9ng
4cWcnuwxRFDcVL68dbvn2CirUFNMf9uKzM0KCKMVvyVZ0IFXQiJzcoTGK/qvYi3xD7CMaGOWMh7x
3+8j9WlLf6yQUEfNEzoLFhggoGyZzonqLUQbelY6G+qiI/NDMaI7il1krsU7WdQc2D9ZqtszDWZC
TuMJPqYwxYb4oxZLRFNrYLvgM1ZuJxMKGzkIKauiG50tHOb6O4TgQ87yqTU/jxsfprd3oRtARGSy
oxJHF2E0D4fXuukk5hSf4U90GMlUQDpsjDIlW+hgDdeZEoexRTUgovhRz6mpKMoI5RGIorDLXS6q
jI1z/3JAa4D+FUhqGjUjSFEAUwSSOIdsvgLpQywher9rEl16suhtCq39+ph9Dh3bIPAaVtQOwRG7
CvxRsF07HQIYZkHsk6CqCKLDGTEs78t/U92xM2/MQgRgwiYwIEdwXXqK8ICmEeaQuUFNtNFv4nlp
6CucUbYTgm8SDLI7T5Tt911Nx5zSRDnXx7MTCef6r2UJHfcLcYdbscXSwdIp7BuMHjKtc3CxbjNC
hRuVWkKCAMKPmDzh75m2Cz9lC3ZIS1tpkTbo4D+b78YaJTEWA70pZKsPpG1sHXKjKkKyLz4sEUwS
lYbEcuKeQq34iClqR9XPxtCZSVDzIl4h30JFk4Coa2O3APK7KJ6M6fU04OAytnN9HHlOHIeyRMtW
9QdnpaYREm1Q4zE0W3xXqS+kTeVzB6ea1bmeLwZs56PIeXLyPgys8mlIeeMP87XhyBGNGPBdPj5E
2U+u491nvxEXLV3Fr6DOzDUCIDxHNCmt8sozF3FvOYbIERHyFCYzx1olnTZlITAOTCfjVe/goLbu
ZdMQ1mcWRWm69mZkVrGEri/fx2YEyCVuZMzn0PbyGi9RL0QqAG2T4zUmm2Zxp8tSKyvA8BoILzdT
zxH1vxI46UdnxEx5P8wCmPuu7lmg2BExvDV756OdARZE+ChSOlxiK0/RC2fGYD516F7NwCJZgmz8
g5aargSjsoqW2ZP4RXOQDmDtfEavc/o5Tx+ny9ZHokgOxiuhn/ebmOIZoHPvuqkDl7RTTN2OSZz5
E8c5o6R9a+aapiZ+yBoqXeAph1U2NJhYQuciQdDkLgDGD1flzzs6vO779hSIAmUdC6M7h6zWaUdL
xJ+Ubb95GrXZl+CmLVjquoLSg8y5YiYW11Xw0+tq61CYzoI0Afmf4lSr4jY93Y/pqR3kwEt2tP6b
/hebEgF9X9JHJDJJTSVB6JLzynXpGlba0WWRU/JVF27+QuJizI6plnUWV6HaNHEOBqSWalMNe/2M
PJuMEi0oH6XUHtR803loekO6ond2Lv8M95beZLmrsLnJ6qih/w3/eH+APvmr1BkJuSTEUKCiSf+0
oCa2Q/hXV7ebqFvhO51Mn9EatcmJlUBTX16/UPz7IQHUju1pZtJYuiL5mGmOkx0ReM3+8HrTR+mr
tp/EaEQ1z306XzLNn/uH7Jk0S8ya53VPjFzCHfVE6E85BdHBlUdaluH/AEjq5+vpgaYukkGC4RsP
8eLS+L+uCDen21Qu63+1F1h5skIFHZdqDHoSR0PuEdW69jePhfY0A4Oy1cpS5sNrmSp/iIP4hH9g
i8PmhpRY95zKs1Ugzr+qe7GEfQlOpPyGGUWC/PHOe43M0KwmNhdFKzjACEcWyNZAUr+BY2gV3QE7
cRvKXhPViODA4w375VFIIFuW0G7tzfy1K0A8d7Fyt6HU4UIbFWNz4PjzFdnjEzG4zQXuEWrVNMT/
pJWQEIvk7oNR0CevYDvcO5rcH4+mN24G3UqbaOr6qRclQK7NPpsjMsqUnIXsMe7tKeo58zKylrHi
G6zG1RRiajvhmGWIKFmpDCWdoMIg2crqmIX/vnHc85hLSAfHRipggXk/aA2p+8mAasc37H/99Dfl
CmdFgcaMRkzWJuzfYNNfeWIhahmFX05lNkjEnypF4tYufAiklAKNwd240vJe89KGyrXIxhSggEeT
s1ftEmABqAlUO1OxheQsMsW5oAYjiAYUIyJxrMjP6zIXlJPucPkDciNn5IT55lA2n24L443fyYAd
pA4T86WEMjqoIjKlvcnQBBoHVTERLX742ugvyY4DJ9ErNnQy25Dpfl1qiEgNHnsl5+SyYT4CiqBs
jUTI4M+MsWxy6j8EoQGhD6dUaRivSm5n5iYgzeNwnS2wWtYZHx2IfH7cRHnS680lf2bVhnyntM8A
H4V7zMQVySOh/4fhAiZrW7rP9c37u2/PIz/zSXFDTiE3TMdPpiEol11grM8A8dbomUmaW31Utcpo
U6FQtQVuRLMmyszOFpCMsyBKu768O1fVeYZYZPSb3ys7HkhunTveJsM5dB/MJgFC5yIdFRSCo+6b
ucj3lynn0JsfZq7D+U5KlqxQIPeJa9PN/jtB4WagRSTAb+r+Tr3arDN/NmQGI/Cg94KnfWbXmOfd
k6V8LA/uqWRaIKKmTf7kRBO4SH+zzCdmbCO6+ceoei5AjyAZHXj7+sGrNWGeqwaWVLlE4Ex2Enm0
I2K1rVnSvxPaGpn/qgWMkeC3BnQ1mJloZ2uT+EM0ahmStgLNFKBiboFF/zF0EgRBYdVFTRtkQRb5
85vvNFKFUo8aiuDY1+XJ8aZ/26w+on7fICTlJZ4G5fCF5v1cFVFQpoiiWTkPy1MoWyBUcusdcZD5
ac0ACfw5z+2erFvoryZtO7ojkldyGY6iVjbLCxmr7gpzCSRHbt59SDa9PWvoEfXXewC5le7ha4bE
74diTUoSQGbRI3q6SHMfgq1ZJNQvJXhxfTNNYFGsDb8724QTw8H1YU2ZXd2bigLIy23SD3E0bv6+
YGOCbreWdGce8tfjZBHzCCuoZZSiS4glURJWqIJSVeRIs/9R83p9Jfvc86415OCzd5YUN2Cjygao
cM8Mu3VsJJg7CRM0Il0T/eoGNAz/7xc1vwkAqI0ZGuJLGLpOquLDUzNXLZ/ZtJsHYAtzajpSRFw5
v0tIMKy10+KYtDu7kiGw/jYHe60cs3aOhB/4q0k0n102VEjYc1YVaFv1o0vs6Wkm06J4n68C7g77
XJPxNN0SvXw7Q7hza3OWyOQe9dMhtyKakbmQXwkA8FXkBLp4gfboch/9LktdvZmrF/VZJfM70ONk
a344jsu+hNS4lGGPOCRk+a468z5He/wqejb7RSHlZToohl3/vtb85tUTbM2Wv7iAgO6TBqno08q6
H+62OG9LZ0OKD6cP+0l6FJoJLTn8XlO/tOskF1Mxa40v90ZHuIyBEyDmLDsg/j5oG9IMLNyKAMUc
8ofeZh/VCdntZT/bBI4+/sdRWcXJGutxKgZqZg/nf6aUniX6TWKp9UWQrIrwmD6taqJ1OW4GvGbP
XcPOqq+RspJoVjayly38gomutBdTsws9kcBmKCX+2V/kyVIDiiyOh+MnXUlRZ6DZddJe+Q8TeILp
cm/ouYh64wJLaZEnSrLZtVOlrTtnaHwtrlgmrpry8Lisp4aa98L1ezr0r9MQj/mhQdLD1QHQQalO
eIHtswvruT43LvmxKzFW0UDX+49hsGFTyVZppL/JjcHVDQs3DiCIqm5q1TJXJRlblSS8GKZiDZJE
hNv6DLgCHHGshglvkKNbBTZHefb6KrTtG1cZhdvooyuaA+MgBxD3WmPPJwCFZBforv/hkztbL/o7
T3c8hTItRsSpYZGpRQ2WwaJxUHzSFTRNagBv6c6boI8hFebCfRAjMIDKZfyt8U58weu3x1gCh4+v
BaybsozYhhTrwSV2wZZo1zjhxTNlXjtOwOFwi54h5aUN1ESR5R5EkmiUOaeWSFX7fwRzcw3oautp
kSjgoUp+wglKO15aySBotkY+80cuTlgRASuOh/c0l1vv9SyIvpFz19NcWZFHVO4MeO62EoMdxXMw
WTk6/VkIYiTp/m7M2ufSTsShwCNVRgwBtWGPjZYIuK23xS+JJGt4QMjKxHqhJYbgazmzNVk6iU0K
a1n3d9XuNxja93jRPoF+eE4N2F6Zt4cSu54du2MW0fAGkUIbMK+PZ86hFb57uuZmzRIjNXJ27SNC
+fsSC91FSM3tadx65jao/o5ZK2deVtnZkUiJlaQQG1pfZMYg0zIJRe+SkO1iVi9o2KCKH1FewoPt
a+TtMHlCu0t18lpJkMVKFT7q2/9vs86TC4fueJax8W38Nf8tHRO0yi27rBSo/+nAOpRKqNGUV3dd
RD+GGBcwv2m0Ij3jAcymfYNolgZyczVYF55uF8kPhQwQrxKhDO/wD2iKKZF7mnNiMtj+yx8T9pVb
xdPj4l0zgQaJ1Qs1NKL75DlFD417G7m3U1bnhpp3PHmiIcFI6jf07gLM0ngV6v8J0V36UAa1nls/
qB8Tc3mlBK62f4gM+ICKP9XXl2MGASfE8PAqchDlI5vcOnbq6jYkWd3xJXq//B16su20ACa5IXzy
+mBMwNbCmbJYz2naeTbcp6PrmhfKMxicF4ksvo/3VkImGL4fscEbQxrahGRncfDVhB93u3rwOahz
2+eISWdquJQPdb7NbMplFDozVspCKvk5On5e5QPZHXnc/KrJBgKzCWO8cB2fJF+PCSoyayafJLEx
9BoCBmtzehkke7CmRFUe6XqXmBvOpQT88VakW3KHo6WcAjAppoh6tjPRcu0IOsUrpN/JGFSUTGWD
tT/1WfaMlh2z8977ZuTH/Lh3FpWcymj37N5J3AguYfS2he3QtQ2JPiTaftdXzti+OSe3lfFOPXxY
3oSlQfnxxF+HMOD12Lrndk5lvUhTcpzBw5nK/i3SbYg4uftncmWoYRdVVlEezFkB76AUd/OBQisa
hUIbOUgG6etd9ENSFWd7XpUap/m0jrFVRczQ9RUrbB12IhOwV6QwK3Md4sQPYhLaS6CK5DPs5Apc
SZpO25IDVjjyVan3Sdb9247KpWv5VwEr5xqArSh0cuejiqvteGU5JSQY0mk/lon/YN6jiWxZK2HC
Q4hHPUbgBobBmpkV4kU/lwnzcUUnpgRWf3dIFTzpc0kb/NaRuA8nyrYbAGXWotdUs9hOmYFhH46V
76SZgNa9lSxUePtu11pICmxpebV2IdCXoecX8kWhROHJKlpWXEaEj2xYW58w281+27eNVJ90mQrX
sI5U/PGCR+0MVnJLvm4braQgJ9ED35FXFF7zzRJlolhKpKrZ+yxMW75s8127gWCl7AeLkRWW6B5v
9RHlo4BUGIhkLYw4CouKqrS9j+Jmtwrgw9wop11tECxCxohEJHJyeRXyNxviuozxJDDpIobz1ct3
oab8vSHB6D68WlYT8XdmLtred4q5uF1wM3uWTaAlYkyywdTofc8NSzbnfu5gLIvtZkuj2rLZpsBf
aVWZuEeGqxdCsiABFPQDXC2WpwG3oXbMuN8pu24sUmq60WeuuHgyaOSGXC1+oetqjY6+mvl2geQq
UiRNDiLydfVGWyjEA9NP8FRDVpOBPI4PgoFN7qv0SuDsKcjO2hss8V+rLGMZyinSz3ruQwK3UOkW
MUj5bGeUCDVqli7M2nBHVhw/x++AfbtROch8oikwcYgoqsS+Y8/xN8QuzN7oyX187wxm6jX3IFSE
OeG7rtSQue2s29fV/QTQprIFLEHOqy+xmyLrnfT+ElntDsYHN9+61loNGMhajoZL+wjvKNknreHO
04UoP2QJ7K+/A3ztzbIba4NjPC2N4di3QP2Pbx74vCwhmXiQjWd63bsbG5hCmI5ZHCSqmv9XcQ4A
+j2fMzHxy1Iv/7tfF67m38xHAgyT4WTfycosLE/t5DFDIhltv97Skq4JecdGynSzEeCOUcqWc4lM
+a8qPJURZmx80pMJzeVlgfPj+d3NMiFEhiyWMEK966VDfUddfveXSFl/MqKnD0TWNtoY7Nhm48jL
9y/0lJWePrjFlCc8jIhuEIFOXmqIjONTo7AWdOFrnPyE+A+2VE0jAaUtzUu75AZX5GolxmTklIeT
vWgyAhiQQwvcjmmS8EDBKKNE4sJIiur+fS5TndI/6sPo1RPUakLQQkPP2XXbOZAszvHEFLdViBc2
6qDMlvHzjCwTATEWcsU8te8whCuVRQM3Lc1Rm8zKPqqXxSEowv0k2h4SJrkVA9Je8/2S4j5FXNBy
9y+tWH1ErdngvNnwI6OuYf29D54nS3+2gZr343Ny5w2mXHi+NI0z8/lQXhl1ZePyjMVKvn6H+JMH
EGF9FZKTtZIJJItUp8GpOcmtE9sS8rEzyF1+e2pkN0SpLTUIBrdJYZUZ4/tiPbhCVVBUsulahXAJ
m+9MZl+Cca2a6UCMqxOw6J+46X8HHe1xNeV+9iRfICAJlBCSL1f4cEPgLPzK3kC6T5B0aQnLX05u
W4qUWh2x1xpp9EGPtr4PtABVTXqryHdOzKiYI72VZuGKpjNcSULdMnRi3XxdSQvSIb6tiia1UgHH
bTq10/7x43wfnSqZrEBoWlxQUbW1DfEDRQvkMWJa5RxW+slIv7GiqGeL5dy8CrzBO+gYbTSz4jUc
RT1SwMrq/dejbnGhu8wZoqx6FzVvwJdmIEsHjymCenJlFAvuqY1x8ifg/IAGAeMODlgt6B5/FdQP
Vx+wRtV9WqcnGUDpVPs/75QO/SVqGfVQCs521xTwbkhb4N/eVU3wz1wnY/syhhwX7xa+G5+JacVs
W+iDafSPHLp3Uhybw49QPjJP1emv+8+MCwyTxjLNTLFDEeaNovo7O0EFLDyXkWptUiO9gdDC4rvO
hZwAHMYWNXH5ZmmMXqrwWKglAJFvWZ7MorDNnzr8GqUUfx5yAXwz5IMpvMQTkxgd2kwGDDyXpcHd
JfF/aOpyzqc4PT58PbhFjPvQpee+U+G8la/gQFSbVqPkwj6VSjTikBCf6oMCD5mrmXbyCQptLXOh
YgdFiBzFcDe6EFhg7PpkM+Hfj+GMKHLjhqxSgnH7O4ViSJLvXFuaGkc99KTdTFIaEUGW+j6HT+uj
451xa6E5ElXAj2Jh1ZaP56RRh4pJpEpY8m+ra4eGqESG0eB4iuOqhWZajAiJ64r8mYdcZFPAb9e6
yzG94yRqKKiFt6m3mcjBud1syXoO2j+aMEUDE9yCFdbJClNA1JWfwHXDb7SRKutrA7fAgc/8vbBa
I9dMuAt5/GXsfmwtyPxqiE7aon+ty5vokS38gx4wxXjNdfGxyDwqAOXqARu6dNUcIizK8xT4LFT1
6yD9/xC37Busr1axsO53v3IdB+d69Snj5O8o1WjALaGSkO6Acx8uePPPJITDIdGTEQ2S7U3eqhYh
aInS9SbWrJ0AokMn+9f6G/S9hxR31CJ27SW8J5XQpUo8+EdQjIhESlnTd68LmsOM68Lf1j6StPut
RQEUPaaikvw9l07H2RX1su3zBE1Uj+J9K7BSydLa2wCOm5xyB2fPW6g3ewrTwdMxxX9zAhyM0l/J
PIDTdSYFH9fV6suBdj/CgOIDp4CbvT44BLYJ3Oo+YM5VlyrYEG74fufrYDtGw8S9nIbPFqSO29Y/
z7/UeRA6GYsTw1HjBIJk1eHNtYyNABmhqQE5xfyVnjkdcvK2bjPHDMqTV9RmSexORpXIxUVE1QwV
O6/QBs4IBZ9MDd6JXTBt9MeW1M+VZD38cOnyECxbmOwnqvyYru4RHdYTADmVYxivRP9t/qJIE5Ur
eVK3rjMOi/hZd8GHb++sXCMvJf2QJK8TScq0b1rzTynMR2lwd9PBhi3sPkx+haIRGEP1xYKuuyzK
HntXxzKH5AQhjcu8tHJCs4MlA8P3PH8jeiV4lgRuwttXqIoj+eXA1I7LiT9b2gGwrSmylfs6oNdU
pWnK1V9dwf9qXiUfE+xkiLjIfa8Hk23zE9lCRbe5D4Tabxjjx+tm77ignN6LJ4kpg0r7e4LRrugb
LB2Sygz6DGsNZ4sCn1K3tWWoRG8d4tw7Pv2VFkeuVbB2eHFGpabjcEFSuxUqMySLbcB78Ch72M4/
MWJbnjRAn0R9NfJ0MMy3ZWNXo2TwoH3AH/0n/p1pj16KLP2/yMGGcrsawO6vt6bV6hCY3uutisbJ
eAMlvuBgyrWhqI7Izd7bM5yKRkMFSCSQ3l+/TyF2nK5GL+slGh8ZwJmtJKcDMegV6xYOICmcJtkB
mSW6Loc9EheM4XKOxZHe6M0EEfSwljTfygWX8KDmMn/8i4+0GuaVHVAE/wOk6JEEJCn3B2PU55iO
MDdp6Wxr9rLaG5pwQGIMeAwxgvapj20DMjUwzG/az9yjj5uCo7Jo/A9EFkZCTFXvDTAkbv/RhQfI
gFkwTkktOad6kM1hfgqVfDLxGL/XsIiTKAs88e1JSnGGE5h1VnXg6jd6KUaz0IQTsOu6lw7opcFy
EK5gmRrPWYkUoCdkacuvo6poJWOohbmAW+6QIKKjAe134DLoazRLTgmBXgHHn42WUnAjUxy/3Eda
nD+kS03BZdaJLMrYATIlM58qiUZMZ2Qgq5TG9Vv/uHM6IVZlm9CukU7xRhge//9j8DFySNLIBSC+
sDrjeROh8OBL/gl/wgVoaHcUpepiLTV6/90sfmEFbz2dgJiifoFo8/3fStkCRHMjgSSdYN3eAgIC
Z46MO8688sJzAa4HgsuxFCQVSb+BAB3++NNXIZ1AALn9lLAVhj1oVR8lCSndQ21127rfkWu6cDt+
Zvrr15yFA8aXLT0WjMGRQR0QRPv2Ew+BfwvoCMYkHIYb7ngapevyqSnz6NpJLMvgCqgCOvGg6eJi
kGRnEtD9BOsso1YUgFFLBpv3L7GL/YOzcAKOmhbNm9O7f6tlbfP85mk1fVE9qFGaPPRfH+o8+kRy
T1B9D9Yw5H4QmhbVnZiIwaeNnwA3UXwOYpRFqeKuPxUV7e8cfPhYn7fQlkjblSV09TLuII9G2dgy
PaslA4zsZIu3R8wDT4Ln1E0JxfXY3Bidxg6rA5+dDBvdmGbTV/zJhrHivEtneO2RtVYHEErP/ipc
Ou/cYxB3r4EzggzU0cHpu075cxqBLJA+KjVSR/wTVsEKMBhs+dKlcNUPXQtU9Fn4lasqzHytXtiN
w28R5Qw5rgpBY89NaRutqx/NkHGdloyNUXggIdYY7h4Y6RGm5DYHsCuOKpIJd0SwwyrajBE+0hHK
tv60snlUNd9Ul3kwXA9fD7v9fKS+dF+dJ2+DVWdjdQ5yXWLSDNcdxCdqiaguDtkxwIhSYsVLao5E
puk46NfVoKavlja23f3Gvrie1G26y3PK6px1lsrsw8e64b7eqdGaCGneQ76D+hoWlDp+da3nYq1J
DDZk8pwjNGvfF3bi2fAbm/lpL1vkmr5XVc0QgBp3ocOrisvh86UX5+6jJznZTh5MmVHwoyb6Rowa
kUROhZDj7Vvf5oFXma63/rEruS5V9ZHn4kEOXyLYu8pW62RzzuYoYVQqHO1NRhBFuL9LZYeXi6qo
6oT1I5P+fyKYKnGPl5oENxKrKgekRICKL+2Z++WEfVKhin/3QB82C+1RYnaSB5WVmm9qP22hWiye
W8oO8ICKnKIe6ae/dQvx1MXOFxzyVTMH3L438PLEmmH0Cl+LBJrbmDYAi1ENsVXUHL1wNxJNeg4f
4vluF6D9lvLHauEcw5Qkh51tD+ignJ01x/oClJ9BRakyG0B5GNmo8HKkHorEylLmI8IkW0T6Crwu
y1f5/2p6pnBVoP85edwZq52bPsSjHxMvomINCRtUmjgYafBMf3SkFGUwzpF7phEZBVAsLa7NoZYJ
Sex3IcNt6EcZUL8I4nzA8pjVCisojU5CEbmT3EDOwAdN5C9dgMWKu/5MRsvMW8sR7fKNOmllyDV5
owTLldmSdcenCZu+e6z6YsRBx3MV7mqr0eGotCXIcWf9SOVJCTQg7ylUhzPtAsuWocIxbLeMVEv7
ipqSHddC7Mnazqgkn49c6/KiFLfZ3OAo5rCIc6hDb3l3N81+iUR41pm/fXeexhkopOvW1yeMy0SB
ek+Iz0yAceokz9S4vy43V6pvP3jisI+uUfq5jOH/aV7Id/9HEPCyKU5D7JQeDMXuvEXic7whXCCg
seb6HToAR53i0k1Kj+ecgICVGE/K7iFpu+JihTczHS3DN3MsSdOVneLap/FHop8kLqTIDfskYtUZ
V2wizHvlpBoAT2u0uIh63/KdxhwB8q/ydBchT+21vMECPlhcbn8olRDLlZ/qu+n/7xIN1xr+ExLH
oD5On8pQVVp1QBua/Dzyyhkge4R+iVkMngVjagbmg5BbeOm7Mqr7fAdNtq11WcaSMgo5bSgcQnMc
bAbSAS2vQuswbnYL1Hg27EvDj86TRBm7ErraVeZX7z3GbXYYwMsa/xDz1pIf1ajvRwyi8DpAq9yM
CiSnx7BgQ7yoV2mThOS81NjRdcLQy/mnxck+rN/WP/T16WoJSTYNhvmlepDS8Pde6EuO1ie7Kv0l
pzUFVfqi4d8cbclo9WziV/4Hqh7QSJi7rNNrOAq+MfSXmdPdjUiVCbSUOwv6y0kkfseSIuZOinxy
XvhCFBsmbZDbOR8x+wVFLy1i42188a8aBgRULvohH5SAWZdg4jd5tXUM55EVoY3coR49sp9XxqZS
sHj5T58DDbh7+7eZLBVVCvZhrt4pMp5ww9ZKGEVvsXSkFmgngS31hbsFLHTLenL+iBKiKfSdC1WP
ecjUj0rwFfsoxZR8RTVQbzE3q9PaJoJrBE+59jgC9Ncx4iG14XeEJ+Hd+05H7F+R9/8Utc1aGpvJ
djceyPKakVMxSaj/xXRF+qBnfc8x4cqKupcAQs0wlG/efW41HTTzMoJMpyjDouDZ9f8Bso/Zo3i6
oMl5Kri59LRv5yvLhVM7MfAOv+NJxlqi/yDWcHa45MQZcvbKI9zK4n5wkSbegfYcdtIT9ZWVBRz8
BjRZEhWrS5jHLSJN9BPlop5dayZs7ASH0ahq37fYJIie9gh/l7mapNrTCSlE9rr7rEPLudxBp8dy
2T7t2LHFpXVd6xPJWcwI4bJvYVf41k1DxCeQYmdOeHDmqy6vN+x58+dxvdCiV0nuYqP4JvVoU14/
gJudilBLqEHG3oa0Jkq8MOjPtF2MScpm0JmGd3vLN+VQpywUl3XuWju35A3pTEjsrhC1Ib4wzXAv
sTywnQwosvJ5kvkON8KCPvoZkWs5GMpcy5V9sLKG0QINhSV2NQpC3QpbLoLxboIRMKlBNWwFD0iR
I1MToF4aBnXFQlfsMi47hwWBy/R7cJJjDn0qvpK/9iz2n849VmUfE3kc7hCZ8Eh6G0Jvze8khs1B
N+zrZ21g1jFrHDuX/JynRdJScZVvAPHBjQezjvdxLk8Nxe5fRouyzWvaIUrFwU19+8R1dVeRQCoR
bVTS6rgKa5ytfojdLbp7J6V26eogzgX91/f5WIP2B6Ibj8vn6vbeS/bQw0HmwCgnSBFlPWp6Zqk7
/vurHAGJbz2an3P6bALAS1Vb2va7QX4ErApfRHx08Kk4vUMoGRswnQLPKsBZS4PKoHzlfA5ZSSTz
xPt5ZeXzwbBfFPgBZnGAkHiIlhzwIOccQLHgB7tMCGuJ/47ITZKZNb834AIeupQFTXH8hy28DK8i
14Z+K1JIaEZ8zQjhWy/egujfHppxoeoExVo+P2IDa5nZfLwJN+VnR7BiuTSuR/AzS4clI193emEX
L29serSv/kZ4vTq2DwbrW9qQ41fBfE5Rjku/uiFaoIlZ67RalJcmp6s+7xVnDF/XorFCxKkmzT2i
oNIj1h5OOgorqMVm4HCQUIFVmzuH3fuuC8pcs2f/esk+g46FTe5//jTmuWj8/imHqe+YCYyBTKxm
PoALbRkSp5uaG6O1wIyi2y3uCVmaBqQOZuDMbweJMbAtY7QKkuNNVycwod1IHO0J3AQn4MgduEXf
Bp6qhpycebiznBuq9dxem++nc9l0DMCSG7/1TmExtiLIE5Fl8dmHoc5L3uQeai1EU+w9hlUTWsAz
X6MW1vENWjvtx04FuuGuZej7XbGxN7PfqkmYsHoz17nMqWVaPDLR7EqYbSbOQaffTSDAZmVCMJYI
T3zD/xvyoRhS8R/FQJYRq25PjhvoXLKESMj6iipk8s2buBhZPEVH1SVVbDhyhuWzLJp7qu/Dvt6m
iGRa5kHSiYiBvCDCDP+mdeomTM7vm0FHmDOTpxgl+2wUs259q/E+jHVw5fXdNtEkHVCiy84UUyX7
d08d9wPHksb2MjbGGxAfV50i0pJ1wXwXOR1m9yqnVIhnCMFIRTfwAR/sKKpOUXW4ofFk/WI9+bCa
wjr/cqGsIke6IlhKBV1TaGaOTuT9PQj6H7+6zQW5ZrmKCPjghyO5CwNkGoj9dYwJ8d+X5KyfQfep
izl1qWsal6tQCUw0IUa02qKRr9MJAhYsAb/hEcW9dec9F88CrSK5DuF/FNHmS6tU0xb+Kx5Wngzn
3QZCsiJUNuAJ+5pcZVZIvJzaVo+Lard+pTdb09XDtQWNMmJIwJHzBICGLfDmmfX1aFyKtmG+uxvF
q9OJE+5wRgmdCkOHcNbl05zc/y4H3+P+coY8FBDUY8Y4lT4k4R+FAfPVySeXBSx2kM+UX6CyETzj
xw3rK3EFct5/ZQNsa+C7LHi/9Wq7GmR2kAe92m2QRzcaI58az6cgQ/dw9v//WI6yZ52r7Oo0MgUu
lmPMKjpxGrF0PLlOdnhwG9vSti5Sq5Jxb3mFHNhTeFpHLiG9brk0WFqzVOfCWuruCsQ/2q+vqqv+
90Q2iCaOGGg6IWZs7Zxgr54ZUatun5WHI6sJ7b8Sxb/gFsurZRFZV+9Y6lBQSs6BbdygxYrxLd3z
PnJCATDJKwvkUhem5kFqITW8O9mWaYDe6XgmHf1ZTG+xe3uG+l2uIokiaXxTvN/U6VGpuYfVIurG
p908dvh7RequjPDbQ0iKHZabBrmk746DLnOnXv5eUIO4uDXIr6/pXiXgAiw8Ii7hpDa41vZEptda
4G75qlJBchL7zQTcyhW6XN7MBmoLJpqg+iCnZGv08429Smh6r4d2VWLX4q54Lm4ZepZdDEZfUOvr
wkHSB6iKcVSoiN2zvaW3sN5WqABN4Eh3yNP9w9tDx8woxvnPQNWD2i+6kNoD3bwhqVzvlfdFd+XA
p10ZomlEvQUjx/SqXIuEAt40dJQdWZzSmtg6HeGCk7prxXRIad9LlK8ovdgjowmpwC2hpHfW8FE0
Q1NHqTsc8SyZyG2M9qjdfhFbeGejhbdyKcsgAwvQ2i0VU8ywTO58BQfO3nTYuK06Gf8bhaanf7O0
AhxxU9nPqiNvHqiCNt135zF2SNaMURvjrUO+N8WZy+ZAOjpKNxFftv7GWNocicDt6YvHYDDcxrFg
jLwWKdLWY9I3GLBS9A+qXvLYz6C6RmJdturyrCLeUc05XbZklN8+sPi7ynNm8j+d0vg4F82hPvqD
XJw7bZRc6UJTqHJpnShvOPqU4OZK5T10k3C6k5Zalch6rDi29O8g5fDx3TIorVqFdRsFCa6IEVoD
+C2GAFq0cabgcHHab1d/6wa/isDyOGobMjXaNeINN+2UKO/WQWueOdGWHEUQEUeQi5YafbaKXe7U
OynaexUBK14+lWJUxxBZZDmIvffcqZcHCz64zXB9N8GBJIQCK0xGj9YXFKFgmu/GHVZSPexIbndV
rQ1X0EMk6TK2mBZn+EQLBLExzaf0SxpdolNQcj4enkhkcpD2egxHMtzG7JZuPvPqoU1TOiayUvU0
1C4HuRm2D3WGeFjjLegqyA6eEyQqHveZh/IAFhOgGxUXWp2qxEisyR4YfkTClY2x9X+c7SdHg6s0
KgtGf7c1OMz90x4AB5VfDsLWluSb5e1eORIKHtj58fio19GxJ/UhPXnsV7dYyLe5Ws48P3R8ntSX
OpNFWb2DliA2nggUQgMO9GKuHxcPNZ7Za7RncnCg1QdmkO4Aj0nIXHE5ghcoX1KbduCykkPE7WPx
6h7Ipg4O+egQai2jEohoNg1Apn4Ns7kbfAs5aEyWyt2sBuwcLPiC2fuqI8V/sGDhXmZ8mgfTKXNj
7GZyyIEhsWCG/O2adcBaUqZ7mMapowx40N/mPq0fwq1093Xqab1B9zft6X/rZsF+4UFrKQhhf+HF
JbX80SOoqfMDVzrXkzsY8QxUnum1JUrcCAj0GfhLps98zNBJ6RX7+CIQvoE8GyPayUo53d1X6QqE
EG2wi6aow5esuqqEMg4gLfg4iqF8pQ/4QMbXQLgsVhx447rmdvGhctJ8dTZN205L/em0FqLsp3SA
6bABfV3LcpXbnTO15e5My9m1aWdflrlYvYE7GqUNcv/8wsFxN5k4f/8JgZh8RUbnTe9nM0RfmpCh
sKWbC8pwh3OlZqKBHRiEvuo9rzQCDerDItD0Bx81aEK28igveg5PZFJph7bfHDTus1A5i8WBXPKn
6OxAkn3Ud1X/OWPL5iImEAbE+15M1H5PqdO4yyK6yitW7SNbl8ws8VjFMrmFFp0Ud6F8zSAYvCAS
be2oxIkqj3mradPMxp7RnRsZC2V/hzqjamiGhikJHParYCvo1VczB74YGH/7m0KiE0s4caQMILNw
n1gBkuB9077f1NmvUdPa5dT8Qnpbsh6zaJcnA6gC1e2Yq2iuntjQTgd4g4Nr1MFJStBeF7WtD35i
/+0V2YjDwhwy9Sl3CQNdyl09IZLCQxwZZSlXfDLQPxeVTSNPjC2WuPv27zBwBHMHGpydWnKweVXk
2NgObZcQy/uDgsl7PJvj5+/SAyOTZKUve6u8SY+G+skQDUaPJPqf5iFBHlfYwU8tEHiEhBWshQWC
i9cAfGMyQJ6gBuYhVYdqwHXpI7NY7wpABRtZYKfeaUFkrLx+8045LQo0BPlorb+uvFOia3WY+Zlo
8APAA64MR1myX5AflQixPjuVpXSbYmHF/kWcDlAjNJE5vJFyDKkHHD7Zx7BojLQLTwRF4mBXRHbN
/GyWvs7KIbcR2N2yavfac/mIyFcVbpiYZ8lXdRE1hgcDWr0u5Elv0bLipCO811AnoYdlyUA0yzyD
kdxL07dOqb+dsRQ+C+Zgxxqwn3hs8L7hXPuIgAsQdZl98lAhDhMILYN0s3zj25Vflsl1XIRKsL49
PCT3OH4hQTZMv5qqWrXt/3pjh0ltj00jbsg1XndpgMX8RX1/fEKdyK2J0dqWJGlaWhpnYTEVJ1ff
FyFytYvYm2xRIe84q1lQmX/UG/NI2dIY40NNv2YAuCBQmqZo40pSitoD0ajn7LS+LDc88GUsMInc
Ylg+PbJ+aFDzcPrD7jbFRuFEhOIxoVjGgCgtFEFe845+UxBLF3Rx1wKQ94iOUz6/hrjZoXOdFuAK
1zdJ853Bkn3j7dxMVJC0lMm7sQXqlw8Eth+pZZ0myJWK/qN4ocSJyeqJp8X7/+kxEn2a7U346me9
XK3TCnFyb6kPbjwn3lRhx2F6vi4ORz/Ug+OVIVpQGUiCMrKgEMxKuDTNy6oOejsDH5uvipwiFvXP
f8ReZknN/eFWSPiVFSgoL3G8KzUpO7jqOnjU/AJV3bxnmZ7kPjqTTu0QZh5LErhP19pOr5fgwkZj
GG0OFdA6Qwu2dT3S10V4JgJp7J2paJ/oifCJSIfNBuKsAILbJ//Yhcdu0NbRtL6zX+zz5lD4wpZH
GZXgmRwwqcyfa/MrT2pXPVqcIkrupu6LYCqiX+UhkZsN19yK3cUtSYlopXmiTwszf35b0xo3eqok
DPPkjGMBZ/YKZ+/S//wDC2RZ8iCK8hrRCstYLj1MqeEECqCRJ2JT5Wnqw3F1nq9dC0bV3CKkrHfI
jgRd1ReaJHu6crb2slE04JpbOv/NLzcEAQG1pNWYwX2cf+jTTYCBZRXs347bVkej6tB9Zlxk8xN6
Brh/rheOml8ZciaFI5SlRY6q7sG3ekBAPEtn5XWBC8pBP77bN7zRZEEY8uHp2xtURlSG7DoZWz2h
g2del4SwxufAsKyA/pFaSKrmja/qHlFeN+DLGXS6Aw4x8/y5AzFkOJsTBmFwjcqIDOhFi3mwtMJv
9Ca/VpGHr7RCju66MDUGRKH4Rwt4Wpb0ytwMpfW16UWQQn6rVC+zYu+52Czs1ANB9Yl0eKVca3fa
NQo7tBisnoykYY2xDevk/YzXXANGaXkjY/H0xGVFiyXgo70PTB4a0d9Zh+Pf/DbcDNtpHjMDhG9w
s8emGDNnAygsouRzQD/AkA7evNzvvdOovvxLbsmP+yA+07N4I2BOxqcBc4BFJJEEC+uLUGj2a7WL
pG0VRv3/Ex6NByMyITBnpO/voC8ZqyDVTrwrOxBzWef3NARDyPE+9vGPqUYQ6FDo1GrjlA6H62EA
55hiPt6s4qOmTYWzURu0lOAc4r9a2pHXn07CHObO0d6JeG3DgvdNHW7/xMO6DKezEx5krZ6dx61E
WkaU4YwaAIt577j4kbhljbPtqucsTpj7PA4DB/qbyu1wIeYcBPqjPhaVXyzmg0kfF0sGHOXqgAuv
GWo0hNIamJ01LyHlw3YIzx0IoQDd0bOEzh+KI6PhOAr9coVzYlHCp7taJn9BRyIS8d2UvzqCrYSH
bReCzVO85hSH4QPWBGfMpTuzf+YdudkBRjRc55EmARhuR4Z7TCYnftxv4KqhNIRxR78INqwftJjo
gP+koPzLbnxSWJZGRw2SsXVQlRqpAjt4UszxJKMMm+cBTrUjs/N2lw88nAAMXBpk9naxzkUAvVvW
S5R3WWxYaQyPyV6mOutAleBuJy7yq6ISSVaCOdWDccJuXl+gRyaRT9ottfGB96hB+CBGDsnW54IY
tgYO5438J5sCdpnGK6PdEs499aV4soLDAramoT0c3sHyFqmGyqBUD+UV0H85E9RnM3JPWP9Wnfwh
OiRUwDDyHlB22QDhHoY6ijE13A7PE09E9VRVJeuO0x82ruVis+DVDfjRE2IzMBVWPfpCcGHHzMDK
Rta6APOJslR+otcIm4MMOLg9ey3YFg1ZMb7YMWyZdog7ruaEffE294LPUf8jwXSMOUWn9yc68p9W
MXe+7ZA+SCyj7M37b6HJa5/z1e8c+gZbOXrRNjWr46YfNBetPRe0VM+hc3/2hB5u9sE4RehKd/qq
NfDV7e3w6SvT296AxWFml/TFG3y7U22L/gAwNGl2Cha3vLCvBlOw3wuhM/4zDdo5xlmQA6GY589G
8Xn6s17mjyXhMuOrC0uFREZ9uYrRqWSZSwQgQYn+w1vDRFAICqoHoOybHKlWarW9GHvf0TXxlgjy
4qpN1GB0gq+L5dRjBSTq3A9/Y7VkHhh39mmVQo4wSiJQ3xSVF+g6QafOlhEs+Vf/N0rx8aaPkxBH
YJl0w+qSdIk0tvROkQDWlhOoDh6xw3AYrJMPVZcIeWY+6GYZk/dCxV8lhWX1ot3tyg02M5+NyhBB
vC/+9oHZdv+SJJLzz/qk2ABzqhuDk8cC4gpFNW3790VBHymnTFA4GtH8yHNINaQfm7CCcjoxSy4h
CPkRc4Bne2qcBRtXLja7XYeNQaCkG+yBnvY+1J1az121Zzl7rgO/RUh1e0a3zN0FWYfE6tjjf/N1
Odxdm0NHd7+LVGDCNMQO0Gok0bcBBYXwuKiJJVDbYKxZH7b8Vy08bWAclC+zYc//IaVOoyQvtzEG
BBfi4lKJ4ryCswCuNHJMbF8c0VSlfE9+JkFGMLswJbsC7DUhdzL0WJG28uvQYd/bPRR4BNAgR7VA
qt2GTJ3axuZnaZZAlIEGfLwG7mc+yIN44jnk90axwXsa6WxtGwfIk7YXYLNCJ24SvUpKDA3q52mV
W3UDB7KXiMZNRvJBHfDLknaqeVScyZPzV7jpxgbPTV2PExXi4tTUNbZAoMEeEaiq/Bu9v+zZeNQg
oS0gg6o5VIV9fSOCtLbro+hCbvKKC0Me4TqpDPS/Gu0p2r0IhbUV79IbXhRztIFbMR04Rf6FsM1q
+kk5VCwRwf7T7aHlg7lrDPhtlZRJX0sFocVu3/GdTT8zwFKx+TzhHcgKbk+I8dJIfkQ8NLRBN15R
vm42Id7dhBE8P46+8HPsLep/yeztACwQ8h+HvpYoEa7qfMFvaC5vv7ARindsZi9eadjAQBsVzqFN
65dc67+Re85p/qhyUrFdwSkBa3TLTpdREtxWLaObOsWkIQGR2m4rck6wEQZfM+MThzlIR+REaDO2
YCva+CgbBKHzfIWMjNciWa4gwZM3loq3L2XWJAYMyk8QrNTeP+zzoRcSCNSofshySXMYPbRaX5jT
xP93x3XD2mlYJz9jFDBnl0ZT1NO5NIvfYjoPli8ZOHpfATI5gJOQku+YptXylef+wPOAKsQCFPxr
Ws1Bpg7HWfa/4LGz6bX7HgD6nrUEA63qDessEdIRy5JklKCFOrHKqR5+98umsIvqU0TjhziUJs5X
vMjOS/p3fwuSfl5vjq6Oij8uvZZMXizWOupw89rJH7zXzk0ehtZmtrTDinUOnFNnV78JHcLoHTTX
jPW2pFaC7KBOsgD4aaJYjs0lOTLFlhdO8gDt2lDCi86qWR8VtbOFRrVYgF1TYdDuw3EEYs2amt/3
48qCOGkTFBXryzFPk7aHb6OYAyzKEqrx17/CJISPeCRjLQ1cIKvHqI4CmjsOYImdsNAFy3hw6V7d
qGvI7qt81daOa3/kTBNnYDXQR2GmyJkh2EP8RxU9KvOPG5+GKA28QImk8k+/TY23X7kFTt+umC+j
3UobuBBtYd6tAyuSO93WDQIXIJQLWd7W95HkCVMMOpRosj2o/cNpVSrU20UOh6YY3sDcYxyjHLK0
6K0MAt42FM6YxXLraD63csXHGkF8cPdjeB2MEa+hkb+uG2LrVIx72VBV6Y6roiyrLfJ1L4J4E/Yr
Uf8jAgRZ09DBzO4XwEm+gAU7WhtrdgzuQtAEGIHr4UPBhD/rU7x4H7H/6couPKRbCDl7FZkoQWQa
ZS2xlSNCG7AWeqFb5CFNqlRUq1drlrv2eUx8sjxBed5fbgoiu6eMkIdq04K1Gys4x+G6vo7MKl6C
bSjerL8K4Ibw3HVilPGwBKn/grQZvIgYP/fOV/8/pIU3rBZzByKGwOS26dRdfsrtuoT7gZN66T5m
9NU7SogMnbelRvSmgpBpTPsLY4KEqKGOIF/W5OW7hdMqt+CgHLTctAamZqID0owEzrIfaWaxnkFv
DtQ6z6KHRJfIesS9UqCJMLvSslutkRyjBwT+QBIUSrCbBeh7B7VkWgMslwfJ7LGCWYhtYEOkFEYC
ev4zNHW2h19Ex5HvH6A21attdF0XtUAHzRgwx0x+mrP+MY1pI7aqCK2uyJ00dOx6uyum6ZQrNDrp
5+5XS/i7gTxXKGQhIDEoa4a6uPvAdWICRJPudhRSfpCWB/DpXHCs9TgiM7vDgxyym8LcjL/ktwJW
oFiCl/mz7TX/6+GaVk6MoQ51ZD/sfz/Bp4D1Pgxmimpng5D+a2ljIe1LqwgdGMEtDVPWF2iKShAv
9LWKlMQqKIY8Z0Cc5Lk3lIttMse/t6GDoBwNaTtKXI3KCeP1c1fPe0p9QI9nsJMFvLeBMRoxBHrX
R2gZywxfpKy+1GqxT/5VVxAIM7g7bUq9fzpwU1M4Ve4ZVbXCugXEkdiyI5/7fo0cSlfR4uve+3+g
aZPMoP02zP/UyDQ9p3pszafdLBZIwWrnJLwI3iVyfn6n+0enUAqouf2Z4QbicT8ypTiscDHbRsp4
FiYebJiWe8Exgy9Yn2ah3nAM39o5pwQh6hxgOgnetfvdYzz1yltFlt95EZXhyYvNAJZxtO/6Z/IT
X3lU6LSg6adXy8MawTlxfTY/QWnmSDvafjNZDhVL8a+IFSFog7BW7P1/0Xc8Agx+Syx8MIr1FcOl
24iSVAMsVLT9W9xpjhvVyYG+TjrNeS5Zz7kuIp+nE36P09yvv3F9p0+SvE8oByOxFjqjX59WUfXj
4MKAYJrQi4wSqcv+g5WHXegTqFUNAf80752GPKtdhldkcqHYmOAlug6w8eDG0pV2PW0JWOT+6I1p
M1eQH1aFL04IwcsOFQvxdYxoQTECfV9khAoKI84upo0wZrXIy5ZaXSSgiIVl5zl6xjO27ORd9W7a
a5maZzbOk4tYOjlvggJtiw4/dD3+iomWFehvucSJT2w8itc+8W0aLpNXUqmgl2P6wMvVnwBqeyKe
EZfI2FnZFMutdRuAbfjebqD4DY2sbtPU4uEO1wuOyckJU/eLsAsGRUmx/xl1pFGQ8CieKBemEFrf
SUc7bwbIaeAQL13regil++20+68VSi74501KqYU3pAImw1hIQCJ4Qwae8iEUD1LpGMtNH/TdWSU3
WDfLLsydMY1QLMFElbWeyRYc/c1VtbzHk93GgTAdi03wql6doUBCfVuuKbNXMFHZYIfSG0JPPa5V
obNioB2iIeJyfJTXhrnIVxBu/+ThvbvI3jBEz8/ZpdODs7jw0K5lvrizyquFBvXzlI4roCpTMjXJ
Ww01z5WAzf3ceKjMIi6yn8jZCRJC6I7SO6EtEygNFnk+dmPOa0f5AnYDZGIadcqHeLwutze3Amar
WEogm7mvVPhB6lCJh1oclw1Vdmno2cCYLG44A74v1L8TeqbbKgWkJiQGC0xKwiyeJCRs6S7vpihE
Ld2LIk/rDY4Rn4HSV4SqurHzgagXx6euTzVR04vXYzZ8eShrG6CL40pehKiDd8leGaUPhRS+VKqy
fhMYZSE+WWx5oB4V4x4nKDrsJUfs6f0KOIy7mnbfsMsjImNXmzCJ7lqBiGwpywSy1mB9wWAoktWx
DIVyfLNUEyEETDqfgk9Yz6qz1PGgJ/BWA2NhV7g2OT+GO3gpxcRfgGDCfNg4i5aHVc3UScHuBXPg
PI4+11cn3e51L7JTrkh7/D1KIrLPjOSHAefiQH2jirW6zdJpu16wutVcLy8dYnoTRjc799TKfOYY
RpMxRoU84E8llbNr4f9m353XjvOlNVBK/cim64To+6jGs7Yn/GVHBEp+EbBeehsy5lXI5xPhPCPY
dFQ5ucMeGrC6F54stHl0FeYaa2axhP/EGBPayqBnClZIDF9UiAcz5sgsLE6N/Cr8ZFy/N79Qzqy/
oMjvz485pchMPpBbNEdT0Qnpgb8YiHEGgOVOJTDBaoDlSEpH1/+SfucFNK/lk249eKxaNAx6Ze5q
TJaQuyp8Ie5uG5Vf2iCF8FDE5kDUuUQHv1wntMacKSjza0ZGdGEKT+vi1Hw57a5yXTwyMuiW66WS
0UjMqdVCyyRxlPRypSQfyUZM1cSW62Hf25JK8Kyzp8lMvrDRdqulWKF2H2tR5Y5ZFc2hEiB5HrLS
lTfCFufBlwado8BFro8TtqW9lmaUXCt9gws5xvIysfXZ9nr1u9XkWG3gHsOd0jK0SBdepJ4HFmAj
X7UzpigK/394EdbfCrQwX9fJKD50waMX0zZXxsGinep9WgHk3xh4CwdvpkSGscVnfqiPaVjynG/L
sTJwh7Xy52SJmRvGEJpYM4TTXr8nsH83Qn9cVY3xxtAK+2KFufVmm296fzCLdlf2RVczrxidEbMK
M3BbyZjCU54sul1T4YrolMESlltuwuGmr/+PjlyQeFAYhIseqshTEUy98PikZyVW3MshvaHC/N+Q
Q/F4Zc4ntNKaa4AbtBcax6GO+6ZMp4wCFlIHUnxcQAoUYfEjJ+qtqhPCLOZgmUkfxx8aoTL1o2Gd
s/oBB+jt9E6liUGo5s7aa+vasa812sxkLqjHk4WDwN9sMQfSupzgdfjUi+j+3zTKSuHhonLawWCo
Oe7CRX4DwGbeaallRJUrucPgrG+9q2v2hXCsfIi404xdqPXc9xSG2zzHOjvdRhFyhGelaChi6Meq
qEKw8YCZhvkggnAcLStiy85qkBAA2vKwGJQVQJ3Lu/dC3C/TvIstHDQVzqAXvWqOJQHlNSr0MaZk
ErCIjplMX2sY17IN9bF13Pgtvww3Wv+upOyl+p0dWPiuscNkvEnt+1fWnz7NdrxcdEiFr6dAFZf3
N4F1lobe/v17CM9tBS6op4A0oTobDqi4hrOdGmTwGcmwVRGpzxnsTDZasCwEnQO4ughFIYdCslZD
Is6YpNDwvlabpn4+Mb2Ggi6VhMeyI/mBqUmT3a4moEQuW2XduQLaQ28K+QjboLHCsvWmhSqh757X
2TbvL8+w+zSfhoYE/SXFpNQSE22BEumsz5kOuItdpPX4MKq1muTsSylPZs9/ifXWmCsCKJVP8tNw
F94eeqZ9E6tWZOWV08IJ5GqIu/vBaQ7jifO3QGjwzz6jBH4oaUpFLAkEBX/9W732R9x7vbNDwNnU
UdBMkzm+Dn/o1E+ECMtdLPQ+9ZOwdJOfBl4PHKqWjkji0YXsROTmhLszWvHcZBwz7oq9ksxm57Kl
gTw+rWUfUEYvAWlgNumYcvHKkDFM/EtBUp/1gD7Azo7WPoCOaj+W+qkKZxRDvVfShUHR+teMzKZl
Pq+0kZJEioEkM9s1XeCS4PFJn/oZp2XpmsjleAttyLWXefGPxIEhVkNtLx8SYqpOa89M+ig2Ujj6
a2OUa2u9kpHs+A3D5xugDaMHybU9C9Nrfez9vLCQcP4c+xomxQrhs8p65dpmbLyDdgkSB5gJGCKx
qhdIqwRdwz3JA9lrlhF4vRLiZUO1/ovUvdLPKr9LTHlTpT80G5XW7FVObXmRzpLV34B7xyaz07Fj
WvvltMf3VUdnxlayD/EJAyq6g5P+gJWTFFS8y1g1H60qS/cIezoQSGxmTzMTBu9Bczj+KcGj1w+A
hev2T1JVmftjBrSPJZ3UMT5FFU+3Hvv/pMR8laHzeIR5EutAQNa3U5+BOqsKfx53kZGgfGPCgEph
WqAKcaAXVw3Jp1iyNH9nXBx1qdcQ8MmM6tQn4fa96sh/JmjTamfq4gge1hN+MGnpvnNO9Wmz3Zer
KGYnRxZpA0BpGaQhZFeqcTvIdAyzRUCp2xZu/3QUS93DK2leSr48mzFUbgsnhFoz0lhDCKME2oA6
0WJ9uFI5haZTIF3xfPCjTpqnWW2+/BeFOKf5OSE5yeG1hKpVSMCf7rtThMz/6eW9uRtAFyDyucIs
YORd5eDvGMgFIFhbl4PhsyznyFD6ujJnOIiW1BeCTkrBrpKaHkBEKcAD5OdgfEWE0Q/fcFNQyVhA
Lbjh7cuNMQEYLNOv54OXf0mXIxJRIA2J/47eOTOTaiRn5KNEc7z4TqSP6rb8BbUAS7BXF5TpKVso
X5OTNg7CXXd+d4N/tNRmN4enDs693QEN3lKQlwMRNBmdeBaMmRyfq+fjCf3kCixoSxkBMnNYdjXz
YScqUkCc/ONaRLflrWOBeOuE1V9q9uHb09hSxQgIQxTHAbBNWeLJmxFt0+UTvI1X1s8s2pqSPIFl
891kOGXOfJxVxRH+W9X88VUPo5n6UXXyQK9p9YVsgy0DIEbMrmBwJRgtJMPrdDIAbWU6DD9ZcqnF
HIrWgIJD/grRT4c512dqyrKyuKVKqLxVVervjRFteQ2dyz3nIvzsKlPPFmY0L6SrFWoHxFhV15By
zJdFJPKGiCCnK5XKAwgE/TzA8vqTYS1IjRXmFyLA5aNAl0d5pJd9P57ZVRiGsvl3A6r6lgBKvCIy
DPVsuwxDgs4BlIY1uXHN6RVXVle0M+w6kHr87kpRRRzS/tzZ36nz9VYE++CviP4zg6yZq8Vt9QQ/
XhtlbXvt2N+hHfwbDs8UsTDjwgqsZKGWhqA1S3uaEY6cs2vtB6pWK9vxYHeJ3IOiOmovYaKVZ6OW
pDWnQEegOnizLgShC+55VBPLbDoEW7C6EkndNOukDdrHd0rY653vq3b648iFkbDZSKGjMa6wCMft
jCkFnJikDWK+xLtn5KnQcT6iQTSUYgc4GrFlR4SowQKX/F9E/CQmJayQ1j2xNzm453E9J6McTpD0
AzMHCwYjOj2xF/F6UaXMbKDjTDS8VUbGsYUQ2K6TK8gAi4xAYXfttlCmA0pf8ZaR1oGd1uyytzzJ
mDSHBWv85dxwdmbx55Q5jrPV1hSRaUQhZB9BrxRrkYVLth+CZ8Axzp+duYSNhhs6HCnLk3MzoGim
MQbBAiOe2j5w5SfJvFmQhR5x9dXNr+vzkzCEFBByhJqBBv2XJBiTPCjvolRxVJzLibqHJLPFqwyn
aSXHElNGaOGOkEeIkVtgNIHYEXmAiEaGDIWL8IlLNnR1adZF8c4bo1b+LWipf7Su025ul3PiadF5
tWrYbFC06xWbSYcisyddTLifBPUvDGcy7CcDLFYFNoPt84zmDTpGUxqjMRswGB9v4Usnv/aw1iMU
bYqDrs5NuaqnqRZjnz1YRsLlXcQqLXIfhHbxTeFtJ6bbCHmQ5qZhA8DMSqXP2lrHrcbDVkIZPa86
uP0MQFjPmMj4DQUEx7RuMsRgw3ShheGE6AkNS7qqGGb6VEgYo1e9ztaN49JmDyFDAruXMAK9OKKw
jopCAWbt9hBcgt10voThD4Efjyc8zN7k4p71KJ6C+Enk34PmBEgIZxtAnL1lZHat9PruN8m7JZy+
sGUiPtUKUuZ/3lyR4Plm5+ywRSs54VFuGAaUp8fnTYoOn6P6UcxF350TXWaNzzbDzhCvAQMwOImI
VTlERnZsRPnjkGNRYualtGnsazROxDxRb+oYuK+f6wSFbPqre11bnLn8csNQcYXQOCk0BLyUemVH
LT7MrcOPeRxVt5PsD8I1rwOyhw4YwXq1nMxIVNN3BU0bZ+JE1kZeLv+64nn554R/TQpD2VKwmaYS
0MOQczE4s/UjyISb7luEHhd+vEaeOwr9AaMU1+xmt7lfQj2WUvsNU4tsPslyQJWJlmFDEaLHCfq6
zMocBcqg2OGD9rYFFWVTVbed8RZhNoWdjI2BM9mFFajUmEnD/ZekEsTUKmFDsB9ALa7CMIgggoKZ
26w7oIAVaaoGowi5bRLtCxinKgk9HFe+Iy8y9fRBBCVl0Nf2xBCYj4fAr1ivewNgHDx2TQ461x3J
ntw9D3Rk5EY3VKqcqhmcbiLrnCNxHiZ48M67WpyQH4ivnJjN41c22o1pV3FQtpLXQ2AnKogegW8P
iFolZvlmzRPW/J97kBd8hKgS3ilDM1+Al9zgQEZ2MKS1+uD2dcFMOUlZiprjCO6H8VpY64LulY2X
vkFow1G6DIPmAkrmsjY4Ao7I7T7EvFLXAZnEz7TUahblOWFQIIwBEFjO2LAhgCkgmQ9mkPi3BeDG
B7tV+ML/4PrVog51g9Jw7Kng2S6qo/m9BytTuNr9AlyhD6fRsA8YX0oni5beJcGpSs0kn58pUZQO
DDH2fjA0hrEQAwcbvqSSeBNwsxdj565MzguDxV6jNCdLjB3+VI/6N269vEZGY+O9ijImsgKUiSHt
lQ1NRWP1W8DjmWWitU/mWdHLLhhd+BKd7iyqMLZ3ZVOJFeO/SPqV3R1+/Gh/iyXzNfzHLz7izSTZ
Cki4klOQHki6KiXtCNdgmuXaTl8PgAonYYj9MFysvKMOvh0yPY+mQYWJfdfzZpvg+xBw6dQP7Si0
3bruU58DaiLZ4v+YuFQtWZnuZGhD2tEiDCZkt8e81+92nfrxq6ILxqCQCD/8dO0qq7ymqh6X37RC
QmVKtP9eI2kkQGNy4uXuxaG21RnAzppM94ZYc2qqYY+K+rQpT6P3bDfeI6SoPiOJtCf+GgJzJIe9
3slGIHHONHQwBYizsvojfaAMnt9552lPm7j/VJwX6ckk22vV5S38XZU0rp16L4cQ02zomyJ3ukGn
sVAQ46XlRTxyYtLbC7AjY4iqUj91QW3pFn7/ukdS0CZVmpOGWBwO3J0KH91o6AnVgmRjwG406MeM
Vz5rEUV4wIvaXqKk6uoGyig/7eiURkw4dkBraCmrrWA+Fcm+nqEOI8HPLQnssd80WtO1Q1pD9Ggh
8EKUzeDSN32hZpxZ1KICNf1qFn6Cd27WPDjdRhPBzGGoYd0frD6tKtzTLT7UT3Ei9meQxEIZDxRU
9yCHCDxGOn52O6NPpg8qa8d1O4XTwwZg5CUGSY5we60PROEefcWIWMnZWwz66HF3ziAD2YQgGz1l
qEOaX/i4YcOMNjcpAmCBKkkkQ7s/ldIlGh6QqkJOLLp/0U/mV8/YIzow03Sg8P+1RCSpVTmr2qQ4
/2UNk6VCZjoS2ellKZbn0GxPYkrmfRAjfP287jmHTI1RwypfFhkwLKt2K6/rqn3RxBahDgQLxO8F
9zyfxlizrDvMxXXdZl/YE6pNCE5iVqrHnCF3L6RHbbsWpdTeKwqtHxLCaScwmLfzIPqaQoVCOy6b
buAJLm2LxnI7f4o5CnB12lJddXGo4TiTBT5+hey/GaFlvYsR6RPqhCOwdlvXSlTnWMeosM/pF9yS
wkOiwgoffnEuUPMqxu44m6+PpOjudg4qC6oMq+TknlX9Oc0bcdAZV08u/DMUpxtYCkpccxtiwoTx
+xfrrtZPK4s/hoolVQxrBeqHNCV5WMVMWhNiBH1D5pIMLXBP2ugXFPkap2EPOzNOgGzAXFSbrjSY
SbqnfzbfehvgQIl0zMqWS9JUw7UmGRUKtlTpQdhgatlgz72SmRU/nBT5ZpR1nYagALFgiuW1Br7U
DUj72tNEvOTRF2Q4NSMNKXAUhbvsh4PjrxDul/Km9Jy2AJrKZKqvm3FHoKizE/ePD6UjRA+eI4a3
nP3KSG/lZYoBshCor4G/Vp2SACwW8n1NrG9SWH42Ek/M/uL/7AyPkYRjtYxutDwiEprF6QXJ0HLl
yePvwQtpe31Z3x/jFrCwf5c0Shexl9Jr2PbbPbQamS4nJLuaE2tyhQQj2dTnOdNgFK+UOHREiOgQ
+WQTkD3MDAEzLpaE2jrNMs+UVXhNo/OZDKTaOM/UKQAkTaEul5bhx1YpV5BFuPSe8Wqa/r7orBj6
tJLGzdDIJD7rCR4baONew0pR+/flobIZL8TiiQ08VJqBn7UMw6FkuSlrrWf/TBglGrosbpwpAJsw
b+AIWBhAn0wBR/nlPX3C3mPVQf0pQwg0wGPgvvwHrjoHD5E9Tn1PN6MivUM4wTjuvk1/+53EK7ws
3l43PiIUSKIuWSX4YNYbmadMtiqYkZT7Kkl5uBbv60C/sKcVrTmN4Fcc4LoddoSLUJwlOdBgkBYj
4fyTIi66G4oGjBSpBiGFMclCaKjlbc4OlMPBUK4zzemIN/5Ay0HKBBCNLQCqnGyi7M6wYKK3ERIQ
aRepui5vDbSk0JrV49usofUr4FJZse0JV8EfMruBfC64HO5gbEp3mF07NI/zD91ZT6+qrppXXhCC
MPtFo4Wo1wbe92zUBp3J4cItyy+D+O0D6QNAZ19Z/f4fMdiryQ7ZSmRpV7MoGQuG3e8sH/o+5SvM
yXgzllQf91U0Gdx6ot5jLJeXM5blysmKiDVtzmNS55TPW/CDoJIeR7ZHq7hdAwDLa8vR3ktHnwi+
cVEmRSN/QjUsAlaHpqWzHQaxO7bttkMVfRnYOe34yyVV3yjUUqOagXa010F95pMXkxerrUMjiJc/
BetUSApxf99/7lm4MD2PLFTDvyXTxTV7No4YSpogNfZy+VA/KUug41ZqiYu5M0xjDrkutpOVK4io
1LLmOXXwiZ38IqVV6IsL6mymqIXi/dVG9lHcPPDqoPo9K0OlwZowJXZymdiX3A1aXJxijzTZNphJ
uVTwpuTXGWd/CJ69zznuA1FUxGVejaTU4aLtsB3Pta53+mkUOwfUnWz2M+tw+v6ISCHsau82jzWi
4HTf3v/h45jBb06AV99KQ+DVwT+Nya7PWQpse+eBf/L0Uik6Rrhi5voU7Y+0/6mH3+WlqKPb5yex
X5VWxYYCz5gY0ur1QUt0UzfjKH535Wvmy742pNF8WW2m1fu74V913mr/kofeQqocVggEajr7m0yc
AfjdzeEnGrmg77eG9Ug9Tsn8ESN39qvYjHTqk6G8ug5/gMN5HE+mt4zZxIGdVzc8uCe9aUnIvOnB
uOH4P/xHqC0CEgYN7cUYlJIeUIIazlSMRIq0Hpd+an6x7xVniUX+J58klXidadsi5YfAmAH0In8k
67SguLEgXOq1Y6vtxVbNpRotzm1MeuVtq8RkXs2vPXL4Bcdc2lW01dRSRJK0zkNQbueZ6IzTRcV9
5yAw0vo4dggOzBgXQVIcgCtK7E7NC8zc6/VnRJCYRJvw9o33HABUq45H8f8oDUfJ9viSz/zPIHsE
SIINFHvkyPstuVX+iV8wPapX/whkFdzQ0CVR6pEQ96+94V9HA8nA2Nry1VsMF7yC/A9zCFygrU9C
IDxNv4zFMqJtARGd0cq6ECshwvNJsMX/wLMOYEemAItvjiUjAqGOnYqAG/WMmRWHtjTcd3VzWRmL
9uvykTx0t3m5z50XJQKuR9xDzrsnMrri+2j7nIfejyluw0NrEnUywpX0g3Jf8Dy/DSPIuVHOF8v0
8CdpnSQv7kltcFoqYFy5UHyXJLWFCkHe55P0W9Kow/Ten5j9W2pmryHaS743NbOByURPWwb8t36J
UJDOSW1kCRw1JTlKukwBxWbmB340dO6HeLeXi/Ur+IRcrTFb9AkjyJzDfT4DLUjl91wVLBXRvbHZ
ZD0mnH+LnMgOXLtedM3d5qvD8hDow4yu7TOYZOGNQ+xuCmT1bCURpJQskzI3BNsroNWVbmPdJJW+
oldrDw/LoMWv+kzAAK4/NkVwNmDNgJ6JjTa1Mr5DGwV2QKN/ZQ1dlYkHE5Q0dRpMgaoCNaSw7TaP
gmzE7qKzQ+GoTOJTu903CTpGFLqbTsFpgG8cPp+P+dOYw11d0RgchG2/BJ4tKhZHJ3jUMrAVNpbT
939+pGQ9kf0e6mf89J2lL6z90Utuz9lVrLXmK4KpPv5nzMafYJPSUElKudXQoy0XYptENg+xBqDf
UrVpAibhEE2OIHDYonRm+2W1GLhqcWpUqo80tFMx3equ4N9nGdSOW0JLMDltEsQ79lLFqKjrrZnm
cKT0gDwTA3sBtCKtO5gL6jLjEWeWcoNAt2mo05OB8XXos9f37ukETcm3j/yPIpiWKEeSaXu/e0ks
rJO2bkwpMpDSeNrWPHJHaFA6bJRlAkqJqcSg5OWlzGWPETulC0ys6+T8XYNytHtPrUfnPbaAKUza
Mj1MYJpwIzR7RRiSP/38ctFVKQBAAVr5PL1xrm5fJYScRUj1svBCd9xD1saIw3iA9rwErKgLBiTd
KUqVTdCS7/EiVC3F4K/z10/s6wumKDPn1cFlRZ/k/imSmWF5xLrj9RPH2wuGovgBZPAOa5swSFtK
iXF/XP80JdhZqI2y1Zuta2jF9uQQVZ9/q90ylbi26V5rwgyQ27DfvkwwGDGNUXXoUUeLfa2BxUzG
WxDAdtyG6filul8Etd3fdLOhKOp1MDfqgEMmmDhl+tfS11vWkxP+Ie4//QFjnCHkDnK39F2gNVUt
uKvS563i8g8FxzuaE+8Cix50hPZWdWYyCGWjAlB6l3AWKIZI60SrY8xXt6Fs6iCr/UQll37qni5o
WRgjRfOdQr9K8xUWhsBVS0/+MsGnvFPksS+qkAyKMdOakX18AfeR16u//gRc6qLLv0rsP7aLG5O9
yor7LUg0KMQQnMBlPBXctZmtpwuf07Z5uXDOo15y2YOA59qCiLY3/mDgLsbC0OzJ2OIhxNkd6SNx
REo2GsFVUXiywlFAne1n9OtJHLkhzaoxQIE5BhnBVO6OVb2IjueMizWKKDGk3UyRKXnQGwCk31/v
0mATJ/6oUqEVIbIJ+CzDuH/e4fKfo1MQC7g7PfIPmEu4W3rDGMKeobxezs8JSgoELWJBQIQg3Yj/
rnTi4GadxYzzRIG3GpswVrJHECQDgqxNoDEMS9JNs37m6jSXdl+b/o5bTW+HBVWcQEFpr6BNueIf
yILB0wpRNI7aRB3BdePFEqEKhthp7y/C+EuFBG6rjM/aEJRlGqpZM+wdidV2n8vHHWj6l4G7YRM4
zSolwvhvvGrPXhhQ9Lh9D19YHVI9ZGKDf/rGPwTmUB51V4zw37u878mehuigw2UiigOmVvRchwvd
7yOsiMsI9fDf8lRTDqk4csjb+oAhElFusz1Vo6krGHXCv+n/NofYThq5z7ho3t+MQGQzN8ZyG94p
BDsnIpQoFPluyfXoJPrK/wsPVz+C0WPAanEP/W5jgnmPM4mEtUwOi6a1vl9YaUYNABwXVaK4yWq1
+9KZ9rt5vq+4sczIDOBdua1g3xlYxD5qswcLCpkkJm7aI+Rw2QciixFbrvieuJPkGrjwpMhaJink
zC7CXrDUItEwouxxOvWZEl/09p3fxZO+EbUtOiU9N3DlvC6EXpGp8IMmOttkBaUzoxCFzDWbJsOu
4dQBReQyVflDj4PuVK7lX+uqfiNgPVkdeEkWhdszTC8sUseb+OPwYu5s0JizWslmIrz88tKUxljB
gOC8yITxnUinXaZREO8memXT5zXXB258ftwclOGOu46Z+z1r72W4M2Y0jGpxQsYq/2ivh9kkwIiK
/l8p4Qj1W3ps2YZ0iEh88gJe5UYApOTUU0D8Gtx6X5g0fPkuP9vbhXubTAZnukhpX5EAZ9Bn1VK2
/Go3wNSohc+ncW0PXMvUGUmtyWr1KEU4xYZUeqfuP/wMxC2HAYxBO29iqz9qw6iXvYokF9+zbRg5
UTAcrW+antRwiM79fS2YlUZRbxz38Sf74OaM3P1GPW3tT8/kPdZfTSl0O32H5v8wLFzrhpJhG3uT
6Z8kfx6Nx8E8JNZnOiO+UfY1hZq0CDbIjNNkAbCdaM5fjOori1GLRUGPjxB0Bjs6fAglB5iT5crL
Ob4vfZsj+hdOTLLSyX2RezxVNvz3rsYzEXg9Mx8DvU1hpF7gbs1YXPkBmHg9IvrH1v5FehvJxoNC
IjZCUlx4D5BR5qrTOHA/ipZR02rFgPjZZYi4l+OAB6gW5O97CHm+FatMICV9E3aCNdgUWM3OCcXD
9cvzn9J6ObOtkfaNDnlrEKbEOxPr3Xz62d3p9mOqk3qQRz9VB6yBO/Fnfc1o7jqzqcq0PWSh1ZvS
oRNeAejP0lLtg3mr4sMy+FsWNB21cZyErvNAbWvewkNBU9KViqaVVncQn4/ESpWQokXzoU/nV8s2
vQCvaNb2QI6Mltqzdnwfc6UrsF7CIsk9LZHCVH8nYLR7udnRmvTsAZDaJQEPvLSUuxeU8cDKWxde
FcKscgH2gk7S2FFd/E38UA62y56fEDkSvDjItn1s4RTfoikA+MBBuK9CLfJP4lyHPAPJRV48AU2k
AsXc10OQyRfQMe9sVAvaMduo1mFuyq5AgVrHt9QcyXv9gz4tchm7RgHRhisLc2DHfwUJchViEuvx
21H7BNKy0cVAewllfDBQwLlVDvmpTecWE91A8ZuLVfb5WUd8YFZ4ZzTNwoECMmzslmUNjRuOpnOa
sL76mBh28KoytxZzJwVKlM9FPGKbTZGoynKiM3dmlSextvZAy0E1IzznCvK505KiFv9EReJ/91fy
bct5PZi8grdwI3L6ao2cRB0jZdV84MS9+lrEltpP6P2IHgrQKHPngegJk7k9y6OVadbM7pyeq+uZ
aGvn24PNp9d4YdkF/uOk8PSsuLdi75y4qCXLHS19Pwgxjr2sManSLESmFnIYDCnVrDMywIMq3Ax9
fr1dj8/7bzGgCHPbqDp4QD8Dr6ctZZgwcgIpKlEt7cipvlUlaEGHmnwCrwCBaBijQrr0EgF2mtKM
qDBdx1mv2T4irj6TkF8XQL1E6L9/Gu9zAN7drLI/VAtnxKF16N3pUPg6BsnC10EufT10hYNaSmJc
Vj1NB+bmywqhgHvtfpi39V751s9sZVtLHn+pJFpRhBt/hQWLkJ+rRncbTdlljAatjrOUNEKPcyhR
4E7cDx581zRi6JMazfsoKBY8yk1pmo60oSEuFFl0SD6SVi9NSPC2pQzmtC0tV62vcBUti+TaZiKq
rjhBC6j1Ql469PKG4CPF1bhQdKQ9VDQq/V01I1f3eKmYeiSWIj2DeaECIDnCTP4HjMMIy5RXgJMU
aIXmsikm8t5vNt1mxjx+HdO5hTe8aA0f4/j4eTshibnbRA18JI6bOH+aqoqekw8nj6mkQGSnkT7e
+bxGY0o/KJ9RIE66ImNHLXLdNUJeHN0gvBAGNlWn3Bm6rfR/UyXd2EoNNoL9T38bGaZiBXksQlG8
I22SGVvQ2lWZAMoNcRKJlk+lMjapcvYzfV5JkN/vJHp4MDNt4D8EK28IqwUIZFoTjJsNv4L9Fq1x
YxrOWTHeilNbRPvyN8/xep15j/zQGyqEahJFAjM6ObOm1LSxVVNOhzc1XMexSFAhrbZ0UU5/Fr6d
81xdxWUM35zE5zPUPeyMUzwVTdP/oPbUcYkCjbf3TqLtNAMU2FqkrVxT43xMiBHBo1O5sbh3xAok
WTno+jSf7fZlJ9Jg+yk09f1USypRKQvz5vsnN3pBMUNoTNXARijaOlaYuBRhvLp+cIJZTtGg5SBu
smhT45oKC4CcKy7IeostbGNiVI8P8IzKUX90PeaGybyKE6a5wNMRxXHIZaGY0UNXM+FM746n3Fsj
pi3h+qBaL1GRWX2qlhqR7EFN/6Z1YUVH7VKxFrt2S+bJ/k6iVKQPC2uTlZY4tGKTv2fzwUUW5w96
OxVrMtyyOr6cAh2r2uTl8O4SrW++nLqzoLQCJAEK/cyxJNgOQRChtHzIx7UtFOkMlFNIDJ7obebc
9IMZLEiFYTx8i2JvHj+63h0s3RzsbzHP2mHRChNTvHR/6APcfYBf7LxgmduP8WJXWDD7AW8BIaeY
riMM8S5aoyjEcExlb4/mcWlRoJYe1hVyS5DcFrPY6UZffZhYEJfhUN9MoQ+MJCNrsWA9CGY4Q2kC
tA3Yz++Rbm7aPAFh6ZGFSV+DcBkXEuqJn4Arz74b4Np0naZ29R8Syznn1jDuk3bnqojEvnKqPD25
+t5QgHfnM5qFoS1ZBQzIN9j5gF2z0NQddANQDiXCbqwochzx5DSf0fWQXswdoRyEHlv9f8LNTEBM
uV2YHabGhHcTkPD8zyaCMiZRik4bGx2LbfrPNOM9ByVjE0Nc30ZvVgBKjmO/oz23mugc1nFfNrW2
wyKADUm4fCXoFISxUTfnkYy5aUXDT67H61MGlv8YezCsM5SEIO5IEHK/rSpPfw2jk0TJqwgiTn9G
IDDha6wPYCRKJGOXHUhU1RfpbjM9d3o/WAD/5wFynoqeXKJ4mBh2xfPVhUYiK+DHAMcfDDlOpnHe
XqDF37C+53V9UyiBVhf5e2xZEwyMfAREFjW0eiZQ+swBuijGUAsLFtKhNWeuqD2ksrwlzXh2F+95
ZBKW5AwvbGZbkxb8XPCKrJvhy9POYl024OnMnfgpW1BlQIcJJAGw4HAQtkOwdQXaJWGig3kL0Soj
Fe3ZijbVvkpjFMMLfgCXi8YTN68TWo2vGp2UZbGHkj2H8hh/5fyzMmnZtmzB7QxpsjcBrl29GQz8
cddK/Oo8b/F0Vl84Mvv1W2v9hZRwlvhivUv7MjGd11W6sNzczR51I7XK8WVy0EplPyyleRAyz6JK
4lqXDx4HVpbFNgc2izHH9tii+8hUUU/BUQ1clJHgubN2N7NDp8LkKWr/gf6Yhi4Ue61GQ/vOb4bw
drSCOWnkbf8fDvFNlNwCilbrn3WKO8XRdpiZ+cLn85X4/nEmRBpHk6Yx2ETxZMRGsx6oPgwdBV65
YkKsahSWrw211B+N9Rul2HcaIMYYo+lG2DELnCfRGt5wRT/R6rcPUtn87CBtRZ1R1P1TCQtZL6LU
6eLTIZb5UVqSuBfHHrJoHIMJ4OEJCFkqb3WL38ioCC/gOGZoHaE6q+KwCJZnRnWOhno48M2RKnsX
cQQ6CkhglcNQCE60225kk5FqiegmVLXIZVYpMMJAHYtx1iZcJCHpHdP4w57oNQC9RspboA5m1Dd3
uLR6vmJr/162e6b8TM0feluR4Sh7tVQ6K7B2orW7Ug8yJFNMA0Svh+mL9jizBA7/jUVK7LiNI8N/
//cRAkxriOsn0MsLgRZ4DlWbZQpy4Bdm56IiBC9mWpYkdqwKSJQ9MnKwIbGj7E03jH5W+JYOXO76
kuDmWBp1q9m840RAmvLGz2UIQITUUJpljKOl7sFgCPoi2nNHTGiZnSJYwb3SQHhOjWgqeomge1ai
Qi+lTMhEH2gZbFjDycb5H13lJfPmytPj7Bu/gVqnmQmbdrmpIIKfknumEa7YVYZvwEyTchHlo6Vp
YrkmK+vsFWkUtn8A3p6IXs6Pu5N6Cc1cnofNWzao8E8azWaNbIFrx2zsmffPougZeWDfErHSXtEQ
1ob0MjHWH14P8ygYOCtG/Bz1x1WzCZ81js1XsvD1IxUNw6SCWC5gFnYKCi9Se+FNUGHsc+WlKIdW
OqYqgeg1kJmVe2F+xwO+epX3Zyo/xp9THB9lmIdxUZo5IJHfIgO7Ni3u5WH5U3T2HAw4o3JsX6jF
VYCZjSRgtMDfLNzCIkpT8KWxhTNA7MvJScDuxHq8zlPxcD4EUd236w95wCHfni8eVBElWzBjtat7
dV4hb8DTfquqaINc2okgg2NyzJ3SuXVLE/gu1/QJ/vS/jpOHo2V0md7TgcKrxlnOk1xrWKt6dyr9
UBZuJFLM2iD8qy1kn5OwW+phgSQk6gzUfm11kX7CibAeaK4oTStU/9KZYPidFSnyKJkISmE8KU3n
ICLtP/S+P2AM8d3XOBUDdGSoqo7ioEivnzN17emRcxY72JmaUKNZTk9x9Qg8ccQJam5KyAykxzGg
xHQVNJPDfi8b0ipaRDqQ6RdjKl9HmZBDTw8iFH/gYBBUyDofJnf+PisXFfiEcm2H57LrkSqjc4KN
6RF2rT2TvoeJb8fornJPmtZrqEQkqssgv9AespeBaXFPuIOQ7SeLYsEgXWBIePu9V4xG2UJi1qLt
O63Mmlx6KREfmWHQFYtqdIudP2KrdwWwVjSrmJ6vENzYlhMkollI55cjSovMcAHwpTHDQVyfykni
AFe0oRQg8ZS3ERUyzyp5aHCprfPRplpptOzB+1Uyp7ciDO67lE4T64fX5aIApWBKc492WoSwxP7X
h/g06FTEv+eEflBsvCfubsJnWStTMI0Hsgpi//bxnDWmCQ03kMe6/VYSCEMy1qcL0Y+IGhdhmMz3
Lwt9A2WFsuotHAtUmN6f1h2cUt44N90sJC3a5o9wwlyAg6xW8H6QxGIe5NHoH2OM7oA5rHfvpZik
kVgFPlsO05w2CLJpCwVufvZxBVR3T+bFa6iuRbTksuMS5lGd0lc6uKjnmlRdyAnK3SLBYJ4ZMUK+
Z5t2dQOxDnUkCqS+9fWjFRIj9GZ5qOO2Nd9h2gtNQC1LexlFSTWTyN39cnpHe6DEyPITRlyQbhWm
+GdO7PyDpaoqYIVQ1lGWyHqFBa05qUlHawGkf9bBq1lcYAZbAWE4qkFIAkda4jDrEC1OZAgiTiXD
sJ6n3kBZKbAt+gMHFGAOF69rvlJZdBLzkUkTMbBWItGmdThHP/gW39shAxjG2vAyahNNFKfn51xu
v5WkIIL5E6YgloGwAzuQEUyR7ZyW9fZxmslBdaNaPcvwdPXXjuh5eXZ0KI43Fu6+B98z8mNbYeQk
i9Jd/IW7csLLtCFT2aE8c4eRslR0o059sBdgufa1T3VLe/hTNByW/2Svuo6dSmPD/vV4khybAKYz
SoklceRb++5fsPau/KopuFWlIX3KFlD1H3whj32JUf0z89PkFdrRU8k2XMjhMazvin/jtsS6z2Us
Sbf+FqpU38gG+VGzaUI5x+lJfQB+KwymMWgCjIVS856GScB+38GdCUpwhuYIM5KBNTeJ4SjdN6M9
BulAvwRLTuZIwkCsKycHPicqmW1V5SfUk8MruDBhRVDuYEr5fDnrEJssBMMyH+gEyvSOWx73GFl3
OQytXJ/+Odg9Bp8dleU9QYzkIe/rEuDVg110DySXV0yRgxidBnVZLUm0vCvKe8jGO7+pEzqysI3F
oICYKnO/kaQdY3NZSA5Nt9mT64HGZ8yDaeLBS1SiV+vHTaj6hzE6AG538FTQFWdhMnP9PFTSyS+s
2btUNPHFHD6EvuchBGRPlppBHGCiMYeBWVRrkWW8k/hZzTF0CRCSeK40v0y/3kli77YZf/IELKYE
dZQYOmPBHGSlgfGzB1Uyy6UZ4VGOebTxKNQycwmzKXinpOvH863J1rbnw5vsuZDMsETADeBkLIGu
xWo96SIAUzDT8iXct82NUD5dIu2BX4WoxaHbt+F/bQhqZHitGS0PJ9AhewHYFRM6aU5PDxAoo8pI
QLtC3IPCjNyQgFgGOqVTDlZT0Oqyg3bRYn+BUbChTh/HLkchCcD5+CDH2zG91FEHo5bsOFdUyExj
d9nnH+WTBA46w1i4a42qA89xUp27JCvdJKRh0qOQ9lUBcG29BJpMudLKbIx+lupnldhAJMsPCMDu
XPcXtrwau3IoeYe+wl/0WVk+asZBQLq/Dd++Yupg4nJW2AeW2xFa1/U0zCXsBwDE4Tko61/fkV6l
vV6k66xvkRy2GY4mz6a6RBFwtkGpmoeUhbeG5A2aUqTi/PlgcHWlHX0hCo9d4xquZOINUozP0MdM
1hdXbguP7bOp32YK2DygWmLdAjRPMnVY52mQs7EE9Cviu9M7/zibWmIifVFrdzvm+9kViN4I7StG
nxN8Y79WEZIJmSPAdWwXpqsaTKpGfFUGDvXl5fyxnfAaob3PR1wTijCpcKYEZItntW9M+O2E5N5s
GYgec0z+PgBJTIQwkq7uudMi6c0q5ZRur94UUjWf60OWq/85LVH+i/3b9n3VYfoCfiLoWhO2+oqG
s0L8n2ikaxzJpsAxphXiIIYb7EMY27gBlEfmjX8EpesPo6U4/HUtH9Dz7OjaXy5Lo6MP4YhVpyXL
zxSG+TFXHCxJQGUm1NFCFrSvz3/LmmN+3MZm6GOVYOiyTqd48K6ZHsXjYS0+G+4qQKGmJKG9vLVN
qqLZf1hO80HZ6jZTX86mOEJpN8hU9hSiIcKuvXp+oThp46cmJIXfq6I/QH7rg4TjEooij2wsan6G
MvTcebFVZKZmvE0ujIw1k5GMWIMxDL0I03/L2eyqqtAX6ESoXWsk4ESzQx7Tuxif7dIrRJ7VBe7f
kpjd++zYq9VGmvhZiwOMuEcTG9K3V3jLbA8MGRmVHkTspnW18KEw+cN2AfzLJpETogxrqIxO6N/6
SXeZCMtlgzCGZ+bW722rqZ4+9ADvTxpy7Ti8ryI3H2q1TJIk/oKZ3QH5b1pzcGxtiCJkQMazIuYs
GnVy7O4faHReUBp81x3sXVwnfQOMoBQSKdCNCba/hziHUJupEarnrZjW0B2IWEJavbWFFVEh8RsO
Lss/azcPnXfWaHyujS5YSWHakJ2wwWhWrq6HUAHEvOgZR6e3+yNY3JnivtJoyylBmyVeq5DicRyh
vHdDjoICmk12FKov1or5os3z2Sf1lvFR10166NFmFE/20az3UjWeHYLZ35DOVJfYGgEnVnsfZCQr
VUxIabp3zF2iNME8M1/SLSrcZpcgKuwrHw13vEH4ku8PnBqKQXRz3HryHoAE3CiuNxBwArt/Usv+
oUVQbgRONNkDgPLxdC2PeksEb2vlcHgaYzMGKZwhbcCtOIbXDk5QtzxTj7b3j4aCF6g5GpCAjPGL
7sw6xi+OKLHzjIc/cNex5/rsrF/mRUUBjngAGkLeISBhdt/efRp7R0gMtlT1kNgh9+4ITtWZz4a+
MhtmvNWOuiujrdqerugeVjqSCPopqGDGOpCOJmoyHTJOoXL/Gkk/45tGVnnA/0drwCFubw2+U4nO
GfWSME4zxlBoU6lPFicLrQFdCY2Ze+y4CI+hBWYCCZsK+W8AMzb3WeAJgPRs3OW7fUFIDmvPBqDS
vV+6qX3MCoqYMYtfYjHrRUFHGYqSC0ybNEM9iT2zrrd1tL7hAC6TvRbxoU1MrKMPekkkqr6d4Hyz
fCKb5Kdzc6UwqNVliXMQQDLC2YN2Fjne8rjRwXABapDD4nTKQjG5bQYgT7eyvcinXs1U/K86mS1x
VcQrYYjwIJ3hhR5go8VKJM8YpX9MdbVNpWG5KxBOm7ndZPJ8Y4z4gEmb7QWOP2O2+LKTO9hM7Quz
xbu1bBTrutI4scKZoH683atcnxB0AtDEN2PaEhMw6FnZ+DAwHTHScNpVwSnT/GWBLUUw/jwXrWzd
9v4tLOIxN02dBN2aMjicc5XWvlZn/oi3xWpy3tbe2R1vEq1v5dbKJES2lPMgRjduFn2UKTw56qaJ
8Hjspwx4gnkppIxoQmLwGl+GhLUGxuV2mpije4C7Ep2CD9TSlQJeLWYlEmVbX67yg+/pFuICAcUU
1WerQWiuOs712zVlSYENsczdUgfErHlx2EQ7IzNUlC0taLVnxqnzUJINNRM9GXLvSFG8TJ+r2D85
MbFSYImme05vT00lEwTHk56CAhWdFKxs5TndlLU5fuSVCT7o9qYZK0VxI6dLWjLziJ2sNueUh5b+
SCGYRmrGpMWJ94StL4WnMPKWHs5z/vuCt06capL8UwLaFacmaVDK/2/IdJX/FJJ8qjA8CDOI9Apb
/EcJgRNFg+pJ7w5SVhht7slvvVcsfkjQ2VdOxkNXKvE7AS4fVZ911wh2TnxhqL+Fi3KbF44EafcT
5HXsZzsrY+LjuHSS503hLOpdWb63vgvoofLard7ofYzPg0Lfnp6v4TCFK2h7KpwCtaHyrEWg3zZ5
+1VAjTpOn78euUeQaykiStaxleyZJQG8kRDrlJSMVyBVMsEQRD5K25MCCUcY4l4lLi+YqELDEJ0B
UiS8Y6tiY0Jk2dLgbPer6SSrIbyuu31UzvUz+5GDQZoVM17cK9Xgs3pLY5FO1U/Y6uccYPJnESqz
Xzi2MBU+C8NRMlc3O6cezRdnW1L+PpNcfb9XETLPoMgsIyY9jFx2rNR+4NLkMhVHm/5uKtnPPCW2
zvuJMQwX6oKiFXtMipNHY4xjVnOike5erVzlvncjVpzC4bl7hkydALYwcntQSw+u2zW38dtP8ujp
1Dx5XWR1YKHqyTtskT65tTS/bWtNR9mfZkryJaqWT/U+NOiDJ0KiCzgZ7CRedbpejiLQAkQpKmhJ
Pd90cwCxeo3refVuyDcZZt3yGK/K+VBlz3mKqCJ1Y6DOOSrUyMrKDNgRIXXfUsz/N5WaUR2QuOJr
JzxqFrUN7VjSkCJ7Rfn573FL3vaREL1HGj+z5Om408QHxgQBiyoH/pbxkg4GbaWVNQn3jZ+7tsdl
VKXHtG/faa4X6VhOG8qPsBRNncKJtqauF+aOp7GXBbIQxmEh3Bx0kzhDdVOT88v7i/KSUg1+cJWt
mKsbSlOOYVm4e3u5S/QUPU/IWujgYObvMJ6JEKi/2wEx64HpyAP8wGeQGzKq5BGBYMeTMFPLcY4o
Kq+Ik6CfZR8jLU6mKPFf1+uD7TAqQocEjNz+VjdmgGQtoxsF9dp7JbH8pqQ94Kkkg/VuODA+35eB
nYA9oAwXshxY8uW/YAmOOY70s0LsCWVS2ahf91rMWcGauIusKAYzgHagxkQB4ydGCNC8Iw9OF4cL
KODqcKVMNtKXrljx/EqhLuvHt9sK3OTFJ0jDDE2MQmLhlLEq+zgXfDEhN3mUf+0NYhHrA/DbKFI3
iaq3yzifiRRMiJ5mA5U25pNP2I9lJf97EqWzpDnIGSnbNuRuI89FwKsD3XCkjQL/wlcKHGvqWMHM
H1Bv0dhBPJJ6rA7BXrfKahh7lQkfKx+aCe4CuHX7v9D/80AGlWO9hjO2hPR5Vf5rlp9/Uq3LW4Nj
nnJCJVQK1tKWpMjgdj8eXi3RPZw2/y0SWFYB3zcyXziSpSJYC127gvZNNz+TuQCN36DPHRYzReul
zoJU18fW8aqN2Y4G6O4eWsyJZmYYrT/l5ks/RSwS6B6vDggxwil/4RXwrJfKtos1U/UQEVBevobp
gkrFncs16/DcB0duB37nRgYYHsios8qrbzH7oQifVLxsdHTn8mbYp5ri22aZIACdxpztc02zEBXJ
s23uBP70dF58GeeqjQ6V1WA+AEuqlWfrEhyU/q7oBFP6x1E3coZrrywDKq7Yjf5sD1KB7dMJW+er
MPDBCGfxelOanTQvVd9mBDFHxyonSbvVuVvUuK/51xLyV8JW49o/N9EVbhsPL4R/zPvjQUcoVyY0
dIEyjof6T66j4JUYSK/t4FZfXwZJQrRvrQuY93y78gc23eW4UrokNneM9WSUePFigi/c5bfkX7eQ
tWqeQeSEW63P89XGFxtY1tBeVZKwQR2akrroZJ+515ZZQONTOHLsYyCUOict6ARv5yEhPu04080U
FkAc71vVIu4QpUABQla89ZuxuTIIMlzcSKVrXb2P6Mv6W1EnAkfrAOvsjTmhKQ9o9M9rQR5+i8Gs
Da2bQigEqPR1dVs+2WoWfNB5WOcUsS0EpCsOqWZne9yxaeObHDzc63dZccEQ5PdmlV2LEIzDlYln
EkjT55pESIOJsWZhAq7kEUuK693Vj2DU7XQzDs3LxGrjVD31cNT/z5zJq4GfPhi/eueN7h8GZAkk
Q19ix/wEnejs5jxqiPcWj/aRR+eFzbdigklDkH7BNTUHXo2GXpUBGRjhhZ4JN9Kga2PBJgqYB+Sf
zRRqB/vT79adXKhhm12deDXxXvG69lFwHzp5iBI3Hrw75BFSkiS+/64jtXqs5bRVkgNcvtp6j/9a
Yhb5NWWG31Y1IcPlYU+mxuQgzLr7Df7uEmBZugej4momLmQMKkPp7fhJ66A2P0AXn9lvj4D/j61Z
BA3r8jXSKSHTXgxJcHmclrBohlYjX5vaH/i59xlXdAmxqbcFrrVQXYah4VycLMUvQSt7YiNtAvs2
RlfUO0aO8gssW2j1H+TpReogZdMma3TV706zEO1FSoODlpwuvkxypgS1xk4EUgYc3kqVBD+L06uv
rLf2xoz8wo8iGswgnw9SEmTBou8sbgWW4AjGfzZw5xUKK0s9L3iqZD1ZWgflpqZyKlcX8nZVoHdf
Er5IXJv8PfXrNmMzy3aHVQijZrl52dtAD/KznsBJJr22j6n0JSjDvrn7WekjBInwmKlRXqXVf2lf
FofPt5zaEAOlcpjzXloE25iZNNBLLRghcBd2zcBQf2NNXvf4rCCi88L42ERffchynJ93BSDgAAXI
Df9chNoei0ULdJPS15Baw8O7WvbA445fflEm7yZhV53mAfmIevUI72aWsIxDbRyxmwHam48KNOkg
gmCAOR71pMaVqPFU8QMSQBJ9qXOdwlQzTZwyf3IjqspLj4bOfx6BTIa1/u8yjOqzEAEG2RA4mZTs
dFefruM35O2aEqcNRVD5lUCz7+Mdi7HpDrcFBezm88+YydLLHgni3yH5oxVDSAFgBoMMM9vebYjL
3W7ifGolkZLV5j4i+CmOjSKxQSbWxGdml6JR+qEGqUEy7nnG2NUdwT0t9uYcSMLpPeQsXpmj0qY7
4dFPHJiAOhF9MU+gJbY1aye2rVkrTGqsAgpMjtpWjCa8nhQkt95G6Egfs1OgKWm2qc2L732VpoJX
VOi9xoDodQKsrnwh29dvbMJdx5frEo+yXVkCK0JpwJDZhcpTlFHaMDV6nIMpx8D2sX7yv3xhyvyE
ade/nV9pagWRIGf7Lv+vFYSRnIsDO0OVsK8uOqMGc4RFlwXiqG+KAHcC9Qij39SKgC7n1/oPoxrT
8+nu1Lodje3Fl1z9n+znBexY/kH7LI8eVQp/D2mFa6GGPb7naJik8fbN9nrtP/OkDFhNONrq+bCE
hrcfTGhfhHvUuwCO4RFNllMaJaBxiTAzo263i+IttqKBkA/EJgePxTF9SIHKCBu0ygjVlK3oYGUa
sIukNnUQ1uR7v31LDmRxUlO/TGX42Wf0Voe/FC+uA6JIusGiaz9j4qxueAKX8sXI/f86MZvmyAPl
RlcG1U9vkpVCqExKgCbNM1S/uPvs90DLEB+IwncuHaTokq4np+Gni81bOF2VYWpoF6QPWNJiVSqE
PaK3Tri4YHrhlPX9zjCIYQBbTywHtf4FgtmIWVvTI1gB18ILUsoIzMD/glgNmtnsgyfe0RW29+nI
WCP2pBiDXLSrXjbxFcLKSTQ+4bbOSdn83awehYMld0ZEgHPc/T5Cj9GSjB4J8MEIAv0nNITw1kd7
DSZnykI1tXe2/Lwzul/y3hjQG9CDsguQ8kNtSz2kKKlJS8Lo7n+c9uOC5uV6DMd1Ejn4cLzFAyJe
OcJArbwnJVJubLjZ/5I5844QTJiE8puIYLzCRhtfb1B+f9HTqWVB77onEbdUhuvyTEqlaKpD6Qh9
zb6BVChGGdwuzUTKi2ZuaB0tQpoVg3M1v/kzyktyVnoNNLBycuw0eiB+L4K0lMUXjMk3pOZyDIlG
lV2YqZAl0vMSBB++9brsM87eFgTKk1wQnIODcgVfOIKYjSEsV+uBD0KrN/h9On5JMU5SqpM1+2OM
idFvP+KaACIGf9dIACLzGkyUmPKE9AXYtTZQby6Xuf919roUV+lugXLE+BYh+Mz9gugRogN/wDLT
zuIaQDiFe8E0g1u8N+exEHoHN5H68p+cELcbeQz056Z86BrRB+pni81huzwKQEsxpRQWaNVBSedg
5NrkwqRBs5TpEYjecO7b4mGfloMquA5dVhEh37TeHyfxh5N1j1xeVUxgsr8+yQzukATdEvK9sFKV
VdTHZALfszEyBE1cWAt91kTwQi6R0uSDdHyPDLaxtGyjj9iDmyMPcA7+msyT3EeoNmVe7ur5aOq8
ZesCGFRXjUssEq6UOKwFeqGf/AS5fFX8PfB3a44ICu0O+RpS8UM8wqtyEiivPBZB+3lC7RQBglYT
MLeWBi/tUoPybZruunraes3REZ65277qVR2DBn4rz73SkOd90QCePNuGBlAsZQtNKs8XMgqTXyJ3
y+0o+5p/ER7mP+aYWuaOjs+lk545ZUYYL2LSdPPS4zGtRcp2q6Gms7zwtoUdQ28NHLxVp9sXLz7v
wE5sBJ/s0uDNdrBAJBlGMIxe7B536lk17TJwNcbbomTCKo5qFcNcvOvE1CmurOEof5ZPvjmltdqv
M0Pqt0H8kQ34/Uyu4XKAj9XI512K9MlaMbpVoSQy2LV6UDXm9xTnw8lrzq3PvIUcQsEJb5D1Ncfe
3pdFrQ5EFP27sz69K7WZazM1o840BzxdMAlFQ1FHZKw0mCVpFJIelukYeoWOROycxqn27VMffcMS
ZAMw2EUqvgRBpTWuiAabTYnZpcDhc3DA86w5gqeohy2K3nByr+qxeogYR0g1meSbv64aPfJVAe3m
yr+sklg5kdukRb9EiIiZiqOrZCxvD8y/EXu7Wsvm2rZk5I4YCppZ6hoGmCVAThJhVsziumdbmTB/
oTPDL6487obIBaVkHiBOG0vjXgxwDMYNIzKCDBLeV0roQDMZNp4dlrv2AbRjbXzIQ0QKViyhp83O
eaHzbDrx1JvF765+Orv7F5TZU7i9bD0HqFCG83n7j72XRZRz0bSDnblfAAeeRsPSKIjKvellQNOY
y+Ez0ZYwSnpV3Kjf21zwynJflL2C5udmM8eI6ZFPCx7wJm3eq8WdQdNCyC8YluzTv//MIWvB97mq
TlSSqQx0QMFFgI2lqnNeItBd6fanqtp9EsneJcwjarBNVOrWOjzqAu/+d3AM6HmXWyL7LbrqKlXV
8rhpw/2mwSZcyFPRTHvsK0bBleCKOOuWxdWNpzSyXA48biKAKU/ImgV5N/oJUARKWsnlw6dsajh8
yikOKS/esFvKF1bvSnk0xClKXJsIPb+kGjrfLZYKMFq7Z66hFELyZlCW3vnxDag8jgmhsKMLXXLc
dtATHf3bLZR+eUNpuNUS29JmbqRSVYZq7qrJJlD/hLdYy4AgQImvd+bme/jiPMWr7I4UVUhm0kx1
tkUFhgPDOADJkoOSpZ5aZwQIW/mVn4VDXr9RSx9VJz5sMfONyaxJHoPNbVEcA+wjhyg3JdrgTuZR
769ddro/SzCZTvGcyPkgaFiZ0HMcwZIVM0iDCzBkQfaDcgaLErf3l4Ya1Uim7iuRgqXFj/S838bz
GU9qrNBZFHGp4ek70DI6fvnkPa3t33cIIwiKZ5cBAuNJTxGKbYG1ODiQUEGZLCb5iOqRk8ofQdms
iDFv9osES/gxzVno9NLJqNnrqiSn9dqsTHM2SA+RErjw2F7wASshJQ/IFoDLXqYQbwyNbmqxoUhW
cMeaddBhQ7qEKBa1MHrl8zZAxwwcdXcTv1JOUcjnKkKoiCelGOKRNffNEM8OTi8RnKgJChKr+LTB
IXLu2g9SjcKE/3YCmJNcs+t9OKKwFW7ISb0BXp0ncfCsD2HFKM7qP3n+3K6Trcrn/jv1KJ7kE3Sy
KDSW4jTWvZ15g3svaPcm9EEyg82Ncd/EMr+BFHDnk0ZDUN2si8IznCWHL5JoORMTdxyF0ieKt51Y
sJjdiz6mTRdN8RzCfkiF09UtjFQbB3ol1RZTz1WTHvlAYteCZMzx/7Z4fYn0IbfLhAtX+WYfKQh6
hq8ifhyuDJOOFhDFkc8bJaqVLsycLaqeSQhfa5EfPoIpGtZShdANg64wfNlC5VqAVGHpwrhwCKLB
cXNitVL8huUuS5U+kfgltKjMGh/Oexlw5V82G8Gr4LVHg+kAaWJtMQiD3PhQGEHalIBTZnJoQmBz
hcbfWHIUM0cXZC00upX9w7eI2zTIaLbkgRc2u1wlyD7jmqRNi+/Fr7BofVGkZpu2c7suZk1+A7dE
V8nrYgBMkPitBUQNzieaI4Tvkp5mCcU1gx93oFzIF3Ije0fOUtKylik//uACvpWGyDOecSwdREW/
Et+Z8F/OgZtkKw/b6qB30BEHlzoDUq4+9NSIGuS7OWmM2AUg1AWtPllnpvV5EWQiffbJmj9XZyUN
K2OzOl9CtcR4VRIKqAB3agRMdGnesbZ//meNxEc0W2ZUelBP/DvCbFJFRnCI+jCoy3L9akgpZT/4
LfIJj5ifeHkoNNtSZSIfvhzxDVeofgNLWHnG4il6Cb24rfxrdJNwbglycZNi1hx2CuQbKJv7YxN0
Hm+vEH9tOAV2JmXvlkM38TErwyPvrmuUGfZiKvG2B/dqOPtI4O5rxXv0VSApz6SdQzfMwF/yzhV2
ipeIxzNzqYjqA1rxdCxOkW3OypL/hLV13lQ1bTOke94GQlqvAKuW8hyW7TVVuv2QgAiyBZR946Ky
6hnsDXxmJHw3KMqrw7MjZJqhUis88ZNlBuU9fDQ86KGwSavKQRYJccOOvgep06zYNH1PzRMK550y
hih9CVoZ8sY9LGqhnYRVVXI765wLhZP1/vipNcSoWJJqfHk0sM3QuwiAstksqpJsYaqL0A4D8iEQ
sNKIYQsGnll8s7J4QDOhe5vc+DmtOH3WboCpOaB4Em+5bk8asETYloYvO/pTbnqL5gWeJKXnSRs8
LQyNmAzstRSK9J3e5M0W0iV7tVwjDY40C1QN4Q+AncoInw+9feUx8jptT/wZqZgIZG5EqGdnJFYC
/wK7n+8E6EikJgxqhU9ueXsht6qoYpRYGA9DhW4aq0tmnKJY7AAcdzgg8lEIX6Af2/f4d9h8Qi0l
ThmHXhLbXo7Og5CK37LNCMCJizp7Q2gVaz/F+KOk8BW0xVrBrpsQlo504fJIjjyTqAfMr8AVFoME
a5iQOkaWoviAy7S9UozNB3KWazD/zEOgoVEpoOuTMZMebWtTY0nDb7pNbEImTAQ/AEgxGpyeENDG
jD/0aG1mxAMhfbVpowBSJ4B23AXPd7R/6n4SZwkqlFkl8Vc5+kJAOrUg88+XKu99N9eMT/H2xyJY
Ouk70EOeQqesMMuJpHA+4P9s9KXhkRMDhfap+hmvIO/Y3KEpTESg4QUKDC8U2bupTtvqzE4RMQVH
Y6SgLL87QWdqkp4cl2gQ+Ry1eDA61F1DdddDpMnc1Nh3ep7iMv2zpUG8Y64CxUiBQLfxRit7cB0Q
FvEO72pW4NUo9S5olUyr7TTjNWwtUDYh2MzmYy91kZ2QiVpZ424y82/B/LeZmXXmPmddHwNU5CVl
3uYbuvKf1eWnUPbFMO69ay2PQpcKaBqjAmg7uH5cck9jzdBYYKNgrkwIRG08BTWpsFU0DBEB74d3
h5S7l55whyaizjvKQtbN75hciyWH75GnJ7vxM0sREFdApG018ZBut4R2mYvZHb+UVfxUy6M5ZFwj
PtZUw1cPNJ9NlhzUBJJTXNo7toLnrSKU910llm9kr+/T4OdjF/3iZVSMz/Rnyx/gI0WSN0t4Wg+p
atIxUqN9YbYkcYXWXjSYurvMGG6oZ6MM6PxgfAqSrOYCNLpfG6xpSyLIXh6mp+RZ3+HP4uWs4bll
BOtAknrEMdfFNwj3JtLeTRTTjaISQjhDJeOxx+F3XLj/iQ4WoPRq0aeiIOlfQZHmxHWUkUucAvyP
I+oLG/08sGqxmDwwIVqPY+fIinZ345FRqaDHQLA3Vu9cOI0EDX8mFHs108i5d0ftVWHiVWT9Vr4x
BjcEgCIFC6kZbqTcYLBTAzrcMtUVYhSZAjAgwge/wd/s5yIxTgVNI9a/cLuEirGS8bg35XMV0O6R
6LQQkkfxoxpaBsDXVpMU302JG2kKbzlPDcaZitPo87EzZ4z/rNYLv+DrWJm5KDXTh+irsXBtxoy/
Hda1kaNsFd7h8DuW/sz/Kuk8IDxD85DNT5q3q2VNV3KU1CgU01v+3RYPumNSKjyD2M9XWO/MB4Ih
rU1GlwbOc/cO+ajyyyWgJffYaU4DY6ipRr2cBd6ukzN/ZEQV9ej+e//aFHlCgdekyICyJETa4ECw
j04GylE0ymD81t8AijR/6moGC4dcbjifE5uAwlQrJJA5TbIAJF+Fa8RqfjKzM/Vbby+rWjhPNAqw
f+2xXNa0Lue1IoGq8u9M8E4ejSRpAS15jo2acZmNlkMSfEHMzaZXA0D7py1xue+VmO954Hv5BNOu
n7lymnsccTQgCAnyWT4mQHvg+Z3iIIdwfPOdpOhl9Bg5jl69fb0N7fFI7Fv1KcmEbZeQ8UUgx5Ac
EktA45wCfI/T0UnY77ESn8VjS5UXuuxNHUdvjP8mBgj1g+ONOTGqWF6MV3s8mmqSZJQ4EqPd/8UH
fQZXqzSeSeQ9URx1WbVwGCiv3Uu0irozPoVsy5K1KGRs3Pvl05zMrqP3bqQIkpO2ULRyVIQDUEes
iFAAjDCm8DcbMUxomOALUhKU1s5wuWrFelMqtAaXR56Np9lpU597KffyEY4m6fRl1dMJbM/7xBAT
EgVog7tpnSkKA4+x8N0kNZUpEzAkgm2Upm0vLwku1B+bLR6W/NdAWp8fcVHmDQbxtxFcaqReZrKV
E9qazrrYNI6GjcSFtX6flGxCPuxcPcj7btImMBE0fbN99Dkj9/UcEZc/0KPnAeD7JkTyHsN3ikHD
0zliZX9vA17ZqeMyPiRq3YBaKAAbCQ+CJWPXYd08twUNtolj1hqFEXaAhCHAgfzs1qnIsnaad6BO
Ieb8cRbNZfdEJgpuWmeYJvCR1uZFvYbCB0iRM9HbCenftZOmRDH3snXZnHBWI3g7Cnu0hcl3orQ+
IQhAml8yp3Oeo1FUjP8/2K+nEwwNbfUC3IQKsSIbkbmYof8aCze8J/EH78/NlKjOvtChoF68byK6
hvOo0vsGXr0qr2tGQzcjmF9KGfgnZJipCcG81eaxWWQE1Z56vJotmqaCRFMF6zhIeStufiRaOwzj
GOpQ/X/1VxlTv/C2JPmw/+Lt0to2gX5WzE+xMV/qfuTsEJiZwJrW/Jf6yNeI2WmZGgD/yOiRAIX3
P/FMazEEpcmimEcpubC2gDmGjD7bTi8AWSpCbYuAydni6FQFH8nr2YHaCvjuxPl18RuZz8tUnnPi
T9lB/uR6DXlkufJtuyFYu8U6GBcUm489LiB3o3PYUjjrFzbNTubzb+P2u+XGWVr9nEJ9vkWeGGZi
QbK5zvsXFfBlTVJqHBGTtj2UsmsQVJebsKbXC1A3NXKJWZGIPNMAQKRP6/kk4lmpMal0OI812cCp
vldGM/sPmieWchIMwI2A+/gnr6a12bZoCIBb33D1ORA6skz54JG6EKfz3EoF8165eaf35vzUGcqJ
djx2IUmIUvihmuYh4i0ELL4GPT1ba1EpJ2YgjioEC4I41nmLiJRnJQ+wxhFzvLY0zmarr7FYULf5
qjJBLxV0PG7LRdvR5q2mLXWS+B/jCjqPy1T0MnxkuRFPf8rzWrpKxfK3pmXFQtcpMQK33M2kHQWx
NPPRUZOvYRMMvaASS2GAZ7asTfGf8FOWVKknBNrftNsk7+c82WgQyLjWfaDdqL45+zfy+Ju0o/68
kQUy0uVO/eoS6yS0nlAWUS/Ns+IkY1IdECt/J1Bkk09Okoapd6rAAwUi7ztGb1I9yrXh/+ScjyWq
ELwMUPTSsVVb8xj7NQiVaH9sU4ygEePxY409lC1Sm2JyPHGopjZEi+dbdN0TS/kyL8Hgc7hl1U52
C7iX2U1zD+29Ws7umDgehm0UxJSO9nhEZmGFhnU6ZzPah5CGKsqDjt0P8hYfFwhSvTIldtd+ogCg
tA1iQp9OZHMqsyfUbieqip8/QYaPzDPj0eoag6cg32hy0KgugW2pdr/6RNO/Odm9aeT2T3Z4wcm5
UKUd0Y1nMlGJgubx8QB9YBc6C+3pr3NeH1q3dncpbwK8vpyliBYs5ohSw5HqP9VRwLminLV8gcDq
Ecl2HyttgzoryBFPjxn5lzGqYPUsWS1VWH08WF9dw7RtLDUK3Wzur1byfe9nCFRhlrOzUx4uNlIS
BNQT1cwee7dUtac67muwesYo7eCtkk8+Ce6E+X5xuPtmnCV6YsIhbZpCTkdTkQDjZxJdUPqQf3wO
qTuSGv9TIJ2VQIV2XcZOSXm9ZPz0+hsHmUF9BTlKQBbWncNNYihqH8ie8bxeIlYeTDCzDJ3YQgJ2
Eod6YcsL1JEGDgVHQMDjniJY14Dj/eiPW6iZfmWL2CxJmS6zEBvju8mqghi20oxYthHAjY/TGqN8
te4qQJyTKRlfAB4nm0S9Bxv3azhEE0Zz+zmpf0NEQmhx7qLtzJ3BA69E9MaJjsRmZwNWJQiLil7A
WmN3oQRA6Uz/872DRWJFLfmN9lCdP+K9Ax6q/TqHFCzgfYpJ42Z86bBjjmfx7d2z0YwfGQXgk3PK
tppmLCQqhwB4BQFREpVs72DrJfFr982hD8dHN0zKb5b4E/Saar9YSmZsrLqhEbhjMY9GHlsanJO6
xCFxcLukA3Orx+N4odQceOiW1OsNpAa3sz77xn6iQ2HHq9YafPUnRsaSDhQ02EJ4HeOLB1zrTLnm
sZkm7lXc/H7F1aKq4vgtB0kewBO3/wZXyS8t2v+iuHLIeN8I0Q7uZ+3zw6NnuOs34zXPRGWkWcfX
vpG8dpq61VEo80TKt8/JTIZjHMPayEnf7YZrQaSo4KJJ7Ns+9mrwTHirR3uGbSrhV0EvVROruQ0o
X0v3k35rESmEvL4Im6CTadzQkdre/Av5g8ZF/LtIDNSuSkHHF9AopSJmG3KWBEv3Uy2GSjhxevy0
Y1e4Ry9NI2uY1+IF1+FFEXVUENPqozbNa8a5XS9+yr4oe/xC5crfiaYI10HfNUQBE6tjUnQFexBP
DycO2PmfuFqBlEsZ+jU8CBAmDQfEKthoJyWtHycBN6CGSxi1n4SD00ugFGFjRJMDMV2YCjq9IHrA
/hIdpqKyUMqBeikY5jpVT0duEzE++760WrmC7HhVVIakmBzFCaNoA1wqLUadum/cfMImlXRMSvuh
w1UNtyovUyUnhAUr8pRYaFvSaRh/hYF4n9wrCyIZVnfLVMNnaa6J4VmA7uikanldnd1u7iJkE2hc
Ya3MjKtVUiFIwe2SvnmxCdoW9ugymPpzgwq3M1z72KDSMxl0SVmEGb7nkTNjIxFKzMNhxnnTTFoo
OlaxKQW1C/Dob6r1CFIeVo5yZ/IaOvej/3tE9/rSiK+2wU1kLr6eY8hbO5wA8LRJr8LVnXaqgQtW
SBQTchsAMRefyaoSpRnJnkP1kl+sYK6a1c2pE2pWuU9nfRAgIHnuWYZFUtYVBaf/AKesM1bm0Hr6
oGzZcS6HJpu+z12SrXFMHRsa0ER7VPnNDwFkFS80N67Trjy6TKour45SAmQDG3LJMgKJnSTpJ6cb
uczHPtHQ++l0pk4PW+V7/lHcjV6FB6+0AkoQg+CyPLuUPmLIthf7vwylCukLiDNiXqWU5kTuxwtv
D6k8koHbPeJEem7lNNx1+59F9pUa28M+YUFhL1Ytdwj94Qt8cHqk9X+Xlc9BXjQ81y2X6a56qbzy
owfCNrK25ZfGRShYptseM9Nuu1AmUhzoeU9Bo+fPjhGSocRGs5p4JQlWjgR8CUGoSglJPcMPvR/7
VgzvztQLF53PAsxXEFhz0pBh/juxEXYaiWwMkWo4MzV22hSg7z9gef9tGAbgrN9ebEDKcHs6STeY
Mu0vlTYqBKN4KHsaUp8SroFn12IxrkPEHra4CmTmwoLEhpzaHh5cAV0fpwTS8x/87+5qnA9pJVoK
UjEyCkjsTasT7nY4YLQKkGlhjUIxAYHo2eyNwUJ7Xvs4hEzTxRS2aL3lJ0iX12QC2tyb5MsyUFEu
QW5tD6DuDFwr00c/yig1C1ctrE+ZgJSBHDJeW5ZLD8cR0e91L5UQFi4jBzbXOjpZlDYZ6gXh2tAX
SSb+OE4+iDIhilXBT93Of/khkOZQaeohrx+LHADDYcq7wa2eAGglbX0YzZmU7jyYMX4n2CMOUbNg
0UGBuwRtK5d6DgGRD3s2w+/CKwRhUAyVG941e7eyxg0qqF/idresq+pOG+pxHRkX1QEClYm+8/U6
OIuxT7UF9vRgv69eCnKLM1cBt+HE38cYSf053GMaFuLF2cWhG0/K45UV+k/SpfUWhbN5YOm56eev
/iVEDoUEaLZUgsTjzaW67bgUiSyEdToX7KeYskuYquo4fwgCK1SfjN3xWotFB9jZmskRia6TCIC1
dY2Ws43T3doNTLK8TgNkOsbuwwRhJuplVavhxAYthIA8Yv9HQcJEmVgfOykDAjPnqKVD+CRBvoQH
KXv+5P6eDHgFlVrt5nqpdMd10vU36S5qQvy2VdXrjvSbWlSNxAhg3i2JRp07ruPOfcTZXolMHBa+
ji/2QorGoaQAQlwH9dhqorNthgEd9c/jpEdfAhD04iHXuBiq3aXIJNJl7yy8a+6ww+xfznLuWdv/
Wk7b8VBOeDElVFS6hKNRQI2WkzF5CIZEBq0wGad+t+j2z7CGcA/MBM/cfCPG2T+hemYEQ5kF2mBe
kxrQvj1o2zf9F1fLCvIEjgb34F7emO3EZoRAX1k1hFFXEDC6bg3/D7+iCNWZzHykk/QILbyM8rPA
Npn6X8mw8wn6HjdI4yr1PSkqWoY6+j8ONLgFGTFrWEYdRLXrClH6fp2SN//YeJE0L9iqHOiAC4uA
zAw8793I1VlaCbniyrmX4PEYuCMWKfmyF6lmT+VfP1p0oAxjNagJ6xKDUndZt1NWsVxmO706tSZA
tfl/Jpx4DDNxiER3IpYQMMkdDIT44HEwhXi093L9PADzflFPNPWq34fovriNyIwmDk6T3oUy2kgS
fqMg8q1oON/jfHFbpQgy1iQCjHw2imYdmHoPYG9nrr3b95BtFEQBbypX1FX3GoePe8FlP/oPEjmU
H36VyAEOFVm4BM+Ay7Mpoi/EIUH+FJ9OIAgOV5RqYhhkln5HHy0CEb3mbB8r1eTsKrdiLwy15NlT
NgloZKABwpl0SFowO4jeKkfNOE3S9TRS7kJr0Nc5O/UpwW8himz+0VuBJKvsdU+lsfRoi7O3NjC6
W7DrE1agxobdObf8I9DqRgf9XJVX3MIs9//L7GQopJUurdrMs7WsxDn72u6fFEJgyw/e+JRzlIAJ
GK8BFoxMIpDHzu5gwfqrG8UmvbBQdki8x1fyIwlUmWn5T65zeQdpGZovxNNwS58XS+PqvdKpbg+0
Fj9YMJlv6Fd8ExkjlucV+Ik1oh0MFaQZiLx+4t8XXaSgYHAtDYzzxUrh3puAoLo8nZcl4iyaL0U3
/ZftY8xdK2rl2MWSCYUuV6PmBoMOTSH6FKq1m8++FEeCW5D85CO4jwBE2zKKs5WXxHY+Lv9xbbvr
qfdZi20BLFkLTvHMhKNXPBElY5IefmB3MDVvHxzZVGw9UW9/Sb0xN8afYqwMEX+MObaWpL2dHi59
Awd4sLFKMNAAlVe0w7e+6gR46bRyE5xdwKfjWkSPE/jAtavNZjkerXhFSQ6cnLe3vRPMRdCttghX
NF3Mc2siMGNT7xLcLc4KowzY+enjSBn/5Y2lZGNTWC2zKzSaMlwP3z5kUr/fXyuzxVfHpouTYtC/
ekEsCRdmHuhaztYKJs6e/Dk9KVGAdYVt865z0xxaLcF3fsO+J/Y5PzNBmV/VtV0zvQ4oU1XkBlpj
8ghfak/bJLl2giFW16HLi0lkenXAolI9240Bt4tNio6r/S+QFghOw3VGk67an+6Jk3zHhae9EQ6D
wYMN67rS+SDkY5lYIuomToTGiXURkKUEl+HgpGTxuRz6qjFo/eKq3Tj0X3PIy4h2vnvaDhDSAWhJ
ayo7EZVhAXTZBHft0y4HtcCcluts9DiG5fmA2dYKE2Oud4jevt4Js9bSZP1efwIMFtbhvfyzLL67
O6AETZUYjA1oibLTbPBjwmDzgq+12C/T5qRKB0LCJ7sXz4uXiixAJ0JIz/QPxvzcDl67UMVHxhSg
fvz5C9Oqn/A3SjTsPW/fM3ANstJyGhpMy5oukUfuyolEQUvI5pyvTnt18b5jSihTxiUZ4Tn3da9R
HmheR3ggeSBKbVeqVtTBEz3t8TjVy3jVPzr+B839NJI9Sk2rje8d2aazfbOszcGwAyNVDx2vnMA9
y6Zo/cLxToAy17VZ+vDQYIGgFMSvWJlAfNyhhKyAJk/7hi+zxjAS4Fv1NB+m+96gAVi7ICORYw0E
tog6tNFfGLvQT4YT/wRujG0WDjCE2r/0EZ454Qtf/m/4nheGUiMI6mgP3SDDSElHbj1mu2zI3oo5
0NUqO6tedmH2UGfyWOGE9DCKwnnKcSWyudvWydbhbVKMSai9VqjDz8iNOZijnsuPzEbPyuRp2Qz7
T1Ej86naIpKPrkS1ymVmz4UKCWgCHqC25zZPYaAKF43jGYYIBOcM7YZtQFcAeN91lxyGz+Vx9AEN
50ghyoPqU6Wx+CTYeC32Q0guXnUKVdvkJzUcKcbSXE7iT5cU3gRK3VTp7EgxU9cHRH5IYeUbzbfK
WThXLueGDMO0V17D64x58wG7YI2dJlV6eE087bMFGTiUiTv23DsmJsCuHxlsCRKBAyWpBwine1Ln
zqyYT94Kkt3CdAhFYtH00QgJgpASP0I7y9zofuSXqluO+7E0paP1rCKJhpoy79D+ACwdKck07ZtV
oEy4qFN3jkzCOEvgD0r6EJcKuQT7k1sXPc41jlKL40ig06lgVSRcePFgX4WmTEmnLlkwzFj5yYci
GX83gW0fYmXakvHDGoQlvCiGYc1M1AxIPSQHpTT/JhK9zKM7gq2pAW5LsaeOhoz0/XYZcObVjuAl
A/Kn97lfivMPecwYIA1BXyWWLMpvpwBL1jAZZZ0xv3VebapoLE0eE/0JiyXs7rRZmJxmjNCqyr5R
wTqfEbB/I8PxnStpRYKOePJmui3uYcYZOqoqp6nmB0IIGVuDFCRC85se9FtCrj6/JvLYr/xBu3qb
DmyzbALGNFa5tgX/j2UrAnQWtlP7jXJkW5JHtneYTPMu1fGcU3Z27g+RW4qxziHoH/miq922e783
iZM4DcISkmD475GIiiiSxNpWnl/1RaNUWSKPLAiMUS/KB8L6nrdOSwpD83ogw5vBuiq493ceCKDO
5d4sXIAgFvngycos2fOrJuNWvG3MSYKmmaxifM01fmHJ/J5Ej/82kPkmK1TBEyosV0dgDdDCWgiU
AiVX9qVOxrPahNaOkEluk8MvlqKfBtNXqJayuCAyQfajRXoK229YfkbBCgM3aFBlkz8O9UJ22bsF
4N8S4RS9H4x06uOn/QaHgBf7oPqM2sSwTdCyzmqv8Yrg0S7OY93rkMZAwNYq7hYOImhRbNUrqAuz
G0jeubByvd4LWDEX988M/TjeXLTx8catrmMGpcOOHlNVT69bYdCvGyldmTVboDGIOV9cybLyeVCp
I8XlBEHLVlcyvD5D2uifeoFa/nlc5afAz8BUNLQwYZxRP8aUSrpU68Q+q8bxfX9MxaHeLdqeDcnZ
5453Vdo7TGGBvVuBmlMVMwqCBR7k6miCFnvuxpOzIDJ+sfWIEWyzgrA5UgdCo3brmbhvmk2dPecy
dniP+7e0c3Ns2GPN4PZkunV659wwVrFq8rBs+1Nh3Nd4nGb59voPtsmKCLolXiZwF+X7xMoNAfsA
zscptlt1z+YeBHOJdsnAWE3lw8U2yVJvF9ypbPK7O2GNClnTvJLgfGg7sl0/b5rHy5lp2XXpZx3d
WvFcRVyIOw0p5xlF9pDzJPC0+8JLI1MX+6QT6t16qcqcOxapnVhj+rtInQ1d4176iqjjRWXrPExb
t/jZBg3Hb9f5TUdo7WmMtRQaGK+yNyNWipm0tQGKKgqGTjtJHge9p4SytvGfDTYf0n6+PjuEUhoq
yv2H+JkGwKwr1l+R4j6JDJECFy+jGa2Aj4SU/j5ZNc0dn0WV5c5jQkrLHECQ14qdT5NR/MqjmwLd
Q45qsVP7f3KeJMGhjorrM7ntpJzoGr9fD0j2HzFdecyTLWOsda+bmR21I6SfFU7dHwRYphFQtk1O
bzloi32hBCGM2l+r7kVng8S+ewHhg2Yao3sCPZmfNtt5zCPfS1IBv4LBxkeI1Yo99Z2nEHaChGPB
Ttjnl9m7sEazfbG3wP8ptyMeUL0cM2Lox0phVg/mmzqVEFmoi0dBZ0vCHRtJj9Vq9M1OM0nH52kW
gs1cX8tdGsOURnbEJjSs2A0OtD6Jlnf7vW6kfugy6TSDNjwCF8W9V6ViKfcwhoyZDrXbIdBn9H7Q
xI4UxfgGCppe55nhcRBgja4OglYTzvWRRueTSIwWiy3qU0ZQhQstcPBv1Zu1Xb1SxD+BIwdKIne7
L/7hvrQFHEfeOzH0HiA7F6rxicyi2ol7cybEVu1qzccAfuHByuYvBDbyr9s1J4k2Pzqg5PvSBQaD
/qN5ggMYeuQ43MkVa4CHOGhKOmf6JBXJps1kEO32+pvAklCONlcT4L1qdUIWoACTjuQ2BpEQamy4
eA69+iBQ/EdDTP4ODUKzc+lDaLZH9fs7g4mLgwaZFdsw3NNLRkgmKfobAM+lAF5ZBs+b1OR0iBmH
Umsgl/FODVXZCXV9Leuhm2TmDDnIOeuGIfadeNm/X88XRkOZ+CtR2zvofjJlNydrnSgEIaohVAv2
2OT/bdh0jVMkhXfoPl4AY7yA8/a6qXgCvJofhDn+v0wshcDKVZm3IGj0og9KI2upUm1YMvnsiqbJ
pSxPJ+T4Hwra9RT+Ura/i28kWXH3Gg+IbkACsKyKr/EQkHc56xdr4dEnij2WVP2Y4RslHY/T4oPM
cxVv1aMbY5A9myvD+N0RFR3rfdSB2WCKgpLzo/JEVYF5pYmAjDChc6CHdlywu4Xf8XzWqMVqiHzf
7zwneuKVR6nNYOUNcotJtgwmYG6SfvJAPEBuxXRSnGYQ/azGyBji2hpvEIexZGZ98379HSWtMNOB
sXSnEYq6787+inxuY2O+9fkO/I80tbqCYW/sHZkfwchWKQTlUuYzVAd2NL38p3HD2DJAeOtnkq3O
nu5Wb/+1cS5nsKFBl41ykFg1O/wvRHlAqBmAbcM51V/pN0MT10RVjXTlBScw0TOqkiAyGqIou0K2
iaKd3nW7wcvPjbKCmoadVIwxbzGH6pof9ZbLVXkidYXz1FkFWwsyvCYc96U8rJvL1ifLClW2pmCq
3/bO+h0rTuuaQaQinFhSFfyL2DE2XHGwGh6n3i+9aSpxKQSho9Q0hGgqMs57uhGs3pN3QTB6NyOQ
NqZujjrlTSxlLSOmkGcrUiwjadJdghHDTbNXPANcvj+fv7fFmB2Xl4+6lpIEQH2Jnjfk7YTfcf/z
ARzfuLakpBDjg+rHDzrql6ZCYk/npKk6JTd71tkw4BxPjj0sNbGO0eBh+AQARkhhcD2Bz29iFq1w
u/ey+KMqxRZgZWtKGMtNBW0ixDQCcbLLWsafXYMKbmll9tYMqcHwJJn2NcLADosUdGiYfGXPVb4u
+nsfJjPHUcS9NiV9/uxcl7QqSGffSfpOserTRJXi9tnR8MUmeNjPr74tEMnWXNNKklb34nLa2OP0
9paE7MTQp2btrLVhuT0jGmKNvibORvwNCWGYbqt09YkaPK+X0MWIiYnX3HDUlEqkc1CNxXPviy18
FhkoBlVWAhuErwOTT7gEBzhS/NeAmwhYYRjtbwr0Nm2LParDLHazf8BfPl6tlY0/P708Ieshz5q1
LRHIkcouaoh4p3b+DaVPK5scfJ+4ZZj0jD2ctaFsxXcT8wNaJif5VhJPx4ulw8Um3v12E7EnWazY
ZaRnHnTPfMNm/7lncqbb3PM/cpzlQDO6rRalcJofCsaWZHU6nfOgMEotgEaB4pSWfKNjZceBLWEz
8Bt+pQJ8mFsglfp8GFpEWR2pAQNDl4WphWU4fUdsY7WJmlo8F9QtnIPtXH0aJ8oCOBXkJMHwy1jC
b6B3CcZBpf4AJXWD7y9Y8bWN5kOzzSnoHyoFnQZB3hjGvLH+mW0PaxgzIU5QvgCoLSz25K8FRKrU
aPAUFK5jx8vJkBcz2mJ5R4xuIlLUZqT5Pr9hctMdcLjlBYsNc5gEnbDiroKQU1XXQsvNDkwezbda
hW7mZ2zGucFNsrCAKFVUtWKxzVVdkquJpKb572UvPHUYyFEFHx3StChIV6Mjh07N4Mfi+ZaxvFvN
NOiVu5CY2Osqeu6c4nn+Ax+WMISGbz67GpRqCi1SNarUrey4qYcg3bX9q62R3jIqAU1d1ZLoH12k
6iuPdC8bts3SUXafFPRZwkfsjXRH+cvliFRbeX40UYXx1E1XDQvZFk5oWdvR873RC0Z0cg3jkAyg
+Qgj72MpP6Pb0qqIb+ngnaHNxAH4twmhl15LlI44a3/e8lzUgLQVMQV+mtLZhuZT3bG9if0+LhC4
tO80EGMlCgFsz1EcIy1EFanJ4HV2ZFaPih8IW2LLIOdr8aTHBCkqTXnM9vneCVraZGwc0Ws6/Yy3
lS7mJu2EH7HnyPm5q90P810nHgAaLbpB3PKvJycstQXhVwZlN2q56u9tmhAxQvND/Eb2Iohg8IMr
vJhYsYsvsq/Oj1h3KuWY/4HjeBPmMUwmHuMjL5CGgz8ga/dxjPMXeNkJ98yWtp20K5gJBaLsiIZf
o92qX19qF0P4HyiJ5oX9+5PBrwmKcWIiU5uDpBLiaGPT+aQAZJwKXqqSGhe09e+zR0VjlAHoNNPJ
2Unf44qPxW3QMUQG9kzP4RjcepRxrTp8JXo8Dwc03L1AqgrpRqDVgjz8mJ/kTwnJwVaKXqK9iRXi
xmsn2vN90Id3VP4w35ebRcCzdVu8qwh4OmVGzj0q/ztgNuamcSeks4MRcL+axkU+SJVTAQ0IIPIU
uD00XdyBqAwaHzWLhhLNMaT/MJx3epaTq2peIClXYzgqScu7S3JsTXI1Rk8B6dBnSjJRpiEbS60Q
Deq1sTCkAoQFXDKTjykj6ltjynj7XBNN5/FVWZPyTam0tp0zKBCGbmhYzB2xEyjj0Yh5j7KPPA3f
7HkwIbLM6BafOkqosYPiA/BAQEZveZzxWMQUJEQj56KMcK+jP9NCM3rmVdZ8JddOn5BFwIm0X516
Tfl0VqsGcifXBtsWkbGA8E/61GSMlvETm+wHvYSuosUoysS1P1EjAL2VsRzXa6GEEkSi09XdP1QK
maxeCesSevQvZp6uoLiMY/+qP3qwZou9Qjs7cU/SLPptZQ/mEPYVPz2FBAxCe++vsBaWWFFA7MH/
j8Z8mcVrHr9aMH49v1crdcOwuyUsxDq8SbBfPco0gKqysN/OpP/OVh+NH8u6X0uZOExzEvr3umPB
duwafChIiEBCl+4MwR8kstY/ZGEShgBq7gMGuUnUB3dlwYTEUpa/KDeluma7k5hIMqx+KxrYTxgr
6+NguxqZ8L8QIkbsdX9d5RzJi/T0aM4/MSNU28+T5a1qc0HRaypiWkUkNLN8rnADo/pN94Qri5A+
5BDrHLZ0qF49b7Jt+YXa+eDQh3zLd5WKjSynM39I+FDG8rZLWiyf5YZZWMbsDDn79z8YzKgCkBXr
Y/7GLTzUATeMdiXpmkl6IzNDkjNs23ArzTRbxwxK8pWJ2F6cJuXHfLCC9oDoXB1uB5zU6JtoTbY4
Bm0/1UIvykQEH7oxG8PTCzexZ8UZXfvNDEW1JpFP34P99+8pBBUzwXNsUt1RuWmS5BJN5X9VOF1/
k1Vihcb5pTPk0+20env4GxvILoDlCm/IfzACNvGWH5toFMTjzUh1DmHYEJtfT2/9Pc8PduyJOEHu
CUI0Sg2BCTeBC+hLNTONcS5adECHvb+8RbZYGxT7BW2BxuxugxviOIasDl4ASJ+FzRiNkTLMUFBi
FQ+rUvFTLzPmK8+Lw/fzMvO3q0IOd57v/wZHrH2GX7arzjSDpFN/cnqAel0d4TXXPTkFFgJfoK+9
QWA8VElrIxDNg/TSlg6sPSmiSfk8INPrY0dreisDZRuKTPHRGVr3jf+rL/UvZuoKOH0+zF0DdZOv
f5lFl7yzhanVJNpuk3F3Wb3+Q956m1nZ6JqybCkG/iJk7jGmwphp+GWY2xIY56jwrreUi8hSWGfH
vwjwnGtBtX449Df6hXmNWOJKle/Xsr/LAjQo2y2aWjgoo3Rq8t9RMANez0pD6ugJF4OzUwtHinL5
GdZh0qgY3LlZ7PVQsN0EKUZF9DQ4gObudXR+lrCOXHU50r5zG1SFlv3/JBjr3Nrnsajl4A5DyerX
y1Xk5FFvtNfifE2zrvqJgRUt4NiAh4McI93RAS5cSlDJW8ZCEM0Usy3Up4YoS15TpxdD6iRgqr6B
tj/2YVrjIB/Nh0Z10tkp1a02QJeANiQPn7KTQhZdNz0nbsJyObsGgz/tmwpZZLSyzRXbQqO9vebm
QLzGhIxqfNsPyjiZdbHFWwodFaDzsCwA7H6iNuWQTUh6OA5/fdymhNXSS2XW/GBeGLQ0LAAsEg6C
MaMBJ4Z9bifXzue+mPt7wWMffFk5J7jBz43vXyHTp3I84kgsx/eWv49NyHB7csAqYZiB3ofW5wwE
nr1KTQ58pqnjLVoS6iYq1TzKx53zOp+3UGJzhP9bti7+hcaMgVariGrboUiLXFdMd5aq8jLSa/Jk
6YXP85NNu7I0sIqKdtB3OVOj/bulJEdBi0O0miWBoJV211g3cNyGKL84/KDrQu44h86CpPNJqoQa
ZbeVzExiNzXhpVJllEqHRtrkf/FXWx6H8KBj1c4+wogncigxAPLNKBDD0Q0lqwb5GCAcOPeusJVs
/MzirkkjtnvHpaglbIzjxeMN0Bep1rRBuaiQqpG9AVd/0Ny9c67+l6Bhzwt3U5j0sXWhH7qwSB98
9STJSh/fejikWPz6bKs3lIEoKhPghKCExTQ/b8tpazBjdGfc92ci1h4PdMEaWxwo0FmSEyzJevSw
NrUj1DvRkAPwsUuJTI+wgXtvmBFEn9w891GjjHtXPhIAueSHUwuz2ODl6NORjUe6KAR8sXXEyHZ9
/fptgEPz5q5C1Zty75zJD8PqhFSHRyRcdOzHXSxJC/CPxnf4bZxa1OrgV/l4xz+m2Z4TiskJfs0i
qrtx1Zp1WAnDqctP5U32cwebZ98rJe1qVTWIzo8N4yn6Ui+VrVuImRiGAvFbrMnL87iXUVg3rvUz
hBx75RsQA916n/BEmDIxJ+k+fgvUOSQ02LJ9DNxUfG+LiIG3d2taRa2DxLPFJpLTBCpZL2MH0uaN
CHGfUmtaI9ySZ8kYnc/cAIMvof3uGHnYh4qbFm9lZYVAjSIOiBe60QLFKniqePOGVRvx7LI1af2z
ZqwL3eEQgf3rvKrrZwkWDFm1cpMOba06WfkBLLPuXZ6MFLUZp+GdZJPJXUO4Lm84nciNG+OvEvEF
fdBMFebKVlccAULYFvMJYzQ6XiDrASF7GuDn03jwax3RJzfiTptmKm3gUJkZnGHRr/pCZHamKssO
RlaN32cuNFEI+ofT9qsN3QNBO+giI/BradbErk5DMGVIEsgB2sOR8DedfwUolM8jJyetE91n1+G8
R9e5JAK1BAe2rHnIVfpTD6hIPMG/GvfPge9wQEhgdttrFCmvHfRWNrjjsQquyYqN6hVH3pKM1o4x
6LXKrz2aY8BuwEiNfO9ivSzDsFsGgheKS1Kwlp492YofzIrh3TxkPcC4CiAPZSL30+0511dF/wR3
FyUd3XBXVQ3Lt5P8xdYTE/cG0Fvd84+03SVidgVGi+ogBtK7n7wogJ/5iUlCJZODl5JOj45HExj6
oLyKi9OTQ24MSEb0O73rcG+o6DY0bevGDpV9HHjIbMGYUPARHTYp33PBT9Dr15y/pDr00OFdWK2/
VP6v2eZK4PXyhodJqzpGwbsM+lEW99rFHKGKMfOYlojatexQ1aZupngt47hMhW7zH6SOJoAMYdFF
KAt1dzZDd9GJz/X4+da7mpYNuD1ooNOBiuzIdQaF3Zzfeillv01kTFnzG1FssB7qhHSW6ZdhC/F+
rELsl9XH0UnWOmTIRIYYVP1ubCg1ZnSqXbvNE/V8Typ0iM0kx1m1tj51bCGfgO6NxJwluxN4BYHw
m2Zq8vhLw2Z9+pa3h25LcjMC5ECA2zsSsIgm/QZR5dIeYXCfP2lJAnA9JZda79re2dIs8Vm9otEl
9cCLJURW4ein9W31+ZYreFs1lcDN84n88Z8v4z9k3BqiFK8TO5MchIuqjXvd6EZid5h7vFgHdraP
BbV5PaCP7lPyBJN5Y1VdTkQlnjTf7kgLxSA+D4dMQOWbJZXCHj5n9Snvpm1Zp8VAcvbtdPawsPCx
IzYtxckJ/b6ppKzHitXCq14BdsxeEv25Kc2LV0Fgp0TgtAVjDA0BAWufVEzW5orqrZaq9pkyAMuU
py+dufLn01TPRVqAI8Er0pHz0zymKhok0LKuD42GHRQSy8uk94N2bbMwWJOBtFu+U9MmrEhTnfnQ
MzOLjdZ7mYOnyD32ASoV0moKiqNTmrlxsJTbOze7UkknXE0JSpNRzpHQWpZZHPJVN4WL4TB1RUpk
r8ja0Szbx0ZywABxYRAllhQcfKS5dRoCcs/hw8tU/iWayl5c4zgs9vrtYlbFwnAvGGRkioYIKMQS
Hhi+r4AYRUdQ4YGtUM9mYlYY+XDtifFImsu5X1twBPcKQvewGG9T5SBPUav2dyzuThRxPH5h85e9
6v0+i/IdJblix6X0H5zqETwWPvzR6AF0o/xqHG3yX48+Tig+j0jZg0WvUrYJE+wJ369uh3AdrPf7
TEMxx5MbGDQZPHSF+RGsa3p/JUmZzVTLvPuC0fPgesS5SJcSnat2GN93x1ZXNQM38LNFVhKKaF6U
mVJtwuA0PfaPKO5ZPn5R0dt0dhBPcWd7jsERmzlarvw58Q69moYYULgPXG3IeoW6wN0kcpYTUie2
rq+Hyy9x4fNoyqZ9RM6j8VqoLCdh87x+jsrFWmZ7Ic5/gf2mjVcO82ugGvc62rdP3ncQrjvDM7Bg
ccmzA+UUvOYcOwxBo28uKbmeHMxqS66/gnkCO9pWQ1cfaGZJfKgMx/PhX9DI3rUhBkxoJYpqBUEh
O9vIEJTRYwQDehux3jQw2EqYe26NfkVEjuDM5lB33b6i/8V6+IOycj7NhXIg4kL7UpRc54V/EsAO
pflcBL7aOqaG4imTsxhFAHW/ld2CzObHvK1kD8biMoKm5stM8gcIDxmkdw5qpaJFtb1QQZEiCr+o
fQdC/ZjFff5J/G8Kq3lLgLKCe1I3sats3VTQoQ04z5SwpL4WXaiixO8YuI5UDs+GoyFz4/Z/XoUk
st7xGCVD9bESLKZ4zWvjI3UEX5/0UJJjaRZXrnANPrnaKL3+fRD3SfptLb24xqGWOoe+FFLQWnDN
GSwauZek/em2ZQ/lB9B2B8kdDGCpT4v4C2yWbreUlUMQFSc54zuXjo1hDWbIn/InGND3HOLcuKuN
AO1cKX9RKhnFYhq36PR/BQMXHeRv/4JSMyV85Rha+QIAbCMXwflJTH4vhtlMZZD7sVMdELlwFaK4
4A3VxDCp9ae1cWH8Z/D2gxRCurihISlLCCLKbbb4FY/zFNqvxh7xa7KuJ3nuwSEQovbFZ8wzzAPc
b6Db8kuKzgpEsLZyDimW7p8IluDvOsltjBuiBUMmsl9BgC+mnrHdKmTwmO7iZcLfw9hw44UevFM1
/8liPaGVE10LBc/yMijdQDaonTPdrzLL2fSXhQTcaMR7nQvfL4xXOa6U2c7jCH+05RCsQCrCPO4R
WoAaLeMy3mbUmBVI5lyB8nnLWDlag/6L7my3qbPJ/ch6wM0Gy9AabaPPSRX6k2J0l5UKtwEpQaWg
lU51wQXDQlVP6rMoFwYvRza2KoQuj0NS0FIyA54gOa4tQ3+g9F7SVqoZRuOkcHZD2sApy1QanLIJ
SdU7uYLHEi/gxNJbOoRlWOWkZpRAfoiubEvTINkUbhRrbFtsLZSthA5SAmF6SIATikuK7IElLprC
vnC20XKqGcy4534FASCS2a2FeqGQeKKX4eM9h9toxZmvFsmMonRJaHSVzyRE1O0wuZzCOnL8LWR8
Et3r9NqdqCgdkdVMK613WQ2TsWJHhiWZ4gWkA4U87pEO0E2ZD9FWyuWLcWvS+xQrUIp9U+sgx0wA
B9IObsdm4TdNEmLstiMf14p2p1/5VTILBW/UQJbl0siB1749VMqgdKBCUDtNqAdF+uYWqwRSg+9v
kWVV6U1s1cJuDCiNb8ny/92qbZhi2C9svyzYpkx38o86DDHn+U3rebKbFb54B4COR878wQePD5HX
0m+XSOtV3DpwP7uWoWtLBMeHMTHG6yJw9Rx9w8vQgF6chg/1hVzlcH1/LNxTrRI10rz+DBnsI3fJ
3Oj4hfJUzQPebRfkq/ojHdZTjUVRryPXzwskMqa35DLvs09rxAhZn/v/t9EvlPQSpP5KutRcEMaH
HONCC89qBsc+xYwK77atdXfgSc7ej9NOh3p4I9Lls7Ci/gfGju2mcHhnbNJeE1POkOjXWjCm6Fea
5so27wXTREoOHNuJPiki3xWjOkClgQOLtygOBQVzcRtPmkgD/vM+9njf9UYdnhzf0lQTFJWAxqg7
1idCgj8vrVXQhInvlPHLUfeoOxepjbjU8Ye1oGV13sAJECZgme+AjQm6BIcYWpNhyUe/1yJfcGEs
fDf3rR/HbcXkwICMnjWFAsOzeALhUQR9oFJoasPZuuxVSvb2gOYEC93xawdodt0ddOun23IdoSM3
HALQ5qehrgXrhpwf1azrOHDig0HJdK4L7oEH8bgzB9nLNTxpO+PL3wSaWA7CKTn4+CbPuOy2/bvQ
EOSbK6UL184fwAP+NBsdTpcHoHdzMNZx25pFDoTYcCU57TVlLwXbw8sXDB1CE+62FqHUDf6lYJJL
lo80AqkhIMgL+fyfsUmLQihq4BCT0KjX0xqNlPPshsXwF45x+lUO2TZuewYmVDHpI9XKAi/N96iI
Tl+uylhJ+xGk9iLdvOQhU+GfqDVQdqV/9GS/P+wgE/renB4LtOaruxhj6GfzR/DIYY1xyasNZn9j
CEqO1xGqBymUaJIOY1IX7zDLbUnJuEH2Sf/R3UrqKCPt0AebY3iUT631jQzp7ror+e0EymfZ82bn
wOJqA31LhyCV4ZyILIqcBejWGe63V+to4OwRNfV2nk1c5wGB+cvQ7TdiwwgiUTfJ8o6zyys7Mp89
7gyccEqyzJq7fvflM+uMVfKKRQKEPAj1b0RZpjouEal9Gc4USPVT2ntU9wpHXlId9MhXEIXklKzS
x14qzG8DjpoVlcg+w0gZ3Doa2aAVDzBOLF+/9iZPmauev0Zuk5GaJS7B86VOcrKb75uL5QnyOPy4
xXTH4ct8ub7vzrHtTn08cFMV2mrzba37cZyomiFQg9CJneHW0N38IqE6N47XT7G05j1/wvsC1puX
lSZPas2Jjaff7SGaz+9Ubq9nun3oiw8XioX148QSIFabnvLI2N9dr5hO8j6YtjfIJ6QIHoJRN4Dv
SfFQeiDlba7SYGxkowUnnPfA+XObfr6d9+TU/CjDixuaGSjXsARsoFC64VvhptSTPdqb3gflhif5
hpIokt0EqZhhmjhIhhnwjlUznZF9dJLAPSxVBMu/vfavxzgps2JOuoAWe1gUjU+iDsPUSWMkkjKx
MaedxgE5T/lnQkwjIhFfTeikE1Q/TejZrTd6YgpmTGOI6q+cP5T2B3DiRyJ1hegTONA5GKvAx+8V
ySwdeGTlPtjv6khRoIEOocd5gYzWlBirtkkSuNOFy61BKN4DYHBcuwzEvt/I7DhFANUo+N2LTSn+
mRKe1LH2Xsn7GCBw+hjV0WFCgwtQcWwb6zmMC42AehkTykDSs/Z0b9/ATVbtkbEsCvIzqyHFqU5p
sIhsOKDym/EbSjYjPpHznULkX85DGTHCdFouoTLyegOZKU7ADFaMLBvgyksXXsqNoS12m7MlxGTS
iG9qOLXD+QOaDQPtFfewxqueRR/J2dJFPrG3w0+Y6tp+tV6f/J/BTcM4qeIClMlbccHWnkJ8cczE
Kwg2J5ZqwB/OC+8SHCc3nF4zPiAlCZC800jQKtcLqX48mmKoBtPchEW+qPoa662b3K2jQIYkIX1p
L2c05ODe104xM5CR9igAan/KJJSOtc4ZqIW/QNxrXsAGSsTs0XqhpaBucSA9uavxA23EghNKiNG/
aHbK62p4zuvsc2PAinaqvnsl3/pbzbi0vjoA00dfvZXRtp/2If+aW9hstaAXd++f2eGuEdtFiHQS
WWJ/vsXBfoYRoWKVjCrZGLp3xxU7BBQvTK4krvovTEwyEkNg1QrloZsGB+bbE8sv9pFuufuj+agG
wCD+Knun/yE/o9LK17dEoyqjfhPCjM0lFeb9Qf7/E1/vXq0d03VuP3M7dgpqM+MN1hDmyTaQkuuj
Y83qgP4gmSbkkXUfb+RFCb/SmaQ4yGrTR+rzLebCvOuzw+cCndEJ8mqYa4GbMr6ojKEWKNpv/jdh
HpylVi6guVS75vVn+/e9af6sxyNpNHLPSMs4LLsuB1+Nvh+iR032xsDpGh9UrK3qwTcr2E/e1P7Z
YhpF1ZnHSGYjtf5pzZpM925vJW1zW6doF9Jl8RhA1LJGiJdeHvlv7230vdInL0zS3d4gCVx6mDOm
1DHVma9sAwR0oqDu/RxL07SthEPB0NoTdZgWrM0q5j0jfQ5nwkhHwhFzQTbroNwP1BuMc1a69Aj9
uv62wcMOwUvpgEoDDIE7y1hU/Wp9n1QXz+t6FvMrSqWkZQj7JU7JS/IvJkR+pDsu2MNH3Vcvjoqz
W6BBO5lWzyEmIkOOBcgHOli92LKDKGj1lKWtNptN27m2U+n0Ovr27g8XA0Pue4KxlV5+SMVnMeiD
gQzMkrdRya3nes3/lLiikGfDey7Qr6Zp0TpWIar0qdId9C2MihkI428KFIAFIBTvbDHbpu+WgcpL
zrl7rBDj5FQKoBdM6ycm5aa7H9QnhdpCbthRBgp7uSA+q4z21gfoYQ2nchVd5I9IAKonxMjz+SEY
HRYzg+LkndgrmiQ43a5VCie5jkCrlDjW5W+mKVSph4vU4w0+eCPnfRW3Az029s0T8NUDbxcSS/RF
1NQgCN4Io5Xg4dvjWA7veyGnhQaKImt72b9JA1xyW5fF/qSwChkMHW3NeKm11IFIZjf627mIrn1k
gCKhDIDsZMTBNeSlKDCkyKtIIIfqilE/WwL+HpN0LxhJEuHpKb9T/bczT1wDFdFy2jqtoa4XPiyo
4pvMOf8RLMq7H7fHXdnrfTuqgx4N0Zlpt6fh/I3sBLoLtlm6gW2x8UPnvcwNoZkH9LN0tMRM56Yc
Eg3aKSfXjVvWoA9tGuztizL+nXXKLQ4p5fstpBu5A6N5TmiqMc3E5YBsedY9jBxpuquCa0cRemTg
lzZcrlj0+l60LIK4rSHRgzqUgT/j4wD7UnJrRwThop5dM5tHg9uZH1RLXBTU7CKdajnkEyn6AUe4
GZ5DcLR+rjP9ATOGAgP5KWUmj5AynCN70Rs9BLYorM00o++9Wma1mO0rX4u+6KcWvn4+5X3+WH61
w8jmwr3i0Ucq9HYTeZF64GNSCbDk5WVVq7jug5maS4i0PCrmkH80pGS6IUwHKR3R/CdTP5BY3nJZ
zj6zjOqTJxlWbKEYO9zkE6URnL+ZaDZX9DeUtKi583nws5GERx6Pg2oZ0AmyJ+Q7iMaw6Rj+M9Wf
HUyhFXguYrNTm5y9nIsMFeslBxEIGtS7I3E+zN5FAw9C3Fqior5JEp1tGG5ILbiCE04kFE0B/GPA
j4UBTCpjCmbAeQKuoE6gT3NnSF8j3oU/6OTY/sJm5OT+mpsLq6wPXejMsel6fu5O2S0B6R5asaKb
4kMIiJgC2VC+/Ro5iMo4PuN4w8HrqPWKmZ2OhJlmeBz88Za1Oyv3IyBJtn/vbP9CaBCfrarg+Yze
ZiWKiuHldVWzEovX7mC3/73/BQoDI7MJ6++iMPR9Mp1Zp7QVP4I/22NOpANp/9wtfc7hZ8rnRnem
f6OaPtVtiPo0m/xADZwmKRnlRkXVJwtAjt3N+fp7uNkFj2V9gCcnzfmk68Lvzx5NrhgX9lwbI399
uEf0VUrfZwXCJ9XzQ4VUFFTvsFspXnFYQmmATKxeGQLuxYyxOl1pFkJSd15D9sD95w3jfXMJnES+
RwIrf4G27IpJErlAS1hebL106VjxZ3XgQSNWm8yTcybzPgp572TKMNFau7vgJRVqsD0PzjHgMe55
GhIrKHH6qBNzJGCBD3sohi6bC/AGGeJz3onEZPyFoo/yojOnztmflxmV8fE9x27rLHSaN0koxJ5z
SKzswIURcIf3W7ppq4MRF2TIbDUznc1BPl3zO97Gh5sLPMiQ9Ib5X0QHPoc5IUP9aklCLzljjLhg
5d3KxVOcYZWrnvT9VZiCxvA++36qv0WjdOF4iKmSPiWuZe9t0di8T0zoqMPs2CpgyTBIEHQkJ4WF
7SsrSv7aK3XHu5PKGc5r69FLH/KG23QlPNXA/FyuF6KnuLLi13NSCZQuy24N5C9DnEfIg2OJN+vq
ZgEEBfBnxwrC9HVZ6gBtRrNVvpizhUbhwnvc6o4NSgjLcTf6gufTXvEQTsWPfMJOIX0PlEtZeTxn
sjhwIqNZZ9+aAO67MspO6AFSgf7UejXEFAIBMp74QJTIQQTSEGVnoLbT07fZmkqygPNNbx0NA1+T
dsZlpduQGTW0JjDvGkrblVYy3yP/AhvERvzxVGB/lKs1lYm5MmP1VGrRbCTY/TvE4PHxBiAVw1Wk
a/gjEG6rMYJpWG/H0pcW+RMJwROkdtWG+XBbgWUnV9IcS8C3wrP1xP2oRM281PHMDF2csfhEihQ9
tRi/9XgsAKHJPKl5ptyIU+w1R3OkU9H6hVvdrHeoPXwkOuOltxK0aEfljCz4Z1aR+HHYkvABqJHk
CCP/xIK3/jhhnzmGnHh3NUpxyAqnUoK6TqRAmOzJdSra3Mq45kz83bdLvbfOUbXrr8zXzxQEw5wr
r51alQ0lKjYcUyNrJJ0cdX8rRdyQfw0CBp4LGgL9cCsvAPCA8997Gy+hYAm7yKDzHuVSX+R1ehld
MvmBUWw/jRyd7yY+yfntXaSndsXjf3774MZ2FfbWHLtTu4JiK2KFzwub2l8owjvGeTfjcSFCTdju
R3MWBtYPDbIpG//UA8hKx8bVoOpW4ylV5mbI0fl16PrvDMRw8B9FXf4/gJiYq6yuunKPJc7aooPV
g97ZzoHIbIV6ZJCCnnjkhMNLZFspjZmy6V+pYK0cfxMKnxyR3Vpp9FfmhS220Ik5Yr/VtvmRF0U6
gxz3/TvS645yWBMXSG8NIMRlboDzhL3kAvCBBDpd6MqfIEiTViA39I7P8XZbpmPFhlKdSaI+xRrA
i1a8y+64UQiJPO3wOTFCXmmomQVScVe45QF9oQBHy0u6F6UqkH9uQutwj+GDoWL+zd7v2dQaoMAP
k7z+BmzVBmXafXYT+7zAA5Usymf5S4Y8VJyKkUfcjjFRCPAxRvjco/YdmLVEugmnYN3xOS1z+sdh
f54jDSx1m5fjWvIBcMvMnNXY0jFmfJ7Jqi91DBCH6IcqYz4cVTibFGiQO3EVyor1ssCBGpb8PgIx
8ctX8iSp6qdP5n0Ky1IbR/qBJewmJCgV2LNc9Q/zPBHRLR9bOr/WCgnsejDl6AO36OR4adcga0hL
8bIr4tubWUBkg/q2kg9OTR6yU31LupgI4YkZWXv6AyeLBQJ220HzM+f3ggYTcOBh9Ut4HtSG0U4z
G4M1TM2JDPKAa/hvcSTOXjW2AH0wosO6Sgt3JwZtMUOGR3y7NhnvnaTPUBjb2rtbnr15gUd12tSz
aDgPzwAN5u3OZhIKTBv1XX6AGbcSrHkpWRX6CBcBlZTzlvkWhm+NPS6lqfKzC+qC+Re+X+J/dpmk
lj8GEZNls/iVfgh9y12Z9w4DBy5m5nsgFW9dXPE9sFCpdo+YtL75j5DFmL7YSrAc9Uay/dmT1Y5M
A2YNofAVRBo2ZYv8osz/qGQhEq7bfN3UAeRXNZSw2Z+pObNY+jkwRr5/KFRChESZzjBO+FuS9Sod
+4ZXoT3mlbNSCFiMoDk/bzhQHI9gQhjYn+vO0ZW+O5YXq44tgGfeXbF72D9M5TIxYl0CiqxVncHQ
Ccwe/+KRXVbJrqxW/ki7/H5/hpADRudFEvvBOzELxnYGCOC/CttBOU4GWQeX7Aaa4LiyQEMKEm6H
AJ/mpVOU/dL4SROlY0KSVDugz3vSA1hSkOT+lppGFHycjJQFbrxlbV+zMNRvERJK6zjd2XNdrWLC
Ac4jRClUPXOowXtvuS6D4LYaYqqosOMrVfXkFSjcaYQOZ7kzFj9jdYFWE/+lpQLouOHuD10YHkZZ
K9xvxOCWvdMl/h659wDqxdXKsWB+hAeOdr3dcDaoacx7AOYGpK/IeaDipNFA95HjoLf8PZC4J3Me
P2+KJbYg4otbQ4cmJtGEL/F3f3ms5wTIsYXYOfWH4C7FkaeXlgM2qDEL2nOxuT2i2aWjYf95eHAj
j2NUWq/r0JhTP3IgpnBa7/y5sO/Trxs/5UYAzcZ9qRo0jablgVjMWT6idDCCrE2c9G6yQFocfbQ9
8o5u43ymcIr1oTpjZtduZcpdttm4DP+4aHStVTunnGXlwUQxhIwj+gduaDKegerrN9gTAh0ha2ce
E0DOfnWKmpxwLSd9m+2Uwracs7fn7dWU7NoysbsXnNNe0So3UZ3FM0eM6BjVzfo0jHA3Akrxl2YT
/VGIH7EFb1uuhtGab/703WYnQTJYt2l10yNIQtfu7aUV9vKRsAj8m7FYDrpB9uF+o8SXjamvKzEZ
VI7IbCjZnJ+nWn6feqPcPs1ywFot3tlJ3NaeebG5g1GCNAEFax0Ex9vkPD2Ra2gw1v37pA3NYJuc
Wwx7O3WC9j8BHw+grgAITt4LNOZ/h3a2wxde89S+wlm9lAgisUqr64RJf+XB56QIPETFnoKAw8jn
Q//qq/pQguP+Svsu4VPqQXmhZJRZNA5h4FEI4hQ6Ma+d/Cpbr65ZAVUhBVlcwYhB011y5Hc7Vhzk
/hoMwfXppHpLzNbCdb17q3bNnIXx8GzfyOOzY6p2n9xqQYGDnvKLsbxQPj3zSFgWOE+GcQkn0oaW
hmIQQZFQq90t+aAgHmsJITrwjGRrzuemiQN2pwOROtPMJvPWQxqXgQi7Ha6xJx+FhNgSRsmt54VP
WaGylRVyi/9BRb7PzS3jvgJwV/ZWnnwI94BTwBZrFG+LGn86m+2kdtZpyhKp+2l++3ygea4+Tf/R
Hy3bNvWPkJtjGh2u1L31S2paPBYe3l6iNFCAtdS71GDUMpIFGssGGnxRclIlt8SNnrpXXzE8nK++
+iyS5IqQ2TZYVIEVjq7UXgbrGuNJhmpY/1iwnmLX4dCNLbYqQAod5x+ZeEt2HxmKylieZfnhOUrE
Yc9lY4BzGuCeMIn88W2uh3xh54whl8/4h+k3U5wKBTVRsI6PBYT/v15xmuJTjER7564AZO7q6eA4
NhZzr+scnSIZ52oCF39jIoLl/CO5TQnnoydmLm48fAYYXIiU+lN2wau3rN648rjADI9atP3JyRxi
IMRyGwouhXrr6cGRutD+4h/+9t748cRyhbJ6UV2ZfIbH7f3pU7uYkRjwEvjHDnvwzZCRhHJ9Qrbt
BnUMNPtJFF/9wVF2MaAY7oJ8LG9h6orqJayW5WODPLw35qXAHVBiBy+rk0BurjM/43vc871+HPsO
KJaGk5mJwxjhTEX0m50NRovhNvmQ5H+JDWTKGm/1paJ6NYD81u1GpdZ/VtpVByByETZY5U4x3lMO
ZVOVTW0OCOU22pRvkJrnY0BhIvVld+p0BUn3K+UEqtU4iV6gWtgqGBeEBdBlcLuyuHBBsk/pb2Pq
4YUa6ZCyBBo6/wuCPdKWoZyf7+ljLPnphciZJdBMbUrwygxACDMyc9E9gpqf+4rgpKCyhPqn0PCi
/HUHQNOMSYV4tDHW+FHBlW9P+OZtHjYoTWela7/0iPVSI2YvqAoc0FQADZ4xZ73wrXKcup4d3YhB
WbklegxnOXY+BPafTvSU1HCogAeQcN8Y0DNahfYTJkQOW8Ca9yV2DDDVZCO2AieILdRhyBQrgt51
9T962Ks61r6g8P2o+5Mk/Xe+S0d0YpslxlUJJYSVuasT8oQQ96nzk6lpzLRDknZ2zPVhGyx69Eax
WIZ50c3uiJf+yoUfL7gmHz61uK56t5hWgmwM0orgkBxyXMwTaKIh3j5VbSBySTFDK7MSnv6j+Q9C
8lc3JJumi+WU9IPWLcsWo3xdK1uiL6GTuW9KJBSB2ibHDK08eyHYg8UPRsXRGlETflJyLbp/vBjh
uKdxaSszkCzFhhRufY9XuSYdfyhG5pqxT4pAfzBRMZU9nt6nfa5CTUtUM0uf93Pz1LKXodzaibsp
6lt8Jbgds/lVoJc2b7WddD0G1eIZ1qMFyqll2ARjN6tT2Jz999v12OqbQVwd1qgZeFRz1MB5P7N/
vn99apapOT0QvBXQKI7z58AscdCOx9arF9PR+6HS0441gNFwGjjBpVpjrsUTzZltbMVDGw7qAuP6
zuLvi+VH9hDVa6Soqtqu8HjbFanrX/M2xNXize7Tw9XLASSLB3MoAZPUrHn/BqHWiNyt2s9tAfha
YdaWizGYzYSF2ZF5q0ErcDKBmctFnT3lUWYxupyyu+M9waX9DVVTMOBb+p7R5wQgDOrtmczTyrJZ
puqei/MMhZRyQdynSD2XKgZIRi+wll+LqI5gl48bzQC1GIi2UwchN3SpoLAqwY2QX2TVAKT096tu
A3gbN0n++wZlFNWtTFqVknEsKNn/AWvOpJJQoKOulP7VvtFMpDz3kTo5LijgY5SvK/MVhtmm+NyC
tnZsf9dxYr4w77+F7Z0s054d/80/9PEM3JNz9fJeq3hnzlrmai7h4RyWpo6QPeAHu4EhejOKwLaK
lCh5j6sgkIaFs271N1zF82h/QkZzB8M4S03C5FzniHhSwHwO79ExQOKIfUqBK1c1/eTxz5/TUjRA
/zr76X6AOjeVnxVoa2eWMAe0U0o1O9ie4XgWdQVtbPMuP4HN6Y6EEH24sUnTKoMocaTyXrPY+lA9
aefJBCbqfwnRxzk9iqQHXGVbC9uDyr294i1M2077Qkq+ltupwD0FwY1MeTKERI1WWMAt4AdJwjj2
re/iEWgkgBIRBS4x8XwpcTYzanyTU1GFUTDLDapVZ0rrDr7EuqeuYMINjopbOHQ0k+0YALfk3I9V
S6cfond3rexxjkl4xBMfmA81TXYRIXPVrYaHEss+HW+rX/v7B6O/SvDS+2FTZ3Z/QvZLPT//4lKD
Mdrgx70V6knYNOSiJjbie7KpwYN0Po3I3+SAIx0VaUQRJFymP0z61Ls/Q0PHpvubpl28A4t+gX7U
+BJrPa9MAbtIUMdFzhEuo0D0Xj7SXQE952bvN6y85n0ISBect3rX55Nt0J38TwDpNM17ZLhQPlt9
KTJfD1sIWci1GMUTTqC2FzJumpW+sNj/SkVGdvCr8weTXTqE+Df5GfQ1MmcB8BXVWU2gckBJYdoB
TbzH3S0k+MIcwKouGdEZQja30IlCUySvJo0GADaC9cXIXbx5k+Um/J6Yh/dvRzxb089XyfWcMJ9G
rLHFlisVWNaqeyQjVnTqf+Jls4gf0u9hOYf9bIDsRW/fNiShtIDsU06Nf9hPrUG+tYrW8g0ColIx
XNI7cnNCwc/2LXGNmTuQCrWMCMEhFS34ACdsa+lt6vBH6noDiBN3/J7K0GcY0Aku4QAou4bm9lOL
lfkhJO1b+PKT548hppJNGg6llRX8UCD+PayzkcyO1rRs62q4H7yMkEI9H/48/wNbbYfDmsj5fEn1
/UG0mEoJadmzOJ/2DVQ84eRsZMIak6/Q1I4XWMgNlqiH4wVzUbsZJC3foZ1rsriBtfYZlbGszyIg
+elKK9nND89v3TdWk2tEj24SIdgM2Z2BIxTzg0/B8GXxxToPhAAiSLy7YEi7MBjkEWvLmuFjmEOw
beJHJcv8dgLBQZ+s0cgZBi0xchVmEtohUJ8/WX60ZT+m2R2oquiMY1WmSuR0lnW5bAPa12hbO6GR
3h0k1DwHwGX/p1koEHYDNIZKigspT3a70MMC2GJcT7BKuDv3CcwWEq3bAFOCT5mGWkolTJkx6Api
5wt7UeJrIC3E+vVYvRc1zuo1fErbs4ZGC9NxdJLcmdMp+ZZgYcomQ5WTIhKWuzMosuc/j4HEad6t
oB/WIfxaqQbHKqIsPJMZovmGFmIICLAXH6QK+wDN+qQTeh5ohZoTnpmnvYDE3xaNxYe3zbxMXTQG
tc85PsjZtGv+dlDXdT5EFa7oPTI+LP1YVpvFntPFM0lDEMj18hxPCA1wjGqpJ7kJSfhyTy1gZfN7
g4HPduedS97AzYj4ofjjlmmTpzUxn/0ojCwEj2S4R+K/n5m0ZZx38c/4aVKhS+sqip3n81nEgrLM
1Hmvi/CeVycHbdBJ/BrL1wgKjtqy+4/BU37DiC6Pi+CyU2OBqp38JXITfUvrWbvJYsRckwNfTIhJ
OmicqAAQP5qYwKL+d8W9zw++4nu73TzMZ28j4wtEPxnAvSf24nxI5hE8u/89zADnh/aZuzv3wWyl
EKSXGrQ70mMIAVKeEj+ehYW1o4DJlnRxf5A94M/RM1/zNBZge6uwew2h863UxVmAQgLHxZt9Rhzy
znAOD7izZaX8P8qjOV7nnnWHSUGxnzpDr5156t8/+XxNkAAsHVccWKyxLSJv4ysfqcopk5+Wp3aP
Mp1rcMBhO42sXZQB8MwCruEpteW13dk49tb9ij40jiK8LPNUkoTSVnG6YUOz8i548UxRDb0frr9w
S6+pDshqHu++JWtnRa3OWZBm2z0RM16Bap/gsRAyq9m+Ow0sL+SyKgSGbgucRVK5izRIkIeczq85
QeDD6Ef45W0/elFsFK48ZnyU1e8cXtKTymVRLyFPWIC0VOofc1kLkwiYypt/HWGas26aTxK3+NtV
0S9GBRS8VN+Qy3iHqiZQIGuphL9GBVhx379kb8yBLqKCQBYawjNDjF1nUIaL5n6XXxB7ZBzn4Wte
GMV7sOBz1qJHeuJLFC6ecbWBLuSdU21Rz7BDuPY8FDRjQArfiliox2K1gxEiqvaTVdm03syl/9Av
JG1MMp84DGzPIbG9KucjaG4ri5Lbn+qXFwnm6miFZ+ebOaPrPf1dU77iQz8aJncZ8RDENQKdKC89
cCCkl5l0jrsp5njoXl9fN08iuTrZfZdDfK2JD2tCS57HJKjaziLx+c4s5xbXMI3Dh9Q+zxeK9Fs9
rG55f5OtZx/qcndO+wLp0ewXu3LVaTDnyBYbD/UJov4MWD8W7nstjkDslqQ4S4JJuX3eDy1S2OdP
46DGfgc8s/LAfZa+eHF1Z4AgnUL4xQ6Y8q95rDxf4hHWdLX07Vx9xJ600yfdKd5qgIBpIrmaW1dK
LB4FbpnPqvrbjofcTPrCLrOZ7lLxlxUaA3YgDBDyuz+qLa+5BnQ0FzFxebyiwIPfpgjzozQkjkwB
kMo0r0lZ53VNSnTiaNOAHf7k+OJ0dxfOX2HgII8F/71gpOryf0T+FjQtJyESc8lEbUWN1QyL9znb
HPpu/tPBqZjPs3tDxGRDp+4sLmG1UmefZM+69O5votYp4CjVEtw60b+BjmiI577moBZVQ7y1/8Pv
fF1wF1CvgImu52tDd/io7OSg+0xOjPIGmhuYHXziURAKMoAHGRxrSodGdOoZjMgJ6vvOiKIWOhMt
HzCBO9IqRe4oZDZMFRk52eEcOi3RTBarlDthBzJr4MagrrwcX1ZRWkkTMmyleizPscNynByqmqQO
mNmnMz0gumu3FAXg78gyKC0Ng5fplXGM3QBo5cwk8hQLU/bv3uFnozOA+/gQ3DksrHdQ1NcHGWO9
8mAN91zWk/7P7v5e+OOJkgYC0gLCLp5YRs++ZsHUtLhbxqYh6JQOEg1tWmGjmiXkv6Ja2KaSg0bu
WtlvC1qbiR/cPXc00aWF08OrKJvc/am7RmQapnv89dL93QN13qPqvJjlpZdnkWWZhq2O5bL/h8eC
CWcKP9BTuOv/6ftl2F/sKNckoiD2xbl7dAYUJ+yX/OV0ZsdVUkst7bvEIXHIMyFMVKFAkk75GeFT
ST+JpGCYNk9kHflbXH3lRMv+3WzgBRnoF2nh9Oep0IkMKyztOaeHwotviD494eQMLqgXylxZvlWv
SzVX0/3SaPtCWAvY22WFQS0OScsXND9TYTxr4fhY9T6UcBs+e+heuUYPeCw6h3SA+/81/kEwcdVk
yHMT9sKo5vfATKD8emt3AKOaGyiwyG1lHgyq9cHhVirkPm3sjjSAHB7MpF+G8aPSwtOaL2J222Z5
ZiN5HP/dEKmeUWJXHKtj9mUb0jnm1cCI0iFby6jvU9gZ3N/6c3TICcN4Jm5qrWimTTkX//duzuJi
JYnUKbWEADINF6QF+r8Q8L1fYVzVbNzc8HBVoAsQiUFSO+21waCPq8OghNkNPSvMr1c4NkI4Bz9l
nbnOAwRR7mKMfni1AafN136V1Q5w6/iCqXNITDJelnf/IqwFNbnm5ZMhMqqFmfa79nl7WNJLuGNl
UJjpnBdm1O8x6gnnhsrt1DIVE3QQyTdTZfVfKg/QnEf8WKFnjLnYy9p4JJB1Y87VDZVPFXtEPaZr
204K9D90Sbn47pq2gAkGABOAEgnHp67FQ5FrrZ7t4+wfw/jlgJvIVQtS25YDUTkKsFMDGtuRJs89
xq9168QBgyZbymtff+5AbgpwmeXZ4Bp3Be27SduZ044r3cHQYme5evOWyfHq4QzUztYryHOhtU2Z
LI7EH6StfKsjfFXbY+IEKEjI17hytGsws5CuG7pMNL4dasApZRqNERHUycpucgJZQR1xBdcypbeR
UVLZD+9gL4R/GZE+SBNdN/vx6VlECIyeA3xsu+er+zztpkB3+ffUi7nwKROiiqOZIaUzJtbixU4r
eBIMe9kgAX8sIqBJSYDUN/ydi9sWBffiopMZYxEpyWtHpKFFFqkMGNWdm19MR9xPBSv/HR4ftXIq
p0mRX77B83LUDDCZrdKYTTG401AhIzO+kczBnKx59GId4Rxh4QgKXtsVhCqMLpKfzEQf60HH9fs3
BWbmlB9SNXNMfj5dbLwci8hGJTuE4MGgQdmsGofGWQ7MwAdS9q9BG02LxeTs5eDnAzzznggTLdNF
cCAMTI/G8Ku6kZXaJmvdju7XyfqRaAYPNGsu9Iln6WAKO4PPCzD1k+B0ozw882P2yBBuoDUTTWtb
i18SuvVkJ9cK/bpUTy10Lr1m+N1YOgdewwoMDDVpEtSn9XDW78BGIgTWC54c1AYTRm5tbcVmDzv1
sGJ34nCgF9LU6cJogUJEZIJ8Sq7dttiuGFZvYYQA4jY/5RrCsoxqco0k7mMGDKTwIzdH5gQUIU61
5bR/K8Wpqc8JNgmwLxVc5N0Gwfj5mPIZcDCPjcuUQI1BuZXfwcBvmqbtYGIoG9DOFO/H8J/aVwGX
FG1LDiwA6thVlEfc/fnWP2qi1KS9e1Y02jytFHndBDfnMNLpmsd6GlDe53LrZdRaK6In8fjZMJI0
THFwvYJNxsdiaABr5R9y4lW83ioIYeIsYcVZkRLtq8G6b/M+OB2Gg/P98x1iPNEU1qMWkNADwXOH
q9m778TPU2DsYMmOc0kNxOMd5AgpXRafDPbgKuBprXiq6DphaqPfqC1LoNGfwQVRNqSBgBuv7XXg
2HvMVDg4vFZpNCa6G7NNqnHJY0D3qP9knCERBB2JurIU/eSYo3LDg8ZZY2bjmbxS2CvhdZI22HIU
nj/aOTDPCLFZyhm8XGtOglIfRwfuTAYxVIKWgWG+FgUIGo5zHCr6BKqdL/KZTXDl+RWp5hSvNVrP
x3vjagiN93A/EAmE1o4SkHAJneRQooBxmyCNuq82nFb2+DoU7rtp6pg2bf8nW+SPShNUirros1c1
VQAss88ST++PwIOYrvZMzaA58aJWNg/ZG8VoDmgEx3Xey2bQMQRWUJgUs6BBzi0sFIG4YDY7uWZR
5a3swF5NYJINJIyOSsoQRKrMRriP67HnN4GFKKafXuIZkWofLj0OYJ52lRI/GEaCWViwGOiQkAj0
xaKphXHMhyjfrsooVBc0E+f/XeEjX+u36Ffmt1wepNCNBWhWiKPJS6cKJoWtt/lRwZsZza5oRZzb
t+5oV8SWWixR+xgJJ0FrqUE6e6pNIOaCVrCiDDwFwsTtVsreNpIYxnqMRM6LpCCe9KJ1zLMXszs6
cKyvcGtq5f1lRoL+GfkmCJ02iCP+F7wCa0WNJpKvQ9tjjDGOVWKur4PVeybWQbSzChxFUKhLxv0F
RwXtIMrO6r+0wdlqbFss6r6zmfyU7JJWOD9VLY2pIzB76eWfRpvcNPW+tmC2nUYfXR94K2cnQ/1T
kaVRD0vAz61N+yKvAHKhhReQ+KjMF+rDyGymqm1VpxBP6oHMPKoAuRaVu/Er/OgMqGGb5Gw0lG65
QIrN578QzpDN1hod3OMcPGVkUCSsWdd29T2LsHemXSuwlBPPHvEjh/g2W5Ebi2wfc4JXBiMbmKBA
KioQt2SflIURPSUj1p8K6nW5SqYWf08DJcKnStiWtySTjPexugG43RbOcutFtu77OG3JxB3NZG25
Jno9Ij+RjswVWaaBBKnmZY62bVAsvIyWkzYD6VErcJcaW4KNRQyLVdsubxR+W0oSlzn13PcPY+Xg
taOkthzyX2kZk+56OtHUEKGLTo+cQscmxUauMFWvADOPbARWEgUg3oS/RHEqHq1gxpOMooJrkZh6
T93INEoPjyNPz6Ocqs+kviwB8enzEJ36m78FYCuYMthluO7x84+hbbJxYOZrqRMmaqLrqA8p7g30
o78FyfHKJTUH+LxcZWJLy0oj5/7BW5irOdzvaBlP/5FTKMqUmhTa4V4MhmnqFKXkdTDQrXGFsU8k
pIJacOCkeZKLTany4wLVW5JZG5lQdzmkeLKPPqJy9dkUggLMqvngFLAe5uX57HL+URWAkCiA22t9
34Sh7AuBbTD2KYuTflMHjRLm1v/hqSv6Bk1vI/1kuZLyRDwYBKQtwLpKskJYaGDdy17s5CogL6Bl
YwyFzHooPlmNJBvS9500IDlwbHqg0v8IuU7iMgNJc1XqE1LeeaHGyBJtxQ7ZuqtzGPkGdjxV5CJM
9vGebq7kpYUBMZgqbglXpsSWvohjCJpcNUZL4S6zes6LPc82WrorXNQQA3e/+qyJ2MHU+ZvUmXxa
XvkMe7ETpJTtPQhoFrZ/Gx0RQXrJMF0qi+vyD7Exa5WUPFac6kecsl5dHFySaP3PxHIarENlXsH+
noePPHobzPLVlXGd+0wng0LmU0rHLQ7TYeMogAlzO84Q/mbcPNC3h/ceDDGioG1RMun/Q948NJbK
QBbOGSZ1SFzvu1KLlKC15sqpu+QyjjPxCq46zsOvktt4wGCmHIoASO3S3szl5WelfwL4B3A7nn+l
10GyDXGUNRPqgeyUTUB1XrKL9uGO5M3dE4JXGd7+hC3jt+GP9FjWruNjwpakt57BFXtDaO0JHXT0
4BU15E/T/mORYaL14rYF/9yKXHQ3ERkoNWsxy04oaAPXdsCTUOMiB4OGDWaQKsQEq6JGpD+W9LEn
5apNECHehsRAXJ7KlmdUxhuIgshloTHbUope9pSOiJJT9oJgHptlKXfPSxzQw7mcnk0gOnngl+uZ
ycGEEGSfRwSdPai3VWHeaIEF/lPC16x7F65MInDCN8YdSMlEVLWKh28tMjlJtWyETVPmz0OpjfO0
OMxhPn3/qvXEc71AKTndR04+idqY9E0gtHNi2fOGG4JkrMpiDJBoogbq08aHCa7bhV9no7b9IK8W
9W8U0lvB7U4zy4UYB5/RKl0g++2iUrh/vUejI102AbEs1nPU+/hNAtNSMIdq4lEnccD1tgmT1Hpm
hojrAkx0iFYDma2GHpXv339j8xJ48NfwCDKh1K7c0kFQZVpX2CE5+Hu46wVaksIvHyjBPjVSxpLa
g0luVvbCKpcPp2vVXDRXUG+rFOFoMhktGKJGR0T+ZafDCtcY5H/p+hzwixzEfvX80mL8HnRrMA3q
1iW7B/s+XDF5qxMD0HT243HbGqytUpFl+ZPdySzPjqCcrwPhJf6+ZQ2ESwT8z14gwKxrGAwtMy3N
fw5EQU9F3hfBcFaxJ5/gzjePetOinqwt8Uv1fVWY4J/xgwwtdTAoT2fXfFPX/C/sE/4byFZL3JBN
VIWJUbAhFZ1vuZSGJLI9SVz0WFN0ADDEJi6X0pXt7RkiLhO8aMT6SajqWC8frFRedfVTP0QN7nQC
4PI/HQmoff4JEE+AIOEsEaEp6kZv8rEkCLMgqZ9dg9p29oVM8s+kCkawpJZZ1KLrgi3oHTe7Bex2
3s4BrFaYwPG49rqME/wE2JBtRUAilOFtut1V04uaRJ4lsSb1A7ptm+RsqEV+SYiqNY3gTjf6pLFx
gDxuWqYSG0wg7D9q332p+OjNq8Q5DAQtqdlv01W9iJI3ucUtoCSodwKoB6U1WNkk+EJilmoir7Xj
+DxnSusGGMNQjyIYhvKBLDgLPhZw8GpSkPPgRXXcxt5u719j0qPbANa6CT8zmGhsFYuaToMWdw3i
kmIeaZ9gA7ZczmQih3ZjAheLohCoeBdqVmWI/PajnfUiINV0YqfRVhHoEr/cHxg66/McR4GryXcx
2mRgCltsq39nwPoblHJqXfXZAYF7gz4Qr1iTlkYTrVBrp+akeAfNAJdHLcBxUxS6baxRRkt7ktK8
77pkOu3EWLNgViJxe/DzN8Np2rGOaedaHVYnBQxDYM4PdBjvLEzqWtfr5LSOZnkNzQiU4tm2U+48
ENzLqdnjHwZpEWoOSrfT4qSsubYwUlJMvr+NKy6xhWqTYrviqCzuxr6JaxWcECNRFzHoOkNNDVdI
xDrClhWfqUYEh/MxWeQGwzsAZKI5lqTy4lALjztkNunFJya/VZjaLot1RnHYeTD2cYVsXbtwOOAm
9omVXThdL58jIyFJA1cRdMxqVL3cxaGccUqcwDp10OL53NKjkoCngrMIYr0s35jis5XXKmV0IauO
k/3KEqff1oLHgKS/S01s+bBo3DsECwC682WSfMKOMLTKS6rUNiaGxHnfFgUaRklM+EShnXvpLkM9
lEvVLJ1TF6rVxdG5KzV76uSaBhrLFmxyxmGXHcr/XGcAgHlm7qg65hdqU2WtkgWC8n+M8y0DFOSG
3GsUbYckqQHp7ygMNVf+8QXGCQuuXkBS3SP+qI2Pm6z5csIg/QYrziMqgt9Fquk6w+fVnhNnhGss
MBgJEazWn5oij4+C2D8+VZ6klwtAY4DZuJxvEb/o9l+DhF2MVz2y85/IbZZOJIhU1PsIsbLUjleT
Tb0zRKq2yoZ/Gb85/5ThPFGZtjx2OB8wPWcKnzGSJsTCRtluQd2wZIXf37onaWfkyV6czvq8twqp
yrym4P255doPo2vuK4umVvNzjWLKm+S4nkRPh1nDyaSkJCmXRDtuwblADA4XkPBvn7zEFgOavXkL
nafpSQ9dX/2ixghMCCLs+9WdshaHAYLLvJV6A755UUJtnP/AnWLYu493qL54YA0pqLPSeSOv+aeX
ZdGcxLexbSwN9BSO8kveWCx3wi0oCT5c/5ZMxYrClGxy3J0hTOShgHAHtBj6oCgE24ClFfsLEjrz
2S25hTfXGZ909Ist8w/DqeQpqEIKo5zmnJYue/ZAbm9ngJLiYfRf7cAFbcmkvKrxeMIfdI5diiWD
LRiSynKr8V2QhRbGhbROj9OWNPwucJFKE6qwIy6db++Wvf+ktTfINXFxkD3cv0XHMWsiM0ecGUJR
9nt/cu/1fcOymYaYAauwFP9oppNvm353vFJoWzMfq4gJ1CLRNWRdlO3OqNu1zYe5nY3ancC+iLY5
eGywb1ZjXO9FuBpl8Dbpkp05ul3GaBiS9+2kHnl9z8rwWMvTyT30wUYTpe5WSA0eK7u3InBw0MUo
XxOVX2SH1WZ+zWUA1LCW0cI/yYT8vAbLNnz+y9Y4ytKzyPFo1lNz7wgIgSQQv5yNxzQYyhE5macD
G8vI4ZeIQLoue0D0ms9ypsWal017vqSQX/rCKaqkBdCnttJhPK4RmDpQjoGqFe6a7mGqdEg/D0tW
SBjczJOC+1yM8VVeSaVlQAWdDKTLVg8wYw0480h2xONjCuqmphBtFdvXhYwIUFwPkd9dH5b9VITz
sK0UJuYzDU8H9eOZvtuoENrz58nsYsDBxvg+4S58kvVrasdJozUJHob9hbqqG4txKipZoHuCGqkr
ZdOxpYOPm1Uo35vrX0196NzQVFjtfVoraFwYrMnp29LLhFCGTS3rbA51SjL1pjmcoZs4p7EQn5LB
5B4DGa6nOQeOJYkhlajEWEiNZqN+YOYKMmalSyNGbhKiNg8sZXlEjaJBZx9bpYLUX3NcesBV5xOd
ljvwGrXjFqAS+GBDxVQD6odCn+0ywhoM8SeAyUJSra5uVu78N1nTLu3QZ5hIic8N+MfdMHg8jzsV
VO5RihK6ekFnHliCHhvRo7Q4kH4+JIxm7S3Iy92tNxtu+wmGqP5CovZEWSrY2PExlIOBYZkAcoUd
bam8azkzWUxL8TEdXQgFZN1D8YdKszQ9GYbtfIoEGcZeGd1xGH5bIULKWO5RFXEjwFEESAkG0qfC
FesljNArat50u/fytoiIYvYmntNLvy6lF6LNnGfHbSZaoPKN2ZMbai2Wn3O5m6oSeWq0FEoc3y4j
0ZzH0qDq3yHZQ5h870APrd/KfLeiNB3j8xCREcTloO/rtSCkYh0iHoUEg7py7Y5+uHdEMJo1XGpF
hv8C5AMdoFzkFE+MBpAcdKuPtLswoR4l3HOft2Y5YuvxysB5GBryyiD6EQprnGL93COKT26kQFEt
9/tQJBh9pKMRD3hs+MKA8k9P37auwtajZ0MNLIXaoWC2ZiIlrzuqyED+Z9RC9glrN9oCoDaDAUqx
5RR3ur2th1aOV93/JRYSPy4qR5h+Sn1l6qeTrpQPFk8M1CJvoTTquNm/0LeRQ2AxABQ1fqoAJ919
Nr2EwJNejuNLBbYA1saT/3koO3BD3WDXvvvn611NSnjXeAFNiR6yz4fYiToVtoEf+9XKAo0CHru1
WSSVD13IChcV5bscvGFIU3zNdtIJPY7tJdvyxQX2KFE7BmtB03CnJv8WdY+DEyrXnkArETxp46Z5
FXPMA9bG/o2ICoi8iNKhQ0zLXawYIWrZnAD3Oc8Wms1JS81PAkrMt2Ltrs+Hg/P6Nj22rvM2PPaw
Gd9NVkiBSxVwHj8JUwGEj5ULH9ZM1itPAKPiBPQ9Q2s2N08C27TDpFd8JksvYQ7svwEJgWPKzSkt
NOOq70ql3YGQ58oXu48lbXsDCibCLSqp2SYAPR/9mv8UCgfX+f66x12YqggNv49p2vw5VmymS6Ez
vl06B+TqKrmpDv4Lgd/ectpLq0/0gdiaPOTZSM31WJjgTEiqXz9etwQRJMMSzdc3YITa7XQpVdmB
gaeDzwwT6QOYaNBwGQjyQ+wEdFdt+odoYUkIenLUfCDtnJ4kPEqu+Zm6ejAcOS4iActOyl31KHXJ
ZwSg2KTb5Vje0ZVG8eyV3i55EDZ2UOotpTimWna3thEel/sBURolshvGPvrx/N67Dltcn63ahDKm
vxPxjRlK14K4l5oN2wManuUozYsAodFj+qRjU0Q+E+ZClPmEYXl3LxV01je775C2Op8XUE3xem4J
Uf3g+j1Ot0Rm0WsnJ2Zl21Ayv6cnYB8FFz1BrS1UNV8I9jepRef1U/bgqb0Q9j6Q4pHd5MuvbZRm
DcCkemzN1A7vbL5+RDsweb0sk6iKrW2up5e9IAaUtcBeH9UOKVJ5ZkRmYegvZ5vMyvVS3+iph8KC
VFou8hROXNkj1UfxmT3DpRHJ6wouAQ4Zad/+ucnLbnisKQaFFMG9yk3YafbuT2oJpRlPBXmzpwQa
HBLtrJDmqipWEeW2thGMmY5ZBzQpI91vb/JfDMRykntc+OYbzqZNWOTnBd8Gq6RU2ihGhJOG5UaI
Qqt/Sj5NwplGmhoLPrfAKHvJCa/MhfGdHqW4oVWnaC24xIMlABaDNpWKCX52XWEpK+AZg/Pw0XMP
QVHVGIXymnDrhru0v5gy4y/2/771yq9tWEqv5ivw3TxRARIoKUyp/eT7Njf+YssXpQwd0TWUJsPQ
6B/IU25Ebm54xhBOwEaiPSZcOqXhZ/tbcB86LhafiZi0cuU5zNRbX5VyFKG81SQPIFFASKocLuzS
Nl3dfBMj1kcNC8kEtO3DHgp6NsDhRkKaO07x3evU7gAB0o2uA3uwmF+A/bpSq2D0bErCVaxggQ3w
Hgo5sgLzokN6dhfb3HYRPxRZOXbyLUmKAL4KUZuWd+CAjXp7q44nQnfXHuv8VKCfS7ZPp7WPzeV3
X1ooeXEr2glAyy+ps84jdb3PyxlYqkR9zrFbUoowzuZVdnXvNX5lJAaSdvUB4H1ar96d/wbZ5Ltj
MYV0JlyzIV0aSuHG0zkG07u0vE2QH/PDYvi8NIE36MNOLszWLsgyO7wJHuVf3wRXPZ9bhLfC+I44
T+SISD4kX5ZSlVc006TtDkRd/8ZGjZ/ILB1AkPG3EpzQiwRZrC2Hh7UrQIpKTiz3t8fb3NX9tY01
ec7OqV2rTeKD/4scAIaBWTZr9M/B+s61LSJIDhoRjvEXZhbocYwHF8UxsKACMLvuBc46d/+H1db5
RD4iZZjH/1uNNO/pIY0DfkQZLZg9x97tOrnpr+ra/Y3c6TeZqBLu8rIO9Occ0Gh5ibYQSrCu0e1s
sOlEKVInSL6I5qLNbNwnPldtv2ueee3JwDi+Gz0yAflS7VJZvUBF0IUqHPD6kim6+RPUdrSmBnCV
f0FIJbtkemSnZoSe8/bvkGQhdRoa9Alex1oTM22GvQ5aPtcz1xVE3JFnI7bTcXTGNDoz8JCGcWVH
VJkdhCisq7EL8HjYYV/Yl6BQZ1ow5e+sHiit8EtKIHDdQNW8TEYZ3r6FHr1VHwXM/S4HOvgM3RA+
1AHD7bj2JMdWPh5qtM5nfDEFvPLXjlI1HgP2FaKDSA6zyt48+J9RSY/qSJjX9d8bhQ0K4Jt8nf4w
xDRY+reP+CUNlVgvIhyBYGhdAXYPlt+BfBDnQAuu0yuLLRXnBcvPiCh/Vv6zn4vGAvkTEV+vasVo
Sde2hRggQN7NBs4RZG3rMun3DZ7WgZjWFUtapDDWx4LJJSmkuEF7MSy6gtJcjQdgkkzR059cx+vD
WUGqpkbgnUHbpPejEHGbODLNewEIsUEHLffWpG09qRWt9lSeIEebKjYI4AUdiZo/G45uhQfJs5up
AqagWelQrdFRNghWwxJaqsUjBUbtx/18hyvn1n+2m/h3YTjr/gY+SsJFCBVnL7M4qlOgz10Y5o/5
n8D16ShaAnuiHodqgQXEcX0ux2zZEXwvwo3IILPtbw6yPFAzgNNkzmzQupqPGZmjcM3nDQ7ImB7c
kgiSiLM0LCJKiX2Fd8W3FjB5jnlLm/K1xhRXsvHY5CHc8gTs9NqKKXvXhV0DdH+YTdR0Wy2CTG2x
xaNS9R+ESk0y2U990V8u4V/8CdP7nXDWZMhIsp7vkMNr67sD5mlduShzJcm3PiLUj0FHLKu7ni4C
Lq4KS5bAxo/pAvV6Hm7ctwbb25C86NdsvHrXrTnTuwdIEwz5Ta/bYS5FwltEP5i9RvVBIXkaeLPQ
cuDnKYAwgD52ienBMUvwS8zU1norxK5R8DcHDEzXs2PayoKlxCY5gnxGYaEmi+7hPgcjd8h6g2qU
srKwW2YjkoK0NACoewIW6E68Vh+VSY3SXoaB074kUc/MTcTlbMkpgW7lqxSCZjhYobQ6d3TRNcfi
vF0upUVoXBp+HT5gIDiirJeSvQB+3MsLQGd+yABj/oMtWcsAkbbPH0ep/Ap6Zj0EtwBMfn4jewBe
ov76Euxqb1UoXKbq/fcb8k2GYSfytESAA6Fa7hfgR/fT1T+tFjNLk2IWwQIK9+XcE7WQATyxD2zB
pXgrfDMxZTEoP1qD97paW4hWG5GJTNFVXxWMF5oq6uNC80J/Oc7uYBeetKIXF/0ENsDPh9Fh0Gek
0HONYcJUDdI8jfYFiECMS79lO876X++0OKhuhzVh3hpCEty43ss67Pbg+nhognb3YjS/GWcs9by3
EneFj4/HIRNwsU+rFmLfEYeiRzZhY7fug6hryJDrvtjS6vv3TWwKXCIdvYXN+VS3mtC/lUugsoo+
n2AKopujE649IFIIUPfuYhnti4adoVjPaxXY1gJ1bMa0Ku7pKA9s0HmiM5oXltnrp4CNh/dNyO6t
jwkGYyYlZ1DI0k0ZO81s/ee9cbYclFj/AGHEb4BBYKAN+FR87tzJ54gyDlozc/EUbcUJYTTPIkBd
6bszHCf22TujF9K8IkP9JvOed5bcQBA/tHMxZTlBMP7YshCtdB92bBjTRk1vMbKOqnkhP29/WqV5
J0lpmyzBdSB1+byrgO30Z08gCmRB8YX7ZfGS1ZT8WXByF3u+pfHrIqfsnpJbI0FayeL1eXSBOlfh
+YDIAa6mDDkTQWYjd+Ok881Wf+p8xTSC+o3z8mZUGPZxgS1R2pvBzFi8piI9MXmk6hpQvwO3YZq7
Ve+VVYMcu+lZQuYezwi8WmPUj5E81m0IK2kiX25PniPphdklo9ZTWU442dh+zblSYmt4EeyPP9e8
uxbfQXiBaUQBjq3c4BSeTBGQtSLPpuV8poVZ6cmW+RSZPdUXh2f3favULxV60OP0P6n7XW0RsW9t
T8VSC0D8HWB0hKaubz6ZULYWLbsQd8KXPXOgvoyR2hNRpOsHPeuYo823IvBaHrjWvAR7wFCLauR5
179AiVnjfyE/HcDnSR+N/JGyMDQ0xw4lDMeo5QoBRtUQLoYHIiq6gzY1RUo83ECCo7orRpgPIeS8
f531aA9Ksxd92fMxd+4Gb1MyEXzO+LMJHtdid036jFU4C161a4zKeKXX54b86iTpGJWKZNf0pstS
LsJ3byqmTFKRIegcYupLlo0drvTJRfafu3US1nM+r1hihwE1SggAlzJs3bgXdAaqZ6I0Itb4COLk
JRcvcTrGrJV5XD9TFeoTv/DVWTujqu1daZNyTcbVQ6huhaj3hrwgBs+xT+pF28yqzwsuwZGDfooW
bMf+eUTGxh+Ony7zsAos9Hey9qMqzh8DU77+khlJF/c8guRb9Gc1SDKnOoBf0N1wA+Ezr6mDaYfs
zp5pdBfnuRIMMy7FxMdggBPxTlBr6hqw0RU7hzalTJ4Efy7HGTRhPDu4t65NpgNZtuCtQ37eOblh
gsw42F1uO54rwuAgHKvfO/qgd0PyYjvK/iVxK5VsG1mb7cwmRA/hT81FPdOoOcIXMY1GLkztMPVF
/giy/mdd6P8XcK8opa/A8C3EgMHc70YJbA5PsSyjeX9Ov5XrK6Ouub1wRLzjv4uqW0VcEL+NSHX9
8yK2LU7R31Ej3Y+bSbURLgyhK0sXAZexcBW4pFmfesFvq4b1Hg2bupMS2cyFyHesmZ4p/90yS9rj
gMRPOsRraclR/noe8DTK98OFRt3LCx5Xt57LcuGBesTWFt24Ml8plFYgXaNx8dGlAfmAPdpDrpaZ
VCzji5FMEp2zQ3yD0FK6+hpYknJOMAaZ3iHYhZW6qyDcJzuJ2k5Jq3ijmj4+/bC21Lyf3S4J0DQ2
prWsc8VW7u2Y58jDb+terUh0JYGJ8Am6A8EbptJzvBXxmGxH+8uNTv6k88akFe3e46gR7Qk8qY7A
iOVcwGo4Gq7Ri2USgy0NcS2te9iInlBgAx61AVSelgHVgftbQS0NIewSZLX3BCt53CDQ9ydGNVt0
hcJtiQPPdNGbZ//Go1iELnw2XIhaZv9MQxtzjHe0qyvbvweAaj4ZmbkUBx7vPHzEoDNGVZYwM77f
w87MShX18aknVfNXClCH79RnlOu7rQ2TX/cAq3qH6jl1UD/ya26T8AVQSYjOuTxxZBR9blfS/Bnt
fTpUzuH/ty0Z6pe5Z9Gq/yIC5wkyLOLTeF8uttJQY5t+iTJIs/3tf6qKxEqtQ/A34pAkmbmne1aD
0J9DRLL+aFLcHuPUqzkK22VX0ahHWDpBCcnyptGy0F6bmYVnq/bus605xwv8p0vdl5X6SkRVZQyy
ryocqURkOu2XC6w9GLfSWlm7jGZhLBYTKujLbMzQjz+Z50mVHFXDjzZjKXYA3yJshYZ0Wx+A+CSl
453gOaVtNzLBJwJw+3R2U+EVrUDO/fiiQKyEgGrrHQn2EqhU6BBYLOb8ZtXJ/HV0o/vPKszJc9H8
B1rxaPaHG921S2B04b1hw0aBvARyfJ6d8So78H/EoIwIzUXAWafGrHeBazwEonXgacByOR8RW1qs
XbVmyoTVzC4dLDr6m04rgzdd1cFnv15L4Nqe7nIgP+ioeC1rNmAfoagC0PiVrOK9mNUeT/m9dXt2
ybiuvpno2XMv1bjo9LNfYFYBrJANyC16CiElOzVxm4DhxJpceBv1iUdKtoDw7gS4dfY45pJcrkB3
hJpj34HgrLbAX5J/xatMzMpyKdD0p51UkT5snVW1PMNXDkVtIipguf6U00JKYVHWPxbYdQjG2y3a
ltaPYCOfJ5iUKTW798JQEs0kHZXVIsGGMXzEQrNdN8BShKSUOQHh73kYjMs3r9afRwfda7P4c0uH
lr1tfmPxPsZg9q9Veqglf6H4Vc2pBgcvTGYaqS+NEfuMA/2crRp49GKnNiMaqlxYuOPwBF9BCsvC
8uLtPDG4/QqqHzSTiU36CRmPE4OfWCzRoThYW0VVSE+SOOJIYeucDyOvXn9wwMZMltnQfyRhBdeG
9Jdck15ctS/vb/C3bPe3f/XQV3OJXSC2UDHzEV2woRr/iNz7S/pTc856r4r2WwpXAnJq2nNtpYaa
oPZivObwbRCbkxtykeIU/wdVJ/RsWROImZD4tyDazOWIQMjOtwiqeBjb6ZVg6AAfM+nSDA1HzIbE
TfydymPptyr4f2DjSlqvozEjRbK07weKLcssxQ7ofzVbkYtVj8q4Jt1qfC1l9uuNbx10pyGfJr+4
H8ebew4SYrPgR1E0wtZFIm+8oYFu9um6rcb5+ZZKZDT1tcep8KYkS4nVhZ0zPDKwAwe7cjwc4ZUQ
p//PHQDlRr4ydMPUD9vv2xLrHMaTBgnUqhGBQe69Ajny31aBsvI4GOHE7+kg95sCXRuHc7i4GQ8d
siLo9BxaeihJc7GObYdrg0oLJ54flYh6ZxOggDOzE95dPaIUh3sIa3OnOJdnj7G77UfvtFrEdg+9
RsthrLcjnfVB8lDcCxEzNqbynhxUzmzAAOlHodrtGPNgii28fUmmJGXM2OPKfKcmaQ6b8MhgEDji
3ARVWSWPZcxBcPpeRRoIg6YwoXJCm4BeBjG1/n/DGHx5qM2QY/dEsO5qKgyYBfjxpxkm0T3X6hzD
rNYBcHEvxpXjLmDCFYjXGVCU6wnd3URE15g5nho4T0plVQUyPUFbSPqcxvUd2jlp7Nu50mhjfZ/O
8/VRxl9Uhq5k6HD2yvGRgoaSlJd4axS6zAayLZbxtmGs2EaahFqX5nnJBE8dchYJ9LKHXfDP8fNT
a9wlvvk/59ERjehYbq9nNKddZWvDK2D9VWfb9UXvLG8eEW3HDKPwOBET2ecerX1RUic4mKW1Do/K
SG/qXyIs2YC2mICVOh3MFtzxK1pYzsnv4LmX+I0+cnDq6Vn7Q0ucwlDEwH74N9bOWk9OOv+Igmwy
XrMYLX4CPp5JrH2dTavRoiQo6Oi4R6zQxs9tXCWj30q1b1EgNo9IdpcfmFO7pkcRrPj8QLRJ6Dsd
hdHfpVVdB8G9j65nN0hRq0brBe/y7IKmItTGt7CF6YsHSmWUQ27Ivd1EC6ys/vJXJI0jMoJp6XFP
qk/P3YEw1uwPfvLK1CVHCp7nY3kd0yXCIWOizKSNUwegxNuuY8U3CL+KUGXPxRG1KZlGBB4xQQh8
NQjavuyurLf8BZqiuJLRXR8jG6pOEvBeuHTHNnOErs0nGXRx1g9PhJ0ZYY7FhClrcyWwcr1iXKpJ
htiJkpo6hE7j+D6oFX9VwbSAGQ8+Qta1ofuq7KALwdYa9LDz0IuMWW7VrNgdGeQCqSGm1oI/20tM
/m6hUn4Nk8cqkcXq6RUyR9CA0XZVrrQId44wjpWUpKChNVd9ZY7sGBwtTSXafddDzmLkhQcm9Lil
YBJ6GPkNEofSLziDDYlYomydJOFZ+VKTNu1p14eiHWsCbJggEqJIDf2x3feGA6He+r5OAE381M6F
lnM6JxQbOE2pjmPX9P9Uxgf7f+vyZNCfC5NIlD3oR3y91ThB8f/I/73UO9G4dmhMJK1IgbMbu/X5
c0BSKTmdWU8kKHs0ly7HcoM9ckoi1BgZ0qw+pDC7Yvjytc12rNXef65oUKeVNHWNF+4ZwQ1jok0c
z/weTdHxOU59rydb4SaMlwF+rtPwSAwfXlFybzkO0UWuRJCmQyvz2N3m19XtyOzrf+U+zmRFE63q
kfdIasyfJzRHCU4ZKkclFOAasK9DF5TGN0mRliTzojk4NZxNhlVIiaCkdzXAHPpR0QUYtJRwsg0Z
Ck7xr67RXwh++mL56ZZ0+jeD/XAxHV0j8ONn3CwyhRFoN4r8FWpQ0rKsCqF9EjZrgqViFgoMAqVD
5FtGLli5p7m8U8o87FLlMQ5p10h5RfOM8vydAXc+21BCVJOta7iVzgXxaRcKvmGMDL3lMOoR/i6z
MGJN76v4QXQPhuFdnpqpTdfOIypwqGiKrtSdKpAw0UEWSPrBvp2PApNRqeSjiLw3mfkaUTIOvCxd
CJtlmS5dxRmiyx9ozzHzcqtfwaCugs1q7DVoloBgXnQo2OPzjQHPI0Mc5u1V1xIO+oN1u4qmyzz6
/puLR9Jr4ZfRvtVRK0tzwqmEL1QGNNYWXzZQ/v62mCoRV3t4q9o8todjuPUI2jNAh5OsCGJR6nP5
a7FBDe9etUIiZ+Wos9JikshM8t6WeXCykNvJpLwq+F39RG0EXFMcdfaxsJmNtT0rZQnBRV85Ej5M
cd18optTgspzU2dMa6mO5q3NIEVN+nVgf7qZpWGRrMEzt2QBFUVaRnhgw6IbTI6206sZ6mI1lViS
p1rRRuzfP4xn72Tx+XB29E6WGZQkKjys+b71MN987ecM7U4D/xSnhqkt+NeGQqXWnTOYM8nOjfcy
BbMuvnOOVTMLsbmsLsvjFXmSIk/0qsf2LU/jPGgG84l/9/DI8nKRrR+nYfCM43k8+iG92mb9gHzu
0IJo2vhrG6OfxEEf660vdOX9RR31JMd45HN3X//JEgkes5lQW1q7Rqs4AaeCZjSI+Xzi+/nWeeZI
k1mokHSasB/AlXAzjDVzym7FKncarPh5ufIxxQt85ghuDDBPyGD9VcHfmFX1Ch5Tlc/SBHai+tbm
YsnmUY/O5iaviwLNWTwWlUJx9iTh/ZWB9gUhag5gW29i06XW1//gPyPyaXZ80WAvX+tdN84gWKKP
OXXK52lnim/GRzOkEhGfXm8Bzwv33Akq4Xz0pNOiealX65hg/1/Ehy/J8DdiTUVOd1zwYNtCoAJL
ZQpj93AbIJneZjFsjkAl+DXJhUFw4yDf101GZfyAaIWZ/nlAUlEn+k0RRZIyYSCvS9fzvkIFRJqt
iB3Nkg44we/ZSq6qviSzMMTcxBRNzptSwsnstZ6yGP2CUD9z7YIXAnfqlOXOR03Sag1xqEy3xG8G
WG2hcdoUGnTngvT/H8+9ies+BAM5dvmtlIGGmCtG6Rp182SP9FK5YseUoLV+8J2AU/b44xm2kxX6
E1xzKN5pQcpM67tcb5EMFBqC5ut8/dpyJTf9paY3VEi+5N+A2a9Rj1aW3EI0/4pgic6fH7Alo5F3
PJunWezSKeN/bAcb/s0CVMVfLg6vqY7THXvnE375xyZxTupzeoWPaE8dBu6UJyJy2l/mPxY5q6qt
ubf4107IhMfmHbjfwNd2i6vTKtr78H9ZhGJ/5TFzBcg8It3M+fjMvn2+XawFzEB/grJoXu4bZY4X
qNegah5TMUVdGVzCqMXNk+ojq2oxeoT8ImdEcn04QGIV0VVPH1C3CtnuLsnlNmYLGYAS+IoNyCfh
0Wm3M8hut5u/YL8gUn0dspbpvtCah8YSv3RWqL3HSmCrZNFbSU2gAENaKxjLYXKHsUlgWupUXDG+
v09AXiP68OFXoWTzZCOiJaUPs761Fg0s5NvUyQQ2nSl4ViPIVLr4ft1MpmC7KGRyZbquIIvyLRJI
+m8flyiJHY8MnJgknlvqU+6lqmureLtfY7Dv4P0n68AwaK1zWOAeJXfuRlS5yd1vyZ5Eu8HDTk0c
4aJuON4+MeqPE5rXub7m7coPAdRSoG6UwGldpLG+IUWHGFrYWCs7co2cBXPMVwW/xf7Idob1L76+
BwYY+xUW/xN+rIFz6i1HwR1ISe+KHOpDHVwN5ThMJAphqnaA0euWU5QutDWfmJs+OuhWCcxsAXns
jaVRvUwUO0mJPvJSZeNhHFFGSQLZfL7sUsrLRBAUJ8OWpbJWwbewsapb7uiVZtl+MxsGvC59OwuG
sCDXFhhV2BSGcEF759LV4mDaidxgotQyaigEYvkf4SWOAe1GdjoWEC7jcZoSYrFEZTCgYrD0PSm6
6TAemrZYYzEP1qJgxm9BD/D5ANghpCY1nPibhd2DXUq1BxzGPp047Z4SHez26zimbRdu4ngwEuoZ
gcQfFBfE+XCGjWjRkmHNmvLX4q3fsr7B7kpj6Dv+S8cMTCVqXGJnxTyvXVmqmEzmZEMMD2M8RIGu
purrYm9oNM4mfzmRyOI1gul3xAe2s5mSLEWrl9TNYTGKUCas6Voi4aJIMgppXfBWI+ARoM7tCWpW
6neOVwWKbStjtTBdXsSoOl0WUfFSEyHxPmWgJcIgrihBQF+ZokwHHZr8UOICOWl1qJQQQct3gQvl
lX6MAYymxOk5k7MloGofPpLPHIHS/Ptpj76+ER5GD61PYuPeqI1YpGZmE0r5TgYN4zq3DKotBnA5
JRz9p76tnmQ6/i6GEtqrJGVgtjA3liuMmPAeH6XtwKBnvxf8+5wx0B8TWLDuzqCfObKVEzHy1uz7
IeahDn5QbbUytER8/FtRXP5A0auL+wO5Pm4Wi+AeXrqzZqrqtzu+AuKzWdGiqyJUbBrhYJoOlLJC
pVg5tsYyxGqTJocgF5nFxQJy8R4BKEEYTgy7tImAQ+8+O78gnZ86DLfc2D3lwX5Q8nETtqxr92sA
CkNWjlTfOorQvltK+42cHvvPH2FO6GV62Rf5U17hDfVEHmk88a3Erj8iXviiqlliGrs7/+8JJf5U
b08Y4ckwvHGPV4Qj+UF6siMLTuhmGQaqjhYdzDTSQEa96ji318MPNqSqeO03zTtle3o4BEe43pEb
2N2W5W6yXQcSt0NTgTCvVLmpsDgXCxrBDrOkS6mzqnGsN/OI4rOob2/Xfm+M99DwDesw7sAVUWgr
v89/lMX63EgsgzIUDrIwK6jFO+a7I9WM/pr1gyiSKaI8Qvee+YWOHr5hKZyW2y3l2yJybk2viVA5
jJXW8mZFQ94tBeiJjDHKJGw23qT6AWc876HG8vIWnR4cxD1orGO3D6+h41WrrcGUVDwrk2KZnuPn
emuMh0LXeZETBBmWHAEXzEhHWTgAxKYZjYrYhHdwP0XaKCGzqKwXdjIKdTwYgyeBbEflOzIw1Rnv
ZYENpnXZkY06XmcI0fEhIT52tirEJX+cd4Yfvma4SK/KrrgAi+kBlCAybkzAP3rJxcDaTWwJCgU/
76xgBA+Te+LGzH+J3y2QfZ68p05ApEegaoeFJzXfddXqaj0HfRNUFlPuetpMUe/MJyK7o2dGt2Qj
9+6Yrdz44LfFxmRcOzFdaaK7IDCfNFFfV9Cjlrb0PDqoMUthWu92kDyglbfNSlABdfPU80CxX0e/
epgLmwcBlhmrccIhwikxCxQRWjjDiHNBvn5dpBru/ZkI7gfSk2LaOInTHXnwel28e/34Hs1ai9Kc
Tv9r7/ckc8P2C/3U4n4wO/uEPDmPdUgMnUNh6gIn5Sysx3c1iYTdGstVtvj2QfWKYdjetTzfgN1m
TxeyCO6MRee5KmSE9witzhisAEJ1zxH380fpXDLE8bcFzMmmIBBe96D9FIbgKQMtz0qXYO6BXKSu
fjdAUXsQrztkTeVSRcH4u0XaqChvfiiNQjXhefqIlvs/8Hzirz/nYGC5zAfGfBlWqhLwGpJsjISL
Ozg4rZ2bU4MYA2ex2k5btaWXO3gHARpXF2ohJwovMBYVLrbOtZt+lYsnqinxEuY8qcDUpilCMzLl
ueVa0UTWNY74rLPrfFbIYip3fGCIwz8zvG/uMU1IuOUGlGMDVHGqK4B2VDbMB9L7/dnnpSXn/Y8o
Cik0LIBhwghO6FBHy+/EIvVv18w6oswuedNQk77gIhd+v5Qs816rJ5qcB5xuK4OtjIiNTQyi0URA
HteIb4XqD+LbHdoxK51xY0AoxRUzNLDAgbzuQ22PHwFgFduTEsV6wGFC2RA4753LegfomaUnY80G
C3Sk8FU4BJRm/53t15kOr/OvQsc3I/kXZP98Hk3uBpSFowDhM0ohNsGS86GGr8mlm5KFBwGgZe0S
PRnshYllCZKmxcPD1RVxDn+03th5Ghtp5DwP0OswrbfwVpspuFgjL9z4jW49MTtMwYaqLWOEU2NR
km5WwZDNIe2IaSU6Q/P8wLqRpN+6GvLzzLFKl1OW4lEdTWr6gk9FKDIyXkxA8dtou/VGxuW9kx3i
fpGuKE575YKVGbMBVT3ho7QjYd6PYizCXV6pWTN++4Y+MDo61f2ye4ooLtUBWgiv1v4YVUiGp5XO
04/mLPZY0fksmGnErWjBSSL3ZqYkU54gRMKoWNKL55kWlGFqJOQMshIGm0m8/94JdGtLUZHNB7lJ
FJsaYC2tPbrUH4TIwLAnMWtFoCHV0LggNNqWUm3ifpfpvoT9o2SdFkJDXD562/B2jXZezAIv7PfW
CRYWMyrvmHVX9LNSndRi2GiaggO6CEg8rVXYIBBUeotiD3MY/taGNWRCJeroX2KXYpg0uSf6WsMI
ZCXHLO7wqq2do1aknWbhw6zrxpVoZXOs5PId1HItCJfuQWOOvzEp4whVoEBZh3HQecZEFqLdOkzn
ES2iNO1kUG5CQjFasAiuQeqEZbdlOn1uuUZYkhFWXRx+rYqcSfRKFpaUzDu45Bt2ALt+k/Y4N90z
/z2hq/WyhsVTtBHRMdOwv8B2HDjjLB2dbeKV/Sdan+uaCE7o4cKGHCqUEz/mdYoBIrfLOYuN9dFF
/duF+Fp7sIjNgCOs6EVluSZ7JvfGIYjDmNLfPKg/7ATb1r2Ir46QUC5KW7F0WGKEhR8Gn6Qm+qLw
9JA7hj0q5n6f99ux9N89hzNp72vzBuWmXF8azJufLrneJPBB3B+qUkHZKFeVLXcplqiFQ0URBQ0T
o0Ro5ezyE4w8nVt5nsuKYMUbqa7/EaUO1mhTqxKez2mtqyI8R8izy/n0XSDvFrsfsWIWiKlfqJRC
9AzKH6CzygVMHpDG+lMYHQ/aEn/Yom4IMLMo2X8BrJKk15j0129ufWryg5F45jmS5rmx8viVLedM
M7gGq66Ne5Ui+Lsm8tNyXdANObern06v4nhJvGaBq9AgLg1by4IwLCScXBmmy5Lmpmyta4N3ceKu
UpCE6yDr5d2uEKapyt5oi/SDTripvwgTUJJMw7K4/uc+1ZSV0tuwNq8b2ig3Jt74kqvWIBxg0dsk
B1a1cA/l3ZG4MX8MUPgO1L8w66PqILyn47LKnW7kVxKQPOy0nGZ6XdQsGFavkGBxajw9dWT6H7Vc
38Sc+kTA+R0JTSSjvGx/QY1txcUAYdcHMc2Ti06kx97ERGqcborJESzyIamnxVuly8o+PZtgNLIp
Vl6qVBnrntRbjLHEr8+pIap+Gm4BJIx4mFawzRjfEkeRyPc0lNcG8ITXiOnBNzpPLCJRWSoQkCRS
rB85nD8GRvAG8Adz+IaOqqPwykhwSZ+OK8pAR90yatDHZQ5zkYDIHKuGej38+sXzYii8H4FDEvbD
yg94bJSyBhMbH6uieb+rQo7Mqwz9XVBSzNPiqgF9inVUYvUHtsllCB3LIoNFr7fIQZl9+NuK+Mb0
g2dPR1YOsW6HCh99U0vKzqCfLLk7V28z4k9oS4rxFvaz9btPKxkJcQba2e5nF6Y9TmCnjzpXrJOY
IqywoMUHc02ypXEaTdStBXmC+S53JJKOWtjP7SRIxdzb6M8FlaLukabwW+6PY0cWiT2//BA2Tzwr
pdVArSSAZ5aViRkU5RQ1YaQ0e0CDXRVXGuBhYBuXOniPj1XMIGaE6Xcgctk5QJF79mXhwhZ8vBol
9PfWbdhwnUHPe1AvoZhPIUk+LHF3ewTwZL4InrGrrrrD0cjhoTmfg0Sz4MYGCwSC/IEqlksDfBFf
MfdDpu7YLltZUSlHd5CasXLAcDxVrno9umTfpWvJglIsHBpkOvKWPF74DP7IdkK8OieLDDAbMgsC
EzNu0PYaXl1vD7VWWLobbVkwEtirvG31y85uvOr5MKizped2n74b8Dh2fAmorv2IZz40zUWehuET
/eguWepD+EA0TZKQ8T/abHy7XNHAwgoQpdgAEkQXzAzUDQs4b5AP23EkkL+rHVs85sUy5qAONXsQ
qg1ZVgDXHVLErys41U4KVF48XBn0VWxVN1pduaUiDtDChtIVweaGvTkxLbUxiO9m3rl0EDLIdT7b
NFKoGgJFvs935TcqfFEZk8CYNpYQS8/v4sRugt/mSIaayChtSDkxbfvlo5xKTTVY/Ufum5C9ESLr
jnEr3z44i4CjYaCFrWg305BJzuiu8qI60rMZ67+7GDuhr2fcZA0A6C6uBVU1U8bqMqTuYLXqvTu2
3I578wxii1+FBmKYIVbdGBYBDQC0Mb/aLozw1DY8GShU5qeQ1IVqNLciluPl4FXVXYjyKO9m3GAI
OsLUHbgZFTC7vIsqZPUga2lPy5/1Q/T0NQqmRqRy7Ws2aEGi8z5ANaqnUcdtkDD/aCx7DW1LS1ov
oHk3n9B7+2cme/KHghjqG9WX+BD5MFmM4uaf1wxRFKL3HhRaTqVjvA/rNmfWwuGTdro6LPcj4AZu
0txYjYtZfIgNQUWR+zmY3aJ7Rv0f00//77BR4iDQxDvMqnCPJcb+/YJXDSxEW8qY1Cpr4aa8NVnr
ZGLNtbtdNPML2fdki/fkVXv1KWEE/tb3mj8oxiVQS5ncU15YW2d3rz52qbdNdnjn3k6IxeSjYECK
CZlAfrF4/c+tpmIT09XWw9ThPqdEX/Az15yIRvck2wGEIzc4PisdrG6wpzYz0fyg/bXmfnaN1FnK
4LxAAPgVWY24h3dtGjaXO1pPIC10Ai+uxnuSF6Thhxs2uSNqXTjoJVQKDEzUGu3EnkJHp1quI6NY
OwIRV4QWocdIvJbW9JFumjxEDcEL8+UHi9l3q+KD68iNeddAvkVyzCtXWircOKs5dm1EMscVldQQ
rr8lMZr1Q9wVHdDxWOysmHgB65BK1SBSv/s6kFAVR1x2G8tn4yHNAJou+f7PIFaiycPoKo8cLPdv
ROA18naVt88HrGC+CWw8hD6Uxjiwf0pciiY+u0ZfYaWtsRtwjQvQ5NYzwY5c4fFhHuaPcmNmCsLW
H6OuaJvGkh6G98EU02HoRumFADltAczsh5NaULDV0s+9kSORxsNaPBzlp2guHD5HeJhYhakIQwzv
HwUAF+b9cD0ToXGdYGJxctVUUTRAbPiJ1wciycut7MSIMewRPoSdRTLKyiv9eU9a1XMl/EMXY0FZ
q8zPxm3UaBEOZqJICsORgZ9R5Y2sp3Afpw3LR/+ip0iEHX7PiCBqBfl9r9Mi63B9UOQJ/gxWjDtM
VPzWegErZKv81NZuOOEoLobxHMAX9PvZy3rsFbWu1woLi0xJWkgvIv5aEjxp6M3uGq3lI/Ck9Mlk
ipMD8oi8GpLbeQGVY/AKcNx4nNhyyW5rFHkJuZlI5izqPLruZxEf7xSFn6xW0Mg8mt5rjB8uN/yj
tLFpG2OAnI/NYO6GxKE+t79voIE/UrgQ5DDiwuGRbNdM1yNxcGO8R0JiDX3CQLw+SN0UesiHYYol
kGpWtZu8IxbRMVRj6vFZeNuxTyoo/Q7t/CfdgqsKeBeNkv9EM9lpIvrkc89441C6UlSexVzHLI4c
zsfadpKx3N1ng0YYPIa0pWTuuoex4tcGFc87uiAhJF7V29icfbDZEVpY7luJdA5BTZuKY/OKVDHK
r9dsYE0+dDLlJVI5FtfOljt3Tc3DmhcBFktsow5s553tEzSNih3WVOYvnzyRPNFVZvoXUsbn2HzG
j7ueTp+vXyunoNd0Ucwxo7l96CpJVzAf3Lg2cYuvivdtqvFNK2D7J0EWfM8qeZOdyK5GPTLLZTe6
6ZDJ+dwC1mN1f3YXBPwVxoUp0GuozBKSNUG4pMsHO6g7v+YTxNLnJMoLbb/80zQbtGIZDJ8+x3l6
dPPvAbgPIgaTbIZ8J+fG4ax/ME5FvtA1j1+MIQBFzwbxQZtwiBGMMlq1M/xBTQb6g4P2SfqNoUJu
sX+pJ8uCo+60lB8BPgVseVX0nP6+cIJyhVcjyHbYC2dn/4IHfbCeDD9JpCMdCtfK7s2/u4rLprQ7
/N3pEjtZnFqfRu0o22+IR5NmY1ot3E9GJQhQjs/Fr1lxKW/8mqT0vjMchf8XMKXDMACTT6ZtaFX1
NQxHmabdfb56TYB+t972skfAO6ETLXOEEvQEQ7uU0+2iSTv/bWCHopl8rbIurtNhhgYz/cIkk6Jv
PZcwnKxaDLT+pvIg9RrfviPclq3ejEE+nOZ4x+Z/QwcPTTrNBgTr1D1ptB9ew8TUmkDHncXTZwwY
z1Cfa2e9tDIYIYX9W+qQu6OZYgSRezAbw9w5cGr7R4rwIzP1CGUD4UYBcHAPiDmU3jcMfHl8/Mco
tzsgXUbiZ5ufjZEQSuzr88WgFrJY1MG/1RcbClroO9qi8qsCMW4dE1jxpALG1/jt0lRJZOubluVK
sI9ObXuSHbxh6E0WvP7l1FpX5zaZpT+YzDMTk2XhYoHcCEch75A/qrYMCBHRAIY2SsLG4U/x0/Ta
bdPjWo2nH1Rwm0Q7CL2E0C7fpBNdzMsuVDZ09BDHsn+f2VbOsH17qt04RxAHuRw6rVQFyaLC5j+N
KNt9HyiGoLAsgepGmVPXVzwK4HuP/RFVim+Xp9pgPNHoxTjbXXfwRzgMy35PL1th5ENl8q/bc/M/
6DYwrFjqdsXjs+pOPmq22tNk0rMFFYCLLDY2sykn/yl4M11fhEg7kNVzh3Cgve9jlCdCH8lW4uUH
e9tYqL5ptDQQ/7YiDkr2QqGZp/LIZeIoQhZQqbH3IxBFj2GIQoebCMBLWAO2HtqmuoDjDSGIF4EB
Qu3dc9j1Z9QBCeKjMeoGrus1I7yVNdPQ6nRdDOdswMzgNfcsHl+ybPHAdSH29Bo6/bp1K6G5HpzI
0RUUNuEWe7kl27mu4JOk/UKpZJ8FJtHMU7RZF+r362xxZ2RGzHf12Uq60yajxq7zNHoqqIPHdhFX
j3NyqIXA6rQHeRZ4R3om/G93wCSWvv2RMo0DEinyVjYl1arZMztIKZ8sdHdvtOFixpKsi9DeQqgG
N5zyYgVo1IdTeq7hFifsMeE6CjW+EdylA046LZFub5ua4IFHUxYmDrXglVL/0D711f+hrHiibgek
BcSgDRE9AD9bLSPyABqZZVAfGMWrcmX/jsZU2wnUsQwdL2VTtv+/UDK/SasS2XvIl6XqDHlTUjuE
Px4/3iDswCK57JnXnUasR8F6K5HuJPxmrKnZobEymamhmirXflUyvR0LHmrBesy3JENRi3yrEAkn
yR0BA+YG/AAbiA5P1YWEra2tudKG/SZToPn77cVQaVwOGo3tYY2p88TQsVQ2brBoTNsa40zsCkLW
2pINEagOp12Em4Ioc3BEdBaEkrZqplg031WtA0t/RB3+dlnwiZDRdqO902oKunSrcaQwOsdPPma6
BtTCerZnhyubq8YOTLlXX4lD+3EUZNshsH8Njj+frsJBtsIa/LGM/FUPSbH7bFpeQ10fBmuJQ6YH
ff9pkwxfrjWKtjUTDwBVfMRFzC4E5G2OVUEhVdY88DyjMPgUsOfCF1iKqtH7SzpjHX8SiPmPqrdy
tf4SqM/SdHMTB7YUzDzXPPfAlAvXQ+xYK2AbW/0CX6CekqHdWlSteYgzOkZahE5ZnclbdlfSRqw9
UGWJg7GlN6QcRPWLC3g4lXbGE5y/5qLqplD9xmFJGeFR8nIgWBUvoRGpjeIMSn43fO12kMsueFS8
Ldm89FAqpHPfqnzWH0zsNtu9ww7snCN+LBMt+iUAjAFHl3n5Gh68jJP02w4vmx1hRWLo2keRnpqo
IL6GaEzj3yAO7vvqQnCq7SkoILc6l/G0yi+7rbMGF14zaTwfouMDnX7o8WY/2Wc8PWWxY+jZlZaq
NQZe1AyiJfcWIguoCGYa6iggEE5XAA8SYB/4RVvT+5j2L7wDqkLRpq2CjG6lCQiEy5TORmSbS3//
WCOZKr+c3hIRSRiLjmd2NVxKWQOy0ZJKPP228a30PtwLuZbdP3M+6e7QqhRKdWEP23w9uPPoqjjk
prZhqSmXQc6Eua+9XEfZlNfuI5b668Wdqth18stl5wiqQjOJGWSYmLcGuLavMKlFF7m3qWtB9VLR
uIu2HPrg5rT3YKiR5NAt1EikGD6XPJx9zht5Rxzzg/PBVKVmD4bUT36BNEvFVYztwib1c3qtPDK+
CgOrYhon5D79on6621cDi7vYuZfigvqKZsJEvHY730XzY/8MCvWWhV1R3vK8LHKnnDZulXp0dPmn
Hr9HJeMM5zgI0iACGvOS8VfPYTfyIw4MeeSP36PA8WOr34MxPg1Li1F+omhYcy55vuRO9zkfCdYZ
Pkg6Q6QBxPywm34VHjSEwZJ+fm/E1gxm374D8RRnJcuNYdy95Ic5kyatZumJqv7eQAMlI4TJ6qKp
DEykvFixa5Q1Z5zkqIPPteMonxdl7i+Ts9LJvxGwigHnbE6DQuuOczzPHtG+rec377POk/4QWzzy
W+6YUQLH6EjZPGlxnvS/slteYGP4sAnnokhHsNwIHgc78+YktSbeAy6kouVF27qn6TtwGFilqkJP
QVFe0bgiJyzVdk7N4FKcMZqpQzj6RaOxRgF+QK9tm7HPObDRQ56p2GyQqKzmy47CMaiNLvwTQqrY
wxCzt5H2K01vBhC9pP/eORNCBDbrL7WVRAe9WNs3pw8T8HYq84qPhXvWSb6v2yFoh/abQXuNOGyu
91fB3W3TVOJ0SWj6+S2+/BuWrMDmrdNzPf7EmzMkAKEDE1h1Ykq6NLJDHTIf923B9I/XaDoU+Ag6
HnylxpvjMZ3WMDVDJ00wSKyTvBtGK/LFXvCexPxgAjwwGJ4CcDiK7uaRdxxe0baBStQfHLPYKIYU
yObBBsEK/l/d+sg4u8nt2uU+7WKhxDeLrpiQWhVlsKX6K52xEo+xpCUiaJGcmNabvcm5wqttSlx+
7Lw0cv1hEis1Ko8UMV+LxP2o/OjPBAtErCZbF7lzFrBcZdyO1iSVczRjlRl0JS25ayQU1BXm9AHS
tHvGihtTPQFBoYgazDmBkOpfG5YjCQIV3TVdDwfaufmZo1MhBpiwKfhwQpQflEjrxQUTqBLR8+L7
xPWQ3QBTzGY/TBs2m9ncmuSsCQe7mDaXKIg3WZWT9D7iAlbA0c+P1DbRvAYZ3NZ8sNKBYDtqFW1D
XRKUpNIR5BccJTp+g83kr/G5o3NTPaPL2733ShGLgKZvQUMjwjvx9Drbc2zJlhoy1zCl33R3nwzu
A0wLsyzk9xFiQJL9fOouFu4IAqjFGfZqbamn0rJwuKtFt368EpY4RQjA5s224R2F5EtDl1Bmmx6+
huqIbIFt3nMdsXEmqtXRcAP8aiD2Xh7vqlmEM0neW6+TkLvkxs3sRiv8oMJbz9VMockxW7PiN4Kd
wE8fjS0168IGE/pNKpc5M9Hso/q7VkI9qwSgE7WsxpKDauG5f03Md/lA2Cfr+guzskehXKIK+8rN
LijLAaD+yO7F4U3+2TSNNgwT6yuqmeaF4RI6BcNtuF71gvx3YuLVYREfY11ByekiOel5+MC+vqds
Ro33yXnB+SWxtpKyw1Gb7FWoqbJbmprD6PbIIxTLicrLiAsZsUycDDoXexhprzC3mc76zRweFj2T
fFGkJygvsIpqxcgWSt435+aeLZjGyitv/FEJGXl6yBXO0L4SqXSYLWmre6EAfSJ7y1IHJ25fG3PQ
V3Zlgex0Z5AbYHmX0b6idfoyo/gUG0dVI1XpsBeHcJQHCPIynXxKsahol7+6X8vhqD2xEMifnccJ
HhAkQksvVeMMQJHfcZWrWqYqi1tuz3rn8OUyDknndcOYJ9xfd1iSvmfaeoBv9kwLYdSVT/D24Wlf
raAIm+rxtBAOWDVxJEzNXD/cGr2HlN0uH4hHQwi+ZVxiDpr6vwy7gpGZl7K7UK54ibabxbgRo/Lx
A0ZSR+uM0K/E0iv8iGpUgCW134ua08scYpev7BHaaiYfwXGxrmxwDGwUTgvMsDgoeJBUYE4Cy8ys
wIq7O02MAGchOejB7lH78fLGUwdi5zkqdPxDQN4zwzy83uS0ximrwU4ZIqyto77nub+LeczgwT1z
Wi0stBCS63A1T8W7cf+GIpj7mwyFgBWiZ/CgC13SiDQHCBLKoTepuzLW5qyPZwDpI4ihJAAwGC+Z
2I95G5pp7iYRtMlaF1d16f35osnspaCg2CBRbxIbJSNEY3zpCyuFT3S+cYIVETCEFl9wdMpQQ1oy
JCcqv0sSfgZjFTuMSBhQQovdtFWOpVO0O1AApn6/1ECG57W9Hf5rfzYdLWRiTTeqrXbZT1ROBgzS
cD+eyEVpXL0Ar43QmROllafqk+kfs5D8xNHJFCAlYMgchj458pSn2G6eTRSnYTR2ZQ5YOFcTeAhd
baSYGlj2op9YrIzsNyp2HcLQIvQdaqqQD0usl3aGtRjxVDcHb+ExFG9eKpv59TYbtotT06MB4Da4
lyUCeNY2kKlVKPf1iqY1uswGYj6FpMSmNyvLTKVwf5Z+2W2zzQIb8xs83FZDAdMZI5kJNUEqmeS5
MGUcus75XMIguOU0qtNKLllfQfbYKiTblMJNGdO2BByc9fad3fka6fCpUN73HgHz9nhcAnAMBgcM
jOZ0XMb3kM1lvdU6nP9FXzCO9zkFGBW3VtQVTLx0m8HTxU/FSHeWaOrWRigVa9SsDzJjGqkOXtP1
NIiq3nKMc/ypbBpv+oCAlcYOi2wwC2dWxJ0627RZNUYVWVrWmRy3VihBQZj15kFEzmH+x1U6GqB+
fgZUrLQnovXH81pnqluXu7ltQa/2BgY1+6odojMGwrj3oPGgPnk+XrMkrOgYjPv3b0dg1r6QUvym
nBB1aJ2XXe5WL1I2aRYakWIb68cx2RmohqArvlY6PJQm1pNFgFPOz0kVZpyhGMdjje7bIgEsxmFI
A6HKLgRA3S0rioTIMOTyU6B8gOEPtLzDY3DsWnkr1KBfJyzZkV4fZ2xuyLRU816MaTsBsESsr1Nt
oxvUPwVJSC5TZTVgeu8EYHheeQGlVpn0RJ41fJmpXJ4YsPZPEME57pOrjL83K9wEvrvFH8j8He+4
193L0iyUgy93LbANFVSYFjlykUDZ/yMbt5vcEKZk4n/wRIMq+SS10e0Pqe8LCncEQ9ZMTb1pJ73d
SnOaqyU867V2u0xvWv7t+j6xcgQzrGz30Tjf5otPkiGjjYXoYFt5Cl+Xu+yyB5F9cv+MDOoExozo
im/v36zfNpne6E75Zt7z8eeLCIm7x9xdoBWQCzPKMd65Ja3gd533Sa+12SUQvk23JKa+yPjyyaFr
dEEakXnGwZOO5vqY3PJ61xiqFH1nZoJ+n31eyBXbuhoY5ewZJh7koXLjTiNhXdt8ERuvRKXASU/m
IbweEm74wpu8AiLPrHh9Yd/F4xt24d4qWX9EplDXO0AOd900WVwFyos9sbP+kIRqdgzsR5oUrJle
BG1r6QoYRAG1zUd1Rv7yeIABtUCLVxxocheKteMCursoi3wcWhF//PWBqwoQDApVt1GQeE1UpvNQ
xNeEPWbcKuSj41OSN5OXbI6Byr+eq/upkr5JJ79VbQCtInuna3jnCmjZqYkGCzofcDHG6+KxXHKW
g7q+t2bXE8d7nupCklGjBNEhmCGNyryyI1CVj84Q/DKTwztLEa8vfE/y7FvxvZOzawfRpJQPa5Jr
BV7spWxVH/c1xpTLRpmENDXOWFo/qqeGdUslqh2vToV2ENiBU4+ZzChm5VZGHhu5Yhf7/EgcjSDp
XBOqtanXRnTjzJMfBSgbLdnpfqY6m3Bofqk01xTwcwSuKcPPdL4FKhR61RyNOuh9DCVnlxibQYeS
kHDvKV3pZkDz9L939Pn7rLI1miBpjOaxLdloWg7SjjtKSO/pBUvlph2sAEjRitFDNcA/W+WelCiB
3lPtu18xzL+6PYEREyhVC2AvAtCzT7cQiXNXEIs/rK3MHuaMyZZd9EII9CjBOz7As78+v4CGw+av
QGAXwtx/A940Hj+DrhuSyvJHHlJ5KdhYWFXkcvxZjjKKKILjY4nsfzsVm+NLCnk06wgS3dNoYZpf
H0+9UMVutUwwVgnLLlblxEje10q3zzzIpvMdGHPw3ByIqFG2aj+AAXY5rnVl0WszwQrhtIiiGhyP
C2A40kk9Q5BSig1y8RudUcL8J9R0ZrD6bNw3VMWey5rgYfwRpNivvAOqSFktdqR1P7SohNDXXDWh
EqwGTqrbWucLGHV9BdQuwTRsxAhKfWTyOE0IVPDrA7nQ1Zo/s5c7vAoncYBXjQSxb/+D7p+Tu78N
5kCfasCdK75Os8OFsBIv7P+uvH+flGKHA6pOSV0pT9ysJytZ3o/TihCaMR/DS8mV4CN2n/4cPTYQ
WMaG3RclDkKmg0bx6jY4x1thonpt8RR8Ejuhg15niwzxYjDIqKlD6C24zfrprYxyJFHBQvcieQYo
60+GptpeUpLyU6VnPuZOrF5ZOOYNA80jHELntmsu3CfOr/n4YkvZHlCMBYycT1GhWfGXdmQ5JcmM
JM/rCBhcY6H/H43NIEtBQL0zPP7ksUOl+0YXs63zCTtUMvOHZxL45MVpa5eJnE+qEP8za/WNT18U
3w9f2BtpPcGeuO8WibB0UVt/RqHbndN48AfutX1pHu2/r9kJy1+N7uRx+NWF/FFR3px/aUnaPIqX
QQsOUjIL+MqWuv6/9vehVvq4ajW2IWjRyTrwUw80ZY3+vNtmYjqrrhG+TFxjhNXH6no3Vq/0D8tH
EpjiWrOp8CPY8Luwa+g0FDydZslRFjxz+U7zAIh9aDMjhNG1XL3rpQZFYz9T0ty68cdxuaq4d4qm
iPkzMBAWbhgUIq87Su/X9hjhhaMB206ZNg2wFNDBBSKwVWO9lvbi14rASkW8xuBwCp5/t7aKteHw
YxZyvxeR35vZUWt+zgBZ4H8GXpE1VfYILqM7d8SksUPPgviPd9TR84o79/r28B467vA0Fme4KEjI
Afoc5YvOFn4DiDGkl1yQJKzPbF3gn5JFB2y8IQHabIS7fqFZ4W/qHeWeLxbZS2RBorAg+5LsY5gr
GFQLMB7WkSXLqOh4GMFf6XEn/BrKIZLMrhUWH/cSz8lNKIVUVvb3/FzHVMJ4GP+uPUdlY4lE1/B2
L833BMCzoTOioxcL+JTcWEZUJEqFDHBpu06/l/g7vf2NoCru8bXmEkRBREzL5+HRaVOi2mPQhmGX
2+FuzW7qJqxTRj2VqRgUt4AJ9aVwj8lmYXXsnUK76oNY9GUb6StV/oyblMc9xVNq4UsBXCNDml2r
5gZHdBLizleprFtTM3AO9ieLJ7nRjxzuSMMwb76LxZiV/xcR0xBO4dZmAFczLB2I+8AYi5R/UhP/
ioPwrH7ycdBEAplJ9zjk8hW7KCJjvHLWtNecwhQ9BgdXyM+mHKGEUmGljWJCW4yvzqCj9ikCDK6+
03eMaRRj4Izgl8XdiuO8F6xc5yTU6ae417PinB5bIRYubggctCVDRXNbVBs+GCnCQZ6byFn7KFJe
NkL0TwP7Ud0Eml+IkghDV1cx4uaQfXM10IAx5lGKhgFShKVhqtdzh6MJ4yuNKnB8doJWU4CPI4o0
k8TX+MGHLdDff7qe2TK+PU66rlfYeBlEvzgTi3R/+hzZTxAUgh4u1kT7u08wYzwUAlNxR5kOW8u1
cGpXBpiTrzbV8l+myLw8sBiaVAwEthjUzAOe0GMQf4IH81UBcBzVT0P4LmHcTydnrPPrTKKAObZ8
8s9FRz7hUBUw7HNl8zhJEWuwJH0alCUyJovzk49uuQ2oQmsoUQM53FcwLUln6G3lBZtb1K4pA+/k
KunQNBU5VusdwIs3cQKlrI49e6cIMHCJOjbd4GXmfCR6rM7W0n0TmF106KGQz+gcVjbwuw46aPq9
D7LkKJh2+eJpRjnNafSCQvMSOHaaBvRNu7Mzfs4vkTjt3dIc4K4i41ADiF/05hmgKF/QrYiC4ii8
L0NfeEJfkvd4/5dqviDvtGTX8ICmUnzrLrQgNmCxDlrBW5Xj+NLMpFN4gUmWX+aqL7zP7ClWxE/M
iq+208ZojJk1JjwrnlRONS0ybt3NuwQnL62AU25D7+JvByAxWCNtiEzoetcXf+K2NijADdir70JC
Q0P4aoFNnBtLpd/jxddghv9Fj5eS1LT6bh0kLjnUoA0TQMF1kUFZhA/YmNFtx81nhmUK9YsM0oXi
uSMM6ocSAT3sUFpIijpZsPaX2xIu0wyGM/KzlvxwrBjNlrssBTM/4WRBW4Oz3BGNOiE3Q24YAkRM
9AMAssHpnb4EYklCDO+ra7LP1xQS/nDGpxX9hopCrZAKDUVD8ji2CDg4oD6U8BQy5oWYIYE/FUA4
rroZV6tnCVtff1/9ooRew4Z9Uk440rrx/ssZVRNK2pBI0pTl9mhv6yUzaNCVEfxY/F+u2webbqnj
w7lN5Eh9/LW0cekBe7wqwTiGCe7+MIRj6SW9b3rA/kjU5oG8o47Te/Jn/6WA1vnHl+ohFfKtVRFk
Ffxhhbo2Kjeuc78sBHD3W2BLmeSMVZQIqcDF8+gOQpOVG6oxu7E17Ce3TTHdvokv2ZUwJFRJ2Iho
JXTmbRbXvL9FJ3ysRaCu6PKHtxWAQs1lQN0t4SL+kW7/CIHpyy7GzZkSM9i1uvGI0ZVnm+0cB3s/
yCTZob7MKqotqo4XXaBij5PHCY8Uq15bHENyspN5kOkWPJrohJghFeMinS8mQY/4NSLy7D53Q3Me
dsOloKXc2B12os85lUQMVjAARkzqhaJvdwSjNb5rMR7nnyW9BxxQfqWm4TPlvn/L2Ab6iWCkNfow
4h/Kn4AUwf6a14sbac/tt1i9Xft5Ey5NqGLFlRPtVK0oo4abwzO1bmlTrABPcGt75pGfBiPeLLpG
fhsBAtl3ikM5P+dcX654uTxCx+eqlgtjI8bLd5KVVyUo/zega6gF5bPyBPC01CdVRFv2BTl57A+o
FJBDRNa5JRnjbqnA+a6ztoj2YKOG5cNX3paFrQBThFg2mMG5FbWnqs3XrWF6Xfhi0szFJPIqkXXs
sOCTf1fj6RxcomORA/xYW72AtNdijJ1TcTCmjiUjK5HVPUqtVhOCKwX1T6d+MW+I2dHrzigogwLm
s9KEyd3b442QyApGiHFg+GuIGgl/jDwOWuvM/TBOihr3CEdJhESv6O41neYijqFhbHKg9gDmWIBP
CnEcddUmpaXDMY3Uj93FpJGimfiLeNf2C9/mbq/qgqqq0wWv2aCDo73Jd2X1nC3HJNJywzKbF6AF
HSNVLXGUk7aMlcCAbzmJpgi1e0igUSZT2gIQDHhZxHNRoyd6zYCXEshb2xSxx1iGJk4z/OQKRSq1
MsYId55swDE+0zhISb6SzImnpnwx0RGa7H4qnn42tiByJky5LLHWgy/dH7KFJj0AxOJdNcfu0/1m
g5bntPBKmNmQVN5oJiMguAcg4ylN1O/+GLswWhwToOYpqnvqAl6UkHVqSMp8oLnljXGwEON+eDyY
nQpLsZ04klGyl7xihkTs6FHhKe12gqGPQBMUFouMVlbaIreW//2djHCcYxStmqAnqe54/AJTrCpr
Cu7mkNgfHI7DdfdlUiz0dK6qv2ydH461kSrXJfpr7DKXck/ukbYZjjTND/iNvDb/Hha+gJiKud+k
inLJm5PY4JF9ZUoX5lkxyjTlOof/yIi6fmbZfPS4CMbGNPya45RBWvjmvJYVOYpYFELtUgat23AR
Ai9nbbAc9C5HwlfivsOkl1jZ69BGr5vD1EG6pcEX1ow1tXD/pOy2DcCqtJRshYpEniGapTQdvNpm
ULyNbgI+vxfuqes9T8ZwAf6xwT97VGl3TTj2/X7646yGlkZqgO2HpGdzIcEQ0VBgZenuliquSU1B
9ajCba4GAybqlTzUKtj+2Q2CR3M/Rs4SJIa1VSiTwfbmiPTSiXvlShnSbCJqOaf6aFCfsomQtSw/
6tQ7E69xZlaZmHyYloriSYvezyl2eVHYAQ2US5MGWzKWqk1n/DF0EbpyCXfzCxeslgJocXpOodE8
DRHOwqn3BHyx8lzUU25yqOGt10xS1qPUWdFYxqTqyEnUXIRWMaxbOS4mNHnKrZqIZRR4lnr9kdeP
yaCCfuRJymBY8El3AmpR8LFKlbD6LHOdkeNZyZTQN6VIKvhI6lVAtJltoXXazsuWxouSKCQJn97s
x5CV+y40x6V5In661NtY1c569QabgAc4F1WOkrfpYuMh4sN4zl92WUR09DfkmfeGqsf7KiW8bHlP
1ZQ4GwgHMK3FZrSNL5u6B8OysGjnLvbjnjagAIExl88NpcPVi/tbt4/0IAH3sFA4fTYl9Hb89/5N
k+yyVRmkRtngyPvFxoeQ9et/Is6i0HXXPbL2gwIXsMZAslJbXSvRELLl64v0MrFn67KA+SEEf4K8
u/pskwCWrmZNwVcOT25ELKZf2wokDHEvhCE6wxD7dO/MQEj5KBu90dS5aF53J8qVYWY2wC8BwpWn
14wDB5dytsviOpNBPnwqs5oI68Lkfz8Ex6jU/c/tf9a33ykJJcpJUsMrtVNZlPz00kSkaXNNTvty
cZcS7jrAiPOLZymfOq0KIORT6Szi+XnQR86xYe5TsFyrzshrfe+3YdRUkz9gtEWjlQ21o4yGAF8H
nxVyk83h7e5ke4ei3OcMYJ8pkEZSzUNpVOOSpyOe0DcM/fA9sS/cKrD7ALbFn2PWA2b7snDv8jdg
kK11zI7ZBD96Kqqo5c+W7tJkfvmMowhaTWbZhAhAcD8SPdFxvHHmn291O87txQkTL87zBiHJsRgz
0DnTo0Afh5L6UDPrFnij/oUwHyRi3ovcnNGyd3ItHpXPBEpDqGrclHWwXwD6Imrei1AGJBxSrGni
mNbkGdAt5/NXNG75tUlI/UHT1LeQ5g+E6W8BxjtyFs1j9T74/GOSD6vtcSTSBX4MqoMFl6bMnc0F
5x5ICFh6DJCN5IkOUcGasjILZpwTVsyhrFf2kOf9oKLqtJdz8GP9Pk7b5NEpisXH6vWgSejg5yk/
B9OlIGY8JbipLgXcglBpBxiQOx9Wd3OxcZ79c6i6T6S+NzEuxj/0OltP/G2+oQTnMcqnCdB6hNI5
ESiA8IMTjLn+9tDVNKsjsmwX7/QQH3DYCTiOYu2qnBRDPlf/OvXWkY/NB7IO7CypBawZDRRz1C2u
9elv7TklcktomfBZDo1J/4I6x6t3MzluL0hijubshF3rO2fkulO4vS0bibwyv5G4HdaM8FzZkGXe
G2dlHJ6+Ws5oLr97dFw43l5eqqEXj4V7YfabfO6ZbJIiYZwMPjZHY8yr/4Ooom/yGj3zA1Z6+a6I
lKRkhQxDF2inoYKzXS1fTVmqq6U702jkxVaXnwNISMexcRy4eAhr8YTyKdTwAVoGLtjkNWnOUwMR
qBJoCcTWLKrjGzzEenRKTJxzxczvD1ePqklsjedb+oASNGp6NC8VI40DndGlk7pBB7spP5Cyns8w
J9uYVEr5zTnSIO1TVu5hjMbwfZMnX1TmKZQdRoD6QkW4tcIs53iLbEh5MhjzJGeldEOlYZTqCUz3
3R/sxDCzi7LATbZYnwRmpijFnm98BpBn3bfNO65Vnlf0fd7/hASQ3ZZzrV8z9Fcc8z2zjGCMuNNv
2k6EUxfoVOSFtHbjlGDeOtnyIWtqHuge8uwLnXfuI4HkbL63FoZg656TRUOx4LdEx3SDN9jBhPwC
/b3sEmdQJIHr4Nod3wRihP9yvIRmTEqD55EesHGmcS+wVaMcw4pzxrgGILDyzbE8A+M6nnCz1HB5
ROAFV3/sKM9bMNoGKOea72bkSIxOmH0q1Q5yif4DwMf5URU/MePRw0cKBy+uqFt5gfboljEXh69J
vHocpVyD/6qShiDfLddojT0yA53Hp5eoUo+GdmH6VQ0nuHy8C94yGSlWPumPK5NTWYpbe3p+ezeC
Qfzvlm7B1EqvYVO6Qdfg63ae6UxohAllm8Rol4CdJkrrW+uxY4P7+mAYw2Zc/79u3TsGFvW9NAEg
eZGXIDK4goX0I2WBq+3ab/IHnBORZItnF2O65QzrZNy4RhfNsC+ddiAu7V7LgY06FTOR8CAiMKWJ
pTsW4Rdpxp/UXyx01iXns9hmT5G4w5byTBNNXQabmfZ67Cxl9LFPUJuNOEvb01FEW713v1ryMSxw
iY6TTfVr+VBMTLn2Z0fvro+gqy4+97SdXHD35uH9rDd4jvwx40jXoz3gCa6sazlF2ctiZbdHMbS/
cwtGc3Rntr5H1YVzd2chdT57cHCdHLrGFJjBX8r7jA/dWD0pJdxpLVlNfxY7OlUxsCL+cpAr5TAX
RqKjFeCeVcQpLQtm3LGnIJ9Ebd9qSEEw3FQn/F5dA34ET1RHU2O3aTL6FS6VgxrQj+aX7iPNdPsE
uoquCHQngSnYXsZUVoABX9EQGuoz37reIfOsQ0wvxtS67PPo7WZWgQkNvvnydXcbLXJCE0AuTGoY
TFM7tEB3/GH6c2QsR8N4B/fS+keyUbt/I/9cKT+zH7uIvgDYuQPClWDoMsbG2idFHJzMsmNj+H4U
OcZ5ou7mtRVQGcctPyW5LE2tOKKe5zYH6WsSF57N9rgTlVm3KBYcSJMJVa8IsJhCr6wfQm1MqXyi
bEskTgJmRE/VWsWF4/woqtQRsp84FsE5VnmXwp16XMEYZ/xrZSNa1P5hPCEUaubKK7iyofh7p2bp
hcFNdtNlNru3jJ7PJWaoKkrz/Cb6Ft3yCGL25mTn+yxx+OMQC0m6gr8yIgC60/PCL3IBLzcYBZ9Z
G8piidz30+rG5YEyapGSRQ12a4F6OJXGsJi6zK4UtoXNKzOWjMnbQTFmPhNSErHMkiXDhLM7s4WD
Jh+is58TcH60EYtQkWAOu3A3xnOsXicCvskdQxlay/Fc07uAPGp1unpMMOhzySZH1KxI8ZrMWG3A
p4PT3FcjOYitSG9bisSSN5sWJHypjY8bPRDYTguYoV0+NdRVoRa4o3WwF4EQeDo0kf2/k4X/WF1+
gJSmMaxyese0aE3Yc605Nf/ejSMsx4B8SoWHbwWz3Onr9xhovPWoQFofW8koKHmrA8EZtRNLoYLT
kwzLnQt1z3nNFoGLfkKTRenPGe620aEmCrMgOjwhVqVyY7cVYyMl4DO/QfETtAX3hyjnunOhHgi0
7FpGuCRgWz+w/D5yAKLHOGhVb6WyhdF/entHCA8VACAjD7RkIsy51485Y5mbedsvPwN3WWuObZV/
4skqOvqy25BlgEA9nHSjViixpUrRiEdvUUfAcYViQNaEPZyz8okaM5zUNQVPS3UMnprMrFBprmQ4
Y3zDzX2N0CkoQUw7dieTgPbZ0jCurK2APnAeudsrdwCkBaYaZ03DRxiOzgUmgFYmcoy13XiX61FW
HX1FDDmjTSpbLjRCB0oLK9IDaVaqhVy4R7ofKXoVc5EANxysiUcCMA5Lze12lWPES9D8bf/vkdMw
Qry2ghXoI8+ujDOSnq+2fUVTLFCw7qCc2/OzSLLH5UFF/T+1QkR9iTH/ugnrZhINhSXDjf1ou15M
g+0pe7HCuQpe5n652Yfa/MUxNmWVBqicYQqPCfdj0/W4zu/rBT8GLVGEC950PSE1nVToTgVffpWB
iWCVZZagjZlUvNOK+sQIOhQ9x6ZouLydxVrJiJfBIlr9FFePi/DcrZEJdtGZwd60NhIPkNVmErap
mSfjTWniZUpaG7Cahx/5HTnQnjgDwEfp27wVMC43ONqSApIhCwxxZaL1qJhDwJOS9wYcTm48ad/6
Dq+laxgc5KO0a5UKOKjHLKQ+Rm23ULC3Vu/BuTwnOYzCcfXPaTo8LipvrFgKLvaand53Ji90jjpy
o3Pvy9EVo+vwo0vv/ZRDToMgRaqD3LZ6UQ3fpwopKzz+fOWEncGO17NNMlcCyqJbCn8j5hJ0914J
fp4gkmMUTbnqQqfRRF5Hm/rRbvRpi/u+CxkzMe1/koo0T3DU/1//2302djWsYhCI7ZF4r3tKArva
3DCQzBD1/ErKhyKRMBXq6VVvaPBWp8MnCuZNYJyDj8mWTg21FgLhpDgA+cDIimH4W2lm9eqFN2Zr
3MfJdidoGu1gn5ex18LUoaTefmKpxiemhE4LU2okjpDE13xNxnU22iJYBuOlez6S2KorEMl5OyBA
8MN98VCE9ESOrSShDJ27ReEJWRioZVAgMaDZZTFbEfSc3BxLhjW81rdrs2kkGg79pCd+WLqjnw1l
tkC46dUGqBB8Uuoz1+MGYNc6CXq7kH606agc6nha+M+nsN/lV8plm99WeDm0SHSGbJKIqe7LP38h
Sbbf7HB0nYJieKGBeQmjjMhVqVj86TVidQSZca9xkNy3lCL6QMnkSRK9+odsRLQkeD2FmGKLHGzE
r/zkScswI9PTEtshQUsrA0I6zHMScxUNO3r+ajGIezPKOsb4irWq67kZKazerZVaIrHUDfChQnxv
qLThxKTDoG8afFMTCvaV7eFUtU9YXXkNL7joh48ZJG1WJCSt0mbSCjtP57M/2xPVjyCxyNV1UpDm
0cnnSUDmFKLY1sKBH+DAwiAHHXF8wVtqYX+ea0PX+LvjSZDxmHbCDiq/Y9JHpGIyV7wZdoyy3xzZ
fZW9ZU+w069J8z0NmIMCEeMnybMQVcvipFUmChkY4883EzM1j/VwVyrgAg7egsGIi1110+34GS2t
tZR/1hoMN945hAcCEsGwH+TUzanUos2VBUzEjwN2TpW5UdwY0EMgfdsUIZK2azjNq25EcORNHIY5
4mhEtmFKMl/4cmYwP7IsJzBiP+Ir8+c5Mm0n6hXGXzpZXapJ/5hqSFjlwAimckGVTjCiQr4Kjmnp
pY8UjCWDkOc+uFfic5Dy/P4hzUNFywSRUdnWaXguQOU0WY0LSivnC9gDLt2/fSVEQ2wSl0Q71VYf
B67zEtt9n99z7vpccn7W929dMz8V1zaRS4kibYh0MnSERHiqRawO2DxnMEYIvPvoF2kzN9yzvJwr
5M1GF/EEBTlKnlsO1kcx8PyzisOzqG6S4UX76IsvHt546jO5xhiiNFRmTnrimwO8X+mEwX7w4dyG
26Yg0p5Z8+lW+cY6wjOAHo0HVVCMHycC8uze8I65bnD0gcgm2AoXQn0lLJTn7LjoqOLA9mRXOz1r
sau4xcxhWTDIcyQDtkXlsjM2I2WEPIHBudrKPUiDYlthSuKzBisHyVCdjJKsRtFnwvPcR1ULRj7I
yAxCkr4aaY4SmmiNPvXNQ6fK/BOeE1PV2GrQnbs+cdo1zN2rcNxnNAPyclThJtm6QvEnEW29RTqC
YVbEywWJBXtPY7rIuoKFSyHV89DyUdf3vcHROZ1C4XUB1hc2jTCOaDOfgjCkPQ6jUmrqMj2KTIeU
on0j8XGxiAoVYYK5W+Et5lSUwKFW3DfvCH3fALPx6gV1hS1f6qiqBEug5xm3a+ZhtL/inG+c1ekR
1flFbnE/zsr2GxaSRqEyGEPh68Ax5Tj3YCTv87at0QB7wilj8WxVAnNOLcSwP4XonwpOvfRYzbIQ
lvtJq082NlL134WIJuDJnpeRPcJu96J1Oicd1fOwWYfcWpsvxeHawv8HGhB+jVxRVa2sPMjvhIVC
xLmd64d8ytW2bIJKQuEIj+1aZTcCKJaWekf4sAkAy/2t4sq30rNWaX9jrLMS+sf1BpzcqtPFGDxU
e1CjSpsWspdQfBDBbRoqvbop44Wss3qTUMDYF90ooIZPrFXNReud5OfOZPkacE/Pof8gn+sJFTpa
tr2+9/h4SEsUd8cp3NhbTqIZzp8IpmTJPWJvR+1N2/O+cvND9hwpsrpTM2DVcZrtsORyvO5FuHK4
28x8Z/XcFNpJ0EWCJwU4nYC69li6pxsR7ZcF1GJGCHcxa95qHR6gyxh1bQwPifzBIa3lolYNmrOE
L1EbZq6FFrRroWdNPaH9uTsKVR+XufG4zxyzg0JguxVKseHHyPb8X9NQdFZ+RfL56N4HNH8nIIPe
nrVxpMR6BQLGp0O4/enX2zPNksZvISt//Ye+Hj0taf7eJKLFiymaRTiaBhrDJ9orWMAIVPRF1SnD
FthO7VdhTNz3MaljOCgwpS25lUh47uw4diFdnG0AV/Xh9abV2YcAget92FgXn3GMO4BzGmua9sqo
ZDsx8RipzaYTpZwCrabTXq96W0gBZTFZDLzd8TQXs3L3ceQDzAMBPPQyqvZCrC6gg/u9ZiJiGTru
2nehymHkVArwZgdh8dvO5XMjkLnXYVF3EaL256rHChJEQwgehhBjujohuKMQf6Z3NiqeQY5DBJTz
4mXTwFofL08GswatsEuDNDq+NMYMRHK323eeuMy+40ZU23hxpwm37ITa3BaMnwQZwctQiHnc705w
ySeERSVr9T/zW4mFENM+MqA6ts3xAnHskD+MuLiesIfPk5G/cIOu2Ug8APFdnOXUqhYZ6WH0II2v
QqufyIGujdF3jTA6BAI019Hu/8RA5ZV8DffN9wjWJK6DNApf7l0VU1jv/3XyC8pg66A0CFlmZIDW
k3PWwwuKS+iGeijEQaz6SL9swB24ruSLjr6/t7ocyP1+QYbUxBsYH0F1fekDN7Tp9UnVfVRiIiBP
wkQJxmg8jhUOdHnDq3HdG0DAJsthUWVaFyqiQ2xEtuxfb567YnF0ytBcL6+DYplfdHfG+dWuP3Oe
Mj3dg6oqUc8qzHuJgeDlKjSmPE8RGHkjaYNNqnh/ZWXi+1FJu5EheWubd5P4y9vaxyBkFYSq+9Hz
Be2Y5g0LCalvZR94gtRo2Y/bILb03qgZZOQbdG1fp8kfFYRcvDS/X6PbB7wvAt0MeqBh5KnOEPbJ
+xiqMU68IiO2+DGPo1hgmmkzPZuvcapzVfIfqKog6WigVyrtUw5RBgC4A4yK+SLJzyqv0p5uJu+D
VOfs8Arp1kUA3NBtXxde0k2QXC2XatmUvu7TlqYSXbrgfC3izikZoJch7Doboj5GfTaA/rFC74Vm
WZEKcQlNTcrNq0fI5c4IeJjhdfY0pBRQN6AyhiVnFdRDsIX5qIQ+yu+uNTutCP5Z/7aA6Hxd+j6T
rQxuhaMSO2zjxhIpe3kHoJl4LTJO+e0CKcrTVIAL4hB0p9dXJKXzvnTzaGOTSsL8fnd+zQv93sqz
chHxRO/q1ikNvRO+F8RQ89m74ZE01swC4dE99gkl4JVOTTaNYdT3AQACluw8hu63qw6ViUKDHiqk
vvHQetWtqZyALrGiJjx06uXiQWOQEUUPKwTbNbUJ6A0zgm8r3UldpI5GXr+CA5fRI1N/Korvf1kk
BfvndcWWL+FNkBkVa1d5SA7dpMoLQlO+IkIGHdtB4UlC3bQu9c6whLoigciqJW0i/YNqVvxaRO26
E/kckesyJSEDnqnLKte0Gms4Ev+0S8qiYZyNXNAnWXO6BL5g2ptRHmVa4tTzAmcxJM82hOCgDYse
ryG1aFhl86MZIk2EAev7Ne4eAyxmKMTg6xcg7hqoFwSarsqfrneUx4rSH2E4IQvK6ZVG5R9oKx49
4HCR9WZXNzTmp4/i62JadycDTLq2W1YK2RbsdkNN7VHOfvvcR7szMW6z1lR+weXvc/TnlNhEtNQA
8UluyStaKlGZ668elSY4oJP73Io49DEQGtiO577TXr00AbjV6IVtC8QYDIIv/Lx/1dLjzkZerbYV
X0OB/341jvGmtNqvhy0pPupgxyMN/Ro7flogrbd+GqO73snZHANutFtW1sYZza0SCaaAZfW23rNz
WBQBz6u9QcS8cCcFDkSHdPbX78G8XTrGQGrHuG+BEZwUk3+PM8lZjLjDyYIg8w8p0BRrfNj+44OQ
sEOxuoub+1jcOoKvuklbb+d0NA3cnbTWZhj7gPMeLe2OyK1xrx9ag8UkQhFsHjKwZ1zDQ18Txwif
csEux8vkjZMb9ItFm0MYNf52Ne7qmWt+g6a7WJ42QfWIRbLUbh4+r3CdmLzDrvJ14HWXaSzDsZWU
ovGGPcJVynmCVRQ44dC5curJMLEp/wzYa2w8yvWT1q0BlHv4r5rm9jkMFZgROi3i+dgg+78nLbzX
sMu6FuTf7c2usJh+7t7Z3lEQr+um6IzQT8xo8L2pF4MAPt1/+g7P7Qji8m3pxMB0cDYQN/5zth8P
vwMzprGnzHLRz4b4HXV5mHJX9m0jTGmW4arvjXVOj/VazRwACaroMozqwqyPFqPAPB35XEzwUKWP
Y70DrXB02kXGGOCUsMLQ3tysWTEgLDjyqZec5KzEFPn2Opkt+fkprg5MIljqVfpDWrNoY4gM21UA
HvsDpo93L69/LwQPx/lrv+Nr0HZr5RjX8uBcPsZit3rN7i712NnenVIVZ9xxR1+ipBe/nyvitAME
BIuL6oeiWbD40mVfAi7RjjjQ3qZvOHjdYm5vhfNgJZx8AKKg9Yt0PMElNi3oIT49h0pL7Q+ThkAw
opKdL8Go1hCDkYx+yzLYxoAY7RofwabFdkJCdt3NrDLDFhVNXRE/btIx3HCKweL4f3DTbrd2fzzu
9hBaIi94HgCc4iZONxgijZ2k9oi9E1uTF3Uuk8PIeWCpz4gX3JY/2S6GlyR4/Y+KWHlSUd3H/6CY
/DO7RNUzLVsGJqKUHpNQNEutiKsf7FC8ATV4JaxdvzZXaxSondsz0qgCWdOWlDCx/QxUZxHrFeZe
eT9g7/a0/B8fnvymSb85xw9Bej1LqR4z30UqXA8jzixfkF3cewDhcGyDjntLHZ5ZJ4dn653BSoZu
H4qIOIKeRX7SDIJr6xUs/35K2i7qI7lLNDprpmg2OpFmm+MeApfb5kvTSfNmVgWJ0Gl+pcX9B5kq
PYExvsqnUsiEGsLJC9YnmmOYdbtrnWSAITCvXCCAQzXx74oom1ZHh7AMc/ceP4cKr2XZBaZYFT8L
t0ON8k+P0L7FI6Vo3HrJuwa/wA9JcZL4lbCT4Gl4XtHCSS+kcv7qvnfTgB++qHcd+h6wQp7JhP8D
HcQPqyIVQ8aSwKp8b+ZniXwNQZAZ3U3uEeBhekPMw59H+Xo+bcbiPpHDX3/LGRgW541ONNb6go9Q
/6jor+uo9ZkVinpBFxKMupD1SRkYo0fvuPOarOwGSME82/TKbS4Dv49SV6lhfphZDNVsrPvZ3MDZ
H4zaVPSR8cD4JLADmc0oNkWSIJ+fabwMXf9qW3kzqfjfhyJIb1PLEkLXpd3Ehhb00lMSYN9k0+9n
0K2Hf8duKOp2lTfPRShTdUigbtDUL5J7eJC8KQpJesOMko6q7Gmi5VIadihXIRLNZtC7c74sOGXy
ye2Dakq0YyiLA+qa7wswNAJy+IOnZfQpTqald/eK95PU+TdmpkpWxwYyhepbsNcS7SGcvQRA9Jb2
g1XGlMz/ddDpNbH4snBTrH7vGQuvxixfi91JQLrs82wW+aktEwAp4E7z06YUepvikPqb32j122q7
r/22lBlU5vg+rhCCRARjaVZGH+uv2o2h4JdEPVHwtPOudE5G+blMfowZd2ODC+V8kGgaIDCna34Z
I4U+NZqkKzRpShslZVtMVHa13DG3XRYCeEhnciX28xJyuz4fJ1Ym7B6HSvWOXPKG1ymQ7YXrH04f
t6VI85riG/tgAc7TXQFJ1NRbVYWnMhDGLPaXHmj1U8AxvCfXFaUuV9hcfcRntWet1tCq6Kj9zI1b
eE3G0CvHBi7autujVq5dJxE2tX/AqCDBX7KKK07AnZz+7WhYI1BvEn7Bfdcyr+R9+4QFyCG2RoRV
c5jhIzMf2rixN16tSHFRv4KvpxCJtF2mgcOCvTxm89D6kJhJcHlc7syCqP/NvuFFANp1vn0hm9Sw
o4aKEJBL77abJvlZvp8F7tYjphadkq0HLQR9OuLl6xKXDMHUOxisnHDaY81E7QKw9jWRP/Mr50oi
tRpJ9iTHQ2+kNDoGs+i6CO8icLGml3jekMLEeHykTW7kZMPvGE7wHRe+uXtev+nnHULaQG0zHMhv
USql9lrxj6TiUBbrz8B4HLGSE1S/Qvowga+nRR9QG68XhfkWH0mjZjTMJTGrrub6Czm3KBrGoeHT
1ildEHfUMe7bTM/9Th7DEhw4f4Y6qyQZcnNF/wFimTZslfZNwv5vN4vboS9zyNrpxN7YwWDoQF5X
fjqJvzhGY7rOOsJS8jKUXF54iyQvlXMNUGIx/RDdG25owWHNFiFqpL/ra7QtxhfSaOMfHseVXPbj
dQzW7h/7hV8l5ZFTTpYb86CZ0rouqnxak+0kupgnQHQrUGo0Fm59plaDhshlhb92Qed8Xw0jASqT
sNqX6+OXILNnil2Qjh3Gtl+hB6Wil/UK2CpcCeyS2GLuZJttFrGaxcHi27AwHoJBSFxcEKgCrFro
UFOKNmDd28giQbYfkEigboeaZTFGlhMX8uKjsn2ntLbpxcnaJmux1oQt1qNBYYmxfp515ZWb5WzC
d7B6pqawDXF+83a+GH1zMbyly9Sx4THLopto4tv9H9yGjG7iG+FwSNgRtAXFeDCyJ98wjWs316N6
dZpSAi9t32bj/J084iVwnI/isCKqtGsuYizFo8SUOn6/WhW2M/gVoRxxcb16bbcPqX7J/VFawjbz
j0TVLKQOG42h/y8pTxnh9qNHe91/f5lSdYIUtQ1UIDpTLE3I9zLijak7zWvjpA8n8gahjTHMHQ3K
dQ6iv1LLE7xxdBvcLkYKCicPfggD4kPf16X5SSztoWMhJxHjxtOzYazeLlZaZC2xESYEglnidS49
q4bNfM0L/zPzv8yV1Ks2IBohr3CZFf6IIgyF/wX5JXdNTAwk99wH7pJStKOE8fYFjHG3EpAgbe2c
ozfM0gsQcXSoKV0aT24euOb09uA5UucZRHZtvkt9HXjQvWHfLao/pAmrluwHKqgcF4dcgoZS76ag
iIxCEhj2TMUyCXW+S33WHCxaEiIf+SDOm2Cmc0dumsI8kMSzKdS5se4+nydZwjA4rgE6M263NjwJ
kcNsIP9R+gsX4Ie8yTckzfm4/Lhosi1c0+HC8OTK6cAZfg6zYn9KPqhlP4/Iulk1mUPJIkwEhqqB
Pp4FJyfbto+WAm3Os+WhkmoV6Szwbt2KbvB857HALQvphCqUAzCPfBViZspBttFkcd6xeo2PIuR8
XN74ktiYCXbQZQEZBoY8M0IsjagdPEyoNu+PbbqUMgv73hP1y6iZ120fcoMhO4vwFopf2KL/cbjC
6RHgcV1TLIVkupk9Z/l7yrP/D1VP9aHh6gczCCt7pBHD/ULL/Y20lOzXgJEABvQPTru0uLj/Tstx
E5ZuUFqadtqQeCqzxfZfJNif5cj4vKkCwqvFJPEkdNQShNX5NVTher1nKmZS6teFcDk+PBkpjCwx
ECn5zapmI5z5dHXrnMUQ6umhhqzffNR37LBNXFn3/p34qNbl6qqnOVZweE9KuQ8NwI+b5adXFNZx
t91DiOPAbUiGXEHqARTFobhXPHki6ESlG/IttR5Z32KrLpbU7IKYfaRGGZWN2nvKmALY8cb4R/lY
aszh+aOgYoK5cgJT9jthXmIkbLmgwvYozAsD0rr5YNBVM4/S5m7xQQXoOyzl8cc2TOe8wC7SfZaL
XSdpDr3iTbeOIagGqES1fFzKUbvX2pI3pf2mEyq5iDlWpaC03/VW/NCj6gxBEH07FHaO1r9p8WoB
ofgVQo5Q+ZNzCtQL1qWVQ3R1agBlQK/TEopGOv/CiFARzO9ipqLKIKHjmm9TGJmNN8edEhJtX5BD
KJWkZRnDBTkV5HMNk90Rzc90IEZI9I8ij6JaTsRPtSvDIty15FlqHqTT7y0K45H0v8ZyGuspmsiF
BJOxw34B348zf5F7i7S9O6pSpPULZLqClh9GEHhqtIxSG1ZR/gObwEcGDN0WyHzDX2BhdAsDIUni
d/npA/tMqcPHiGfxOlXjiR/OaebIdKmQ8U5tyJevmcCqtXBFtHd5/0QHOvTif/McR3JYR+/zQZT3
61TLqzDqaS+aqURs3C0d2y2+XbwnZvAZMrDGzLp23Dd3aimyb4KwLF4Fn9BOgcte/yYK4kTkqyAu
N78NsXmmP9sne0nRqVMmMfEwLTayqA/rA4GVthi+HfBSpJtRJXjQz3cjGbG+y8st/tQ7G6QztUCm
EMrG3U2Wpw0IEeoJyawdbNiMQByYJwKtimqvYJQITzGAypr4I5Bxxsb0zfDCI+D6x/QeS87s4FW4
LhK338a4k4wlVwkUcMiCGCagaw4ITycExevLDau/ffLibrwVNEb3ncNUeYp4srCuR3U9bH/8LrfC
k3UpXPAV+SBgb7eFskrqDUdlElBQoxiABUjNeiAMvAoKnEuSXR3ghj/7/BZgQrGkOhchdJ9Tovu+
loRtat99QtfeZQkOSj/zbrTk1N+jTF8E8uk1wni5t5zXN/i+Iqi9dPiOTK/DiV/Uk7shTin5UQzZ
vSZqwKYfRfb2RuxNLhP+h47g/cAQnNtfqvGhRuyKlwCMv5QlwpC3ltyuA1LZFo0VQnyG+9Y5t8o8
KHbZv1ZeqRukmB7Xzf4acgaB4C9yKll1vR3ppnLStu/Zwl7tDWi3XeBbU7hWRimmTGkVOlZxsmv0
5OSOWuxnhR2rTwTtpvEYFBKPP/L7lB6QiKYYOEwD0H255Kz1Jxk5ZK9nkehJwgJyC4GgvrzP5bbV
RRQDwjxbQqQNtU3beFH6GxIFnzNQKBxuEvjbWQpcZrG//iJQKvgDdcMNSjzYAy38oDs20HGK+CNJ
7RUGVvCz1Hs04r1oUY+OlXoBN2KgotQHx92hMnYVNjExEQzfNZKJY+M7iSHC+c3/+ABMlkCd92oA
nndY3YUYhumHmJxt7XQ80HteSH/lv8DMdP3BYkNkqABgar6X6kJ5L1a/PSJK7ELg4ydVRHWc0ztJ
zUYFclotLNivQ9LAozD8+r+x6r2vv9s5Hcrv4F5hG1elrT63XlL+88yA2fSWrXpE0/8pbeFWRoOo
oUS0PAspGVnaveuVAp5QAINnihhzJaVWZjsLEejW4BiCsheP/Xpadb0oDqMipfWMtBx7ABqR+GzC
FVcNzjmVUe536rv3M+X9nqqQWEu1eqjLjlgajCIrfnUn6LfbHHnCzHyFtL3or/0KWznsueBg3BBn
hOjp/klhGCS5GiGytn+6jyg5f5+EHN/yeB4AA15DlaA8mWuWVT3DjxLzf8daVsxgCZIXFum6QTgF
c/A5XDui7g6H1ptkJ59sKu5UeaX1H4x94OfDkj1E6M6cnlEXOTk3S13E8/rH5MhNDw17/ZckUO+2
cOgWtfIHNO6NLp+Tyyf0uzAeTjFjWZjlzBKxI9LjUfvQgNN2NWSLsne0oz9kBTv8feA7NAcu38wv
JspCV3TyWA8orDXaAaRIwJ1W/cLvqIqgPT2rHQKJuu2eCJdZGWxUur9owo1sT+Rpjp18pH0GSfzE
NsWQwc9hrruftZV6cOwouRNZNohhJpIkQAnQmRHU3E2Tqg8YawhKtb0QYkhXSMzJJV6IM0Zk+Sq0
XaztvwYife+2YM3m0iI5uqWaN4ltDg/F6SoryAcfpa5wTPMlrz8yve5x3iyzm7Y7lyBSVsVsGnYY
3Ecu7qQNgq03xPHa3kn2FRT2Coe2flN8607BMAJAFAOasQuDRbP7IyhPiy3FYE0RUOjGO0bgYf9L
AdeKt5fmHcmwttz3q+xWmgH5SSoKAMkPqnWj8+gD/5zleMSOzylMr0z+0O1tDloCwuH50jqgzt/p
BPpjy1q0OghSScWokt3nCl/xLjwdPsmeDAKBBbZxbh1kjOfihb18kcbMWdVOc4+20yqVci2jprg1
yN1ux6W8ZbpOv5wIf7KlYtY/YrmQ7H70/XGBcZcRa0NrIQtIHfFmdobvj5/S341bNc+Zb8KRj+O3
Y7NJbnM3Gks8rOlMHrMnn/k3mDE6v6Z2Tt+7ilqdZ3TZAQStv5FAQDT3EPF7s+7ySo1iacMNM0uk
MxRyoZRLatFQ8NNz4p+6z80U8fJq8oGwOP6PDLq5sFWyW8Bdd7i/m1s09CzUHj6E/669kOJq19hn
Sj70Fs1xj1Yn3Vj7OVrBO27gH7tX1Uqa4V4GjlZV4ESI0qU+L1sqbq0AkAjKgcepHOc/Q0+50fcf
jSNoVGMCS/4mc8X7r9yVNjmkVmR7dK/fK/iXwhhhHIJ8g4RyXwC2sE0U/OaSGtf7MnxRhJJRegok
cDttYxucQTvF/eG7fMhcPrtbifpMCM7FOOzK86mORkTsP3RtNNXslEeQoECjAlAY/z1G9F5b0Dqu
5OxyaDGUw3C2ijSwBdR1BNeYtXzGdKviweMBqAA4BuPGvVf5e26HEFT+WrFrdaStkLLFSUbJQ+c1
rvQMRYZaXL+o2SWEy7AE2P/U5GAWiIiuD5FmZIEWESQR/Zdj2x3az7aDE+520Xf8lKnde0zwSUZC
9YnB6J4JCtisaICPHFGlfOCq1pXBJZSTu60uRicLMMrCrspjW4QymVQ1+lAwnO7LpqFhLC9Xvj/5
nM6eqGInO8yGckPtAT5n5X5PfgwBd4D+I2xA2xN+Z5GOvm6xVr5rH6fj/F2UcQXs3zxHj95ac4ZE
whsEgQ/macqwGunOuQKg4Wv6ONlR/VVioHdM4Egwb1Bcb7tycIT8pr4qsCRbF1faxbGWkXlhYl5v
jvJoorzTqx/mEvpM7Oi7kRWs2tjpfWkeMxMKzHDllgIKH6LtikmoAIIbsGINm8coxxb+0hPrnoX0
dsk4lpgEZarXoRaFw21vmhJv6nuAGhvBEP7yh/Lx2xRpOK3vve+BS7qRce2EJX0Be77UlGZfNUjT
9Y+lKohPA23DiVsidrsZgTrz+bYEvUCeoBqb4UnOPNArM0YVDQOyupTLkNg2jna8pwUfPjuomtM0
zIn68qRU23+3Tt5nIGD5Bn2/urM+0SDOI1ROQhCm6bhnds0Rzy63bNGn7FaBvcH5VbYQP3k7GaON
z39ptwTmoGaLKUZGozn5cTJIckMp5mFKVWCG7Gqjk+0fdw4J7ELohByzgb8f/isJ9WneBLWEhCRx
ale0/yGTjHAU8R7pY/t6thxjUqWD0uZXJyCrLvnJey7lfxrqyLWLkfVJDyzoqqogYsLXqb9kEz+p
3jKWnzDyXJwV0lvti4DGa1hszeLzldvOfOhxbyckBnzusGOfcSgVVN3pHCFTplf1N3t8rRLCrwtT
o4r5c9hfbCI2XX5iwuhClW4AN8SOgd9NOtuM1YjaM7/DqIV/qRfJ/Q45MY7Iff4OOBEkJudpIAvk
AV0EGNVBGB6Ksn9Yoj7M8Lc1axWVRQhdEQmxYXvqLk6252zuoe3rxB+sOyoZoq7P+m9Ls9+ozj0S
W+W2sl3Pk704N0wZ4ZbIfT41sJiKeoFa6FPmcuemTCKSTBlXsLJpSFMlV8D5iYbEmNpKod6U9Qd8
QhfXkrjDPOZHCwLmKb3rjbmoLOq89ASGcOH8b7vJ2kr+4wzDLzAKt/y3Q4sSsJpYKXp0OQ44+sHE
QK5tGpIFMp0L56/QTBpo48Y0AGBnmyOR2QbKgUuQXvJpS8ToqEcH5g0eDcDThP9OK+Frkh1u4w8g
WjqO/Rdu9Z+Nk793dSavuYtWmLwEKxnGCnaDETlwEbcqr49o2sxsS/vJTQWfDw0VmgIEbQBSXWCW
oo7CY+tKEe2C0J9yDH9BXrEUFXGLNhpRajfKgk8pRXSZW0vFWIQ1dyqxHq48mhYS3Xz7EUnNBMiX
gF9L0y1FumKKAA7RmFuHspHdA34u8KvgZiSQ9KOQ7WJIRiuwPaC8wAgL3/HKRsJjNY4rHORlP7h/
rtqobT5p2FVpIp1bAum+/RvcbbkfxUE5Lkp8hNALQVPuV9BRPHNUHiu/muSaCIqm+iy0aWGkAjdk
2bZGi4R7J8YmVTblYI8gTgk+G4ieD3T+fwOVczAaXS2zuM5Mzpx21dwOdOe5s8VqXLUfdhuPsxmW
8dAPbttUp3zV5NKN88ceMt9yjwISLbm/SlaRYgaO6CD5JE2R+aDSvn7ztEiOYoT4+dlQ5tSO6CuG
3quRZEpRoRvAYtErpsGuOhYByyjTuH12zY1ZnUnCEWQmgLshMxe4yOCzFKn+Ot9QQCMZVjpUAYkK
QEFVAQwYrycGQysBjSvdwuLSXAbYgK03CvYcKQvkZC5JaA+xd9ab7TYEJ5loWC+W3PpfuN7n0vTU
fKL9U1JFry3+KaApOSO88lBYroJqvVDLJIS4lKGIfTWipyXgTRfS02hBZFEW+cnFZE+mMAlrtsrB
Kg4Esb6dJdkwuxh1DFMwKBCvDQeejc7BmH3IKP62ubQ+aIItseuNjFb2KZikC2JOIe3O4cpaDxuF
/158fhZl6izvZAh2kKLcfbKyju9ZuXhKWP8XUQqN0dkWwPGie2DAftd9Wdjvl+waZzaeZ0Fk0+ye
ELSpnvpXXoPrjP8SlB2JcmVvFZxfbRiMOOgXtm8eJL8u2Hdz0/XBFq8sJeuzk8rJ55GymrozrvLx
8DMj1Bo7A9vPxqHO+F3yTkFv/oRzLIB3h1QbmwVJmQXWAnjPPdiAqsn3RshfbZ2vOR1ay48Vxg6T
dq43e69Zu//jS+H2MmhGkg8grpCZFVXIQiGmYsEZ6c1gdUw15H0WNvvephAOBzdltyr2KOU6Ooan
72dmT8IRSCkWAmXNlCbk2TCfktbkldqoElpIMyHuWJzJBGUwfR75lmr+dRl6fyVWATfg7yCp39ju
sAGKBdhRqQs50NZpMfc8AxszgVu3C5WSBYtBjkKdT+vZz0gF9VV8gbME41KQ206GSLNMJljtqhGM
iyhLEUnHJhrbAWwq0DREEy1nFnGw3PArp2zDrCj6AbAvJDcj5RXB6sCSJEhmsONJIQslWGfoTQ7J
04J2ukoXFbekZ1JWdYYi8Oysml7uRtacaIuxwoFbIY9N+rgEUuIslfw6GWzskx1Y/2VY2+fop61v
A61FHM9pVOztud7XmsIyigB8i4hw+B0Q2Vrv7gAS+wnor5SFF+7zV8dRfGLqCO321BKlacjh2zAZ
HkMxb45F93oESYlIMN5NntCDky4a45e3eeS+ArO73enwKnPRRB6fukm41/wY04NBWi2uqoM6fdnP
b0Vh5sBabArf0NJAi6OGq83wAc3liLdtgc2g/Msm2EsaiQhWd06+VkUjGMSU86F177+vfclRiAEe
3eDSXYjhnnljgTLIdSaGOUkZc02++SmdJYaWDzHK1WRnM6ylDBod97bh6t2sZndNd10a9aze0umX
2gn73Un7dltTJ/pL1azzcxCffm+6Zj939WcNvsfyYmJbQufKH0ipcfg6WZY7s8hBKlEGTkz8Dkpt
tMeDhLj8ub/3+TSKSuCHS+66fYYO0qodFAxiBoi2Csv10x1gR5O2ZHtA5L0DbGH9TYXU0acHPIaJ
hECklW/rYBITECBUMfcki4hz/IGPzd405907oRwPHSOEgyeBBhuwcOORsoeeid+upmrUt6rWwrre
1Mz4cb7wr5sabss4Qm/IDLK4keRz7P++C7uERazsEjgFA4R4Rpe80jPGYOWCAK7ywHSpfSHsihqC
20MaoD95QqatB6htZ/WlkBoCdvwdhaVqEcJOSpLZXtNXPssqrGXrZTRIj3aYXNwWP8VwLgqADBhb
m6j+Bt0n3vSJRSQPiIcguI2YDJj+3usNsfpw/qOdxsJbCR5wyrWCc1hWtn9TwcKt5mzKnHqZCSDU
Wtss10E2fTYJn3tgt2GizWi0Q7kg8mkWBB9eCkbxat5IIZpDR8BQiDlL9na3mf7Ohpc/nYyeO/a3
IfxAEau1bSnIGrhbhEowhZs8pMKMRQf0GChAkmooH5J5VJt9agGVYdxxUM9R4i38mDG4cpAGSy1G
HO7AvNKnJKwWYta9qbqNubpwErSEwzPAPDJABYq2zSuXLRU+ZPgTpbTORyStbY1VwIbjxqphSpd+
1UPQgJU0HAXkHx2ozCmBjsW7YAozWfZaxrAIjYCpimSS7otDZhAFj0apwssotrZovuqhOTyA/j7K
fM4RerGG6DiHDBNsC4B7d6tKGo3/C4csG7ycuIxaTGGd/SsxU+3PeaZRuStzcONSxffAHxn4GjA2
eAoPftP87lQ+mjOZJ4FC8KYCxN5PeU4T8qJ6Q65B2y+eQi2cHlfuyG1tBbUh1V7Pf3TUe9nL9BB3
IMCk+8tn+FFJz1Ci3TOmqKoJD0r/jIVD7lrIkET9zZCHV7jaK32VDePhhQ/yHZ38saCGp7cnSTEI
Lj7A7x5Wiea1prxDrH/VasCgDSDCEHIG/5JsnolMF9nTmj70ef5cj00n0stMPi8UIiYU1og68fv2
6C8gYiPiM723UHkIR4TbR8h5f2ld4T6LNsMpbyhoxlaRMQFinrUPJO/7+4iCLRYcT7zC6Oyj5PKt
7kaLJV8ug/rXmdk84uMJ/6w6vYZfEuBuB85VrT29muknpDcGaHazejC34KTXtOvj3aD94qooSytC
akIlMLAUKId9z1Q2kWpNPVOiqLVFB3R1Wyg707s5JFdunOrlKYV/HL+g60v5RvLIzZhI6qyEg+6K
lGgXdFUzwyDNsxdH1IfCsvyr/9PZZDW/wdcer24qByzwNshly4FNTnnGZ5ronWF/iygyZXFyROVa
UiL2NFOWAI6PGb2vaGlZM5NCMIPP27Rku9sBf3Ssk+GNFGKAy5rqnPl6o6qSvi9Qw5uPTBtE8JLQ
midFGQ8LEBoqsNFqdjRKgM22haZ8IQc4OMvb+mKAFCjVdBO+1UYxR1X8rYmTQ9zZb10WNxA4zPgx
zVE0LQPdR0Hdqro8+WXel8+cPaYr6W/ObRN2eCfgclD0/ibOXMAfxODYr8M1/eSxalOUt5tOL/tY
9hRNslzL2hKZ8ahPrbQlDOSX5HGCP29LZ2iQtJ8A11iy4rpZBfoSkpLljLcJ5+cZEcTzAKqBsSPi
oKPlSj52KHD9xZwgnP4Z1eGE2lNdf+Y6BG8UCLR8dAK52PoHeegVMI6ZoYKlEAVlYyeAklZImJeS
5yhMI5hWzVUumTGy0Pi6DQZmq9gERAvd1AnzUU/qiLRjWruWh2ad7vFyDEFuRnY5sV6ZXfmmcDdC
6L7K0D7NwrEw32Blyrrk5Ah9HXvNs683LomIgNYsVxHeTxfeinL1X1KegpXUZdc+1xlQlwz/XRuO
MSoX7KW6H3irj6mYzwcAYmvnHY3kxFixv+l1fORbFRNDX+n8Mp9k2xavn5vGBMLtEKPIjcwFx2CX
EHzHbyGRgSPGz3D/bCZISQ2vgxYoJ6cyS9yDpSm6FanItwa+EagjrmuKFRth2YiJUg3X1OPEv2yr
4c7Jo7igNREcN7aVm+2WpP1Z1AGmjYF+r8uk8wiD/KqAdf0aF631hubqGm+l9qHbqKz5Znf/k1Fn
DWs6JrIAlBYBu4faZm0FzGARE23fHW1pvRdGVlViCERGwWbcMuheQl/mbGvLDupP8A5qnEnjm349
yOGOpx9A5Btta3tBKqxO7ze4mEKbeeH1ibrQzsf9bGXUbfwA5uf++QIRpA+X7lpKkw2GkyKj/F79
DfYHhzOCrkd/q8g7r8PontSWP2mk7TmXAEtgEf5DP6qoo9sg5q6ip2sSiBBN3CiLaSSaAosJ666A
X+ruvmP/1WOXGBDXEFC9ovBzZ7UzHqjuy/b75cL6toPbYuniklrzflqSVI2rsBRaXg5/rbfwOV5p
R+iHKHHD3HjghlIxoEoKZCfJ3oFo1HhDNY29FVIIn+N5bI8hyGimvnG5Xq/2hlCob5MURrq18oKt
140T044L91yDpjOKR7VcODob1rLqCGKf79tSXCctg5ODZ77/2O0sPuN2c/nO7Z1LAxg+RsIg0E7+
CUzIXMcZxxinsOHsoLiJcK1/psuoKvkuC/GFhyjjp8K60l/3UwAf1xTh1cVR8If9maSURFWKRkOd
stuVne6AWBtfdQep61O4a7VXo0evrh5TNbktMD1YMLw4f1XJq+ST11y6R1LjaGPvn8MF8Ix0vpnB
6i1heHv97s2Xwwky2HRosWJxHr7qVMZMiJtzqqCJ86r65nNEpreH0goP7o1Rqqp0YWZ78gTnkghX
xvJENPyLrg2iJGZB1RFfylm+dhNMjBNV1Rg786jOP0DCu+tMo4eZaLAzV74zoj/3vvXZZXDZ5F37
DPZQWH5pIYoKRuzrtu5z8Qf9msw/dl+49od0ms2wTHEZTid8mF0M3r4RCzw4GeaG3Yb0KFf8Niue
om7WmhXRKI8ea3s77rEUoWaaJfbBWRkslPVCNqdN0IarZE7RRTiptNXPfbfuD9WdxiAJMvG2pj2V
n/EOe9bWNM2kXeILWRZzDXk9HqTwUHZgHAM1ad7QcvEsIhwJWGKh6hUXWQA3ztNoRcvSUIwoeJyC
gMUxtNkYGSDf8eqyfHUR+GH7R2dfoYJtGlhx/8gU876jJsP9IXbahjJMeCYbyW8bz1q6UgjJdYQK
CI8ur1yFyqSRtqf4Vnli94usYEWR7pPcRgMQgoGMoa7B1TtXqcgUl8Hb4ZIOq/4H9RdBmIS5+9rQ
kEAs+0tRgg4iX6zN+OGJb+GrtSmXHzBaz5Pb83UdFsgCeryYBZzeTnMAqZmzogTrRJkxr0baRAgw
sUclkkxXh0Fhx5Jk1nbxY7BGo5kkWdee6ZzMHV5H7yqeH9IMXqk1hf8qLe0Nwp2i1UEE8MMk5IJW
OCEc77q/9LQz70qxtVsorLdKCvEOxphmFb+gdTkz9DcS9MEgKxQH739K5zhzAyGCzBStuA3s3APn
lASkZ6TFL2K5Cfprg7EYNk8RoVZKPw+h5Sje4SaD+Hww2Yjt+/wBq6V3Hecn2NNtf8lqf6n5RbiX
AzGtIeuB/5sJNWXzvWN0h/dfIw/GB+I45LmMVbuzglqlepSptle3BWyR/ajGkmZQC9+Cy56Zi+Gf
LIMsXGXr2BYQtz6JrNOYVp/S2eFctm9VosxF9ezT3QQ7oyYwaV+weiaM7EXumDT4X27J6SEAsYQI
Tv+mg1SVIc/2HegFyXunbbuz0+yF9k1sF2+fjoq623hYdGpXNyrjE2eITgwhbnGOCisL18oHACeF
3aHP+Il2xiujsh/wkISQR2JqntJCYbJrIoGjj0zAqRuhyVnvMrr1l4gCpIaPyVOjE047tCKtE4Q/
rzHXWmC4nHV3oSSF8zojSpnCBi1RAkFtEV4kcsIzTkjwYzBSwN3pmHMgSH2GhACmxsGzkGgoHcj1
xqLseFSJjyeArqFxc+/GbrmUT85GDLAwyNiuaRhfLhtYebvacxKWqFUmOiDxfzf8nRWcfPRMO+to
mQsQUmYTMf6wAj7KJLEV/tsPg0hmDGqgytP0N+n176kP8zQ18n87ZCp0Ew0B/0GD5g81Cip52WlZ
Y6BhV/ZG7DsIjMhgdcwNLTMbDjMjCQUBXVfymZM2y3mZx4tY1JFtb47buxSWjgMI8BfMscxERRwT
zgcfjkPZBWNhFp+IaA/GnV7b+Hx56K5dEaEWiBkSfjkp4Ghaf39F6skmb0uVD727f0r0LjZRMGTu
EQDOhGUUTbcy4YXRNPDaPOadsAb776iVd7yK5irZG44pOCvXh+zvpaBybx7WpKWMOBjozW/EQzIG
PG2/I6qn0r//eRe7ltFvXhEYUxLu8VskQ0Q4GO5nJi0hNQwUS0DEKVS1JM0SI+R9I7+EJB3GuF1A
UbbHYhXlDLDxs8W8Em4jhEwf99BE6gE1mi3kJ4uth5CBEx+9vt9MPuYqHh54eWDK205s15zbLIkb
+jOMQTfens6w759PZJPI4+XB1YzQkU2tbd+9bv8NiMa3zkt/t1HMIpRHXfg1ojsSlUt6+k8aXkbI
wmc/1Loy/BBCIAqCwdBNPHfKJDBDwJktlntqB8Cajwig/x1PnTcGXScCHPvDTrJ7ez9WZt8/TfMp
J3D8s3FFzrgfRYvpG6FmnPkU6rpbYsWV4N53u9oKYfnIA33nHKvW7TJ/ezEc/wgOoypPPJJQClXI
ikPM/wfeVmOliCNb0wYbl7GCIVbAhbdz129QEbbHxn6HWGiFUuz6Q/IgSBss5WYZOgoGgNicKnLX
jCpWPaa5KyIZAlLn1wnNeXwu9Wl9TgPVV6mhSqEqushYoYy/VIpWIiSUt8QwxjCbovnmzRx4ea1a
k0V0Rh3CZIvzC1anpYZ+ccwKiYQDBTCmavneROA+foT/02Z2tgEbT33RJx/H7jGfHID/gJat3vt6
ZHWQeMEQ8XRqPkucCangh8I0qGpVFQbzrMxJ7uQRcf+/Gq4x0zmmAgJ/EaBSaml4AJ5TMGG3rgBs
2s/s5qqCp3zx7kqzv6fSfDMeHzf0zY6tF7pDZB1nogkSsep4FsVkYSWR8TV2zXb0nNwdMbb1+NWz
ctsdmxjX05cDo0mG5tG57smL5qgAYuCfCgB8PlqriC6cGalK/swYvi+22rUabI5W4+JHbkfgBdBZ
uoYM5Tt6S6LnqVDoXpmnECSmvu7hQj6LOVYcujCEcceLjE27kaAiRClN25rc+adWtCUs9JIHFqZz
xM/HveNizXVa71h2StfVUOlTeq87qalxh1+QYq+ywjJhxkJBgQSIYKDQ6zMRyXwg+Nkpw1lMhc7a
AcSWFcf73UAPrT3CzU+HsqIX0kmxNDAw+t0Qh5PcoimMbvfhmAVJQKm/Nlz8ygXhtdONgb7k3Jpr
uzFgsQYIPZAwIlrArmI3WBEryhMhhT4viRwhBeWKDQW2SML/hJPG7F9x65hMe8Vu1WVUrDy80tAi
kK50pXdO26tS8jUG76OtpqCuKKxaG1Sha2pwzKLfiQhT8sSW5rnDuifhAepYSXEzkPxfat/2gmB6
Rq8xjAfgyl7oBDxhApEyje1Chjb8wq0pw7D3Ru3I8ipOfsxf1eMnCuO4LstdD2MtFFKq52q0Wtfy
peiYcnLfDsjnlS8f2G+hRSKAVSUgCSINltoX2KA0hLDNRXPUec82a48J2qAnV3NIUiD4pBCPyma0
7h7n2XbvqxFCWzT40FtWpi5DOzlQOCFff6Dh6/DUGwRj5pOzgaVBYoNRGUo/gCKZXZgrlXqh7RXw
WUhP6N+2Y11yIFX40//XiaL+1ISieJSNVjyYfpAW691Rzi1BPzIkeZwkzMrX2NG/XVmyMSkGk64W
9alS2M+tIbAkBAJnuWqNwUnGmcBXM1RdzD2frChN5xk+YNasQtBIpUx62CHJALAqCrCmbWxEbNbr
y6o7AzIHwgkb0up/Ltjq7iFbmcaI+oDwn9GPq1OLWLqk2C/2Tk/R1xmkzFxjdMhaNJ0Zw2ADmrVl
FbIA2MKNDHoP2p9yid6MBpbQ0+COrztngF/tY7WyhNCEs99LJEza7A3O84bLsi2NAvG1e37Jyuvm
Y1u4XJesLvcsZZrPXog5OrCHg0p6jzUOXkT1XTCXRHyeu75RvDqb2y9thI8lcrSvqv6yIF+CPB8z
6GxcK8dQ/PjaKnNxqGLZTSgAGSWV9A7eyjCv8fdAR/WuERNw+6xTWpGjhqxQkxTl18O8h2EF/lWc
h0gJNnavIbKT2vlR0I0Ip4XLJNAXkghB6nw5tZhk5WwnDUVAO8oG4jJnpTRz1Pr+P4u3GU18OvWH
aCHABgspAFAvVXXhvxajoMwutOgulwbZnw7k0V6fCSttx5Wh4s3tdZ9Mh3eUBBh6sOlQ3be+bFdF
6vb8LyR9ci/KPioQX4ah/d6JddQaqtukIAZDMADpxpBueacv25LXhKLaCPVmEonpV7R7j7bpYs8g
ouAdcZWiGfFjlGRdlxO922nvv8JSMlFPqnSvr7zphLGAT1q0KWfIRgJ8JSMci654QymMLHAoUn0i
SUNThDD2N1wpy1wYPg3KNOAngFyiK5SogGayAkmOv+1VRfFhz8UBu4KV6poYrHT/cVX7IUcp4TKu
6BRVWs1qaXv1cdeRpQxDqFJOm+XavzldHL8rfIVMlfDiPbgCIHkkUulRt93H6p8z+5IvBXcUG7zm
87o3xQxRsWxdxfe3g2DLLMkQ140YPWlHHCwfxadvQE1bTmhVMWxwOWpwuXtHz51/XjTAdak7K3Nh
C1kcz+5N+87NbvrQHP0RxxoTREdPiFvdXFACPvJ6vI83NhrcLOhHD7CZdzfLAaV2+Up/DKRiQXLS
gkbjyJpQa5387t97ldbiJd7YRUmV75BbK3NIG3hILARKcGMKQmW++rRaSOYaiD5MzRoA5tJO9Lfe
rfE6tWgH5rS55UphyGB1aA8xJOvwX2nmHzJZaxX6/agPXO8sTqC0D2ceycwg5ktxyNsmqCgCaizQ
REV0gKYvnLKKeNIsKbSwBlOL0ieL16P9HzQPmt03+XPXWTUjQPLUCb3sLaOvNB3AvC75pzqzyae2
lA9vjGbu3V2FPWgpS8nat9yoKMoEwb/NTAowpRpHiI2vrPt8v5hY9drG5gNB7bhqSgsEcdItfvk/
KpMHgXj97oQRHMRpUK33PI/DnlxIpnCqnfxMYSg4+dJnXbyD02xT+DhlZdErrAC4OAKTDUTP1x+D
NFFMefHtsjwmKVPNj1b1qF32edBGR23ngKmSwPpUwDgNA/pxxSqYIJYGZQILp/90q/Yo4FA0F+MG
sMvHugybH0tefoJvw7dkbGXvubI2EV5neFsoA9aW9ObZEXF3M4uwl5Oom2EbQhOduL+BhVLrvVJC
BdxdAY8SpQjFSEMPEXYObzElvCNu4dJJc43LX8bvC8N+GRMhwwv1qmhruPo0De6SKuShXTfbbqHZ
Ol30OpwF2hPIevFYZd1Pvul0rlk0quzVNwSSUiqB6d7u1b+q+Fzi40heYzs+ftj6PsO2redEdiHd
6JPpQrKuG12aEGBuGqQ0NcEHQGXTxxouHLcQFK5H9K7Rxx9Oys0gf3B9V+CZteiNdCBT1bECJ+K4
BMhdV/4vV4LH3IwkZdRZiST8pSvOSVExuRV/6MWHHVUjdVti2L00c7nB6vwQSjbK/wX4A1O/ox5c
RgHJskQH/Y1PzxAySBAlaFEGmuXbxEavXYBdLcmhR08ZMo2cpPmRYAn+Qv5kgfTmg922XLDiK4LM
TTxsTShmLALlYoj9Da53kNUz1DU90G3ATxdDUcbheQLWl/2ER5yyANxq9mjgoBlQR4u5+oP2mGv1
GRQ7b+D6DRrrm8vrg7q4TtR7UTtAGBuSl3bHP2rXuhjjnTawopNOALCNQnry5SdCwFwqi5cvCTA5
dDKzEdgFmMfY3OC4JnH2dKhu6I1+AJUswtqW1RSopigOpcEp4CPydkqIMliEVdUBot6waN+KsxIV
MbB9flSP94CwRekZHsqMPi0O5LpvKZgbVQkx/0urhSHSC7+EHdd5oc0CMvnVQdAC+AyfPSH7jRLy
FB5ETDTGAw6V7oj4NoyhJfoLXe6VwM9om42l3ERPe077v3E1i/qjQal7/xoUcjjynYsROzeZRKeo
QBoP9VxYDoB/PTQ06ChqZbOiaZ4SLOY/p/s/2y2IrUbJHnHvFC56tk/AoxwScHS5bCeJRK7XLts4
OMOPahZhlYsQcIuASWRjhf7IWr25cIzuCVDfN0+/fRBrVP48nMfiWSXA1twoVP0qRc/+qjXEaFYg
vfPDUdMcIR2KlitAcXb5GKVsOHn5WKHQM97xLEdPypfltsmU92VUJDrox2/ZUr6So/qfofeJXiFX
9sRdMRnd1sxfrFYNUFo4t3R27A17tKFo3ki3MyWC2Bd7gmjmy29S9o8t+8nP7aB3all3bkbTirwH
SXpLtCVeg9NviC7qSr/j/O/qPXhaM+qDAUBhQ/2sFWqz0Bv+oqOUoPC+t/s3+oPLMZeYlLYR3zBQ
6sOHGxuE2of15EAgGt6c0QS+ue+dD60OjeQqQlsBPN54lU4WLpfgsIskIr7HPQM21pct/dSWsIHr
u3D355CNsPikXkVdZcX+ufxO+f/n2HKNTu7/FPOqOiC3oxE1W4zSoafdILn54GBMmLaudOE34xbo
W6Ks9OUlTEqUtbcuz6OiRPuF+GV8+k4zcdi/P9fBWoVGnoAd60Ana1pbRBvOs+skzjTwwrWZfNfQ
r/NYcIn63FiWcAk/cqb6dMmO2pGZqxJn4Hh2/9qva/z8RokfJxiSXz0m8UyDEx39fmmgGq4gkDb9
uBwmFOP2gp7CuX4tE1CBgTDQYRNWjMKuzUepgYdqVHbLoFMIDPbDrvIW5UbCzbWZ79ShfvS1sZPu
2vcj5F/nY2MBWAhsEcjSS9Gd2heGo9UwCe3YjHJdEZGVixwUZaBG6WYb/u87ckZUz6oKKpxP2Waa
ccZvRpVKdPrThn/IdTIO7q1d2hQz8yzoaxFdNsFdVx+rbNc5o4OZY8fJwCrRCQ0woKVtAsMedgBx
wXOAU5nQIPMLCtkBokPGJ9NXhWlSUFSZnOZHYXbMSd8KT8h90G1oapFg4erGFgiGigvg1A0defsT
Zl5kpQiSEW4EYtxPf33eg0jcXKuNalt2yP8QpR5iLm54RAS+wr5EEsiJSRAHI9kXyaXMKINakAZS
Iy6Jb3MErGTJWTxHEe5o56Xchx1qGB1n425bl6O+kUWP1qQ/sISIyTIIiRDTx0Kjignp7EUq8iJz
Qf4vpv0hoCWXzpmh8G9tZ2uEVkm2pp14mzgGrjDR65DeWXzcLlQ+pGQI8681L/e1cSmWugw3W9Uq
beVjtPUn9fUyBY10wSvU1rNl5eb9aMajf0Tjmfnl/gnwwZIQIzmLQXOi9XH7iVfIX/sOrMBRR1rK
2IZcM36ueuAQiTQ7nZAbhpAZZha02+eCVs8VLjqjrnMBGqALhiXn6NRgEvvPgpQ9wqhEK0WozCYl
FrySX7xTNEaJ0ufMckimY67j3/DNR+agwBu74tJlyHLzncGo8VdrdA2zNzfAseNXO1h0xYt7DVTX
X1yrxQSd1TR7eRwTp/WcB/WacZYYoAlNz0aO0SbXecUQnU/uWWVBtjP19+sGW6PFsJuoDvycV95b
/OS3FE84gCCDb5PcMZ2mItokVyDQPhgb2QjLM0GtyeWjdKbsDmdF5oXiMjr4+ZB8sUXnDh0eTUgC
dQzzZ1lTG5TZV0S0Rl+3fMhe0aawWp0uPTX15Wpwcw4SdfBlQMy73snlBiTU7i6lpVZ690aO+huA
MHTj+71Ptw4YFQPq1wPRQs3uDC0H+vEFWeOFc8AmbIE1RC1+0G51w0SGPWYVS1hXC5w5fm9alYgu
LhTHM/xIp7R+8BnwqxEDrYAd0CNhwtR0/qrcTeyHWFKRT6AAnbN13mGpnUGHgxyroQ2MZTjoWtcF
oBKP2X2lohczVGd5aHfE+Ul2mwUlfJc5DldXMX/4lqHrZpMe8LeSEeiRJLDeEulBEYdTjWjr1G96
V6jHt89FuHCr4yCO45jF4Lcqko75efgMAHWBRk/9HsXOPow7Y0OpCP1RquLbE0AwrRNHg40KlZOu
ZPITJ9VM0H7944JQBzi1x3WfXqnsZnV12B7VGCDQzX6XYA/SKbNF/3pY4CorIFMfNv080BqDW4uh
nuLQ9aHf0Fa+p+k3Gp+KLweOLRBNyLi2aMPfpG2XWz4jJnr3Qm92MVlmn8duq7uMo/o0/MfIF2dl
ZTH1VAwGyvd52mdp3aQqoDb6dQX6ioJtbbszg3W1LrfWIp+gbHEHAivxrCI34YIzTvL0qo46ydi/
a55Fcqu0Bk2vANQY7RIH36S8rHDmUXNl2iZPCWtyifOfUINO0DGf3lpdanNA9gGbfkcJ10/facdD
sGIeO8jgOkSsPElN5nFldQTY+Jhm8+V1TSNQ5V1WyrqKXLZ3irBSK08tIKxErxAa17U3SFLPLjA2
O3nYw5uOAJyNR49NKQL739CUAUz/NkR9No0oo2qM250UxRSutEvwIUzPi9HnDebveZwF63xPdxTF
0N/tQ+OU1N3E0CT5HgRwDoEP6+D1DvAckoHA+RvydxFWdz5vmSw+gy1VtlXfM1H1/JMzfeC1aqTQ
5pkCag//MnW6gFajZviZpDN7c1CALo1iVN0grMuPb49ccQ737zh8qKrJSuQcAaSQ2JtjYHaezcp0
vS7g9A+x+6W7B2zv5oc8iejQWgODDdRdDKE+lkUOQ9+ugnDWtiEWU/e/Df4rstDUoyWT5st7aKQZ
gU9Fd9zx/xcHw7SlZ5gPdsbVd/iOh/BmNJ15nB9/xNW4DRKEH70qM1P5aB3XxNPfeUnTvPLFNmbs
+kxpldFgdRXahhH/YTPryGxG3QYG0KaYq+o/9ANZMQgcnyT/XA/BnkUyGwurenrCujPBqRvtW0PW
XvIbnsvWjE9YQRnAs1uDKOh8kV/zO4izcO83iADWS36Njp8tTsntzuozIRLEXGjYiCjFZUYDroh0
Oawg7bL7VxeEe3U2xuLWaXOFUHGHwvvRsTNjDmJv+KXZqPQDkRZLR0RnDu1VhxyyS+pKy2h5lmpz
JWf0lYFDKmrQX+yWnJBjwsREDe9i9NQSeGkfciAJT8UX7HDDhXq3tMQRI2AX5fVLlTpAghhNzq8x
we6d2icAl37eGQ0fmpFR8Yakto03XGFu1+7haTHgN+TK6gCxYfqewQsdbsCBMa2++J82i9ZnZB6R
hHCHnXZARubAPAErzGEi2UZU5t8wWAtiIZQMVc2tZyMlg791a2Mwl2ieLC8R0QAV8n2VLp3hDy53
ORXG+6yHm/2OwKFEKFHzCeXhLD4jguw34LA4IsZBccnlszZlXjvhs94TP8EME9vH+Ct1K1GNnWFw
IQHEYJi9FKIxGgvsY7rIsopkWh8/i0TmL3EYU5Y9mWpY/NZAL30sd6wFOlrsO3dEw50v8BaJZSSq
8ry9TniOEO0k+utctlKG68U6FzTEYwa7jrUib71Yi/YZap62Bf1acDSU6CbSu7ZZIpcPSAXaAe91
Pj2RcS5HoANxalu7KDNtJqR3PS5+lzoJqkUV/GqPQKow96QrJcf+F50jVylbRDoGxpPKBOvK70Ss
juVi2Hho7nDRAWL0+YcPHPI9Aj7A9yIDFffniiXNFqSK5rwA39kUgE9/vQKukdhatM60m5PLyp2C
Uef+WKHmFg/EEAn5TAsWuRZyQeBJvEVUFQuHKbYlJqByH1tzHaAH2nDHQMShdFx5tWtyoPSYFrZ5
Ht6D7iMjBE6wzfubvPWV/NzvP8q12YUmjJaT+j/Hpfn7B45QhzHvaHEcPGptOAwJ5kw1NWKviB9z
1HBjrdiKmhRj4X/0DgKZ/dcUAB41r4xih7JsVE+4vKatVzxomLAYdX/r9Xlb/J7JC6RCa+dSmupj
h2wQMOYsVCcsZwfgg7WoVpE4NZIae+AMJ1h22MtAC7US4Qo2J2VKDWAKUhv7a9kdCtxZD22WuhKl
qpnzJwT80GVenDFZzfmZeki13R+/SzWqulsOFE/GHRw7jX0uZCtwMauIznyKUiEmByGrU8aCJvt8
JL963lu+0jxS9Q1qh1+PMZ8Su3Z/v7VKXs23ET8W1M4x6Co+9P0M3P/DxVd6sHJNCZQZZXHU8/DT
Yj5NQ1UEY4ZrBz1TOeJl210fZOXoCjxTt8YdPaLGRiWcK/N0DMv2k7fiVLDu488YxusUMS5ll7Cc
2uRFw9FaZYn/gv397ZHeIVNzUC5KCAg3DUzTU5YLUaZlgvhg4sXLgED1uzWctHCF5UGq1HkRsxDp
zEoikh/IbYhxlr03oEy+0VE8XR41ydIe+6MwT6ZK4/e2CH5uecjo5XQBzYAfnEoiHYC0UtnQHG0z
mQookXLI+p6Lkqk7Gd4HQZIwgPgZxy1oV+hX7shFfSKf3O+lV/SA9pCMcah6JemnLVJKP8QZSnQ3
REccfXToY2IKXxWwVva6sn/+ioe4AdBT4Vq33KSdS2XGt67lLjbb+dkrEtWp6p9LBhRJpBTC4IFR
AkQSnPpqdFsqDmvqehabYapzB21Bq1paCg417BTe6ADflE7AGS7jtyHYktrA39FKFVnrMBFyobgF
+fSXxrpmNWd4r9bdtg+k0ePUTXyx+ROQqlgg6DyrqmeoQb0P6iLPMe70Cf4Swm+3xxBeHCghl4aT
eYunVZ1Zn6uO/b8b6PWuXcYTgErMHi8cZ6cGCpjtZH5L0jUcbTjypP//HVFjfIQWxn3w/K6KURjY
gR7mtCVkFSONPQ9C7R6n3UviNj1S99o3xGrrk1aAPzQb5JE7LZ4OH6HCwxDc7GAFEv3SbtT8Mx0t
dGeOFZ9CKuTb6+7Cg4+P8WwMN9FIwlxMekOrLmQKbR+HnkWGWQC7gIeO3DGadnhVB548NYYyt9MU
ZycSdvRcSUvZPLH63uyGfW59zulPJjObMyikSBUC9QjSVLJxcJlLNvdo7DPic7DcPirXSc59NfQR
PTlTXGuzHgdTEoF3ixe4ISoGnUCWBEg6uC60mKNiYme8eAfTzliaEVYSOWC5LoMa28bq9Sw4uSjI
+PrS+nxfsNyPcpv575uCkOY1kOStPcFWwtGWSjN0FlGDOcOGrkwi3KsPLsaOMwr13XhXtu0py/IK
o36IdIBVBF4Bc+4k6qKau2CC508pXZGcZ7bHCCDSJ/gW6yKiMUdR87S2sY0mL6vtSbfxQrq3bfHy
y1JRwOw6EHzi77dqIaiJc1XtnLaH7x5Pb9zKSPGVzQTPf7bLsA5jGfy63iW/BI2E3Q8eOMqco0zd
NcXJn+oaVlT6bmXtGfUJzCMT0IC3mfUTk4GctaKKg8GuPSFl4be9Bp59ckM6iuHtq+k7tDU90eqt
afUujsTZ3pKVvItntJ/eYDD9YpPj6Q3rdDNTzC0fXVDJv2cQWtNS9Q13qg1QnPvzyNGhHyKOWt0z
u0TVqbqF6kFGW0xSl5xQPDEoCGzjlTcz34Jx0F126Wedx9eT6KN0XGRkK6hIst8mE2gqrscYNiwy
66Yr60FmILySfMbV2x2XE/LeMVtnNABdnAO8pzsw0K9BcLpXl71o8dHVcKtNig0xTkNwNbcUUO4k
CVyCBwfyq5lG5Zw96uXfi1qaDXEcp67NxG6xhtCSFxc5WaTVNMtRKSA3al8r94aUl+bwAfI0cF+H
6vGvtwj7J5EW4QtuUaJtfHAftgB09fZI1ffMvBggIdx8hcPiUDNmhFUeN2UqV30RXX5ue5rMh8os
TUXTVJGVZQC0NN13pVSEwf41Gt6VqzPKTR0wLTH4KCjTMUmUhwf2f7S7wD6C/WXFRmDELXaE/vPS
tYfoQpXXuuMUK+dlW6IP1DDLDyT9t1SmDU+OrFM1YE4yofPfpIq2nqFpkw0L4EEahGOG2UXPTtuh
iVS6df0v4xiGCVo/97enZbEBP5HLj68MLGkdEQ4dzireCPbFbIVSXllCbkc/tD4522sZfQbEexwQ
XEiW/jBlRV3Yl0kdiY+3FmXkBHn1iFQxV8SEgM1myoqXuiJaYC+MDY8HQ2K76X23xDKixfE1Mr4L
GW2VAd8w4f8nFO3O8DWA29MRyGosrPiI2rI2n/pBU8O3zE3ZKTV9bT/wsLQ2zxsBE3DnKGmtuLtW
o8VRhydwwkbXXJskopF03ZktEqEw/IzQIqrFK6/A9qrwDY7vQ7P0epO8CyTUUY2ZXdgzuNzOKOpF
c9iICKhletUBhV5jvto0k2e5ag3iIdeC1i+qHTyWY0AslBXKwmbbe9r6Ch9YLOJPvrNPj1zliyfY
EWOEbbSI04HYykA+NCv82/HV2A4EQVFXww8Kmq1Fry9r7j6cZIoEi+Vf0vr9pXPc7Gsv6LmycHo0
GmYDaiNBgQCaVQ8LAze5PdhckxztZw9QLsakh8989uSvphGhcsdXV1oi0Vne+vwS8SPWoNQ/j+rn
6r5mG4BNCmVHFATZNTfFRKKFdteQ87DoyJagGDyGc5eDiG1uAWfy5ZZCDK/4Bnuz3KI4P2d87mjP
Ec8ym3NJj+JTWhOSI+rG4f1iNeQY2hFELQruhLJJVK05lGqIQ88ArLcVCgHanez2ZAMLLNN7gGpN
rf6tnRkZW54WAAgt1v8GZFxme+XnaBhikg/Ywre15NUad5blhreF2tLPjFcprWFCuFiFB48MLGWk
ZXiZk3wmxmmmPnT9hdDxZ+G5q7juQoIPdtH17PSg1iIthS+dpgREH5kPIgD28plRUK6ANSiADV8y
pMed39QVQ1aXDwZXrCuyNYpO0+ybIjLV7Kj8CCMiMDEGzaVplVmT18wQZDquheDJ+mWRctoIVfhl
vpU31Nh2prQ74o/I1aDS2Yb1MINCuPVgIwhaQM/j1q9bqhJygpFsH45f1F9JOBJRNY78CuBCciOa
+MaRTdEo2PWIlrz046HtIWO1vLGvZuatS2idWrdtzbfHySAVKFnsy22xrvceia+G56q2FuUtkyY1
itaxPnjm1xjt7Wp71as8C8w3gIB5LtVSLU2tSKEqZfUEq0wxp+f+BIA29ac+iOyvZVrjU+QwDiHv
EhrdKtappmVEXIFF5l9JmeSVUoBu1LVEUDIUkY2FBxrwIrdAo+ToVJyAmfND7EwxubxI/H4I02KK
Oqyo/l9oqtKMx+RT8E7sjVetJJcfq0dwectlGWyJoBVi5AMt7dnwBqESCFO8M6esUObHSWBTDrSG
bwSf7nsOogt7QE8F5nPNytEuU5a7XzKP26oE89Cm9cOicsMaTdEly3oo1D69Nq/nVGZmkJr+5868
yb5iu0bx64xcUKI/LotvQcZhcIohE5pZbq71jAligZ7/9XDzyLAspDpRMnF5wmREibrgD3lW6fqg
e0bdYfbxveSPzQByMNHXzipO+N6LcPVqF9Pr15xDY3OEW/5T59B6x14ta3UVZdnmdohbW+9J80OS
ziK+Mmld+0lUxCxE2alNbSmIxu/EBklyeYJxsuZq+KgIFFCDqknami9KpERzNn/c1ZCg9aMO79Hq
AbcVpiNwQdgzQehETKQ3UJfEr6kgXM/61mPRnX7IvNsmHQu1NSJjrLQ1Ntcjio1ukRw66V5+oLlj
/Q6kMI7xnckjYfMJDY1xZT5z3+aTcbwWZcvlkfb9ONDonp1htQr/Ma6TX3Se1zVTgbybbWHupVcR
NrxYPhSBuL/WrdiMuzLUNIWOTAGI7PcMcGKIBpbPGV5I+aFaI/WI9vzLbS2zpBKgohHCqFZ83y9V
Yh5d8lGcUzCy+J1QkQ4xo2gH8U0K+/5LpRQ3Y/EoJML/AHysKqsMdqPkjX7mqy/LRFZZ/inyURFG
B3ziS7q9G1UYry9g4cKoth7mU6nFoH+L/JRPssmnC3mww4D9uqvW0bY89Cr4VX8LaZckdSGSBJT6
etJ4RvokMvUuvAghVPD31cheC8UtOk9jZrKX5ri2tYYPZSQKayuEFM2qhIVq4tCyRWxvhdJ9PFH3
tgocb/nUDV1MHYIC2RiB2wNiBUtjAM5wXQN2G/b7tblV2stfrl98lNucaE4rt9cWxlikevPwlKdw
+L3x2/X3FzIS/gpdKJSTLJ12xRcXtOXgpm7zowkfZvb2jUOfD0bn8vccVn6umzoyH2le1pjhI7Rr
vcPNJt8NM++U6E4vu51TGOydK9sf04MShSxA55CM2ApaRVwuUuOyaOcaeKVMgBPOE+kTnaxF93vL
oE90nesrtXLUz/cFzifHkzvcS1QTsjM99azSQvoZLlUNJHhqaeV5pG0YLGzy0cCQ8PLdqbw9JuS9
lcKDbDXbz7C6KqtvDExF6BGc1mhl7PIR90LsUBRWHcFq8yCBVS/GWyOoWORfEKlK37edcmvVBBeB
cZ9yCB0L4l7Hc+pUo+pl0urwH6EqmwNt9kpRY5yaqWGN45+3ywgULf8T9ieTvZW5hrtSZ6qXRtQb
MdohRQpsgjtamTcqCMXOqtAG4IcJP7vepBudqX4KLcjLRrny4o8rn1MdWcJrusvg9k61Jvi9kn87
9/KHfec+ynFTvN5PoJLVO4fCKnptF5sey27Al68XdnOtb1t4A+094PCVciE26gvcU3F4ZpyM1L9G
rTbmjoN20ZTVg0jgYT5NdhqbSddhMlG8phorUDamUU9RNYYRaLXThFVDWf44fs5EzKKXp/reeDBt
gueJ3IM69IRfTulxBTzntGv7n8z6KgCiUzaD4aeYHN5T4bQZi3GVF4/9emgn1JVoYTx55mQUrNLB
bIy3YiGQSlGXX1B3ZtgalPprq+9ObJcjwRzqzYLdWL+ff+F9k3o+QoePemX9k3qNdn3v1eJdx3mf
OTNMfaaYiao7af3fb+qEAfHXTtwFiQX4emiwYRhZygrvw99g2RcD433H6N2t7sVILmGfq5k6eIdd
vqLaNE2JO7BjVH8tBGX5QZA48zwlCY0fMvJ6mJZku3eIqhupbfFPehDE0ND4viN4wzD50BxuYqdS
C6j0OsQ3T6DCqMjC1TYKTHm9+eNTQmwVOhnDqLOg9yFWoN9X/Pt8yqQcvN0yal7yd4fEOXdJ2Ah+
F1VdetoQuMeZK8s3HpnZVYkQ9EZiqVTXmOFKpZEWFAs5HJ44VyBNH1Lxut1XIOWLxOhZP+us9Ocj
TocC+EaN1E6IgNpK6FxDn4Rrt7WOMUOzc8/sL/LjClYOu/fX5O8HhNAEvJoHAwI0atzYUo8JH7aj
jyFOo1F/713WR80vQAxbVLxSHOruvU9yzQFBVOrx2t//e6R8NjEq52FY5GjuMo+aKTuRXvrxfVC1
Y/HEIVQ3VPAPm3WK647RqbhdvgyDSerlejhZBWzkAer0oKko05GhOBLpArbdvPZwALdWRR3kjQQd
5q0roo7MDNuS9YgsRl1xFG77bE6capIuWK5+P4jkxOyZnFio8wJJFoEcvnZk4NWsZMPXz48yRtxi
Arw8Lu6Arrl9SXEdX/AlWzt3C/M4Qk+vCc0W2pIuF6UBP1/q/zAA9ofMF1LGTIkFu3s+MGhtVcZB
sJxyBBuSdQ+FrIPZQ95xCi4Z3qP1/FcbRc0VL9mhKsL4c0x2pAHXYxi6C8MZIdY7MY2MfYiOBHCg
tMoIAatw02REEnpwrTSHaN5AYxmOUFtOju6a0WGhQ0hfPrRhF1sxOwSG7mqqaCfJM4Y03ZMOvhvi
EAK/ngp+KHiOxDi9degrXm1KMlH3kgDDssb9ev95I0ksmi79XhKsd+062XNZ5SdNtGx6R3f8uRBI
qJXGedd7vWFNHa44ViYNrtrP7Ne+sO7bMeKQO5G0XSkezy06z9kgsfrCjWN40LkY2Q0ntgaj251N
yVxOdWeO6Erj+8KLS+InA7q9Y/aSujbk5EebCfqSV3bb/LSzeGhr7Jp9LFH0wCnluUU2c/MQgR9r
L1e2JXEh91e5ClfU8NJ+/GyIMx0HRFGUnuguAL5ozrdL1MtfInF/hCBPLg2q8CIX9u01WMp/oHZk
sbF/qYMcNdcDib1gMH0DS/llc/1EmGS32QhLM4FJVdgbvz3MHcfP/YLe0EY0ioFn5ziYvheiXSnv
r6NpJAf9TKtpYeQdWL+EEyaMr0N/S9qqe3Jya9gwnqvaAxSWhr3I17TYwpJuGLuQJaWer+UDkiaP
rUGgma34ZNAq1kjXsU4iEIP7yEMaZ2OsfrXMT3e33Oaab8aL9xUGgqjF/ER9NcsX3jTNL3oVi/U1
zeTF/TKbhKRKQGZM+Iwtds8lZn3qSn6ITcx4k6SeUixivuV3kB9nroRydBRRoJRcT1R84z5rDw+1
H87yjyTSBn9SyNhiXesfWvdTW1p6htK/knrgUFnd1pjcYRfgS8M3r+Quw8QIvMxBfdL/xJ9ilTeg
RqBBMtLoui9FsS/9EyaThOGMRCi9RU0lCagS82+q3qn/4ARbNxAHsQy2k10blJAhRSa2gt+cyRZ8
L+849tPpPm8KnoamgLlXSbtugz0df2oO6wEq+mCzNEn1QzgtKPfqX7XJWd/EvN2JP04kWqxmldaT
RLQJ7GvR3keejWYEgSUNB17zqgX6rw2fcX7xAsdvxXKGS/N8yfcRuYNtrB95/94o78UkIzzJ6xRl
HLUtlGNqOeJjA7yPdStlgbKEA2/a+UUCMpVq1dZvqMqw1POI8nO/3WDCyKd7peW2MH2NVtf33n4L
WqGHOcwyqmo8YaYxHd2aFFN2AYc/MxXRkkVqRb5KUSs/gCyhOEBPFCRuvdxzer6H5+2T487S9Q82
D+r6IQBUPvmltwsREfFNh9DLCgHKMEQiB6mxyVWU/SyR/FNLYzGWmvVWSLMXdVTousvZv+v0fA7C
MusG7hvvJQ03oDVPAeAsq2SISjbVaJ0VgCIplSUjxOvIqDeH9Egz6yT2m/GhSJbbTPEZiSmiXtEw
73wk5DDDvpqOiQdhw7Nufzg4wVEeBpeV4tWk83ioICsjZj6uF9liylsmnUoVqqP6v0iB9mGky1et
9J3rBavCZ6dhvnmsHpFkm8fKdbj9zeSLCHrrgUvuVl+kAdBFeADhrfWIzkbPo9yW7imI2yx3j8st
172zn78U86OR+eobEYVCnDGXxbaE48P9O1JP8wysMRoNzISLpIuaS7dLDaMvw9RW3rBMNds+F27H
XvHfADueg42RkiAJdo9s32G1jDmUa67fBFerBe0+ZbngYzjy3lNg7RxmoDLIKtvDzH1hG3TWmp40
IitgQvnU+z8W+IrA2ThbPClHatsR1NrjpqeYR+32P+hpRHxz8WIn+8ghDXCFB5sHn5KCMpGWo+YS
m1ZWRDahwLa1JxuVzaAp+nVQSDa3gu68IRz+ByT2BLmSByvwdBETY0c8H8tyA+od7ydZOAJi83iV
M2ZGRaduN3hEVEoestBDqsNnywSX1EuK/BJoDvzmRnDFbeJfFaeenRQZg+yanBce9+LU2EYD2G6t
qGMBNyWKC7PYJrL1aaZ8UiLVma6pl76+C3HOj/ATmMDMC+VzDGufsIN8irt638kZ/jSbublbclq8
kwTpX35jcYwgz6a9TNyHIYQ0wfC+r2q6wHVASL7UNygTah5tWyzZXdCgFpqAWy9M4fzUsv67moLe
hlTIDXZRbqgm/Tzs1N9hqAewDAqKa18UewDllP1g3vDjjqnO8rQ6OCdA6kqhem9yx8LSmHDkzLh7
01CGQ60xeMytlK7O1n/hn9d+2VsRI10qwjQIIqP+3RMWcnwiHYVcHdoDkRjfQGlDaH0shnkDsycM
TUt3v8AdyBf1j9Y6P4Wa723GSocNC9ShRk1vSY8eJU5EL3jWzazFRiB8KPu/1fGH7C108FkFyHBx
yiBgOP8fKWe+nINuRmh6hanr/FPL2spyYQycgitOIzYjzY1dxCrpjF8iRo4zdvokcYUV03lJ+GcR
KRzEqnmOvnwByG36MtKSolb7TwInbk+xm20FrfzAVwnG6zmlujG2rnqSix8zA2AlmA02ek/8IhH9
+4Zh0vUb3DwuyqLUiUKay+l+P4OX1sOKxfxnJDvGJX3pMtjqEbxzUspa5Q8D5qu0Upmhn93Jb5/a
5Og08WPetBUTlz/DHlEb3J3guvAauGSr5AdPT1DeuGOPr4vxTDcTCZoUhB1AlKAYX4uc3YyyhAXc
DovUOgURr3QTWnzZ4CWrOKFmPiE+CKpdv8Ds/gwErSFh6X/DQMmy2caTrKcE4ysKFuxT2rbFZEBg
YSzPGxL6cHH5ZVDWNYI2qfs+jr7thNZAvt8BB4DNvJ67vpsWbiydAlD0L0nej4lyyA8+NwF2Z8rt
5Pk7pQw3Yy8kVWzyDMKgzerofpjbrOgW+K3E0yrX7ah8mko4/7JZ6wNZYP25cSKa26zGWpLmX35E
klmyGLnPJn9Os+RIkC9w2LkEEjk/ueLJE077t+SNZxgpxxt6NPsCNUwfU5Thtturl651m0yDha+F
b/xpAfB7j75H03er1vtJaDQTY1Gx2NqXsN60El2MewSNZNU3msxghXJqYoebu1P4oWBtZGM2h+5E
NJFHGiIH+edtmppdW5sMu82gQhZKfJn6vie+y6YK+6z2WxQH049z0qJ8Yldgaks7FQIQ3krXwyWG
bHcgLU4this4jNkxbHFX/W45Zs9lTN9sm9Wu1Pmsjin6ivy8kYYfEkoRBGr6uE56c2D5hp8QK7Vp
xkBwbhki6L3D2ir6F/ON0qjxNh2VAUb9Pw0nGndNopTxhzpfvNaw2sqkuAyn8YHVrp6uQ7foL9QF
8zBzGS6I6dthrvTL6Nc7u6ua2XPXNaibklyj07cAkLG9Ca03kO8kFEIxKVHufaRpa/ya3+W2kRHI
TCnfLU7akcBkSywrtx99tLWpks6yHshA0UUlf8zQ3ivdUtoK9WMhsYWL92qp9Mdt6dlbTz5uzK/2
K2lJ6o6vXkavoNSgqwhMEpPAeQGZlUWjuEv/MkeayAVHdlwGUTLmsLQz3jGN2OscrQR3iqe9Tv5c
xC5iCwLgV/D48W8scJwTzRVihcFisbzIQ1jZ01iU7rmNeNjV7YB6opqagEnOP1Mi4yDhRfLWFBe4
gCI3YNs9Dg6RWRIIwIu3p+zWssRzw2Uw5tBsnL6NgXZkrq5Q2XhI396IIGV5C9jOLO7VwvBBRtc2
uxuhOnSz0Hh7uFmHxvAefEcD3fXxsbCZHY4J+G3KFQkxIb0eGkQNf+4rjG9BYIJ4Q+cEI0fQvkbo
q/sqJ+QzuLpcU0ymUXcZvbfTqfc9JZQ061Ix+vTAGCy3zvVowp7qSi0LAk75Mj0CuKyOz4WtBaf6
WmBrASxdvVF4xqZuUNSn9ZfszbSxGVjnSlOj1VX4GcDDTp39Qg81X3FRpZYBWKKbPQdmQJfU2Nw9
1qEMNufIPa1HNeW1FHGxheWngKG0WP0GTFAGvaf8N/g3bsbI1yCOwB+DPOvFj7rRz53DYTPg223O
MRSDRNkvnt9wtPZVbjmg+RKB4HniH6CeGgHBxDFcCjDwwN21GUxikupLW9q/Mdg9MRKeC0rwJuVI
pdvqOCh6Y0/2AbFXcraqx8C56Tl8xBPlORqmZfBUtC4dvIFOOrxeTXKiU2gF7A061+Pcljafgxmq
rIOEWElpmM/PdxNMDUQ/58NDhzPAqUsfi76emnFng/HY+jj044A06N+uoO9Y6AwRjmnwsW1bOEj2
5i+PwaHMogY2UKYXcXbca/UX0956BzOv1Lrh+aeEHC9JNVPvPlWoqccPIjRd1PcSBwTJHuw1ZcCX
4yxoboRCsXp9Vderov9Zj6a9jm+iv1uSWwLsfo9sx/04QJ6M/15w3GUAqRhUJAodOB4GHL8Koc85
gBGi01jdhOG5SZiA/FHmz9GXHyGpjBPpuZHyq9fBryoe8IdUOWBEzEyyPn5OQVjuFIYZD9/br6py
aeDcAaBihf/G6LzUQrCDmKj9jMlifZMqXVrB4YAKkOLCo1CjTaOP2TZOzfamlmNDLIPN1kcgNLi+
OHh13dLwPUpA9suZQBrXDk6XUz3NnUJV6kPDiNFESB8EYSasPb2S0iB02dfGgz+7taHz3UzXpbyu
vD0NVrXMgHsxyK3F/8aKA62/jzsB2K/h0kxilQb4iy239s8T08PKhnAPkg68ZtAw2exxyYBxysCo
cPPVX2MLW/5HLJ5A9ItOvJ9hWekzWWyeWDUWU4IXbrJsRApN8bTVxxWATHq5kHd7jZFtK4WsW//e
XEP31+XBhQTnqGVYDvud5SVrGzHicDY9rw7cxMSV3AbZLoPfXg4hljv6WVFIuhvXSf7CkU1yTiAB
JKI7qQQZd8Ub8l5Wz0o3s86k9xye31l2lWGMEMlRs0iGGTHndUUQ363FSRZPdy18A3BGIoIjo+ac
JgvZyXtcGfwL1cQWIYFxUuA3fyJ5ZBA9384uMSnht6HREUzNMoxk3Kk5pxqJbm7VkQyR6hqkyC17
KGOxxodj8XTRKRZn85fqoOTNiyYHtzwk3p20iEwLAmBDyGawxIgV4KpWK6uOpQ6sP/dJu8TgjYfB
F/h59JvRn6zwtImseSB4eV3VSVoUafDidhuhk6xOhxnqehBlhCBdtSUXNNu0vuR5WeOs3OZVTkZZ
HLO0Wn4S5hpxWvkLUCakligqj2wKA3mKkfnU2hr+dNjI750SziaGHA3CtZ+n890MhCaqSsUNdeHU
2CJou3KzmAJk6+O4X/nCPDSuHAMjWtFOAUitE2OI/Ke1GtNuMuAGY8N7Yc9bAHBT8nATmEi8hi1R
CAXAVEMVF+XDq+DzskBZBZjfnpfFHG6wk7zIeyXu04ol9jKdI2PovWAT5Ym1IqWprh8er5NC0Ne6
jPQTFi40PGaxxfxB0B7tRAixzdda5tNGSiULNyRM/MbyBPBnVSvi8cRbkrxIyYAtAjh8GZw0k8FE
vd40x4h6phFU7/DW8wTjYGl85Ry6/tPX2jUDbjQY84DqDMDET070yfHUSeQpxI8MRLzZI3nJ25m4
QEJryfZFiUhk2wW5YhVWZqvY1sQzSexxNpzgSKJyi5ZLGNY24UK7zhnzCHoA9lY5y1IOfX/YF/FI
wRMZO/2FaU9amqB0KBW1O8sMOuu4/clXWLwu/+FeNNwHLJusWfBN8EcxljmEL3Twyh1sbSS+pmcZ
TR4tpsLCMnSdNZjg5RfgsTHTwUd5PcL1h9sYF8yrYKlXLI8A1J2ZWzTr9udwmzxghMWZRn2LIYoJ
JQ40T4rISHVi4vI60lnbOD8bQE4c/IP2N8DKI7u+E00CwPVrjATyAInrwoBwxLKLFuqlFq97g1Zw
FyxKkBcMCf6IPmGjTOuEid6O2Bl1r84qXGMJQg/tt86akl8ZMuRYBO1Wyf/t5iA3LCzg3wAE6Ttq
bjQC/1GOiSRQCzKV/Xm40wXIivJU/iURwbzvFCnvJANsZlp/nJPYbQirE+a0mWFp+si38oo6hm2X
F6iR+ur+j9x6Ix4br7+tWSOf06dtC4sCqetp0whvXaXJZ9+sqQe8PeNdiupCKWVZQ3DsT7mdL1yb
RGsbGSEJjbdRQCC488lAvCXfV/V46c59U7QXCi97BuMY2NJ8CKrnpzrkYJWH2gl+SIeZ/dfRHkUR
MG9wVAino/RdiyVpZ6MZoQWhfP1aTLC4FD1IYg4uPzrNjJUs6J/Msv0jY05ZkS8kxalJ3fxmYXB/
OLIsCUU1xtJTItKM01WaX8Exn1d0WZr3l2E/N2pWNfFazg+mG5yysru/hV7Ho16+PqpaOTQpSfSZ
KMKWITiHEmBaavXeOaohU2KAKm3XkgMmXW2ZQ15UlxlTYWSzRjFnS8cDSqGHcncB8plg018f0Rq4
JcmTTvL9xveWa9lTRdWgParzF7i/Q6MqFOUsVF3p04oXwoMLhz2H7fWs731qyB/fD4JreHc9hk9b
px6bNVllPU9vJCbjzDM6S+7zbdwBC210+h+sXpNmNsqyW1IGHWFS6D+O27RZHS73qosK9ps2pJCy
8bqfk8jtGa0S0v9CdBDYFrnfqA9uI7u7UOtMaoZ+BE/CttI8/UuPXdTs2+4z5+4q9Q1sEMfbGe6h
5IMEYaYoFLSyMBQHVjNsNdFMTF5fX9kK8+4X6eu0UPs3+vqhL8e8El6F9SdxclfWVtLnhjckKmzr
IXrRAfR/tepAIBB2gWVyFBr3KyqZIkG+38md7gAGpg0C2vO+BKIS6MwjK58lYiEpKbHDgD6ZIOQL
m4ZugtbAilXoQSV5EcYpy9Gnzd4J3fWSdtsQgFORPd6LxZaNImk8kCpBvsItKFUNq/NVlRz6EvgS
jq8pl0TauUrv7G1PxpY7KodiouSisqC6EZG5IBtKtPXE/xyC6xzA8KGqKADB/zGQrRZVh6NkRBGf
zKdqx6IgiYelvn27Otp+/AtEUO7YtRPQtuKwHKJkh8PJ8w3v8GUQoQliv5Uj/wB3G+/rQUJuPnlF
lkBOs6xHstYXluOTfijrxZOW8kuhQ+91e5T/CsZCgX8EWNH0YBJsU9Db12TIz0rFvjnA6CuxOycW
v6djV0oz3z8PETU0TVt0Hgasj8HH3UFGaxvfLXmU1VqHpDP5n2cksDt38joJlcR6aZ1thFomwhVe
XrO8wxwRAb/KkrKifPfFYjy4HA6OujC6liYUiPSUxNQjbHYgCUposfzxOk4hIc51g8LiVxxGvRFU
2QVhG70vVOmVVMaMpuKXn+wFocVQeYTm0WALDz1jbTTfZsK4kDSG+HLZNtY1971GnS5xA321em1H
VfEU1OjxluR1cGjYfLnEeAQrsNCzYbO/94lh9/BfwyGVehoFH1hFQ1bm94zCiTM6IUCn4xYsmfNY
eXiT45xx2Iih61qWAxedXggcj3OKuISinXXonovDApSLQ8FsQfOMkYg3YQsmaLfcwt88yqTtV9V9
O8lb666XvHhlOT7GJdV3EDhO+11/1ASHmAgqKIWxQyrNRVHyF4i9N852A7QR+oH40MlZe3Gh2Wbk
18mWNREgPITbJGx8QLNdsG1xb+5xVghQVJHbYEARYu0OTCePXJ/YLCNVzJuS5gGH4fVZuNDidgWJ
DW+0Xupo7laSdSop7L/dNrS9BwTVAMJtvYOiB8RFFKFwlroZfFcm5sjraNVzFaLxqtQUeSr8Phus
8Srq9Dru+zHg3lkflYgk19MY1Orlim2x0mFyxR6hm5Gk5NLYT8lvDUMaxZe/0QXbdgakaRiMM3l9
w+5fQfw/hdwBWTNy2QarIt/Te26g1k27IvvHuZyJJZY5Fqmn6nDny9Gt9JOwrEiK+IldLRx16odX
JFflvS2AbFRd+NHVNWrpRMU45jLjK2Ed0eFE1kNrEsdyPxGRyZreVJo6ixUgxy9VToC0CaUW+JCH
hFzqTv2rhr4aJSng9IEUXLCNsw75cVNVguLsoGuLWDGlQOZmLXuti4ZwHRKWQCqO93wV2ychST7N
8vBSRpLX+stkUeKU5rA4klE7A5oSC/cXiJXAOA3sa/x8q3D3o8nqBXseebsb2uRhepnPqmdei9Az
bIIGqzWBldhmr6Gm1GK2Yj0wQ5cb7yDp94jGLXY4qwSNVQl7cu2iU0B+CeaYlSVIWibBjKUdyfHh
hM4vAAI+5iwRDK2jG9NZxTGbc77cpKSqPNFuZAd3Z9vJ3tbdXD7n7uGcJoPcXvrzDb/9NI3WSKrR
UYIXCxvYV6T10JaxwsZvhxGGBN8huHKCF256lTc/6wXeYluLNsNfp2DiKP149Ssa/jubp/jYIDdL
1AqsgWvk8FqCSmW9C0EkzA2Bqyw6S5MldNLhLsldWvYJ2m3tB4EFbkb8yAkq2Mt7XzmP7FxRELiF
+eO2SbvIn3/+Cr4RjKCjh1+r3S0Ss7LkXzqpMIcbLDI0oY5KDvUF4+h4jhCiEaAzleswVBThZlyh
YY+nHssMf5ERxPh0ITmy/DtClifdVp5kM9r460ko0JfDxOqbUj1eAa29SDysDM2Fhhv6OWu89ntf
ZPeVfZmSr0f3E4RJSNOkk0Tnw7CdvnzHslH2Q03BMR5ERc038Fa5ZPJVizxfWmEoNIzXXdMHrlQK
4ZkuxcvdEzZjxNao3kFhCClMkYfew/1pKbNa2pxWg7TiUIGzO4qEPUeQMxYLtS/GyFUSi5SCrEMv
p+PeAHif/WdFqXGVQh+d3prWoM0FfECalUoZd/1F83lpn1MCJZWAKG1ELqIPe3WvhqzSNo9Udn+B
oc9+7+0XCA0mxXvG3ZQFxTvyHP7TX1CjHgM1L4om8fObHmyWUnf+RNiee8LbneulxjOpLarW3Bra
pDVeeXcnov+vzX4vTnb2s++JIly9gHTnYIxfZ2dN4PD/9DLTzIP5rdq2aD63MjD2t/akQim7+cRT
hud58Vaw6VfoaTVcGKYDbUCX9p0Yq9DJ2J6Y2+UMmXDRoQTjKtDNSkdA7nv63fg9TIpg8rL9BKmX
t3HfeiymqGxH3RUOMjIGkbQj6TAQN7tUvQW6aJGO//cz48ZXs5tBnXaVx84ZKO/3getdtt0nuZWZ
elGhznztg8Xb7jiXmtAzzpVSpoJ7D4AYT6O9Z+/TMz9AB0vCrFTRe/JdntqEQv5Pv6s+UAEyXscr
wsAI6zZvYYpEQqV3KmC7F9td9ep9OXOg+ENvrAWRN4iKVXH8vXAVmxNatLYVh2OdA4LbWcuQQnlF
VGI1p7VuipAutVItWy8U0OrhN5TK05M7aovfJ1HKLT8yIU79il3kXtPPyrtRo1IzfBZjXOILHCOQ
VTPdjqYIHPFB8KprDXKO2pu5wHM9a8mv7qSCHsy+/ErhdZEs/hT+i8oSfpG7SBlYLG+4lCB6jN2q
2vE//03CNWjce1jqp8yxGWicnNM9K81ehg0uB+3xhm/6vwmibqyWJdrrVvedkbK+YAd9uQ/fy0FT
InUhy3WvsyzlQsXir6/97/ttYkSKg7cxr9wKNDtfsqDToyxx+2qD0HQdjJjasUrZEZEvMoDoVPBy
yhC3L073N/FTc+sMy/W1MBcWQtx5AEXF5Hdjytfm1U35yaEifQB4iGiMwpxyu9ga/v7Ghea+SKdO
U+NjFrktyqIAXM77DZ6GYVODULtfEmOSGD8OTZJez/5fYKbFdXAtBnw57u4ayBoh6SPAiF51JsKH
7c5rRIpjRafwfqBQFZjQlfvZnbwp81ONsD3iC+GGfRKGnHP18WK8C9P3FEZNr+55Nj08YMELdZH7
sIxHt9H98utf6wNLPU0FSdTuriAmuJOYoN+gvYmHzOauRXHq2ROfdYQzWqhezoP7hOsZPHxzwQgf
fJCMJNJHAKEtty15Tlpd94VmIFRpclY114DFlwhNX9k+ksdGgbmEfS4KvGl662wC95mQpwC4L+Ar
86bm6FmE3mDvb8hRy3sYwrXOWgSE3HIoq+HqbdC8COGIz4SrWJKNYKx9l4KRa7vw0HzJeg0XerGl
yasGh73k/yRTUJr/0I9TjHR/20n6WQ2l5y3uedb+44o5hGNoZK9OY6hieHXLaN7K6Bt+CluuBjus
m9uHByDsSa8CXNGWQ0KaVBYHlL32skq4yw7YL9eR/SVRZKTuMTBDNtWcSMbz0ztNgZUGAybzX4Dt
zDgavVBoQiwfSoNMBqom2Umoku20qNTkWKc0vFxF6/iACkPYQg7f6qlQjLS+3SZHVyQpwds33Avo
FsG1WJESrQmwKjQdWLxabOvvTvD9ykhSL1lGc9AX8ahEqOg+t71UwYA0aYqgYnu6pbAuo8k4XEv0
xttOKuqD2Uywa07ATtjs1Agnnc+rLAtu/ImJU1YCjoKQHFJZ0ONOzBy8K5pOMg8CsSWK3vyk2oPf
TmszIQEyb/qnt9WhqSdJ1u0/F4JPE/Eudsys4XOlPwYkTwA9GQCfasUCaA69lu4i5keWeKobC2Q1
v7Izvyyknjjgj3X3IKXcC82BPTk3wazpi5/2GuyAenGNUg4jXp8nOXpQCosepreIWOHUGnfIssFU
CRZl6XDEDGFBBPHHrqT3VH9YYO4+uGHzrOl9V5V07oq7UUF9rznytn2hP4leYCAGyK129xGM6g9/
G/NmXdhzufjQ1z4Zb43jcPeqX3j2BG3OMYaCKvF0lbZfMU1yVsDevJAQprB5m2Ee7P3Pl/eMAUT3
HID6PWNwA1felShEj+LDVy9uc45P5TExdt2z8AtvmDKMPuR6hN5kHhzUXdXeGY3HusNQP5QGKH1S
CdbV4fvMq+09UTnjhwIkdCAplu5q4EOgjbJD5KtU4dqdQXdPRotaSMj/ry3p3UQ2Npusw/SK9B/x
zP6YVk9/NglfrJ/2JrpbO7J8YyYX+wVxjnLFdjvFP9wcSNvlK8s/NZmHlApkmgixPDAK0Dm+rowr
Cl87AqpDUzyAwe1bhWdWoEldsYy8bnwge4zNw7KbcEpkSPBYIC3QsvdNSFdjegsS/CLIF+OGa624
R4rL9AXiHqatD6FCxQweDgPpcgyGa5pSGlzzq4gGyGV7B0OvhWyidcwPH4ovFc2za+0bOBIoWToy
D5q25D/JsolIOnv6w3v9Th1SaUuxxP/vwDw4jeK7hM9+AlfTgaQu9pefylPLFZMQQU/OrF0cOiUF
7O0Y6UoeROIhCCGyuGuqFOiSRsxixpVSnSO+n4gCoMTMb6a0hiLD/DDOix6K+vwASdIDwZHxjAvU
8zKshwGyJ35KJvarDTwtW2NDp+/y/seEgoNl+yb2jdZgov5mu9843KhVQtOPqFvaB30Ksxq3OVzF
OfHCEBEyd8Y7NZyv80Xvfn1ls30dBOwWBl3Tug+cwB1HLnS2iQjm7qjZpS2F1cfTKdYI/uljdk1w
F0spDnaCSOz3AqEBt4qMzwqnprs3JmB6lcZsYM0Azh9dpwcm7hVVYZQ+GIooZWJC/Zq+m6l51nN7
Zz/czfOMaZBDunGbho8s+Lw9da/pCw51fjPvVkWaKtD7H9Y/JP3wyOs/Tmd79wLcVFlTrXcdZnd5
+nNFhOh0PG/ShLmmFUMGDdoh0AEtIaHvdiGJWa+AndklY75jS5ZiJuivGtpGzjebXv/mO9AQZ1P9
A1wM4HIEmbko0QRHC/fmXBD51ViOVXD6XujqEQy7G5zPNguNaKu3DkRe7gzh8nMU2vW7FrWk0zVw
JoAKK0hgN+UPjz8vvDR+TOeMmniwPnE8IxcMMJ0bJBZAwoGAWF6udnA+1+CIUFphmPgzia1D7WYo
D3LDqW/xfVr8ZOU6UA+f0cwsMZsiGH3AR6aEC5hYZJ+xAHeAb+quvqhGIhY6uAO2fgFg0g3OyMCt
EPcdKGFLFDvT6au27z0VCE98MuY/fFUPUB0xUwU4dSJ7ktESoQMgJ264Ig0UIy9T3oeLsSd0Uw2z
M4CUvTLJC0JTPJw8pQTfcJL5NQbR3N3nDFy1vgYR8RL3VCuqVwCbU7AizSlVeRrB+CZMBob0NLsE
S7ThgpCLxu+n/EEsvqpuvcpVmb/8PxrUI+ipLAVvIHEMixVnxc4aOVWJJUMwWMBbrpwaV1vNbykO
es6WONn2pdaPnCsYwPE8OSFca+UY+Zb5Sj1MecsDiXgxVjzE+vKLqJPkaTRWZBfc07+vqZ0YAh2l
Lo0fYBrY4f7mmOQ5ZgAAdiTBZGreqCoJdymAviXNRRspuxa6czdPFKNiTNJPcNQKlo9vV9GmZU/I
hHbKiYOPnbok0U/M/Me9ooKpKXFNjnW2G3Rz79a6UrJH7sTwNu5+SXJLxakhPfz+/CBOeXBVAddu
qLoq++fedecQgfskiDAAX27+oZ8QnyO7DhrX/r0GAk6AM251KoNen8JSJ6GCHEafgkhyB+AbpBaz
MwsCxu+RUTnNk8eqtITl5CVjrBMWz8tN+U8fZfIk4mzGPK2mPPX4057MJ8c+Q+4P8TjQgjfYr4V9
YYcoCepUr3IQPw6lg/mTZvPk/M4IvGI4uF4mMazgf+LwqT0ifTWTcSL/3E5L6/l8wr5YjgZ0PMAq
URuIBIcFfXFilmr+t9tepdBiKdpxYDlTOL92crv4PLb8FoXN/CSp8nIpWUrUYOOVkVolkE39ZumH
QyWhyY7jnOY4FVREOm6L4hmmCzyiqvg4D4C7CY4evnsWJ0TD6X2ZVfn38iR0SKCHvW1vJkXefj4B
6DZRrOnUTRvTHncB0HmyXLr4bzSiBGmiHVCorfdbObv7H4ZSYCkBYGlltLJa+ggrP91lEIEr4c7M
x40GIFQWXBP0YEtEmxG7OD8Ic+08TmYVdoTFvPPHNm/x6lPIPMUqROw4DhvDoj3DnK81X3ONF5Sv
d6N8/nnVcS1fsm/klCyMCXXwRmNEXHqUdAPz1EkQOnMzVMugVkDZMFJzmMRl5hDeZ+yPxuPh+6ix
vImdlZn8XTIBKAV/LHnMyskpYnki5oveVouQz86GmKkojwoV0r5YxIbRoKLQzmvdcf2CU+8rGmCQ
kS8k4Kul2mG345Y+SDafi1hrBn/BG7zRAaogqMoxFdvQi99lMj+WTyauafwHecthHJPLJh6CJFP+
AV/4W+K2MihkVRLfxZVdQhBiIZ/ni6V8Eh0R9hs+83JtmfM/1ZNg+RDl4jKn9c9j3zdOtQlPUi/T
IFLovKWEovbtaCxw2Rt/fkFHLiN871np6JIGqOKq6kRiFYONIaAfgX/ujE4ZKcnoZ3iCtA/dHdxK
S0qKqSJ2gF1BpzBgsF6HTG1aRPIW7TpMumS7jJ+NgvJQKRmer76ayDTmBqwCxJU9U1uk7hYY9/S8
mjXP0DUSik7AZnzaiolfurev7CVbTQZLV4R920rc3bZ7DvAyCnj3B//rLXfPmhVjECuihXt4bUkl
P+9bbiqLJwgkCH3kRaQuaPvT1ZPZpc5kf1N61tJIccEMLJ0VGj3X9uTTsOwCrdJXDPnyWNbz4k51
dmkrbloJ0cl08yfFdpWnFazfQ0ZTae0sExaK1r04HLUw+Deo7WDh3i636Kg8iAqQCUjvqTRY5gzB
rPZyDsf85+WBgEumQSv1iWynPWQiW2Lr9n9u/dsmSPjnjfw9aEwhfYkY7jEOaz/5Hk/2IpzjTMes
1jlAsUxx3qcwqK3eTZ+ZnhAcjNGGONYbP9r4LmfMq21228i35aSP7csWHwuGDZLhUTucDbOCLnEo
NogAd9nSaP9ZlHcCO3JWYYyeo9Fvz9CRFJvirwVd7UbmdNKDhm/5ujcuHo9B66U/Cj3QgaOiLpex
GGDtAKDRneJLoAIbQ7sgyq6xfu7qdX9iA9JLRG/x4As5vZU6sDFZO67y6M2tK8UeqUuGjNLlbdkt
HRPULb0VwvohpEPD6lmDVbVVdXsCmzOF81qB5Xx1xqW9hpaJP4NFgQYQ19ASVT7ccE5thTGlTj5u
HKgEPewSVgx+b0NJ//htX0n/0w+ibW72LwTl4kdZn0vsMg3t3GPl6wDm1dptarErarczmoNQm9Xi
yGC2QdypkYUi4ljNAVjNstsNGokWasl3QILiBs4vgHDMfys06xOiIrx/Z3IIHhIqJkpJaJNZXXfl
HXBdQFamqQjypkmlgSfZPYfRLwBC0DQVfpCa9/3J/JuX+A2QchG9WigaOYWpdF3oIyIWS4vdzey8
0RdGPtaTpoghVhz8IR3seT1fh+N7wVii+gFq2D4UkswGGcsMU0VKXO6PHhiytprdVtD5DWO5+rrF
URnOqjbYu1VFfVyvF31lwibvjARqm1XBe1Ebg7D0BsCwgLyMf0GCBmDianBeTaMMWgcjQ2plQK2T
H+DaA6vpvB0JD5NS9jQnQUt4b5wMoWWwNJOcIuhcbU2Fz7hOGrjanykHctv5opr3ou+IVnsXuoAr
EQKeShxR7T67slvnPjoOWjy3UGJzj9HtsZYeAwx4w80kygsKHs5X2hjeqyPy63nFJan8QxXRXmJF
Zotu88IFBIH6/aDJPOevi1G4+43JtdEV159dEH07OSrWkxJSgF/8Tkdz8YlbD9+boAq8lBMIFVv7
H6MTR4eJyC9AGAjkQY//y5JKzpk97oBYs8eQouiQC6eh5m1SY2H+sWo59ZrtqNXpWuZ54BYh5OoU
0Nlq8Nfpq6OwMljOICrxxdmyvKQKEi0i1gOXWMUh7oMI5cIYPPRgWSr3+Sx28geqLqqWylJf7fMH
HF3fI/S2gcM8dCHanmErdIfRV/qm3oTgmbK2EO3f54YBxzq8Tl5sykpzsdK4EJWHMQsEm4qR03AC
tuGiNYQ/dSbSrPCh0hFZY1Lct1TicWnbM4/wJr/1iHutaGNMJOmmCqQA1Il4ABvGQf7BTMyOo9aT
nMqoaw1zBLo0qJtmW6/FXPHNRKRqpZ3lVQItuvS7AQj9cpNZQCwBBJ52mYQk+9tw1y7akBwByP3v
mASu+RM8UXeh8L4pXhHX3BZanBktLVcr0vFlVYY8mzeuHCw7I4qgDzCE1fDbVDNkUQlWhtPXXGQ+
4ZV+X8QTYm5h6mx53B5i7dHZ3mMHKwrcVSIiK+kyZAuBp3UwW51Y9tV0m6QSnb+j2eMTxygR6Osv
lizP7nA7vHAWjIyoABnI3Db3QI/z2u3wM5zYgDzY2tVE6DFUT13u+a9aVBrKu8hnr2QcqCayJRT0
YC4KT40y/KCWnTcdysNvMm09mBXaf9dnkMpQybJfmzpCJ/sQ5ME/8vJYOdsEBRWk2nITptJqXfak
lxo7U4Ekk9lKHblmykGWDgxtV78eeshClsFdI8bcERbe8Y4FLpWTNbtqxraysBXbbbv2WOyibF4U
kP2FhD3VZ/Ifnr7R4nencsijtFJqXFd0+V3IH78VrRIc3ziFqyrmhO6TxbCdl+piKqzCxy+T0bku
j4G+kc5Kj7FxXltqH2sAXwIdxLgCDug9VEG7eSlNuo7O2NJAKtB4MtFvwKYOT2+EeeKOS4wA19OL
a/BxPM+shSO/Pp8lsKOmw1RnK65MrN6x0l2EWAQEcKwI/blcuVe5rH+l0jJDm+hgSXJsJK8ZkJYO
TBXPAqMU2jCY59Ya1CeihcOq6MJHCzvdChtu5QfE5CnohacjXsSQhm63abbCHk9Tqsp/ZaZcLGaB
LYV5vIXakT9g8E83wXhlXiaCBbxPXZXim0EgDUmd8btU//7qczArKR4eDVogBPZ5oIRMCRUqUCJI
PG+y0dMLm7RYi7tzBOuwTWBcj7Qfkq4qQmcil5FsLajaGnkvX+3gIGcxNw7TC8hEozuG5KbD2/4W
H3stqLYffPlwHAfJlDKwcCh3bQ3dlzrd1veDoJCu9AJWaVbDYtxq6x5BEigmuOGCiWVCSKeP5cAQ
Ja/Auu8PKQ93LstFRlv9gpJMrxaqYixhgL+wJVM6FEZAPPkMQZympTaUWYnmp99iVHaUJUNxROod
a9DZLXQPKGAXO08M3wAsfxzz/Wqdrv0uiLfyeubHnbppoei6TxxhchvSHUxXLPsKpMZ817+BDuun
n1wUoX4LyrKqYFUZIq10CAIkmdoFUdNtQW+uBJvKUOX3xa/esR5O1bdzLiJLDgtJe07Qi0gjOXcs
jEPI+NmT+Y7FMqqCcTELanL4QuuRgUvTjzogwZ9GxCTtSgsaKAev7GwkMVdGYUG0MpYFVAl+h9mj
Ai+8k+UEH73xzV6GusKt5Dh6aylKHa0UcLA6R3Zo/VpNRSq4gaO+eoXP/Pxqu6DtmD5AoSAvxovH
oyRLBxdmbve3jReqFlg3KBXuvhFKfvUzdQHXEvnF5hxjywRSbcVzugE47y8xdWIKIFepsQoJ1spY
VwnJS+siL7Be554qaIAFdKZE2vD3F6C4Ll9w12ZITdCDxk0NlRrOAUB89iTtrSx/sDzXNoBSs7Rr
zPsMyUwp3L9XvwEzH5lemOeiK7PZ8qlCeRZSx8SHBfnFtBf2y5dW2Arc5dWDFP0woEWO1EUbqzw3
do/N5cf2e/1WWc+mvL25G+twbSBXZxIaKMgu33+LY1lH5a0Dx0mB/Ottz1WHgToI4Ek7+v1RYe7w
g5sJGyjZ3ITyG7UJr07qw1xKYGMwVCxTeQszoJB2fPaRbw5qFf6dHaNABZr9h+TSspCghwzWPMvD
6SP8ht0uHc5P6o+iEtc6OqYM1n6GowCkS5rBnbqPi0EQt4H+qPTiPD4SSaPQMv1JlTJVlU0aEc2t
KFftoEC3kiQd8PW1FGTpBHcKuvHeTrNf6hmDdIugNr83JdEsmjSLpZ7kCq3c5rPfvcdL+s4XTQ1Z
lHIt/UQ1IkE4jlvFDaU3wm3oxcm51ZCec+KHJtGF3p5S9wfebqsQjIeC5jjugbSnsxMprIHLESkP
WxWTUeiwkdHKQVDeMRHtHgg2HulycgiFzf1/9c/q0xPf5XluW+P7C34HqQGESEE7vDwSl2OKJOe3
OrQm1oIMbyZwHbNyChXa8nElObVUldlISOevlSYe72UZfnST8JxpvXiJrqOx6Nq/zI5B/UmVlqj6
6ygNDLrtIVkoer951P23sgwsf1UliBdNTvuZ9P61b5emHMHwuD7L3eGdIE54NQh4EGyIXfgST7BN
7s+m3P5yDEjh/JISUpMTGMsDldOMpvMlmWuLkBdzTO9DjTVlgCSSPpcZ4UEigEtwoXKiYdAkGmVj
8BekceFRuPX0uJQ4Y26Hyo7QU2/E7rbqsrmwLWf3bXFgJIIYcqBH3pTXyvNghkcUD1DHzXuJxlNR
I5y2wno66ILYK+LB7vNRSCYG+L9y1IMYJ5hw55FqtHcASh7AQNYLbKdr6Cg+t0ZET6mItQTLvIf9
z/eQiYO/Yx1Y2WE6+aTITWAshGb5ipNRPy6mMcAitlhZr93OFFkwM7G7OpYqmYrHJYw400Pm6BrV
D+C4Az5do5muS+sXwF5pkJuTR70aPEKrltrzxuJ3SJkb2U9GMhYm9tO5fD45qITUAULGqcwF01hj
xQ71PNxrJCUXL/rDVtY2KKBj7/xn7ryP2U16vnBo9DSDMtoboD0rEck5BQfS5hpwrdho7ZpZBFwz
XcE83IOcm1gZe5i2u5MlwVR4PfqLSiyfP35VpacpRBb/OjsPOJggxdLdfYR4h04/4UqQmIca0sjN
WsxLM62fZrux9+lSoeKVd0QkWYw/YNyEYGVkQa19OS6KDF4f4s6UYCZmy7my2QmHtSyw/Z8vYY/L
IlP5vnKbrRGuu/YBTecreO9V7/NiWWK/miWe4dLPZMssnOsVw2gXbKa8FOJrnRnll5puYcXdKa+H
nKaMiOu6d+kW1O7AbzyrJL4oJ+nWz7VwIOHTdrw34rWxeAtAgllrsle3jzmGFdS1HVWZKILs7LG4
zOO3k4Vc9ykRvPrmVzSiRVdax+mM69JlaDqzXH0E+K7e2K1PSCe1Unlpszuaa0Ie4Se8rUAqrxf0
p3x+51e/9r5tkQkRW2z8B/jWP4xaNMJ8cGZud+Q4Uot9LoNKzRPtxZrzEXOfS+NxOhhhpNFfgHFt
TWk8NZWlIqlPHGmNdDaLKutkiocjDvnyep9JVImhYTLeaRJxR7Uuc949E+9PHM+71yujfeACDKjV
gk2EgZ24dEPgzK3JQ6uujp5jygQV+UmcmEBfavW8jQF+f6byYqMAoTZbDNmBpr+jd1ZOTkYF32gl
HkND15EsS2JL5jB1ZmFLYEXG4x/iZ4qzpT5stuoT+CwSoRkLbQ/0omV4/JiHfXsAQl5JFAEbKCj8
fk0QL/+Jxk1td8FyL5s21JW4LBYyQ3jGu4n698EVju5Yjt3cZ6znXhCYF0gcpnT7nwCABwyLIR+L
Me9GYvw1xIA7THDHY87KbjbI2rktKC/pDeKJXsvR1mPW5xC1tHcqMWCG74TrBldSHW2rLohUp3zw
BsJpdN/nTz9rzgCF3z0DG6/5SQ+LfvsLfIF7zxbHUKOjR4++wDasL498InSXiJKH+YOTuLpe/Ms9
SNfMXVZ/FhcEBLFr592Kqr/AjuaflUaZyFpSu2MDVPbvUnB0WPOKx5v393hNhbznCMgQr0q3sW4v
9M7fuTrDbbSr64ruxvCDEKeXcCliUShiTTUd4GpFzPgyknG5Dt9w7sUYQ0NzBmkAspwsHmEGAMj1
zIgJPDc9Fe9ODtxiicekhafxplYicRPzY7ATdCy6JUWJewnWE3310abvLQMce2jVCKgTynUQr58x
7+OsUHPLAq9+fC+PTOPeHsAT1MTPMX57dtsG+iuN+aytvT0ednDlHNxBh+fYksYQCAShtnAvcbqv
j+5yDTXVracfTLYvLn4sxzjy4l99R8JX1JpHKTL4rVA5EmmEVm/2lAD6fuEV8rADx3lgxaohaZ1P
Owt+MYVPMpdYXpieqbq5HN61VzANee1XjTD+4JIh02amCpUdjGlBkbf0Eqw0KRE/hfPb/JQ2EUuo
+wYHEiFrihSnwops57jcYeUxuC9i1G7Mcfbljr/qlI9rg+xGxVS4v4/qsBJUNYD/OeG5eeE7aX1h
CkY9Z6Bk+FNhy6HCPWmMWpKXC8PrfOKefUrYwtptW3rkNzogAYVFGj093DebAeyCUvf6W6+D+L5M
gCX4K6EfQzYMLzwlLIOWZNf22KFghVrH2eTCctSoO45FWEWDqYOdre0c/6HYjnKGz+SpVeRjFXi7
l56twPZz72YRoR1ujIOLSUcm7tWvprmyM5Jz3yUB3ntw50FJq3lO26ewx2mfoy4iAhedVWcy0uc6
Fp5hT4U8pzv7X6fcghVgtRKUi/wYWaAhAifhQe1tgP4H0Kk2AWw6vbjQ4ShB1sbBg0Hx33SzxaYW
pAkGp2SUtB7UnTifJXYxSdWBOC7bpuFLGTSyEZrs2CYnGEIP/S/OpOG78flSJZ6ugpXPjPE24D6I
nrkXTMFP1V0ECNtMl/zvgaeofsf+UhI1erfaWhjVoRr+EB04klF/7HlzmyNYx5k/3vs++V6C8udu
y0ldUS7Xf6854/Hbchnr5Ait7AHi0wpHL4BYP+zEflGphtkLM32oZc51dbQ7ZnvUITN0PERU2UdH
kHIXCYniOmlrk+XuJLDjTtsLOW1dNOSF+3gfRjoEWvSqfYIPsMzTnbuuM4fm4d4eLS0gDD3s/hB/
w8ultLDjVdQIBrWvahoBaQmubvsiUDgcPqFDlZwKOndpvNu3NydnDKYr32X1MJAYb++W4e8fic1b
mLIBtF37qCRKsqF/1NPpULaxqgp2TBiZInRErj8ISf7I4wG9PNKbVIcbzqSoJZwGJtZb7y0YrkBQ
iN5/hLKWAXRMXvRnKuh8icQVbkFOdCC8R1Y9TIuKnYUqiCTQIfRz1FeYRhGIkCNb7m0lTnUnE57L
lA+SGZbnI85SVN2xqtAsvMDGLcjYvk/ALSFXBpav3eirgtd5UOwC1x9lqS22RIW7Zv1V7epS98Gc
YSqBRUFU1XUjEOaYaMypvKZyP6eqrdN5VyI2Le9QKKVHaQwYsQLHibDEL+MBxZpE4Qr+wSipJ+gq
3EfGidke2WhfCXouHU58EWzG7khXfAXRCbodu2+yYWnPl52KDNlcxhVlowzSIDXHRmoB360my7A0
G/XY7Gs9wv3ZIGojBIn+5AMeRsqSbIDdlHPkYsWU/SRmQo6QFGGMUwRzwU0OZk1pTCsFVNhzBaOq
on+kavku78huuBNwK3YCF7CiIWwoy5mBKlqFq7KP0lreCDptr7ThwV8KoOF4LYxZO1KTKGqOAhjn
zu2oi+Bn5dSl67p2qFFxzMVEQwAjQQMfRWyYrdFqVBaoOgly3YAv26EJDh4637Kb064yFaC1n5kb
CczNcqDldMOzth/0VaP+OgOA3aZqTAHtYcEibMyzEFaXrIMvHDrzXYetjPTRWWXBJuNMoHm3V95L
Yb1ZLszQg41j8/74zaMVTQVpJlRtdZUS8mKoj1O1YthXPY7hBVfhp1gFZAyZTkrGOZc6TvKh+xay
QI6bbRsHgQz1Q1xrWlKn9EquBIHXdmanhZKYi4Qvo/s8uScfR+Dx0HEwIco8Ff+YmMxyeMB6+z0r
YpSocGIx1+J38JfFFqbeR5v/LReA6l1oAIgukAczlmWWe/AlMDnOx2+3UxJ/N4TWVArxRHr3c8CF
vHwr7WnjRhCwDMetYZVttRo0xl1j1SGnaoGIIn6WGKjcp7Nlkty8BRRmJhSnkUZ/hci051dlPF1P
Jv9XUNDElDIXBsWb/C0fJW2jeI0K2NpNUTTKa2ujVo9XznX1887e1Z43sy5OlD/q9IjLnHQT1nMi
Yc8NJrWl5QGg6MboBkjHcjIGfLdFlh8RG0ZOY12EJbA2/3GS1EiBrWCY5l3ra5+tZUU17oDXGBi1
OjH5vqIU89BmrtbE0ghuLQ6m0wql+AhWWUZJCIz3jUw8biC7BwJ0X/Ckg20khxUW6JBkyRHgqHTN
BzTv469/1LIS0OlgwxFJim58eY0vl8ssoqLm3ODHMaNvjZyokYVYAWrLAhSemQw1Rar67i0eLdZg
i2lHOjArNhZZsBN4FUXyPRPjPzdKlJecNyMJ5dlm+0XqWofe+vro4C7DNlgimaIHDQzTfq/VouDE
wJnUdwKBEC0C584on2TFVVYME7lXs7gboP6jxgFbYeHfjLovrGBnVf8V4k8m64sqmZXUHDtRgJSR
wU80SYV7lxeGb2awhi89qpXflKwpWzQbbMqjF8M4rDnFLn2jgR5k6TnHFF1rqL6Mh2DR/Ciwqc3u
nTT/OmkycBCMAf+SAsxObkE/5wwOJmb/wD4AWt45rbFt5XcluezMjYf6X8Ddmcc6BExe/3ehGAPQ
i4ke3orDV1CGFCtwu8bnMHHafZi8890YwmUbCsBIFijiioXHCaYvCmO1fqANQmb5X2m5sp5rV7HG
HKqGE8k6g37sHL8OzVLtFWabpKyPRerqf2v5K5DH/rHBKnNIan+opCMppUgIuSKbOJ85IUSLOM8v
UnuLTqXa8dWqF1CWhxTTdgWo2t8F5y6hwOLkdxBS7V6/UaEIkuOSEkzNYdrwSQoyr9qJBk96Vgnd
H4FMV+UGCgXisMcesWEIwSP188SVYOH4UvgIdt97siKAPd5T3i6HFDsY6X0uxux7P1F2clmJmhDB
PoBlLIxHes5htZLVPBi2QaBZyx9tFwl1BBmwca708cpK/axgovgLWT8Fj+I7oE7B3h9ydN3wX/Xf
eyKHdoWg4rlYrllvKhpGNrE7BWOC6dVmbQ2N4EWNoOKzFbX/dj7XfN1sQBrXW2Sq47Ybn+ok3CwJ
JtSsQdJ4hlidv1AsnaGj/X6EC3E+qeLx5BFK6KkmUStKEZqZHe+LszYTWWhDZFJ8nZJdGhGUtfQV
c3UvvFhnXC0OiTstcyfWNzwKqwJBNFuH+xB/89eHimfJi+SbNXXv/OhPJ1TmyCxcF9IDcaVSfDFy
4yVdHhh+Txv+yZz5Y7aSIBd4NjSuLCNrak/g6YzhkmJusRnJxo8j42JJqj9oyUYEMYpcvwsglvZN
W4sO5GGvODoAO12YxCspcqcW6wUh1Lly15+Ln+zZyhLnKz8lj5YKJAeu2JcyaKX1w3xjXIdGVv6F
yvZHHLA2VKpmrM5mD/Zk2Cw8BdRzNEk3OK0ddolVgPQZERkXWRQsXvy/p5shT1OgSrRdlG0mBQvH
AgTD+0FfmNmFs/a6vxojL0SnoGjnE6gpfqepaLBqockGBNNd0jzk6viBSbwJXLLRRnGZ3Q8e9XjI
5WUqg7skEbJ9CF9LqPbiLAvGkzIk+Mg8CT001QMeTLAplj/kVRVEuO4TQHy1zuCL0R4SjPdk2nS3
o066jr/SjBcIOpFEvmTNIMeqihYmvGRVrL3rcMKWMWfVRFoELGy1pPn+f90e++M7DCWzNCwJrSzv
TRtg0nvwDUSGdYCzYXk4SuB+gWXN2wjfBd9d6qcaJaI/g1Qi4Njafi8meE9EQGHSRqUS14TOeL/3
j6AX8tNTBogVQuTdhKYxwdMOpLnSlEwejo2cACfa8/2yY3yqK6kCgBAfP0hrkIJ8/P/ZVZmxcJUK
K32bAK/J/4g0RxhcRn1xYG9e6kJ27gTZzIfSyWVxzU/kIOu21vXwS+HPLRxK3txXtNzS7sjxn8Bd
m/eh2Ln5XpO4cylH7OairnoyJ9JWSv1HZAwZ1mBoiP0aMlkBUY+YuWXfUG/SpTNYnbcbeh4MxDgj
l8wncE+VfRlwug5hwLDSuBiKU06r1RMCdIIuOVO/ILyYCTrG7HGnB1gComYTZgXNbOQo+4Tl46ht
PUtlRB/bkpVcpXqbhxF/RLxRr1l28HEHL9B041O46V9ve6lutOZYmjPl2oZ+S/XBnmVGjOUrAcFs
FsD9vWe3Q2lyKTLw9jIhXQE2Sl1JEqIAGp9rArkub9WHgY03uVWOEL8yZGmQd/Aw2CwJr5ZwpZbI
H1CrLZxZSy5DFfnoJ/1D3Am6XxsDiXutRl1U7t/yst9s/sKew/ikPfaHkJN//Or8gOaVoANwYjGn
VneHl6eFdKT393NyrO3oHLNpOEwDawFPiTIeHTLXiz++sVRA1RoDZHf3ULIjHdSl3rPNU8fwCivY
Ajn+T4aElRfcUuZoSlSldkoeVqAp8gk0mrbC1gaVM/JxErWYXgeDjgNXNR+ciQxHUMcU72wlCa8+
j4HkYJIox3+2FBKCTNoKRrq5KSdG71EhFcdoVJF/vnUnNqWPuKXQNtQogA5KnWiEtNfGX907uceB
5mKuo8UHCOYXwi1MKy7+Y1IWqeqD+4+nQ6DWL+BhROpglr1D22pxMNjwneHanb+HarHAiYZtU3rZ
BpC9B/wLcKx5abiRhX676A6buJpWX0fKRj/7CO45+ADEQZ3bONUqnUxeI2Kdl3UueTaqo2b3C3Sf
9PomH8cs0O/tuIwcSwkTOgB3sfVcHFNor4RJzz7ivW7U6RBU9FcEpJ7bdeqX/gTakCfZLkAEnrcc
DoU1jl1RSq+Ky1s44ONivnaMmxF0RnmkYX/bB5bQPruwf6cc28dYo5zJ1RpBlITbu3PGmUhp8Fyu
QZsz5fe2nUHNb6IxyacEyrXg8yiamGVWVJAAlfcI3KhxAPDTCkqUu8l4ClLKGecGsNEJWfKbhxpB
sOD0kYkYo77bPbgVgpZL6mWnFIhPGaQr48t9/+3DpUw7tZLKtxnAGAViUum3bxArXgfZlCiqphmZ
TKqscsGHsHha7jL64GEGGIrM7/qMnwmE9QzLOXuROfGBp4hZ5cbVgIFNSH8fyQo36hFBneNpIi5S
ONa1ek2LJPTkpUv11/43p17EDf3rEh/fGpEvSdEBkrefhx3ZFh4ihRR4jAHgWv9fQdcv1s5BQ+9V
C6dA2L0CZHCynkcr8hjQdRQseFdOklkdOhLDmnFoauzBqGkXkoWFINIJ2DKvrALekEwFw5csD/cT
7Haw2aBvnKSu4Yl8GC8SGZRG0SDCCjpmVOw0ankitj4+QqEH0RWHN0JpPaYWZuoHamYPR9tngsJx
/LxpQ5K8XlRjam3+cEUn91KFA/cHlML9OLEz6Fh8C3sKF1vZUpQESHT51YOo/urPEmaBL1q+BnE1
iyXXg+uybPijEja/s4PD8KEyNEEeqGVUiHoIto1bFjndMG08q4sPCb8HGlPqCKk4fBhIWX7u+H4M
mdsMdgnrn970M1RwALJPfPqKOxwKZGknwer6Uvhw/PonEOs0SclZGpTKbO0EXEpp2nzY7Adi/8HN
mLeHX6GnGECbMfZOdBnpMsqW2tEvmju+gCsxP0qpJWxzRpdROB6p7NONs4ZbNjrCboxwwYkSQIRU
Ar8JC0SgNCIPM3UNGg+YGE3kiDSpdvsuwQgf2X5YCjYOp+YeD7qN6Tv5rsVcRdyzwAiWUvDygSN8
ye7OAUiAHV8mofDnliCYgi4Q8EYX0/R8Kyt5Ao6T+pq0jKQ+qdHdqN4oYLtf7eR1ZEwQIhXqmpIQ
hm9XYloDz6+YoaWwqhPfvZflRDF73OlKbwQRrUNmc7mVF4EYiuM1aMffOV3HDDGd7OcDc6SZkmib
aYEXMUvto3TcWH+roiRcG/B7qF1kg3NtYMwgRwMsvpk4esdvJbG7Og/YKRVsL9//TsqC+5wsnKOK
xfFYmM6iLerce6VmmhlqiZwger99Mavp0/AgUzD5FM1oLUFYdyIqNMlMwsUDcIP1AisYBsQwqegb
+nUG06uhKtdPI+slKOYAkQZQe9PUu6l8MQjrhXGDiQ+PjgkOS+7C7UTKtq+rDSo5PxwUXmEP7ENE
1XS9au5s9QQVWJShocgbJUYh4fnIDkN1koQlbGTT4X5Fpnpwg+LUvQnmjbwlmIR2iOhhSG7LkX9H
peaSSIb+r7BX5O2qPbN//dFy+DLmwH35/XwgnXmpyM7naUxCMk5SKYESBokQ7t3s2LxAKWxTRGVc
iZJ4xAFy58bugqWuFWxBBZL1sjaT/AaJHrfLYN8+je8+F1AcfcOSmvl8Y/rzck5hAKLMLFL37uIH
zdYu85Ude6JOf89uu35jEpoV8WM6x7QgkvJshmhbWtYBtsizdqwB7z0hH/kAy6Fg7W4LEIJmLdK3
iytPW9+iRGmqjFiim588/oYvDDCD3yWzsQ8g6UnMz8+39ObCK65hwiLwknYMP0qWfzhkJti3rIDw
GFvdm+nht7fkwKfh3ObF4A9nVM6ffnCr+RWNT9m8gYhYONzBtTmL2va+JcJrnuwma64Au97JjaLF
+2QA8hHRY+ZOcvBrVlEoSZHY2ASLxEiJT6A4ktLi49UeNlUeq9mtgFYUHeKWqtmX/tc0+sUHp9pq
u0/svwOH5J8mIelaVIceSph4F1QGudvwsM4ap7PpXwJI5o7O6+nu8bNMjVUbdcfu7Gs4rtB11GVr
/LjQW1Cv7MqAEuVp/VTKH/oFmoFcXNvZMUviygDmCSNVA1JPbPnG4UH8Zh9LDScJ6ooBZ8OkMbRh
D1d3OuVI3psHBpYCGXogKkivI8DNoJXgIIKXSS4NmvbskxzJLgOR3v3dGdrkWnDRIjAOzy0hoPCz
UwofVwVzEY3hm9REJYoU8MPQmYv81rX11zw2XVUGWPThnmkRf/AZvL+60f6LdvRJA0EmjxKiimH9
kO77Drr14BSSewRf/ErkFv4awm4La3fyXxW8MFXA2lBwZ2uwHfPSB+kZQlNn4HfTFt/vCU67yulz
EOj6yDdKnfV2eNKTqMVz51X1XOuGXnZuPiUaCDZRymsPN2yCcJ6ycu7XaW4VPuRGrTiy7ooYMkLf
XK2I1aiM/skTWpf68ce9054QHpo2MlxfMGtfLagNV9m8ytezIc6zDzmrptmkX/evTKcFCpgVcF5U
6/TUzXJ/T0DqpruAMx4sjiMXQ4Y8lOZ1nNt4grk3rQD79YXG5/Fan8Bqa7IHuc95YIM0jBgGHe0a
IubCZHyVsVoxlr8+nqMjbmxJM7Id1fwgvIp8ww1QsaD95V02KcthfwDA+CrjrZ1HAGfomXuocpvK
XIsn4Dou2FGxZwPJ5VNW0LrQnhQk8jBIRc9wbDndmarJMMP33YDugV7i0P197ZJMR2AyybAD9ReT
OxvZ4rguY7OW215JBBHn9qUN7isiAc+0BlzOoKd9bwL+7hkN9cu8/0z0CoUVkxYrRbITsaN54xpV
VRAPKNjgFvBuUmQ9y+k6w0v2UZA9GQ8EJFeeFvvJhKBjiPAQqoXSBd/SS0fCqDSAb8TdCCqTF9FU
X7jXWOj2YJMMMFTfRQgEhylnFoSgnYZ4Huu9dSg36kn5frbsJRB694Jcsq7Sm2vxJyDE8eK52vW1
S2RcZK043iWy8AFj0YVYa/iJRgdP/NGmoxgBjkfFDVxkcn/mkYUUVnzZ1K4zLAw+ucxpL/wSnXGi
1m0mRDx/MsrVEU9+Ay7ngqOAMFrIQbuiNurpJQ0kFZuEoYfU8QHiHOLcX5F1Pr/xovQvWLBzo44/
AzoUYh2VsDNRBvzWAtdjlFhHE4OdpFQc0YNjKk+Ip8++cJ8gtLqEzmjFOZ14/ql3dccsIVX2BY2J
YBlZIHVx3xdY2Qkw59ypyNqVq5SqKdEEUIgOLFbGaZzrOfT12+brvZLtS8zvDXI410FsTwIHkbx2
AltTpaAPEvWpSPtAHEbPzroNO8gE/5Ow+cpWgR22OVAK/IaDyeVoqsd/GRY7URx0vU81W/YRm+y8
g56FV+URx3eN4lxpVPhS47lUkkj80b3RPhyC2U2NyE6Qj6NtiJTOiuK3xwt4vD3gCpp/dtnaY+IB
axn6ALbhyVaeDk8U+yfgfqt36+Zoc+aE7eRJ7Wzyqy0XGKuw8XnmG9DcoN6HZFc6hdA7ebR2+rWr
SGNwEPtBeoE3K+FQ8DINXWxr5nEGPkvTZvEDzEzpA7fE1P1WriGPMWz47BpI+1lG6Brs/eEk1OW5
IsWK1gV+CfuNK2CaH5pyF24HnUn7syoGVmGGzWOqbUtfT/d82L0pz3fwWdpAvbD8Vo2Xh7QPPhRR
DGgdQ3laZogr55WYnKoSvKKGQMRTOwiKsqx0OfStWdtDbMf6SWJV7GsMOAaOGCbrz524ZjG84OFH
DpqRnINbi0q6KmNK/Zj8+jPesziLGKg1gxuUaiALZF/VgXnHKQwhCI1VVJ9RIPZ4NCJhXAJdCjgs
cdt4rlOTpU7QLyDaa1PxtibJG3a9Go5QAIZcCKodd34uDxcwdyuVxMojuK/tI3ICglrbOYvrPC2b
2De/7DzOvzTNVY3d+WMftlgjkpvoOuPQQggOj7DcF4EsBoKt19AdggqrPp5BaBb05D+6iIX30Xlc
qIobgPyIGqgTfpUp/looqRQgn++GLLSQZSkhzIpQSDFH9Ev6VKuWbVpZGPLQGcglZR4TnZMUdLjS
rVbaWQt6c3riekeFzxlFCHb/sCVWgmyu2KRU6NvKmcDSfUvmw+q+Kgl2XuCvPYJ9OptdTiBSn6A4
gDoMjEeZAoRfddS9PknhpZqyk/Sa6MZzL/XbCCuRLUZ83WD0TNKEv6hJ8QY6zgI7zN0Al6Tt286E
zknpACHw29huplf0zDtJ4CKbHLythWgrty7BAjEVJOBFHuODoAJ3ps/UWRVYWHtACamFMlCZLiQC
QszdV4JTf37qYrrCZKFZlijyOWlzcbxodpBbezCmpq/FV5aN6GiHOe5PwNv2ukQKogz1atDNTfe3
VdI5ULVjx8iyPNpUOOG39Cq+nDf1NwQuYgqaZ7bgozotovZWFoq43EZ7HmawMFul/9fdRcR9wbO3
SqquGqPbaiGnvSp0HUftlgv0JvvL9iJNOwHSMClyhEIC3mlJYe1SD1rLYdwdmkWKaDmHEiLA81YK
nwsBG8J1y/CTCr7ojkIdJjBzpMQRzcNKJgEDt45e4NLFmPukxkw8DumFYuxifH4OpFS09CuH3FzS
vlJrKSVTADoH+zF6wMKBKMoitXpAvlFtnq9e9+vU8X1c6llSUZfjM6G8atdGx0yyqt16rSJmCXEf
HDLIjhbwjqa91l7S4vbDd+nqJFG7DnjipIn2Kat/+s5wFpvdNzxd7hqaLBx5zjIvDPOGzbji6PMm
KWNETIajrjR50IgGMOZNy2sxnv7IbGPIBGmGf5C5kiQQDyNl0p9w6bsX0QPIUXGtrQ86RTLbO9JE
wBK77zdyvrOla7EUKq6O6XOYf/x/SOgoyuFkOEsPxo1nXN4sGNqvo5tJJn7O5p1tnYG+oriHgU7h
evvNJaAdHBeSMqK9TK2TrUCopf2einL3w4Ar8iBUCZb0ig5tMn7xtf7r0qjCyehdUvPSeisUDmS2
pfKsCUhKLs1AIqReq78JD1kVjG/88wLts5rHix6vxz3fQtkJ0L4SZEE+RoDNMfh5rQW+w8Nr2X1V
06CklXgiI0qWoyr6eeyFKfwU1oDqnD+vlK6ZDtnxUPJzkNSxraSJAQjTHbR3kNsyCPBqscn5ZrIu
wvyb8CC/oimGZv+5gNJdNUNOkXVrg5NxJLGBRBrvn3jrYnaAjVVc35C1QMjJi4UC5JeUOt+VF3qD
Ufx3psUfMb7el+KaUj7t/fhRmM4oBhbVGvnp4wgfAbGdo5HWSgYxF6dg0xJNX9ECFOlm/IQsBmUr
j8J9a7lbyYGi5B09gPrclXLiCTicn/XGn/2pC0x9EOkDyBXDWOmPz++3PHRnOxBV0ChD5AWZkAeL
+WqmGKHuFFH6WBm3gmUqOcXzeAwB3ySu2MhrMV0Idwd5SLPrwOJPQxQasmbkhBKMGX8rJn6TE2JR
8BSYcE+juIQ5PuCuPrwiZDmU2b6Jp1ChpFdTmzdx3tLt9SBA9g4YVpN5i94j5KOEwIiiTn1Hnx+G
aScCn/s7v4kawmfm887g/MN+RvB/EEbbSo18BJe5TbiwYo4yS4Nl7ul+G8YHh5e3mmvK6erdIjo7
NdFlE5KlIkduL4S/AmWCeo9MVpkKJ9ZX8eeAbaaWXQx8Rdr4Wn7v+ivBeXBS0sZdZWKa5hbh+NuW
iH7rqj+VjrJqOHD1NfJI3pW/1Wpxr42fuDfcfIldLloYrcUjpBWlK4XVi727wBoWcq+lcFBA+e+q
IScLUycTColw7XmBMxmHEnjd89yezblvl12TK8nvTgi0AY5D9cRoEtW7yJSMDIC53Qr+DkgcjAqf
IVMIbdxOF24Pt+zvxofhV3QgbUSObzKISUwfovSmnzbkoZee5G9v4CHAdA01H6ovP/liZHXkar0K
veabi14sTvCbHch275hUynVZ30s+UVcyYE40g95+7n1d8NaSQ7vT9Pd7nE0NZRLX5oEMnFCTOt3W
7Knim2TaPSErkW14zHwh81BD/L3CBjYJTjgQ0SXlbd4efozdYe+fW7BhhPFUhXTPw9HlIqGYdlBw
HWkpWfNoumGRQWVPjBDmKESYZZGqp1PhvqTbggnjEK32XzU6OdFEXHdHOOLATrx2oM7qPuzz7r2c
k3aZpkb4VfcJDzLvCs9mpS0HE2kaIESouTZicROuolow4WsThdxeDk+chxKbr74y5FjOWVtif5wJ
nfu1++mVcPrEQKRqaa9pgmuCI06CCEKju9kzs5flU/1aqnZrGkxMdZ7hQKjL6VD6D9FXcw8aSZK4
bg9N4Lihd1vFk2jwrXQJWptGyGsOkicm9rSzwkjuDhzTdiFZ/NMRRiJVa8P+Nc8JNF7Dm8R/wSrm
hU++8VW+vAOYAbiq8B3wemVKHL9Fzn6R+jWqXLUm5dRgslLgcGUavBubDEHNGVhnfpnXFEj+/YpW
EbGTI6baCSoZ7W0t0Oxnbw92VHTQC30MpdsFkrNTrclJodPdeauizYRVcL0KoD78DxM0ng1s+6lg
AIyFdlWgZW8e+jOWxB46AgUZpqTcTziF0koe1UJauqo4d/qXBq7Dv5EWF66o4o0HaDhqFOyHGYd4
SLeqVT4LJA4AY9Zy+kdczrNpLah45BE0pDI5HO4pi+31h1WPmCtN08wDytwZu6xBU4pzXOwNZlNr
POvEwuf4UndzFRBrhg/1vYsorTTqyvMNqJy2k8FzN0JKx7QO2ZB/1D7sQKtFtSMWKQWoYX6ldQrH
WKT1RxxUUmISAzXA/i5HjpIq3MoAzXDjSK6NjSA3lHwPg8fBvY3dripT88Eytprfi6cm1cZfAJ0+
+s8nJtKCQKGoUPFPHwPambg+DHzLVjfWSaN+Gx0lsFrAi6/WY0H1+W64HmTwSllmbURLD5Q/SLm6
h6USgVorS9rp6Frcho7Esvc170URLIDCXm50+YfYh1pCulVH3ytzcQ4JoxJeVPY0skB1h44FvQuQ
KRxn/0sPv0PpR/4mQxAcQvFc4wRV9DbVPNefu7RyRsIQId6OfdXElqgWSNufxFlQgjXvSwO5JdXR
/gA6eWE3aD08jhBQfDM0l00+5TemojpjARiTPKK5ObjYQ0n7dyc7AInd7vRNNHCCG6RL1owYvwDO
z7FTP11Ge9E+khEbThp9Egbv4l2tOy0cs3QdEPHOTjn87kKhhp/bAbBKJPWKVLB3IBAb38bHBG1S
7qwXRvP1YsraJFCGGEIzTrODTlVpLk3CBV3V8uWnFq267AkBju+qjSaYz2ac/ctL9+GsIyt7Tm0v
Eg0YJwDvRcJtfMjfQSyAf/S1L4FeHOF3uC1P1X83MPJB4pGxgmo4I+SkB99nKe8eT5TclWrPvtV3
2a7By/qo5fq7DcVW2yajV5eeXmk+1zx2LIDOSGh9PZBfxcr3AcEzN1z/aO8Iea0e4F/1kB3r4/kO
pBaCGznHJd1N59EIMC0k4+eTaPYBktejIPUpCo8B/AOgaAUezeSt9FtT9BwQWenuqu1DKT2Z5Sie
FNHOcsZQq1S1OnDfSIzHDzXw4vcSrENWo2wgFZf7vbocBViQ+DpghYcNBTGchns6TRxVlr63VciX
urlqy0yprazZP4/iKhCDkMjylfNahGVaLSG/B1bF3LwTFXdQ98KNIPMTOGBg4MxUq4uNTe96iRJh
HZ8nj4LGajY5VwnZwM6c4t7uKfog9RqO1vkp7pkZQxwk5XqqV2EEmZh0819pITRLTVOPqbxP+2JN
VaU/0nqAOPze6gZ3DWUE7zcFQvg3vJYCm1UORzbNB2jiXyb5aEmdAJKxzpvD/WyWFj9WLi8BV45J
94raY7t/amTkMce5aZF1Yc87mEaLOKEvjYHU35+zgORE7/Zv4OcpEHaEOqAeWRgH0ucpe1Qyl/7p
NMQ29irHWfZ1+lKBUTQHwyKGa2QrsLIgjlW6pbFoRYSZJcO1Vj1+DlORsZu0JPKAuEt8mCzjO7HJ
2ZMN3P65XlJMcUY4yAre0khQrwq0tJzjn+T9VxCSl4HupcJ0hI6Vor0CVDgmTFtwqaG9VLdbNHxA
7HpgTHZO3k4nI2S7n2ZH0QiI5NnVTDUer+TjPt8ox5514GITti8qmPzFCeDKaAnvMEede0SgYFPs
fogW4ePdItghLx7Yr2kuHvDtXBwPMNp3QIOO4mU/gqODj7n+VpgDAE1ZX23ryIouy7BI6YwCIaZP
UjWSpdIR5AP35BbwANfkFMVttAd+YzRxmWH0NmFjybf9GdglkTsQJt5XXNjG2SSsxXC8GJLcM+Ys
zNpCEDUA9lpJxq+6GlS3S+Zg0Wypgy3aWvj0j2Rfp/8vsbl40SlnunAM9casnPRKMH9Vp3P5urRh
ZoYFaHBp8tLA50rJM/HQu+/Vl03jhpzOZtCMfhN5Vlv3OWBHp28RzepkG3BWUD4yTyl1VHXlZ+x2
FDrYCd+RGROoz0K/NwLydt9j7VoY602jxkFGwiMyOQKMGPRrR4cl0uNmnXnEF5T6tZyo9w9FK1Py
vVN668mSiQKjnrTO2+Lp1Yrnu9qc47wV5NEGFXwfa8a9AQnlKPymBR6ajCThXwBPr74i55lDWsiO
lZAdlc+RZIs9dX8JW+EX7rBMM2qtJKKlb+t+apE6DmmukQglwOX/Sto9reXfTOdra2QvT4APB5xf
PAAAsrwY4p1BzaFC6j2XaNHn4lAZ9IO6nL8b50DCUAZNJ8l31ynJXYAr4ciMUtJRB4KzloNFMbJ/
yvGUY0WbFKtoz6kJRqUBD1A1gdYsknzI4IEC/6bI5y0SlqR1uYqGcjItBFt2BxqEiCq1oNONGxXH
rcaQKpXJ6CsZfa1Io0fvx/i1vRI8TmQX5qmUJCHLgIDDaQTxR+ySoBkySmNj6DGPw66lFTfHeMgJ
Nwbe0EH6IryYlipXr3leGTkTc/SiLw6m/rAJMIGLjQhOkIg3X05JMxcl/WPJ9MW8G/YDT7O0NcoV
19S8L2EzWuylViIRno3PrI32xNWOcDPbCIKgY83YFIiXQZFfzrzATEtQaNYQljfWo6vKU4/Isd25
+WpD62MdZQVgdmQTB06OPYI72euXJMBsobNiMZJSieXqW7E5qtU5zpYHK8RrSqeaDOga1FnM7MN0
UoRGslZ9E/Xpj7jBJK28YiUJQXlwitwYLMb4piIQBJu5j0PizzyaM7Yww0d/e+cBg6vvntP2kqzv
+DD2+7Vs1ibzJOKOceUqhoqGqaz5twKAxwxOnwx17krrfHHmBXZFGoPp9jVA6+WVGpj1iFLGYlsV
JdirGL2cVF+M7D27YlPyzC/04pExtr8JVvegfC1evPBSSKKyPw7Wo2GlhHW10spwPfu8bDZ8Hm4h
E0OOOM9yILFUdlZoojX9NlK+7C+XQwSDJfc5vFw/xPbMk9zkMx+KdlUk2HhIDA9BV3ACvA70ozlw
W4YC39jieXvHVmnd7HWFLQWw2/AsP13fEolL6anJmFDlQxPeCUy6WUeel8jBoT8WbHaAE27GsbUu
pD/WzfGnd7GiFgZ4qdWNY5tA48FRtsqHjL/XrdDBKanlE3X2NHOMPo67m54iwelhDKnjuuZU9PHk
RX495Kb29Htc0U6nn79B+RvPsTQMtHin4LizyLSfCdtnpIVFSAKJ7Iabvw5vXsEom7h4YKCEUpVu
F3nmqxWW5Ecrkwd2BBmC38SHnKeGtBNchOEoJAQMOh6v2sdZoPWC+93M4Sct+nLgJQcDe6Iz4FC2
FIV+db7AoOQA4ACQ554+QOSukQbMfhjV65ljPWhO8yGWJJBOHxRkWBG1ZxYAJFFA8HGIZOtM56G/
V2c2+pbsoHjuVOQwUIbpqWL/PVjWeXg1pjHdfx4l8t7dQ5whb72M7KTVkkID7o2ayzocib7EoSCy
7BFa3p7rlGAruRKC8h0rRefUoeg2ktAr+kI05sA/3e/QnyXMvfXnl+PKUoeR3Iu+Vu899wvjA8h2
gZQTv/O9HNKDxGv6zWluEzBLhFlKdx0JQp2fu9ZJHNVD6RXgGbPV1UK3V1bByj90EBYCnS6aHRRG
h3A4mhr7c54ZadEfV0FfKyaJvWEcrKQU/Pln7v9rSnzvjYsaDJJUoq4KJsOf0gnzmbvXkRrwWCcP
6hKMYPc4ZloU1ihs6OLUgo5Rb6x7dzM5B8nr2vqh+ZYCOk8c//ukO0qvU/SWlqeg5nZ0WbyBln2m
VVP7aofEcHVLSHxcwZvyIGL3OfIAgwrXdzvuP9XMnLxs06UJONLnE0LgSOeq4fNAfal71h+8Gvhw
iT89wTPwqfkZLMxmG7yelf2Nv7ff0NCr8lFR4zLr4ZFZB+BynjvOj8VNglpLWKMLrhVMsh4wZS7k
frUYcq5PiGaBrBBkXUS0aMRDixBOB5z5W55KAdLChygmhGZSVIBX5FS/ZnlDLEYgV51mBpSS269o
0riXfBnnTOfo+lBPLxIcz7zctiITQgjpZ1KNCS8gXfl71dzL154YW9otejE+nwpBcreadyMQykq5
luROS0u0t5qmGcp2M5pYC7k+A1rFoyk26JvnRe2xmg2xB1prof/i/PG1YgjXcSuvDTJ/S25JRAW8
HExFDZ9yBs6eXFe1YN4dRZ/dB7l9ZTYpl08m4oMpuJ3jd0kuSgU3EGf3l0eJxXG1Yutom9lhTGse
9zpEHUMUpd+wptUi/lOhld4m1g9zUfot7eKQnyH9s3ZIwqU6rcFiCpfoAWaqt/7m3tmtxQN2L1Tc
tPvaOHpHftHcyKu1dphjQNYI1Kvkrh8JLW7FQAJPW7vznbnUMoSCrvFVFncEC3LZ+yjuJ3wAf28n
HAqUQ8SVlxCspXQlqJ3RakP003cpoK8Dl02N4qVvXrKcpHq8r0kdOEI+hCYGl0PYgbVvNuzvvhwg
dNCZSPcydWANGoAFYPc3uUhpScqC1HjjO2Fi2n1YG6u9gcGVfoqZChTurGNrHLJp9f0E+E1xttyQ
Yk2uyV315aUYMeWujgE1W2vx9WcjTDpdckL2M+nVqkhQyoQ7rART9HICCgzoehHYfwVMTJJVcK1F
RY8cqlxezQzPPxW0ff0MVCGdhsnMqhSvVjFKOm3A7CIt2L034oLDCwgBmd5iyYjOXXruhIvyDHb2
MRPURzMxajMGWKMMJQnZ7b7YXmBFxABFVc5fwQits+UZUB+CFj/kgFtl6vbP2f/iPMjOUZRAk0Cw
mlf/vh9ODw9pnDjpdaq0AexWOMaRzUFE6/IwlPQQUz1xYlHoORlQ3Tf6J2pkA5raxjo5m8/1Dmeh
xZpkWWL6o8Cc+YNNXzm+oJ+paex5p0gVtkpKma/WVNX0iaw82auDXBNx/hLWtLF91K2EQ4Ey9aL1
celwt+5LctHV0WX8lkc7GV3pZtYZvCrNcpRBXcPuvJMMxeTswFJ1f9NsHmAEFeaFlstz0CvTJNOS
BEWU8iK1hpryJZhG/Hngt4gluB8EfheX6OFCMFJlo13IZeCtvLl4aubDgNMSkICcbBlK3kzqHZ9Z
5eZJCG88u0tYHahZW2i77XTQsU0iCQTJcS/khuHAbeBajooR4MOIWZXIyuEpbJvPtGrX34TVeiev
yDesIYjqqq+SwGWBMLiotsxn55iKZVKl4ZrjRXP0Fq1K4GclaacbSepQ8tlpGab8T+su9TT3O0W9
dYqpZAaGIgumcP/OCsKLzuZ2bwp4RXGBtuI7YHApr6gbSv063NRsZ/8dcwrlIvzecLihORetRee5
7CBqbxYRPxiRJMhY8eYjofF00raEK1PRg2kTULL9Gfy231c7gqB5nam0qWvwctNlICPSs38lhd8u
TxwNBYPq6HmpQqQzDqMtslfXD8bUvIdtcAxbcrOXajRafsSet4pnIQ4kKOVTLe/ck4wC2TET9/j/
90W9fXl3Xn9BldvYsrpwXf+GasIbzsQFEYt2WihklpdH2NcPTA1YuvQoTK0eFvJyoo89W6jAFeUO
ppr0STtiaB+ophy+7Pu6Smoc/duRceZ2IK8eagv60uh0olNcfDrUV2gHILXFiGy5kz2RpoPvJTKK
PhHfj/2kJQhgbr5FmqDZhl2kLzLTHHR7l26UqmhpP3bvhq+MTcnco6SMqFWhbwqZDxaGBMWbtBpW
IbReblVpwMLjzVDk8sQYXynZ70SSTe4SM843KZ2ZV+tkXReDS/5LeCpJl2L4ZEisz60PhuCdd9WS
qaSGWGnT14VEbTtQzzzGIU1lXDuBvTGhqV7Ve8p/FkYNh5zID9YL72R1ZLzESxJZmyeOXhkDulPn
/6PNjTybn2dBEXXiFbidBwUO+Ge2g0ZCzS9+lm2ZBx+n6RXCdg8ekDwjXwANmV8W9LZVq2MN8C6m
Bxkh6dSrsiioFgJu127tntfQ9SwWK1ujI6eWhyMqxlR5QTnGPvUy0+eI7yQGpfnyheL1bsF2vgH4
FoOVBj7Q/0T9TEYHjcYt2qlmKJsd9HCzJS8Hk2GE4wym0OtD2FZ9IhTVMbbx5soeBvktEeb3u/H+
sPjjBr5XtDt6GyIXMUK6x2eQ1w9JKJzxLZLAxWlU/+zpYYH3wbAjc5wSgU3f6qOFdMpa62t8361B
2ATblOQCJnNgRzvQXb8WgR2yh/Cr3Qdm3n9rBFyNEhrfXfikiTea7ViuqLsfXddYeCCSl+WKcGka
ywy+3VsKPO1H1j2byf95PVeEHz8chwji0tc4N343EgGlQuX8TzMc8tNCaMkXWXVde3BC+sQVQjhz
CEZD20gjOB8DYu3ErufNPlBnxAffK/tcu/tEWsZjPa6L5KXjuarI6pytNPKDPOga5RmPr3wbWYFK
VuiWNsa2W9Mjp/N7G1q2PwdeQWF3Z0TuRFdqFQbsC/rcScyUWsyg8QrhCl4XYxOZ3Q8ZTfWkx7+g
hcTvNM2dSifQfJqCOnP3IbPJ8uR9y0SMsxX4CPwFp1wGR+Y22q7NDWG+N+8t2CpjGg6ZKDqacm0u
2xfaLl+trntFNnehaa+CXXnmrsu9UHJ3yQcBgDnGy1BMYEuTF5NuJiZwe47xNdyFbj0E/ODoGllx
gSCyI73fN462UylRCHw66p1+P7Vhc/BnUJfzeJnLACS2o6pSBinN48TlriJQ/IFXIM9gU4lY0Rd4
EypEx5uBb/dV1XEWFdn+TMs+a/2+VChWSDtlklJHRqwoLhCX6EUNQIekgLqLXPwHtzL0BPA1QTPW
kN04Zu+xhrpdqgVsNK8/z0o+Tkl0yrQaa5alNxdXM9f9WVRkg0EgohaWOd1SH8BGtPp9LxiqYreY
9jETd1Gji+uh4Uw9HDbJGi78Ik0KI4HTxq2izckwlEA3hjWhlBlPCtqh4R4OxyKKc2kgPiX0vLNm
5IuMZw+PYB6/kIEsejUjZvhdCBlh1sNLSNPuCYvrbvzrTw4BFF/EjaGu7g3Ni8jgo7CM4EmbaeEi
pub5FnhxHpvomLQGWhqHlaZk1zaHuIOUb57d5CHJU1PNYFmdSLa6fzPp3wd1OOObC8vT31ajx+YJ
COe0MiPkn0pptK/Vnxd5aXNwEsOScHtDn4Uf51y1Gj71E7ad9PZhdl5EOI0IIAQCzRE2IRKn+HeP
Id9mR8VQeGlJi9MSu0dR6lDsbbuJj1QEXrlb5r97lxExESXr5A5cANSlZq7THHZEvtp6aSBJ0S5Y
bMZuh3rdbnwrwPIA0GtuzyDDhDwmN+dXDOdUYRT/bAvufYIIvZTCdO9Rq3GTP9yJ1CZzh9oHr64a
cL7e3Xn80NvR7s483K1SN2aRKJrrg5wqeWpp5qzw+T/vfUrogJdQrpaptpy404ad4RwQuAavzrln
Dm78OVRwjMyuhyD5wxWcH2MmlNU5EoB1kr8DBH0zUCxMyWSFP1s/8GmCtYT5rmhTTKrcuhIl5y5n
Rj60bKTEn0yX6tFfw6/UhfVSbbxlnPc5JmYwlSAXSp1JJU+nsA/mEVHbiij5QJHKEiP5NQEheG9L
qOXjzE6RvDTKKZ2Z/nqprDhLwH9TlCxMKl7xCrMiAt/crg+pIEx7Z3cwIB0cDE9cMwZnuRVKNFLk
g2psLuaPIh4At4fTPMpQrwBTtYlkbDJanJ6WSfIcNuk3ij5AE4NXmb2MhsQ0H/bqqi2eXRDCMYQf
2bjmYQSXA23RFrZAbdy7q0j2cLyniY6/onqU0oGjVmeJRvfcv6AnSzfHsVX1v/wpB7d5y3IQiAGL
tU68LygjK57s4xRRqQcd2BptEblx8kIgkSOtltGDnPVU2Ya4adM6iWI35tFKm6Wv3JPYxjyq4Aj3
0S61r4MaM/uktBD+2mAZYkkLE+HzMBsCMkUnemXcI+uc3rTNmY3FJJO+ROs62ONAEUH1W7Nt75MP
cX03S8/2ZTsudjxyndg28kmqcbzQYWDqJcSv3f5NVuqBRtHNWFMMnegimhsdfaQTjnC2TYhhG/GM
fuKjybAu0C178HuZBBxK5xBAVk3HM75jRVcKOYPKxkWuIwQWWTQQZxBPJi9Wm/IXdLk1YysRczyr
PzWxTwhc4dxfsi66BWaYjzjD03A/Spd01hBmKoDnwQ1N9Y4VkWq0pc0QFNELQ0Ma/bGH9so8HJu+
kHd2PNoDLAlU8T7xwr+HGxfiJumSEbj50wEDlP1nyPiU50H3w5sqnq/AkNk6wbly8g0m/ooXrJm6
ntLnFs4rUTpiZX1+Hu0AGRjcyF6uDD2ILzGz6f5MufU61gVUWorwG/Xt/AFztaE/FgTK9bW9RpuG
x6HR7Vq3DuaAqBJMuHQn5mBNjotCHP4dMjafxDSuPYYlOpunNYo4hSnWTgin9w2ZXVn4OQ49Inu7
Nj/liMKmnYW5mSqSnUKu3cwP8bNHinOVNHSsnxxrvqfJg0De8fgfd3WAHmIIt5cSrKES4B8UZnPw
B3gJEuPFVqpzRxVfjj0U3x9MPmKelQvrK9APUCPpxIsmwvsRHS2qz9u0D/mlsa833GSpJVZzm4za
Wmp6wvS6IBPE85uNMktsY40ncFVJ3bGKLc9s9w1AUC2O6yBzaSbfmN2ViScHnjrivu32BKAgDyKT
OrPY0cC7AinN6yAZUQYK1N60BdOluBgPMRnjqVk9CtgCueSofxemrNBXv4o+fJClOxZ6nzDKNycm
vaoyCpQDPM+bM/NYUhtGRWIpKnKi7jrTUpSj2foJ9IkRTrbBp55qWGKiYmEh0HxSXA8hoHHLG6m4
0hscI7H+sq2lG+mYYpLeZzmcE1tl4mgU2HGZixxBbQJYDeF3Nsm/qIN4q56CM9roaQmSL+0Mchej
hM5jFU9guRiRt3/RyFOyNbNbrTcGm+FObfTNSMmqH0spI0iCTR9k2u9AJ8b9yJGzcUV4l+8ilWDw
21QLl9dS9hAG6/drhuUigFIsdwdc8GFmbEDrxO36JjorQq9T9/vFDdjU8ohHhZzap4KbyJYYs5Ue
4lWxRk+s7DoMy3KfyoxJjmVhz1WfDC4MUngV1w0xAJNAUsU38VJpW/t2T+CI4VBe4TMD/HgBTkTP
GiXIQ7AbCJv1uLoHHt3OipV5m/8y/uJp7pUFtB9/DNVi4XIYYvsMck16MbffusWqUYf1plqOkz+t
Gqp0FdeQIegEvXhCEwYjAzzAGYhOZhSaDADmPc1p1qV0OxsYislKqmcbdyb99Vd27wKC2zNzunH4
GOQWlLc9kbNeAhM2TY2npnHj+cZk7J47DeKfiy+EHHexfWKQyPeDHjLyt7W9Ze27M7u9jyrzD/Mz
hz5rEQiN3qwbbNaGgXoK5Ts5/whwOtBg56KUpLsMXTCxHIq3Xzqnog29CKJ9JBFop0JdqcF6gFRc
W2FxoVSU4v6AYVWlKEK9euwTNDzXIKY54LIzIpvymqy4wBcn+XIf8syu9E+e5JJMo8EyuZ3XPTzs
9zlyqV3+5GteMcRbuQjo8ihhSGDxu+tX6n/hBqhLkzW96Jn0iSreLtmxPXXyMJMAER0ljYwP84a2
ejSZn30k7SFaMSyg/bxkDJL/JU0qzkmSl3wQfsKXZ09twkHBzaAEkAal+i/YdMN+sCSFiBXkjcTW
8M1aKtv0KO2xjK2bqjMnQPVI31e70b4Oi3mgjwfmtRnz7KTuoHcLaVWsqBRB1ljz3ue//V1tLd4u
iFVJ9kM9ZejCOYJJ/XwMN4ybLAaHsqg1MyRgJMkW8d9UBxyxqq6KkTqQz0fDGDcjnQjEcRrnUBTb
LMzodH8I5Wg8SzPUU3UbolfAic2KI1Z/KWvRPOwlHO74mfqbGVP6nGzXUUh6V8hs0jNUd083psdm
ytvmxrmVvJQCVcRKC5eqY+eA167Temi6Lo0CGkCOf0E7jko25H1fnEBtqEZZYKTvvjxtTboQ1/6i
J+kMkaDe0aFCRekKLDHUwfGp0svNtmQNbA16fy0peb0DJE5rk7xTXgyrnHkagfLVrh/TtdBY0Jbw
Hjn5bSuTozsH2Q8s2jiLAvuvyZ23pMMbpmCJTQsgQCqFql1fqGfBElprkHdBkCUgET9hZX+YD6TW
iNDuHQ8r88d/bTyDH11HzIrl8dCbi30v0zh2mkA3/crsfB89dVNHY1xtQTPURvsigc0yroxBt1rV
i/dGg7XYwFLT3twXfWt8vSbrGQ7qT8xs7qRZqLU7LDCd9jITOZFJ2ZcBaKzGeK8d5a1UVIQioYBG
RxOtYSkU/YAqMKv8UnWy6L8Z935aNIR8zXheBpbmijYbWOEr4w4F4ie0XRtalslvauGcJa8g74yR
FSRxFg4eBeR2wTVBh4xLyGHdTTH6mQhgTxa0GYsK+V6q9sw8Vqt+2LSZaqt9nvlpJmddceBfwUG5
uoKuIoMa8hY3TWZl0I7EQS3v6GvjtVKVfsAHOC4iJ9+ihdPisSaq4l4DLnkQ3JYfWq0km/rRdrNY
qCUKEM/Avt4eMGFlXQgwK4+II50mOOdUYnf0AIkS0V3p3XhXbO/7a79t+tWjBBTwFff846ioV4kS
V3U/r5S7gWqhEn/IfIQCtGYNTRpzWrC1oaa0eSl5KBCiqbe6EfDohBmiEigByFgMWo0dw0lidIJu
FwRwibjhiw4x0coq3POi4oE1zcl0nLGF5uvfnB7UTWCHHHBJisLxACJvkW2HCujQZo56fMvMN4IG
byWwILIQcQUPWCPO0iaeuf15Gd3wfyyNrJmcwEHYMl8+8HIDand0Sgj/fUZuzsY/SsJvry3p05AI
9F6ci1ci5tn7HA1dHLidord2umXexMDKEu3SYjENhN1gzgjJ6lq+1epHCt3TkE+Ulmqa5e/mU/LO
5vB3UiuydYKRW9VT7kDytyYndro2bTB8wSotCbGyYxlyM+//zA2wNCndwWuLT62mhQBo21Seiypn
OkeQXP5Z582QS2NqVkP0NPkxfRwZBW3iXIqIbjgy5Fq+UJPcoJOcpYgEZ4bnQXV/fTi/lvN+yjc4
Xcy0lmbConLhK4z438nOgaKSzkloCT8T8iTjRRWDXcV650zedRhboxGE+0nUWzqVEPQrbu56ChPz
pzLmNJ0hveczVsGeQ9ddoWl2SpmHr1wQcWRB02dItQaxy9rNKQnI12TxuQwA0t53/IuV3fI9LxX7
sLVRjMdPfi41nECXiPBvqgmgJG/DsESTG5540sCpTDs3JBH/Fnx/c5U+h1YGSVjlhDO4ISMJyV6h
sfkRBmtr6VuWjT9cP+VQyX0GgB96cqKOVbv7F5jWv5rWJRj/jjdVk14uK7YKhE+dmqP17mV7Q1WX
7vcCcYdWgIjWicUKnfZkwq9oP3nrk6yQTdm2vQJRn/9cz4UU7xC+AVHFmlUf5WTgvvERHwBWEoDX
CQ3U2q1quyoN28XkluVRmFVokf4wzenoXhit41FSqWGqlKVenhCakNp57VgkFXf/aom25Ai6OIOr
GHJygdoMvo+zhxaY/DIArUX5CIq/0NF3JDiBFN/z/42Ou7knSxcCjUCkGVr82prSbS4F3ZcIbfdg
JC53pTKw/mdwUgF9GIEZJXtPkFh9EV7e98fvpr7IUDVreJc4AxbxYyCIbZMfDwDGYzQi7Ap75yr/
CW/ESGgkhzhlox5GVbglS6Rkcn2lCnoo9rzKF9uKpMy6il8Ksiwed1dSWvYg4PqXSX9bkeS1houp
XMX8V8aRJ+DgvuG4zpJJT/utHn3OCwjMsA01zTq5SDBPTCvQGhsj83PtfVus+qzlLmPwNiugRN41
HpW+RYxkDBp/FSORSnRKychTgQ+8tq5lEcZtFfkxlwzNK66+ozwCY1tvbxPkjVhvSzjPLlmp55Va
oF4Uur+OlcTX2qaCs45MjzaSLdOAkruIR9PdRV5RnDH49XUSpcSSQtkPljPOn7t4BdOrO3qTvOFA
DgUUu43XeQPLyCu1NroO/YF2J38eMUtj8JL542+l8AobLahE5TZncU8XOUbpyvp/V9NBDPgf2Ohb
1kuwXKRHOw4z9jnBdH7/tepPmHxtrabsZWK/2h40vdZpEq+jTfZAgsQ13T6F1vP+08OJRFxMf/dw
By+CNYYZgy5oCuQeGt/1zr8P7/h1LssFBKryZokhZVH4ibBhpWNbOzPL3vmIk2ceeI1XBOECtPT1
A0EXiEqGtqTeaD1qYAK52HlALsmdY/ITgRFhBBrkHjTqIDd7yh46cvZHBJ5r2ZSvW4nHLHdRGO6f
7ALcwZJ5WVtHh0LuGtFgHgi09dNyFBqXspHyW5oVw/f/jKZO9UhamCD2qlpn+fzxZ2rB+OONXeoI
W0HhSEJdfcu6MMJJdioFDc61TYRSPAFTkrbv0zm2j5K+ZTvN9q8cFuPZbuCFPzQbHoRinibKNIR7
VVlcXNJMl16IBgDgFr1y+nEX1of2I8FFXtESLPn8aVRbacuMZ55++okfVbLUwNqLPT3YCyhkna2R
kwsVVI0l5I09BNSEJCPVsvzQQJEsIhFzulzv7+/jv9Aa4fSHa/KsbShvJkE26N9tFadVvASMoKoA
59YPdGI041yiPGqXfLoB7R8oWREl1ibqp0E1NV2i/D7Zp0Si+/6kCHfDdQLwl/dpenSvkG43sbJW
llg95nDBjctpsJ3OQHNY1O2i+YLlN35C9UHBDFELa/riBZsrl71CnCX+R8OwoMfdPACsDjBv8HiJ
5QbJ2W3voEkfew5/hV0otEATwI1OOSrEfXxQI+lPpF5TFgIC9HP2k2C1sDMR1V/mbK4R1ot6oNX1
ZLs8gonHzYsOxC3paS/IZVYVG1MUGuli43YQ57p+e4Ht1Cf6M8KB4qe9qrVU5YQIELGnOmoccv5F
OiBsxPmcN/v4dRiEk8CRifed7rJ9+NnK4fiVHwcjbY98C+gCd4UBUTTUG/7a/s54i93B0NuiF3ct
OkhK9fh6f3LTPRDmckdbh4HVabY5Q2Ee65YIHnOp8dzqFTEuGAYOULsm69rPBnDw41+t1LNhdFI0
Oj2LqrlypAom+BCMiAJPu/02t7MVq579EvQNFn1hhrL0i0GG4+Z5zAG5QVfbBD/YmBUG5hMk7d8Q
vrhAgRfs9v+bAmgng9lwHmuTc2LKkcwrYn2SXQBpwFu0u2A7aPFftXZuecO3tVZrtap5lIEp8H0l
vt/R0l0hQptYYLJPsWS0m9GOMlvildc7fc1VTJl/0TeV/cp4Fw4xMEldDn1OrLs79fZv/DTCOa6b
6Y+tWOEyJmnInO6upIPenWE7zjoJo319txk4iQ2Kmrynf5hoLucNFtkVGA5IiPrhcC/dBKPQle4J
fwbcZEhqifHdpIxNXb+TqUHDp5VvzCjhaTtr7SPVuRDFPB3w3AbzpJh3ucF3T+6bmHYUVpuDAgrW
cDrwE3jAut4miakGLyQKY0JVk+NydIXdBFOsQV8mdLybfRXjNo5+VqcHyB/8MbpTnYptfyBt3y+O
IueUyBPAg+vtdSb27+qUtDIS30KEviopWZGSu4gDqA70mp3+V9tQyNdneHfhqLQ8d8j9MJyv2OoN
MKM1zGRh+SGWvfGx2lgPL8mfuNxuHlw91rwbYr8NFzeQIO6Up3zgV3jZt2f3Pekopuq9BH+qMF3s
jyqUr5cU1Vm1xWPAsqufsSFj0Gj6XmjwE8WY548VOvrV1ShjO6BsIuIjfYrC/Ol/qEMx5PKiGcHn
CWcn/LJ6txZmslgQX9R90+q/nG2hxcbK70loCV7CSLMax4ovCpy90VJZ1Z8DMZ+14o+0PC/tpMzd
t040aef+XU9iOKdVH3L8MIy+3tuClvLJYeKHYLNcQLS0aLQWbIbEUp4khzfsxfvFszqWAgyXnF0r
iAczAXzbVEMkAw45pEKSabu9VRqtNcvxcXru/0Itr4hZU0/mPPDC1Z0/Go9lDUEzBWwTLcbgdOyn
++R2U6eKwlbGY/0+Dm6wGP9/K6Ugz3V2TGL2Q2TnUz/S0a57ppswJYU1vhp/+lhMYB2X/HDPUm4/
Aiwn32k2V/V/sd48l11rD5y60MIyMUbqF7Tw9SgWRbtnMeIVNZ+qwZY3s+GLRSMbDB4grAWgBmSP
NBMKMLdtAwkxkNNKPrl1MKaOoBTX0owYxQu3Ho9h2Zplle7XOeOlzoa3DfRMHa6ouRkWUlOQNsih
hmCdktC8PT3rw/trEIZXN3aDHNxd7Arv8Mq+3CMTqshR425rROOfVOUwW6XUUHnIohtwLUnpvnsU
gywBTGu/P+a/oft4N0ZSdf0a16gfSKpb8cI1cOktVqkZrZkL7fWA3XZdclfb/pQVs/rZB6OX/5md
Qcy6oQ4yyB2TJR5OEcQBJEbxI8y9KGGvJysvjD/KgPmoIuM0FfhVqThStgkqFM6Mlf0Fr/MF9jlb
6PoUzm5yGeLYUTL5+Z3JclT8gAXMW2CQgYI+wmnloFaqs6CwLdXRgv9Qqm5FCrJLhj6uWHzNLUbI
TI2RYAsCkx+39dQg0uvBUdp4RIgJQge2+949QY98n/HOgG3daWGIhR5wf3RR/jZtwKjU+fFq57tr
JRCTvsF96nx/nj/MxLQcrQIS2SNC4h8rxIPod4511omTO2aucvI11rE6lyQ2M/5ttU4WW2AMeH8K
0MBKM4KofVYzhboxswRcsSpzbfnYREgcICE/dKaM6329ikNhyzH/4h/RM/Va6aFcYGWarOt6Nqqb
tvKk2KBEJD/7c1HJaVSzkEz4bmYkhzMBgsIdcLH44pcwLtl40qZtUJqYC5WpPmJdZ4HtM5AL3Gzo
2K3WtcYLyJgdaXBv2CRfaTkg+cY1ThM4j9KodDWdJPG7tyvoqKoHlm4Q4LOKCDDtFPicb2hKInMj
q8JMiurdFZavGrIW/heIIolqcc8T2Y+pn0Q9GCintO/ox9ST9jM/3BJOm920LD+ui2LuoEqxje2E
MNSP65myGYczP8gnTPtN2sozuP+363Ze+T/JXArzugX2O9VlLkCvcLsoGUZPQhYw+QgsdA37cI3P
qnv5+e9bMsOzf3HM6VrBReTsdyVtuTRqY1z6goR8Bple9IPigwqim68qk5UGBvbkF1AB+qmgC27i
5MpvAerA93s6B3ixK93xiqj4m5ui+cC1Ge/U/2FAQEC2TkGo+PoDoDl6fZ0Iw+QcE1qdX0bK4SAG
/umcQNrjGJtE6BD7aDlhEe5V+00abAZR52Aw4hEvQOA+LQq0IfoHkeNtKT7a83cnHXL9nQ3MWbtv
3AbC/XYpuWTChgwM1hic7Ct1wo8xHUfpVKjakBH/KHXX+EQwVlOHB9qkgavAPZYAKbfH80EksR/z
B3hy3g6+LTcAvG6tJUkCB6N+Qa7W50Mh089HEKGXSYA24NgTkvOvuM+YW1nhvfQEizh8prxAPrM1
1d0o3DZpfIoT7hb3EqKyxfuRgZF0eemKsR/u+p1vbIw7kAFoYQrJWAWX9pmeI9b7NGVCy/kmTKui
rZn2TcDCCmU8W+RlvFUmErwhoR6KfjFRRUiz3MbzBWFNYkoKEIN23ZujHrXTVMEEQE+kruHLUtCw
DlQVBvtnvqD3WEIbzhvatGSLrkzhvfUKdLPjww28PzwDoKQILK6n/r4p6LCbfMs0inFtJa4Wnt4p
r3R8mVy+PWNL50IKeaQ/9+7yL1UwS6BOTw7qb8bV49DBQMRye8OvRBX1pjNTJIR3UIVclOPyM/1M
Ps4zU4XgqZqqB8pQuLskYcuM2W1qUxP1gLMP544JOoFXXJyxhSgxUD8ZHT7kO74ks1Pfb/x68aem
LAHwwqeGeWHSIWAcgxudTLTAudB4PxNGnfdYKcNjEyO21fMJruqOYeMYypR8Mzn/nWVi4jZ7Ttma
CIUcluTdjeE30cXBe6rdvRFqQQtiHOGCLu5VN8r3/LX21LgdgXQW5NBav0CjyhBwtv+a3TFeVI/T
6CEpCFzlzhdakko7A+pttEyCHhiAhK7DSgHNWmykmSPprWu4ZIHHbQAkjt7cRw3nximHGJz4Uru7
ZrISNKCxgU3YGZdW0CA+VI7k0q9PjNkWxwwJUNfH1M+wFemm46LRYxWA+1ZF4xoOF1VGDHazhhLx
CFIRpkFFWSbQoPEg3lSZegPnDDvq02HAQC5C/k1zDKa6AKrmWlFzkILMCKsMmVFeyW+qx06B3Lot
T9m5m7dSTIdbRy9ypfPdn+n3dc/L606Hl6YbTAr3H0WXQxJs3ywYxnHRqGZRhimcpztcwUvV1iRE
6Wg2325dhgyjYQlq4x7m6mPvz+1LucaA7NUD+1b7D7uGGsStlUJnb53R59ZgYTvGUCG7OBuuYC3V
GRaTFoc/9hxxkFli7UFxyJO6Vw54X+8SyE8mzlXfnvf6an8H5NT/XjdPsgDFdcBLpdwluqzHsf+y
PTMfNGFudQfyM7keZ8Dxj5uAREvMVMID5XRuzTBZSA/o69jhRNpDVm4OtobYMtyAgr2rB1VjsO+b
Xd1+XhXuzNNSTW3X56TjGZVT7caU6WWkm08yrh2x+mKrIspaHj5ysP2POrfy/jSQDPG/trWmzzV/
AAMtBaOLQjy3u1XXPTFG2qT/Tejc9sOIZ701NOg/JSKu9oUm03zVWd+XPaFdO6DsO0S54ETKoc3j
5LEKHXKXTLhJDXks6ohGn5bi+Y7TvVM+tAjMVm+8QW9vIFokAOaiq0RYrB2y/A5/AnDpVeRQyP/c
GmgLQo9KyzffvzEwD2VI2Wd/oZngIvmH4MqUKSPtq2R9BPtnS9xlJQv7HQCYdb3vpmFi7HOWDF1x
QUgm92qJfQ77GTQPhGWbzxxJAXkGRP07XVhJMCVD5KBUQSbPz5nmbpSM2d/Oo7yCGnC68Yi7BoY/
VHQjYVpoAUwwXTCLE4Z1j1LN71OCDVTkvXGx3ffHEzXq77+R+hNps2uvhBPiRZ4AcRoEVam7dIYO
ANJnST3FoFxw6WsGATIByabqjLGuFz0z9yjKqBNN4/qNT/gR9lk8/L9GX720+mS05FntoFTIb8rV
JReA0F4E1p2mwp9bl2KMz4DHgSTM7IgOH30tVfcQZsgdNteILCbxf1H5lI3P0juPNIAbGcaTth0E
b9gxpsSNJuZ+8QfLYFVBhS+1XMf6nOq7oaPunN0bZcqAi9jA+RcZ4zGx1Ux7bMbxC9EBa4zLLrDg
7y1OY39nUX+Iia/u0u41CEpebxZeCnQ9Hu6Jor5wPk1RiQwTyGfMI3yDhyaw0GMH4SL98OKqTNjy
tBtaegu6XnYrxmbWhFlOr+im4+Ejc9xOon3mmYcxshWW1sOrB88IzATjhlJxXL/P0kXfz7W04vaj
zLZkjL6VFn14/DAHmP10xOC3hfJO1V225dxyjVdxwg078It6bw0mfQR1dyIZTdwkLS5iQ4Lef4AQ
0o/zQWHhTp6JpeaDZdwbccySjGdDMGeEO/QswrhwwVrrSmuuH38ekyGtsK69lOpbZ0slEmzPrQGx
6vfH7MyVLoEfEAF+h8leUXR8SoIWWLtLjgPdjc3lZyklJ3o5UF1dp+zbsU3nI/gOkDh2FU/K99c1
99gf//zl6V/mrOtRUxNN5Xr+im7NtA/VV5MEzruSRWqK05ofMPZeei4FtUSWPjjJ/R3w0utaf8EL
8SqKH6X/CmxK3kTSGeSbR/r3wH+lWbKiYHM5mdHguvBRaIWbpr/B9qaNF/FsRXKryaclKcm4tQB7
xk933H94aWYcJnhhjue0ktyP2Lv2XPeM2ACHzGj/MVEVOG935Ti39d+9naELMzq2EInAqcPtU33i
KbbqAGYv0SNxlqygYzHCndTOTBABw8gTUbQnRD7b4olZntUZ9mimFY6ErZRFXEjN3Aw15Heg3txS
RH2NG6+FlY6gEtsw/JDmmOL+Lbsz56IGRO8KZxQuDBKMU02eGtdqbRajG3XCMBCAng4toCcDaKq3
YYvTxIvrWRWOPL59fL9NfRgTWU5JON4fjkidH6Rt1mtJeTrKfdWkY9A/ghzmIPiwEePqoOBNuZS7
NjwkFvN15lVsRqnu8lhcT1aQf2Ygui3f/4o0xLztVi3fArR/rNtshbLDcaTLVe6nhWDDJ00TiHuz
e6yka+UXf/C4tNEfvyaHiiSUCrLAN+uivknKeMP9nnQmqI0oTxBGnuGEI31KMn71L9a7vQH8+0Cw
BAzdTbnDaLmh1H3qI4/cAhGlcU3ewARLxlguYjsBy5esPXxUoCcs73prXDaBbKKBuAjVPPCoO1rM
4Nfrf+sjEZCf+QiRoPLlJi5xPyIoKVU7Hzq3LYvYOHt+BAVgL54N6748q+PVrE74mtr3Gxy3kM1F
jrZVazQNPTmwhduPSfhqGPqxcji5hLUXmWA6Af2DPXdOIpW+LsdDV43KTxst14nFVj9bmNPM+1X9
pSdpZiZFzt/KDliA5ecK2NZxoBTdIMe5e4dosPwyLOIMyJTPd4s2ClpEkz1al7QmYT6pLe8Jgf7x
QYVFN580D3kI//IZop8p/xxENohamJmWJf1YhwjbwxPM3s4fVGrleL1HrmWNh0UBcp8RGKnSWxDG
mPTzX8ToHzYiLHWz84CVMzPielVt1QuZxgzfoTVKrqxXytvw9xoxt2QuBElrB6wgC8uJyPnLLvPt
PaKHt/f9bhVOZE+/jP5FStwx4NPnpecykc/vebi1/1rpMKFLexYMHp5Raxp2MM0Y5Q5qPNOAuhSv
rIyizP28PKrIHJ7/wMvGNucCW/87uuIeWTiurv5sCglnfSueSexpHMiWu6CwxzERZXTDQuSR/aTi
99lf/78pPXw9jClqZS/zGbCytupE4g2ztBJ192t0tJNzTs4muYaVKiPFIxr/HqfrZppgO9uZ4DHo
+Ed75OSPpuMjeCvKYSuIJXulB6qIODV2eQop16A2oidzSyffnu0uVIpg53dMEbbe0LfEI0SKi1oM
o/AIYdC29J1AQsvotl6t7bzaztC4shdDpwaXwu87oEnlfZicYqmfPLQincWSYwoAof/e3g0pdOzl
2t7L6BhvMZO9/Rmlo4MgNjSoMtZ9oqMcKXxbYGBfUxOvn5I6Esqhe4dYxNAr2o2c8lcHVkddVxO6
emIcwpkIv2oFWqGheulS+SngPZ8Zw38b+fHWMrF2ghdhZVxMJoc43q4HONWKVjHEp6GyqdhBJoKr
+QhfYk8E2ND9hhwd+d7QrMQaOOo6MQzVnPtor/XYV+TRQQP1PEACsC970iTJ3r10lavD1nYytWX4
mDoVzeGG3xO660XD+E16cC1mw0juI6sl70ek3qg/gg6Sf+sjmekVvUcETBomghPO7ZrOvo/EbBqV
tLS2dbI1KVoeQilAFxTY6cwLjsyOhl/9SwmQZxvsmeaWPm1g96dAljw3g8urg0fDWIAVNcZnpKhm
vFAIxVPg7gt338TnV3L5x9vmuPSbNO9VX06KLzJCReW2+A9nRu6Imb8T/CxKlHsXo8CerFhrZ5mB
ghq2XIi6jlU9Mm0Ix7EFOISEsIc8hvTZSYWnJUUs546TpQ3dSPzH7CQhzB3wpvtvXWvWE8XJ3QwA
ZRh50ExsD5EGeGogmbQozNS5IUU0+K5/zbjCf7E/ecq5PvsO3tIvPy/UB3aXfhbw0uayic47znT2
rc+u+ec3JC44OTDiBb2sdVHhZxpOvfNFO4sR0jgLQbW/h71mX7tZd8umm2GM3C2F/QxmgBLl5fq3
pK3U2GDoHUQ7J52blLjIoNkGYTi8CSubd62gBBLoj1wVfh8ur06zkBU6ACRMa8+yzTJzpQiq7noZ
oi+ZFKyuRbquDEA+jk+7f75Qa/sUPod553c0+cvTfw/vNSP9hMelu4aLg5tSi+O3t3QIZdRENbTL
LeRDifdsmwZI2GthwP2blw6XFhr8AM/zapiqYtmuBiwTpNGU8WnjS1LpE6mB6+qcmzwtpnXEyOVw
zrDUFZDTZH/bU1xGy5CO+iXju98pIFsK7zSxyCxZwu89UtkxtK5qfTrJOg9XcDT7/oReSgfm9ezr
Avt1ENqCCcgEpjNTXKcpzQtjeaI5RnsKGmb+kfQoWoCKmCqrqCtWyvx3SlpnVK5e5CYgrptE15ox
nsLrF6s7E8tAmlRaGvy1rq/xDsvlGeK+91tya0/3p5xV342CHJzq8bS2tvv6ViPP0VzPB1zj5eIp
lTNjFqMvdVZxH7+9v0MF+rFysIr4RNYmXPzmJOrXYi9GBaAIWAi74rcdLoTyFHlJWDpPYBwmMCpu
TCkZUR4CvxhOikUAe+GzpGa/4weXkLb/lOnXSvW1vyfOxBJXoXfCyTQupbIde5NnCOKHwgKcMviE
wrz5FRLKYXEDHKQMM0RmxYOKji2oWQMtIjq1jV1Cl0z8Tby6MjJkPQdHOXKyASoI4KxQaIqKVcDO
6K5EFHa8YjA6YiIkTAv4znVVCoV2HtWdADlo7DeHldW+btDPgsMkwcmAzlrjXJdWeA8UpEVXmsIB
4x4eRDTYE/L3+DsWrBa+66gKZBKfYA4JlbafTDoURPe/VJX3rcYDfljGMQLmoOO0l0iVrCvUiJTF
0zD9/vIaO4cbfww2hwKQ+Ov09vW67vyjYCCyJ0o6uGknY7ZdBscpGfbLkQWntgtGB9ymJiYJaV4G
OhSnFFisdUVYEQFFmJamhE5iP+GUM3RLoH47mQdYeEoWYqSu327Z9BG4aFDl97d8TqI3MZb8rzo+
Ntf4nn0A0aVHqWFE0t4ZoSHZEutzDEwMAhI548IXDbbXDRPJsuyZMC+nfZDcdocwaRRWlnxCbwGc
bCXt4rW5NU06fnTPVg8ZbPD16O1w5JTXOutKfhI6+tFX6m79XeJ+/EJkXIkIraRT1BiHwXpUeS+f
kNbBXMAns83H+R3HWPYL9NWAb9CWhkeXWFH8HVmOTsjBlXmDi8Zb6MKI0f9GHst90boG9wrJurr0
ehTjJX1SbHhHH7X/omvGiGieHD5EYg/j9hO/FRgEkkv6lR/lGd9m5H/bLpjOns57lXW5vpr86e+M
IL7XggmLKbEw/ck8Lu7bJQUHXZVCQJOX6jxewxJH1D3GFl+sTqDLSAn1Zv1S1huPI+RYfd1gYLUb
LpQk666ckcdgq97h8+qEtAF4MR9SBIBeS8hzJ/dnPZ5FfoI/9+u9074KB6BPeP7HKUFKMt8X2b3g
Y3SW8mb1CkLG01e3vPlsBAmRrmaKqea5PKXI8fsqtg9NCxyPx+cvTvbFLx9yxwwFwLcYWULs0cjT
MKQfoGOWxT+s5UrFfjH7SvewbtsJLEJNn1T8h4iV4FuqLD4MI6ZjYYYB3H9fhiibdLgvOP30+OWw
sFn8Gh0sdCT4wPjg8uqF/eQtJsyjjg0bPd0Zeuiy+jmW1BURb/IPeL3F6CfD3qcecZQNJ7FfY3k+
SD6iCJ0pxTJOYp/iWcSmhXxWhjwbPowwxVYeSOP3Ie/IHBqB1dRzT3rVBfYIsaaqYmJvtsc7JatU
K7dlvhx0LGAklWTUBVSFenxxpYlkTPzEL53D+APECoL17bXa3oR7lNlD4e9eNj5vNfASxG5P8MO1
yD2hSi4A55IVvQ/VrmTJM7HxOTgK3IRV84Tu6ZNsBaq9dpcHPruQ8pnE4sAt5U5N/1qVMT4v5qFx
nuzE/pDNztfekZF2vBAJ336+KuP97yEV22IaL7jSEAsdrLU2q0Tx+6V4pfztZGa/YoH++79e9rV/
eBasbMVCz7x7pBftY/MlUKxZT4RN0xfN8f7Ote2Bowfqz+b31Tzrshsf/sr7TyBfVb80foEHpYak
KYe5OAbn1we7jiQcCjTt1md2WvnXsmt9S5J2IO3D605YMmxAHqOT2cWtgK1iet1cOtFEsfFuCQ3t
DZWDBJPOD72p01RrWsfri5iJBxeZQOhjbqVMMZui5JBHYyojfEmaf+SE9BHvJhbfOvlSkGkKywsn
RiQhJg2x0IzB3+HtleoQQbMeJ+7ZTkw3nSel7yXZ54dSqbuV1P730gK6coagWP8eeBio1Z9Hm1B0
Wa9Dw9x5eDekdrhFEPr+Gigj6hFD/Y+PaLXFvyU6VyeJYVexrJOmFwOw6jBm4H0NyESeMYlIgpjC
aQltYqkI9bgzE5O2y+bixsIEsr0l9XgXCYoUaRbL1+AUh2R8FIG9hxEB2jDmji+HQ3xIUvXkXZsM
hf9yQyErhY01HBlwoYcPMUP50SbOiyi7Tpsxhly2PqF54U63HG9GmHkvMeYSHUwfcROoBYeIhEg1
CthIWMMEDtykpJCLMN5wegfRyA9ZdwrTZ61VAtkls3VaF7CqVMyxYeXS80CqS1Ki5dkKtJ5uGDyJ
bsSNAiympnOzRiC+T7rymxnXyws3jKSLgxzd5d+46Hf1B+8BSxfTBhB8Bfmv+fqE/yf8q2pw9Tkw
Ff7S5yUdNIeZj6vvWbzGKyMa9DdZzS7OSofHdy5mCyg+5zimfKZWO+6eiGgomvigbF2YAMn3LWzG
+lfttLYO+ACzfmCEhW9JDFsgtJJ1MHs+X35VUXMuk4aF+zukrcGXnY1DOKBDWSfodn73iRILU4Vi
IDtaHKW1om3t/yPdihSSWwHXhdRVS8IN1vj5rcGSMrImGjKgLBiS4lmVSm2gVbYFa4+sOKk1Rm0m
ISB99NHVJuflTphNw64rBXQQX2W54Wsg+jyTT6hSOXOErQm3fTGbWI1l5OSbEts6djFyyeD2nkI3
uc6RcIry8GNcY8C14bQq53FqorMAz/MY1EfO5HIn9X0T4zWxp/92FgtAyiWSHn79n8j4AOFv9FLq
/aQIGnHrIsuiE1XjIYIhd/Sk631fCAvB/SLNO1ITTBWwLIl2QCHXx5hkR2uKfTsZcaZe5+E8lWro
n7DAPWUBp1Jkr9BH90ED66d0z3dQCaxHGsNZFaxgIxqUlci1Tgn0Tly1cmmmtEtmJEiBzw5EGen8
JdxYxWB9+OJI6jWUeVHw+cLjBLfXKo0rgtgJXFiJ2feEcOZew6hab8HYDDYWvLWR8MWGs3AtHcUe
VK+v0jS/0AhZPeVkjOnmO5CuFJPKjJsorAPvh6ZK6ITkfOkguQCq5zPgRuw9jEZqBo9GVNB2ow1Y
h4dzzkyZAsA5x2Dh9UPClUJWY9LZHWw8UCfmtq28Jg25DOnlaciY/cb5VKbIT1QQLUUp9ziSCHjk
/YjM9OLn+elQ/SdVnLpEej00PnQvGOu3urJhBDtxkkOz89l/4xGS4vlQGo6e4FWyrVkpByAKRgKb
ahEg0fvULmcEghIZ5lRus4kWjnX75RU+19Gb6s0EW3aggxrL8Rx7/y4QhwbujYv5WwChkVi/u14K
RSvY91trNNgafktH0n2pvoXmEJJXCkGQAvqFTCHC/Yl9uvskMwzuxfog3XEfv6ZT2/blEaT+/Lbf
pO/D4TW4p74BbPPnKtiMTirVDQ+FP4N2B62uKgbMj85owJYE4ZxIv673BeAIfTajX12RxT1CPbmN
xK0sd4zOhMjePhb/Ct8YRVRmkvQrfzvbAyobKC6C/KoXL3g1Jk+GU36WqnqFqyitPc/t2XgFFqOb
acq0oDMmsGVnWMHpfv39NMdMj2EjyHC7dkYwCTveniMepr/piwKr2szYOvsfg37sQBnUD2GTbrX9
KQonDvUe2VC9BRoTEesCZpyXfzf6HNl1q0U9eMrqagJm6Nv77b8OSCk2SU+S4qLbbKn3B1R+J4iH
QQM6WGMprDg69RpdngjzQegA2akZNIVhXblTua/n/1TY+toyTyIyrfIXJbS8cfEOiqwWGZsvvPiG
ciCFXt3wTeaJhR2NwAcTLu+ckg2bm8wNvyTtPDyOxvXayhRCvrNbVQt+kwxl6nNZu/3l0R/CCbYQ
92fzqF1tAcYwYOAXYfp4bQ92nFcrtmy2mK6cAndRBngzXdCCXhZotr3/jFcC2i1b3q1VLf+XJKpn
dmus1Uu99Erii/Zb3i6Gb+C+DT2oJwGml3d+oBWO/Zm8sIQAMb46DFXIMOaUOdcvQIR3FHPclQ+g
MBLAb1z73gDQcZOT4PV5rHbNjcUUD9bSpMl5dvidoYbwB7GwxgD9clJAde+nnyai4B0q0qplai9g
8ZeJhs4jpswp9d6ni70HiFCtBk8/g71BviEF5jZIu9MHGICTEyoNZyzcuFiQ36yzOrfvCoaNL0fl
hLdGd3UThY8t4Y2/qOOv/+fH8+gAXRDH3u6pz98sIwaw3P2en3we8J/UE2uPprTkdEXgFYS6KKjx
69tjw/vH0qKmJBCtbAhThrE21XuDMpUQarJ5e6Vx4KQB8mLb0Q8i/uHbvBo+U5p5GPEW+6YP4d5M
3MzF+f3odzTmheenhuWLgsEBbG8bZYEtemxGXCVzaWmUsCObjXev92BXwFC8/kFehpjQb9JwMXpC
VRnw4HhQ2V4+UiE0J88tPUhWgQ3KweC6L0U+y/Nu/UfbqTPKlfR0xpGpd/FI8NS2jNhzPIUD+dOE
reFcDuBvy7ilwboaOQx/pt6LVl+6DRrVLo2PZcitllCdihfCwahY7kPAm76Q8XvMuMdZ7ivSrKVG
Z3l9NPtOZyFaJcZQqp7i0iYRFsfz//X8tm6MR8lZipT53iRW9KCjo9eyT0BVN5TmPkEow8hpf48a
T8t76tafafHq5KCU8i8dPuyWaNAtylawoUVvAHm40dbxoD3IqRs/3fFMgqEbY/swZXWJOuGEqUA8
q6z+hlb3hi1M81u4Npmlxaq9OAgHnQucsNi5GkP3VjPksQjbwO7CsqHx5d7/Bb0DXJeWjpXnj5TX
w7wkj1eS3p3w7hHZq9hbXhS5M5DzHRLyOyhTKfk2k3UDE2ysgd8+9jE+7JQBqXm5o0FktaDwBPdP
pPGHK3Ct9QELoOQQ3EdCU8QFAH5UgEY9cOtRNs+ewb3lnsBqJ3LB0VQ2jLUY0sXMknfBXdLfJ2u1
ti7G7FQRY2tXEL+WUqG7hP6mKiIQ7SnfQCf9ezLmruFz/aXy3zdEn3/cV0PYsYcmSPdgvyHjUKEV
5NVDGdZ2jtHng24cidggc1eHpOn9UWHpQUORetPV+VZCc89W4QRnii+S0rQCFXD1xGUrN2imGabt
Jp/RFmX2MQ9xD5vZr3z8GgA6cayMuD8zFlzMsTjy0dH/d5xvvsbqmgyLKSmbhDh3kxMsHnxsM88G
4HorqwOvkcfFfWjbg5dhuiI7Os9oxszwr2Tg3EvnA5ieShfj9kh0uG3f6U2c/n2PLj8f5XxS6D1a
FVrhsivzxFXZljlsLQRFl2LiTeysV2Mnl6QUS2hXFtgZeO4G60Ch1t0juyls4Wx/7pZlt9RurN2Y
7j66Nk0ZcZ8FZaYvTzBR3qLcr7jr8CbmWAF3iX9MZ/o+YWCyEiCv7SbqhtpNPYPlX8b3pYT8TNp4
V83XytDaPB69KhLaEXWlfcxAcDCqLsa8NguohydXLkGxj9uoXdiGAR7pk24Ci99qePR97/pmsSEZ
SoWTuM0CfP4X2e4V82tZy9TOfmtv4NvHEJFCNmU225PKPWYeKb6fz1z5t1pakZC8sPlBgHgT2Duw
YNQWebTUJIUXgT4Vp1cojf+YTtLdPyr+X1EB6LotdCOdeLmLvLRuwPqmmHjYgpeUz+blz6z0SiuY
WaW+lnK/r9jEMP3o5h3p/y58af5zPbKdTEBxDdAAqxt1GZInrtN3lw3WDuzDDioJKWz1i9SglbiR
MS9v2yxyH2MS/KgpV5ELBCDGewDY9aQMYoiX/2dNAVl3AQxqTdfhXDdVwgVDphKYMigF3O40zs3n
8g1nPMeu79z4l5WbtQo2sYFCTewjNhVQFL2W6jp404p2Z5hJ0XCT7Y0Pf9ZqfA8IuHbsODoduR9B
ny6N99VIivNsgMps0BZmT6XwceUS6O1JSgW1Xk0yk6v3Q4VwH5Qn91F9f1Asxusnmke719q3QEjS
9/FwvnUkLluamITL0FkAydTfevktMio67vu1bEbR1X3vcfRXGh4JtWukYlKSim2PtZiCPxeaM2BY
Bxz3srPChKPJSPO6lZP4IXgAJ827gqcFlDmGiS5RZJvDAHGf7F8sKTySppwOtYh+7oLCMXuYFhYH
7fG0AA4X4nYcN8FatUjicyU21NL6eJ+ttEkU0dqIKFlzVMnEeBCK7jgqn6Z2u/SD8JfQ652l5zag
xsQcK3sllVkwA5srJK9hBM6jL1fxeg+vCbFprCYBCSBKrPMJwzEs72hSdr1MnbjzHr81S/+X53JK
4n7Qbm50dW6TD2N048jPF10Gc7vAdcW0k9/dzEkRsIQNoQ3934yHrUitCqhpbsXeDXwfRD6xj07e
cVEtagCOnySZt0+bNcO1T6B8bdHxr02lmdl2HxjLDOO5LQJKb68tq4iBVGMk+dPhQENI9yRcCTdm
amLLhJqmF9JyG2xX1FcdeCgJVDvEl0gOGtf6DHJnaVUcFXma+X3xlUGsiWIdtpqqz+mLKkD8Of7H
uH4nCpHVkszlPbuMYAW7X0olemt19L5xx5L7nkM99RzvibdnVdg+fk8dzTQv69d152uWztJ5HP6S
Jx5nmSS30ZPGDWf32yllklBKdFSq4GiiZgeFnIA2QV2tED7naAcs4jmEfF3iedKhAia3GRxxr7Nj
pqs0N7b8RgvWQVKRds0v4rqDUGqG9TNn7KbPTOCKJIru+bVVgqmOLB+aqPRsP7wIB4q4icQHVDG0
J8C8V0ivmBsVpaCqkpMzEyOGhE6SEO2/ALOtYahZhEnTDAoIQXifP+JpdXPfQlP3sYdm3cEjc3VT
N3kXiz/xx8COXw0NK8Rmcujn7aBc/Q3zUb8dUTP2lGGoyTIS851Bt3+PLHUuk5y+ESwKCUUGUwRG
CE2cRspBg1E8AGq/j3JVDE4crw8EZdpuc719f4jYBsM6J0srpQ/0fUp/XrePpMW0cAni8zjCGO5/
1NAsBVdX36KeWtlapUTT5JLZ+bI6gpH1zY2Y4j8jqdeCpCLRW116u2/zP2q5zgCP2JVyRRuz7g39
30KlPWkUj7CxTPgeleUNTaecKCVOdYWVH8lKJDxjoUJPvnabGJ6tvmCukWEX6cZZ/xBGkOn8IC1J
VHNmft/k4LT7CzcVSnlGJKDHVizkCN+/cjCxzxe5Y89FLfGlPMqSmp6tolDiH62cAbPIYQYeGKFw
C7KTze3auBSF9QzY6BdFxsKnBFnUj8YcNRO4J6GZwN4O71UWEA4P0pfOQlH9eiqXpiiZCjJhR4eD
x+mwCblCMKRp9mBwOVBINf98acSRuWORmxUtfSgcCM5L7oX162eKwF1F9kSTHDt3ryQFUuhRxU0R
I9B/xvtIqj2U/eWFcAgAUrdsrEkGwvNQeBwQ7Rqr6m7Sg3kQfaxeukXa5GCFLPNfoISNiGcsg9FP
XjcY7dCcgBt4ErLcNKcKwANYb99LYMNKHQb1S5hiZ2Z4Rrg2cZT4JgZdvQzazJrQireqhF8X/wFK
PHsI/Y/sYYSOOnuxSZ6trbrRQoVWCYO7EkSijIX+0LRWjk4NaPmd5jTaQsbvpoze2u4csXvyKi9N
kuDsNhqnQb/l+hLq+VgPKKi0NJnEd6P3hydvBemF5CCP/TiQVWmYNVlczHQkN2Uo2eHr/nOO7avC
8NFGYA2Xl15bHtlu8ygRX3P4eI5zM4h0+GMjz4F4VsctcsEgs7n64YTKjG2wCgaUFd+jOZ09vJOB
NYdDHm7+GQOTt/G4g4HCxWvoYQf0GlWHdEMUgQJGrRNEzn9KlaT0QLNc+8joHxuOxtGrFH1+Lg61
gvX/JKv65MuAARWPIPzUaHCks3nNYSqr2Z/e+iPawoXymk2CLNv5kCY34PCNHtQ1BeDxLEg1Tad0
XA0Cr63E6p2ZxeCBVVTFBzvFGb/Wyap7OqbSNr0F+f32LXxf5z0L6B883cgI0SOBUAFw9Qpxf/+R
GlsyZPx8qaUVn1sVujrRq2nubE2Q7AOApnw7AWi79d7cJSUOz5jF4w3GoAs9K7XarZBGtSS63B0p
dBWXqHMzyhZokR+s/7zFgMFrqByJOz4I4guZ/mL8+JEHDbyeL+cmv025sEDTXzp9AynzqajZEqPD
3wCNOq23iOdnbj7kxXNtKhw5kuk4KyAj0bSmvJJl9/KgXSGrl5Aoq4AI1H3xrvJcpVOqyX0wpGgW
jh+AuU+wraYMnOjg5HvwpKGBRNyyafowXxxhbBR+mhckXoTreMAzwqFgBltLdIXB5Afhl5OxYA/P
LCkYOgtWvpz+CEyzYj8WFBl9WATbr0bDLdJ4+9gFp92rwgKbYFyECRnjWaiWV0T3R/S5innlOPh4
jEOJG1vT6qclLK2ronpkgCA/0kztS1T6b+kxlJLZIvB+YDonA/IwNP8Ul+lbeN0V/GWY9B2oQpU9
AZTC4/zfuqy4a+uVwPOe32PPAZGvIcmdRdPxUGz8wlINAAYa3ugWeE4FHe2d/RApLGa02P6Z1yE4
qeAPm8qCbjrNKh1D+yU6BHRi83jPI9V7Vg+kJWyBQvGOJMRM9mDOixz0IduNsQxm9bRsUFziVBrj
ud2v08bo51ndVnnRhU7EbyHfQBqnMUVVFVO0TzOB/UT4P340KGfyYyCbxLu6dlTS6BBzXbhXHl3m
oCVMmM4vBVKK1OtqER/hq1VWciPEKWWNjvvIuS9hW3NuVXQnBcIU08wq6N3ggrmwJGTKo5FRULr/
VxZKRvQ8qMyamYY7PMqQDQdysfkvma5emx0d17mLcTAhDxrspJXLGr7FTGzWfyFf9IrG9/UOjUfg
1ybPFDc+WYqWxAtY5MGdN5yGjfitJFnEmPEWQHGz45928AYJdiQoajMBK/60J1aQt+dxsiPxSbK4
qhiEXId9eCZdTVinNCv+ePE/MYqk1pe0u4WAjc9M/yKVbFcHlmv9pJ6khhspmyw04VsphjR67qM/
O+LHSR1V3oho7eYWrXqgIv1KzVGBqn6cLNOmpZEoGjCIQqFDvd3nWAv8HudGlsq8t7Fyue9l/dJG
oA+IiCVu4UPJTHGnrcEo5Q5enZiZBSyevSJNIc6NgS9wanLke3nj5yH3rFRMpDUyIk0cCpKQ9x5f
cWf6MvOc5f+QK0M31HZGX0ieaTIeDcClkoDE/LcAHLy8GLdaPdcJIpR1Hq78mcqwNvlqkUwUACOu
i86/znggUfJPGidKCz15AmKTGlO6eHB5W1baLzrwGdYIlSW78PWjRYrIHBDq9ulY2uIEIAiAo9S+
K/EuWyXpk9+YsRDw+/MaZJcB5q4JZvlO88N7Y022J7pKxSooeuBGlCrIEV0vkqt0K3ntnP3kDLlU
v6aTH+AbC9Ezbf8bW/6ThiyFflC9uLYa/dSrYtcRhL7xY4RZVnEhM85u/YU5X7CtlibtFVBVts1S
kFnS5Z6fPH2druHEpMfvaBs4bp9+W4rNEjJy4SXBuxOKvddWi2l6KyOXLHttqUCywbxMlu9jG15S
LRwgz2zPnTI/e0TQyXIhVsGzVELKetzbVI9c5nV54LDdsMLDy23dLM545OCEtZv2zBJ0b5qhtsFQ
yzGFz904qM793KX40MPfbXDz7wQMRU9vCTzpxTpEFSSPIsj4Gh0FthLSRbRw+8ZuHvVYpnecRPRN
MGUFZjxkPTpyG3g0xRDri6QoD7VcvhAYz84EQp+MUr/hc9SRBHedvhugnEKpM9QU5tclaaOjW1I1
OWGvB13MRHagzpuW8NPhNhkaLL620rlfJbEUL7ktcyE1YAaiGQoe6sAgrwJmEIBekJNBsViMDdAZ
eVLikoS9Oe/bLTGTptLp/p+oJBdTQSQaPWvkNxt7mMZe2AoGCV4Xd+x61LM0/OCUv7wl9lE+C8lU
dtnXR7/nM+RmgqS/kjyt3JNIlGFE/vaJn4KZf8ue1ihE7QGQ6k6wJUXj2cy2FJ+wj6cB6G5bLeVH
Exa2AcsUR9P1k/yI7cgrVgV/VKq3OnqdicHiAqni2CWT2NEiyLKmjPUm4kqKJw78rhl0riweDBXj
wapZDG/4vLbDODqXfOEjoBa12V+GX/x52q1HkLY36W2dPOwJIZDhdYhXrvrrtWBde79pYlZh0AQE
q0j+nakHmd/1iGnN5QbcorZD9/bbqNmBf3K1+eQFUVl1eTNc/DrrWNmyLd5P3oEFBL/5N8ktRd7b
7CdNgzgW3bSPtxvo7T8jUE6KqfU6F1FH2at9IP9WraZmMfsu38QuOXs4eGiOt0g10fwUKQq4Q0cL
vatgjPP+w/x0xi4jkYwGzynKwyFKSVXjfXiDBqkDCl8xjJy96QLnanRquJjntVtN8rRaiZHWVpAG
v1CzhRtwvB2h+ucDW2VIy8O/U9bQ7vd+85qwIGpGkRgqc+ISthYEUew/ZzvHuHdw2Y6N6cSyQLjU
0tV1Es0Yv0W1XZsPE0TlOPWkOdYwBvwevxB6wyDBXNKpkQ6YwoClkNVypunMTGRmhl0EJ9FBy7cS
KENTnEMhCwVuwyhRC3XPwOz0ezfftgLofkGi8fRQeGW3JXclJEDZ5+1R/9UDMBo4bGlA7TMsTJn0
ferBVe4Z/dAEg9Zb0zHkw42s39FZIckT4QzYS0a5ehJMpVV96xNooou2fVDr9t6B8Rob3y5aqkcz
GVqAH7IoqD3pfSbGE/WYfL45V4haIhqQPj7xxk7uZxG5tcH94LSPteeUxbr4L+U6/0Iy9Bmlzp5p
lJ3ncTl6urj84iSc7Y4eT2qNZSCGRkTJGCUMkUrxgsgTygRM6xrHvqAAjlR0AKvuV1fMugzJEBas
mTz+WEuBoOtN+Y/lPyNn2Pyz3PK6Tu5yUnEfP8kWbcmTrOZ6uQbQHt+RrkSs1nlXwi6sx8SbsKZ8
nJlNFmtc1TOgSf7u/n7r4lNt/mftVdTf/oF5v+uhr9ObKR6rG1KbS1Ml2VeQxK8iSRdzu0O2oE7D
MaLGJbbR6wCUrxteIEI8BeLYAW53UQNXr87RBZAsZwq7nVkiUv0og4+rn6nPdx2dX6IHmflZ1nAZ
Y5V58DdvQ6zMnyyZUMr35TbEwyn2m2ZcFsKEEFmPTxlGxxLdMmmLmk27Fo0emYMFOuziKQA1evzs
KHlCpANbN9P1TEvRtB7Tw+VQMuSFbcqBqWdK/WU5xw/ZcsaFO+YlEuA4hHorC4J5RhRPQpMoVGUP
8RlADHd3bHDAgBszjid5Nk8EPEmP5aZiKTFNxpDrxMqRj4RxZsdiXNlluRt/D02eAnxqhRFEr8Re
gJ5IFmmMNYSkD8T4l7+x+UIAdybGyEjH0zE4MeiS1AhU2evnYsjkdDUoBLtHe9I9kqSP+pl3pnPc
fbUwSm/XV9498XW8rCT8Vn9mQ5XhyhwsI/vq7hygLbadatI+DMT+Y99bKVTyXJFhpjUKdrtT+KER
quXnFACdGipB40qesxxPmuDMWRk4DRqo+a8ZMZo0xeRC8cpAWekkfTLNNAEDPfbzBYPBg4VrQQzo
YtTV0nIesYIkEuC7TpQ7KrACWiiZs7z1A8h/gl9XnBGJi0EKdZcdljeMvQtr2hcuAoU/+Sw+lwr1
i1mTi22U86NNraAEhM55jDII0Ug57XWYWAnHoijmg7Hwp31zU6Dh/aMbbjdVibTcnD1q2QLTbsrO
zjyUV3GA0zj7wiyuNZ7TOFKfYNorZ1E7UiT/QH9OoIfGLXkOaCGbchvwbk9/8qo49p/CcFBt6pAA
MNupwKjZOU32k+Qi5nPXJSVvSJ05VC5AITnxEsEvEfDk4AY1YoQMHtLGvehbj1pzv2GwUfj55f7x
ojWi8sB5yPv9BciT7zDN87dEKTWTDWtWBdJDrEkTnCF4Lqs4+KUqJNmRZ4Q1Hnr0V0owQ+lNDeON
D78ZK2HOI5AMFzHeao9rLly/3+teNZZRZ5BQhy4j2tbK+/JDj4ZHxz2oT2nmz9kncL2R5ps0tQCA
tTZS5wQ4wdcNMB5yy2jwDBN3kRhVc6NYADnLzPkBi88E/LR1gi/U+7ZytbcC8A6ZmR0IY6HhN2UX
gIWate0Z23Fn2OFgKip/MpCP1JA7K9N0aseiPlZ/YNPgGxkksobsBWV83RVUjJikZPEKVZBaHfPL
9PlcsVw0g+9MyK86KyOTSIojQ4k/dnxNiU/Ym1nsfcqXeHRH8sjxqN3mL/0h5edR0EaUBy4QgIX1
NO1c5oti0gpqVG5l0hWZJknpJYPqmzXK385CX6pAT7cV7r0ZCl2OVJmbUx67tciOoVGjdPzl1/t1
6sWn2F86NxxIevTJ0GH1j1KUYdhm7yVpcw+mblW0/EGYmVEdpROjuq12rGwdJ6pxXoJE1qE/G0KF
+FeTPcR4TgkD/CSl8kTNto9y+R5fsCipijW+FFfR3uvT8ugmhIZ/djC5WyVfcOdVR/krEzz6yftS
t2UhGXNxKo4BjQWbgi1bevrk4RuMoBNkE326EQFm8YX8UuB3hNceMRvOxXClUc7G49oUApiRIU/M
jOh+9/CdAkd8RbRYAhp0KQLTvTqCNGcBAtlJX2Di4yoU5WTbBTdsHT4nNWy6qQQAV/guXlhJyPd3
bKM8OnYb9sfuXMkx/9wMCUBoMIte5aEtpmJwPzJOUAmC/1S9hbKH03MvKiml67exOBYfGNVPwEJd
jbHTqAPFoK5f8LkHWKJhcRe2RHk1AZ0AE9kSASbWyfxvH05Zd5p84i1mmV5CB5mwQwM1M6A/F4iE
u1ff/FHQDPNgU2eUCOmgwOHKU89mG6CjGVB/72wXvXHR/CD37t+cSGydKqFWuwmnqXtH8DXsaof6
eaYuuxBUwcB+hw0biT84uNw7K1jffSKNJsYk2wXJveDpY6xI0RVn5LO6d0fb14jkeXDtTD+cLcq/
YriJlQsmg1bpht7WiaZF1Yb1baxybBxnuFBWCej4P7mr/8J9FtD+wu9n9TkR2+Q8TyOmQENbAMnI
8qFY6nBEk5T/UEhCan4AuSNtd4K5T0DvAMU8TKV8QnzsDU+epmvOv2x9JgXF8QOpvYm/B3fh3kCG
04VkkuuNjF1teJsTWGKxWRBFy9oDrzlDXu8yYCg8PfvIma6eCoOwrPrKMcWTqg5lbiB0DftNqy1Q
mtR3k+XsOvgMlq+6NWdnST2RrpQSUxojsz9Xzs9fr0WWf/zBmfZm2xzqKOSn0cOJMo0ybB+g41Fe
Bi8PKQelTHrw3UNWJutuEMzFHQqV8RryWGvr3MxAi5mgux7IvknUNFSGIMFIG+hmUuTgmMpYlHyI
nPZSv0uWhXBT31qv9i6UlLBZibMfcRD+ZN9H8pj8dvPSl+v2N8HoHVnYtUD+a2xZ4ZoUeSnD9fSS
8fk0ZVlPghsm34a9fgLOdJsaUtpm3Kheuq0twTPYJs0sRCigCG5gE+ze0xPxPk6OeggAZs03lcMV
5emyO0o5lYdFYr32C9oLa/0tYgkwxfnOTxDcRXgwayGXP++/468LrJTZLmCzT/r0G0tsNwVbz47x
iuVfFH0qdoz0GE+aT2xFgAh1nneLxILM7jny7L4rui6VYRgeBmxELR4QZE+88fPZE90Ti3mhNPvb
Cy4IJF9xsUjWYN39VoXxt7+I51K6ERYaPNoFibu9LGFZA4w+FpOijAhx9wQBfDJPSeSYEFlc9zpu
OhdL7vJYpSzreX/P2ZrIoiLYfuK+BcslL/bYzYtqMXWcuKUaQFVNaJrDoMezkzm9V6XGVuwV8f7p
DokiqzOsYo0OoZkHAvWLRxZJPuLsmWZUeFDrnAKslqqyfnItCJTa2j8TxdjcEWfXYY2TZLwe70ax
qkDj9ALpTw119vgKzqpi1koVZB8i2pQIg0MprZBuowMhjNJcJTpZx/EtGao6iSiy6QcoTcTzkGNw
BoaxCzQks6KClrKJbg1U1BAZrBSrQW3FEMrVimOHPC/70W7vTEK22CSXt1B+kD02fLHBD9dge0x0
uRZrNX610RwLOcFz7CRd6LhpfJKxYulOvk1tHDJ0S1ghQuNA5NOu+vYZwJvzaIcDLN7DBnuYBngT
VDAwY1tG1y+ZfenjJTw77BrinuSVqHDZNW+/ApyuecYx1ElYttWt7R35LXT75cqRnwF589xaqqUM
5BXlthPFJrkAhRFi5Jsq6wAA29TniGz/0McQ1DTbMST/p6lqpCjbwcVG+LpNvnz0qwEk+xuMA3Gm
7bXfWU0hPuZLVVXNlgPJEIm6HMLw7PXj9jSMTFnVYDoWbcykIwlZqSTu0ROE88UhKbEjmxnu/VTz
E2pnXUbkgiMp3A+xvk+qhH2arRVDJMyZv8i8zC3yJrtS6kR+/OjtKYfEKHPKzWVDTDMt7p0NDQYV
Vjb7go3uegURb8oTanwqFL9um1e41nURn/YAbkGe5eflH7wZ74qSO01zC4jBFVx6+Z3DQJnSXy1w
b/xMyXIPpIynLHLfvywNrIRADMQXQmGMVsnYYZE1OTb45MQ2zX244nIpoCrUQUPUSB4EE/iXrPvS
dAbw/JQ9abRUnBMtEWWlUNQ8SVRcmB8k0o0KjcIbbeX1BYeevNT4V2mv0GBFhX2htQ6X+3fyZcyI
HFwJDiAYz0RnYwxEAKfebLpUqdpNk7PFw7mLw1bL2NHv4FJoe1gB9UdCuQVg/+h9kJLvEa4lmxB7
4BEFleLrGwvqdQDfsRgzKNb7zPDZZlGQ04CvOYA6QkEmQTouHHMH4ZOmdN45z10gKMwbbyl0MPOT
AxKfZT/Z85iZ9HLi/OpcOiNiwjncMn5ZP4+wtkIKyxd+wKHceC5H/rgJ/XlJFf66hx4onDmLVI3/
Yxr1GbmYwPndjVtfLOeVzi9kYd4yyGpUEAHastXqddsMi7qv6LPmR3l0X+qyTIWU1F9vuWTm8xNp
dJmXyvrD24CujxyW+AlVa0cARRQ6rwZNO1dKc0gv1fZsYhm/04xtAKcnMw+z3cvuv/nGPePEhTui
3jrZyApIq7X1GRGpkf1bxfD8ECOoV+DavpIGeKZW3V2ngHpRiplOqiWqwNf7pInPBlE7hQIGNp3d
TvUQ6HbfTzsa4dnw3c4PGhjMPFt10ozFJYZI0i2fxvlNM+d4pN2rBgccrGZuG00/ylQQewKoX8A8
8N1KT+VR6cFLW83gmRqaEtiaIZvmmNNVepfqMDF66M3RfFftYil3mJfnnxVPD5it7iCT1BmlLEl4
s0ks6SCmVAd7Ju77l9Ur5BUgjeN9VuWRx9ZYonNFP3YeKt5G9VpETMrl0P5jGM1id1GjfOwCr0ou
uCEsdvUo1Tn8+7F5vszbWYiGXe2gcGwzfg/yc/x3qwdke2P7jCh2fk3Bf8Ek1EAUWAUeW0o3NgpQ
MU+nq3d9vijsQvw1m6FETydsZ3W/z2oRbg2BHyWwHboIIKaEh6FF204TgYB9q/ezBkzw/j1HRUU/
gadiC3tEhUz3BdmsUmUvYNmMnsXcPThSi5ND+V42vjij/4ausHbyKA33Xv1diy9hqhZxXjuJ2+3p
G3Zf+C0EbahqI1MeBPXg3k+QiA/deZaMTSxg3MIgaIyaN9gUZfx1iP2yjuC0pgkd+0cQdteyok6G
0y8eJ8COl/hhms9rX/uyL/cz9typDhOQFqU9q2dOPG4bE7Px/qBkIOAEyNlqNrhxdAZt671SirRw
9VkxlsdjBDUfRqTHRZ3nh98gVgTjASicCAZDRsbb+k61vlzuY0EHLiQLKix1qA24JI1iEk870oLb
afIopJ+CRb2Wby+8F/P+ak1LbZow5mJtJmkOzhU3g+r7yQi/HXQQu0mnXr395G0hlVJ4rKcIDp+B
Ic4ixGQ3lmJreghE2m9mvWclnROwnYoNWL0oyvzy0p8QHrJj6yas+HJ3sDB/cG/uhfnqm3K8TzZb
fQW3gl2evhp9FYDRb1UerkcC3ejiNYDsyzVG4ds29/Nv9tq6kkRioTuyZ4vAUDu8mnHtluAuJNSq
GuaNZuG7BdndK1157OMMhmqYU7r3Pm0fV45m3+bbI7zLOyijA52rpfEUicMGEqH/82ppbrPe7RGr
mM48zSh6SzvTCFI1YmyWipo6mM+maFOedh0Q2bwa94iRX/vs3YB8Eyz85ZxlRBZ/u3lCZgBg3JL1
mFfPzK2ZmJhU8ISobUTSWRTQNtQpJfN7zBRobnfdW3wEuBA94f7mEHUOodxRavn/0zMZ6Ynt1D1g
XZm220M4ycq34yGQWztYoUI77viCtuiCPsJT0FXVjHdQsx1dXoKnPKb7uVu7XFbV3YvbM4qxcijx
Kr1cP8f6RHF76CsTP738vfuLBWkq6Fj+ILx0uSSBLQ7Ynk3HBbb74SyhnGlEx8Jnoabh3l+WlHI7
XoGekTTEhnm3axKSLb916n/nytioqpkBQByBOBD2Sa0FvMjF/4aHiqQaiyYO9NwLrEnj0tcw+VeV
t/Mkr6cuiVKGOv/9XlS+W5SoHHKXj0KhOYvDpfFVpL4Jo6H64F8sYvilugpwG/TProadYGzXiyvd
r2kv0/ZQevi2bUKC1KLCGqS+qno9rVwFpFTWfUxokZ0sm5NNFfx5onCBPjC8UXr9DnHAQRXewxth
mzHhLKDW8eJlgRA5uLRpca1aD28O04+n/8W5PY4xQdPF4LOCd/0NqBjt/RVXEBmosqhsoJVI5w4X
BRlbT23N2S5Eq/qD9WqJLElL40xTzPkQ2o8IzbmXb3Yv48uiDN6651PHK7/lyXLWtgvNdvln2TWg
nGjGmZg9HO+3w9KsRkYPVtoEHwjsk61oXUcc4hJG74e49WLTGwWrxBLHAY4IgxOu7eT66b/AtJ6s
oereliFAesDUDSkxwgj7ggdIKVn3mzvFxdgzr/vw6MqksI5Al69d/7PLAvCPdzyX0KFlP5irrUl/
ZxPeXXS683LHVG7KCp5dgdXS/0zOQAlPauNNWtS1acnlA2+FDGVxFkbF6zdobeG8daLxGJ8ndi32
sX/W/Y2zHA8HtygWms8rnp07rj4tUWiWrZaC/KisWdi+XFkiMr7dHvykV/r0auv/D3DefCtVhuql
VvHNStDk5QaEW7Xvlk/cvqS5y7gPBCU9jUDjYEm31GwiULgF+Dp1I6UpGbG+FW5Egqh6vjeOpn8n
8VTyp7yMFKgBR1aFG7Q5Ld6ExqYkRX6XfqEZZaG99D7mpU63Alq0+UWUW/z1INLvsqAOn1luYdrS
HeOpptoGaJ6OsrM12vFWrXBW2oN1z58YgqubQVVm3MD1E3ROB0QdMxRA0B3Wm+IBsWdXe2YfLCvx
3yKMr7reDjHrF/EhwtM1SDs4J+o/qXss3n/ud+LZ4oOxtUAS3Z0gRP5/6dAOxzoNDOOrN2mXBAYV
Yyobikgg7G0TVErna9BlWRxZwfNz06nb5JLz3UuQN34EB7ZSf6wZ9qMmckxdAuRgaGe3j9g9rinW
Ya++VAdBSMTUn8x+CHXMYVVIhGsHAj9BWmkKK+pN0ll6BuTMpRIskTxLNDp8C8Xr2CwSc7s+sWcw
EHhmz2gIrzih2D0Cx6VyDwcddPGuk79X2DKbpSjtE+AAUqHXJdqkw8sS2yLzibo1r+koyvleY+h7
O+7tNMvwUz1rY9S6JhGkLC0DiQUHIftK/zqPwB/Xr8PJht+BFu5zMG69gRO47k2Q/6gnEKTD0Ifx
2yv9gpGisHXxSaZRMQdz6WmeA+kZjkcjZWIC4jvGMGZsMY69WbiIWirOeely+3wKSsXetagHAZnP
0HluJbsZ0RECTPwKIC1C3PpMwEO42ADUSBavCvXmxT/zUOLr6ahnVzEL37NbciS+Dmf2o25mg9u2
e8eP3d52xx9McJS0lo7FhMlj366WwAcnFMG7KNfIr6xzAABPxwtGDzUuZA3oRe4FDTMtWgIlnnOG
2xC1F8cnNu62tV33UvaPm2rgF2DO8AkpKtymWC4bgukvsmgDmhKWb66U9otZ/sSFoH3SxMFtpcdA
BFrvmb4Xus2wi3AmkzB42OjIlqoG5vvppZ6OVKBwnSW6vdNYbyFiVy8PCZ/unHQYcNoogEJnz/hB
ap2v28O2ie3C2rEunRWBDHjEdgREc+1jhLU8RZ/t4gFKdDss9awSBxLwCHfWAG6EvqyDoaYtHlw9
Fd1umoX1RZI6wpIlpyZdf+a93qJCECbUDDtWb7chMys1U3mQbfSUZ8//iirBJxzMfUlOTIl+v0eD
nEulTi+aTA/3lxEOkL40AOYNrHV4VS+1ahRRlaXHpJixgCaVDj8Rn8oCs1+BcjVon2jn8fMEyGwM
y6s2TqcD4FJGUAu540WA2u6urYPHsTaQMoYu4aA5rzaYGdcUo37Uu9xncXHJzv8lftydoIfo1NCr
hrMmcuetV/RX2ztGUW3/Fco4YVwDg4kjpDO085vk/VbwJ2YeatfQD0vat7E+B9IL+bCcEKetcFYl
Ah3+zf+U6V/eDHU1g51IEH9gqGHSAg/OTAgQV90koRtg9fYrvmO1wv2VwjmE1+8+u434YVO9Iyzs
kTcQCjZPZuqq5EegOzL1G0C70urhXzIaqlpyJBD7skzPslJ7gemLXBBORKV4xyzb14eg6ZLxBpaB
TDXjQM2p1XzFLdkxuXubOmdeNWbG/7GuWlP9ZCdvf0h36juJeZ1JrcUy+htvJtG8O7g+c3lJpkaY
Pauc90sXHKA0Q1NnS589y6490ThPrZvWONqfaXDMIfzFNHcNt1blHIjPyaXFlaNpFVqlRJEpZavX
ZncHfrkEgCRnkaeos9M/9vCoGaR6wIxA3VyFvs/2dnqPRyL8TWTTQJvtJIp4ATFIVvkEbOO8CeCd
5xVG5soKOhgclJP6HvzndsjMHGeaKZ5MeB2KY4O8WaMzv5iTqKuEAANRvQ3xxUiQvDUc78VTuzn7
NW6ES1ITT7sjTdi1oHcu+vSp50zRrSBQ3afX9Y54rzbhrYMm/sF2bgIiFp6Oc/Fzh162vfV63XWQ
OzDTiKb1Tun6CpQd7W19KsKB9xOPLiVJCl5RCdqY1CLf6DZ1DMsCO7HzaLVERDHBQw+U5GLeTcCp
mqClUN86elVSoJTndiSdkEsv2Z0GypNIFAvuJJjQ5m/Ip7pM+fhzf5ZshvxIxb5EFlMbCFfH5S+I
0RvU/3czCEi89mlLevZ9DtfCbIZ4x+R/NFte1ygM8S1EoKQKcIq7Zd1aAvqth/phGEfYVYOP2//0
1VTciGuPbjMu9QBUz3VBrpX9fS5X/rtl4lNIt5djDbIIUjv/FQtflfnTqo+ouLWXRXM/R8Jrg+TS
HfLwTfY6oOUm/0OFjQzfKq977gLM00lRKa4g+KA9L6OHPdBzMB9t5/DazzIzlKHO+Hr002QRigD6
17EBkAh3cNbZ/XWrjFyYg2wOeqIoWc/n7/a4mkYgH+C9R2UfKORWpB66U5x6wNS2vCRytKDqboCa
Ztb8q5xDepxzKT06LT6kCBNNFNhGCzf9LvFGNymkoT1bwiUedoqveefrAV8F0yKRXOgb+raNRJAy
YRvb2NVph4h2uKUHg5soXeBRoWYBU4ZdcAqFfpvpVsq3ug2mDfS5A/cS7X1lleJnLr6O4kkNLcGR
ew4Ml2mqJHgKXae98KXkja3UYBDEP5ijFPo1MKD54sWNmyWeK0MXnJNohVvge593UxUX1/Jj6Gz7
uljf0osoH1F2Yebm5sV9Tpvg2dmPnFNRU0/YA0X70pwGWIEHB8EJXVcCBcOtyoiUDRqOIx+a83dP
1uhLD3imQx8dqUJi6YLKf4v9ORqwB22+TOZths57qlrnE2NH7u2jJxd2yr3j3MO0IBgrDVztnCgr
hCx/JYBCbwD+Pq9EFH7KQ+JYYfPRhSCXWlPF9PAfbS7jS9Zv2OQDKwL/YotjTEzAyDF/vmtcNCHU
2AgNE+UgJGifI8oYXsUZm7kFv25TCRbYvbQrPjQVBBVD+fziJljpJ/GTChVh9213D5VME9M3MA+m
HDBCek/IzB34VnS09ZIHlBtY6ntVlkHK76/mvLiJwsE3o6O37W9FaPPWN/Ave8w3EGH4MZKc6jCj
VIbMZVmKlVaw9xHq1HB+C1OA6rYkiLRMilGASOyJd6/6Ww/IedRSUijrbxpeQYvLExL27k6bj8LJ
6ZosuwMbHzRjRImGQu3tiNjMHYY+rcioUp6zgv7bDEATgsd1AJLNv3qL1sg0eh09g/8kMWe1Dcx8
k44junpn/hrKN1M+jEDXx97esAIhc/Fv/E2VtqBc2WlZpSN0Fn7ehz/fe6y6ojrRkzHVZetW2kJA
i8H4GJrZFFDAKvW3Fch5ZKM187LlhA5a0XMt1BFrULg3h1aYTm2krhLeQu6lWVJ7bY0A0j67oDQv
aKsTGWHqQlte8qubnYX9b7JZbQpaCN4UvtPQFNGkoPVZrGhcG+fdZymDelcOj6oplBzz4DayZ9f0
rqKzaMtJtZ7Ho+RgbRIRECCEsB3sffDkdKYkQ6T1pc1UA80oQxzeLKBbia9FhCpT+g7LLkOiELiH
dpG3yLYD3gB81+IuYWAsfekXdf337C01pguZuwtizmQtfFUqLwD18QJA61Ed3IkWfiVhLLJFX4Cs
j3HmSMhpMQ/UbpTvP49z/8I5WUhv2FGBcIJUKoyTBGzXJo+79zqRAAa43SpK9MOT66hld0IdeaN2
0Jj2POS3rg2KHA0AzrUtroUcCVXWbpBsgYkRJgxlA6mGTRMkvf12Ih1lu5Z6LbfZ+RCqGLzo/vZ1
qs5+bDhzU6YYe7D9uR64brVO55bgct8XuwOk3verZHf00YrmzGRSkcw+sCgzfeqySOPDJ0On4t9B
3/BdFGxZCZFuO0TepRogsod4iphbURnRHwuXCoULp95jV4JCVuMbj4dXO1QozaX4VncxDPN0cIFp
GQFOl4rRnWGY/hVCr7pHfYWLNwxnx83SE5hcCU4x4IeeEmFPW3THvqXaqt7TLrQXAX05w8eG/Gl3
tXBtX1YjkVJgh4FMYdx3Z3UCgvST5GVvmGCzuDwSiQ11plTln70D2xwJclGILLJP+IkFtbAfqc83
5Ka5iK9AATvFbQdt/1B/45W8HMzrEdvwLJ1rKEwlX88NWqgDOhmWAGIBGEYJwRNTSBtQyqdIA1e2
oZv9CLuUBL7SBbApk+H9/o/UAF/NlWisvqBrIr/cbNqYyqg3eJ6X7idnsuCQc/o28JjC58pGFSac
K4HNyH2/oJGBgbV+yqOpNtudo6Db8EJGKbgPe+OUiKdwnMa1FnlyuzcBXvSC9jjZ6O/SnCcxPGKo
eF3lQwjdHQbBHhc+uZhF5Eaw5qeOgUBO3zXh/n1LhIKxSRqrTk71Q3p7l3s9Uut5nFbF5e/8BJQb
VPWojNk8ah3d6DvmagO7VpYztBhJUx+/FSEgXVW8TEdPlD6wVPV8D7vAEp97SrP8lwKsoGXWEDsc
4Ly9d09yi4AjhHyUOwvKLQkzUfQF+iydhcjejB3PX02I5TNa4lw9XplO4bM3/tNcMr4HLnhaxQEl
w1tHtIXqb0/T+01NrZZbUKI3+sSko4d8OA2SX15pEkXjzRfVBiRwXS5wAZ8+Gt7DsPsDfHOySpud
i42ldZxxc6TAjI738mVyEG0Q36/mq36EcDk8t4Yk4rRUI6y6SRu3UX7tedhRx1xe9PuQD2W4+NVX
PMGNXozXlUkmLnFQJFee1/2p7/2BF3ZrAP/7jPuxLYDeziHgggXRwtsFK9gL02YmlnAU7qPveQKV
u7T4byQIXUXCyXeZqvqIM5HOSP4fkr8dfg/2G1goY0gYLGpJpSu2Ji6TLhd8kQkDNnNrAXgy1Bc/
5cLbVvwVU7YRHc2dLpVZPDtMTTRDXGigzBcG+iSK8XgEVRMosHIT+rPyicemARvI0hd6IqL3qQoS
zpS/JercG+yYIgYWTeEzz99acBSUknRh9QFe1NFVOnQPHt5N1YMGsQomLMEuDp0rgH2ClIvsHQTk
kjDIdxCQZqYoEVJzS9fxQeZ4yTxeqSH31cmyhmUMRb/vw6DVE9G2Hm9kNqWfGVoRWLjMPc7vQTZ7
xLrHPOG6ZeCPea8kRztz/rj6qvkLItKpHqkITxc0P0216GxYX7cYeAjlXsKWepfm1XUoCkgKMxLJ
cpadb6QnZ9vEkW42GMNmplgM3s68cRHLIiMLckzerV+d+LODT8ymJRX/lKFmmpIX1Tu00/wfY+bz
IM1ytD5+kkbK5XKqEGZHmTwH13zSm0JTGr45cBCUPyukkuj8qNHMQ1qiJaSX9Mp70OV+DL85/xpL
ike2783ZHldQDsJuGBb1E6x8g2/G1eAbZh312pDi5Rxn/yrIQWDolTk3QgGiU689sJavYHRN9koX
Ec6xOVG/YjfgitQl2cXdrFOpIXULBWS+WoVyqIaKZHtpRwLB/pvkZ6JUKgmtm8BOTmC9zVtoaZ3B
QyyWt0bhe2O7cLG3EPRGEel8f2xtuoPeNKErkDyWxC8qYWwrwTeDrpLybChygjJRZBZim7O2BMnk
HXegrnQc3sU8fBl6+/lH3lOI09ioNZb6v2lJNeiKdp3xq/RC2pNUzaRCpvskyPGp2v6UVfFyjuQc
N1gDDelhlwggmYjGpmMhc1Tn0TzIfOcB4R2gxxQEhHqbZSKv9/ijZu71cuk07sixqlSqJzTeXHlb
y0kO5h7mVy3F17/sBtMxEXUJfegFS+nnBYaUOPNii2YFNnXXB0ho5aM9DF9izASuf1Ui1InU1ZwD
p72QZzh1FnHcDu1gyk0e/YFv7W9Q0NEv7uh1BhFDvlAJ4K3QcuzoREFgbrWJ+4Rb7EznnSpLxtyY
4JeIgqhrQeamWrPDQbaojIGvxgE6mwpGK1wKQs8BOW1Cc2wF2IZkAYKKOP6XoIjT8ATKeCdnGQnK
AO6e7XCoQi7j7HCQ0eGZIKztHrH2foZwEBKA5A6onmUh0zGyCoSsGpbuOOsxYHg8yAPr29cfVr7G
HrdJQLPsXvH3nImEL71JFTpGP1fnmfw/EQKsqTWkYikRLENsfKYgOeTphCkW5WtNVHv5iO/j6LgW
HDEVYIDLsx9Pd7fKqL74tbOKT2dE8dzju881og3BD9GVCzevvRf3RSDoqE1E4oxRZSda4oHf2LUQ
PDhQBoarbKW69OzluozgzQiM4nK8rtn/WE4aSsoka88wwR7p4b/x1/VHSz9DssQVsBlCOx9lOJ5H
iuAm2jZ/Ku2Tz2QIhwxEeSD4UK2hEdfZSgtnOripRRnb93xmbG02uv188RCotN/mX4k4v6pepRXc
Z3DjeP5GaaOdK3jvcbAUB0P9q7Kz9LWoNgc67hiCQnlO8xG+rsOXdmMs/1y3OJCgAcM3GL1SvMn1
3w5iGBc+5fegw2q0pVX+UN+mU2or2UL7lxR9ZhTIXNFUhfOroXI0pxZPyUQ1duSSxjeYmCdNsOWu
bBC92XmBT+gazYzHTD5yjPdrcZU2k7G7a/Bq4aiMeC56a8RzLZhW1lm8Q3tWUP0gnrq5dSh+oQ8h
LrElkvNtmjTwSd5VZVcmAmHrqys13ICGDBP7+49V/3cl+6MB1PFQJ7sSluPcWVWxQoD/Swn5sSAF
4i59r9592BgmUTboS/IemLHC3eHTBCMC43c/TYepFLXmFHXvJ5+vggwyKKtfj+cVTHENJpIdIBaM
Af4p4lnqquLkm6JCK67sMoCAn+qMzPuMeeLcBooo5SvEB+Nq4hSE0FrWz0Xf69fSDbuJYkqzH6la
/GtMII+KFdji6bc16PH3nFXRO8+BocQtcH92+jUEGRCKuGJv3UCe39zHgFwRwPiDmx1yRkMNlC5u
cF/eDBMP3NpL4elMff86aX5N7H/sG0lNh6aJuRBSHUDj6TdJ5k1p/8tEw72mhZGdsoAjTA1YJjZg
x+mkhCxUVC++pRjPfg5i+5GlcmzkQnJRmd7Gj69/WCHFkgov6UrRo2H7T/JOStByqGwBTWCGE34X
2H6wOwBJX9ekwIFhzNreLRDr7YAaPklyKoG+u+A8b/SGbRpdhK1HNcKLflVJZzdxvMym5Xzhd3Z3
05PezT9hCOUlCH2KPoHMjop94v8o/C0cfm8Gla3bhuVJL3HfpjO+BUQPbwgpJt1oELfDC2F3Kqoi
L0gAAiWNGVkjxHYAIIk/KeXKJJxvVZJ/S58xGo5EXNJR0GQLZSGTxuKBY3nYHFOrV8nDf1K/shUB
yFZtqflyy0kKxALcUxAtBunsb7IZOGYUcc63Xe9hQG7vOl/pd9pJUhOQzGoMmHRU87uLWlW5i/xa
HWZALgBU2qYa/BdRL+T/jML+7PlsuPnVkWRXTt0tlta1c87p69qe8rS4SWzDSp9g+dTtsXTGKbnE
0Tsx8blivxSsWAd9l1qXDS26Gc2sWCk1lE3CoanbEFOSUyxxe+NrgGCr0zS1EKPnhyY/2DVdG1hf
+72k17YEn9HPWuT7hYvBcZWdwMIuldqSjuPjiJBmqjzXj+8y8uxWTZyuigCIj8fubCoJyqVcxQlu
+RDOAfCzoBaBMMb/x6dZQed6fzr8V6+P8l+m1BQBuVHz76/wqxko3yNhbTZou9grOeUCfMz5aTrF
c6ttatxYH6gdSid68VkPVDriL3wouKN4k9M1MLXucsvx6SgAd5bj+7my1PaDh/yYHMronjrhqEvz
bf0DSyfdT1Mbefo6zXTrLLhC1MpsXVzUrgHLyyYJgE5TYE+QvOZaqlKRYRqFelwekr6NnmRym7cE
8qRtTyNt5dMZDtYki2gxKSt5YwBuLCt3v3U4CwqH6FonzNo+3XwaJrhExl4jLdDdPZ33juvSTLCW
spaRYQeScaj1g6xR1UnLf9tfj+a19p4qXup0jfLPWHBBcW9jIKr6A/yaY07FxHfFOW+SRgu8riEf
0N3+Ayo6coi26pEiA0ucleFRHWcO6+SENlEik+gmq0P4VaoOBDM9sx4GaOeHbs2d5tIe8Wnw0v8k
hZplk+59kQLtT2nnrtw2cT54mIzoeckQOmxG0aAZFxAsXI6MVwzNLXl567nU+uBDruBKS2QjEK9k
7moiEHfr/johqtJKEqG/mLH76HaASDYNODsFpmyWb8Ys5gmBzqBAAMd1BMwfJEvN83KfdfmWTADP
eNNprzjNIWg4HA9Jquw9gL4bfnXlu2EjacoMlXscypIX7tkZv1Dho41qE6VyC7aPpR6XhcPvT01v
6YnXp5mMxNzKB8Cp5VXRx2BfRjRyBd684/E8N7lGjGKmOuU26ceO0CTxcDc+W7LqNb+zxrv7p40/
ZrAF9UMlQu9AXcacUHsSCdjmxaMpKvxuXdIdRhT3VtBqJbN6msuiyDr6K5kEBVW6Tc+BbB63Lb3N
hv1o2zCkAf94DeNp0dDWPFQcvB18rYxOuNgQ7zTM+hawTmcOATN887RvHRuUr1Le+xKvN3EB7PyD
NwloKlcxsUJ9Xgr1BHoQt+v4BjrC3NFhF/z6gFxc9+GtnOp3+W6melvHOt4vBrNPKHWBKnK/BFAu
5egEdkl/opxTVWdIHIaODx4LeuPhwYA56Lz8noew7cRQdRJCzRIfKuEpBapyCU+jHgZh1Jw3HXWu
FMQ4Lvjlzgy9MqUGbbThHqIdYXnCiR4BD1kfKG0IGvB3ka4a+UkgSj+cdpNivo43IcKzNxo52YiD
yVG7kLW+SSwj0Pzxq/PZl0NEKS74jsJMksT52wSymXWgfkcz6CLUUPRUOskhdnSLjes+YJAaaH9K
AEzeS2vOkUOfV4OLFDj9c34f+20UEBR2NAz9oKbd5roFaLCyN6zQB+g1ppPDtIv/F5YH8Rii36Sk
A1W0q7YIn3Nj1OwSqUQqF81gEQR6Rp5OZSzU545A9bC1ZF1demLRC2cZxriP1maoJov8zQGG1/DN
+DYDpcmN3hDabg4ejXHIk1SvI3L3TdrUX+8wnRADX4GSs9gQregdPPNt6SYOnzxbT6wNEw2kxCyv
opqf3zKawCfUh0X8n7ftn4q7E7l+4RY72h7HCrG75U3K0xpsjg8C9QLgvXHojayrwzCsKpN6IuEG
e9B83n/KN7EOjeQayFZaMBrdtdKt1DvPk7tlJKnVm1KNxpldYiO/Z1cu2DXfWsuHIfcGXhvzhSjI
EuZbPeheEAYEFOClovJeGC4dxj5PkliMkSroMHDhZVYKCwaqwXMT7bXPkx0dMKRvSNnHRggM34Ra
3YNPEqRAYdk0F3w4nPjEGcJrWz18u4K42Cru1VxMAUrq+UHVt4KoeO9+C/g94ZGO6xr+cUZs9Ai3
uSYzn2Gf+HojeDZVLw9WC5bR5wp5JHnDwmpxoBOh/vDw1G2NxjtCBBYtWWrAcoKRUONlGq8M6Ot8
bcOIkRIVYfbk8dt2GuJVO2MfgvRx84b3S4TB0mAhGUssUc5p/MfzIa98nGyTas7UxnQcyJysC46X
9nOvdJ3K3bss3RSJa49yRaVbRZsoVsanXp7NYtgpREL7ZZBcnFuDxM1Yh15DJNCfzWTRVZ3hk/6B
jWGe/+T0u4Dd8Un9ROfE0k2Ii5vhYXRcAPn9lJoJt7TK0sFg4eLD3FO63ZLwDgoy6gUaGlvHk8+4
nd70EuLdqC31U6kJJkbsGENmlL50k1FGVD/2utnctXHqF2ByQGKF96sCo/VLobCh99HSnIwAZxxp
3OLFYEWResdKrZ7aVXgu6++vckCJqlgsRogFJRcoD3kHwMJomIRjbCmrX8IQYfJ812lmaaNsGaZz
4jmi5LrDsKUjHZlPiOqnPm3HvSAU24CVI6/79JUSU/RaCDKvZggB3mgAv0pXHZnNe/tqBEn/Evlz
jkFFTwsGpBjJl5DAVrrzBqGQvfAQhtiiQKFIPaTqW34EP39fpqkH6AVuSWcjMcDsPfm5gFCGnLru
0eu1sLpqJd1DOskn/+z4wZrPTipWVsbCF0Vi2EaUT/q9uPLfOUHHyfgZMSI6xYTTsn13C6jMgaPB
+Sepf8r47jUIgf5paIxhKsLfhQPo0ZUnvgZrOTbYOPkh1waPLELbpV8/xaI5iQwOt0lCoITdItJr
5//S8N4WoZuDFxdEK4ORsAT2ekboSux6Lo1IQDV4uyb3+t1MgqVh2jxp0JUuCwHj7Ss7AiMPbMd2
6IC3/HMTXz5eXgLSd/lfsB7vPlygfRcdq2RmQ1+/VVJk1yofdNMxxGtwL8oGx2Qc3tE8H9H3cWnh
bzRdIxBtLNFjGP7SqjJlAVNpUyYON7ioXWxNDgiDrjQiaO6a3FT4zuUS5WCKWAjnPYMXKYEItoFJ
1Y3ch1ZrOQ2T5+M0OlIvIu0B2ggXmD7gk/teeRH9Jy8clu6kDYuVc9TXouC/o09ZrASA/Nw/8Um3
px2I4JkqhvsUxBQ2aqp7Z4Rjr7qWwNmwOe8cPeh+eHDsT6zWPQzO8ioW7l3Q5xzkRUSncBvv2PJn
wXChSnbYnyZuWvcUnVKFt3ny04jB54g4Ye00tL2ePq8way2clWW5lYHXrpbYDt/UeSAg+s23Itct
YVPwRwmJnY+LnUVpUHvLMPA5nhtJIM9fwjNiD+QMsyHGcElE6RaQVtOl9j20ukbLkg9rYlVVfGmN
SzipAucD083QbXOrC7BLhBgnbbiTC258lxRhfUROfVAm7Eador+SsbsyeikLisZBQiqYKUawETK+
8by/lM5pbvqX6su/C8yQ+fQojd6Vf+qRI35Afod93/Gad+uy36PP/XQB2dLUlr6YPfsS061CXrFj
KP7bBQnBebVq6QFEgejbmNMHYnQQF6Ys0bcbqyjWmXnGO7TUhtR4Klo7abt/VsVQoaFvqZErp1vK
P4PTDaOcgkvjiHpVl4JPXf9AyrDeKUqO/rMZJUzA6mGM6n9JBbAmVH5MYDTExREKjBwZfc312A3J
TTIY0xLFk1N2qMEpfVMElNQU9SZToZhrA970tU3lkSm9yxhFqn0QiE6xLYFPGgv2FUYDkLjDAzUu
IQuDAS1sCTLe35Je9cXuo+qWETCuXUwBSa3rRJ1dirxYfPLEFG2nmqfHjhvPLp1GcV2nMrTM0adx
rVws6y7VdxE4OnznOiJ+p5GsKYgZzn+3x9TAlKzLHuy6suUZrq0wZbwo3SB7Zu/XrM0PwI4962fA
9Sghmsj3GOEYMp38x/heB8lSHfvFqQBIOl1QDeezD8j6krjN78TG4VD4ECmTJKtNigewDMyeqW4k
53Qd05KRsym+HM0FhPZkBUqT9i9nOsUCANTTmPj2jM2zUgz0qWeonvx6zZSx6VNUX7drWeyK+EdC
lXOhm4c67xUkCd1QOMGg5Y3ADdtZoBVeWQfGs5ggV2A1AoXqkAwEHq+MwSIaJTj0Z+MpCxriN24n
3RAuBtqWgtTEhRu9rtyULYB+YytYqWZi9yNhuhAnErEXks/BUp/cvC9Q6sH4OQmIhmaLMegXeu7A
UbNZlq/SerArk9YHNDR26YffvZrDvcnA4DuJSZU9jOuA37VJW5sSlxmwPLIUMXbGuhynf3jXMGVd
tXHBgzKWPk+N7Hlwn8bDj8OxMD6FpFdtvjHn95O32lEzs4vs4XsE+DRZZaY2iwwPzSM2AE41hIi2
l1ZgLKK4b+hOKxCTLDUtrTmLCZgctcnpHTOuMHygjIqiShchPGWTAQLdS3umJRgTRbney/ZYmK1k
R1eW1Gq+e8SNc1DjuPfWTwX+jmEbbCPk8BBg29cTLhDOBdCkSokHGABhbKThLREkPM+qUT0b9BhN
1mFIplzgNAeEvPS0qeNZWc1DElazPzPnx4CbM3IyKsEzOMKLFDSHLofcgSVNv9+gymSWrIYpxppD
anQsOXbtml5R7sf9XSB1fzaShesmpSME6YB6xCnk4k1fnGJuN4EE0B8MuW8tqCtQ08kpMxXdr4cu
sJqYgDkuR7iNRRjAEL1zXdnKZKq1daszFSIwJdtUDrX83y3XUpvhAS3VVSkHDYMdD7oEWEXPSRJw
cni+b8tQTI81M68Aj33S3GUbeGa247YguXevfnaFq5PRgOBN/0oNFmWP2AGt0ar5qvfXKk0x6z0O
CF2t9/y7VWhUlyJO+K1bTTT6DewuazKSyUe277ZBOrj/eKAMHnpcs86IDKxGZvxg6ew2OYcHyWIg
wnbouOMesY4eQPR35FyL1bpTWLbbQRlc/w6fAN5scg2BaGE9vquSah5PirACt5FVQgWf4dLcMarP
Ypn38+x3gSabwfXgTj7uSloFwRSqWswQikfXEEBEFUT9vgMaekq2rOlYZXSD1gmGraUEglhHKkVz
i3mkOXIdq2R1CofOb3GWvH3HWeiFpicDYCD4EDNC/n+1PI9yJpUlxTmVOQnZYwoGmhKozNCp8Z+7
/PToEKKhwXItt3rj4ybQOwLqMkAzOaw2VTUAtsxdtvrZtcRoR3CKCDG+eXJTpo9f3m0G7opqbJE0
RxYF/2NVdzlIMu9SKcPTVSlGR9s95PeGyiG0ix8YHoeoUCc+NNqqBM0SfDgmegXJg4nCp/nLcM2h
BJxxcLiqiVd1iW96GPrKo588d9/xF6iHbjNWfSoV8FW9ApkeE97ofJjylytf1zKsFYBeLFO6zEQZ
1fFQKKGRw5R32wsgQEscQTOYnGkXIO1gBebFERkg9nHm5/fncQju3K/HNqhq2RJKdw3ddvVmtHPW
zmosjk/DWVBi/bB+hvv95VH8UAkrr7MAEuKMNuITazO3SylLO2A6xSOQ+SDVsTnb1lmTwvmqvVcK
JZ4MoBA+4aHCqCS8vBTY7negKkwGbODSbo7WHqI9+KjQAUw/kMUSX6ic1akZgmuR77z2Mz0DyLOx
4K+GyHPJp9RzWK2b89e6XMU7DuKMJTw1RV1UN9rEbHafQ3cyP7t+DeZ5C1gjm0kxavLT/ncUOUTD
jbBym26Q9+R4RIM20QHKSt3zIFoPC6IJ7/uXxwhImYnWCwLXU7I+ka31MalkZRcsa2NP+EGP4nIP
3zgRgf4dqXs1Of1CPI1bPqaps4UZYkQt6Uhxr78KWQ5gs/vYOcvb0f7r1W0l7NzJKWs6QFHiq5tk
zNPQFUJGYmhTmC3LoCoI0UFstpJe+XVUpU+btzfw1EVwIeCJyqE3W+5ULuMhcQ1X5z/3ObJ/fjlk
MroPOtM5kFgHuwo5gya0trmcLZYUrlwzZVqiU7Nw5ZvWWSksZtvTFvcEKDuEYYuqWXo7SImn644/
4Re+fbvjUJrfUkssa/m2qMeYnrjCVg5JTGw+O7rYyS8rCDZK3W4gFM/pNC8TvWlx+XdVn2MXKtKK
HxCyAJSPU1fEFJRQ0pQkIRa5Zh+wlIz0NHahBqINhaJEys8tHtgXL4JIlG4zHxsGuib647+a/N2x
j9Hr6g5HOEgoguBu3nPYxUDPt0bZDr4qfkA3OHJg1N863weN+WpzOSaKteMuu9BdZS+4+rWkQLsH
mX/awSi/O68VzKjUCPV9hk8l8Gw7HeoJs2JtE19fFI5SmS1wJ+QU3i3RAyiB0lJm/N9aAz0kEmY4
5HRw/2CeJc0FWJjfNenhWewrrYxS/Qr0CchUGcI799g7cDb3Ze4w/bdQlNNyoR9/IrPNlaRboGJM
0ybJWm/zh2dCeVsCFOUwKqagMJ7NCW6+6JZqHfYVq2MHi01Q58VdpCnlG6q9tyqYwZbrXG2F+1+K
Gj/BIHm35jlhyEQ66b/Lb5NoMtsZR+31fGS/JFXxJl+dbv/wMZt8WBD6aIHfxCqynLYOlhs5j2Jy
P81phlpa4LhkYQ7a4e1Q3StM+bBMzE14ozEOXaUYF/zh5jnToadSXu1+Zp86Koh7EOA87Df9ZuYZ
LdcxXwVc0AOCjIs2vnbTOKsfYyFt+x0c+ANI/vmLGcvDJXhy4wjbrZnzxJBH64xSMpYFlIYzhDFT
GLcpvtD60yT3SR2LJ2TS9+T3AtTlLLNKIi299natGEau0dJ8mx4yXrqDyEidqauxxlsNnNvX0rSj
p3DXepVj8+8OfyvjVX+x159tMwhD/EnPksRpKll4EVCFfbKcS7pdAiHKP/ANgqbi+XUEeQFmaNo/
Ke3fE6rc3lmwHj/qJ+AI+2H4Z5IDoQzhAZ0MNqmEqyjGmjGLgCsmdiKdjRHY9jdrnYBlaFRPJiNv
JBTesIXJ+DmSWQeNtXFVwA+y7kASMLqtdPhIt68lTiLj6W6wInEs4fctyiXictEpLNxiVdTyzFvg
eFDQYw2QxJ/2HWwvRAZ6K3U6LmHMNn3oKw2fAF9FV6e7lyME7fl24SArF31+18Qbh3Rg3lwenEIy
LTK6WUtxSkde8Tm/P0UxX6Xi1TdOJ2OuHx8UzMMMpmaYJ05EwNCwBK67ortfcIvA9aZUZovc2cvx
71UHEmMtAtGupqpnHfSk0Uz8lqNUsqdjkoNxoCYVSDIvhb79IdKVrByX+jOY9RBwMtjISsShiRcF
tRQ3xnF69YcELvbRZ0RIQmn2j0NV6M7BysR0opUGtgG/oui9eAsACmnyv+aAJHyFAJBv6LwJbF98
SO08RZnuWn6kRhpHX4ab4ox+6TJA7AlaTZmssBTP746S2Bq+6FF2DbZvEdDdIkuqaAurjoJKjmTQ
LYLU4NI8OZJrIM/b971tTLumI1hRsFcBxEPzUG67UUuwsPaVH7iEH1DBzeG9srGXxvNrcIoPavNE
SOTxtDdy/2YQWn5z0UyHyuYnZMA0BJoVqCtyLX+nzmCshTWq1VuNaErd1dkRb7jq7GFIeHF3PJ7Y
VqqdBUd8hgPdQr6fHHTLIg0ATNmoxIbQhtOPd2dDvE2bKW7QxA1jW4HHkxU2pkjLDuHQJBRefoyQ
hCykJeYm6vXR8jJ0sWrw5eMBBSVghb8n7zP/XFJQmEtRIeTKxyPglTlGUPO7OOH7qWqTN7yGqDzx
dYEYjo+4Fd6QhOTKUQEKTbt45BDqCEfjOmjqh6xoFDigGoRpYn7IQ5E1Q5XahIp6GNnZRaS3cOje
QFWM3R4QVcm4u981Jf+2NQ1xIU/fLyT4ci/cxj5Kv/NGusdJrJVASI3bbx9crRgw1xks0uDCzOW5
XN+wJW/SoOYxs5h/uLJQIJQE8lKz5vZVU9Su4UEuOD89jsgGzBuU73rH2rccSFqxtOonHuuwafIA
F6cATdN0I1CQEPprdAfbq0+BIb/pcye1s7TVHc62mNss+QrcVCHk3MTQ2DO0qDBeAFGWzykNe+A7
9+9y4DJ8VoXzkC4kmCm40/2CiHfx/TcPIKuln6eoc/XwEuWpEIgpORSuYrvJ2MSxrQnW0RNa5bA1
yT9/czYIrtaJdsvfNwzH1Gn0yFQ/0o02eM2kmR9ihdWvpPMNXQuRGuFuLSKZ5NrAAM4Axt/u2HiQ
0EWZdbskU8qCpERMJh6FGsaHlLs1018y4Ysdtqdbu0Ff9um9TuMhUKV+rkLArbp4pw6pXH7bzU4s
SYh2hjxJwMH+5q3ZdPjSjAIIkPOPIv/NnfoHGKPugs1mYBJNoIqUCuZ1rgfmRNiFavOuJmrhvSsd
Ti+zg8CCaERofie6aGwLdEBPqi/joyDka6RNyW4BS/rJuvJepp0/jiN9+Cz9O9PcUqT5wNi07bcI
rAWRndmfgTEkeXk2CYJ03pRGtk72Wy+cSB9aqKwHXxtE767T6dctwtvlU+8Y0GyLovsqRbAscwnZ
MDjxOS9rhT+YtpfK6yaozRNHQ+Nhf6eDnOpTaFQVzYUQEzd3g0jrpgSQ/ke1BPMf3nrwhAbuUA79
d34sCs5g/Gm01lwXr/zJLusetujtKqGe+45Pjl44wyo0sqlU3Fr21lDmuRyVqAJ/vO1qxDFRTSne
afC4X2aSzI87iGorWw7S3D/m0Y+uYVm4uDpUsJ37nYCer/PsIlRSL5S4fwFASDdV45wEbc+vH+v4
W3ARzTf1tolBWogMWRHzK0cj5qaPg+bIhhR1nAVfZNSYVx6kGXMt8/bHOHroa0/kgqbXCDqsuCpN
mJD6GjVD49qt1Jf9hoAmy6mGLJIFt6NB0knkPyCqiTlcndSVH5NTvnbJBwk4B3Q9V1yZz2i3SPbY
7vjHJLOi+1Urr84yht+tSTHKHkGq3O9AF2Ofw6QnRb1q6QdBpZ0TzmgO/o86bqzmrbzT8D24F+BF
a7bs2MY/bwH0j75HvNdnQMNDq3WTXvNijyC1JIQbNIPqW3fOnxsEIXPmjSrsY5Sco3bsjQB4KML5
vFyuHlZKGeaZRPHZqXehE/WEpqT+Xg6xA4yM0hO/KRaFho8aj6HyzMvz4krWwjG/rVLHahzBUTyt
RZT5Z53HOtSt1Y248NuKXVZ7A83GUWP0SrXaswrIlsEiibWLI7hNEjlzYgW5+Nx2gjYu4FBdVSDa
RfC64xenGTgHC3STKDuZD/BTqmY2kZq+dO3Jurj8WFbWvAKeaiO3hO37Q+9MeJjzuUzoDulKMqMw
bisx/p7168vMCdNpkNqqm2V3W/PvAhN6ASzJV9JBBVfvPIg2D+WHLmlTlNBqcPyNLbFC5xc2j4Br
IOpd1vJMj53yiqcnS+JL6gIYKfcxcADYeImOF8wCt32IW46lSiaf877/9YdBCRReShMG+oEDJwEz
aoelT7JDNtbnu5A+Dy1DYSBER3lQ+Yc3cITzBYMjzT6q0g/IRdgjZVQqnXpnL+6yYe0zKp9MD6GE
lwztZ5YFZrsKbNL4Lfp04U+7uNXXscDjZl5HW/8I3Gj1N/boLMD7v/GFEHCvyNBteNurWEN/6Wtc
M1bN9IzlxjvaGgknv9CcLzWQSkAYX+Lz88zMzrbixbojJSBx9aBbD1SAVlR9Angll+dSWVZ3armN
fweKBf58z0RCdA6GFT7t6rGTpvsJGf9pmzfIqWsU11B04x1eN4PdvEkw1zsmfgcpm6Rbli3mGpcL
SL+WHwK8MjqlYMFVJYWm0krT0C9gemGsHlHXbJmi1eMvluzebMci90avOW7mTPcZV6cd57iaCDz2
KjXbCSIa9jcnlrjIiIhufQ08KGBfRdaOM/arbeIj/jOOmroa0oP/FccssgX4Ijpc7FapAm/9ETYN
gtQni25S5a3DKERJkAat75i9+NOdFGgJ6BIwMP4LOW76pwX2U15Oj24xU4Xu4KmGR1KtxLtNpuyP
mnpzORydBxzxVUc3qFMKPlcqCFwffqYtYDr3lIMKnrzLz+E7DbotPfMePnLjPOsHrcca5pI3Mw1i
N71oEB3GKAxzd+zROy/wSlqtelmQSocCRY49hGyMUEGu5brThDKM3JI45aQRwsjI43EgLc/0a2Jy
RjIsvT61yTfHISvipay4YcmS+LqPWON4KB2UKvSWmKH1PPq1pG+kxo5JudYvq8vdmoZqX7fvH0K9
03DKWfZH0Dudp2W5iVVUsH2aOkh//1hq7lwnjNXBLqpH4F8wMIAa+Sxy7DyRcN7h/bhcIFs/YKDc
raqctr4TgDZY4nYzKqRt+c6paphbFROFtIqpZ+xZri20GwXWj92ZQwHD/qmWswx+MVpLbUauw0/1
YOupOjwNlP+hU1h/0DWbjvl2KImzTjyGFYh1rKqWjjnHEqduEIOeUQVAW+ORvaca6JXnIbdoJVwG
R9vmT3js00DwfKqyIjr0BF3wjbb4NHLUJQmzxA7tGdeYFu10AkM61yW/Laa+7BkkWQV+oVHcE5dT
JwR4B7rlB/kXpUTxTotD7FnIPi1Jee5J4JMklATPRiemXFLufP/IQcWMgS9uCPqRENTSGUY9kisW
hRdVZIXtoWLZY7pKHeTDdXaR1Cjem2T9QZDzTLP6iMMLtoVOJtKLWW6/bUfEnUcorxzVJ2UNS4Ub
O8eULPt46KWpU50dbruL0xyIudci0itY2HMhty1Zqc6CWgEAEss/TbZxScw+ws27lVk58leWBL43
5dEss1BDIBfKwif9Kf+YJp11fsEHtAF3ANbpBgn1ouaoY5y5rh8kM2Ozjp/06Rh/pR/LOEMAAu49
3Nl3XiTAiDORyYbYMRR1I+vivBGUi8/zvPYdi3Mxn1ipd0ZeWLgeCeoGFj9svup7nV6K9hFZ4dTG
lAKCCqrTvXV0Ljy5IB+92EAmv6XMMdEw7WRjvFr6ReBvqsODd/jsDfqKQGj4MRh61FrF/fRQol+k
XrilB1NgLkh8Vk3LdgZ4wQSvEZVx3WRKwbUJN43u3fa6vqPWpRIC00jg0YzpiBYsvF0TFW3Y4mAB
rqmAMYziie8S6S4zkRFQuhUPGmqDuXlgR9r7OtE3g9Z8He4wmtwjNgjlITcWzX2TqvolaFSs5vAp
ubfSN365LVK4fY/xYyEUD715jMqPQ+7yqh+RgQ3/wZtnrD9EUMOfvvyhniUnpYvf7bI+zFO0ghb5
iPLQjIjh4oXXvuUKaxQqY58TsuwwPi4WoDVpuIsbbA+wDFhgyOZymAWo3/MB1gNDB8aSK6Rii++V
0iLsW9QrBwmKaMarLrGQe5dmUhDQFRi6e5kOHZPnjqfOG3BzQKmNS0yGR3NLfOkhe7S6lWS5TclW
cAyCGKUfDLDuOih5c1MzbCr5Is5XHOcqJoRV+c2+tM6RcY+ZRKUF5HQyOMmHl8yvPJSTkEzztDCE
FS1iYstW6HvbEJ0pJ9+LnxaF0BvI4oTsLe+LxJ1EWv72TFQ4KF4GvOE4X62kcyFa4DZaXj08oZN3
c1nE5Y1KiIbUq3Smthq0sSmZ0UkJgCy+z8eRlp0g6gIOurCa4iQzwaRDGdR1Q8eXi3TY1GrG8xDr
UbgbJB2YsLG0fYu2kVsuhyOnzhMygFNSnqXlbDPzD4dyLqKeb1EDTPNpH+mJaEaUJBqSm9ThXNx4
Sp7OqhjmD0BsR8JmpQt2wb648uxTTnGCUsZALfjqtqhp0dC5aEhBle7xejEuhG4a6Gy30t/fw82I
L8JVgHCYvA1RfqG6wr3s11GjXKKPhcWInWCwh+ISowsQ4+AlQJJu7v/gSwIDPFI4cDgL2MgjxigI
28KGdqQZp0dCKk9R1eejqJ2S27VD8pbLVfIfusUSrcwJEVB/rX5i2Ws/RYn9hX14e/N5M/idrYEs
0YOYxcbmsXDqJWm8VMqTa1T6dAK7WASQvx48/yxojTxCU5rXfhnXgHU6BEzmgulomsA6q2D4ZLiC
rK1muCPESZxOIWABcjqIRF8RxJDt9bPYbVT6M8+yi/35K7aeIFpbravKTbA1Q+ZwXskbfFd0NTXj
J1Td7LTMUm9NigOErNbSJ11m9OLTwwxvzrIm4dcV/lGgyeHjY5mC+VGKUgyPHMWrpl6cC6mNj2mp
B7CJYVO3Fxt6aQ9SWNSbYY7NscRuFGd42wpYDHiUTbEVvZj29uGgp4ExYSkwPDWUwFxvjhzTOqvf
ASIouT2yCpMFJLwf1zfW+fnlejTkDz5P6Lvt11KHpfdeGzHZmbG3GkBeQKMLZaTbhsQVMwINhIfM
Iet5qWIW3ky++57JNFG1ucp9FmcXAFJjXT4Dx3UUjTsi41K4R+G+jPDpSIrYcC9z2YvusLapU9SW
wYOaiuGp77f4NE5HOVDhm01TKgEVSC9lU2+SrvlzTKf42INCTGcJXpuGMZHRdR/42Bvh2+vXh4AW
P+qClAEt1mSoYT8LPBXhFBD+gTjlFRSGaMqBOQEplaP/t3ur0NH6LM/ThIE1bq2aFewzWc6QGmXp
Iq035NQtXNWVJDCbbbPJ2MPz96xud7Lc88d+j5s/Q9vD3C3+HtwIHChgevvVkaop3PhewOghXs0W
niFPVC0rA/rS4NnxrVFhqqX80EITwRu1zyBeDsijJ40UZFmVIrCKeXsOzxryBs2vjx090UHAvJKv
TtNRCe0W1/T+sZKlTqsjoLQo/HK2RDVr1izBOkKWWUCOvPeU4HTlR/Ein6ORO4yQgjeGCR+1x3G3
nOb75y8yyrn0vOJucEz+apIF8xsr5RowiblJ8ssuekiQP0xlAydMPIJE5ZvVw9OgraJiCxpFAB/a
wR8Q1q5OHoQI8BH62/V6ysBdFl6twKP82TAGx7KHHXTKsHP9WSdET7rRhDcbceY5fHAMTN23hd8/
R75RJdsYiY02RA3i6DIo3PM46skqB61X3o0f37EU16D2ead5GM9L5oDgPzqU5gIr2cmt+AJqsCy8
m1Az1CKd8ugCa1goC2Pi+CKP9C0ppVfeNCK9LQ4uBz3u8lhjpgAkb7b37Rq51Y/wlYE+uM+N2Erm
7h+5j2nWhKi8LRjCapwqfPj+Ht3SN7dltTxeNrZnsEx9Dv52rvkRwxFtKDx1aht2SVohVEgSe7YR
2JOxrmAKT8JpY57fn4fw8y+0a2HV1csFU+rcJJ4pS6JTZziJ4yo82Ra7TNpksuhHJMAF+fa4YU7o
w1lUi/OjKRMKsKedSzOwuUpqzIQhwNFdm4NqkKK4n+cFefCC7jDrbkDt3ysUDz3DaiKTIze3oPOu
rPqMusVeUWYPtTBCxUleqaFIcPnIVS22hURryh7/f6PMfhDGpnrmXW7CYjshRhwFLBCwZUV6Bk+L
NU0j87qX4WQYy01rU04FreR0Q3+QEcWktKpE5fM7ACte/sy/LuNHIlSHth1yah2eOqHlnVxZQYPN
1h/Sgl7URrAolqK8ZEZpoQMipbLc/exsd+cePFqLMS3Sj5FSuq8R+eQ2lxT1ptEksnE3+YUrleTC
latnw0J6UwlK+XshseGp/Gs1iZefiIQmugAUDVNocH1CDFNa+Nk8iB9zEZd1Qw4Y88qeHVEqTZo8
wx8yamFPF4TcXElVSYSQDJrtNz7S1404vmUgMQqCimgBy/LD/kBvLkiRmOwBh5slXTtbxgAgSD4e
0AxDpI1BFfxJqdQQL4hz8OXUYHuAC0JJkEHOCsMqI2i+AUgdq7ZQarPEIleT+pbie9JKs+F24uNb
1rNxL9fRFTgFuegiOX3w0/FZYPUJWXOySL32exwkrNBrbX+VzAavdGtOZZDTKDD7W/U2Fj4Gl2gr
gs+/2vY5chqe9r6ahY1BWdk+9hvJAcOB+EshZZRmml87DLeO3K9zzcjIP0Z1yADYW/u7L57/90H6
pt7R1Dp/2qGMKE50ErKqIbG1C1vxfnwpyxiQh4ELXpdpLtopzd6Rb0Wdfd6jLlY0x1irdR8TZf5K
1T6N9q0ESSD9KXEjER63jObTndTo1PI4s4cBcVABkrX2k23/8Uf0ukqtKUl7vvwjoBszSuoy/kNM
M80RRIzpcTkVfH+HN4AVvsfzWn+ozGeZKrgVqMuf6Aljfjt2g+xPJV1uEADw/vDNrz7NAmD9HTAf
HTC16OMGIaiID6Cs0g/Y7TPFnAaKhUuEnBg72frG+LRbP5Dwux3lma4Antut1sL0dGS9ZS1JtHX/
ANks9pOFcciLZ4bbM3TpCxO2RwNQur93oe4mMU8jrgWlJe4Cqih7BtfdudcjXKzhVABWUsLFKlfZ
7JLW35UcPx9HsbZd2iZkxR/gjtaB5CLNaBcGPmxDTqhAYaFx9J9agb47J2eaWkXbr9XJHWCXup9t
A/TVb+V5V9Het6FmU9Uy9Zo/quzuz4xPcveVdahn7nVAZ2SYx5Mv1AyXL5q+z7HdhAN3IteUqjc2
AsWkaxXXXKKX+dTyWnggE9wUgvfhp9JCb8oA/zum/q7unR/z6bqnApub8GkP0r11s4ZF1Gw6D8Zu
yyNaSLOvsNoGSqyFmTSiw8XBjaQRb1JJFK7QrQX6JUf3YXTHI6a8jTBwpZpN0FtPnqJXrOAECk9R
7KxrrlFEktiKs32klDPe2w3D06U+Wiyuh4XJKsajlSmdo6l/JBzVTeFIIds1UlyjfjCs8y/V00wL
Ykwj3Pucw/tsN6FV3gU+DbfGM8HtUoYlzT//ige/Mtb/GI/Ck2UPDTGyY4nH/Ksfi7E7lHnsXECM
o3HGvvBmRnNWKlrCG04I8v+AAtdddbsSUBtKdrjpsBu7WiVivu3q4Gcon93OQiCxoInsUGx/dGUP
Kez4oHxBHhiSHdQv5t0NgP+h/uF6Y8AwEdoN/sEp9CoX8D0SfAeSNMtJ/3YgAujnXEOyEPz01eZ1
KMCU7HzbEmINkbPaBc7GjDCxe1NYJ7fnhRSFLVSZApkwuZ2pAZQWejCnE76uK+TLXLqIqv3M5Am2
QiY7qsIyBntNCX0RaQ12xwn3EfiWUIPWSsDN3Hd8ppQFgWJOkm74Edtbj3gWgD/Wzxn9/zkHiOEM
mLS1QmId+XFxc5azYV4M7obhzSgRxe7F7CNPJqUxVpSkge14S9jMwStfiz/qZs5jx+TEG2dqvexj
tYqK3afzthbhXqEOZvFBXWRjNRMLgcH7ujEUgEE6lU7VJ7KeFdnYbu/sVxuBjMPincjGxVlkU+D4
bsDN72TdbEYsRp5eHFVxf9jGFKEu34ylBxSREuzRqgxs9ivs6byB0RxuA1DUPFjjYtbdIY7nAVom
zxplU54Bv/hCNZ5L0H6mjjVp12ac07Qeqax1mPKDsL1kqqQfGRcf2OYOMADluwf76O8BUiMzI4cE
n8NxbSJ+W/WKJcB1quGFdIeH166wNF7JTOkJdKmSilzScuwrbNNu3Bvk9GPIn/9cyw2JpFrB5sd3
ry9tsrVwZ0Dz8WqYdpapjAvT8o5ypHf4yw4m06iVC7akjJdBU5jlDqW2gOho1ydwtT4qRct9Ar7Y
jLxFLb6MOnkZvG+xnBTol9FBeCR/mrvwr/20irYdrtA/65JVp652SDcl74GkeYS+IS7rAsrVZeHn
4FlkY7DfSfosirxxo/MimCEad/gk/zj6kajVNYW64Mtn/FjeaHo/OhWecdo0jVQhaYKqm4l6MayB
Ha372UcMuAmm+YK1YFEapZjVlWjqADu5ngkgCKKtZSN8lgoSdSdADR/HxyQ8+1HpPeTlD6jPPR9W
qyB3nNzDNKcf0JVrbB7UA1k4fgUwjIIWcojNLekZtfvxXRbDmc1cqg7c/wR/tGp3NEQefau7aCGm
yKUyFldCs9v/kr5tUYnhL1VxKHfGUvvuPSpg/dU5fTU9Elwcs1mMkwZXGlLSbUU/Vs92YEEpqgHO
K8zGhphZ7PEkKuP2dkfuKaHfsu5Lv3NdHbP1RZjPRlnBdRWqU3C7T5LKGVmNyUxEqeWrp3GrsAl4
xa1bPI3aAb/m/vixWU33eUaknFk74red04RWq1FlgRoX1kiUT0SDy57Ip/xrwG58aN1RnWWTnB5N
K2TkU9ztC43TRrzXneEFNXf6buKO0p9GQkBoRT1QaJVWr3J88u/wt2hkkil50mO8cnGg2SvKextN
HjNDkoB7cf+lnF5ye3fglIbjqW0+7ueGUaCt9gSmAYHvl5ZOIfN0X+r5sOD1tUM1m7+QOn9V2ROg
rHHnOfyoQfJG8Cwd3qMQkJ7PqgH8QQEdr7VodrL1G+dE1wZyMHMnTXyMBeI7iVif3YGB1yhc1Pj8
wpzK5oRaMImBBd2igf5vAzBWi0416Wxzlh3mMptYcnPTQLBClM+IFQHI4kf3rjlDoMfzUe3ZDsmJ
90YNQLFbf75a2y8HIC8Y7YK1EaLk8ci6XRynX/aqBeqFDF5NDwTYNRFHspP9HkrURLQNxcfCalTe
k399zIybRkoBbD2zeHXVmu+ZH24Him/n4WLGJA4DPzjqwZ0jzNtIRULlLqdyuh8+C+H7mOCkY5GK
D6xWUNw7YjmjpRZJ4rM42xqRGObxVSvCV3/n4u+95cxb7miLt0KjNW43k/5V7tsShJ5R0IMiL9tY
pDKEbtm0F1gQHKAoj0AoCoEanIWKrrxaDUXFzaZDCQtxTumGzDudtWMzlKcrM765oqgkbzze9CuA
YspSctffCiabdDH6HpFkAlaj9gO0l6p9MIZD0bVC9gelNen8oMWZGzyr76yJl6ubB/OkcYxtVQpx
croYMstS7MMJaWnMTUwi6JZI5YZxPyM+jpEFvYlk6Cqx/t9r/f31pxXAOXVwBbWPIRl2BozD0nKp
qhq+CyRj5+pO3Ze80l0ECoNJI+Phx65dWMzUAiRr51ddpxV906eOXwbX1vFEGeyjVqS4K9n4xvyl
aAWS2PoO0tea+snmdPj1xRk+IB4j++hm2dBeRS48OoMd2DyCYtoR3TqkWZG5YIHnCC3AkgyaBwqk
I8NoNW+zTbupKDitlHjpZAWFVzJ6BZJ++lIRwOf3oobmtLg/kmwS+5cye7gsXkP6rblni9HkV9ox
oNfBkmI1zTPGCj/TMRmk0IWoebQgm10gJs18+fj0uF2wp9+UAi9qS8lY/+ay+DzrHoaDmQjm+J9o
XTgDA6Q5CCC96UfislkiIlHwnMGwdngeujy7KEpkwPoylseXfUDxJU9nuPeVzPaDXjhAhQxZTGFl
LWOr0M+LtvzBEZrPrOmPuypsS8AULmkUN2HiAeR4IvdRyXFTfKQIWAP0xqnSvPhRDCvJ4aUrBGg4
DPVcLFXxyiZzl4X/Ut5QNMNKGTb5cSzaB4gh9M5oQeMtANQQd/hGnCE1cwwpziOtnDHQt5OHfnO6
MMMvEw6gWdC+lqDy9Mv2ivIIesnPJl/w0BsPMLItO7BcSFzhcswPLC13kgVTgh1kQTa4UhhB+kOf
vAXigJ+cw3jt0RSkmWn5UIhBukoAUAN46VpOt6oIsCGJKS/fBp0hutFwMe0wRH9K49A/vw9Q52Ow
2G9lt5WTuHFk1n7sMFtzQRKUPeLE/rzCQLmdPyt46FLbWBg6P26sk7/CpY95pk04hT+VFPce+ZnZ
3GQVNr6QbXXU4+kZIu0RYw0hX2ICm9jGs/r+qcNRJ9hUl28F4hTDYPJ7/T5aL2Y4MVuCp3oxxHLY
kKETc4ER/eE0epM7Q38jz95VIssrS4ein+E2c6Z5l+c0HZo4qj+nPsXcZgxVCFiSCKkBstU3JTie
HMV4d3BPYinJ1aPVLXo6OAsttxb1DDMlAgmHbTVZ2aUN2Hh4yH/3AtndzBSMKZIEI3LqDLpGhIMv
er1712QCaVjLD37SgARlUOtJZ9LMRWjd3zxmVzbfP+S4/EwbArL1w4B5CEQ5PHUYxADGF8LFYQc2
ntZqSCH1j1VpeBsk4wbLka3uHiZGKhZXmjLo1YNCZJPlC5JHAJ/LC9Y3UyCzz+YJsvaqkXVmiC4S
M6JQD2H8Xr9mkKjD8VONx6TE9oz1YHDpDd45S3kqNb4QE5ThqE8yibPn5Bwd4GzIVipAKGU5oQxt
OHPg1I7/hIBwUh9dzIsT2VvwOUEPErU2gTzgB21CuhqFvpBm7cN+qvUARRF3nGpn1b1p0b2DapAE
bIkyv35DRGA5+7q97Q+wRViSHNJscZP4morvN7mXd8YqYOE8EAxBN2wgrKxop+cTAthkUAVaPPMX
WZ20esDibZ/EO0WdQupO/FqMaj33eugOgaF2QtvjigYg/wM3FuQ1R2XIcxxNPe/BUsTaomz4cH+l
8Jy9n+tdY6oMbKwYXQd1jmy+Obo/6moHenwro6lJO1tmnloBa2JsEUirK2OnYgAN2OTZSIfoypPf
E4cFSOc/i6MjsqpSz+uv2K5po28pHLC11EZDS/1+nD3IU1f8LFK3oqDxxMaH50scP+ltHcX8uUE2
jUivxIRYGYRpU0RPVu1eBR94IypT4VnOzOjBoU7bsnYrnlkeNurG9/guhx6xX7hjZrZqT+PzijtM
e6sBhtMXlnXuLEa5Z1FxlGBBY/RBNmBJtQFjGszo8vcaYbCOeXj5NjVgAyWtGLtCbpR5iBklJ/kD
C5/HJyTptnq3iulC/TsmQ9Im/Wvf5SCHNTnYh+JEo91VR9ZSoLf4eA1K+GhFwRNJrM1iSNfpXyet
uUYr4Ex7ZX8rifZSA00VgqahKlqijV/Oml0zYK4mN3dTq2CU9zWFTcjLDoj/FN5ntEDJpYkudYEj
QZ7oDZ1BFQp+hNYlpKw4MWM+ju40kYEFzzIo/r020GsOw1+yXpZQBky1j+JqRuSMSaPBsnkDLcm1
RwJLnUcEI1eMY2DuOohRKivH6zQ/T/tAd8b3qZWCj2lYn6aY8nvP2iyOcltc+rwtxiySgJmfryYF
O9/3Bwk1BbTdV/iVkRcWTf+dt8kAFeoUFfKSAwlLS8vg9dRuXwTyt9cFn4DLnDazkT2aeksPpE0c
88w1a6iod6pXt/KTUY6LIRKmt7ZQ4v34Hu1WFqTAhsSriRuW50F7y3si8nGhXdiliDQPuwP9897t
t+nRA46iulDCq8tpSTOOCM+VQN6Tr8ZuTTRxLF9y1aEOGh2/abIgLrM7ZAQjZ4bcvlYZS2Fnqhcy
2X/0yb2BtMv3WwarX3ceHuZq5hylpCqftr4c+z8sGrJ55d0Ke4WZloUIpRPJfJClOGyGFm9nZF0d
Q8uiod8cLw5dLoYEVHxRYK5KcXukwti7OMn8ZVDU+SNEIxUoBbb/Wz05Yh8uQ0eMhCnuoQA3uOrR
jSYYdc4xS/TjP1Ut2I7SSa7YbFWpzHIa8wU5ltqpYhYUi0YYtzy2sxJmIPjHPqUvTpVU/L9oiVRt
43+cj2IkWgAGjvA62Uu/ELwofdhOmtOgfmWqXERBMuoLE96HVmlRMyj7UrQSWAqkp00S8vs17VwC
b7tYtV4np8Y6/94nygeanvL7qtYejO7JNQ65L291WSZBSxH5eu0Vt3iuuKJxBq7Ecf7r7aO1MIul
PSGL73tWtmQ4Z1kmzPAUhD67SDRXZI8MPEVvkMQOvdSnYcZtzL7C+4IvqTQBjrkOasv47Ruoz8J6
cFCy2w7b5bvXqy0xA0NkxlAhTAgPtmbwUdkpTUNV6dB9czOyLMBB8/No9CsY5Ug9G3Ogc8tS3iQS
LDyHWWF5XdBGdV0Z/JuZZgS5PjCOcCx55YV6halQKWmWNXuRi3V9E14Syp9cfCL7WIHdmZ91r1dr
/j7Ebnbv4PXBoZOhsnh8tDcwMKAFrOfoeEP9rb66zVjxtCIluJGll0xjd7yawQ3WCnicSGxWTlJ8
Gc2iT/mrIYwpImoW3XcqSfEP2Ln/IxXhyvu1Plw1n9oP/WocmjyzQCo00Kb9+zd9abUGG54qMyLr
wIP/zfS57rVqX1JKHX1bzS1kkI1oHPUJxan1eMtOpaed88pBQEsT/zBUzKJuL+D3sS3V7zuNkg0y
QzUzqqLAqGzc9pK/3fjUSJuKd9BkKoKKOXDosTZinS+gRvbhizRY991AtLWmadj7oZpK2fAgn9md
IhXbugsEEEsWShZvVUicoI1EsMm0GFlEq4duwjiTPfnoLqAInTDvyb5AxotmTYxiBAVSAvlgIkfC
+uvaEfvJyuIeoVVXl3kI48R/JaOlDXS69jmRDq8Iq329V9Y7H/kRVLVPxJpcw0jkQekiI9u2PMin
Kgf7rHuYTyI82g07VMkY0ueaLwgQZ+9SFerKaUxNtiZceLxfxbGj9D83LZYyn2co+piQFQAkVVI+
qaTYf8UxXPqnO7Pn0wB3R6FCT9FnotQ+ROQ1aToC39+URCm6kOjm/O4XgcqQ7FT1wpWX6/QhqO83
1NH8f2NonNnyppv9UFOhFbVLqMuCnjiRUGJw37Y0ut2CWuawHU7XibaskuOzQXEoaBQ2fcSJpFyf
BSeMQimbAEaKrClUwTo0KamQdXCVv0t9MYY6HkWWcX5SfKjrGpU0jiQS1PFrU8mJ4DD14566NzqP
Ci8xlBfGimW5ny0ELyvEL3kWE8/SVGpSRM193R5wcWCi4XoB5kDOj11d6rzHBzj2Ol774aDy9CN7
v1QsmagbSM/DRBdwpsSRzhirfpR489zNH9RYjjVCtOO9J9Am8vd0fNxS/bwyIx/Jgpjc5f3SLEOx
RLyQE+sgujpm2ctYzPBed7dBG678sI74/AoKJMbq/hxirerBYdtpHe8wU71A8aojJmmlrinex6++
xGuXKHu8zKcU99OFaCU5Eqt+1OE2VHGQ9LW0YVVR/LdIdVTIJvKZtNPgbAORDMPvXcj94lNfpl8j
yUQFX0KR9nx8HqIKyW1/s/aqLCfWfa/FsA/m15TX5asHSlr5PnybUwCj7goNSBAzUroNVPk/Y6fI
jwldF0SYt5U0pNtUeqHq68z6cOe2I9lHg4tRMpRgh+YHDDuhW3aOCxF9K3N64jldHiSZ7LnyiDks
ldZUlQqN6bLG5ql39lL1b6SYKO3VU+h8FfaV7qnrEdnxEmE4rVJroT3Xbx9gZZ8/WGybb8r1Y3aU
3q9BqwQxpaeWMHMFQ3izuS4N7trAdrhBJ3dMEQyQgDuuLk95MErLW3m419o7xIfW823rayNmVPuE
TvDqRxJZ4bQJ8VTwsmwrfcClMT3IrJal++uG6+8OeqfP8J+pmsD9T87MrQQje5QusEFc7vhfFkxR
mzz4slSSqWwGz7IkBzaqJUdDgcP2E/V51YQm+loPEzq4rbaZrQdY6442byW1hML+AOinXTadho6d
LC74A4C0+XjOjsisNH+Ld1c4ijTQuBcr3GVzAHYdON5raDOD5QNXp/IEqHu62YZtLvkifIm21IBH
5Ph1mu9TN0aKdrBOHRUcRqL5CK1n7/KMelH0AzgTxyT1yDlurpbmXVksjxV8PfFqpZ0Dvscm4sEj
q67OWquzlPdHXbo3j0cNFhlCi2Wpf0ao3F6afD++xVqVtZR6T0ABCChcn5wdArdWC3gb3rNUHDA4
mtedTThpVgk8J95WH0TODhN+ZbhHFV4Yt1zuQoUnXksigWr5Q1Wi8zWT8H1DtV/eC4LxdRKsTf9l
VndJEvx/dRmsSHiEwk26TW4RnmuzMgTUAxa/1vsNHhNN6pmglYMMsQlMo+PuCxSNkBsO05qVA5HM
6Bhk4Rbs1bcqP46xNdbOhaqFq2oXGYDG2vMaV6irLPN+VsgUAgjed6QIM7rKSP/vcW9KEvVfCugH
J12EmAJgFEcl7T8wZQMW7euo06Fn5CaytEq1smFoKwuNx4qrSd6voI2k4optZPFn9C27ZZo7OxUf
RO+OkkJVGjYsU14rjNYbykBn1R67uanhLbCtV+jmYJMaNKFIMk+WAhMYQCEJO/1LGfqB+QUXdG42
524I4teLv3L5ycuXDuKdbi09oUg14HwuwNMblrA7K7IwTE3VtabJfvGfPonPzZaMJzKlY+RgN0mO
MuFWBiTj5MxiBJFQLqmyZmR3KouqSsLnTrC4TEYOPtklDSZskDNlpWrse2Ud1SRKVRJ5+UPyBzkK
HVi3CMw1JqG4Z+r5Q037Rcm+OwI1WYLyjmbVCwd1X6ASJ95I1mxfdlqhoTMZfFusnlBXz1VSHsoA
dE5kbpNk620opxrlEcnKsz/UC7H0bOma5A6vRYkJn6CSgCypccL6+SIKrQg8tyFJ34QGKzoTeFTv
VqPE9dDZL9oK1qzR6l6gXAKEwWj0+cgfUNhgqTk8QcC5MJrwL8AS1OSCoEs9kE/k/9GTGmHoiDZE
Brnfh4KfQCEPG6XzjreXhlLrIaVdsKZU3kBokwxBcETlzeMAvhvDmk+zGz29Eg8JLJ8KPom0eFmV
rHqIkme8Hl+j/dGcq2wGJrfVxUtm+zcgyjkTs8cRyHuTlAWZUBwwCK7eNcYsevX/8Nta8YcgW5jA
JIMmSYy686XrrnJLupyQCTr8vcwy8tt2v9HpTn2kVODFjhMyo3oL2Ra2gcGVXHiWHRsLQyHYYFPl
j40VkN2/aofyZqo7GAdlTSVKxRkuyzfgdakZet88qaU5DqmiU8dzeRca0EL5+geMaeCPM3nAcHn0
+IKOY7mQjFgv8h1ELrsjEM/XC0HndqyBj/8k/zlq6bhvDZhVdB7DRDPrBo0c3Sb1AhCZV4q10iQc
Nq5A8ewtXrshEPtCiqg6cONPh0fzkZe+6Q6r/FEQObQ5q1NflUIvLC99aZnI5ye8f7btSBO3dv1F
vPNZQ5CYi9rcfQ3bxjbcBbnrgTVeEysTI40jjxIHONaBKwUT6Xzcb8c5niD+97B6atfipHqvKhWS
Vgi6KdGp67RAsxIGhjulpBbXOamsxay6aaT3narmEqqn/DHpnEAviiW9dCaqxk+BOgIPb085+UGV
/1PGMLibnKhBE1+4UwV9uMT/DfvENkD5izScOxhFoed7MVS7nkwiRu4J8p/yRC4N42iYkoCuhsnL
EXA76MfFBeTgJtehMhcRkrozGjle5jtubkZWYgeqSNR9gIET3J3buZ+Pi19MRc4lwMaSCoLlN7OJ
hjneRiuEfEW/h5qR2PHcUGWSKi0Tm5nfq0C2gCYbaQNeDYi8yFFIuBKHuP7afCC7CbbLzx5F/pyl
Ve6OyFt6qaZtzKJCq9dXNWLeQ0o5lQz1ynHteSwvjDBEGBYkuF0BKslNajOBqfDqK87SfM3h2p3q
zBegIBBSrldW2FIJ5Va2nZWkzT4HeC3h6ZSM/HI5uRUjaQheDh7u0GDdk+ZLLDUuTzDPK9IiqBBj
VUKt88nr6G41algSF+gQAyMV8a8odKyKtgyxCwZMTSgBksirOFaOGsYu+v2Z6E4ROuzPAF0p+Exr
vdr67SENlrW4DRwVk8qE9mAY15xPW76UZ5zyV+kx5Lt3xkmYzQGgf12zVBoTfWL2OcR95m6PzdeQ
LuNdBRofVeYpDPfeqy5WgvRPEw+L4zVTvgJ2YchCBOVsirwpjAlZ10jfCaC7C3PkPeOGZxzId0I5
Qes41f3OJ34aZRXYdOyMVo0cv8f2sUcg9CjJSDcUbaQVKlwf0nqTpMpSFXvq+Ky7dipFdlpySWiw
gUuJ71nGwGMeIU07ReKVz6+u/LY/3zXPWjN3BT+rjskzQG54Q7KmUTsno2ZVqBSdXrhu1L+4FDFV
SNeKtQ+RhkUYwCN10rZeGCWZqhVblFiZxrFTEILeGmuXlH8kiOQ3lVjaOrX0jUbJ4pslKX1lR3Mv
0egR99DAKdPDTUxeOU7gGLHGuhtvEmqKrW3xa493MAk5jN6WHV8l7rrXPzrzMj7lP+KjVtstPTe0
CXxkvg6cvfs60lM4HDTYCmI2Dod1YdK9Ov7r5V7/fpjppBFwVRAcdTJ3uV/9bjX1RZMRg8TxHWfR
8V6zctAMrb+45C7flqjt2zySpnW0X9JIeA+Srs0OTUg4v3nviYgomJXlgPL75f+lPD2cDy4DHQzh
6G1SWNneohcRRo88TOJPcrAG048trSOJnTtFysYkFTO/wtYQFo0WUZdXMD435hmxcdKi8l/SYppZ
apdrG54gRR2YiexAN/UbA81TCxhe5G4H1Cw5xFqV6zUc8GGDKCj1/lC51if/9v+sxsg1eJuOXlYb
WBg5gplQpNHa/YXKAjMsj5LzkoLRZbyh/lmnc/rx6MwB4XJFiA/0rGGqzYBdsEXWFyvqlppVVFTG
9jthXipxYAE8s70iGPrXCy/ubpbaWL/FGcCQ5x4+opzlLqGrG3ZRHoWHpqWalIanWGCNRYVR2iNL
h3Bt+1Fwx/nqOwZ5vyPYOLPaPm2OS6N3T3qbmAzoqMWradUC1eh4+kC/YMbc1PQPth8uQmOI7CdW
RjFUN4dkzqPy5IFAxoy8XK2mk2IkBknFTs4zy9DaGgBs+WFnuMDb64NgLzDlSLJl1Om3YVtSGygw
AiBOmZCnwA8cYHT7hgU/OUhA6hUFRm9pw4n94HbqPz/6JRaScb/brcX2IOUPwLCLHSMKb4O+j5A9
O9bkMX69uobsFjZbO2cuNu9O0LBJM5FlLNHwNAJuQfs2Ay3H7af1G4f52C2jeM/jchp/TImGnMRt
UZAVPe5HBNeklpHRWBeHcuieMOeehphbUODq4W/payl89E2b/HUxacGYYPXMlvahHjo2xXsda6SJ
kU8MOXdN2XzwiSsJhea7JsVshsJUJ+hnVwccYuehLGjLrk8sTyr4eildGMjFXdZyDuG0U+1Omp4O
aBAlRErFN8AwIiQAZHFKDhPFdLUXBiyiy+oKEa6dnSS+BR1uPw0up9ANLkGPymsT83ZPQ3AdswXo
8ml9+sKoMZhqAKlh1KUpEMs48/dSxYV/HBFT51Wbr6HbWpgB43NBFfrZl0eGxWlHI9XpGXlU2sT8
17IZ/2k1cyiB/fHNMT/vt//PCzzSD0KwpsW2Smsl0Fe3aTvOle0L32OKOtvSiRt7viS7iVcKg5eZ
ZpWkXIrJsXMd1kbfjyjCYcawBYkFZmCmT+c3EgbivUOWOdwOEVK4MZEyjjDGNOKSdJdM3/JYZics
BD11gHPKC7JkMeXiSAIUDC7f1yu7VTab76eXFu+sI2JCbO/UHh3w6jVpsp2ydAzODTdJI01yfupE
tGkewiDvRGtMPy0lI7yEsnMQ4nlOEGW9yX/65v/GZomC7xzrFk5nHRG7QODzo+oZOl8M66jF/dVe
dXa5WRrQt24FDu1vSZkCMGqglSoSeALWzMRNYE+PUydKta5MfGvPGxIJ6ytrvonEgHH/MsRudI7p
fCPRs+/5A+TsPHBaWWySThSOyZpxafnk7k5oRO7GO4c/b2khulqQW121NEeaQtuOdzDEPNd9YoBp
xC1CTaBNJ4mseIRJbh0hPO4p9wYrir6X1OZgqvmicOZd8CFJ2AQNRU8FW8fCgI3lTaJVg1t3zfy+
G6WaOs7JtnQBa5Rw/Pq8aMo6eVf1qU4X98UinIDl+eLF5YkyBC0tUxS+a3sn5FdG+FbLGqhj3yE3
Zc2RNRKix2XFusx5fL/3puwBgadLTV8KthM80mTZeUgmnEp+e1IjmrbkOXmkF1DtonugQdYKdYxP
HjnqPv9DzUT9kRvMiwlNR6cmP7UC8LOpyVn0LFpQpe4mc1RfN+IcJJYqc5MbuEDs1f5Sfww3Pyxc
2R7gtXb8CYWFYPLWpMMYD1tsW3ZqnKKspDLYMt+5AWXGWKnfkuy9sJ7s/1XojyiIZNZDS1rR9iJO
G6J7peccH4olhwhzM1padg3WJqbhh+V3vKARfynh9Z6/GYwTQPcZQvBXq9Jba0Yh48F/x3HC4PPN
lW8FkA0z3+ZIW8eGUQkTgyv2uQPlmIJif3hCSAbm1olQ5lLVQWopI/iqJNUZW3FgKr8GABpW28Zk
a8lBWXrdUy21YoYfpELGZySbxchCPHG5Ogn2QEe4wftptFm/ZstD75PZbdCkQccJF0N2Vwd5elWv
izyNlSQNOyPuYwpqgNDTeqYBl8ewfBcS6mLkw1er6d6JCmQ9mkXISY9sIcUGh7inqVo9A3WqONFq
leigq854CaPgYe8zFhDfZMJdoEOvIaB8FIuFeXZ3+rxjbCOYLrAIJvFboplDFAM+1YFRkjmHuHck
UjMMMuRmCJA1hA75IsUxL2qd6K46H9K6flWf19YFVYuCgA8tNMtqEXE9ToNyyLXjnwuYdWXbqyaf
82yn1YS7uyPWq7GHmqGiZfC9dD0cEn6IcaGjET3k5WLFHiCnbbR9ImSvPjS3FYOBjNPzo08sWo1s
LGBwLf+OvinYNEp5/EZQz6uA2+wUWIEKbhFhRhU3vIuCsjCNRLD2Nc8iW5eiKlp/jJziMGbmNvLP
RzLE2doeQuHV2ST35bqJOcwMXHHrtnEnMJM8jbtsTQioSj4Rj1JoWGg3iO+XW9MdZpk+MMHK2I77
WoY4lgzBddWuKw9cLLKLq5T52IhOsW1kS7/gcP42iW5N3LxOJ7aLom3K5KKT3QFOFAJvCUiWo8GD
aP3EKxS5Uahd9TJhfSpG/SQG8Te21qYjN7PKmj0f//xFS85UGWhi3aCXCNb9GfzsRJDNfHb4aTRe
T9CtPN4/oGJARo9H4WCWtKCMlXIzGgGFjvFakALOkhJeV5zta9wZOmAbYVdem4V5RtOF58bF4PuB
WiCKKb/4h1ekyqfq+5FW//34uHqEXF5s0WExxaTBIVeQZuDWQ0AhI5JTZnwelOudAO9B5UD1WYKa
hD7XcHC2xtxZoZRt7yfgo5EqV6sj+4XJMODCcb1xOCFaFo4PsXC/P2sWbImuN/K4AG5vKVraiFIt
bC3RUgfKEF3Y1geAmKqf8FLZ0Azm25PUA6KOaFG+wCmHD0GEv9FAR9mqnLsJ1wBuQIDTZIeYapsm
MPGOxCzfvEmw0BDn2/atcOwKaR6kSPmRK8Eq1huK39s4KxagMIYHSG6paOcqcy46+ZwvEQ/pj0Ne
gWgvS5rJgi3JRHS/4qxOgrLiRrWYl6rkeItIyDxDiConBsSUaJrsc2gWiY2EPJ27dyBzuDXWcuQA
22vfTFDup0feMiRU/0TCd2RQ/Lx8md0ljhgLt9mw6/4guWjXgIgWfx4kZJHLGy2gt38twvTjyTnL
ZbXEsKhyctE62Vw3tUo0PjMOH9mA06Ufh+t/FaOgswZ1luhWd6lAK2skD/din2r8j97SY7zDJO4i
YcbdF6ui0943emUjzAW/8Zl8ydzNmpxMJueNJ6wqaNPXYBfRY/XTdP1ztvVCl7ITHomOUJ3Z6/1b
atmNcK+5UUTGE1eCH/MxIkCSugiIMgGV0eUifrIoZ4ADDD3hHCzsHkuCv4+v5pSx8dQdmdnRwRTY
ejwIwI4hxH47wszXmRQscgbx85R0dz7Ys3tZ/5oHsqlVbDHutFe5A+utybbzWf4Ty/XEfEc7iwhZ
SH9E24jZtuUcdN21QEwFbOWejB5gOSQKiEDynxy1j27p5t0n3eL9vIEcFc9aX44TItfvghYlwiwJ
83NcSOjFm7PfoaiH+3dDKSSiSbsD73pH6m1kbZQYtu9Oa5LOi4cKRbrk8dcnJEmShvCpgAIDhkKO
nBTKpDr7Ilzf5yj+/CaQmMoqdE6zS458fv2iQVTIl6OLQ2MBvTHBpGkeVveXBSkw78IJ+sQ/iavG
phs2qYU2idQ2gLcy3bGjq2+n4oZMoWEqRzqnoLCQ95nDYB9/OH8+0CHH3b3GkQ+OeOBNUUv07qnZ
Y2GE7jBALAnHks854zj0Yv+S1224l6qIuxwEeQCZlBWWEgFo2qUCSLkaC80618gdpNNdCmr3c409
XDPrbAwxHopN8njKmDX4xYNCmduj0Yv+tutfkaheXyQU4ot3SVxvvIQgd0cfyuF258ZRuQtOmP4Z
7cEmn5nKOi1K//cZ/0dsP5BabmOsRX+KExYFimrtDweHwQow6rtsRLOy0RD1u4+WYC+C7wtsCe1i
lCuwdSGYD+60ZYffZ6prWiVg0FHl4abSRWc9ZyPCZcuYffZxxHf79nWh2u12tuOmV6gyJk8JMCAa
dB456mWiSLJUd584Vy7+b54QNLrOTaw8PUFZGaZ6TRUocsWOwqcFcLqvH7l5Y1/22jAu6eo2i9PZ
xCI6twGAM54QBOMxdyfIhW9idQHvbFdHFw/Nw6tjH8k8J7e/s39w1TP0tPehAwZnsXUh73LwECB2
AcNFwOKIqCsJD7zI1P3SH0pAE3CHbcYNH28fiLqLMM3pk3+ggCafVueSwkB/JzMLdctgG/05ShyZ
MRMiQvDI5IU83d17krKD0lqunxcyLLOe15egfY6ucnqufocq4S49vhmXZHbVG3JQMXLHwo2V+rX4
ixOW2X5rRh22epYF2wMF35zzj/96TH4T6EeZdHUtL8boA4MamHFsqzTy5e2k7inqZhGEF6szGIEz
VQmdPZvbWUPriFTV7zeo2tXMh3FmoiS0LOyu2+E5hjRpjMaZie1qJHqG2ad6W/WE+FfLq1oF2/NE
wGC0OLGWc5+OFLN1fxnawFfWj+QyOGMjY2bpON53iBd99qupxmLjzHY9Ko8WryM6Xv7lyxNIpZhK
GL0FqISpxGoDF340nowMbcaUbHisNtD/wyr9MswoT4sNgB63KxbJd4HhCw616ZwT8FO/R4ozCH2c
YI1N3hwKamnp0/thv+ktnprxGTguKrSlKJIlaygMyzV59DTMp1TWP0EQ6dZPsZqnSuRQMPKSVoLM
d1aZxxRHb8nNxkni92r1a6qd7ex4Wo+qP/8WMF6WnRR7nmofs7ADODgdfynOwOHLxip0uZAMGM+M
HfY3PCVZ6Od7JlDZXnUyjY3rmNKFVpHuLTts3Nly/ZbOvv0GRyXDSJ4Husvx/pCPDmdKgAeWtlw2
Vcy2q+v4xf4gPm7aNJK9J6K34q2MWd0MObi3JMzhDCSFbd266R8l84XLZ6hSem+6qyKS/eSJZE1G
gpyqYnpgG4IRzhM3wstTS1R/yy9c9k+9Ux07K8lnxs0vpED/TF39EC2BXLL/KfaVCNR7dmGHFP+n
c+I7yLxAHH5h8j7oExWWRdioJgxhKLhrbaDdn9AcdBXtP3on8qEN65utNn5CRxhDaYPqNJPO9TAi
/+7NtXrJ4PYIqH2jpCIH4f6KXvPsLP6Vd+nXHwUDjOHrFiMclxDXP3QIdqrBb5298G3PfyF5aTcD
6WhixNQkGwTI1mb6IDTdC7iyotIpu3OQYKab0fV/qcXffvVGbFQacHRrAikV9K7yBF8H+E91NJ20
st2JVRSAIeTC+q4y1+4NZqrxjr3fr/IvYZ0P91O8gM4vrq/L89oW7Yca8fshkIcdx9pLfXe3Zj0u
5YPsQn6bQtq9DA1Y7WlayCaxN2Gwa2O6obIuk67QWV48MJ9uYJ/kBUI/zkbeM+pJEIWzQ900Hzt6
p+Zz983Q25+9TkZG5dMe7/RMbcRyA6W8iNycasqyjC/OIMzcbi8CzLhBLbaOvFo0Eg9plpPsnEWu
F+nMgRe1Gfhs3W6PrD962it9Lm6YdBlBOaV1q3E04r2cLHdMiJ8c4jvyXy8sUFdmdl3+XyXkLbLp
MbYyiI2rhyy3+rjXlv8m5tQK7pfpZ3HubytMXjnSrOV3sPhDjfA7eV1ATllgZVfCi1x/w06bSA4u
E0HMvuvdnwiKMnP7+aKzHX6yvAlz1CA/ylAvS+L4gNkG4JEJm6Lpg0lOv+x8awlGYq1bE9k61IXG
OKFheFTTC3asEIv2dSuGN41QHaALW/SIpMnEfjSo7eJ9Oi9vwJKVkqYIIpxISFjjvJVUz1qUfVG6
CFLM0cXZy1hO57J5rW1Puq+8SgBEnb2SjROf0+rDiqE3qZP1RrEOPdqJJwZQzNnqxBOxEkds3f5W
vosZEIKuDdvuPTI2JkDtHX82aO434DC5Lkb0yt68pLSUlp3e+Jej59Dje2KpZ5rw7q/XCbisDVB4
3kfZp4TIUU2azmOTVIrUIms6B04J/ZxOtPJE9QS1SnX2VhR5uqQNAr2YnmOXEOh8IEaYvLlO2P5M
I7hBWyrrL9QzwFj1w0M1R9xvNbYvNrE3N0Hmoqkg95FZ5wpBoeLOsJ606N0EX0csv4W2Yu2wHvQ3
yR3gW9W+hA8knwEWcm52sbFGVuHwifKyJBzcjJzkRMcxOWqLmXf5ADcj9JUeCekAZj4/hxGzprpf
MVsLkZLmiGUv86AThRhy9SJruBDLZu4Fqi0ksAFs704SCDd0q0ZfQlhUzQv3Q51qsYaGOhA2ugiV
juim9WdglCjT9qYl3BJYQtGZiNovUZiVZ00rgwqnlELg5qqzScbFXBovWkU58hV062czH7n6UuN4
S3/nBR/C7MUj2pz2i0WS80Cd6hycFWA5cxKsOpR5yOcm+f5/tav3Q+OUtLrKZd/4rRmGvsm/+aYm
iv3stkUankXfDsXvLVLLBQ7TjtQ4tpLtX0hKbG4i7IPGNB766VX44Ieu7Ek6dWWVL8yevBFAb/NK
SuveKOrGIdbnODpim+dJ16ldddqaq46KflIQtMx2h2XVwGnXP3Oo+urAXWRl9ff6q7YL4jwuq44u
64SBaTTptF/jkaDNC0ZndaARYEBWh0TceCbQGMftYlWx33ejZWHop+ok5ajlCahsvyKwRNOVOumB
vEpYxVEJZVd5ac97+itxU2xj5wUj5NtdzWKhLT7O32ptW6yJl7Dbo4I6tcfCTE+JhUWxWHNk5Gh1
M+ZpR30CZmXpnFvSLlwRGbfVpIyCDbBPcCBT42DBOUoX5/4Y6cJsuMCOs9H4g/6LcW0QNkRJPCIJ
lHp1QEyEYOOVRVlFslpdmJO9HMsKzZiu7F99JcdiSogXaPxLNMYYNIQOzdSx0qK61WpsjLHEiYNn
0NSezWWUL9n7Aji0v3OyEOChUZJl8ZjFgrneTI0RBJmHfZOFC7rrJI2cCx1pRzcVtdL/RP4joclr
rTt1fBMf3KnmafOkdIfHP3sRoVFCKn1w8Fm2gwgQYBjXPKpcP9JY0qyUJLPXC/uo5YiiWBbb7Kyu
U/trqqc7E8ELHPrnLF/COWMttk5sH66/qgYUGO7VKGBoxfMkEyeKVk+6jkHspkCL/NHSX4zMcnOX
KCMpl5FkTbyfsn1UkFcw8hVPOeDYwmcor5YRnorXZoCG45rzA4wdjOHC3CsDcE47uHZ4siUsbrsL
fWFz46e8bJ/b7uYtxSo7qxNeO/e9amFcasASIpBIozvtYVu6xThV9OgXmjsLZAWGYrj4HnNFuQw1
e/g/aOPxsNoutzBfIc51NLGerb7anR6wzOT7Oc4IYFJTH7y3x99JjowvjQ8pg1hsqurZELnj3ML0
PapwhDhkvGc0PmvhZkeymsSnH8vMpM9S/gmgGjU1KOoo27GI7jQIpyHqgQFVWVHh65K1YFf2ipSf
OzvvSQ5L5D0PqN5aKYwCD4C6VcsswulYSp4Gr7gk8H/8kPQZpcXMppyuZPEoi90O5JPB0tPjbY8q
pDkYZ66P7dFDRI2Mci//Osg1pUZpBqUtr26bIveV6V2+OGK5KLs2ujz5ORXJ/nUs0IyQoYLexhA3
Gchvxj8XNipgK6oWYATstPflLHcxV7h7CYGLuELrS8Eyc+QIDIOWXKhV6OYIfQDZiM0FYiR+x9Kg
gUr610CI/F8utlndt+hnO813cxXCLhHaAMalT1OK4FUm9ze5b66wDTilb+gDF/iVfGhOWbYtQavb
yTZXIXKwYlzkI2sKSioIXd5VZu50IXHW0dGTRhbEMNCNwM1Qw50syWmj4JUkq+oaISal0UMzOwpd
2KJFC93FB+4GKoF25pWw1zFN6hi4BiCPuelYXpgzzJoWO7yA+YmhwYtSvWrfC4P/IKxSJApGkZAB
SmXNbWrKg39BWyQA+r1HERaR3dHObHM/AM2BNv9EoJyyAm3NMaUFs6/YFeZX3qJ1oB7j1UppjMWm
RGHgUu7aYUYxYP5gE1K/kpYbopGhOtzEIlPK6tIsb3WDW05NSoOZ+S7SxrQR92IzpZdmAZZG3mYp
6XACiS5j7EpH4mN/q6VvYlm/3/B4rs8++JEDaCP+UUusu36kz41nyfhYiHubVLWIJvDV+nSjDcVl
bHYE9VG12k/+q5hR5NHXb7iiFPeh323Q9oIdHWAxoVYAxTWZcXNUAg3lZ7XhYuAvFH5Je6QS1K9b
JDa756vNp2az+/sx4uFxh9GdLYSgb5nK+mNOaM5zcYui0m00OqvRJMzjw+GzjceixNv0YA+EN6qK
t7VWK/GvZJm1ggrUHU7upK1v6oGt6kU64sC5EMyCu7sTroDPB+z/WnwzaBkzrXcA1KirxrgZVgHC
au1I+PKwmJeIqAO8FMxLYWZc8L3qv+23Xe2yyBawLhOvjFoO0zVdoHQIpip/4EnI2wWRgKHYivfc
zdYmj7fthC5SpsvAyueFAp3IpRxkD+QkTxTBuxqJjCA2g6/EVgBgXdB5voW15ZzQnsdMQsy109Aa
etYzWAJmgejcKzO3nHYvRaGmUOY4YMaVWPfZZQBJTtFQFAarKA81PaO0D+B+KryMcESauK2HzQHq
yVzcGqyBhySy4WAAjxZmNX3sCn2ZnWPvHZVM25E72dAqZ2Lw5mqvfHxJnk2FFeZw1mdDRZdlJ1jD
xwH+LiEtgck0tfBGGcISp8WMC1JSRXsegnk0ZyLgGeLhpRgOjr9CDIZuFbayko7RG0mABv4uuOno
GIOevePXXsxyniVJGL7owwZF6N67GtRedMuMAS4Nlejgmr9nYnWdcuMZgRqZpBWGVZ5D9hd6Otzk
t3R2u2drPfe2siB6UTM7e85ZrYE8GqNaxkErsCs2TJP/KX8nfHPGz9sDqaM59icZ16VbyUIbBGEy
vX0PfRd6J+NTFhR4GdkujL5FeiXparkkwNnXsPJroTTLUIgvEfB6pwr37IfD7DlT59RGDBrnT0uB
LG95bL7o7r3E3mXc5clJPcOaxRQfGlAKI9JQQ8MWWJx5u+7PSWbCYbCfsQi5z1e8IwJxC5rtAg7R
d/dbzjSXJ8Q/yGvOqP0tgKJ29GzQngdiTi2L6WJMQ9m7NO0GQRpPdYLCL07w/ZC7ayrcbUpzWS1Z
Rs6FvoVSWDClXs7h1bo5SlWuS42cgNcd4+gvDTpaSjcc9nfViDbK+G12KJ+mgEVgmDRRRlBYGyAh
atJamlnUhpWGsKlhyfmS6HY9PxdqwLQjJD2sSi4ERU17Yo7IEHnPBcbLmJbO31Sc+FO6lzxdbIeW
6B+F3BRN81SJUq6cAISxGCMaRgeMgf7l3UOh31MMiC6JSUV5Gjy+mzBt9+TWcmjOrPy3WEujauKx
qrzI09JOS3dtt41EssxQZHn63fqSiObI4DHTxvCYg0w+bsl/4ByO07yuSxe9yZ5oTm8Yws3r2iDd
QAZQG/TbhwYyWXrzhlwSeOiDCdLdRN5pfa4D7CcljkwdAwF/FNqnO/yKc724PlrU3Hpzh1prpUuT
QDIZlle5QeHZFuN4ZthFVqi7nxsYmP/aiMpjOtMdsh19uEphiqWcpW/olAUXotG5w1ISMJUzM+WH
aCB1KrYXJQri1Bq2vFOgOGP5RAqPNHrFg6j32rmfE4yadLfYyBYxhtbFaKHdWH/pjUleB5BhsbAX
ZWq6ZHx5g20YN3IzPdXkBUxW65iC52ypiKdSDJB3/raAYKKljLusRhLWT4GXsX8pGi3HYcy3sK+j
0s1oZipy42+t2bsGcsZ7eFEh/GnRzPfTk5gZmCspmREh1OwYUUvZGyRVZTr6F97loGNBseYC+f4k
qdAKwbhRgXxXJnlZyuckUl9wGykhOfaNS0sYxy3/hncuz22WAu8ZZ10TlZvgFHuVz137zVvdttpQ
a9ozHk34IORuvD956/ru06g3U0jynQEgNHy+YyoksAPafeuP3IA5ZmWDwuj2VgkfvqEwhlQlnslc
oi3HnvKsxuXjsxedgYYpXSNazLUXWv+QYBNabuHWrqrzL6M8rLJoxGEGi8Oy/aavOAAupHRm47Vp
v+5Y8aKlOHEbP+m2T9dWIHPKLZ6XRpw+qEC9yZj/nCi65hovHnLZzdq+L9Zm7eR4Ba3nJYTjpE7G
xDJZfvBoNwq1DvJcPFVsCcHr8Uc3IHi+Yb5QIXQNc8wuXiqkAJ/D5reXSOcMbmYJxuwXy9tphjzN
6p8WG8S+mJYUzx5QSzU9c3w7OuGaAszl9hce48f5SPHy+qdCeUCMU4EhTDePTUiPm63QcjCjmpae
tK2tV23yYZaAlIh96+0eOiAwLE1tBJnlqodWwNH8R1iWbvqAQll/3YK9zIyiWV54GTBAcoqD2Pf8
CuncvsB4IrB/MuJuY1JdbyxS4bB0rWcoRlIkOIj5tbZGGYhi2pCvRSB6uifWVSBVTRrES7QzRDJL
49KT1NUYAd9/WGvT7vz0CIuFHt/MH23MHwIrkDLV49zIqCEk1cQQ5/+13wERW5VUERi4c5IcJbOX
w8iQNlgO2z5VBRoVcs6C3YextwbFJHoBiiIG+jKax3JiP3DJ1Qx7Qqta24igtDdXJZcGf1Aj9ikZ
xTlrA+L57JK1Vd2H8TfwFbobROqj2CiV5uFKd7ErxFy1UAqLIyB4JsNjbilbunVXevDZpjnAhK6P
934yBVUE5RMlkqt0CkZJy3OYrqQtGIpoU0mlPkxXRyFiLVsxkysiZ7JMiCCVldYSXoAMLvFWixFs
IWYp509ZTEX2ASqKN/lt1AficskcFP1rbkNHKIqcVs6+Rhl9+/Qn5e4K+4sLMu4Aq45Rfl2fEZEM
/K8DRNvs1P2han0A39/ZOs+hHrc0GJr7x0S2lFEJZUTuSTYcDGuMr1Y639tUHX/QM57Vs6cfukBJ
/mptbBZySqERq7M1gd8Y8n1gsYMWnRpWe4m0KYxHA+pjrQHXYyPglI9Ql79AWm1Fr/g71YQE3r/y
hTrnUcTYEP4NrQgcKIukFO2l5pCDwJbh3ejtz/JikUJrdytGp3bxtDo/nG85RkLUc8dPslm9EDyD
OmB/AzGfKmAnp75atfAaoO9w3HXK2ND+EKxK64X/2XG/z+n/U6mhMPKfBWuc0W9D9weQ1p317z5g
AlYT+ISmRoVMqVp1P/3l+1hUWisSyI9kIbB6Q0CnfoDJISMma7TXj1onV8s+nF43QuovcFUB9WRY
8ZH3F9lMOFOwqEuiqVVeR1s/cMdL5m09cVjNcA0H3nchah1c2e1iVASSEOwwNL/8tdYf3sOlOeia
crTT65zVrhuX8uFRsNzPedzoB2C+5diy9lGwEZce7NHVBmJ+UlRVamnx7qo/XlT1aN0Sci5NQqJz
dVXo1opT4sP6QMldwMJUc8vp/VKvtisFdLoiPhqEpl47aK4tEgyeicbz4EJxE4yRJV/fAVPne3np
zR1XOw/x0FmK2BXNG/SIzmn0lpbvI/a5HqGuESR7IM6pIIkaZPcFGW+W5e6VWRxArOJJzc3iUeoi
M4PeGt8oHAtafMCwoTcAtfFuCtmwMSGqOOImNxK5lDOsvBThJBOqVIwEiGRtB0HUHOhFf1fLdJGu
+OnSVtfydrAifj7wJGUqfBK+pDyamYtYCUan3SCeTVz9hYVKTQqOaM3oxuI+9SvWQf1I+BubaM9+
t5Dr7N8ZEdf4vDQCgdl6xeZQENQgProGuRmQeqQAKOjrti6onbr/o88Z5RPxAZMVqyj2E3cX4h0O
9et1dv3GqQ0x2bds6dnolreq2mKt3D4gmDRYX5fHdVuojQ2PwCwlHylJ54UKGJ2CmrqTpDKWKXYK
atYrBvoT8xrTokpDqnDn6YxqoSUWQHVs17XgR1gnw34aqAj/TTlr8gP86qLoRPYFtAIjARPjCM//
igLrokFKwB7wST+VlOnFPvS89i1UR2BhHKadVhZ6lmqLrJ5Ot693QstVzMRF0/Cwp4xJIfSnVrFr
kz6rtFZ9NpsnB/2s7gUaeL5uiNAVYYsSx/0aue4Qf6DpX9qGmuwE8aqd2CExdYNKZT9bVAp4LzzH
bdzWRaGP1JQ1Zm4PkFp9mDcgqRnyDucSBYqL+u7wk2bjpQtzNBgU1z/WeSTGRG0OCV1rdYu7ehmR
tUqV7BVJBsDFf/A8RrOLv3fAlZej8GVOqqaH6/xpj38A09rH/hoA/aEPWZpuBWNdW1egN878SZCL
O9OqhusWWKs15XiIdVJcgy4KDkEbpWfRkl2jiANXbg7C+D7mtEJxcaQPT2su3iHAcPsUneUsK72I
9M2WMpyIaLrJGEoly5oJMODouDUSX1RyqWfrAS7GRLwDgBnhttE0A8ccpQmlH8Wb6ADQMnE8Gpby
wKuNqz3irfhmozZTNK8XZh5m6UwIqFSTBs+GEqZhTnzMQKxHaWA2gkPUcD5eNSIobKZSVJBLnXZD
Fciqa2u3c41heOy+BoHFvHLo3YG6E1rAMrp4/NMq1mkZjKyvzPmwpCNk0tz/WCFn8qVaVPiJpJ/g
S/qvGRzJSVSzr4RdGTXaHNdngB4gs3aq2ftI61QM5O+YUzLiadtcxK2INI/UfDS61tGl/Ftrb7ah
CoT9jybzmSfYQ5rQWnpACpLpfSBJyb6AHOQnldz4m2YykafBJtKWxvm7wOkDW8R+rNWR+aLLHM0q
bVgIBpO4Z34YqOm4FRf9ivexH188IHGdtvhQVuRsytZIOIZ6SrNBWOPFYm8149jPKWkVYRSXWrA8
17CWGEDRXMbJBrkRRuD+nPRlQ03QXZPNwxUysF7toqnu/pBxKhyUYvF1eLwv6UJ841RB1i6PTZ2H
I50nH7VSzBMHhXV3eTLVALQWefRxi5S8Y2iTx41vwfPtax045ksMHwPMe4BCOnhzOXwjuauTCJxW
cGTPBe6/S9c1jDSrPB48DnOALLT3TCeKj95Y4bnMHovxDWLuZsuNcBXOYxMXwqCy9m+XZjdD/Ayz
imhaO+alzOqPx8cRb5N5apyXypKAgb33Wju41LnkK5VjHUFgdENwCMZbW4V8LeujYnCM8Vjgmxvv
KJGYL73qzryEGrgPIoHOlrh7ZeSOmmRz6Yag1VwqT2uqskNpffsvfM9Ssa2wPrGmE4WJ/JyuV2PR
YExMeOVmbPkW4tJRpMznZ20rIVGpJ4hlypS8Av+P3dqnoF+8HIfIwu2MWMz0SDfe1PcP3Lk/OM1B
fRCILK7Lc9ghDsyw81mjka4mw6iRdXGxw/OQD0K3QchfYDxvS9REnkTZj3X+LkOR2mod939N0WZs
Dm3ujAeLo/nLJ5/kyChHPS88BJ63NdAWDnpBS0mODOD8n2+X4IRl+ktys7Y3MHqsryuSX5ulQZwj
33ejFOFQ5iqhvjdiMxJ74iVZZPPMy0Anc/XOls8weFDE9r2lHNA/Ih2+x95n4/JKUsxhGa3O8JSL
Ixfl9v86VS6Duuu9g0g0Siy23tlF5mb9+O4DI4iVenRi64fVXJxvKd9KYmCokewOeqCnRBlzz/XQ
8O86KYLLjd5VIcQjStglRbsOFtqBX6IvfDuA4nuTif7ghyvpkNE/lflnns6SfF4SvAm3v74udwnV
ypMPMgVudLoRjDAB5yHKidxeHvaw3zVT3pvNETSkknuktA1e/nzAPKrMmgSrG1FXsVHcUGOFJSnh
vuqROU7S9SshUSWKCKwMN5SfFUxFVRlJttjAvAxpK/r6sGh7GWGqj084uwsUS4LdbKDlZTG/ErX5
1Dkt27oR2SYZ8Z8wYW2WiRSSk33Aej4yeWWQ7hNz45DYZUDGmjZKnd0sXkJfXGlZh8CznFWv4319
XxobnUaHWtunNA1FreC1xowQOuBXbVzd7b1tju/qIeNz76keKCCYt7rzg/p6+brq9AH9joRdoszI
d+XunODo+fCJidkwB8zjqWJx1zCCkacvBz0NgRUEzQsP348yOXZuuO4BCW8wmgRSvI8T55LDl4OF
9642IQMcHUDwNQtSnckzkNamO1gF/NlGPwzALw55nXvJ0pLUcipc/ibQofIZEqywzkMG9hiZfYnM
03tvi6xrwlo314GggStbZs4YbC++QGz3td40yV5qntfYHfLPsH0XT5epPK8mbjxIVUk7JWjVUWpm
WilUjNkTxXxOqpsooiyCaE5s6gyPPQ1Is/GfTbRIYDcb9+1ekG5ud2aRsBgTiWirgsUDR47zSJar
ZceDkAi6p2WTEByAzlz/IqCpdU1n2Q+0OjlnzG4LsZiFyuRocPoW244GvhsLLDehB9EIVuT3w8dX
ca+pIUopZFrtTbC8FIgaZfv26JWOirLk4rZ7NPDnN3naQqbkuNESOGqiIUJXczh/K9Frf1989VXP
kxPE7CWh6orYjXbPA3mN5TtFopPKJtVlXmpdFmVqQo/eBXrNSyQQ/l1eJLG/t725YK4Um2qZKzSC
np9vlimvWtKmYNb+I5/yGi2v4e9xxjZPJgLby1EOUutu29Zm6fU5QbEMlwXxZmdeuJy5Ok2a6xs4
km44Q0EAQZ7NQ4s/bbZ6TxFrp3Hy0YCnK/Rl/qMuN6r0Noa4xT3piwZyt/ZreS2W67dQHTfFArdo
mvCY2QZBNhBHJAR4/s796zI/mLV/rXBFwwr0kDswVyW3/3kBUYcEZQ325f6t3xM+1awYNYYJW+vw
lwFawAIa9nMJqPwwRp/IEn99FziQOizwkm7k2z/xqunMWRNXUKkAjcUwr8Ca03L/COFzd/uWmydu
SWr134RtmMbejSohzt3WDzy44F7PI5IrESJEwpb/MvUidSrnk1fMJ4esJB/HqlXhDQdjLcvFM6fd
ayLzwEItJJcnja976elWxYjWY2ROGoJDcE9jZIFdW6uKVU7XecggLybk7z/bZORq3cbvfmNNRn4w
QTfcH6pMg7juEPZiLte+1oAr2dvpVjP2qWyMahGoNG/9+5dYUqS8Qnb0/rTJPuWorccFmkCI2lLv
eWzK7k+VbaUQoYQD487lEbAkl0AyopSdF5N4Jh8m/pZzj3He7AcFWKnVkooP6p/IRlo8R7ki9KZW
JncRm9+FTCe76YVLTHu1K/LxsEdwrKfOkbS6hUOL+bLL3UCxyL0ObeZasosyGCH0O1VetdwzVp/U
jiFzMluge97L0bme8K6sH8TPRj6+OAYd5B+c1QgqRB+Hn2r1tTa1N7PjAe2nylra6ISD+56u9quB
fAf/KjWcMHvFQNaNaJdKgFz6W7TyEeCpeotmKfaXeZL9C2uuWDoCGF54Olljy7LbD/KW8Bd68ZYB
2cyUwwzt4twOxuX5ypxrvELM/a93zdHzQZ0Fdi912KDLiVFLSa68cKaXYGr9yy1ufL33Xp0+kh2D
bt5xkuDX11cz0MCUXNxiEug2ASmx3EzaC8L4Ek+K098rj/cCLddJmEZHk/l8O1aU85SqVgJpVvOc
e5F9u0oLaFQoKVYJabBJ1JEPItLQUCmehzXhYbVjxMJ6GwcDvYQlNLzxdKDzWFSwUVTqm9VldF4y
/P/C2hR4c50YfWyQKw6EDDXh0ykKwNeFLtroWiJKvV1tFi1o4YSjWyU+q/YkCkPnOIAkNtBpD7Gj
9ZfxVspIYrS+vCyTss525WTo2MuoZpMNFBCNax/ZOflg2ytrDwYaRxKGlq7sTlnlltZHB5wRJkHL
YyhiLadoNcr747og/54ok1OlzC42ggdr6nvFX1cinLtOTiNLuug/QhTSdCppSE/D3w0T7BWhbz4n
3iCrZyZ4mjkASTtfPOm2p3PGv/aoFDkQPU6sRacWZB5DXYphJWYXFHOjAqxMvnyLEMygvrkmjlX2
U3Crmj6WZ1FuMFiH/v6FC5IUEZnZc3hqclhpBHZdj8X2khkp8gcgJC05oxl2SWFqsqiuSg3uo9Gs
DBrW361vtoTiNAbYI4IHv3bq9A13ZvZI2OAWdBmE2PTNbaTNQNJrUbVtoAuIHq+AyuJfL8p8c40j
2AgNXEA3td66q3jFySzSVcneoFvnQwHaXQW4kYO4s5f0hpay3SNzGMbTl6ERfIXlPUTYqPCLJ9as
+k4dWNL9/5DOcB3hUJxKLMaSWYoMSMsIpbI5JQP/yU6aVwnN2BZ3JDnU52+y3pxX+jiVqz0C3jPg
fXs5u20992mo7n2vAnh18dQH6lSw1mJwl8eJJ109w3wk+EZETelX7z3nUPBaDEDw8uoG17cGjnXc
IWD/G0zU007w2y+kE9ucoVUQxc8LDINiomW/lQed6ohVz6smhuerquB7Wjc7NgOAZR6+9ksqIHPP
ojGwQPseDvg9TZkSddmVddlZuTOOAhPUAGH8xjhNEn+crV9UzKgT5lrZqbVpQUmg2dDfBN31B3eS
jWdnaiorFPPSthdko08eV/MDF+oLdxka4eZXt5N4xgqItxEOcVU0zR2YzGihtn3yc3ZKhjpMi1sD
b+2P2NyyUIWEHK4PhojgkryQY2vOogWhF/k+F4boGdt/dFAYxVJni8+KAXLNBVesHsiRqHaSzVFd
hLb99Lq6UK+ZHWaBxlnHFv/khHa/fJ/aoA6XOFIvxhekxz1a3i/YwmrccLpw0qT1FyZHoeyw2VfH
rkXTCo4eckbD4yFDNDPumEMroPKtD276BFhEF+AAClQDSUvNsDhvUB9btQ/o7qJQR7G24c8h/yro
N6wiPMpH82nNq7nirLkvPD6TxZOz9Wwa/wuMybzSS83jARwrF3KyY823UDhren3ajOKo71+Btcg2
GRM/JmzIPv2f6fVbLdqArl2dcZjHhwO5DeNsPyETdMfVqtZufG24KfzrapHwhNrZkQ6xTStG6K/b
PfoCRrP2WUSxg+xLa6xTW5pYp/uDdmhAuge3Bnh9NkmCG4KBkDjTQFLPCYiI436ROcDwWblWFuCn
4yWGEKv9GAEyf2exodb5ShiWx5wT4qzSDHPniaDb5Rc8eS5Z3hKynPkBeiKkcStr2bM7uMQNm2RW
95N5AHpKTV/0FfVY28ntwgnb3TkUzAslCGMccDZiZ1MmfQO5BNTmCz7h7i/rol+BRRnBTcmr9GbF
5Si3oWjKYiylI4oxWAHS1e0xQ9ibFZR7gGamEdUbQPKikka4Bukvi6YD7iClFWYWgaiGDArkrEJ1
rlddtYJqoydJ05M77suvbv1coo9eOyPbuZk3xWPHdSkUqtESxr9Hea3L3dTV/s+d4kYPsK7Mc/+o
T23Q9NEMLpzHtRhPdirEJFSGD70adF/pBAV8XRQbbTc0lgvHucrBOU5akpOmyUi80+Yjqy3xIo5Q
8ANbh7bUfg5BS4ihdm3FF0AejoO9TUkk+nF0wfY65ml7VvMRkKQttHcQfXX0MA+M/vicVGsOqiUA
anzS98F3Oh9b0XgSQwZgESALz8d0JN6EDLKJ6nLShfAohVocPfI8PHMcgpBgdI+VytGhNyI58V8Y
EGkHDc53+NyPbneOOHzoX8p3TWEKz0AEbFEhyjikC9J3NqHwvpXmQvL63SAxUTVn6kU+qFD0hgtl
1MqCAbWbSA2CB2HkjlGU9DQkMEcLwXNIlgxmaghRzLkcp84QZqX9ENKQdZNMo1X08AcRhkaR3YNR
MmUu31PCLIMraunEydV3mh8xsQnhIw7EFdZPHx5RDNAbkXUt/GEFQpWO/ay/RJTpUs1K3L8tFyLV
CoiU71qmf1YhoWgRtNqMls+OTfFH96CI6UvSgiWABy/XcaeW8QVWmSTAHa/fh00A0II6vLu0Wq8d
TrS1eKmKtDVxtlTUL+slr+LmabmH3eTqTTSPqvJLlGLFntLs64Tfbq2H2MxwUeKPyW3GeNy/m1ce
pe/ot0Pbn/bLEftzewEx8gibVct9ghBU4bDkypL0U0ClnSMEIR5qFa7GiPg6Y7VwTobEkbre4jr3
lapMS+4m/+tdlylO41SX3tP36SfPyJHJ9SqiBr/xSTHHnwgGMyMnt1M30ww+Dh23zCJFwx56N1AL
juqIvobDH3e7KrDpW0KcYDm7BAMHjCXr+9PcQJPjsQtB0h14rtOx5EKVSVjiTwIQ3XqVXlkXx1uU
3ptAoqMVe6RiCxoiqcK0zDqeOItp1o5Ze1da93IUwgWXfQ90A6E8tAfNjWSgG4dUeqSBt2XEOpio
id6zVwBesQoS3EMrbNTi/JX7G6pBHxplmkT7vALnDzuyBu+ru2ZV0lnN3ung2w8B5qZ/3yn+dkrK
hpg7jrJ5GADF1cXOjXgaP+PehCut/aJAJvZ2hDoWRrpmrX0Sr/RmLMXWJ5d9MmgxVQnJ8oomta06
cmPz7bCv9/p4iHtdRMFigo++2TiWrvMP90oLVzuEl8TsH5hL5xVB0sXncD8NXoy62YV5fuEgGsxy
4zRRDJB/7k6KE11WgzR0oLSoymo6e4lrMVASxM4NY7r9J5tHhtS/SJ9gPAf+9j+AprOzYCJT59sO
SwSP9R1OGkJc2P6r7EilGBMsnh/7bwJuV2ALxTjSZsJMwEUtdsThQIf6egvI0dGhACxVkBoTmd2d
vqesCL1opJ7Xnc8Rx06OkrCoM3rMPVuE6YrJUzEh7g2N189HRvPmOVeyTfKhnYPbCdG/V7ngtlcV
oLZH3erhsIGiUsrPgNIq9MUk9c+1XS6jqVPQCW1spLgdy6cOpqMuxMpeGHqo4xlJtfcyGZWcP9FI
wditF1XTPk6pUhcGfxrjXQ1zJeu3EQGuZF8EzMBZ7H9vn4hT1IrgozqCBRDwOjt6H5x4OgaYVJeX
cTG4/KWSqfY9MrAl0pwqgGmbE1vDesRb9HNto4JkWm2L+ndyIjwcv0R3DGiKkGa00+L0JO1jMJ38
v08eEOWbkP5yXjt2tTJXkIh/LAYZJiBHAGSS+2yGrgpz9y6GL3wRnZPmvGMWbNGhVyAhoQ6WL4CO
/0D3A9ok98/ZyQH/q+c4Y8Bh0yVuwUByr90N0D8d40Vo5qTY+xQDluzQhpAt45M65Z6OKEmIWoGu
BhWd1/J/YvZShgOVm6kUrbBuOgtDS63GPc2NH/WRE6/ebEbxFl63q7jIriJFjvDD2oWWek5/i91H
XVizg6E2jT/N9+k10t+Qsq6xHZ+ROAfGViHrELsF+JhmmrnIRkNXr5hFjitrc/X2zEDhR0YV2IKz
Aag6cOJ2mvQcXOgZ3bVeNEsBwU8XowedKuHlHcRawJ2FZOSQzFVfOjFmrgD0bD7QOF/FN4+mz9fp
5XkKiTbxlCO0J2fTevSLCJpPcEL6JKqzQGqjdpI8Ea7iudvI2FGHqKWMU/REOkisDgnhQzdxRsSE
Df+OX+qHkldY3xNvFJmy1gqZs3E7z+4NQEfOjw2f+rZYe/FfkyJ3fRbmRub7qzmrhPsfunjys+X7
hby7wsAtvxKBcyI5p7ehfwJp2c8C+2nOX58r/il53E/EeXedqU5S913pknINepkvYbWxYSj/w0oe
8xI5u0KhpL8uvx8jm0ZQ2POwkuwVJGfypgAzGe0f/F4EMvswlhhetI6Fq2tzuzb0R5B+bxDe9nkS
QfBHnHfuokiq7Q2ZNtCOsXFs5qpUcmhiQ5Njb4CjhkW3P/ETm1UHnMGJtl7ktlyUOSqG16DNUcBC
P7IQw9WCfjTs+Mc+Jz+EaT4Lob0cOsfkN8QKx+Jjxp8pvB7zZpQa0eATA7hIA7HALkejJbPJXRqS
qaXBXvKEBU1nZo5f1Fp7TAZHkjwDnX/KOMD/ONyuY5F1xrWAtF08EwrnrKSpRsRduKDaIaxCOlh3
bgT6AyiDlpIUIgJybkdXCfreiI5i2jnnh8HAasTbW1c2R7fxmy1fsT8QRHqaDl+wTPgLITKVDpo4
eMLBl4wl9wa5X610SyAOmsFVHMUn2QdvVWRoCmIxMDWNhgefpxkQCC1/V8coPA3DmhZRH7t2DY6Q
CewWxn61D1rdJzx4Wz0D2DEbjh+8nBWCsr7bmrOQcrJrUGmTcpBkEeFynF8pH6zbqCtT61cu0YZR
qzz+G5O/V6WjPaAY/IiT67kmz9X+DP/wyqvvdHkYJJpz+gPOl2W4BIznV5x3dQWSOvDb4CpufxPe
docQn+4qDCJ+uc1pYQ5BZisinRQLSQxZwrVEe7LR/5hd867ah9BdjN7P2PfEMw2GTauFIqdwjjBV
OQMuediKjYTMVDAplvwffFfQ3eCRFOFAQK6vjRVo1oYublNylRo8S7HutmASrXFuZduk8U9/aCCE
qiqzJXVBQG+0Jwg16ATtJ0VHr6hgg+He8jMZ5hX2O4gaKM75wO0lDw0knd4X53hRWXMLdq4Dw/gL
7LiaPic68Amvb28cEK/l8Tw0D1U5SqPuZ0I7RdC/36dUHtjejWW1xUdYyzplSlxBDuYRmKM5ahws
Bc6H/LuN3MGmp0OVlyqPW7ZKeD2gXWwukYqGMTZl7h+pD1LjocaRavyNZYdHz7rmVSRYLMlfRZeI
hcpS7KnvAUgdkyDvHh75s52v0QJ7Xr1nq4rDIRA8KXa4NOiMwrpF6GZl4Yd8A8xf9noqiZqp4n9z
rrnwsF36uT+3GhN1Z+MzvV2JDpw3wTNpG/My38bPaJ6/3pi6eQe4k7prF/1LxureCOyG592XU5CU
2E+ABzXZ9eKvSVGXHXKVe+joKCBkf82cxJoLKEBDAWXKf435xVPYn4Yl0gfDPxPy3UTSo2m+KcW/
k35JFgt48gKFmbGkGZps1R1LYwTy/O4Y1/wkL8BWJnGCRNQLoEUbAFIifRkGYVIVN3j9ohKcnDgV
KVIALggyct2jfq1Vkg6euwNI4SaqxnAzTHf5r3l4prJDxYdwObPv5CqziF0+HxTAyZLW4/a87s9Q
kqqHD6d4WhMWIWM9zpQtoNA2Sd6taImdk0tFI4JM6PPSCpQfwLGvlQ4+dc6IaKbhAha9uXVYlvX6
U11TvA7Cg8C+liEzGe3KJPk7a3S3gvAOnwTRZms/9FKD+w8sNaRwjylwWAqIAv0kbVI8As6/XmBl
X5CoL6hkTGWFuhSITCm/qi32OJG0Wu2FVgfjLCiDvWHmsZIBgW9p2iBK4U13Hjr6k5/33nFPDsGn
bu0qEk+CIKDMJ21xy9ddCiis9sKUu6T6Lsj6fbC1zx0Dl6YeFMlPaVQtxqFfNCHCxL0wSeUTH0Yg
mHNfmVr4dBM1ChtJSiJ9DRynnkKsylszrxT5Ax/IZydEF4IoLSPLqTTbIibPjyqHEU/mnVRgWDZL
JOC+pViR8SzUGOBmW9gSFQ8Hg4ig+7wNA+nhAVtOBxxSizF4AmCJZhaXxhs5eNVx6RxWIW3Jtjfu
Nn4f2sEPA41Wxx3aCfFMN7/qcSdsHlKkbnOtTVPZ+udtpU79jODYLfh7d8k/55EXbHBlEIzbyFzq
xO+nmKvyFfP5HgdR+F0AmGaEJRjzLytyoxRg9k3wu50ehcvmt86LuKDnTXakSUGok1H/+OMhRvzQ
+hDYkzPycTUI+XgKWK7IUeBoFbQ98+LOkuMFZaSZi/Na6Z/M7OtkEqyZ4OOjG2lv43O7CYgt9jG3
xkC9RJH581x2sa+6byTw7z5D+bNHftZgSLk7tIQcgdMFlyz5Xds1rS+oxdNQZrVBm7BplsW9DZBW
76MtkabblsDH9J51CgrpbWzEHnUVLhmQY3+c2pKnsMIKZ6Wo70npakU6VS5u/mxxbeqxk90FpBnG
VmwIoHinM2nOXKD3FzlkKb+/oAzZYUg8JadLQvteXV+NintlvtyAH57CTQQjuEc3W4iZHxp4f7I+
ofn1i3WvJqO2tSTgwdbUsV7qH15doYep12BlBcwwTBSOenHgSd+ID6ZZ+Zmh+BWHej5oJufzzMFJ
uieREJfrtJuYtqC5gdrONKdjl1s6uXdk/UXyTAX2z+oFPATT5a9Hl8RX1TjJJran0+x5MmvDQuwx
FXyyLNDHX8MQQflXSy9a0SKht4vA09utCcK+o++z2quc6rXJSttod7yqcmfeg3dyamM3aw51WZeV
P5ybcfaMaDwZXCBXEGY9V6AaKAOLRwHt3ohpLYlVxIsJd/+73lrKAUI9SAiis3b+nxK/T5oo1KDn
pH9/vYsYZbV7dvQ196hA/JMC3sG3anILDfTyxgk8B4r/klsz5PudBIbIAW1/SA/d9oQmse1MNk8F
M2rL7mGA1bRV4I9Pdo6JIbFfcqr7YaQkMJU/MVkBnraVQymUzphvDMrkqR5xSs4sCgkw9DzzUKZV
e6BD/jwCu8kbT5fabkm7Rl96o8BhHQmq2i2Ft7JOfczdnaGaQepinYqV4N3W1L1BB54dyVYHtF+i
O+303vZPE3y0DYcrfXB5WzPP6pyyzrHN4QFBaGpBcNLkWiactBF3uO9LYwmFqOcJV7VTL7C6md4j
q/Qe2OsP+fG5iHh9nxWdl20zHc+r2wzaJrG54cXrSDXqmSaTmss/NHPSJR6QnVCX7nbCMMpIxpyQ
5ParzQJtJtn86IYFr16ZnhHxyQ9ZOfr3/bPhSM60uS8XfSQBS7bDe2dSifzx5MX/koDWclJ/BbzR
cZrElHu7tWsGZvHTshSUeXHtuyxeOFb0J9tB1ON8Rnc3QeAdDH0TxjA5jDzHWoqgIZPUmjh49Q52
TxsScKXFCjrJpBqEKaxThdk4QA9xKo8pk00y9YsRf++YjhiVlzArWwpWy+93fAc9mNns2henk1vG
K/I1xwv8cRxA5Iyg1zbqt/ilCCLFF5XmFd9Hm2G2J4mbwMrefsuNZu8BnPfaOEkMLQi8/Ngz2NHg
/7sPhGBfrzFGXN++WcyqkEVtSmQp3guthVLiPVGJqDMiGrfLMvrqJ0P+cJ/tuKw2Sc68n7YY5ji+
p5S4SEpfo8LK+0+xiOWGx9odWU7SI6XvpPgWxGMYuuDWHu9D/rJvYDxgOytMCDqwvwBPQhanOmoF
Ml+Mlp+P7YVOoW0j98RuAvhfiXkrTg3Y/gnaM/o3IT1MaymgFhcsxOEp8G1EsZQaPZ3Skyn5BKIO
sQsWy/9rLs4kBtA8IO3F8cjVQrZJ13dh9soopUsHRCzbC5rLYIyjpOsgvxMPK4HG7B+1ZTzGrfzn
hRmXeGRssY0jvA9sCM7Bhftjwq1qMTddTb1yKjmC8CTjtW4h0rKZWmIKsCZo4WJJ0UI7cvs7O+2C
gbemj8+0rJE27yVnX5M8hDop0BpTm7aAumN+TKluR5uOxO3Bk2fgVlNrQvhXI0uZTph9mFkpBgLD
g42SMtPgG1+EtUTUUKvamEZmmBywgtvLWVQwwm+yizRqO/yMaYFqCuiDAAI88hrsty12ANPQuCrl
qKKLSzn9cPEauYVDljNNhQ4oq9NcWasJriYCxLqyelJb/3yIyiAcYjPSb2xHvFky+rwptlEB7fk7
KyhLqBNAKsfoISC2QEd/vNXlUvNhPBWQcnrEWzba2+x3TiLXltB2+nu4I5rTtwZBsMFLh+GXc/gW
QfDBCNpxkDtUmCi8G+spWW7huoqAcC0gNv1DvzF0JpQI8sIN1T6FaUTMkTz4hnOlnYkkHa0S8H69
BvQwj8YEO6rA9Gp+TtIAd06fGYuOJip6yk+eS0KYa+pKaVEd0iJrT+wiPtEGziKVkrJG4TVvXuaV
6KaHZpW1B1f8wqXRFa2Jbcefzlh8crE6AJ5/CuoVY4JE5Hdj1Ya3LNi2XBOFD6JhokFoqiDRcIl3
33llCRUg9n0LI+d5YnFXApLiyQV5n1JXbCXXucinisdTb9oxYPVcqUgj7bwEtniNFBvw+Bl8aYM2
Bse7s207vJAmG4usOpJTes7h9rKCO5a6NODxLaDtrtq1r9Gox5pU49outljS54k/lp4l31ujqrNI
7ocU8Cw9mBng+3rOQ8rJNb853S+1fQJfQcdHqOUz1SkbKPiZQaXH8AxN954RlbAyvDjo0yOBB0Sm
tJVUN2K8ew0v15UNXMrvkelcIY3YvNPER6L0YkZmovmO39CyyrUJp8CSEq4ys3TU1yTHXwo00A96
zct8jgD3WTZE2+OHBlO7zGGRK6DOZJ6CU+qt8k6iwgSR2TGZm7lnruHhxiLQEjPAwjQp9ptqifcf
R3H4FewAlUvBUHuTeaLv14uQoPJ54NOutfz5qA7tUTjS8vejdG4haJF/9xUs1rAYffPed/ouEz9R
L0fb09K+fiTYZTnHv9pmV75H3rlVatDElsZfe6Hb+U8Ew8/EPHQlsVrYG/dCBiGK5gGlQ3Zm37U2
NL2PW8/tw5US7MF1ehhIWsAfEaChKY1SIFx2R3pcMcGhEq3+4dDuKOrnh3x1rPrnqIp+izV52gLi
W9a/PgU+ND251bG3gLPqXuqCrdqZLc4ehl0Ghp7jyuO3ff+lqyyqf6yj94HFl3iBeGCXANH8mrEO
jhoiRunKNTpcXQFWhsEa+4VJoRxLQ3bxo7kGniu10Yv6WJhQ1DJff2EtVFbkxrBKzTa33bD3h3Xh
YWAdsYlZHRJZxkVN09PkXcsoSyabrRv3Xgn5Of3QY8fCDySRUqDZOeJf7T3jBUEWuNKxSoebeo0g
iPTCX6i+wktZwpfcbXs1/3D1ZicNgHkp3CQxmxpaSm0sC5jKXVOEWBptTOKQvk0GpZHjpdZ8OcBa
XTHlKU6SqoY1/qcHLbae6HhFWQWvJKs5Mjxwv6osbh/ncT1AQ3O0RNN/Mp43hx6eo5XHNfNs3fzr
28vFu3c7DZjvO8B5CgCmVWl2Un1vdt+QE1xAIt1i2stJfwDzL69Hy8dh1zGPkI09Ui4EZCm9dewz
kfHqCJKRwPuKHvtnjYCDJBSlsmndvzT1iK9iAJWqhoYNfbTNckNdYUbZA5smVmAOV9uY8bwTs18V
XjHYbjjiyUs/JGbhmZlB+KQUCCbo4La6VUX/68S5J6qLerTMywFJQ9y3w+7Rxks28Axr3i+tb7rV
DSNbo3VMQ0CR8WVEz2FNvwBhI8O2exOQWi+wc5l9e4qmtmMY7Y8IxhZlefJMEqEOQ88jYa8DPPrZ
ykOBotjFLVqEVEjrripCfg6U47VyOqnTMPSRYU1MJHgXPA15xbGA7pnU6zOQ7bcgerPjXf8gNBXI
3JNuztnhx8ICwW6sWkthIeNgYp/1vGANSN57qLWl9oxpy6stKwnGVs8/wNNxHxlwFZrryY8KIHYD
uCy1TaXBu/4HfcwpSKLub/PhsZPP8sHt10S9zgOo5SpXB356nWqB+x9gZmaMrWnWpn94CYL8LsqP
rIM6FFMEcY0ZputJgMfEvwqTW+eAErT2BuW9a2e/zUhmhvpoi2md7etbuUhkVhxp0rzmQz/9/uvs
l6ClTNCNEnJpN5HcqHItwzl5Kcs6Aapvv0oKptki5rr5aBvczqkHCcCEU3Sy54GTPVRk0YbKoG89
/aLks2pGeBELE6pdyj6fyQ0OnoE986Zld39VIIy5tLnSwT98Fh3ZwzxKvtp6h8mekvhzQzKrzPDJ
fchPrQ0aCXZ5L3Qhg4WnIbWyw2XDKrm2q85mc3mjnZGbmxfvR+Kz9Yv1ArHF6HEf4WCh0dtwwG84
IizHZwtDcXlFpo3Ukr0MyFf934E16FSjJvBlhIlPmq8g5tcH4z97A3QdCLTKI+vB1J2k6dUQ+xE4
EFpdFHOrq1ztK3TuoHbd6XmONzMc7fYjXs0mtQc6CVXsd2MLU+Z2ugLmsO+xj3nMFqwRr4hPslXW
UjSku/M7Kn6tkUlpTUHTe4bJiofx6PLv1+XHBG4/Vp2mqzHzzpoD9uhWZH1xCZpO7De6P1tf3dpR
TZlyNUuFsZhaNkuh+v/1j93k/vBSwEFvrMkAWiLlO8UTRuiXpDfKeRFKefcK46ipH+zaswRtLAjh
zhuvz+9qhyGIxitJH1BBtJJdUY0NefkMOKNBQjjFP2/MV0/jQ84EcMDIOfECpsrzOdYAvdQE3jkj
0Ek9eilYVKcAWxtgUfqumHSlVDgsorGtNCyZtWv3/EMdU/Eeq+2LU708r1CqRM99i/xNKHc+/ObT
kDI5GVRpWTbDHhoFe7YjMhChLZHAR3n46kZUj80UkNpBTUaeznNSzYu5gJXj33eWQ/OddlcBuy3L
BYcrqR91/EH0JPupDItG7cuFXTRolbirdDVMbrLngInJyjaTm6ZNy7qQ8YI5mH5cQHftWI0ONKLH
8Soh0o5XWTbv59B1MgaxDUyO89cOa3oNDzSZS7DabaUzD2IEfhSA2e0x389VJouYXXX/+7FTaWww
8KfFAr+LvyfUHSVQXzq3ntaYrr6vV9kPInnMqfgP8b0ZgrwT6BKYCgEHVPjmEJQy1fahbTyFXo07
4PIfTcuJByVEQYedx/lOkkhirhZ+k/tq5Gr/SMrnAmxV89CVMWllm9Khb54R+lA6S7d2xfAtUCA5
tY0rnvVHkw4dS7USsUjYc50g++IOnpnd6fqSpU40OtyklGyctCexC4H2DBedPEyBoYLPCuVHGXNE
vEyUahjhFzHcmNKQAfQOqnkza+Ag1RYObLvRB053E8lWOauv+ZkCdRJnrvxj50SUzPYWCKMeg166
sYdrvSotmz2LSeSqxJCd+uivDMgXXthEhATSEECOs3trz0PeAY3C0/3UkAdwo42VfYzMDDvkuNeO
7kLidxKA/NN6Kj4G1lbtAj6CdohxLjkpdDOcNCKbMYrE8kjxWfJln+WyedJd06TTCACGnkr+apob
FakHx2LQcmVpUnix6yKjuS4ZadUrsBmkeJZJwYiyoxCMoUBd7c2jXYjNdT1EXsYSNt+lTD9ChuML
uHSdPI5QmbNm8GRP9uwzGZ4Z2toJo8Xu5Ry/eRSFzPCiy5uGxNJsv+6QwmMFJFWRgjD17dOuBSCG
+kSByUyqGiry1PzUkIuNrmB+UjqwiXsO+YtVHsCP7x8tu1qeaVBI01tX6/yHvyCPrdsv7U6c7fUf
Zx53/VzaSTATjmsjoFKJkw61DhydrGNwkekaSU+ZZ/VECUWHDZXmo9XFuwPN1HCLnXewxPpmgMex
+ixnsw/5ll8Th/mFRm7JNx+ODgJrUD7CcoGDcMK37QY8jYWUikQK6AtMhtqWmk9XY/sJQ6wCtahE
xw1vEiA0nGRt3R7H7JLz8h2KQGnOBpGU+6E/6pEis/h7AVX5Z3VXyRabbxZoFUuEqLpUfIBLHQy8
d2UySbic7v5iykCp05UOf4evXZ85jjGIltIxV1sNxKqBD3zkWD+/S//oRIh2rBK88e4qF4Ii1t8r
SuUAOmCSuJBCMteqgcxFq1+1dSGm8dlo8XIMJrylY4wloPz4s90rgKEyacC4vuB0cW/++99DYusE
SuI/OjsAXqMO2P6Dc6AcZOKzx+P68UmVuL4Aj1EGCx/k+aybl67v1gjYgKtJqBIR/26oKft8rG3e
sh3BS+yidLmsUYbi61+ul8hj20HghT1ktQ2k76hVl4lmQ7c3FOKrvtP2Ieo9Iy66qNo3biEnv/fa
WXo/UcWQ8hne0iuY8+/Uy5/8mbVotnVsGeEL4uQnh/W4I327GFqzhFhLGxFCLLo/i494ZcPevMBc
3ssZsiwP0eKaYk0YbtmXcimoSlgVUlo0IqJlBjXvclEMq9Ob8DVme7bEQjnwNP5ggnybEn64O/cu
6CcTlDN/VpeWmeRSjGz+UcFk3h7v1KIidTX7RxrTavuno8uiCV4NJmpfhdwyaCW2MH0+7BuS9d1e
pFguGgZOlHuOkuZhMShhbm2TQkybabfPDFH0FQjMzxEP+iaCPu3GHNVM0Rg6iJUT4C9qApGuubEj
YItu9YGB+RwwmLk/mmF4cnMuoKRT7SqStKqKYCZgn1UBzDKcm+5yDq+9Anzzb+RBhM5rIdFMZsCP
Rqn5obUKvJ2lFQOSMe48icI4BwxeMQMgkdWkJqPEnAiUa8sd069TJanoQsW8sszI+Jnyr8sPzj48
NRnREHHy+IzLI3t3S0uou6x3kwTaVyupngIR2uuBvk0avZ6sVxFnzPg9EuwyYefUJNIaHt/bj3Jd
N+lMak/ZBN4dYav5EV20uUuqLYXQKRzVrDQ2ID+xNpYcXQH42pEVOF1BGkklOwZvZRzJ86RxgKw9
Hlf0hErVghE3LtXDRjtgoY/p9GmdumeO88pl1K8A0c4H41sfZBm0XrB3OOnd3ojPJ1/kR7f56eOu
Bg96MKsGHXppJieRI3aPfgnTerJhGovGnjR9Ab92ZAAEk/gUu4ez0anjYXiIwtbZmh0t5qM96rrV
4tTJb6rdr0dKgQPL6yYmcCcE7+aO302ws4EDtB3w0SAocvY3U3RZzdvfeXp5jtL1pWAVbAtCiLnS
57zmNYTTD44Rhcb9GtKkIGsHPVRUaX4opUIlHWTDD89MqPJiYKO9u3tkBlI9ekII9bs62iGZOQKV
qpAG9rhvhn1UT55hOaTaf1su5vo55d1hBzpFQLvzLwNIgQ1Ecz+G7GBGPYXW+66BtfsJmciG/rso
z2fayDSHR+xLJDs0cPbVICoT/xvPorZd31MMa9TKtNKVjek581YLQFEPA/Vby4goHmwyfwCLwxFt
scrE9UvDzEtf1NjQe/RsLrMM98LoWWLzvI286n/ZtHVz1gpv9P2d/aR2a4iys9CxCznX/+rBYimA
srcW6XOBkDx+sby979P5f5QpgNftul3m5EKQ4xh5lmEX1Vhos9yPEf/EM7JP/qKF9GSJ4XaTDmTx
5uWXXt8GakLOcG4f56mo3doZnO9FWXthqUKguH+yMfKuSA2Yr5LVPjUUjoPwuj3Y9umzEkHMKtFz
4e0Qu+tk24ablHh/aYfww103y2WWURUCoMs5t564Zf7g1+ia9eTD2UAVuwvP1ajTLbOJGRqD1gL+
pk63EpVEh0iG3flPrcYXCw4FJm24s9CMX6F1cPk53HqjbaueDcptmNywD4U4b///1xROJX4143hq
BPpWorcmZsYSD2tkwEfeJen4wAg6uKqhQTRxZLH/R+KxdjIgqAof+Xb28v1q4EIA+XepSFXobqI5
tfyttaQl2b6uPPPxQpcbjVGJ1BnPtVZXPYh6rMxPcbfAkzeqDNWBFhqwa3QL/zmeWJ/iaKRWKwPU
4loBXIzHMME4+9ylA1GMG51kxdaxqQrVr9pNixUvi+JXVqZC1/wLqs6RmRd82SXQDS9Oa5PtC7in
BvQBXpbOGJq5+QYUiU2/ZzlPOfWjSxddg81FSOFvAsxXGWmpi9wx/C26rmuta3Wa+PYSVKNTtSXB
09QddHHSNqvXOrYbVAXpZsQzdbcK/KcEcY0RPVIjBVrtPwnrso43VaM8jp809aogi51lnACOB4e8
fPQwxBlUagCBRkb8CBVkELPJaECqPPuWHKsQbJ/N+mCGHl/E/12UTL8K1EKeFhyDUtdQmowvRMIb
2M6oKS7OLfa672HwupBKqXL3CTLBUqQdtS56Q/KjrXmIlP/vgkMTmGeoOdQjH9Z7aTfGUTT+93v8
Zvwjn+iDhRWL/r6dmg2Ii8J+jhfa9OYrdid26se+JurYoyi7kDsOHcl8+O+TpJncu+T2u0bc7Mg0
ks+/XLOHMkIn3CSmCVPtFRvGcB4icYjL2Niwfw/xeONXT7daiRsjxk08toY3A3qmdDcX71Kus3+q
GA6lYQgaI3mEcU9+XRXRHhfLlZxkUTBf9RRF9pOgnwCWQCuPSwT3kKwayrWdHXXgQVZDzO5LXFv3
TL9PAQNBx0BhcUDMEoeLJVHqeo6ALnUy5oFl1FRsjYQRfqI8rDs/pQnv0+EaUXg0ZlZ+cfmoFVu3
/7XfVWdv9ymisHGFDYX4LBBs/2cS+Y2p8uKVnXrBBKazPHA5j9unHIffEIJfPGYsUaaCc/0eQI2+
NOzi4FGynBVQmdW3Fb/wbjaI3wJIbs0EJt2J4gDNHIcD9ppRTqoIIdkQlFmHrc9jHg8h03fbnss6
x43UMeM/JtRNfxAFvVe/7UPNdEYwByxVbKddHUl+moU0LVK523L7Z2Eyzp8ksdCigTKlEvZqWncr
pJw/7nwfSHO7F6ey1qeUmahYzLdG4OWuhuTdMvRO50WeZ/GJGcx6ZatlGJECgPAC5bI1RxB6nUiC
EpfChqfPQoe1IYiKd2SlSU3WYd/ZQBYxQtlW83h8VoAhuN/dTpYOFW//WteyYQyOqxUNqdZ4HvGY
QdC6JmqSmrFpnyPHqOK79iu4SVYl4YRxsbzpBzTRTUC2/iMG6ERTxJE+36G8j3MG2I0MRnKn8yge
tyrQj6IUQiCOYuvl+4jJDHskOe001ivlkvy1FNefx1eGvlqyw7iiQrKUECaTFJNCJnPgTFNHKDte
R/iitauLpjfnkvuOr1tAJvA8GLHynS2fJhvgy6wBzIMgO7KXJZ6U11k4FjK8Jazo89MDWY8CcslS
IKFDoRLL05WieB7Ho2yFzbZb0m1SLjLYo0/fU4QktxbVkImLqM1ar1RBrgMm4uQVB0hBr58qUqRc
XpiXf912Deogd7RWwWYabPEGK1lAXA44Zubv5+cboot62Ll1AprRgHdyQcNkD3TxUqJjRpHRljt8
jGnKDzHxm4R9BpT4GFz6zR0YB/MF5A3qwuvzcLeGQfWtNaM69Iu8St+tsOuB9SUvUCrj4LiogB3M
QzkJyybdPsnjKkaX+X0Ol4bc0O5F5F2A6V+iH75ag1Z9Rr23MRtcisYmHMuNriWqLA3Cxyw13EKp
xVZQIvY/CSRCdnv++PgehPCXG5aNq0gr6eoZGhXNART9X02vHFz8My1mE55VGpcf/4R8GCzD/e1P
8dHkpASiTQ0fUN8zC0w4Lja4WLIGV6cr3Qj54KuyWPHOj5Bl+CU/fTh7ahSau+9mwrFb60XXeW7+
kuT9MgdzUhxiFCXW6yYCEEIDW3BQOB0Ddfq/dcRfU7C/Xs0FIaCxWC9ey4be/LIny9fAyObTUdTh
qrzptbNzk7C2BqMvte6rG2AyrXndCT0nKDA4M/3JlkbZhLG7fSOwzq7ZRuXgkNtsg3fyhBqfrUy2
8pZzZgRoOeXKq6eQ9S61/oF7WboN0dakkWlP0gUFAkOYI1wob9KYJnVj0JrRQtFibNy8wS1ddhgU
yy7orep+YIg5y1JE8SQhSeam4Y4TG7nnmbIzAjeuC4EEjE8C7tHcW/h464h4/cPDz5Umlm7ViPmC
paahJCnA8B//fLxn3cxCT693+zjApZbu+zOosZEwAwopjknZXh52zWUcO46aq1A8DqiD511Comsh
CLyvu+xCQUNd7gM1ygUN0/6xShZiJiTrx8o8nfyVbQPMcKykGrwTSvc4wF9v2KLl6+iJFcb6Tfrl
Hk7R1aIxFDSdXYSkBRRGcJWHfei6u6q5giyi0dT32VvFs/KQo0Pgek3yI1MCEhbzP8d2bpDFL5T+
WqReQK32a6U8/syYSMH1BUncwqX/PhJ7s/MQgoYAbzMF1NcjVhp6s4ScBFr0HXhRcFCFUG88I2zv
99ElfKEm9vW84yUB65122wHrGgbZcDra5+UKp9N+eyADHXq8jWr1cxtd6pivGiNLovoqefEUfOUF
lCQrkt4cwl6Xd28c0rgi6Y6B3jaAt+J5uVZ38LuIJCcVCwAE81jAYg/XWr+YzIk/+6SP/nplgQq1
RgY9LrxNHyMlnWjmQLH5tHiNM4/O8DmWKDaMiHabH76F8I2/z8o2ZmDlTKKli/7QucvTw2a29V99
hhbUX1qVCMDGnPAPAdr3bw4SMr7XMkD0uErENT9l8E9/KZx6GpqpJbiKYyAltk2YvK+3FVOcvK+i
KQDDPC7kYJinGW07/3lloUYPy0fsxqhMkjugdC/raPFlLixEc29f+G0SvxlA4o6VrcnVUJcyI/46
6dtPMRhgMA6cpYTaD9AEz7Be/w3IxCdXghOZ08L12qq/+OMDPsDPNfyhjjHo1gplWi9GxxJTPEX4
t/AOQ6bh+cBNUSNcyC+lGHnrXETIXtyJMIwp4d6Rpt2QK44LSQkHNdDjiBkhS0rxJEFAGG5UEqLr
4ZG11qkZAvCV6kTLxvHlyyq3Thn4npMPrFEWKbwlcaCfLTzHjZKNK2OrcWharTwP2OglGIF2pF8p
Eey5S/VG2bR11DWCu5tZWFD2PS1s2QXQIDERJjeRzIIB+6+AhS7W5mXETAWhGzVSJZnYV+6U0qoB
Vc2JXPSvW0wWBpMWxDuqhBh4rQznCp04UAruNAuG3JPxDhq7vGnEcyviXKwwAffLs8Fe9iMITRYx
0x6To1UEqMaosQ3/sjV7sy02x2meqggH0Rxt5llOX2pxI+DToL+j7TCCTcBUkZ/w70YIArbWbrG7
/sdWoaYEmZ33tAi26873d/cMaPUog00Nh/X4iwKC+p5fNBlDc1Kp/7gmZqldjF+aeKwFWXTViSTY
l6u6Vjzo9lpltG20bJ0c36gmYKXt4AcY6dBkrE3TLGumI7EbHZ9fmJWxORRUQTTYNZthM1ymsxTk
fmrKHxlwrZ/P094CnmwH+dLRJuRRA54u/nSX65IpvnskX5PW3go21tMzb5hLZUr+tWSkKzoSzg0v
fkou/RPJ7DHMjXRzUa8VLF8EIemQjZtMvV7vNJCOLNRoXbMS9VzoKNe9ojvkzsgy/hM3r6rqWt/b
sbUX/E2cz2JCt196QC7elZFtOKx9yMwEanZsWQ7PL7YcXrHSY8RWsM4oE0ntc72RzWBjsPPAiCcs
HMUSUUlL3qdblePgtrMMwnD8P4HZJ39AQ2WnsOhB9Tohn4ky9IR/JRQHMMrRGJq85mHdqWl0s7Xj
hxHlBKJv8jRpFZnKx5z9FGHpdYiBuF/F3XCyt7XkeNwkAzcMUqmqtgVzun3MNsG2cMNcyk16YG5q
emqpiMSDzG3vXZAu8UHQ0idcM6smkAKCpdNiq5skqlDA6Vx/bA2e7Or7pPebIIveNVbweQva2DbS
3xv1LALu3TC9ZJdSrhdZt0uMxHEDHqNLSGuqUdAJGcQOcIULp9ZLKUH0bk/4Y5INF4QizqN/4d+v
Mqfr4kABuZRJf/EWP/I/EHPvPrOPeOWcPq8nLK5zHJIVP4cfuL9q1LBccbPtfRIbRXcbqBE+KW8H
MHBkhcw0w2FyUAsmWoQ9DsfKJ+Y+vT/n1oKIAetFy6R1w9gBdG/GlNctVa45ClOnhfinMWQVndpU
TjsUD6Aha3QloJLqNtAz+XEMZcl3/VYyb3t3xt5UADxXESGDZVFuKtCcSqj3CizATk6aaT0syke1
YvDLlAHenYvtTE/3tTqDsq98lwRJpqGVIttRO2uUJAPSgMKZC6k4Mc13bSJhH1aVVtBFDmggnLWZ
pSdADSLkCsE5Il8Eis5QFX+/WFiPiHcW7gA036jmkJ/Lk13Hx9yL8lITs+OfFjk3DZQ39qT+owLS
937iEXezUDZG3I8bdLMUxMjP8Dvo790roadWRA8crrl4KZtswctbMTQyXZH9RsXXpqfX6CznzBSc
sCmPbLdvo6ukacXuk862lagRXvNUlyEQWN0sXhv9oYZHwoGUGthBdVyEZx+AOTJ/bZzP64QtfUha
SjjPG9BJEoPSi+xMh+Z9IjFyVgx6jhoMnkJhT2urFsTJJxcSlTusBJ6wvQySgFBN005Z1UVJTj8W
jLvt0xJ25UT5/hIenUixCoKLyeYcnP4WXVhIpQEMLjs8qf9z7k4OWR0pdF4QJyS5MYAZ65LNc+5a
AFfvZWnHda+hwlzWphOrHSUxQebPQxnqo1I9qBW3+gmLpl4sDhBmH3OXEGDDNp+gaoy0g7nICCpM
4CR7IhEQC5ZKShUiQa03kS6armgTxAyWMCBCV+D6F+mMI0qE1LpuL4PKx/OINFyPL+tkc6aZEx0z
Rb900VW16Hyj2iKebUbqRG9CbMW10IjqTXicBjtKxMDIer7xuSKdpKS7aR9k8DlH5V897r+FHdPe
wlNX6wObvm2wjuu28L1x1rnVIoPLellXMEJ7EvsIae5NJXbHPnfKYxQVPfsskc58Hd68kntaQ47v
8x+sC5fp6AUS5ed8pSugA4RhJ4ADmCOkA2094ERJC1GxtYMosCOZ3HirwmBr1NCOTeX4k5qaoiJX
LpBbItFvoMQErpfFSmZYEGRHNU2EG7ga0QTcr/3e9WoEhiqcJ8RP9+UDOVfLfaMYoKsa984Njvwo
JaFxaRfK5zpJ+orjhrl3f8eoID/cRi3VXIBiJqRhOFA/P6g5KAxPZ44EUwClyUHI7A/b7CWFWCMA
5hGgpY1jWFtr/iuWTWTPFLeApQkdERLsXe0566D/SSRZmAeWMb8xtbW2ztFB54lv5xOBRRriTWgl
rIM98hLlVeAZKhtZZbUIIkcdwALy8u3r1T5PpnVLUXFhBPMW8q+mPuJ0VWaoXTvy23KyW+iOz0Rd
4Lz6DD2x5QdzJSt5WNTxYKcBzrn2aSai0O7dti/5SzjL7l0ej282kSlOuyeqsyI/iTkaf4hbl5fG
ZAX5K4TNkyc/zB57sPS1st2x6EwySlD5NRxyoLEO7xr2FIPv+2774dau/vuyRaXa7XWX7NsSyRm3
pW3ejLy1h0OXk+0H6bQuJ7LYSQblhkLRAas9ZgkAIvodjphia4b/exP1GwVFxYYLIx80KTK0XqiW
VHOj700PSekI6EE/CoBKChh1YwgzW+ljPtSx0FkYxRD22Dz7cKRXZlOZQWAEP1L3d3sH6xRxs4hq
7JTMqYl56+KRs9oPHWxlUPi0RPnVZmMR62a23M6ezfS+6+7pOBrDplXNgZqVnCQ6vKggxxmmhNzo
eeZix3o7FOmKV9VEsbEjtxHQECRc6T3n3Bs83qx/EcjBBE6WiFw9yLgu+OQn5MTReeNp+SSLjCAl
496rE1yCaG/iFxNagEucLVvfZi0N6iD16iX2w3DiLoEtKmSO+M4PnoyvpzTnTu7Ae67Q+E8vzgz9
8RRAu6kAqjIz+N76sK1UkKJc9z9KdqU6jELounHZB8FlJFPR9upNNUkUhPE8Iq4y2AxQrLoJ7t0o
4o78SZSrZUzTojLkBCyUM/u1l/HuHyTBJttTvuLUm7ApFoBRLTQhsOD6BzcJeMOfutgzj2L9u9LS
SCoecwok4a18OGZa3v7tZgdnEyo9bVbsdqzsMSq3zwKdM/xNCqmm/Wi4IyY1fODqgSojDkCIyZw/
5CAoX8wCBVX5a64vU4tyU2GH30mjuG2eTvwuwvmVgFC9tywd9fMbTkjO1ATKbYiODiHbTaAymIb/
Kolpgg3xtYRYHE8w/UEe5yXna7mgjX5kQ+phz9Ehn7g8WwC6xuCuVo5gKTLvVJeGOG8L3LPPNWBp
AAqOSJmIHakk2Q/nZsRv4lHNEOFeG1HUhQJ5wBjFAle/Ns1VTxx4BmQlpqMccYteF4/mJeuP4o9F
FYyKcTJ4X4WdxY3rVE3dlLlcFVe0Itq8IXZJU8d21vBRRosmmiThUkWg7gEAyqb7y6dvP1fDzNSJ
IoWzHw/Jn4Bt/BhJxRCfnOX5No5LdH5JAWSs0jUcDG7aLWIt1/dVXBAnYEZNcZWDgbFPPfl53CCm
wZgaZ+wGT0YEX+8q2MYrSWCKjt0RsIMase2lxWjEAbItsAima+gL5WqN/W3oOCzWwfxEX06bN2H5
MdQLkqoSRt5HY4bBJS5WKp7iOU6wxIab5MpS9YMStmJwVkMNAtnC7yxDmLUnbun+C5etZXrqZ9t/
+ODh5aK24p7/HiJLCGLN32dI1tYCPvLn2MOGt8mYI0fxvIbnJqdND7Ik8a8O3M6WAIobVghbaUvf
OQ3Wsg//VMhyTF20yDNh0+nmfdaI0MdDDqgivr3NSF7fEalCZMXwM3M0P1+a+9fvdLcdC6reUTec
G/Oae+pA+GkUSZj5rnrFtHP+RCJCYyIDUVQyUyDR/sGID8mbNUAsr1fprzM49XRI/E71so7ekkA9
eibSIESQ/1Y35ZhfHb8emUUlKPtWVH2onUYKcid9SOsyrFwvUzSgfUH9VLyOzljTTt28eVTANt1l
hSQSOJd3I9bwIKXXDOU16MnP8y9zGo58amB4ORef/u3Be83E7mQNfSUnpvVDmr3CEiX9U26FNVlS
UGtrHtqWCPnndkEGWy3OOTee74/AnpeDwLTIDMogt2N3mjh/eyphciLwHCzXtmR7uMKqShms0iaU
YjMWOeYwN4+plUuD6OQL41UYe5PUM9pjS9IjvlAEXqaAFJG94rz5Zswh4B4E9TqobhfQpf1l3x4+
aFZ96hcllAF+aRZz7FVrCPTrG6elbZoUOl2y7DNTOrVODLbk3G0wt92/oFEblR4ISNbUZeCa1aYh
SdrCHjMuO46xcpUX0D1X8G2ZtqmeLfbziRTdVBMWcLtYCEuZTmcOstwIBAcZEY6oxXIOL+LsdpDx
0BB4HqOpNLYtBQ5oNIieh1UKmKEEIzNb76H51lPsC8GX9Uy4PFyDE24dRSGtBPfBVkBFK5S8WmN5
CaKD8smV82jLsA295pjMNBxpHHKV5IDlaUt14w+sZSWAYS/3hU6Mjj4PqSo28TwLQM4MEgFpYlX8
dXxbpKblXZ5tIDUGoJu7538qXNQDyTDDzvK0lSOLja+lQ+YMoi7wOImcmRD5C9D6oqggAQDItvCH
T9GgIr1/DZaBV0Ew//8/LDLgiMRZehB28n9YKc6lwEonAuC5SBCNNSfmTyI9TBwyIUQ2vXkBmYrz
VokVDwAYCjlr4WcDE4Xqr9eoQxtELRpP7+208TNFB+WGYvn5I5Dp0qYJU7qTBKjeug3UzhDgk9Y3
A+JbHWYSN1Xp9BrcrwuhXsTtlQF3yHSrXHtY9jsFrVV2ih87JoUiIa4j/wqq9Khx3AWOEygUxhhS
V/Vw0UL4HV5GgSw47snMZZIgn2NfZmzAoZTCGb6C5QJBN0FaLW88S7gV3NoNlBEomD4Zc9/eI8Gq
k+wsjfhFmd/PPzTgZVZ/pxWndE6mAvMVi/JrdOukrrJTkF0dVyXi3wMUihrqs6ktVeq74PbOLw6X
WLJGU+DX9xC0afDakIFtp96r/D9+YWhEJRGFV4AziG7Bdi5hG7knz6+msqqr8LfhsctyarqO6Pap
Wrpis2R2xuk1j6iB/cGKpPu8bC99sH+DsT6L8FE45HVlSVSbS3AuSF8sM9SCWAnjOvdZT3r17Al6
Xwr+Pk3QpXBQm8ln6F34845HW2lwWM/QPoYR0OErCI+v4vxMJif/9w4BFUbjo/R8DsLmltdNzfL1
ZIZbl423pb274DcNVOuDRwhTZpN6x/FlvBujvcRb0Jvtapge8/A65AzM5yy22u+DrgN5uVvb5xOu
5SGAxuoKg8D2Wad/9ncv7GvY4Q6RncHRWHUa8LWlT9GyxIfsmWwCusDO+Ee0oykt7O33bk88hLD/
jERAy2j9hhqdDUH9VjZWfh8kkXQmoIcfrf5QkeWtomOn4hiQPTNEMmRDDRjnSM3lrUsvdf6oPrAV
vU6CFVVFokjOC42Vm/Ybr2YAzcoezcfb8eUQD8ygg/oAy4Wiw4rYR63INejwHqKMj1DLaaxiJzFE
gQAGNqq3wndTnHR1BeiH/TNTsXdt2Z4SlM/NpEGvyQ3rkaLUiZrAoa9VER7wkO+BE4FBPow1q2eo
5LAm9sTO7gzH0ZQA7VRPDmasHW9iamMhTCYsdQLmrSdAiBn55xLnldzHlkSLQTS/0YZzX3FTxutX
Fj/rYPlBu841d5IRPBJVxYYeO1AGvzsYKex5VYEGOWn0PE/7z0DP9cSghvBS5jtRSaXFn7bSOINy
RbV/7bV0X289jUv7vvKg2bcoLNuZAc7sw6srZ2uOACJgr4m8KbNMfFNbtOBuSiHxKSxTLt6U20rK
D1W3VvVLg7M9sUSUjkZL9J6SKyUeWrTNnYxAarzqFUOgGLZQY9yENzAFu259WHD1a/or36Kut535
zOczih/cI2VA5RYDWm93XIi7WaBz9rwaGvw6uJItp/djVpDs2+AIBvtKMuyir3s3jhtZdXYZi2T7
wpqzroYxT724o5Ee+6w3dU4f48153BAJMKyopB5JB6U3OSUAOOfAFbWmzwoBbz6BH7dBIk1b9qg2
hscBe6MAItDq0HFE77Dwvmi8mYEAU9dmxj8DJc0GuOLdtzFoYqWFgXJZX2B4o9JitA1LO3DPTdPW
Op6tGLgox4QZQpc895qT/3cbvy2nQkt3KgA9Pv5d0NgOSimJBqRdZmFEXuxvFXSeXsyu5dnM8swQ
6muTSVARt9pYtVDccFfz2WwgskBDHdYvOXirV60PSM0OP+/QVz5q9XGoI6e5BCKcIYMogyqvYmRV
30b37vUzADXN0V67jPSYomHvkVqoRHpyT+eQdfTxjOCLQwsmpdtUoVs64ML/QQLlNYQr2Mj232Jr
9ukYQgGsbdNcD0ZLvVkB3P3wSUOkoprj/HM4BEeOKKbH9EQUPRM6doUOUrGYWrK1cwK4NW4hVgXO
AE/ilSmPbheb0e5HnjFuduudw7Itoc5OVTHPUvHZne72Wh1vUk1EiVplpPiEJO3j2WTC5icuqKHJ
EJKcjV94HDF3VN5Q7IEa/TRZwIIiQyhNIa79DQU4SN2+5ZXiLw/fHWok9hmgGJmDVQ4pCynYqJcq
AaHkyMy+hg9suDYiv591qYsM8fT4ZgfvMUxJJkrljhwtYVulbVRguxg4JOkm986Im9Okp3HmeQB2
iZEAGwtrhRq+7lU1hMr8Bx2HOfzxSXuqmu6pkUJ+1yv522UqcnMYod4/zdH8r5LSgnzlUDHBmNPm
S5du3jpSXrtIASWqa84JvkD6fNqg7geDOtpitlofznzABTkgmsBgfi32aAee5dDsR9NtTng29ACj
6G4qgbAS9CWjg1YR/etAVxz4S1XhR3nwI5q+4qt08Th42TNDEw00d4pn3K2kM5OcYIyGSk+QP1s4
/xsYYHjlFdlDpkbJSOsS4ha3QGkAIsaJcNi7SD6d36vdx7qqQvkHwei3HvxiK7Qq0oterijKfpg/
1VDK7/ICl5dQizT0Qpc3regDB3QQTe6u46VA15SUrSoccJ04rxcGfF7PIShmySXqGuGOEDZ54vxJ
y4JRqBrk0Mc7ZT2Naj/Q7bJngUyq0Dnje2W8R66fvnac48fCbtL3rZtiP/kelmgtxu3JcMjGVgPf
z+mESTcXvCM/0IXaETvLFppMzCdFyb5UWjshc4o49OmAPy+Hcus7xwhWSkiGGgsY3xlE+XQd2xw4
v7VIR9Q/c0/ZH1/RLbX9IqbCzmdxOdS7S9XanlvZZMA1GaXpYkvDUfnQgSs4aMsLgDAsOJ9cnaon
udj8//MZoKK2A9Se8yqAo8slomO290G161ClZFqUunJvfRg0zbUkaGRy7dS/l6V+IJLIy/YW5LE1
N9sA9ZQS2BljEzhxxGq4jsz0/QecI+MB5MzKSOaUNcn+mYiSNkyt/c6voLVSd4HSchm/131wl+uz
TTvVAbamnEwC47cq5bXVbSBXeJfVOg+jcS1+zdqyGHEH7GEvcW320LV0L0ene1WrntcLIWEP/pQb
36huxelz58hqpY7rmFt98KTij234A3ov4RJL87xXxDhRhdQq7bTHWpqfNOCagF/AdfZmK4VoA5Vc
kDbND1Ns+smbzex7B05uBDORtVIsX/FoJ1RmT7ti88ZMtapxsmOAxHSvjjrUxgCLbhhwRudIVjnm
DRYk8gCM8ruT7wYU2ECLyG+tLFssQ3idAb9bYFpEMmBr/fluSOgbg6rHJFFqOPMusjIsit7AgHM9
JBViVxVUafQw28Vwv6cDes24DpbWT0IxMIOwXCCUvTnzZLc/pZ8YjIEotHtC9NELHJEYxd1mZ4f8
2Tas/tzfQ1cLJGkSyZosNeVtXULeWxPpEyWSJAmxD+ddBl7ki+4Srh9ts6yL1T5wvJCBY7Ya/3jN
MxDeLp5FR/K+M5e0BbO2F2SWCaQheZ2oOBtjlucSzppcHOXuAHx4fInUi+mfVo8d4xAmrh2VZxxu
Sa29OUEpvXcWBQh4id82SjAeapCbc6L+K3gLt/Dxg2Qf07efzw8R0rvyyVZwwLdt2jfY6BZEbPQK
8yVAaxx6iStQlmNEMMeYOhiFxLfse9vf19FgmdIDhj+BKQ6//F0as+T7fKrW+jcruagrXnHkCpYl
ocvdWIrh5jPdWO/NRYo0dAlGzj6tp3ULX0fcw9FJmoj7FrUz1f6jXEyMMMlwKIdri06sA2we0VO5
OxncZmDJ1hXPJCk8RXNzenEqC76+MBS4U5xAXFXkUwUy+pYw1BHQ2J4tRo1ZN5QU7DzYGK4MTQl6
4C7+neJEkwgtc6J5cu73QlRSzPgHEgauvlSeAa65LL93NDo/ru+N8p6dVBHRhGeuyx0878rwIT1U
TUIe+WJstYVtacowYPwCWgQDZQcy9Klg93ByMqgcu45h6GYsy4QdMkKqJsev7lykTnPQaLNo4Z22
Hg==
`protect end_protected
