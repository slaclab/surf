`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
J/2CPEUwld8+lsVZLfA+qextSaLLmdhxiMM55IX72kFvJTNco1vGIpgzw2fUQpwR+bogOz10ysjD
mlWpB4q30w==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
hAQzEmYX9j6Ng+2sJ9WMp2/GTEcdPGQ7ZhGD5PiXNzv130JHl4Fs8QV9Nfsp24XJdJuTaT/Sg21t
p8Tb0u1SKqt0x++DuVIGxyRBuIXpwvs86v5f1swVzbrS72iyqSyW2Y/a4Tqiismk3kf+qvtV2C60
8+uCXI4NPLZLL5esQFE=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aYvUzBCGuiD/JXFbI8KAbBaJtraSIxziVUtvclIlHZqMaJ9kbt1d/V3BLj/aBaCnM1RWXeiGQmL2
ZH3th6fEGFjayXbTm0YPPJXzcoAvPz36JUh9EIHUqryO2Ejo1rU8kxzVH58hj8Nrs7N+PL/lDUV/
kTCvZkVtD3Oy2X45Dwk=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J4B4PB6u909DdPOwVDcvDqhDfqlT1k+7deo6NmaZ2L61dOvt2LHULjgvfytFWo4GL4/Ie0nLKHwy
hfE/k/WCiq34PF7G9BtyqOamDgw6ZnPqI+PVzgS4RnskCX27sIbWOgCh6xv8qcBd8HKRcOMW5F4B
PK6cPsINX5/CzJ32+DFby3jsmFH36ouXeuv1NxnMz8Q9T28kLebB4RN/h9wK6EhMAStN2v4ifbOw
AHbb+t4YR0jl7v9MruX3elAXVjyr2SDVoIUWDrpXNI0RJBwsGlaN9EoT1M9/E3RoUsb9EYiEbp4/
YOq2NmONTH+EQe18ckJoe0VIDYbNX45S5PMoMw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
IKcEDAAtO/fqeeG2ndb+GWV6OxmwWmqle61ZdF+QgyBSHTQtl3LZcoBnRUayFhKSARCNUyUUdi70
pkm0EuRlKBAXiJygieOLL6OMmqQvexz8o4exuXC9J1LzoERE8yQM4vSlnikMLVJ5ojJAqIVPQDA/
PV350XXGl+9bhPIVlz/rW3BuQGnyJLw1B5mRFjYn6QkXND92/hKDJRR4cg6hQqAIATTEjj/OaWQK
nBsNp/tDuPfniiE2Oh9SIBJ8WfqnqIfVESLn2+WEJOlvBUmOgktza3bjrQ9wuWBeUKmwQ2H6VuIm
P+3uEaYyyWjlqHvwcmA48qbPnGhZTMd7o35izQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
sMFy15GYUP/Gn+pgxN3QG2LGVACENfPyezu3kS9nskaiwAnpBRUfUt53SMGX0nQjHkHH375zmtZC
v8sq29iXuyQHAuZLDdvkpdfaPSY/QhRP8frUntmUosQxcQg9XdpkBqqa0er93h4QvgM1K2nGN906
sT05b4ANr5jzLyT4J5tfeZRy/Q6AkYsLOvQgMyB+cIcU+dEkbpJaRcWZrAQ07R0L5tcpe01WyXWn
QxqJgYrh8KFzwouKIZ2gug/3cZ2LTE/TyXSHSkDmrfyY5Wn8f1pRo24qvxy1zTmyozKhl6IwEC/c
veVaSztPsssuu9JOMfdcEORCektTOSO9oYaBlA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 151824)
`pragma protect data_block
VCcSu6a/a696r9Haucx1tTWhaG+SY5/2FewUaTjlQ8AH3cGQSaah3T3pi0UXyKGK+gR7cYYT+xY2
HyHEQHrn/M68+9knI9E+M8ndbI1UZhRbwvgON3ZaejgLV6o2cVXp0C4ZdhQ2YivgvtIiot8Dc57n
sxaINu+2z8ofZwKwsA07Pbg6gNyUqdomcozam3t92OYQ0Z34IAJeP/HcY1VBNRNeukwQl32vXFUu
eRzhvwZQUOQEoE3aU48WcLh4DMJ4c1uhqTJphiP+6iuE7ornaxLC0cPtQyRUx+yVDCufa01+/W72
4dDlyz/hoLU4Ey53T+WDcVCmrEkcwxiT5rD2jA5R/VPI8WVLsqD2B7280Um0boz1ghKEBgEuUY5t
bBBMzrdaJTUazyOk1pnJNGpuiQeNkNBF0XxIhTlBzMg8fjn7cLBy3Ex0TfuegaC/vDmcN8MXQCHG
vR9AhssnJd2vnxwCtPV0GAjsTbrw0fVSM2l81wHuPf0laf/n4eHBu/UzctUo7sCEGhk6b+5/Vfzy
VxRvl6tqCAfMFLtiAy29z8mIG4Bu1LzDpxKvcg/c4HyQaOvBYpZyJbpJDMeArY63XXVA9NZyD7Zp
uwcIsApInfP9ATM799Kn2sv52IdempPSheP/zo6pgZsUbc9q4XHMUOgLcwkp/dVczWTRPLVxqgLV
KxVqRzgWgenyK7W5Dp3unU9ksmQ5DLsURkDcu00WDZ8Vgm4XH0RUZob0oLjZyhFuJOT7qEUK2YAB
TG4PQ1ls5sPlUYqsVGFOc+awHI63i2zcyoyUup8hX6RS0zeqieyd2boc8k9CjMGSRvHZVcKERIBY
iXIcqZkkKljV39cOcrDGtpCFbch3cEsRiIMIId47AiL2Ukm5iCMqjVzcZBCclK4A3RQVURto/85S
2s9kgww5dZSUmLlc7Jg4fuYzYff3UlFjyU9gAY6w/6Kkvczky2fBW4HNXA0D9tZGngrhe8ao6/G0
3sCVadNxKZQng/rlM4XShxswwhEQjbB/ew1dwnv8aqwKzHqa+UB/RY/e0q5XxZfYYXWVqPsew5i/
4l7VY8ObXvOUtFwScsXVb9iW38Y+eDx3h9fmFBBYhfToEULBdZYP9HkUDJ4FI/fWv6NsGUhL7IEr
JbVwdSr3DfBh79V73ytPRRdrvYyS2hiFV0LLjvTjOHdrXWascApdEQNUUY1OSi6k+jeji+Kj1iIM
4lQs6BybM8RvFdQMfYM5osbt9bEno9Jloo6/ataZE+lIJBob9MSL6SDAvRG/3lRxi6fGi85ilxAp
BsL3ATuni3zFoJCzovQbgmKbdM20dtORDFiQJP9CAChBm4oU5CD1vpMk7NDWJdmR+HKbjIm1EEvp
WoLK2k9uG8k4MLdyF8DXtRhFTrSxPURmsBaUTOES+Zy9kED4IvWNWg2XS4S73Kp8K77vXyFw9l0n
tt7dxmId5Sw+2QUyOuQKnbknaMrSqjF+dMU0fbc7F+e22xwlpengplVTcC59O+NR/nIeNuhHtKRH
ENEfemtLg96IwsUdAfV28sgdZ6RyL6tcuuepZo4ziE1vGaO6MwjyRd82EENqQ2ePRNsY96KD2dFb
XjCQBsbTQw3IwY9NL24UbvljYedvrDRPFzJ5KsKiXHSbjQvBcM0X4c5xZGt/JlYng8QsYSejB54e
Rei0A1eQvyIJN2W9nGCowXHmoI25p2viJO1IaHDSCqncwqKR8cwUcctjliZJ77asneasXDTGJIcN
j2pt0KtWcoor/NTIfzDx5PyHNkDYDTYaaFmEKcODFE4NnOiO65H/XFWaOuSPh1aN6Q/1/E40YJlG
couIGPXQj7XWUmmUaw/tjB+nUZfdLpJvY2gNmFNJrJZIGs71ouYVSTukDzpcs3bzAaKl+jQJALdQ
g3zBRctUonlz+VkguZer/prOsCd+4I5M/7VhaeBOynWZaPGvt0uV61RVc0GlBUkp8vl3xy3zqxMP
Uly2XC5JMUaNmYbX2chU2gq84PYSX0YSEu+jeo0//4Mn1tEgR7HcJjlvit4Ix3FgacBF0PYExyK1
9dshGQ7x2ZFW51uP2wS2grvTs5Idio5v3AdsFstZ2ItxgdmBGSah9rjTiv1YnYvrRHiuyiwylzQB
slreKy/NCdd1XTOj6ufV0hwXlanazz7ggje5igLIiWGZpm+I8WSB/QkbTPsZywH3AmWTUSgwx0xB
7ljKqYCzQp3cqpsK53TY9GLLrDgnUkopeM0gPQEOwJRTMGmO2VXnKYysKhBxHSYv83iOIONii0if
Xyx2HmuPpD9T1VoM0Zk6BgALvg7l7fykilU3hci6MqJOTthBgc8kqlTf+MbxVJhUFZ/7ZFUqSwtO
HjFGMLd0KxmGR6v5wIrkNT3k61i8mQhh035jyZtyRwX06mPnS9dT32gx3b4MMIXHilyVDfkh4WFZ
kfMEVzqPRbjPAmGKXBcolmK5aWQDxOhYga7ER5jzlLaNxHNVv8BbfRF83hbAdabEdbfkQABRumt+
fwEFMCg8N5SPqyv5G7sd73VkmF/YKf9BrFDg/8hj4JI0IGfOTPR2hVqz43AJNSCA3HZwvobuH98b
1NqZqHPV0gQ6yS1t20oGp2lh96FPLhWdGiwHC+zCsl95KU17deTkZXqs11y5sX21ICmtTDSNbNe5
CfMxrN8ljdxqPzWVU6MmRzqoiJ0VAOYIQFYdJ2eOLQjoX0ZUgQuuzD262E39UEfEnp3k130T6H+C
HNYSyn9plYfi5Tnx3Q2+lbTJxXXsOKaYmCrpcvX/qyJUs2ixSHvRUnvLhqvvzOXh8E87E5hZMMq6
wh+fGy1ZLoTUmaNtaMFjCf/COIFni3ERZtbZhFg20BI2XMUPdtB726R28n4a+a5RsD3FF3bmdU3P
0UDVqWTUgk3NR/pygdStifGbIm1ZsIPyLpPYwAVKd+Yw1uMglFgW/vTMI2JGsTseYnnZSXIx/5wu
2FZ3o/lyrmP0qiTnx7WrwX9YxEgWXXQtLKv+xNgCZf0nuyONmQFJ3arVplsard8Z5XDJtgXEKBYU
HukJJFYLFNaku46HAgTq/IJva7otCFW7cxcGPKT5Vuti2oXcftG/IqZDSOaxXc21vJN23jUJvRyB
DdoH5K9EQ0xA2CmGZfnvEx9NoqdoF7rIDYwwk9fCoWOgtN43w+7B58rWElcz5zoCh1hCn+fQbNfU
OnjDpAJ7YmnzLoY2k2o/gKL3O2YZKTXyH1L2aeZb9/LjShWM38Panm7IzMM6F/hScIkjSnrX2Ikz
5bgp0sOn0NYTsmSJ68EgSeCKxJ6tOE6HYg+00yrYptkV3TMoUYqiy5bd2b7WHQwv/g5FrVmo9SnF
7ZNqZpxJ9f23vfU2ciN8/vWgSnnvLk0+sjv/HwiDnoGTdZcn3vmsr/gstMMycS2+0IcO5p8y2sDN
pnE3/p2I70OehSt1vGqxcF2GGUTmibp2YMd+2AsEoZT+IDEBNJzUWMT+QPp85U+hPCOj5Eq3/lOT
HSAxQjmsZBYtd9C9Jgezm7SFZmUeGa9uQBnlrJk9K4rdj9d4KzQH85JpxRrK/9JGx2RO9IzJ85Zv
pHgOuUxncTh1UD+jYXGoB6Kdv7yBIuFt8oR7GX3jprgpegJ0xvM1uiL/7vnaaRwTc6jDkOs2NXBt
HQ1g1ihtfUBV13E/lUvOT6UPepW7gTTvbaSji3gCcVwOrh5k+pfbIMVKUGlncxuFRA2/seCmUNGY
UzTq1AaMVVmWkBH25UVTMfPrd1HzGpu9kIFn0GkEaDH+n2NBZa6Rbkqg/sD5eDSaLEcBr+hnbq/Q
Id5z2eLvyVdtF6SBDaKNxNqufcXfpexaeZyKx+/pu4BrPcxrB9nzDL5a41w/3w0zbIesvX7EFP+Z
pSZwkg8M+C8KBbtuGFmD5CF9jmlMTEVCKziFpLVhW3oH1XjSV4X2Gm3Z/xhUf6AzyauvVRWM6TLL
SHTaTRAoxeHIQ1pNf/VEe2cBt60b/HNoUc8Z8JPvBJ8TGImTS646JGPpKzAJ19KtG2liqtHuFlTA
aLPa+3lpFwEbj9RqoWAg+MHGO7eXYhipojLoyy0qAB3k/pRZyzoE+tMsNcrhqs+z7HkejZdrpk2Y
ayCjKmm3N993a8TxpLBl5YMdTxkooi/Hy8uEiducONE2aj0TmbAZJl7LBVCK6kALAMTIGvUG0mv4
xPY+vXrmroBV/NJb2tKDMklfhIR/qpDV+0znCet/WeO7xMnkMuzvPXRSB65CDYQ83l2pDp4rKqGv
WIcVu/CSTvX5G+DYI6wKQ3k4St7kkilaG11fjZG0tA0Vv6EgLGddOkrCNQoA6voRFgt+bDi1Qe8b
NErJ4RBVoI85QY5UscOcVhzu1jnC02Bsbjw/Gu2OslR2xovh0VJFEuONmoWwKbu5FnTVjsyB8hYM
oqB3lZ2R5vk2BFabEhWwOpEck7tAq1AYmf3YHafBr5DjiZKbXKG6jqhZa4gC6BYIOHaw3GOvpEI1
EbVYuomWFUlVOf4nY3Wv85Tho9XnO/OzxXiHwfF7hZyegOmgIsBgWuB6QpePaSIawvkX/NcPq4nh
z69qyRQyJJ8Co/vH860a/Iowr/GWIhB5/qINXRweGdHg+mgZlmkLIyTnV2UjwFsKW5ceOnLMBmtd
Xuanjh/qwye91YB04WyxGaOzZw9UqjSisxAtPp/vg1xnB6zpW36gMxnTZEK7pRdMzRVvwMD+2O50
cRjcL1lzzrkI9EEqfIeOrXNGJnmfqfHo4Q9rVTM782qoKP3piPvmAQiTtEKdLHjncFsyHV5sPfmn
aNzgGUyu40t3//Msjd3HZ/ss4gLdiWBVS0VOPXi1smOLGjd68eI+2qrGiFX9u4lrrHyV6qH5qbE/
sXn01o4j0sRCxu4L1nfCb9pK6LuMFrPnG8q5ye/rOpujxd34Y7Hod0lWpwt741hpGgyVf3VQuovp
MeqcpIrIXPNHIDsn7G43I0mFTZQJQlLGebQ+3vczRkdssumLN8Xy5/DoZO3eitbn+cvzVDfjTy/+
zUugjIlQbEUr2Rc6sVRdr5r820Xk9Y341ow9t3aoGYBc0V89fz58ACZc3mJjWxWFX/QHu49Am/+g
lBlFotPJ9C4l8aCJNi8UXTDmd01QFWOPVa+Ll3x72UIYyJ3IB3ae0xhKzfN7edEbrBgUZKT7ee88
LZNFHGfz9FaM8tfQj/usDY/d5ZwTuxPVY95t49eDvpW+imczcjY0nDgG5c3Op5gCZRoFnx2LmsXT
dYm6RaEE/9mKSXykp2FR7SeRwkM7sTFsx6+h3KXrk2l6xIxMHJe8UBc4JftTtYJ8BYNSEerqnIy6
+9pcGZg3ECDlqvJGzOJRFulJnTbHqPbEEA3nJlJqI3CxB4zG7J0jKgdeRn+EKoycpg5V6+r2e/6K
lLowp8wKTZx+TIGTfV2heTMuPMbkSYE/Xspz5AvS/I1jUzg7VFinFv++uoVYNCulOHDMrP5/puhr
a23olOwfp8CfCfxnby/vL3f1G9e3r5UYzhadj6PMyBwy6gKUI5bfr6f8eOZCosOkPOAUqpgpk+kp
Zt2dS1tFJRzKLoC0g0JaC6FmtMhXDj44HHfYoxp5si9zWnT/6Hb1K0EQj8gD9k7lMQ+jNdgj5Z2Q
TetG2VlsTq0vqosx21JQyw4pUU5afzqsjTg0pkVU7R346GoyxIuyFYbzjdEqFxDw1R+4mnt1wH71
OQIY00s8miQuZ5yqhxunwztcbYOVR99dHmfej/pFLG9OO6LDrkBJBgRjosXQdw+zrC10fOmHFwAS
84X9lCir6d5qbyyVvs0U+ILVm1+jsICczz9gpw5y8Mt4KoRWzQGI5rHv4xFhqW/0vLdSQ3iKOL5Q
dZaZc30V+quK6WR6Xig6d8p5KNKXotG6YFhFr3/OlR9bSOZyhCKCquFAj/LDPv1ZmIASmqZHVdp7
R6i9chbtFDILb6qua6AEFrC06oCqVXl6bngnet5GtPKCuvrp9dfTYwuAFbFUsvPvmAGnl5LXlplv
ex1FOWGKbFE/PJRhhy6n5ZNeO0jj9Stsi8T5WyC/9+/DGgf6aJHalVQudwcQyoLUBeaOt7NXeVLS
IbPZnWHdDeIE133nQtlpuZrXw5fijN8Ohznb/cSywpFzd/AZH4Zq/hHBIkAJmEtUA2wGMoYgmuiF
IoB4sP40XM0l3L0plFZE4gZM0v5eXoddacIQAu+ZdNY/KPfdrC5/M6GPGPpNSBa5lDQimzrJDqRJ
7O9IjWEosqckt3m99D/jrFmwqigE2jgTQ1oU16+873DE02B/7S9cIlgjPi1aE2VberphMzh0t0WO
7OBDOvmfOG03x6ZV6gDzan8FoCZKu/5EZuq3Gsqo7YHX+jYfg+br6Xu9jC/+u2kphJa0nTZR2/9S
HcBuaZJkgTo99AeFlcsCLHvHrkOaQfPcXhpoHUff7BEXKM81qBzMfCPi0gyeW6UsA07JPNoqMgz7
ZW61X4n852oi/d/9tmlWxJuYUTnNk2dAVI3SYNUQBmkdxVYWqCdgKTD6/rFueaLAO9UoXRUqsa52
DZUBASzr7kGlXJC//ext6rykiPFN7OV9AdUnvy9b4PtFSUMA7XAIL9St2PJKqxC9FFW6W5QA8xbb
ADwgHYy+dLjIlWEdxPEjfMJdiFUinzCsuR2lMXZSJmFmjVO9ZgURd6CD1MSHeJ0jD5JenEiO8f+R
jvjK9yh5lmgSYQoIhqwSI1nn5m/wA/NHz/TLn/PTfFiw5Xc6VyoOtE1Pz8n5QrdicO5OtGY11Tzv
uFGF9Hv1wopogYWPXor9U+Rfyn7o4+wsORo16hhYIGbPGa9pF/p9EjqIFFcdC22LY9xoGTjRpS1F
HTX93UPAG+kuNV0ieZIWpnxhAx1YrBmCQYYLsjtGxMYpMMMPFY4dvJdGBDHFGs/nwm4XIqqV5M6X
GS+8F+tP327QzeejDWdpUvsytp+O1GBw6qtGBiEgyE1KXDLSAZ+P2JJqPf5oEF8Zle1DOeEiT2Vp
Hnsz73ywGfQ/XKHa841py5xrdahTjLl9vKI/CmYoY4cEhij5P5B67VR6YLWcJWQciw4qej/Kmnoy
Uy3Rb1bYJOb+ty7WlYFQaCqKO0kka2ag74nHklcIaMEK95n/YN75O8gvq737IiqE9qe/cesM9hWw
u3MSqE4X3RfPl8kq4rQOouYPDi2owOV0nvpwucf0WR+UtpVLxhJHU/4dXmtTyngykFpSHqi5FuQr
TPk8dKWGpvTPpQ+aZKk4cfRnT+/H7MZ2QpManNHBcdffAvVNI6Y/J3URkg18VC1uAWa3fPf7PHuB
rsWbPske2Jb+pM/mworP+6Ghv22QKfeSqSn2nffXADxBP1iqgl6b67CVQMPURS054mjku4nk1CHG
i3EEUBVdMbc3M2y1jJu9n8ZDnQ/KVTNdQFRsWYeiXOyBIoXklNMLPQQSVZWJKcrLxSlF97BCoEsr
RXuuFpzLj/xOKE6K2afQEb5EiZiFJ44IYVfQXtQ14UGq82PWNOlC63wENlJ2AfuTBrO3Aa0KDuvY
K9bTTtgteIZ4lDdVytQaSJqHMSM4l5rG6fRXPfGOheAvV2tVddGbUSdtVWMsr2myAXcoLlRyM1on
5X+kYpqmxopqyjl1FvAReb2RMj/tuxSl9+OKUQP01b44nvFnYiwPyzsHXQXpaZebw7CzmHBGqpH+
O0rXrHy0pRdCOfcH4loLCPDw0vHjVftMH3IrmSQaUE6EK/80+HRvxZTfM0U9qC5gnB+uLDzMfEPj
9ejPhzmMfyYNnBOa5aka2RcgIiFa6RCvq8OzczN1md0aL6TQ7F+Is74po0e//P+Gf2ud5XBvInU9
Zje5CTFKw76JZ2A4t2Mc5OJwy9G86rftXFHFCaN45gTQOCxmkux6nV/NkKL7ccl6I0RnrqWszedx
bjgafvvd1pvR5ab28m0XdAPV25iOPzW23UPO2iMVoqgPdCIiKCWmg6Y4wu4ZbEUyZ7kZrZlTOgrn
bnAkb65E5XhuqvDTxzKRJtU9XYh9z0l+YKw0PSJHVQpOAhDTbq3u7voUyPwqx/qial8NkuoTDTzg
bh1p2MGihmolhjLzn6K9KDJPtepfSQaDHDi9+eDeVvz5BCTq4wsajedInSQ1zrMkZJZTpAMOJpLV
TuazdIfhe01FfhRejBg3Im7ktIKc2ZrV72UsmOLqc3wt2xqTK2PP/EkNygFCID+gr7BncZTBTLkL
xKHpznCsvw+AW5SOSqE+0/0/I1KY+vmq/RNf3DRDQhjwdDhDu8VKNiTRBkGWZALfxZsio6xBAKDN
F7lcHdnaDRRkxKz7oYqYF7C30jPWgkLp51B95foLKZg8FWi2sgnzneZE401qko6z7+fP/lTEixXi
5ar2QYiuTu3ff2l6Ugz5KV5HCn2bvspUh6G3gpWe4T70LxmTmqSokb4nlWog2YHbNZgHAYD4TBwP
fxKdyAo+aPln8OcM7dYlCh+nEkwWMk7U88B8x8wQIozxUe7qvwxDBjdY/gu5xHJO1Oy2lCCMM5ga
6J8MhdJkIRkuojgdcBuT/OSbsfYL3HbGP4KqjXREKJ3mqa5Yxm1t5Qv2kXaib0CSFQPTlXWJX4mN
79kagNDEh+BYYSjoHrKvBPngth12empjGleJcarPwXKZX8xalu6lsdzotHZ6Mqa3OPK4SSqRgGTL
cvhsXDoR8hDG9RQQkvhu2443u46NHKAMan1xk17GvtAIM9jJkt1m+KB3f2QBzI3m3lrqBvC7CvhO
6uxti49m5/hqf9fuEm0YNodmPtR9rvCxurtZvbbMd+fjr39UI8pKlfBmfBhvZfA4zGo6mVuRR+3c
BB5jDn28wHPcIUP3RHpjsRJ1ahAlpoDobEAxLsFmR+7975v5KtOR3lkVCuZhB/civXqcoi+d0d7W
/E1ttXxVi/ULPfLCv+HYq8vDXkpWXtrHuoNN70qGBykerxVoCYqWpuijmpohyHkf6eZ12tXGK87j
TCVd6sUiZWd0FFMbScN6e9wFNCdz2KMvVkAnSuwpJWnbk7ZbL1HsKxEngM9D6A9g/0tJRInQCNNg
aOZOX38/NdGBo8w2NP8L6cRBlDHgF3ZVg+QoUKNKwCuQK+XMA3hNyoEwBLqqaBLvGLprLnDlcojv
fTpypFNkS0cszkXA6Igx4gqq0VDBsMcrlJ9NJUTYfTlP9QsPzSDt9490+MONpzgFc1dqpjkSmY/p
SNqac7RKgYhHTPx6y1B8DGxwn/UFPiPfAe2wyXc/1BGkhoqQhkcA5xIOoNf6loeKgRtOf+SpVvwL
t7HgpO/0gVv8zcrtBTWbap3U1s4DMJ2TIi1CjPOS3ytvhTn6BJM+DTwe5zG1G5+SNJ8HTrg5Y7HG
ukBVnj9WZRP2boZnjJkBjwchrDbyVBsNGnWIewoZXhVOd+AzcHegjgZf1Qjv8o7x/8g/l3OAipAy
CM9IUls7nQ4+JRCc7gabvcP3XqyMMo0X+2OwdBI3hX2UfgUeXpisMtWB66BOQThgJKVdJM5XO5Dw
z7yDkQMv5XwOy0QZp+rqPIlg5fRORNr0VWZLZ45zWR0VOa+Uwh6sD/2eodIpR5rfsh7Wynsuqmql
B7onkVc8NkYmXkoG2W/1jGIH2JGnuHA5tRB09NaPw2hDQ1jwsYC0AiinwJDJcmoObb5kX3yjXr/v
OdZkYIRpFsef+9irGJUJ4ws9FvSb2YXKBPmJMn7x0pc1yP00RndnGT3tcj7NqD+Jmk0/+kZxvEUW
c85N0JenDlDX33MhuLuk1RGlfAtfHmOox/BMCJ5RW3yMtMPj2MgoJH5QlLVqUaOl1zgzFe/uxlB2
nwayOYKn6un+ZXKS0vME1UgvBho/4ZcCa/hpI9QwsfZJVJ6g+teGgAnL5+LYnXoTSoJWsLuIbh4V
dd/SQkadKo5aFTDyxnK+sIp+tt9/PHIojBVArHR4SAgp00Fj4JJfdPm+WD07wGiaRUnNDiB5sFyC
oIUhNX7ggnVQfqXQmQeUZWGQd3jpMD8AHtSpYUI+Vnb0Jp0MtvozGXCGj5SI6pPbO/4JPC4BLqaD
63jHedI4A4pW+TGB/FHgZDEDMMwQ0trB0qysuE5bcszhV7WoYuVMkEgst0kDkbQYW6aBdvoi3zQM
MBr3osQE/qXUpMSq0A18wtqLN1k1xXr1ql8/HvlMyy9I6a+X795UKOYoPW0BZBodltsac5C4BQaw
W3uAUAKqCmNu1dLyvo68eW3i2kqd5Ehcw0ZicyqENK7KfmXI1QfIWZcaLM2ZGm0lRZHAOVi+U5cP
X0WR1Ww5mo8GqZM3LFH39x6QHka2RUafX8fFOMA2bmS3fCc1Ns7Efj6gT/PiU7fYwb9a4rQ36Is4
9qb/lPvXZ47bs7oF+qow7hu2W1GbsdsvQxJf1FsZLpIDaxZ2lD/90H/Hunu6dvLlZ6RxygCKOfjB
7SdxfW4N04GyGUykUVrdc3XRtDV/4JI+5GTe8jPgr/1V0Do4IU3h3do81J4BNX7E3x0PBs0SyOD3
BeMgK832k/s/lwPnUHq2UHxwKg5YKcgcJx3ARoPh7JeEAxdguIoH+sHJq0mugCDL1iuNDiRmAmrc
dOFbJRnVGA57MFUR0UA3250izSOoIcV0Pz2v/o1zYGUGD8QPC7ZzkJle+66tlXL+i43xivPiSoPA
68hgTbki1bqlfGAYzS4sj3wI0ruLXc4DnCSjmC6Hgud6edEJtL9eczijJmszgE4FvBUqkPWo+hRf
8C4YoIMAMB8D79pc7EkPSgOLyBxTHzJ1SXzMvvVxlmNZQDSzo2gZ+s2BR3zRhIDQSe2OEN4Naupa
AiRxNvIikiAzxGn86XlbRcaWxyef1pyAmTMD5pWhztkZfohlLwekDAtWWcSFS3Rze//h/rzQrzLe
bniETcyIuLaWWzUSVpKYyx2T0fFGZF4nf04qptVemRPpQedu05F+MUpjESvpuYzctyHTbPb09Y3A
QDgAEsKG3wPRhWHHJWpYwzlNCCqobxfcp/pBxAQ3dlSQ9BxaO22YKT/AyoTPURGBxyB0wRD89Tfo
ZzD9pd53Z2Sjquzq7+PZcuBNvt4ccs2yAJxUBU9sswo+0S2RgazYy/7bAiAYHfyIVGR7DYq9azE8
BOlx1yZQDyVnMxIdR/FwiTqam+x9NzSAH1lw2GUG7AUuVwcgBbbK6VN/viW2Fv6dyk0rEd8/kUdu
iTf+BLeMhdFzip48ZjdtsXuIprbE41g/1ahVcoKWv6gHo9DJyDRFq9KzkDv+jM2aLuKZgCg58hMw
D6FTtMvoedzs7wDMzcEGIVN8qtsPBfn1ktvepU4j62yQ2eJqHpPBCoLRRbbanjl56hFfXd5UK1oX
mUpBcGscH3r6Fgxh+OA8SpCc7oL1KjRxPyNnyQLvb2i5O6quVnJ7kBl2ZMujqC4ePulYg5NA1paF
DHv78u/Meve2xyQVsDGspidYu3akyqTImm2q2J5XOl4d2UskXpuB9NupBU1MC6h2S28V7n2ffP8x
Oz/whl3pxBX2JuBtwVX89hAyhrt8UD/OqeISCk1jyUoSJO17qUsA6q3d75E/dgaP9OhnjEKKG9UJ
tCnm8hmi3OtzJ0tB7Rmo5/1U47FtdkzN60PVk37jz2Vj3kkoeVKahypUQoc5+3ChVW6X52MAXYLH
Kx1dzkFnrXMdmxTpY0sloAQCO+kf0hL1oX1YJTGqJklFZ/xers2AUyGBWut5Ih6iXz2wopKx/uo2
+2MiKLz55gUlY/mb/HlKDdZz2lZEFGxhyPZASZn9hL2XMwzoj9a6RowvE+fcOqw4/25o25GymMYJ
ktl50zyWk7YUKdv5JkFTnz/lKLLwbGP7T/HGvaQ1djFoMztSNrj6MsSUZHpqrRc8TxuwQqKYE/1q
+XWUHaBDME/VMVWLpbFbjsBkMMnDcupZE8K7rmDtReIq5Ghx9dlWSUTU3mMiHydOASQtvSW8zXvm
iUMXWKhorbd63jMwaLACTcnQlv0DtWaeRPOTuvwQvUPS1mFmTlYBred3dknNGYpbBtqt0XSjL76A
tddRH18qxbigWWD7Hqjcc+1pXB/pizerxQYt8xTdW+nBW6g+4V6nfcidVeYP2VzGU34SuuVeTwoC
PRwpyZ9+19/5E82H39cbS2BGr0wxZDitcOY1oUTBCtLihGvjADCIgU6499oTzNP2ZmDhv/f8wr5L
Hj8Et0YsAOo10WxR3Pbn3O2Texg+Dp7KMLdIX7WNqM5b2YHbjHO7HJ2FLl1Fw/WD0YlD8ua/dHod
3C39PkI3NmPWHz7b9QAmubmcsURNZdqitXRBlMn4Sg3Sin5wamo7zBzNh+WSJ/UjUjc+YRANtlfM
CkbATuptu8B5acA1lDiF/fX/gARdAg/H1b5mmwntRoNXrBvAeWwhGtFsqdjlJvdH8XoS1CdZVwy4
8RuMFjhtu/GTAQZZC3qy1KbPUtoPoYTi+ImADZ/xJ8XTx7quj0kIsRy36UiLXOXq9N4xdRVYpWwm
L3KkJYvRsepsYAfIL2h8hYnvMbu8oRwmGN/R0zCHcl5ZLZ6Zj+5F2nzf/6cBuSC5DUlusz+D8/cB
Xny2sFVSFGPywkHMrtgFpqguzl+4w4qTFR5IjgAEVsne8f8jToz+0N6k5jLj0f1pzEIrousO4BfH
qkz1+yfNgtEyFNUnAcUuCHHOFUtbs0ToTQWfND+BXaXUYo7oVqqbjj1IJ9bF93W/Rl5EaTTlWmZX
oEfOX9Amgz8Uifi+D3Lx6CcUIftGtx0lXxpAb656mSEeIrKSMUhKTHcjtIEi4+yYFs8VD/yZJb+s
CT0Qk0HI6zJhmEf+DOhpJEW7PSizif+AS+rKExsf6Mh7HTsbrnhV4K8txWaWf/wOtwq/zrQLMSh0
l+rxpV1PihXn8sBQSMOFH7/tbi0m8RB35nqNB9i5iIvhskmeiJGbCNrlEl3KCW904Wgn7m78YpyF
Bn33LkVWTz3yRUgyVJNAd9BLq0MKNKZsQ3GZ3GIO1XPRymPC5Emqa7c6X0RYN7pEzzmCFqaZW0Tq
7D7jZwlewMxlVEC+OnOb9hAZrL3s3CZGxoSUB6BpDekyPjtmGugyIEOCnS0VgFCyfcT/WhHuL/Y2
YYoF6LWhlf+NrCGgkJqtCGc4wfapUQ/gavObAD1BK5V1O6QS95Q+HgZE7B2DHJ6meQNdkQIH1EOE
oQsJYVpivaHkirPHys/Oce6qCei+qVdyJYxD6au/lAzrPRinMPJswo6U06dRGB65OxtBwJ/UPGvD
IiLtqOoNo9rE81x3TlKQxznwgF/D6yDzGaKOqVLqwm+Z4gvJr4g5HZni/hQnpwIojz18PeKZjbvM
OHyfVKI0/zc233/72JPepEjpysn/6S7NsvFVt2nlwrRUIeO7RdFVO0cCxvAY7qG66BsEqWlq5E8U
3rh7UoSA/bP1ixg2lfFaOFjs8yeqdcNnUS77nlXms4EwoCfUGzU1lIwPWOh4sixbBhbZeZ9bXhe7
AXWZrPZW6v3M1CuufYuYecxgbudoFm17MSj1LTGFth61avPXhRAXA0cefLHO6f/sW7BGmJvIvKFQ
QpnTOmDD0IAtt4pfAKHchLWbd+xJVnIFdyO9BzXfgmxyr3wpJBOUWTivShgYsZL73MrS36/dXxwH
RafgJo4Ja9eq/2sPLUM9goigDCO47w1iC82sxnuBdcNTBZBn9do+2bkOzfRfBD/Vlyhf1ZFpdUh+
1Tp8DB7lwAhgSqhDU6jHoPpxWgFERg4LR4rd/CtBwcTkIfHsHz/jDH9sV7UKO2jcfczR7XQQoB3e
Jt6LD+FO+9ZreSgb9G1Y87Kbj0Pep3GcRXWQuV2jaTZym+SJWtHem0GMRkcUkjr6Q7McrjM7LGbi
RcMiJwS1n4RdQ9WkA06ofFM6fGeblmyFUrCe58qa3sthkqQPkpkVtcGbD0WUVHw+781gLMUXw9Aw
eDzxkXjqPUKzGP0OKFVQlW7f9C3xe9+Fy3e/n3lBw7+8Xav8pPrUmqVzpty3WqPoZSqEcUObR62z
fXSZrjqkmm287e8LDxhIpfjmgFt8ZJ8M7XedNVgRyoU/3qVcU5qUWKTjN13BTzVCDkVoDmSYKI+n
ikRO/TyW/TTEvVt3mO7cpapWdtrngQ+lms/Mzgc4bnOCPwfRJSuEKo8yGAJysVQtx9PomYfijR3v
ja4WXqg9BAz9O8rvlv2PtST3TYZyon9xrNRy0PtFrj7pqSxx12W1ArmH4L2KHrZZjPZjQJ98FYzJ
4+foKlloOiSm8Kgx2PCGW6Xd93bOwmSCf0q5pxaTiqTQ09rEDmpYkM5CLx0VD3kf2kDxJtg5gowK
rqNN2n2M9NzUsU/FPfufCEHHCvFfbkhcHNBmW28whbSalYgJLUkYOBSoD722BIsr5ef465zXohLo
7M6nJghZcUfeSLSRjk600K6XL+M+zxmAKtx7+E8S78GHmhWfKV00tv6JDhbRZ6aYGjXQB+y/ytb2
sk3w/PNfZCxDBwR2nnWnTC0+rAw/TiRsMVrqPOAn8UaudHAZVKFdaSl3HaGV3a5JM93ywKOjiMyb
5OehRbNYHqMI+0cNEhZmO+O2OjAvGcXSQeudvbxJU9ID9qYkaJ77Maghmhjh0awFbRhe0xffn1Fo
ppH24V0WLlo+ICSkgMXK3N6i5RJPNeoQARsscpMud/v+TaPJWDnN81lc+w8cqL+O4YQrhXa4LUP0
63hUUOmkeCCHSODfwM/Uk+54IKkV0OeI9G+/6xkazGahxRftOBKrFaxqMrrw5aZenC+RZWVTvrko
gV8/CDY5AwXpR2BApE4MZ69ayAnzIAuif/SCPvBTr7DuUeVkwwKAKP6YqhT/1b0iclwiIehbzUDg
fo8IgkAFzIfQThFOMUOpLyySB92Tx5qiGn3DkTdc+XRKxelPbcDUFQTZzFoIo5VXr5AnwXKpf+Qh
kULEoKioSe/dFPA+FlQWb9oBo9BVbqrlkFujh39R1iFsqwl4CI2KHRZMXTc/W49N+3e4IRK1c+XJ
dc4JeeOc2igpWfesAj2UOASm6YI4o6K6PXGl5ZDo5BcLFK6Xj84kJDb/iNj4xOmlzqWiMuFNRkLk
GWlQnsqDEWUgf/5wThT0OuuFpU5OIeboCP6kCAKaRWwwFN3pzo9vuy6ZNKw0vjsQmbkPnXr0ir5J
b/L+MDsVWm52QlPd6LDb1/4lyJJ8US/ypHI8yyS4ScbtrKzUIDIWFhQj2FLbCf096ZKAeslsY4tc
Tb9QNIwrEtG+oU6iPKpd7U7oPHVA9euOwg2SzGyOHZqAeaKpZc7US7zVNfQeS7dQnTXv8eEY6S9A
/zP5rGiG0eV6uHPK8+7egyRsn/dAFhUCRT3ArQatROtDzT5lTe9UV+kOUmlsyE4slaDdgT20gvfi
qUsODYunqpZ6qxCag5jDvqiL+I8riPbULUtVRMYwpEBRn/YbhU21F5ltKdNxetOWkuajCl8A92kf
sarPKBmf45TeuG7Krz9PfVVLARXbFB3ZDsiptPTrJRKdyUmiiI+i/LdT99VBLR8iP+T3r6TUfqnr
SRiGtco5uWE6224COp7teBewYNNBfkDi9knNs45tG/rF/8K+THA+pz9seX+k5Moe3UwsR/P3oPvM
icnT2K9amYjiCtCC1/1IQazwBpv8XdOrxxqiEesc3qLpGCdy557O2HzH4/csCG8yGxhe3kTT9NAH
15vxH2JMK2I+onCh11xUwNZu4hJpoPZZU8YI342IDuQssC7lsRfjWyTq21jLqawt0ywB4qFYPNEw
kKPngOM2sz3Ga9xqSa6TkF1rHsLCa/9QP8mDpOQUAPjlCc9QtxPzga4JqO1LgTMwkEdY2ZZJYwQa
4FFVwrnSEe3ry7s5Tzpoje3OThGVH14rlf+KbtbSEbRuQvia5v2L7FAUbqlvEvs1aUQtZBldAH4L
VYnKOF/nuz8pUfABqLO85iv21vqjZaOxLDR7+dVm1xwsYjh65BT4eD9/dxRkQ+s1iQo4cYcDzLhY
4zIzG3OcVHQ0/xeKJLp7jMXRgYJ9K0xDF6c7m/FHCOAnimm5aG5Ew7bpkpHJCr2Vw/gs4ykuozsf
KY4QqudEbc0DvaordxQ6bT7WQPdorTcvOG26EA9C7XoRHspSDJkk49RbCe4jf0xViMMVlm9YLsoS
VAH2NJngQM+0ZoKP/4W2q+C/yYgk+3QciTF2/5ElhqgpyVcwoFhm1phBwtb0XsPve8hNFzUhtLB4
19N+pRmb0jmlQJNGp7mDx8SVNAhhoYyM0JS7GLInM0zDDP5FNdMWxSMsEvvneOdzVvaJVjxGrfhP
wuKmQE1PvAgmWcibHPTAKwdrod2+l9jDK9ufh7CooaToFbOT3Jp4A9/HDME4namIcoM3tJfjOD+P
spmVd9qzlGQ24ZF8nwUbCeDw+qT2w8rZ3e8xFMN9RkpDwJxQc6bdl3Iw61qzOglWHrV+h1MLYUw3
p8pn4bczNTw2rOVEZGGQylWQGHBslDR5ususnWS+ZJEEOnc0yaf46BSmmIb/XX34hlIWv4OtZCjV
ZflwyWfdu6zaMGohEwfBduxFnzsRvvmAC4bZYSXJ3r7aq9Ctztvaz81QDeTDVI3x4+1Z1OJw2ujB
iOcnzGekgcZiqEsXJrbOSpkB7AeQXpyJ0XKefIvhufZSaBOMVVy3ayr4X/JmL1wvzgZ9uqSZOpxa
D+SQbjGZrdJ96MPiRrEQ2RM5XZ/5+A2F4ISqpCdHeggjWaocHQ9ahQV7TqofCPG4jxxmEKB0daFZ
AfgYMpbZTniz2nHzuVHHxUr8c2mev6/JH+ZW0tpiopFJab6cGh/O0ZWVUOpACIeyHdZHg/HAHGJu
kC4aZxz6Hq7zayPiemZi8cCC5mb6FbxYkfeYeyLLGV0droa/RxjdGBU5tR5pXspidzKNJhAJkk6k
7vrooyahCQcSESS9So4huWAsASQkWkHRHVl9970KiZUvS3/qoXd7DlMl6WDwUnhYtmotQXNQQRbh
KKh2zeK9ITgOwDRK2qQbzUpwr3VFzzQ+4p/nTtfHEjTB8o+woE0MUTPI3L+9X1sPIlKsox2zK7Ih
K5pHZIwy2IeBkqeV/eWnv3S7d0Qpa9FPWMGiuTeS9E22/0JOgEa59SfFsRbdrmCTdRoMC24Q6NAP
HAjCsmfxINkkK9aFjZxMd0qEDncAYUE5UadedQhmm3lJ9jEaXsxXt/yevG6ZgIL19vEdZgWNlv++
8NqIKC8IdlZElGrXm1vudiaN3HXvbredyE9vNHFdSx970vrXLiC7IsPiczoJ3sITpcaYRBm4mSif
DTLC3lx/YVd/+BaLMOuuRDTNibZF0YRlhTjme249GJzCmKRq6kl8CzqCcXPMPM8RcnyjdwPMSWYy
7lBMVHAmzLBP0ssDrLpEbZRdmHSp4vqc1dSC8F/cFzJyM0JvwI+p4kcQnkCcSbHt3e/xElCsAREr
Nyl3YAnP7Ex6owg/LBiMX5fYWiAGGOi2eluOtuMvDUn9ASPqbRgIHrhtUnbVo1LAXn7scdQRX4k1
5cVgpPiTZemHQsOrFZJgI2zXQJUVUdzdmg69X2pRvEDEgm0ss0Pf7P/U5kAPYVNhzqrRt1QHGpkg
VVEGcvFllhVxeWbl1p0WysNBBqeeOQkGEdRaH13Pw8+xKRpm+4NbQin8zPMYmy2RGk8JilqN3r6A
cjePyyyTZYQf3QPnMvEl/eGLcC7mwYFSW2zyxqVW/Y4FacudfVuMqFtmkoQHXOLDS6aWIL/eA9LD
81iClMF+tbwZGaQ6ryRuPpaWV6YZIVfYgVtIbwhQ3rgGPU6lUarrFFWp9gidJM34F+swtY0Oz7nL
D/17nxwZi8HZqsUV5cmtpyi3bToTTVRU4t9GpAvQkAwgs/AX98Rvu4BtFD3Gos2plfE09TSTzrTO
wpRrzepAwPGHE+3/yRak9Awok1wWPWSRQkGJDyvLYttNnQ3/V8LZxP9cxMMFinlEtFVM3lsc7kp0
hyK+MMgx4OuWT2B9+biwoBNly36RpMqlIAfyK6ADNBje8ucByHBOS9gSsHK1m+ZQIqLh54ajzGlJ
j0ycGvQsA1Oo92r7U0k3KeiwETduuh4YOcZO8SOF1muQZyqzf6azuKRbao8WUR47F33VAalWH90v
CP6aj7wjML5jyaxM2gRW/S+AMHCS1HQTUV/WYeYfVyKwyWY1EGw4aH6Etuc/2UcOIaJVH5Y73IBx
F/8AulqsTPFbslFmHcYemnbvt3BEpHPNxSVy+4vRLORs+9BJOYjuCUs5nZQWBKklt20n/X/0m6Iw
/fF7htE1NCvkBCJfyuIA8ZC1OXAQjpJXowPvuiOEBi7afJD4wCQwtPANIFSWiRT8h3zREq+wawc0
JdTtUD+KrwyPiKkYj88s7U1Cu/Cf+KyIx4RK04Bp0zSS55tEUS6QJaGNFisN2sz58hYLNeixmwdx
K93MYeipFIP2E21RUTKMAsurT7trtW9z7Bd4ia9WSgt0hhuKH0G19K4fAurP+AD9tS6Ikg1mKzlN
ob9GwqlEHYQ5tVWx251fX8AQiYloIsZI1px8VHPkvRK+Kkx6/nScGGl4r0BvdvG79Qn0BSde/rwn
0oy0ujJTUDJ1kTZpkNyruGElyh/B9MTob/hE+HCrYp10vWQb83QKnv78YFjEA06xtdCoE5416K8J
2zeWE1VZ5Orm9IXNpSXlwGfQcOr0A4VaBMcTgNqInnY7Zu7hbuYVG0pq0lHlNVoIpFCSEksLZH7x
AlWCSuEHNogdlHKp6aZrD1moHxjGjTHJRQFp6asYnlPSzmOwvFB8nPmEmE9R95Fe3eB4bNp7GyrR
l+NwIPlyGqX9YgnEJDO67KG72OPbvnOkbE4Ef5bPmFIivyLnYXP9fBI2xQ5SnnohRPjXRf7N0Po/
XKfFD0cosqmQbmwpBHi8uWTXrxVEjlG3ZJNY5MxLpVCn/gZVkUuoPFO7TkdML08LZyLo+Aqi9pvR
dFjCjTvDryDC5bfCI8cx/qEdo0qPdlM3dQTdpYqoVKsTbmsnh4tUWq/ZNr8UOHLN7NcHVUpvs7If
3gNjaOK6vcwav4H/z32MmyEzg3k+93Q0UIfd88feI3FOEeGo38jbJbYE671fmfV+0vHY3Yq902kL
vKlDVv8nrF+sXrj93kod5k6lL/I/kRBxM8X34NgP2yevZAlTVi/1v5GNMRdd4wYn0jNNSP54mxrG
sOLoZJACN/3Ai6IGUYpiNafX/kRTcQG4A3H2OIFMRe1NqU/BesCWvLoNrVulwn9Ki9hQ0bhozbnZ
EOavvv9hEoo9pRFlPPyas5UklvlKIFn6+5oJ/HQX7tm+PD01+wwMalSDCWM1hmzo9GThf7w7cTDl
11lJB9UQ5c9DaCZZMoDU4HhalvvmudoIyBPsMjrWi+1gYyQFYpZUBdKixkY7pN1qps6d1pewhAQR
jtSrn38+/nafg4lsOoyYHSfMRqFZIl4hPloKBHU4yPrw5x59KLxMa53PXY67hd6uoIqi8+OVdoV2
UYIr49+Hb8cOYN4RGqL8+oBkbvagLUbroVK01aUxcm5ueK6cA25PHYdh+dH+y4lbREbdqA/WgD0E
sSa/WZSu5yGlCsRc46fzLotb3MwuVcyu8ru37tqr+wEa6UmHweifirKg3PgpSVscjx4C492OtEjv
CQJIfav0VOSj6uGLZwfMvWL3eISQVOnyoH+FXeQDqEvST//WQMw4KND24btXUd0JKAz8UpQb/wTU
qnctJfdfLv/MLwaalfvfIODPtLhtDN71uhLk3OwLWA+BfUQU5u+n/y+OtRH74HUhjG7AOPzMigjP
d4H8GHW9hUqbfwb+fhqiltZOmmasO9D0VXylBY7+0yDSxzeqTe+5FXTeBhoMhbDES7TfRabBm3da
K3Jhg3qeAuCeDG+rMMNFkD22SPF6Rojmoa47L4NrcRzroU0jDEAciyjcfpuGV+oYT9niqIg8wmRD
lRbo+cK5JejkOmY72jxR5okhjKbHeoONPb+oGKw4F6etaCg99zCcuMwK4lkPBs+4s6DYsKaRYd/V
np1IuPk+LUE9/XWq+8AHevegAPYaUIEY0thFP7WEIHE+Vv90vjbaUrwkn543RHxFeWIK3KQVm7Y0
bBmTygEviE85lfcEpThz5NEAO15KT+wcbFybP3d5ZhSYuv4SgMg0ENNVNc7Eq7USMYj8g4Il+upS
YW+oHyeuY/IJMlxgZTpgE4QZoUsCbPEDQu1DEWThaxyvyDFrLAGsz1t/qZJ+QGKjq94OkMGQHycF
YL7RqxIxrMkkndxXLOvy2psEYfiPf91gRWy8roZ1zrkPd9OtH6lr0iUnDtUNI9sHbExRM84UsAP4
H9wthIpg3wKPDqJWdZwp2ku1jEqq76rggU3RHUUhRflVL881/LYQr/1+KHSUl/DJqQV6hzOOKkiT
W+W1Ux10Ow1iwH0KxoxRDrG3N2OLhvdDFHWnwMHW1iBbn7Q/Ky6UKD79CXFx472hFkhbJ9+X3DUB
NLCLUZsRUB9uosQqeMmya/STfcthand2hK8pvokknVBfmiOXxLNzBIiVZ6RUkdceoB5bfbhAVZjB
nE4CGKBfAC68S2XuRpdLbgS8+3ZD6UM06dyTzZPNm1i19JaaPPzb6OC6ejXYSgQrb0v7WVT79kid
7dkSSsHIIU+twb4iA6M1Rq1+xVd/CqZQXiDbK5jIe/hB59+DWCSevKqyLQdMqiVH6tyUbo0E4hDM
Kzb0o3vW5X+R36+gGKnUc+ds9i3hVniQ3ucSqw84Gdx5HFliUNA0BzSE1DUmte30Qd0nT929Rv1j
PIKTUw6CjE9oj2+NJwN9FWqG3jfKcgMVK+1eTS+41ttnRTCJ57oRloIjMKm9zsK+bWbMAne2BzBN
Pcx6YsZAo30/jA1zwX5ueEpCC5dypVyChoGBJ9hX/Bgr1TxTOq+JbGNwMnNGq7wvYLI0+e6yH3Li
O1tnpkRWHiALpMiJZnBfVO8P4WYI3QMMjpFu2gWJkhmaKiY8tmNiaLULqBxEMm2j1eFxwxKgi9q/
WNFZZHT0Upn3dQcdXujOnwMnRNtl82CJOWuo4KxMEtXJU8O6iCcDlwVcghPmY7tg5+orf15cMwT8
+QuwNe4AYVGOuWrmmxUK8JC/yJOWGbjEEd+I+horq67sZeRhfFYSgaJKJMayn3inWFCvu+RINPhZ
MJN+UhyHaGKvjnR8tbU9vCvcQc1hzWwdF6XCMWrSHZWDgwhAAmGnvYDpTmVsZ4DRs88YJ0qTIq03
i0lTu2sl70e8MZaKB2n4YfLP84ViSeKGaGlv8uPJvRLp5J3qk1DHNehfYnnzf02XgR3/4wgSGnjg
xYhfVyE8977j5+PE6o3NDfbGDmwiTpYbgUj6rHPsqCTRdqDuBSg6d0ucIvts6hV7SWhP56ii7OJo
KDs1zrqTQLyQv82uziTYT2+ldF+tFZ68upS0NOFqBtV3Hg4K58P7njPHSfTGwH1YiUrMuxw4QTHi
VxJttwiwFnSbMpdCMBwyj7AsOcW3MzBDm5Cn3IMAO4u2VB1M4EaNsTtHbRsD5hLHe2ZrxveejJBV
I+AsnBGcRk2bdZvh1oqajuQGiv7HScmHBrm5w0BlqIYamz5GUK+OihpolaVScsI7BdN0pO4r2jgs
7qyLDUnRQpR/1seNBSK+b4wKuGFAgOWA4gvSJXA1Dh/vXqpid+a8epNz1sR1JjeAIcs4SEmDZ5BX
VFevQaXPsX8rMfsZF1eN6TwKNS2y6eKpOAahr/HjrprbtUQmTuSeYpa8XfuU84fQ+x2slot89xlH
Kf+eOrphA+eVSPBCLSCPiWp8RgVjUK5QUgbBry8Q9yV5M3Rbr/naU0wGlLs+E91XtdS7WIp5f2xa
4t+jO0nWw99Dixlm3Jdawgvj1r8d6BbspYCxZL0YjnMXUkI5P2XhjaP+DlrCYAdmURjNSA9k5wsr
ssh3pCpf5+fMAlNFTjaPgJzXEU9qLbPrIQkCeoVHj18rLJ4htbizJ0CRsVizH0ogDvS30sB0gP7R
oNQmEJwKre3sphw+2K1W8rfGh+C9DiDgM6fJjG60OGmHlzXA4/e3PMN6zfrzvm7gZBpIU0LMJAcM
IW2d5HWoNbnR8v8wCgB06GL9iv4nEJyBeUHeVpZ70gJ4RSCHyY12kDYvtkh4Af0i0aK197Ygaltp
Y274oxil39JpiUPOykdr7JDbiDunVvV8mDnI6O79FeXWY/Fc3F3rscimSCWXdENFylma4T+m/hwW
BpSplmg44eUr+8/7PRZbTUZMzDttyy5ypgbNu6dIyXKqjeuesNpIrBGLZzhyyRIxQ3pvY9Cie9JZ
3Gt8JrZh6wS5LXApVzZVQmmuE7PJSOof7NMP38O8/K8E5Zc0H0pVcWdn+45wRXc2esJOo91lTTOG
1qh7NhdFs9L7n8kjCT3AwRXOmW7CEXLRisa24Mccyyxj41t21/xsmFsS4KM5mUqPHxUQZodiH8qn
5gpivL49sXSFXN2qihkNmt/3JBToMUF8WyWJjkniEEbshNrJyr47sEuNzvrxYTLEcJevotT+AL2Q
waf8HSq2SOLv6+vEyQS0PtzA2VdcjlVgYYWRnbN+FOc+dL+146vAKO7hqT0pS1TIiOI31om0d+L2
tI5TkZCbpBFTL+hIqwAnsNyfQdXNbyzkvRenB/EpV3EY57rs7RTyc6gUeeK4FwOfrNoW3XP91Emg
vLt8MQrkk22eCT+PV10NGIab5d6aVXHGenwWko8Bn8/0E4M7wkOEvjYj6U9udR304x2Mmh3Z2Iyf
nw+PixquG2Y0uogkOsdFeHp0xPNXR2ES6FUH7bzXKuDTWa2G9NpA3VCkhAd1wMViQLbYYfS5zf+4
3vUGT0pHDRjyabdjBBDnP8ocpDTyrSNbSVQWnnJvWy+i/PDOopm8tENu9iRyj3TZ05kwpwdvS1jd
20CkQkpzzg9GahBw1u9rqxj4OTFMOAmPLV1v5Z5yWpcrtcoqLaejZlgfSgJcVoeJKWadmLJpRQ4W
VBwvYs9+5LtMLl0T3XV/jpi+9pym5VC00jMLYd/L8iK3H4QMs0bMQdJV3836g+2R41VZtaIPA8pw
c1FKSFL7BQLIdgC+J61Uu/SjJ8RL56yMSuD3G5z8DQC3kdILf0G6KY8BOf+i1v8ucLKCeXb/ByW8
4lkj8r3xDrkJwyOd4MNr95qLBlSZJR/a/eCFyEvO/iCLKAw30J3j+sNN83rIs8i1XJK5TjeHAW1Z
ZbaoUOkb3FkJwZB/BBeU4S90mf6ELzHy0k78CvkRdfBVPhJE+Vq538u1mJSZ58IFtObHAH9hk4aB
lU7UxkK7z0yZviz0FcxMHYWyLVmyN3z7QClV6KNnA3DIvFL1eEHXjD4V862aSbr7tvqBVDZegoTP
dQBX9z5CDiCEiRlw1s8OPRXK79UgDqTvA2dOX0ugQceXcw3MhurOYeciVXAh7M0ljjcQeU2YBGxL
on8zypYlMGuornt3IgNkKPTJcYfMTXy3aT/J34gHo7Cys44JU/fvuV2pj+/3UepX4SXjCIRsUexM
Hd/YH6uHKjr7k7dLkD0DtuK5/RqQQd+05DJd8RQDdlEIohPtklzkIsIBPQao39EFQYEa2fkS5FJ4
qnn/hk00p8U5f5V+IiSzi2ZH5pnREd1U+4W7cjfDqyhIkwuH/Sn+Qqbu5O2m/D51LnP0duznlGPh
2bEjHll0hFe4aOwJE4Gy3TL20jEVrJ1gc/tZ/mDp52VruOvpl2b5twR/jptQfHp1T4MHH62+OQER
5iTHpvAugmMMpYLwC5wdbFWh74NOvMMUrlIkudMirPVPV1NBOWiA9mWy32Q4kWNeGj0HxW+gyd7K
T/GuU4cPMascB8w2doC+Ha9oj576Q6JtzHruaUznXPcqVsrAZEKAxnmJG8mnpniWRFMkJCKhWfS3
HkjavgcXzGNSdyhQWY9slI2iYCnEeopBrcgkfObrxqfbdMfAYqa+SyoHdOZgHRptaJS9MKJ3l3Cs
9SuO87F4d25B5lMQS7vcamgaqdH3HgLDIfZ9I+95fBYHtfwBYZeO3IH5zPA6Hrt1KZ/Z1AgEYxOe
f/0eze/1s2hxyeikRSO7tsWIgfmEoMlEzDVxV62/z4ip/UOBWPt5b6FKOjgk8Y8611aM0BJT/Mo3
GF2zdJqVB6cTbenp14UcDAji2fGK84M3i6XBB6DQ98ZG2pZAsFgmfrwIZRKcBEUqNKdfLVUOAxCB
fjIzDR1SY6wqp8EBOv77FrDBmrEsgw3tN3SBO4zXJ4nVH3oco3Cy2RF4zr0WuKV/uLQI3uzhS1Q2
Elz30VnzcC3NLPzgRxrS45b2BSIJhAfKkMd6vBCdbkE9VwbOHOcgpEllhm5LXfMgAhvGQv+COox+
+Hy1ExQNEPLxcURnbd7gQboDkVW5wMwhYxZWxj+jntia4zBep9tN+p0b90sUeP46UnkCIRlYG2Qc
oGDEBAhQqkcZmxmYjtqwWxcqIca1XtWieFqzOcVrsRaJMzU2S4F8E6oi3X2qPGs3EiOsgcP7md+x
4TQ4hnmfqHyl/UfTY537n2T1qjr55j2XaQSRjTROEJK3wVSbPn12sKLc3fLdXTnqFzh+T3RYYgF5
np2UGpYWTWyKl1C1OU2a3g135tNPepRyjkeHO6tlF4au4LFgf4iid6atS+uDnEGmy6CpahVhPMZQ
wxMu+o1YVZSftKTmj2S6Wh6sIOsly3E2PHGN0xH0spuCrHbLJq/3PQCHzCaYqpL6buJwyvmQOlz5
sVpQkJ7K4OSmhytzRGq5jwo4tAPIWF+dVy4TAQukAbqs2vS2ihrczl/HIrNg99+GgxW27fIQmaCC
z017ePWdwKnfFNfnf84GrgCodRBT02f/ZKNNgLQrDo5XlWrKR3kCt3swGVLXw3EF6+8xtmmg/OrB
4Lv9KVtdkzGC2dMHOi+mlffgEi/KeN82ASfUPSMNLoqmtHx+1m/Auw/+Gk/7fpdnz4kfcQuyMBjl
jAtBG7F9ClQDv0LtpB7nCMFj7vnaT3aAf6R2aQjwB2NAaM9qimeHnskE3BK+aZzKyXhbSi1+yMvh
Rvj5cwOHs1nVLNMqvtjIAQigYMSKzU/ZXqg4AUj90K/TXfABjomXU3Bpbj0sm0EzJ2eKKPB4KD87
NXc/rjAd9nBJjZmnm++7kWxFDakGKBF/WfXRtt/6FrNxEg/UeKSxkQJ5E71AEOz0qT+pj0voyVGc
+WMQ14LeN8dsrlMQiLA0W8FNSVtn2oiCMP71mTg9Bi886g62sglkb9UTgrs8uQZySBGjaCLMAqS6
AkiKTy5DVhuL7sPwWHx3KgpR93u/dA/kv5ccbgWR7G9aslpOBfT+4RCnzgKER3QA9yoSgzJ/UYoK
Ym6CSxBmsExl3RETsTJU/WeiDRGUQ951VI0EW1+N2HzTSnJPFSTa+8vWEEJq/+VJdlGqYFpom4II
Llh+PwC5lWH26eYyrdA8mnTKWl82t3XT08xOxQJUUBa7z+uE+JKGRSWp86HLAD9AbdDBtwJ9Nisu
st/M/8ml3YjZU8JFt1w+cXWxapmtk5utUe314AGrsK/77uf/gkQFkOHvNf4dUG2pIE2NHp3nNbVJ
fN/EAbMFtJRnKUPMIMzTwrB+PW5fTk+HJJoaMlWnN+X2ZAL8mpyQ1BkBQ3NtOkhJejJyipAhQ3Dd
p03UYKO1DjyjEVlG1mGLop9u/y9b03rfdfY5gH52DUL4BAoGdpk3Q6fJvrQ0KRMtq0xSJRUoh6kN
o4t+BeVtDmEYCVL/qWEd0RJ2rctAODNNbFWYGsk5aKuW5nxx+P3bUhA8wzMqKnIXVSMtHl1W4yuk
SQu96Xr3CNYk6BYR1UUPx7Ytknu0OFnSdYgTwJ+1019qe2T9/bxX+BLQF1DYjl/AsYedx4VK7E8o
Ux1zAQNTT6QGbaWmKxCG5I6OjcdXsDa9ga09vJcxvtNspJgsXRPuz1kcCB9z5UHETUGaWC+voSbf
UM5xwOrvGwhdYft5y4aG6oieBH3JsMilQBN0ZHnSrbNkQQ0QXIG6AKIPs6mxEsN+Krw0UwQ/QEzH
iWPHwNp86IQtNPSA6Sg7LDMU/wGvo2HPJgjeq4+ObosOfylIq214pTu6G4gxE4jkNOEye/1VK/w0
ms/xA5dUkLJf8wF2kBvsto5DIpQAzYrgp8bKKFW8GexkO27CPWJZLsMkPZF64mAMVrjWR7ed3FrX
SHQ+bEWmeQ+0/MawTEKOBf97VaIwCNEpMaj37DzrsuLmoljuqAZhhiayQLg5cYqrE/LS4t20z0FS
lr+W5YQ4xUM17i6wSXZ3OmFrY7x4y6+Jhl6J3i3iQkqfLRtvCU+ji3+O5L81z3wMF0IDjzn63CMe
DbHsmSfdPATyY7KtlIK0IZF7kscyasIS3siWdDY7W/b9mZveWxK4SG5l8tt61YXjcSkUxOE13Xlt
mGEycYogAn6QjjCsPch9vuTI1SA2aONdmOt7FJ92SWWFtwNZ6RyKLKO4EDD/aqeqFYk2GfFUQakl
mMCn8+NK9IaNazmuS/f1tx6gYM3gaGyR1yQDyobcg1CgjRDMgEU6n4znijx3JBanldbt4+krIGIQ
BOAlqCVoOIpdNZme8WS2koCxgYO+V5wiQqI+duuvDdO28M5jqXhZSzU0tprhTa/6czrim1vAterr
MzitP20NexMQrjXO1wZi+D4wiEz3vckoSlnStpbBViRC3wH2ru0LRc62YCI6ofrnxFZYJP/14e+3
Z6AMga65lsStmYO4pOXv3XkhPxCPorL0SIP/xfyvK06bNuJupxJJ/DMrRr7ZwI0LANOe6Fd6Iu/J
IX07JdnSGIxNV6/uK0nuRVL1heKWgWYdfsbUnWxN2gwHKXC/DYFZyB+QmNVdkKUHhwCEjT/+MLJl
CHONGgAokwKxjKNM9TBEdn+OfNB+04HenzkDkU5S1J1l3QRAH1+cTGUd23Ll4U5eQ4UBYYjl9rrE
k5TR4EkX6DJfWJo3gwAwaMy1N2ZYIITBb4aZQcm8NUwQxA87wkpgotuxocN0aDHkc8nlKWG9WIbD
MPV33AWnohXevskb/tmE3TCn+35PB1rXnt70jq4f+fcJsexnhovQ72MDIaL0KG9Wk9bggFijlZ+n
ZyhPuEkgzGOdG3whFccq6L1ZLkvR2psTAtm2oR4jCar9qWC5hNCNgnXii5AmCNctXj6gy+Imd/Ek
7DNj4nXOwqkhzBs3poz6G3HUR0y+CrQV8VlWcFJSlLDpN5rF7ANx2igZd26ne4+/fp6OoUVhLoaH
l02bDGaucSxO1qICBS4WCB20M+v9ZGkcX/u7xzb5hingcA+aKspHB9jko1Fy1dtHwQFfTKvJu0pC
Ygw+TvMoa/8jtZrgkPnNdPupXOe1wnNuN0WBK5y50WtrWnLlKSkshtpXghqqyZqOrkL4ji+I4yUo
dA+tw5gwhb2OEF2bqyj7T0afLbXJ5ZzSv3xhlUPVEyBT8cjtGRkLg/jPtNzw6H+R8OB3df2IkLs2
8iRmnB3GoHE/8TlBq8KPm6mw3lu7gPyKQ3wkZ2qxVgjNlqjEf2b4yVXSb71mX4DyCBSpCMssZBEU
6she/QVCaza+SASVyPDNWSpl3uq+o11oDZDewVElWqh8Yd3rzt6FeJwfJWpbpHhQjivCihvdu4+n
mCeuMatXdd/UHosmCRuE5B3o7zXo5dug25l1teHrllfKmFCcYPtmxnOIMihuwoN1MJ/p802rgUoW
EQx435Lk50DsL1a3b7J38AMeuirduPXKp6Acfjkw2LSIw+OWoOFqqF4oDz1KjTYIQRiW7efBml3l
vkQOBEss43LhEbzzVPmIoj7iXxkCxR1CMg9DXfpqyF3f2nRReAERNRQIXqwgaLFnGahZoe/6Kycd
ayBqdWme3C+qC4vCjfJWinHJf9hoiDRxEp1ogoGzGYjvERH6eeBjlqXv4FarK4jKFxwabutmWCxE
WkcW61z5h4A4scWpqHYCkl7a+t7QDviF5NtUifcqWgMNXoHlJNnz9C1/u5oAHCRf/0HMIwLy7DaU
/zL1zNCenWdz0M9qqsuf4d4h2RXnYyyD/YPKJCuOYzNoGxEdrHya319XMZyyKZIyKv1LRGEujvNf
GawPkj28A8yKI4r7QXpQBTnkUzSt/KNkf1sdiBvm6SIcgebY8m/+rBcoIu8vzvKLGFH/GlvsH3Dc
5CESxKpf0dLD9CjfcKGDL9HYakU1i82aFMIvo/o4UFyXtNn6W4uEzrNOyGZw17QJ9mLLwE+Oiwi/
v7eZkAK5dHqhJpq83nTYzunY4ZNlbnYr2s5FxrbDYtz054vn6A3+xKzQuIwfm+2XGjbhPgvOzj8r
FOHDuoDfzVTXsFm/KeQXp24YyxOItS6Zvww5QVsRCW5vpVWbmrBo3Mh56IomutvQ3lFkxHMwAvmI
hDvnlpWVid8WyGNKSqCgqZFgnb0Cy0ozZTe8pJRlFxHAJgfcx6/9jECybyO/lWtHhCqskE563y7L
/64hMMZuHZIS6DOSUPSBNbXm2aBLNXQmDNk7Ev2NC2BMIE16hBG+mbPE4dVNay0c75sI24dE5pbC
yC0BCBxtuFYPSTta63OA98sQTsVnoC4RR6BU6jTsUD1KsqU7mhx2ZHVJTdknUrEfIPt05q3zuSRs
G/nhcRnOiJU0fzwfQdczNplKpLCAP26aNG3/gJy6bvrkTMEnYIJJF8HSyzrQk33mJc7XaXobf/mW
awC1BkKBQR6LWD90+AWiZU/a3S7vhkG+rHrtwRFeEPgXBYZTQUiymYvXkDNQj/na2EfOgNyhSATF
NSOTRtJHAxXjUwWGQodwedmVRtzomtfpKYkPfJC5nWZ52eN5nKd+U204H3P9MeKneKiPFEEQSLjs
YlIbxErRotMtInTQ7GEhfMv73IxQKIPO6NaXX8IFsBQOuxzfW/awN2qu/NsjITmylg6MA9fDwZDi
jyOmMsFdmCNJa2QRgocPg8PLxsyydHNrHWN9NeuuwfppAky+hgDcAvKd7YqdKV3VCLZMUC1h+UOp
qO/Sp/9Yc1MpOQNUmkMein5ehBZl5fGhjcPy35VtnLcnMTTRaoWfY+Wg4RYhtCCNwgvmxJSkz9oa
W4xi7wepsloUBl0ko5F8pwSKzhhcW5PGpy+tsQh7JJt41d/0MwbAB/MhhNYD4k2NOxlEWeVnog3T
NetKdN1A1/YOTNeGSNQ5/Yq7sDRI7tV+EoG9wOAG27GATKRNsIcf9AqwlO7/L6IUMDgBOAQadyqh
2PAxi5oPiVuRynWSCkQjioqYa8bT/K5uusZZpXtHzCtPHtoFRJ553WIkpIT3yBgc58MgkoDaQU8F
+IZ2+QLsBUpoyrXbjdzKYnEQRdpV40WnuVPprEnkeMHf4Lu/T4b3zYhz5Ue4ERgDfpc53qAipLz8
CsMtb2QM6pzI3U5p3sau0sSICm9ZF37ThfYrTVZLog+c+VOfjGI4AOQdxUyXXjrfBsdC6ts/2LHu
9sWw6fcpqLpB4qgg3/QIqddk3ZOVRbZ4ztYgaxuRX8hF8sKuYinoGCxNz/sNpdpSPR89ETAM6xWq
TXCV0T4tsYRqZYtY2Xm+vI6IDf5dy44JDs0CPILKf76Q221tnM9c2AXIbVMFuvDg64575Bu11K1c
eDk8ODZP476qk+CyFzxmTkeLxc+MgK1y4FDClHu2MokuECJqnI5Ow39tlZNPIWUVQDImHv5cwhzS
I2RmCrjxcmik4kdTp5ZEQqJLGV3h9H8NTSLj35HI1GwE0xejOFgr1CPFBgyXCAeeLCNrIBobiBuY
6v9yL/Zi9BQQh7fXZNH0DzHtCvqUZF+9u8fIQBjiOdC/kFO4B5xTcK2209c0CVzzTVe1QAQPk7ne
LPmk37sJwF3zdCCRKikYhVoHh2hTANtqW7SVDMZDx2xWGOv0dnFz0L4PygUdRacBrpPMvlI2i40N
ecPZzpGpduZLiL/jWGRw2YunNTNuejsBFuMraMhT1omD2NdpplnyI4z6bY9yaOqY0sYWaeisJvgQ
7Z4KZiLwIpDpnA6wya89iI887QJ4Z/j+G1Bi5mUPenw65d9EO7RX9X7fMx1HEgbZIBm9ggYvSgEL
x44vQCAXZu9KcZGeA5jbhcCmBpnp8u1yJBC83xWh1bZOIeCgx8hE4+6gBJqg/sWkO6OzwsxiB+yl
VuzU7774I9ptNOgfzXxExJp7tmnzhUb+oCUZO8JKHNPxAtqfu88KH8w2ZskeNa4MOwpiBc1rG5nQ
cJgXSwyNuVE/VlOM8gxLy0ahhAK81wgzFAjC7T2wKCbWF7ViqVJ+5R9w0zia4dYROrQ0edLo59wx
EVNLtoZLODRiE+UUujoCf7HNJrCz6DP/ZtOLeIbVfbvHJe3sUiKqGDLcl6djXjE531cOwZYQ/W5L
Eat2h2B+1t8BWp0Ym5vJeHns53P/s/n4yHjnvQB5Hs6zfiEY3qpq6zI15qXJ95UQSEjoPq1XA8G2
b2Ux9wOb0eeLkE6Au0pcrLS55TDzdQFpSj1Ko31ejuCJOq4Agi3aKaQGoHvsfCNFAxt/fPFZWSSi
w04isZKL7p8biGJ5hFouCtrTndGmn9Jml8KwEPI8MgJMP3HTLRhYD+6mmnmaBcyfH2z94fP9RUPh
Ga8XvbOCQ8f0N3VTR9V2P95uk91ljtKxBZctU2PlBBvRabTpxgGCQRj7i2KHJWurQLUSwPl8k03U
NgbGW4twZ6WV8L1WRDDXV105saPoD/8vV96ILyvPrsp+7mC7jIXvDtH7MkdcnxkSQ/uG4tuYTbTc
fRQ67IxU0NYxQz+QTwj4cteE6WLRnm8ryY5Ekq/yGWep75EWZfeA97/pR+n+cxM7InuvcOe/NLkg
uG77UJ+XfZ8B7XjmMm6i/BvVArPGGm/0j4Cum/C1SeKRlP/YqDQ0I84EbuxXDjraNBoBwfHCD3h+
aREI+sFNojx0vr36iqhIJ4eA5091O4Kzanj7FJLUW57RhXuSExPP645xAxOL748kIwQtT6QKoiIm
4TUZkya9n/ddounwP0GNGOUChARnP/W2AJIanW6xTxmLMyQR4TvcfL8vjOMl5C4YTv2uunwy6Ri8
3F5ljI0Um//EFMWnwBc2r/APqtKx6J/bNzePY48+IpeSbUxQbChrlCRIsJsR7KZuevYlxi/0Rj9a
wX+tZZN4ZBoMZ3C6Rp3L36xW1aIo91fhpHnxjtmGXPFex5NVARp6lxRuifEFRy0dWgu1lx5Tx32y
zcVezHsoym4UUEFO23LZzd4KhbefpJtfsp3JhdyW/UDh8eUnWwtft/S5Cim0dZ82QB4rHashrB5g
LjN9ptkkrXaoQy+HmXVvQyQv0V/r5VEMrE9+H+zpFR3l05aFK9vncHJ0e/DuUxqJ3I0Tn0ywYVNh
zKldW9UOcbC7AtWo/xnne/xelFUnv65KfxGnWgHRRtR3HttOJUQrymnZsA15s8L6JLBYnya3Nqb8
NnV5lAUC/Z63Myz+wopOrSdGnC0N1SmM2mV6V+NNOb2gIgR8lLga94cC40izdMOm/UTp8lwuvT2H
q7B3WCyRAZz53BpQW0aMNquWtg1XKVKd0kA1tYyuVomxBUaSUcKQe6+PDEt+bRZp2XyzBazqJIg4
iMBWES1qZqa3SXq69NvUWlDMsjqmpFQO8fb8FykcHA3sIuBPhJQOO2Jv0n/QXiWuSSmL2RTC5RwL
mIARGH31kItyGiA7U2JIWAIISdB69V47faeIpES5CoccNoB51XT/UCVaFThINXa70AnZPXqd/hGX
9dNtJy9qmfbiYCXagNG4GvQXT5onx920iHOurruIAQWR1lHpNtPZID/5gDM4/mT7dpCPicnuJ3pq
rRi71ilrP5cEC1m8Qydgeqjzl6Wgfixel90OxNqm4VLXDbk0Z0ePwvDZjuw7v8l+yCU5x92KEX47
7T4fbfbnhed0WrkJtajOOR1ej1UYw6etok0G025RhuHAlucIBPQTv8XqyyclMAA05r3m9ebUo3JD
8BQa9lrLelDIoAJVSdiDBx9JvzWZkcOix5VnKcpf7M95oXddYbI9mWoa+VwC+62MwEXq0mv5+s+m
msd3lxaUmJVEPi0k97KnwknsCiVfCLg42xttY1t0VeOMvHctcI2kbkmbVF0+0bW5vTN2Yz+tY9GU
g8PMFh3HGAyk37mc4rJps1it5k7sCb3QrWzx9FxoEBt8OLX/a4Mxi2yXozm4n2LSrh75K5cVRA+6
gqEu5Hw/Y1asHvFrgUv0uJ/fTzku8g2+qyIfV/fDLlNayvoT4fRNoWmiBTMiRxoJCfbnu6LHApqs
dkbbt4w3cuzyc9baCutf1QCX2GaTfbkVg64qP8VwQJiKEs9s3duNjOPpAh5mpwlCV8EDnV4Ymv6O
hKMq7jNNgkV+DaZ81jkkGI8ZjUPQ0GAfRpG30eKQaN48CX6nzaY43igrOX7v2lLcLIhOazibVJsc
VU2m23Kv589PrRhlsJy5p4VTeY/GEVmVomWS1y2uYehdfqSZE7RLZeo5qa5hp8fAUjvTxLz9W+4a
NZeYzwr3+PFBSGo8al/mnMGOG6Td+VNEiu4CIJsyRyFgfUpAJVwwY7qwdwZQ3FE3xgQoATo+tLiH
7aI5fOyF/e9C6t29mtuXp304Kt+CO8I7KMXEDShzzoBSgnxW3OUAwbf3iDU0AAFU7i/pQCVwZlZy
gX4mPZ5OmxPI31cgtOTXPq5L8KqDiumL3bAFDd1jJbs9Bhf7I5MytukDD8fhPO3h8LDsVs9Umm6S
cQklgJA+VhnqDR+OXJnYxxVcRAAEV6vjS03Wn+x22szXw1e5ycl/EMZmxovBO6Z6F9WBHdiNd97w
KvhOvcNSZV/Jb08Vd8AbmWYoHXv8zn/WlJrfbKvxYhdH6tFPClBPyxx8GJZqsvwDVAdc+lsxpu5e
JMPYucaIxmHN7h0MLpfRIF+nQVZ6ye4ATO0MVwQ15zZpkb/7Hn5t/2s7ldD9TkgwnAASGw/FBl95
/+E2nmeop4tb2V9VTaW1OmkRVbKjIRkH5mBo4tmo0Cp2+ENfdJF40cxR/AvIxq+o5uXm53YHiXIM
JDXQJ9UHEDF6+VOg47WMak1JHIKoxN7mOQ8l80DX8o4m7sTxe2azc3RrMxet/6gyPs1Zqz9US3W6
G0khfp5Kflxw8oW6TC2NalN5/3vOV1LaRO00o47GpVbi1q0HIPClBS+h+BFOXQCIHGvUSImde40f
Qzzi+wvJni4J5ppMU3uXBZj1byGaywd6cViqd8PZ/sRAYFT8VPF5LbOzJ91uyO2e8i06s4Pk7tVA
M2EHR1x2GlGNYouPcz2FLXftSl+ZGEhDbzQtlM8KvPkOZSKqrUO+oIg28KtKkOXThgus89KUEYCS
RAkH9kkujOYAY4RUTxxCHHXZMaSL3guFFN1sMFY34S/JAV+qNch9X/hfPqH6e9tRvAC6u95JVs0p
GtmgOKjAWB895E2Aaz0knV9st/999eRw8bY3i649qyVfIE3viyn4si2x1e0tqPhB/5g44Hnld5uv
6aTN1YW6ir5TMr2nxlJzl6+cilIU4Vm6p4pNrRlrIzKx3mbgK5govDsHIOhPTl1pRl2rmYq4jblR
AIBtRan/BgPMhzR/NayULC660KG6+U5osGTfyzNlqZj8zeOFrDwDpuAkcJ5c8P7eLb61tMX5fB7s
JyZDtPEq8A7EF8otHGJUA7IWP6wEhrbg0yJkad8cY8lleQMu8VqBFv+N1WvkShlv1wee3P9qZrB7
gQlpOpGhkdhrRiua2i1+r0jaRLoV1sgxWBJcm8VWZQGbIBq8uV4K988s/pPfa/rcxnObq6uicvvk
8PxK9TYgvHuNNf7Ov5ORVq29uMQ9e/2UKgZupKmPeUcnn1h68+nI1W1XudVUn68biBikeShwBxCq
NxLthRRJPt8r1uDkQkFYnk8kzRB8mGloqht/hQfVTdsvhnDE6WAdkSvYuplP7yTQAwcUktyCKene
iH1utknDoMF4pemdZkBMQhJfyyb0eHF10FwBEOL32yZXKuhoN+cAThCaBYOBjYxkpH1hYtGgUJva
1uolnN7BDhLlhPB6/AzLBZWyebu6HlGlXDGFd/eR551tyiJQfjJxhcFyRuGH9M83/PQrsCV9XCG/
HD/3pvv+pZRJ7erxlS73x6tzflvrBvyDYqFusOiE4T3n1HAdio1DyaYoZpoitD+MGNlS0cpfG/al
Q0lZsc/YJej3cVmE5mnvyrsJpSJBsGdwb+9VeqdTm/arzIew9ELbGP7rwex+SZnKRxyihS62pZH9
VCr/du1ceyn72FmzvqmgGfWWESM5bFrWQ4XmQIQkl/TfqSnxB/O91mtazsH3dhYgy5gvoDlu4W8P
sv3KnmFZeOtQsor5DDYyPgVm/4rl1nULjujLsxsjmguGinGGtH6sXguhX9c31wHxyD5w0OcKtln4
XoAeSBydzszNCPXs3ZpNugSAu+3XcutURwuLxV+ZiM1r8X2hucv0+e2dyLQUEDb3bOwPLkzMPHN7
dWXH7PK3tJawRT8nHOWpqnxkQCwpkTv563d2jB8asX2P4gqxX2yaRPHgqSLuOPrZqjQZjtp/Om5V
50j4xtgicgAoi9eWw9pLbXw2/uRdpbYK9eNHTURGWJiU9MNePoyl4QaEfbwAaWg5p31Igtr1uUWx
eEBel3FizVtpikajYXe2hck46WrzKAynOwXV5c6VH5K5OU/+avi7GjWwkjdQakNsgyaWKMkgvJ5C
moKzztvUs0PStoc2gZXg1lA0l/7UBQ1yGsMlOHWI/lV41V02adsfCHPJW3Z1tz49T+XeO3hksM+e
KzLe9me5yxrxPrkomZWFeDE7Wizvswlv8m0mlGt9LafjZYTgACAkFzyHT8Xzgs80fsz9XF+RusNh
eoO3QgfdyAo/oeFrOA79cEagDLgyTH4uhLfoB2G1ORh+BBvPAkWoZXfc167dA+EkQUT2t1jerqrq
qi1J5OnkJUNellVDjHaUD6tk4lkBjNqhfc0q3DMhdWp9u313kenmdowXgAiaUn7RoU4QAVSJsJ2I
a45dAf6LmLdrawkp218vSU+mMnNsb8K8hR/qh2gMiIppmetiMWkSBhaHCgJT6nbZwuNFtXfGWE3e
vkWaWd9/7HGeM1syPGgJ29hSl3oRu6lIRnd/DFwZZ35n1VZLCM6wZ2cqY1LhoKwW821Iuds+IT0z
gwW/UrLuaZfF79TksFs2NhUZ/K4jG/2nR+t49r/cD78jiPASE/Ir1M4+XpodWdvEeoObUOFTqxOc
8F1XFAQYLHZ2l+aMMQ9XsmRZfUbEP+UaXLYqvGMa9VOGXZw+dvrsc2vAyZuwZZzVfsO2t1rrJK2r
83FEhsZg6CZ7T7vjBC/Vbt5RPzgoDmNQ6+cbTAdk/fR7kdsRPe5OX7iGukyFSxYArVU+/LPUhUfP
T6NlYbH3gBFB9CcGeL9G6AIiDem/vLW4eMImLw2FW++vwf3vxw0nlYHjSlTEPyI25ErrknJo3GUN
nv1UQG0MLjtewRmzMLM9Gu9MQe5TWAFvTB8t/FAesQudFFs8xpM6JnRiIDBhPvUCKw4YVIGdTJ9i
9NlyPmuSNjkLTnbo2++cUzyebqXDbeziRO4dD6KXvWQfwFNOMODaw5pgmzsEaU7fTaCwcBmLj0Yz
dCkw6zG0dg7mfbK2jaPRUPGfmbT/pmbYmAMvh90T+PMQZsvYXkWa3p5cJ9UysfeHzoqdWVfmgJOM
GYllH3+wsLt8AEAcwZXPml16PdJ4fe20arba3bqvSbZlx9KcJNjlgF+7+LkjR4A3MbrnIpoV725e
f2anW8vCh2T4V9xRGY4+j8NrC79Chm3LnYo/hOiUUb8Io2p3MCQ2Q12n2dock6OD4Ncfl2R8dnMB
YfwMwVLBDjHb00oo2I/qwyM1JkOjzbc6b5zwHeZMhlOQkIqiAsz8+1T76gkpt0IMSCGq4jpD60Iq
PN2lsr/ZywvpvzytGo9rici4qDILQMjmfsi6XS0dZxXE33pTTHSJVHVdoqefkDn3RCW8cQ7KA5RN
F9eH63wx7HXKRkdyPeftrLCn1SSkB5eb37ThbM5dxStDrQSm0ji0yCES/2s3h4G0HsDZgmRWpKi2
x8Dx14PU8IO6KRWmDvjF4mAzilxr8Ymepup526VMFcu6Wkz7w5ccX7aS4FJzlvkKyVkTS+aYo76P
vYBOAHBSQW1UWqMPuiuiSQRpb7HO79hlNA7kxh+ZAWjMqkVGbTv7UKr2TRoqH7tvMl9DZG144jII
dYKCwWqPILMIAVTDhlHAbsne0mAhdiRwP0uUdf9lA1LuVxjyVIkEE6daFl0+OdoQg/ViNN2AdbCi
togDyNiNumdQpLZOxrnDUDmtym1b0heLHq2fsQwl3GdYi1EWvK9oGHZF7Gg5VsPWYWCC8XEmB4IH
p5UenNN4tB6EcTRYcp/J7AFxuBFFQ9q/tnmC16UYv8QFuLTo/V8XnxJsSQxbEGXqNyqiSkktL6Ld
ePHZT2EkkfW6PPDnXPtWTm3A9zrXIAP1dfO74yY0+zhSfw1bfJmnKIKWyJK8tZmt+C0xGa9WHV9l
RdnhqtZuKGMX+WtNgUVIBP3NyRFASS37YhimxSYkvHmDFyF/UZuj9r49k344B9FQuIFEPKAycXUR
FirlRs8AG5gNH2W/if7soRrF5bKkIkzCoQVKZhA12NZxrxsEkJ41OzLXm382hgmWmXxLLmbi4FPK
yTH/DXkW2hwnErbE0H/QLKhA2xN0pW9IwRGR8/ZS71UfKZBn9YMTyQWXh/1ktgSVu3saIBMKcjhs
o7akozrsWIatgFzPBaBO6Ajx8KAlQ09vdSLCqWZfg3TzRIux/L7g43PuZmcXAWybE2bCa5L6NOTC
9SvssOvfVMlofXg1UZ79aGfeAATSIC5dZiUKx2vK5tSYED+jZaDNeOSRoOFhqa6WM6ZGk042p2BH
8UYrOWQ3H2eIEPIU7FGzxBa6MTZihCodU6K7rrmPaTfD8BKFvpBo8iY+hnhxb3GDUE279P3Dbcj5
n09EJB9LiSeYJRBIGG8LybCPIzKrMY64bpq6G9OzUXeIteKoL7EGAsLB1490L3minPk13kBPKknf
A9H7JPw0gc49I/KhLT/aakKZNbp49rrGP338iXeze8qe486o75sGaK8IdsFFjSCJxpXJ/+ccMoWE
kNZszjctIpCnx2BqvkGNERWlfTo9aF2aKiOETwnx7Je+aRaDenzeXq066xCPiEgVR9dIiKnLmTVn
CkCrJ9sjWh0UipGJpDC4AvIPT8/qUwtNHYR6ujvUanEqaM5FGP6sIz2ALThP+iGPYdAexcSLsxuj
vMI3yNmePzxLQ8t2HMqK30ULRriULewB5P1LvawIAPNaXYbqNK4WXgFMtm6pxcwI1cDlmJh/2tDU
8M9eWqkgInXliFkEfk3mg+U+PSvcJRRoggQdD0ZoVC7rx1zQYDlKYV1UsocSd3H+FwSjNofNJc4d
2P7if0es+O37k+s5pey2qUDQW8zXko4+KS1YViiv0RgrylfG2ap3j+3TaRAHMzJQWVaLu+VC5sB8
cSoTieyPQYrl54ECPe4cjWtV03Q8tZfYE3VzwQZyL71fSE48LYxWIlTjH9UzGsx78nk/c7yGZgjR
f7yPDDspdvU3hEWm7Kks5/HQXacFtZ40MxPeqlGVVN7+8qQfyOBsbdx0QTKx3mtpQcydvklvmtf1
7Gn/adXpowzAiuKiWJCHoDi7Rfc80KaAVlYort3lH5Hjy3JLV3H0Y8YoyKBLDIuhBjC3I5/DtVg8
9UDE0fecw3qp5r+l4BOw1lh2Ie1nbRjmhrjHwY5jBwdrp9J6yX8ubh4WqNXsXN1iWInOAj7VAGKY
/nxWAdHNIxfKsBW1M15etjMSieTs1BsYtLorV7t12zbtEdeRwlMuVB15YW3H83HL3oZJasHOeTHe
B7vxkNKWe/M0Y6Z0+txz3NMg/Lota4uxSuCPXO7kytKWot8HU7QWTqV8jlJ+opVRY/v4qKFcq1TC
i0U7gS2K0PBw3w61p3n763JEsDZm2glpuMoA5KnT4NwmQ4Aw0lFuDMMkmOzozI1DiFws9MOZdlym
xrSmpiWUFMxw4mVi2cOtpZwYG7NnJPUZiNIk1jmv+Han1oFYA4AGPbNfJMWcfhKFdKt5zG1MIqSb
fbjHuEWX5YeOZ4ZGWr1fAeD/eYP0KSoWmbndk57RVJ314wUMum0t0vfkc7msozFgFPNu+eomoUhh
KddjVlxrVqJNjWGYTNCwqzerhaZNjXU5qC6Sr+yxwKtZ5lwbyxk6RvrDQRYlalLPJW9GaUvDVrzB
RYwqmWEry5FKszrjqYFMFSo6RwahkDidJ8sSTKIaqoelDfiRPLidd+robdFy9zIRyl7LolK+gmR+
xtRY+NbE94kvmqH3Vi7fJ8h1iC1QOU6HL8eOu84/AalOLNEe7WQUXU0S+KnBRJtId1QBcwVy8cJe
IF/judep3M0GpzY/qks8g4MpYWu54WA8Mf2NQddekJlsU8S8GKgWRRoZA18WvvidSw6wJ0o23IL6
xadgnbViQYJLBlcC+fnTVq2KiuySbrHrXZigGIfRqDGFz3Fa1iW64UNvaGq6s4pEytTMAeQZ0y6E
ZbnWnsCif9UBj5/Vi/KOrctmQ7M7eNwZa4YLsOn4l0fOQBFtoH+pmsFYmzSx1Yein/YD0Aqrv1u9
0tK8Mz7U/LiZlXw8oHsWPw4ODRiGRzBsQmjUvmpXz+mnRRNIBxSLga0Ns21Ev0uoSrY9X1l35zsJ
1t/K/Vhl/VaDpEjFINvsSynrxPBnv9PPkl+Wpx4PixwwX6GtO1ZN93CPIJjo7WY6iz90wexI373v
0OARfTYxRxXQd1h+Ds+7fpiGDZSlq/ugIrzYSqAON5bnfXzlbIpKCeo1n2FDmWy52Diwh+g/Kv5v
Phc5lTg+QTO3/vkdEuPisVupT38a9AZeHuKDDeV6ydLbQr44oRphY9Z0u6rCfTPikRwogNtur1dy
QY1+bPk8Wvfix1zQlcrmw+jluTcOEU0T+gA3o7D7xaxhx0J2eDoFYQj1Ageku1rv+r8wzoRHDeK4
/fWt+5UG+OM6NmRemAEuXAOn3gTW1jcHjNLNjzq1qu4OtkYPjlrNcXr++Gk0Vm1j7XAIpQ+ya9YJ
Bnh66YI8PBLiKqdDR7QEuQpyS9vx6FaMR256JI2hFswtBfg7IDXM6G6OnxfFtZgnBRvZB5HwN/DQ
htvWXydVnO/HQ3iHBYrn+n9ccYy2E2kX3yw6lqhy3189KAvb70/YOnAAsUH304oMq+sWUtX3Zgvv
yrotq/2g0YcRViB+nebM9y+V3zCL9VVg0XP5hxHJky7q7Iy84rgcP6qX+SrYc08pdpLCZQgCRfTd
QwrL83I9DrylzxCtyeNJs2zICkpd0p8mUb0OoQXFS6pp6HECasVh2lu/E0BBEhBbjSuhAUKf98xX
HKwrkeN85Q0LOd/dxA9owGreIZavPtaKiPjfKV3kOqsjFVyT2Yy/dTZMITZQak0c4P4aeg6u/38N
NAEqNAmKEdCiwbBXFL+0lxvBt6Oxv6lb6p8U9ITwsOK+2TkhWK9U6Knft4gloee8HErlwMCskaya
lNNwgbQtNbFTl2gIVaOU4FGMF9/5rK72ADJnhG7ybmfw30TfkSzKYzikH6EGe+B2Q7RCQ9G8Hxam
1+8DMXUXeG3qRbUAZkGAUw1usJSE+3c/m3op3Dt7zrt6DcV7X6qjHNrJpnYzj3PogVbtLjhbESNN
Vivc0Vfpc2pt0+p4Z1X9C9T5NS40EkHknV696Dyn0cih/VJYRs/SV/SnpFXsGhSOB9De+RpY3Bg+
C93ZMx0hkpE4czbEFuc8QbSMxU9KEPgRegdHk1d3A1EKWpb1M6IQRkyRjtg3A5uzcSErly2T9HYh
BDjlUSClQ97tFUZ6v64PEmDPLw9K27Ez7ke1wf23qvj7Wd5XFFxt9WufUraD2OiqRd8i96n7NJpB
Pt42AxocMZdAnWvwjBwCfl1QLG2RiRm+03+yCKS/vAGVlEzNjWwJH9SzylySjipAVwFiYtyjLUdV
R4PelF3ZZ0pfmwdG2pr44xoIb1knsc1L/EfODzXNwMUEXHaZRIuEmMB8paifz+7tHPN18VF5X4ka
sTJozM6ZYJTzKTWJ5PYTHzfNNIYknIqmjU8WAGb0R/eHOJ53cp1W01IPbywRnhIgYASDhDDVnop8
EAiI3aBcwZmtEu1bCxroPs0DH8G3N8mYYjcX1AWIHgB60KLybWTgfUhhulokiGPd2VdNZXh5r/fz
z05aJE3Sm/ZBx1HUFIHIotTtRd8YgpzZGpJAyJjwSIzv9p6YtEVYFtHADmaEvfwOtWkFKtwLzUNy
3TFGUUThasRTKsld93zPNQtNt4XxfJgEr6ClesrSulOdPiuyB4mTxzVsSZ2CSwNn5ZxNFDwvikMu
tL9OGdDNvzp0NoCCzme8IMOq8gTP6zN7o5j2s0uly1ctpDNbo5STm5eCDTCiXQx8I0kTNY7CZeRv
tfqBx4ct5rhxlpJjJe52lWRbwTX/sfgCR2We9egIYmfKe9SlsJ6BCVS621gp2OeKaZS8ZOHro+Lu
z+jcO/L0dYNNhS3ukQ8/aXe6UtQgnylWlvFOqkvjGc+D664g7FdgIhnp2hOM5mxTLTJtFOQ6t357
K80apaTqvKd7K4MiVbMaWarNXmXxVMHIqpok9N9M4/TCt0xF+SYIdJabJfkKRstIHKNVQazx8yEw
tnsZ62D4Qp47Rgl61Iyz82Rbi4QmdhBMcQm4a3pyJRi9wsT+HguioCq96J4ezE7THKc3F/bz7nhI
n/f7HitMeFhOD2nFxEpK84WSguk+aNFguX4of6oHGMr4QX2cbsr/sfovv6CKggnZcNWHrJYwYc2Q
JUVmaRwDHPwnuhAVuByd9RhWnINRz5jpaxrxFdKhYJyoRsLVR7NeyV++in/XcrCVeE1G5IGb10Yo
EPTBMO1OugO5Hegb6yhehmTu5nDId58Mg0VORIt3jyCBVAFUytzq4vjyj/inoHFPtwJ8Y/BHb74F
82+60Q8K0uoQe52jfmt76hciqpbJ3HmRXqJfBjlasY4UhhYkFsqlKQ4Ku/crjAudBSbKBXa0hcBp
arTXlDEL0xOhMyQ36DobpgllKvV8wElk7ps7KUjf707sOlGh50QQc4oBiLsUFPOSFzo2+fJ02FmB
z8UFOBUDOk4SDQao+1t36i7xvPbqQsNLG/EEn4iEchXl5TtE+PCDDC//K0Oq88G3B7VdgB3hDlTK
IfGAm0sMupUbk/q15xH7hqPKAAtMYkyuJhUmhVlU/FfZ6Igl7gQPBUj2kEgTllICtujooZAvTb8f
oyHV0idE+7pfQsX8PDrrZTT1xl+7o5BZv52TRwF/4MSaIqBm56pgW8WBYX2EpYh8eWy+NgDx5XVG
GQzhQvD0VpXSXPQ6DVWGTDVIzOmWpQZW+yAM/buMonf8Pd9n3U9kwWsCzeTRRa9fmfVN6HLdMmj5
n+KMGSHWBzKUdDROVBikRraLU6emXqRsebIsRdBh5WHgIbqqtr7E5Ilho2cb6OUksWupEFfaOCwb
y/3MUfp031IHTj4g2HppyDGUafOYNyrF4sdLB1m7HSjs4Bbwm8EYxLJi5UcmsPY6ycA9D1Cvn8eV
bi7jNhofrYqS80FITwsjF2qISXKqpbe2RVX/aKnlncPN4Nv4nEI62MabvehAqTUSsdrQbAHCNmVD
ITbASlS1lvJm/MbwVzJE8wFBZzQ8fDjyzVZhqzOBnH6GG4JUEhNDhCDQNkHjZ3BOX+5MI8MemRs0
n6Pw6ogNbYDHZi7BmLa8OjM2nBoRVVYRD50wJPd1Xk+WP2MUro18UhJwmtYHOLl41FS3ko2bBc46
UVnXU+pvogRbe/mS8N+q8k21DnJBJ/g8TNov08JEpwTg3DUutvuxGodQvph1jjJu9WLnBcM2FvOy
SHpVS036MFWGgB+e/Oji4F2oz9ZT0cTL/Z/W3I1gKevadiVHE9Xe3yQehqu5Vps6gvxDkCTCw0lo
U/jY8AOu+0t36ALhFZ+wsGF+kVSxDxR3brZgt1ueRpqQt/rPYFmRIpxJGGtnvmvvj7ZNLn5jA++D
fPx/rmvbVJ0NU7d6NMv2t0MzCCrROkRscU+EMeGqLYde4wtWa+nXGCKqkU3Zr7nphMe4xMC4/Cvp
Wh7jXuudAp24AQRIKI9vSMGnLPhTPfmFcwiVW91s+TkM6FgeGcXrZaeA5Z3YuOqiP1JEeMsErsiV
dHoOmkGc/vKw5YyL8UypDTG+Uz8H3Q4jsn4GnpcjE6oOjJjR9+3bgldLTRMV5cy/qb/sEPOlM2ut
04HqZIogN17oaC2wGBBKA/gt0EdS3dHW8RkAZBT8sjaWbnlLoXDX14GQyEqFq9hnONZkoyyQicD8
XATNEH2tG9IyI4zetgNa5aEujIunYy8A55/u7rLhq94E4ZI1CwbD8AUyG7+fkxzalxPBGVIHlnxV
3xIh9+cn/CC9T2Y2AhIaHeO+tM6400MvcaNSfQ8S+VfSAiG6rZILxslfpK6y04aYEHuB5i+UtSfI
K2zGiWsAkkZkyJEVRSrL7N2fCHsTTGK6HbCWniGBxU42525bkVeAWDSDzltCQviHKyJOVk/KtsKE
foJpholtakdIpMejR9rAoe0CfvOnahey6Uxl2Mv/AxPmeGaSlMfVSc0ypHlumsz1wfZc4lwMTc6+
AdJTDMQXkCCpsP/uRMwtFYf6PnD1lrELCP0wHEFwoavU5CSxtYN0Tzv8e4przhAG7ztXKKEbwLjU
fgh2FUwe89uv7hDXn+h6enE8VUTvFS1g7AQ6KNrqQS4FwoSMST8JwNHK482aHhbvIC/slRwk40fk
IKEoRCxGas6Z7tszlma6swsdoxrWIqIM6vBpGaqgyKfKPH1eZdggg13wC/v/pRCTttBbK6PdyKgT
RkSaZqSj2MtBuhIOOpJV5XVaiIKJUfR1ZNIyfSq8OkPgWCpVKlGepqKUuduELzZ5OrIdEqLSZl/d
RR6M2jHONQHKse9yo6ht0QdElZwBkVn112de9zShAjDuJot9iBamXS5/drkwFZDhAyjh/5zNEaW2
s/VwIJ/P+BfrIuWoezx/d42dIYOrAH/XNmQg59i/I+KOUy9D+r9QEq8EQvweh4Nw7n3zcGK1wMl/
oMPUP+yHMuY4KxMHJAqM0Jhse0t6hmSUbIgvnob0PqhlZjAM1/eTVv2iD7lZaCOKNnCRkvar0nEz
jum++F6W64I3pXox0ylwBIazqbOcAPqQJYt30zwMSzvecsQ+ScaRpDre2tOxdp8ke03JGdC/8yw+
jZXIY6KtBb3UrOR2BKNH2SXvC9/9NT0ftWeJKtS3OAdyxn03NM8QmtZ1x+XsDv15w/j24mI4xAD1
+nx+Qxe8iE8czhJXa9gdh87JUFA9Pd7AEgsIL3c48ITKzw7tvhVd2ELqqbOJyWG80Y1r83ADzYoa
BSpezd0ND6ZFGEwedggjvgplctNiFDsXf/WyCIlQhrwNrmqtJlkSOXVXdWVp7BmjhJzgC98l3JT6
4iqbUXIr1NfyTLA755NBQaFei+LMSMkVR3wrWMWl7whSPcuWDOs9WWhYXfYdcWAGoO7+RxKd7qag
jCDZr/xMERA1WpLd5bfg4W/gnSOB3jBwwrK/HRt2g4Db68y/Js2PjSNqip9tSaanAVOWB6hrfN7S
7dp91PCqimhXRFqcw/kvePm0zH73RIqiYDZJ4seP3yzMFGtH79Q3UDJhXzo5wphbFGX/17mpguZS
I33k1cflXeVJ9C4qewMO4R3NU+ASevA5ICT9S1KgmkLPtl3JEK1obCJO/4thtHZi09s32llEva1J
CczbwQFmSvYJtSeQ+1KHjWrBHBg+qNmCQjVppCRUfoeYt6g+J/IGuI8Hk+xmKXxz3L9lrzUCi1BI
+xDozwYHExTaY4Z2YH6FG7OxEyXrYE3pUAvq+zKS1geshNd6dDtkq5fF5NGQtFvhi0XQUpydBRHl
m24jSYWby3LZ/K5rb7ZXd4tqubH4Z+YRXKOU+aVy52CuWXsEE0Ieo5LBHEakL1v0P5LgcrGDiC8E
Oe2Q5budjV8bu1pjfub78/pUsbJMFjigEUG3vjVA8jzCa2vDj/7b8xbGal5KWJP0cIUPvRU1gqSc
g5UPmD/UWCEqSF8Ixf3tL6MpN/K3jzKcYvH9IgZzrBQwKHNSY7RvsCngFlt17l+BO09Ft98Ah3Oy
zmIVTGa2IgYSrGoOHo6HqX3F1/R8t6FOxfUJT/+kzkxZRgQYvzCTRGMhE9qiWWpnZMrFtvSwmDTb
NJiSn2fp4mQ/ztVdAmWVV2NZe1whlt2NIhcaZsVe17eBrOGcnUJdpbhGchgnMEmFXoprRCrH+X6y
BlfWYliUBRMkdp5CJftf3rUZl0lnOyhtiVelnMgtpwBlWKuIuc6JUXW766Cc0w5bQS0k2e3hVKZm
iM/USNdiI9qHaTApS9taA2WkrkFWvwuuCKlJyn8AfHUu/1rH+ziOT+sQr6C0XdilfGQy65AsySaq
10NdEmRlOPd/z7JW+mTang8yPxpk/mvrEXkQipBpxhauLSvzV/ee2sXr8Gw0WKezq8QZUuCDbtSv
bzyP0WmMB6NeUbg1xnhDsRUaDrpnPs93dIPxwoQlK2v2N3h9qkvsaJfkf5y83jnwBFW5NxLpM6Cf
aRcdlYacakZFwQ/de0FGYhl8lLaGK9fVhbYLUWhbwMEaV5IiaMiF+ZezPovhweDaf77q6E/DOecS
D2ch3R7nHccbk/HiKFsAaxYnwD3/najRWmHY57Lb8iDYkN/qKS/gj5JEPC3hqQBoJaNc422QvZzC
q42f+1pnadGCdBP6wmOFSjRzXMCRTdi0R+Sn4zqxWY2BpjQHbAtD68n3Jc5/OkPx/1HNNlpblImk
r3BqM6nthRc09H/fMhjTsufEGieLYL3ndDcfTIpAcPEOjYqZOc9IAIrUTPSk87WyKxLfvVb+IglH
hMnSB1mO/zGl9LlMrPtBEek7jF0DvEjwgdmNCah7K0bPkplfF6AiKPl6/m1Ua1egAgRaV8JpdKkl
RhH7Tvp65Fkt1wyOAba3g0eYG9unsdyoFpu0McjHv25L9rrsK6YUUlsN/abcQbQa1/tDLqEUznJZ
n9Am8gaF4TAtcyeddAyKzBmnharcSfDr2S/sN9zi9ADfxdzCh/7CiXq/o3pcWabRGt7D+Ta20auZ
XlLQ5yllVPzZ639DfzODPW4hp7LB1zW3rM33MYhX6suMO4I90uiwpFeXScEqzZsF0qrYkSV5MWVY
pCfB9SKJV/KlNu6sbu760OrD3Nrr7mSdP2zaSgV3kORml8k/A8bCPgESvTB7qUhBajdOZD/oxtPy
bQn1AQo7dxU7N8mbebBIajndw37ApzccaxITivQxmzDE7QH2uxeic1ihOP6F7Cq04+iOwEskGtKg
0BYrnN4lwp2NIEzZjNSRRw2eMm9wPMuRSUe5obIAY9oELcFFgaFsgV3db3X5SYMQSZe0WQUe/bXD
3HihmIUj5h0mx40o+QA2d6gli1jcqvakok6Sotn+DPbNrZBfDc+EyNeTiXbcjPYZlFFzLahI81gd
JzGhDXGC/vaJPkp+xeS/jbD/s5BLqUCCt95EYarj1CbD/7f8GPxKeKq4nwIgTb4TozdP0ZAbBUej
UhA+1mTlysY6HdIAe6A3pLY6Y0KABvfqi7QkYKhh1Dko5uzhUOWDFmO/BkkCvFp/ULCtd6GxWCsi
IdjmTzk8FoMEZVLxK+dqIW8QwPN8OIf9/x0nLvq79mCA2NYBehC/y3sn16J0rZni8udK6XfGegws
OG3fdzsJDdw5I8N1W/YuJQ0FVJ/4cLt+dpjSx7KMx3QVVdstkLlTi9LOYjbpSdfT6trFi0FGjqyI
4oJtvD5rev7ytnyIf6Q1PAgx25gcuayOTZ9S/IK/eSaFuO8r0y1vwl8g8INVHCJr8Estgk08z8dF
++SJUd4zE8Hq8Ph4Wh/chJopqBsJW6qTywvjX8iXKveoc8XHHBwW3vu6ClE4Gkbqg+1ktj3FJxOv
Rl+qnMbnn1lKb8+gMgdz+VIPt9TLjFP7Vlw2q9GDHUyv8H8Hi57jeQ2rslS6RfChql2qhOsKbJ+V
hxNeAW/ETGYM3V2kVe1pmsg0HQV03jHWWdlzCkIJbky3thHYHDaHVm+lfZPWmOsbkHpp/Nv6DxYi
BBT6koGpbtgxkfOOT0WzsKiZq8xbWBulGf5Sj5nh7SzvuIoY94sycpf+I/W94loJ187PRhxzfs8C
TgB68SwWJ3Cu/jfzJLwM3Oa/lG1YORGjFcMUqw4eWKhnBqbhFI74C68VeFS7Q3o1tj+jQDdchqWX
nBfPgp50t4EC3HytSRqbJ6KXRI3WogZg3DrtpBeEnuv50mnTxBfrykkY9A0PevdGNyR9XWKx8nid
a9rbuiCi+Bl5Ozal0deQTPZBOvfQM2x70SpLtmK9ecSPsL99Pf5kofWBN882IeDcfn2umDyks2xK
vZxORdhtjvah3My4tVkFqNNsmmHzop+8eehuCYMX2wFLTAiqDKSOR6aXtpNFYclghukXU8PzlROb
xiMLWzJzwhqkNlflGevZaqCXy03rZY4gZb1A5QG2fuKa702W7iVEEqhjSxeCSL3DDWAaEvwIPKo+
tRX8vz6+mVk9RitIB5LkPO3j/h4R3qqBVh1Tvu18bCrqsnCO6Qe+O+lHJ9QpiMJAB21GScF0HFXG
p449rEDzl7GLGHDdUnJNQh3B4c9bjQDx1bYfxs5RedmZ5uyTrtXhgDmxBxJTQAzZx7EbW9+jmNQt
vdoTxSNdPRHONkqdoP0t9nhpy9Tq88PsGNuCwvEc9fR2KuYHq5N1+2lyg7QWfAYJ6HLkD2+meJiB
QGOQYifmFtNkpG56HDp9JYrmhofKLbFqTxwcRHv9ZJU8FfShzlUMDQdysVnRkEB7tx0Om+b4uzTB
dBBTnVDB1KYhhK+1pPhBu0cnR6Ak0VsXSkwxx3b4E7O2zovpMNVwm04F4jyRC+n27UwwHdhtt+T1
U9sov1GS5LIfm7nagksbvNJcoPN48W6gtjDUZumvrYkFAQKqud2CmKxmelSdU5C6WK8HuSMrUK0E
cT0UmN3sz6jZHSC5kN7AT6FVZnsbKogkAULl3pfypsnakpeo5bGqIjDAZHomLgQwIuk+XAoEoc5K
5cye9gv3EKic9CPeg+0EqzkR/A3TGrWDpznqHjthdAeYwxpSEiPXN5mr23E/sN/9MpUGdmRlH1Nk
FXv8bb5TFuoaQJ4wNvTXU3r6gPhoHX+7xzXxqbLCWVuzcfs4XOYDLUgvISYLNkETSiaOgecoEYxX
7XLI0ra1UBxkAmbbGms62WcsSufdS65KprNgsSFc4T5207PUNra6BiWps1477Q2cvHNBJ2yurw9h
DcA81rmpBZiZU1x+d897ddV9hggMu4VrWBoJy6yUVkBvcnY61+Wufy4PaHkAk3QXOyL0SNZM6Wt3
jrJWFSIKQzbEqVCfUsw36JoU3jcXQKLrBQeJd2mt94Bf1Oj66q1y5nrwm/vNkYtdEDBj5vK3YLtX
ijL/IRj4qsZNznzwqOyWwU530R3udqqImkBqzz3whuNpq8wOS8xyXHRcFRAyn6AbLQeyVig3VARM
STVskujty8t8QPfHupQPerwcK8n3I43yNoUfnf8Zm1/skkuobM1IpIjQ9VQdLelVP/oUAb21dUDG
zMKVHuqEdJx7e9jkX9ccRk+PKawS3l8/++T8n7Py73ALYVLs6BZ5zQQcXhZxTwrD2C/AwzVK7E4b
thE/KE+E2drp8Vti9yef75TbMwFivk5FE+VcUoxvb/HN+9eJT0J7qOU/qZCPsJYqhPNHsNe6sUE8
lbk3AO7TQagr5RwiPwMFyXWUPFxSz2ZT4aNlnEWMX5DhTuke+gTj09+w632fWU/c7qVsRn4yyc60
QAhs8v2aXj3H8T+PAC7oezxDEKTwhAD/odYbkATXC2h1qE9V1oS7sXW8PvPvzqqwRd17T37qyhTN
H0MfBRrWAcVPsA4bq7nBQ/dUX7EuPBOPvlgXy8hH4xUVaE50X8ZyIVpla9WN6kKGCx2m6dVyKf9g
Gb/9yWYnHI6aoYtIUgiKwIeGAtSkls9Jl04Lq4K414/ch36XzIk8yYlxX42gd1EZUrZEuRKk8g82
BKxA7pWSJ9HYb27nQYYKHexZaJOvh6xYiZZrJ0EUTVJauDnV790P/BkzPLbtg/bpo2HZtPLBOw5H
zn419wFfDWi8/pUFmkADtTVOH+4kuppwB1VL29tB9OXMC4j1XQkkjqygUJ85OQBNp/MBAeC5+lFi
Sn9gKJHlRBNI1HYYEeopR0CcsmPc6nmo62qI9O80d0zczEM3Z6NuqB/28IshZMlYzBallSHGx6ic
rEa+8L34pjaLiY0b3L1zaGF3ES7zOiTXnvgZNdclR7fDzP1x4PXmA8BQRu1R5x2cUv6g/XeQQ5Mm
dqwLK5KhKBwVaz34C4XWVnaQCM9tWp6amj5hbFQalCXCcapCavdV1peGS+VIyFo6tECvz8Mi0Klj
zYJ8nR3F8UvIMAEvi2F3F80VgNLM5/5vYVGC4VYp46Ddyi8Lt43NlDt9vlcfBSRURBDiA6y1ZBSl
y033a+3m0H8E+BBXK3d5U01Dzezyd6trIgQkWSRJEGH7XD1RP+yIQLtA3OFI4DMgz4n++/BjtXeZ
pkQZ9YEfQQVMCXyUnbjQcDx4tKOl7KHCHj/uKCQK48Q2rlRMak29CdqNLvO8CFZwto7DqGc/QacO
hedbQ/uqWA8CMSMktWP5tHWrYo7RumW5JtwCjQScyNwkn4+0RbDl4xgQvkDUdx7j1S3cOlvLCsFo
TWeqAvhxx/PujFDuzLmeQ0279g19fparPO8t3aXfQnOz98a24TfIlgVS/PnA8YxFIgQZVHx0lzBn
c/seSRxE3d2NZrEQ958WO8nuR+Nwn/SXVjcCm2/uurHI+tMmA9PgGtwfGRgR61bHk3P+c1RYDwSz
QC7Z1E/qocVMdZcOmpxxC0bTLJd47PV3qgCfCauOmHQ4udp9NNbAHnxUpadfgJS2mgU9vgBLxcWa
FnIsZhgINR65X8UDJZNvFFAKFvnnMY750fcwaBvp0GMkSyH5UXBVm8VLCQvFORb82fcBq5Qpb/ol
vxjWfEiSq9kqTCavzib2k8nNFJECpt8zV7P0grbHB3tqpm/m8rjDD9iQBI73zS50QcC0Xc84/0Rt
OrOdv7IW8mtb9Wu756TvTm9vhpbMpff9DagMvLlkMH8bTR8JLY+5qjMHGER4CZKjMMnnGH7LYOKS
dXjUBOkTS7FXd+Bkkqerrab+mat5D3NQGvNanpqv2bwe7+OywDgAn0mSReW7c4nQUOEwO2dMnlF+
LWKTiTWfkBRlcgW65mAULr8LQ+Ye3/0N6OJ5hi/SuDY8AxdcyowMAQMfy6921tDtvkmNJPaOVBuC
u/qu6AfspmxqQVmV5YFjgdkhKedhh21wGNMIRqVpNleNfRSB90JShQmv02hmb7+RD4mjGS+Sm5Wm
RevmIdlY4fO9r3lq/aUGqox2+wtRNkNz+wyIQ8Gs0NyKYBS8enzVxXt+8aHJjzdAdlyu7Hw7dDXD
pHhJzS68ovS5idxRNseJJYwPy9I5SYEhEEzBwq+WzeiPwlMc/20naxz95RSlmw9Cpi69jYVcEiwv
S86Rz3VGldvxhvqhZrck4PyLB8juz2hrapoZmga3lkLpe4SgNoODRMErMrHn1LMYgDAEkNqmTZAN
qj09BHFhpda+l5zdK0AK5M8a6eHX8TQiL65vdoAG7sUNNlms1N8WU1cDhOxNxg79qyFhipObXQrc
Gq23E3mf9DuuQQy2H0olHq5B1a6uEAGPeS//7+iwxw7MtXB64uVd+IxtRCb5XdmtfNMHrl4EYctm
E9EdTEFPG/ref0QI6YDXD4+WduCfBE5IhAmZ5kt0fOdIcfAdjlyGPBrFQb35ax6AJbhdmSZWZWo8
HqPr0Y4dYR1TS5q7z4LwV3ZySepZ6sq1naml4Wqub6Ir0idDbYaEGL3kWvDz3fmDsDwnmFTTer/S
99u4U91VoFv0jnAGmMTPfbMXRJoWFk0upcDFB1FKIyiOMb3m4rglk9wn4s8KRaZt4Zd22URDFOXX
gYAu5ljZ/frrHYldEEL3UPXMTKzhiGmD2GCXgyOrZEcQ/YmhTdTdsyJNI1YuMvx/EGpMbMXSYWyj
aK4t10ivJpDeiMw4S6/kK/hYL6Z5OVRRIibv9kB3RabAhtZk+FTkOubqJMtPznXU704rS15RRv9K
JQCPKEvTfWm80W5ZM7QWZscLm6vjpw051VIKWK6UaGfCsG/QauGnP8/kaXEswAgGMDM2H5ina4Uy
FiV7l6EgfZsO6gC+iHPMPlOHrz1HobBzHOPIBBXFm8Mldnd36vU8Ee4zZo5kESfDBN7lSB1sihTR
hONCtwR5gRz0GzOwt+hgh4L03ReHBKxDA8Ire1NdwGA1An4xkHot60lRfRpvztI8H5eNQCheZUuN
jQ0ZUzqXMWX7kFs9QkjbynjPLjdjb7oy40dwe3GYqua5rPlqMb+Lh7PV6guiV6sDb609tGekGKVc
AI2xyoL6yPnLtVC8h6uOWpFQnLRwBbdN5eElqIFrR0AkfyanGy0KlJgxOcMwcqXB6fDX+6yIgOFr
Utgxlzb46b/vse0ix4SoJ6MQkA4VpnzAcSz4samnQ5kaCyRf5DakkPdctik/dCnV4VYR3ywRFsr5
1pPBvCKFLfSljgc7GALvD3TG3T7ZwY28FvNIpMWZxJyHIfKU3987RTYcxP5KRt4zA5B26QqxKZ7+
BItK9VXG0mE96kDU5+i/WWHlExJosF9IcIECfSgTHD3lmqUK2AvfBIKOGrG6yAe8pdNKEmiGovb1
IHS7hqC2+V2Evmljw1fkMirKt0UFAkZca7Wy9j1jxc83lUQB3Ngq++Rb9TZiebD5LZa89e09G88g
toyrDF2MaC2OOE26go1mMipet7b1PiYvtmpzicUHb+EeofYdTH1cM4ynwKRJ5RekgVtO6wVKjhGG
rqFvbIzDHm0q3gLAdQzP7naL3mXCOtrJXfFNra3G7GAY5Q+NW2EntMK9m8phXXFqNa82ECl/8Uaf
ThuFsqrre8eBI4Q/9TbtRS29sF7hRGQcNkvmPQUu0D1bgnRj5zHDukXj6wswjcGBUnZ2ImND0jek
AHvuKtd5qrQIBQHlJ19DLs16H+upwgCa+XKIHu6fFnCcr+xRA65zmR0VjEI0wG1DYZc6Bf2Lk+zC
fCyNSxwyy66QD1smV4CgAoA1DkJfuU9ilA/wFn83fHMfYyi47Ch1TKoaZ1JHbCuDoPRA3BoTNbVs
UvL5kXn1mZvSA+kpGOok71lKPHhbqxLEzgOziLKDUZFITBAYOFgTg9kN4o079u/ThYBwN9EYTI8h
K/kOBQ/WiJt0t/S+n9njvAphWyjqP0aNq0f1J42eCHQktgATy3hONutS8QR7Apj+IfXjbFiYZRGc
l5pUf1tFjzuhhOYH3wcOp2XVOwDTlAKhdM6MHaTwKBnZ7XXxL1ClPKs8kvNcjsxGdjQsjwOPVPdl
iRe4scLCNwqRz1eTiAyMIYv4FdefLeyQXL2IsOXMXRFlW1wN6kSw17EsAiTOJcObN0OtliGAgkI9
yT29g0byjqiv1FowwAVJw16Eog5isDnT0hqFLIhi+Rbkjfvrwx/OAgx3riXV9Zq8ZJPUBuktJL1w
xiBmJKR49No+fcOO6/uQu1wQOixYWp7U/WgBIsTJ1/spu/6bO0AfCd8f1wZRlDIYLvLdRTJUzmuQ
EdqWY2jCAfkYYZJd8tjGfUgb6jtTNwfw6DrimVsWb/Ff8pjAFTadkdzZ9ZSW74cMLPULgyhozcWU
akp0ZZuZNTrxviEbuekaE/E6zdhZuu3LeMRGvNENQLl5IbhMkGdJ3rQHcJ2vZlSDjSItIsQ3noeg
q1EjCAh/4GP7UZUbRhUuvBPZuOiufXPQ7sDN/7htCNjbd/FJEro0s+t25jBzbEpGEL5AX7JF3RWw
o9OYC5Kd8uAuhH54poI+NIU/wRj33Nb9IgVccFBzJisyEoVkxdiqW+L0XLXhNaNgxHx3TxewGz5Y
uKMIs8oRJoDz33Gzf+7om9wmKEoM8tswYTogtezWXVT5kRuHFhdq1EqkqstmCX/PvrJ66wHSqmh/
EdGCRCMghPdV76wXXG5ZLsdLcXycDJnKZE3o8UdEN2Kf5yzkceAlbx2+u662bqSE4wcUWFrm04Wx
DCdVOPqqQnXrNwJ0Voh8fnfXCMsn7R0HjHTq80HI/IRWYOYkBB0gY2kWBbZMpGLtUAoY9Mf9cAwY
FJymKYWsisBfDk5AdwPsGu0TQb67f2Sq3zFHKqXh7HuuKVLHDEU61yNqKjqAd9u0hBJo3664wvlC
yPjgOZLIFu3dv/XzeOo55PUxDhCj09+e8+uaIDL95ggA08p09yuo2WbtYOCKAHWTTbVrwM311ihm
KAm4hoYLw6h0+O09gGaJTsr6HvOnySppDIhoE5biqF+HABYQlHi60szeNOTBB5hno4kyQ6vmTk8v
91GROvMYUSzFzYQ8yrRbWBswpoi6Tij3cqNizMhcAnaGZQWsXJiA1caSsgaii20zpy3IVmcvRlvX
gsMsEVsxM/YmqbTuoH/m1Ldl/b5KYeZzYLRqzdA/7wMuPW0DzzMoc7oxYeOAdwTN3dXDYgMTblXA
rVj0islFw+qGQHXf79UR5uazJLKTMarE622hSOWLJiK2naNLbxOWxjnxd954IWkxP02fPoFLnMvb
6efpekO4alKz9t2xOB8kJQDW8Mgq0spvIhKSRfwjRk7pKcuIxxtdRI6fsqF4tKaBD6CyjsJWUlX0
3Ohx6docMCDMy02WnWa9m4dZKy25sL7mbRHtPybpRNB9a/X/AUeGD1slssionxtd4+5nkxgkw6fu
cNbtl86zUDc2i+y57Zea1sv6gRONWmA/+IkDMGRsaLHExYMQ/YX+5tIRqJ1qgqqJNxzBZvn8r2DK
tQNEhlzPlUKIDluqOTKdg19LEoriL6tqyrPFwWLcI8l81pus1tl0I7095Wu3Cg0sg36lMJsMSA2E
fOC2SpwCqc7QVuz9LlslByJXSjDc1+/Cuc1xvmWimY01/TgCg8QPQDZGEyf/YG1xVvi/uyz2dEA2
+6JrHjaeNwNNAIUrgnB3z9yTI5EbgaCp+2+KvnW/K9kvfQMcu6uVBOduhVfQ5wpnbWbx2xv/Xju6
nAyG/oPyfZOPu/zkAUJHeWQrMzSDrjAiZ79L8JYglay0UgoUnwTN8L69LcbS3fHrPngi+0/FPgB9
x6+c5yUnyE4QVRyTyIJcl5oSzkJoEOiNEqJWeFbCBJS7Pp3SZaapHWeg8NJp4PdRbQYTWAJyj2FJ
fXVx3oxm4qxbhOk7edP9nA1Lt9nea50pQ/FlZ3BbXZ3mSnQXPYIFLEyoY0PYldhw1CI2Y5SZ+6L2
88229+qmvWHnzbcmV6xrQaNDWt56RropMfoymyTHFVFo3sPbRrKiKafmA2rvRKEwepD9hkKCFBKq
SYWN85uC/HpFyYXvmEUFI4ySEc7RvvkHEvn9hHhrDnkqFrjH7pI7a13P6Y5T9HlaAY0OtzsCpNRE
Y0Ez04UNdNmD9Umd/uk574zdwi9m0LZJJXEVf7fezeIitXuLfWJL4r9fVtjkwSkEFkkHZOEI+v3+
rCE/rJH9GFP9FH6mTyIMTD2PuCq2okHqufEWiZF8rF66ppQim06B2acSMZ5QZX3sEmA8DHB9oYSy
1FSCbWAAV7YqAqBn6Cfp5KloEQIaxv+D/2D8E+S9qsoKVtB2wDytqISppDqQ2h7oA62erFdoFDXC
PEh0FiWOCFAgsEN4wIyKHIJBXpASS9jCHlsi2cNTJSUqvii13AGmzgnRWm1LW15Lt6LOfzweA+SU
SPse9FNswCnt4NL6BqmDLg4OB6DUnX9ZGKlFRg++EpXn2IkYR3w5xWXTAZM9vVVDphIlGdJvlQn6
j1TThGcG6YiJt/wQC3xTQ2Z253ic40aRSoR4IccuHlEGubyYDonTHsNWI7nVKJTU5lBXysqdxzpN
jy4aYU9bsQLF+vJjmQIekcG2Q8gdggTC+Sjm+0LKOzg/Fp7aKDkOD1LQ7Sv4ytDIYGnVO0pRLION
3yf4eMuhvUEg8WVGCI8rdCweawXoyIcA74wC+tNF1wpsEzMSiGDp8CX3j5YBB3ddp/UaxX4gnOJH
E6R2aUninXRw9ou3HCfvMDH/By+WHS6S7PiBOoupirMiWfZ6pHEE6yoyyjQ2WVyfx+vZg0w34H+c
EFoBjhzOt1izyxOsbDGb+9xhog9W/7OMj/b7tKNHwADCnR66hnQGGd5Kho889uNCUCMHKBeC2Deo
jia5VUPDt7KrQYGK2S2zrWX1HPaWvbqBiETO7BW+l9O3YVH6XKp4lmtItoVBXYV4WjSEO/LgENUi
jdJu9Y8AviKZOqDHQ5DjUffKc1vmOYCxcVJKvAwLzxibc8V/8Sp0/KzUrBCzuB/rsVUXcptAhcgk
0OMtEpXX0xgz1njAX17Y7XMS7wtKpNjPGJd1Jp621PaKt/cjUKuFe2afDs6Dwg1Hbv4xBVDlvekH
lN7VdwbL0/6oSOqPAlOZi16OC246T8lwAALYaH0rl3BqQTTsqA85wt0LIj8ZqBhdnkSv0OdAWmPS
in2uQzwwzeDGUaYXVO2tw5DjdKDiN3aWyXkCkA/JF4adWbeLj+K9X8tMK1FvtBIIIVS4oFaSBMdn
mYA1INXmT70k4J+v8vaejtJ2XXCMCVJ2o1THEZSgq9AivBuAb/3baa7MWbr8HbD1CMWkuyGFmjyf
jJrn0uHH+vGbztRKYW4JVNmkRrFfjH0hAGP4nxUANB9Yo0A0fsN5k6Aii8L66rpNPOCBbsozlN1P
JTLiNZhUiCR61e72tyrn0i5O3S4+8I65zzf/OewTQNCcclIeKZiQYkrCGfwwiu4zW1qzKfHkC8a6
BELWUYHlgdl0cNO8Cd85kSEKb3bPGbYxdWnfB6qQ2Xxlz87oWvv304uNAEr75WpyMY5hEcU+3Iya
2ADZB6Rv1iiI1ifovK1LyQshUqx2Ku6rE+2atktOhY5d5scml+VrVq1YC20tFH3Tca34+0mz04nD
PH+x4qihAf1U5pvGwkt/AKRptQQPtdyi/tKLcQpxgwgJAtA/nf20hgf/66pOrpznLXtjAKQ20PNF
hQ8jcDvv5BFPSRHbD3baM2ceywc2A+S4/BO47zvS9ZlljMrGjHgEqjzN/psCXGWBNn0mhZE9ywrC
mtHkfHc3+vqxb6k1jiu2mWI1orj3gbFkMsr6AVOS1YO00YbJ24Il9yS2+38ilvREEs/sc2r7obND
5utdfTxSBYUnaoOeYfElxJout2MZ30KmfgVhy6GcVyyQm6Nfl9POIqY295zx/kT24f1WtKthGRqg
DrfZQQLKJmIvXcU2v5PPsq2nIOg/K/xEvHadUekasyQKyPtKbGoJBYoWJhUWO8uDZgjDM2CNxVH/
sGVP7ED4dCsk9Jhc2QqYKOVXhhiTzMw/A6AF6hL2TTP5HsgRJQFyF7lesFuYY354GO05Y2tofIGF
usj6KwqJJm8PoYc0QODPsfp0FOvjug6qRAXecJ1NvSjKiyBJ2dK44AQ1YxiMakGROESlNNfeIfha
lPaAJGuJ78wQotcgFdtt73iCbqsXzJutUQQBnGVsP8IOxRQHtsw7Y+zm+eKFnAhOzL6AwUTOQhMh
o/YQQgPQTTK11i7UTUfHpqsf5tLhScZIV/q9MLaZ75OSTt+arXVqzAAp0dcXPGYx88h/QSExBBb8
B77Z/ye6Q/VnwMHsS4Kkk6Xuapd983aPDRBKmyHnXpJtfNw6l7Vk65xiLrIyixwpB4XSZqJAwY2e
PR/SgPWjslOHr+fxfFdzr3mdXF+0mCDjChAtjcQcXOxk4bMxjjBcFhMDkG6WIR0jUhneMOd9b6Nk
5aey7U4Ub+tiXIi2MTMVwSeAx82Q24juZyanJSaXS9CGPtOMvNLZ+gxkw5jR2LgmDuxW+1V10jKL
3woAhGndiiyPpPRpkIQfSti3+YLvx3NEoJCH5bO4Li0G0qtytf1IT62Pj50AIypa26YAI0h/vMDp
eSwo2b5i4tsD7qhEPk4MUEsfDUONehiTaxzDQWWKJLj+BXLCh/Qv48xzAaQb4cIGk5iJ0YgnW+Up
Y4Uh2Zxqq0RY4bkiMi4cZht1SN2szpVbkKTUb7RQMF4G2+WbXbEClqFgvYpfICuNncVafzxnJcYa
1Oh0PpP51b2FXDlh6FZuioPmWlmFcoAMGW2wPVlTyIG8BuTYFHR2eY6EGURJclpmoJeFgMbvb9pz
1mDoVkmt28/HiANhH2MbEqZohINBWfctK9t4KtZKXaHiBOeeDSH4YaJvdvuj10yn7IgXLclahjsN
reP85cOROgftrDd4xUrUda0cSVZYGuOJkjXAnOXxmtiU0MGJ2Nc/AzIfYm8fRm2Y5QOlVWttHmnG
394o2VMG/HRh32ThBBC0gjS5HlY6j8w8cOUnXqyyRdSTS5wq1DsQT1p9QWzclB18/yOsi5V+u5F0
Pd5GbG+0uv+8T/XD1j8bB6Ugk+sRQ6sijBnzxgS5mBqNRQFfhAKWsCs26n3YgAZ+DaQIq+BSXqKE
2sMA4c7v2WQcEBIF4G9xIAYyYXKJtdohM+2ZJy7IwE2kH3cOITKlZ8LxSu+ik/z/gtU2NcMFSjPX
DEFANNCcHrbMMGUUrgBks7VM+BKaVqsThxzC1tL4Pxo5LYlpf5xLbkFWMUE+G/SIFrUGlx8fRXhU
D8RXTT5lp5RvFcYxl8GMRC6ilb7vFMlV90Ee0h89E6HZzt2A43d8GzWsqCj8IzEd/JCit9En32bt
SUC35p1KZ7Gi3bhrUK1JvIJ/fzw7qLVvYv2M6ucKt3deJYPqGybmYR1pnRT72CQqTxqyp9C0Dbvw
nAsn8NCgoiixbejnOPl7mfIXMmkYtkmY+Oki0/akGRSwrlbGX85fWi8fiOGjWSfvrupLvGMHB8fm
2fgMTPNueJiISpg61O6c5FfDoK69sJpzwXtjbKhyirGKcM5dLqTZ0MsRSiBCyQ6TSWwS2GtLTJLQ
4KL9ZW/BGXsS1XpVjYO1ujU4BbKZZ2u6Q5OBSQh1UZwFw3ihLh7aGIgiw+aopGQ2xZNWoSdHSSXc
eOhHkRLpIiHinj1idinzdoe8kxYUHhcwFpaQ4Q3hjADzEqmTylDVfYAjI/V7c2ZyswewLMkIesok
r+NQstgamJ4LrcRaxr2ZTMJ3G6nLgblUOOSCBLzYqa1hpWDc2G+up9L2KvxOJmf/OFJx2JW2RZJy
+z7M9F1ojbCUjD1f3xscJTQwxa2JZfNlnkpHgtkQRGY0aDT7TyJh8sXADe3GSD5PzT6fd2E0D4Dn
jlVw5N/sWTAl3kZpJyGepXjJS8waSXLsKMpKbqRMbvVAVpOB3/N+Sf778aSlQtF935F1ncZwkycM
5Ee2lAVm2dklBIZVwde/BtY/QDjC+Djt6dujEJOb9Pe+kHGHiXpDIC9q6FGNhyn7iKFOZh0MoDZK
ayKuqPn3OatDtEZ1zEmllkklbjF/s5vtUZoVTQsbVKPK5hvuUORzDdZYsynEWdZ8mhkkSN5YusP+
VU8cRLyjW9T3qdJ3k9FqyPA/+v22jGfs6RSNyMlFMX7eV7OgU/kiZywgb4WaknDX8np5HGnj3QRt
mvHzwF7i26I1dFLjrICD+a6tLHdzJ3856NQ4GM09xJqq9//Wys+8slFvng6K0KOBQyYVpxeRyVS4
o2jYvLCQvdji+UTkVcVCSyp6s9F6pQkRGSGYwZdRa1XP5fNo5kuEafr108SH7E6lAHFJc7Sbc0KK
KnOliuniTAnBJqZbF2Ug/NqytTHelO0kh6RQRdQmmvWzzaMsPkYhiAvo9YFHYTpjitq4rULeT9Xn
0VWcTk9Yr68MMqV9QXVcRg9Ei3hPzONvbGie+MqpGowwZWGP40x3+sJO9yIetOE/00q6Yhij3X1K
bqxsSxVSMVHDu6nPVU9aDA9ISb9Rw0sA9BzKVkiAzcRPdzfxCkATBUclgKPcyRl2uu8v/WqrJ603
sCld1y8N4K0+B7ZzntCvYPSHjVELR4ZVXxWwiYHMO7+Do0ujhFc94XFhJywuGNf95L+Lq3I0aADg
68GlwmBkKZgNSubgPB1ztSYKkmtqVuMxzabPUxdEBc3dsa5LSVB5Q1KCJUE1GbGJa5BgvHvzhNFe
9QWD683okCJaD6M9jwHRHS+x2ySRRXl7hyeWH657s5szcBbeVQ/S/jM9pvirYuJEVpaqm0XobVWV
A3YmJuC8eFDbnOHDJOIE2MNpn7YFh4QiuGs7JVoJrj4BJyKlKf4F7Xn2D71HwfbdGcxjXNxHRgOl
i1NCzTkI5Nxrd5VNDMXcIW2QZ1mTU63IqHSDhalUaZdjzjZXVXcDcRq8QOCesax66QCjMR2hL9i5
klC+3W5uezPYXFSorZUIwKk84RDBwfw/24kFuqM01iMizdvvhvlK4pDNSg8tdRX2CzRWBYOOKIPF
wKQqE1IyU7q/YXSGipM9VT+4Pc3x7pjKRgXnqgCc1E3WEUaC0ESHy9qnkvi+9D+1FDdCDuEDkWVb
m+h+n+jli9cPYiZCD+KlvnfyCo2bB+9i9S+Qk1175urbp6FG2NzEk9+skcnz6Kto0Wl/dNVDvBvU
3yyTnyfMngfSDh0tnu01CgKX9RLyqumdzzcZiQ5c0EC7hjYJp3LtnROwdHNM71tOVvC927UJBu+E
GkfomPKPQ2WmYCBzPizDiQuN9LMrdL+co8oh1sxL6U1PtRVBKU97Nrc2YhKYH2w7YQZQfdl/4YxJ
+oiZdS6N5I7KyaBmUJCe79xtdEGE7x+3qPYFA3qqiuEzd0pRj+DUI5+blBOX3cmdGIRuE+NQ063l
yrEkskUAyZa+44wCSwgHTHslDX/kpaYRIJAnu7W9/QtH7HbLMbzAX+Zlb6ITbbUXZ/ME7zoLCRHp
1KeZScJjCR2SHuUazABmuwhIYN2rhS7MnWPOv/Xg1jj3TW2DEJVazAyMmQjIr7Dwjzjm69nRTvxi
xh5CJrVwdMXRWO7BB9vlnmAW1QgmmeS8F9lfTnyR46d+TNGQk0/HrqCaTUpa/kLluNmE/D03WcCf
dde4L8ADWlioKg+5co5VFjdh7E36GMvoM1o4MX2wDD2+5ksqZzMDfh1pVbDf8mclyIvXTPmue5Xo
/tvbunqCajOIUzkgpTEsDQoOhgm7tjPIf4Gj8fNyrbAHMiQubSuQfhUx/lE4nOFGFmDircCysTjt
Dcb/TcwUIfSFrwEYdgorwRCPHIqCvWT/tSwNfhTzfC9phN5B0zVZ9I0kEzHdse0V8dynxzM6IW61
QdJPPWqQBcyiKUsZ3HPtUiKSc9c9yYY1DI4CcnJ0+LZvRKpRDkYQV8rD2G0zknvSYZRuYdB3JwLr
6A+V7KBoaYyAWpEw9dDfrNPmSBankFwFFXR+kCjM42EkeEYmkO098+aWuQ9k9UMfewSLzPccr43L
t2TUYqBYx3Iu+kAAgwoDE9pW8ZnypjfkXP4BN8cC92yHVSaCRjXtHfEOAgYYk7Ap91DpHirDyQWx
IRqussiWzSopVaJY06OfbiFOwrpJ4b7uqD9b73TijvJOekPwywD/9m4gm3NPeVMt4TDjrzIE7o+Y
JV59KzASDLVEBHAlPCEUGShNkz+5PYAxl0V3u+/o/ZwOeeTr3eSl9/j53TrVRimvqJA+oGFCyePb
HTxvXLQBrK/Y+U7xaxBVWtdzxehVJsJWfre8HXIK3MivKA9+QgKw3k9q+6Yx8OBs72aivJAArUMp
k/k3Uo4rC9EtYbl3Zv27Rk2EmFmIvRv4Fic+iPrax7gTOMhoMPImlIcdLo0lKwzubvMe+CnDxyDt
l/S2u1BNQ8CBgSxaCs1OOc/hdJH+YU4s39p9FTg03Iw3Fbi+EXafpdVVmUjeVfIBuGRGvk36aGRD
itA+NtT9L4WkkyoFYub6zJ58bxHQ1hiq9QUi0GxujgLhlv8TPW1pi+LwdkDvow36g/egTzcqUgns
JLX6ifFK7LHstJ2UL5qz2H8w8EqGQGLBSKaNNpmHE6SpQVD2a3WM12RMlhhvjdZTwFENzF6+PAL6
AwUetBar18hCqdRs1rEnjft7DQTK0qhCdqRwcLOgNNiq8N6NZZViKMLFUjaVEMjn1AVz1ljDXHKp
OTtUSCV+5zSd7BdBtYr5u68OBAYwuswemqndPpPte7DKzLf7tfYVGKpmg3Chn1+0tPTANcXadulw
kZnXrmygZZoyfqUkGjdrMELPy1LIzQ6uhlPCBiXASph/08QO/csL78JPgfEIE3u5Xw+kUO2gKyuz
BN+nGLfhD7DqlQZuz9AVbCLJOwHieYpgNN5T48GubhKRYpUk5Oq2nvkpBItazQAtaO7fe6Lfa0Gs
aUrc54lhO1j+63ZsIxgkHo7OXChb62PWsHDhtzp1iJ1VC7apY9a5gfJJkNfI6Mbk5uM9qSm+V1No
DRwYFjoaQx/1z7lO23TFiSHyGjE50ByYe7R6kTsrY74BPSpNHmbwCxUACW4TM65ZLyaAldZm21EV
BrlrTn4c0pQu5rgFmGZ0RluGfiHrIhd7chpQLsSyjdSZoPrYV+Zj4DOEPWM8dT99mzdy4duWoZkT
03z6GbnbbwbE19C7hHWfm7RxlPulF7LPrc50ze6uuevV7wlxsHtbJmW/X8aqW7ZDdzfjBfnGSG6J
dVESQUmsdWv1VirRONKOM+/X+cfE783kK64fr8pYPgTzS9HoXpSRdTpYw1KeVgyB5dtqA0uJoV2F
xniF+RfTNA/FQLmXUrOK+vSEez/s13UFDibnUtuT1B9MUBTXiyOFqvqltjfysKtd3H9hmdH7e0uV
tJ/l/za4qmMIn5ki2M3EKZU6mnp5mhJl2ldKd9dp04/uMn+rftXZ+8C6vChC3Q16GPb0gDlhPXUH
qcYn2Gjil52KoVp9sAH3KKxwT228FWwkgXEzOorZNK70FtZ3cs71yyhF0pnmMq2mUghYxAPp9zS5
7s9WqL9UFH3+8Gpk69QFziKHPG5g5fI7lmHSx5VcGEn3d4SrJRVvy2eX4cy7MTUZtVEdWRGc3X8M
G9dJYRoiAomKDXU1+B45YuzNMTes8QySghfFHCnlWc8/w/LFXvfi7vlKJsVnnkGo8YV14eqfWYlN
CL3G6peQdrgvE9RgZjUeT6yB/b0FA1WJiO0z+ReEHjw3xNCiJp2XEzRUv3obpWfG3zURawvva9Bu
DioWhlUemKVV5QO/wti6xt79kHJCvQDVvTAicUCWuEnEZe5zQ3Jx7APXklbxhtpb8qHu/fIeiEID
WCZJ9zIFaRdooDSBsDqr0TO8096zr5pkcKfxmwdHt6jtaZCHDHXm4au6t0OAKgg0Wwlyz1URxoKR
58Vp1YtIrCisyFXLn8+rhyRZLuBCIChibUCoyRxZMwFP44HzAD+AYbN1CfWQK+kiBgf6nPRSSigD
0D3TfGHTqsX/riq3Io1DJhNN/LHr0qHm7hArKbQSzjZmHb5OSQaNc/kpXVALGTDfWVgdq4503h2f
cnmyoW2xUyBW6y3BJ9R7jrmtEI+MQKkuHmFUcoC0xlwaZS9Cn2/zL8Ejj9FiKXvGbtU8HUPfgU6q
80l2nuHl+77acfcn0hY494YOqD8/25BSTkCJxmEOzmfjQvYJM4+9P8J3Vj+IpbM2a2KOtUFJ05Bn
WUdKdbkbRebwa2sr54KHj46n54ylZ7zlDob6vrzJqL46XK3x+GZA6PpQZqqpoy/mlzjXcUh6UPb1
93Th4BbPVs2riB5jHTSXVICo2CqkaJKZAqnoIo1RAkBEeHPR/L0lA1VqvFpIIfOc8lJXBTOTjyzg
IaNddDCa6s6kkI82AtPKBls4+G5rv5rFA4n/IQi5RbdaOYGgi0GVUWvzmKywmGWNgiN6xQ+la0aM
CsumDMgdd0YC+hc/wb4+npezC8HmoVMiaap5/xxSchYTfv8CPx3QOD+RfJl0WfrL2BuAmaDLzhd9
Q7bEAv/cbt8GWCQYedsHrcwASw/z18LvNWpnc9fhayjdY/GqAfazos75RHQFHXXEXqUNukvWhwlL
g1clXEEU+qbzwpATuo2U/1xMShyPl4kCvgLKLAxmbQ3BpIZPwGHelt7j2VAHLTvS0lhGwCSHub20
h1M+MdGMQ6sdv5SNBymFohTx9hWLAC3r5RzWWiKBrvc+YBXIRLrHYmPds+E6KR01sxUIB6xATHvk
thAPx33IE2COEI1kIWyGd3FlfIQ3fqvplAQKAJVm0E7e+hc1WA+jTtPuFSUuVKfDFU/rIm2hrYfh
T0i/FNqZBKiBWVEnYh9RWsokNgkHCSxw39qZJGG1soE129B1v5yGTqatu2kFJNeUzQR9/Q6blkjG
9O6FhyE8l+95mkKHIhNREuaywtDvghPG+SDuMHxF8wk+7dQCoyJTzFiIlAKiQlntDZRcePlYcsfD
YVS+fUV8obbocJpqRYCQW0UuyoeiE/RBtHdrSd7/jThEPK/4hCEGEecn9/YIT9/6U1iAdPDj3BAZ
wvxk5hlJeCsSABycIKCV/yvVJJDZVQj2w+nkCKKwWNDWFBiXSJYpfxCdn3/9p4TXbo9O2GJuMx+f
j/Y2bpsbd05gW847KM4OfLJ8CvjM0PJXjAmNCktwozCfWuMyysH22iCFz3xf08jIdXpBTKQlcP6l
+pubNJv7zWE5tLyYdwjs+eZ4t43DOEz47KiwxC9ng7/Ld/tPS3iZehY689FbvrLH+mswIE/dgw1b
d9Nklhqqh2S01vJFHqN8FZfw/evsIW/Jt0blMoXHxuM9SZLUCcoLm6F9K+XdK3Q/Spg03hblMLW0
Ln1q10faSVjX07HRHk56tYTQmdXHnJY8qThzmpr+caBf5UrtaLbLH0ENOiO88H0A7jk24TGpEOCQ
25s3/Ttru+uaDXu1pgl3L7gELvRCYl2KxrUlLtVr2ncyoO7xR6RVzctljOv6qcxH5Xb6aYPf4yi/
LeJpP7JNRdJA7qmSXiboCRkMr5JsVsvSTtZiowUp3wUJaDuRyzwkfOVFXf28N40QBHUYseJfO2uR
9VSzLXS6bSH9setWSVZ0qxaxU7hhGnuj2AXQh89dU9YI2xqleFBU9BBO7ri6WrZxcfeyOlXVZznJ
HTxgUeUzU9F0TboKGRVOUQrGbqeMMLS5j+BVaO7/95/qDrru399qTCCAbPhR4nBbm3YznKh9J2xg
Hkap0IaRKxPUZGFxij2rnY2x1eb8ZrEO0qMEWe9es+sKUGS/2TTuCQAoFu76JOaFhv09YEfh8Ndj
Mz2Kc0hj6+qeU9DK4m1qbrb58cf9hGlBKL0fcZtO1hNNlMaS9m97yp1qcYngsyp/JleUQv3KMVuD
ckCN+2zxRFP2Km9f+fiBfV5yFYJj1iEMMwWq0AROYdhFnc7DLMfkScAojXqmE9dF2KKk7IbauWNk
FF2utmwiJUgjH1FNmA4SSyzik6qKmdgN4kzAP3pohIBl20wxH0OqKgM3Iw9FO1ABPFskOWIxl8Z5
MNnt59oVtUFYtA4/Ypo24MrWULWMwsZnw3ZbKr5s+g0mUq4tBM5Juer6a7xX5Ef+YB+tZY3S/H35
riaUKoxMB2arQEUQfDT2LK93YABFvcbdivEYKRhmBuQAwwJNU4rGkH3M4XzUTkNTi3oX/JiGQIYe
cswAn4ogklkFeGKF+NJoJEkNIhGcL6AYg520O77WtMoCruzS6hkCtuVffjmbSrYRLj2Z0z4IGimc
kUAZXxqCVqkV5qZWwUQ44TDiVZy0waKKXdhMIZesHz4GbwcqFzshGM3tZelo9gARzMBr7gCyn2FH
AT8E2TRu82EiG3kznfOHBkb5rZBsaGUeE3vOy3r5x/16DcnGWcWQswZy/ohS9L019h/wP6GGzx22
tflUOA/wdkus6aJN10LRkI1DEwSCeasCfvJr5cyLGt2bhDF0UNXxOloS6zo7X+1LdIpJk/bBY38a
B6sfXrm8kwwm/eEmnUax3e+j6eyZIokWZzOC5YkG9oNHEhCuvTlAklLCQSR90GHsORnlP7ZR7jq0
honfU0BoGJzJAr5xh9J468X/krlIs79UpgpmkCjbvuP5YFRNr3lhFsAflxUNvlq2bt9NqKw7epW+
ZOoQpFHuJlzXr8ZguzAqu55lklCdQpn0MMAz2F8quKu1gcD8j2u227LG4iG7FR4AyM1CZ2JN7OCD
XOUzsAhQfgtUuoL08SwRjbC1SdmjOdNV0d4tN/6XibneYzXK0KDjsEyq8lINY+VZ/5xSqbjLtzxd
uw1/SWEP+LolPT0cT6qTcZ/jWMBkC6PoeDCW0NcWx7ILp6M6+Yor/9vr74KuzjZx42nrXNLPa6TQ
jDkqO8xQh+j/6GlKLyHw/bswt7Yu9LSWY/bxGL0IQLw8ESWLJ3G5ufSayTcEOnvPZ3yHpPc856Tm
lMHr3Lb+40EO91u54xxaGxlwIMwR+BixdD9cmSkvW1/BPJyKyl0Ry2fq0bOibWK78tjyFrOatmmf
ClOUtlRjMDwDRBJgZdEdz27BTLa6x+STVBV6uZ/IIQcL4NiGmc2kX8zmElfkPtXI9XML4N4kFJ5R
jxYtIm10AhjRUvUDu67qhlx9GPTNtjFFNxNWzgfFAHo0UoGx2FE2gE9+Tg0orOhDkNCIMpn+nFzg
JAcy20tH1nS9bvRE+wryxPjSWzQpUlN/r6MCMjUjZJb9FTKZL6yTo8G6Hntt7RDZU6q8mMheZrhf
ZSp5yUQmsqkBGBQ4gt4FQ+8b1ds2x05I/yTA9Onxye1nu7+RET7ZV7jKmh8yy29HesP+hpilgH+I
nB7C+xEyYX5HpgjBcIcoWm61vFqxlNf0dmstmw/TZqyJVyyAsIZ/FkTEFE+MiqWCE3Su3r6W7FEq
zQCJo2AVHcbMPVQT/+CSDVlbD2e5T89Z2j9XsJKdu/A8z9AaeNCNiIh1o+0xlEoqdsq+Jc9WwN1E
ZFOiR9p0AI+inkOAsa5C74gKigPvvDWoJntfES6GcvaJGhZq14LDaS/1i8nc2tJxvDXdE6dgxC9V
JQ+lJv+hzPVT4PjED8qRslUgfyM553yQ/Vq8zjoh8Okp6zyKrmj0JFMGrib7Rq+Lj1PSyo5cGFmx
ey76MZ7S3BkpvQ6yHuCH7alKq73dhQG1XDudX/hDQsSeXwzX6BQTawh/2TocK1f4loutiTndyqBv
kfAKZBo9Phar7Enw8+kzTRjslR4Rjo7ew+QUXV6MvjR3Gc52BwtO0IuGwIRWTYUeeXQS3RwrujZA
Os1e03YK2QoLog/WnXH74FZwX8W5QgG6Ui4Mre8JQyZT+tc+027r8KcSZfIJDcjeSCSIx2Cj5/M4
y76j85YhDtnC3p2ux7qjRmNcJ3x6UoObqZijKX+kkHY+bfPAVY0IvfuMsDT7YFNyu2chSSpa/+s8
U7bFlTv6qolgoOQX+aiq3QjmrQma3Ni8tAi9RU1JfvoMkSHLfHWtv6vodJ52kBeI5WSOTR24HSxn
b4wUvwuzoXBD5nTOjFFH6tmlj6gma1rvkWXLzPj3ZglcJvq/+Z0zBRSlMJ637Ex8wqYjR8t3KNXM
e3nAF2I7Duej/oCo2CAHO1xDjJ+x8TUPYom4A2iiXkdusOxLpq3hY84N/dgl/rsBeSZ9dVJLVrxU
TwcQCXZ6aQFw1CmTYxkq8mmyMdgwbQw4/6KZ3ksMO5+ijxdoqerlnAIxyLHHii0dm1Fr6Ossnx8Y
SEjEMDFbuyss+m96CwubS9uBItMyAv9oeeNY+eEuAVEF9Lcnm2xUfIuSfvWfbXvDYtBgfMNICVoX
zgkzzZUIk0K4vd8TjyNnvuGrc/Ts+KIjv2FjZZ+ITg69VZgIIeiXozJaAKpXasfCYyamjON5Z/x+
qKgb1hulM7fNQgcyP5HPPNkQuobHX3nQDhZDMC10tej5SeYWsUVCqPRiER99nrL1kTyBG+0qeGnw
TkZywpaVk3UUAyCgh9o5fcy/bmvp5vPuVRxHKblo5DkKOeVBzDCkzobktckzwX+qMRk7LWBI/ulL
OcL1RAxqPzyDJPUkEVxCKb9dnome6jCSIVs4utGu9KlmBVANpOgDPcpswJC7SLUUtvNcYZDmrKob
cYrRVyUq2gduqRUIA/fmEwRXPQJz5jGXS2ehzH9rXUYiqMUXW5UJJEcpOuz3mer+d1bApw9f6RWn
GhT3imhs6TBejDDnCQJOUf7RsWPG7FhH+tb0ZKDaj+tFKI+wpoAhDuTXUA5FirmQZzQPjL3W+LSW
HlZmmbQW3+KdSmYAs1NsmQE5Fziz4px4ypnE3GzPu7htaNaDqcP7OR6bjE2cZ/WZvj4nmAxWdm3R
HI69/PG50GUnvWwPCpL6sJm7gGEnAj2PITUOIgB5Gmt6HlIzkxywxBxlnUY/Kwp/gJWJC48/ZjIk
RGXJFpYITQTPbivfe8eoC3SjrMBTWuAIinjjqz18gQN2v9a3n3jxYS9wOAgN7FF9jRT1HR3dr09S
Rfn4toYMjstRsBwVDxFdVGCxDadgbEPIua3y2wJWMrSPILhG8ZXZnrBI6YW3o3ZwJHsg87GyILtV
QNP+3cOmT50SClzzrW8RjzB9wp7HTrDUZ/Qr1TSRDZlkHnsGhk/cF/HcsH8dmQiXKN3mzMFlU6Fk
xgmG5fjdsx3CX5k16TQwmUgJ3dQxKFf6LESeyzn5tHFZDZ6JG7ADlCuCFV0j7WVxJhmJlukHFjl4
TDtGYwJzQGG76vZiA40beJhQ7th+fQKjlPIWdtnrJdUwJMA2pTUFx2shT5q+t+Hlx05t2wj860Do
JNm+DNORWv6II1FJTawVThs0eX2sDe0aSUqYJrVX+7gAtFgweIF+N8YVgQLS/Ym57lMCRKC5Os/m
ZkD/9JQdPmkLWhivXBxU88QPYfnH+afvXF/Opf8g4B5lRSBjX3LXFZ68brXZ2TZgFRd73B1kpI72
KXgnUc/0Wn7wNzjxGlYWXyvy9XX6MSQhUlNsO3ZhXJCmPFklXvEqLcmCU5E0GjP1IYAnfKBIJk1Y
yBDvIGC0ilQAKYK1P1nJqRzugP6n5wLcWTJFDR2dfd0taqV+BPV4UeFm+UZO4NPSTh9i2SOCUmxC
v6rjMnihwmlBmEbcHti5O9IPGVSIFSYwQ8K8FhagBkZnfuCWTwIrbG6eWwrHvEv+8Zx6WWsObVNF
befjOBtGOTM6uuyAw5NqEd+g+L3dnedy+DmJHYKKsUpuMl3dEacM7g5jOjQKAbSUn7MtJF0U+2Eb
NJDRwsnW+RKWaPj3Ey/wBNQHQH3ddjNHQSEwT1ER7w+aQTORKPrCyFuahBA+H+VX+08xye3ZuPsC
7xVEdwhU5iRX6d3j+ZY3dIQTJLAUHqPlGNeSmIDit3QJadeS33yULMdioqbFMsBQBbuzE06Cz3d6
0WZBI5kkNUQx6ESYFZ94CBZxZR1aoNUCL3g1BSS1cmeC/Mv6nWJ3nv486JYrDvLOVeupQaBJ+9hX
E9C/AhoUbQ8uidpkusKEl4oYE0W/GuAh2H2P3gUHMaeV89G9MXP1+haqDbn6O+ux7jvO8MZlsidR
Bok5s4LkpdR0jtQAOOjTqEOQx/lY7lZAYHJSM4RKlfDlqsZXteEO3GVxdVezG51svyt3nfV1s5WU
BJqdZzoMnLCo5drjXJascUM2n05JFfjMcWUlBZysXhkNkf71JUpvDU5UIA5mZ9L/TB/6aC09za0T
9LhIYN5EMBrNxGBq5DRZuBv/xqup5phU28JHi+c3ezPLndMj88cNwcnwRRu9LmD2K32b3sSrMDW3
z1DBqtFXu2SOqpoPXn7IAAY2I6d1WKWHqaKhPQltQwThK/8ky3mpfpgR1upC1gjLVogvp+zkoymy
QU/X3ZeF10ZdvFfvF+hoz4ff8VNmhBtQMdHZVb+ZHw1LPzu3Pfc+sXIyKywlwnKTqoJG/bJLC5Vg
m+Agqp1HGmeNuDFYe0aSMYrSbipWdLe4EfyZ5kuU+auCAs4+XZgQJziEYKzM0bmmUGBkSLg6xk7j
/cUDJ8hNEpMluTkjUGFKCg4rK6m1zN4ZgYJ3/FYUDIcKmtFQz4EjxJ92fZxWvqf7JEFPTuumpcFt
MVbeqmHwg3FqIBeCPtx1qUp2m+mtwyFCBbGgvYdVONdtxYF7GbzEaoE9+sDTLXwUjElHN6kBpEIX
L7aMPkJrPNKAEfzUvw8+9e3ixTI7ak059x9NopEPKH4jSJNDA6+5riUs8JnTOKBWM7AgBOmszv7H
CvwQUO9YxJc+3WLYxMyv419DUqFlsJ/GYn4DC4HvKodAtvUBnedpJf463idxzclGaZURgA+bfM+b
TmgZNkDvYzXxdV7HkpQyIwBan444UI822vFIHoz6TRBpkvCJ7lWbmO6A7WnMBJt0N++ht+jLVnKD
tWHsRG+QpSQMRaqqDl00ECvGpo3iJdZ5pr1qke9iYiU8BQJdKn5ETGcc9r1lnm6v8DNLuBjJAHpF
f27SrOYKxjIINsVP3Uxse/CNY3964/lmgZaN24J7l1R0822xWtG1jayyYEPzYsq9OwrM+cobggWN
8hZzsVYVnX+SAuwySnD2A5WVpsj8xxf4SdzscQuhGyIZCzbHToxFpKloH1CqGKsXX/5ddonpYLm2
g6s3jY2rzR1+ir7T7jL9AHAlkyQlj2Q/UAdaqNC8xhPdGotvAbVkCm6s9piUzYteW3nuPwvZM8hj
Xhd6vSSIFIzyQBDzBiH+mmOlGnue8/HMBWALbdDMCq3M6HOI5WGc9drS/NYJmsCbvweAUK6+5jju
RiQSEyw1sbWX8dr+netTrVDajcXfsWpyVmiyF9AdiXofG7bJzSEAjfImSV0RflLzzdgPnuRDX2XR
Nvt84DycycYXLLDoBn48TbV0KCVHOxR43u3mifD8104bwrEv1vmboYGuSpRCZTDnlju8FKFhlfgs
O/gG60qaggTcDvaKOCwriVPQTm4AyDaGyUeKcJ71PyvWdZ7quuE8VZM1MTAIMyFnu9Y0CRsS442R
VmvMLmh/Vp9hYwUM/rTp0BKqjpcEEelAFeX9wIzzPtBZIA9ZUXLeDaS8BQUodkcc5Zl1jVZpeGVo
+hJNRYzsYib0uV10ShzIz1OCYtfkvsvlH11YO5Ujw9EC//KJUb88h0Vp7Ah0v4PyQTssNQ53hnLf
60PpJsydNn4mRmwwteLLZtq0p5iXB4TLODC/JGNYUWr3BF/kaBU1o/E9JHOQKFVDms7WIhONKrH2
e0ntyTj6TyaDksVbOyPFQZQOh0gQO537V6qt6KT2Bw55KRf0o1Zaepjw8cjynj8dzxmOQ0DERAGH
xFJvbOwYbaEbTiiS4nbjav2x3ho/3KpdlDw1fIF7By9VHi2iMvzmv0l2/JiK+QG6AvvJeW3pSkN0
4Yp720jsRcU4+K6F3G0nwia1OugfN0lt8iud1dj4ChL2Nl2Ccq2tN0CJBCMwkCIWkdeDTJpel8r0
75pKoKgNOti6r5xPuBPACt4wbWac8vcXX8esmFqhg0Y7KQyYY9f8au1bAsCbh7PvJQCkZof6ahMz
/E1nR38KHhY404fp+gSdyhoECtSPFA+Sa+oFoOme48gQn+qw6DLApp8G5b1g/ucrV+nwLz7QAzV1
eoOnTChRE96MdrG1VeRuqfgg/OGfaPohX3fh8UYHh+c065epIG5PlXb9D+t8WbN9zrjr/yN9L+mb
SSfNdyLXWrmVbgZbwaAIgzn9HYZbR2w25bPw+RLp8UzAuSlFYFLD3zU5ehTr7tKLu9ckpx3vRIWx
B6Wcc5hnPxq7O6Dz+0u11z6nVdonTqTZFtZGccmdTwo5q2tEtoPrMklJs8R3aixlEYXjkXfjTHx1
/hoSLtj7GQEOfHXF+3jtyh5zs6Jovkcm89zjPjJH861Ulq+BZjlZDlX8Dn4W/zSqLgl4nqNxy0oi
cUgkrSFQORi523/90x0lObIvazwjGCWR5LwJPkNX9zl9wbu1Om+NE9JYxr2yxs62uafS8hsbNu9f
ZOI7AmwsrGR3MovdGYcKiMpkElMsrhwN2Ak4PoyovZfMJjgxJRwgluJw6ZCAgbk+GEvNYlvuzP9e
5WovNKFVlRDwli0kbHxYGQtajEU8EFRscOQ55i7F7ltNen4EDJSiwTNWUjoCOshw2exv2DcEMfBV
GZ2nE/kD6sXXXboq0yOHZ72u+rpmmyVTYIkeCFnMS/D/4LziithY9jxsTwWHP/KcKC5uT0w3bZ6d
Wi04AwLjdrOmgOqpYRpnPjaE0sibgGaurVMOdVZNJRH/UKbDSw9Ci843IZ2iuLDgSXToO8dGnLvp
GuwdWrMFQGQMPcS/4SglcKmibJXcmCdJdiPx4wJ6EUcZnpJu9jFOgIR0lvL1BR02rYMMFvatO+BE
QIXK+RCvgRo2IYJpXUARZbpt5HygsXjHSIBVhi/4zTBg6tViZzWj+vKhcMpsyXaTta0P8RtApuix
5zLyL/rNvIJuF09CvMW9PC0ear0VABYU2h3uBtCyGt90m4JCEVO9gRS8EDmbx/zpQ/bwjDPhEw/8
d8H7l+C/csChSAOjdDs3ypEBwqEg+O+9V7trfkudTNBel9pmHEI2lE3hkU0t+hyiCJQHWz4avEXx
kwdOKti1LmEiXWizX4v/wpZqrtcCgTdJyVpWO5CRgknM8k956rWcODgwQWadRnGl7eKX2kGgmAxk
dLyJTNf5w47jsmQzoDIGeJhMZouhZm2zB5bcQBMCUwFwNjr8J1dRvCM/49E+X129qmXTfcf1gZir
G7ZaWEo7jFRinrewpo4bEogrLxdIf7GxKxXzh0ZwdeegS8lhsA4tYxeWFTfh7Ql++m3wTktnJoQA
pa0TmFzMr8ZXE+cHfWHzhdLHNbrrGRnWLJxZCzk6ia7eXXpUJaf26axWuxoHOdyW/lr1IoRHSuN5
1aI215dQKIEd4hrRZrr1rmQhbQUE7qMcbWfCDdUIHBl/JbLeO4LlilL/6S9aSC5MMh3wz5uJ3EUf
GPteBOY2ucu/bBAGKdLiAR6w47i2flSwdOJRANpCr8UU0xH/8jhz4HtvmGiSO2V7u9n4yoDHtoTb
jAMttK7H9olEulnBGSoGz2jVV8bwG7MRfOkNe2Fs8f1Oo4Fdgi5Z3Lc6vkOV+DDt1O0516EM7JH0
YCOW0rtR9fTOO6J28vnu3FelPJVR3Q3vgBbpbSkfOKhcHWhjD7DteeEkTsFOywoEQT91Epy2JzKk
juSMlKf5efioBAFjrYkRIO376F+DDkHN+oy0BiPMZnFOzrsQNAHlSSXURkqom/kReeiwxm8kwczq
QuYEN5Yg7iv+St5dWo2pLfEqIHOJsMSqnN+BTPhzJ+MCQwT8fK1Nm6oT9t4gAWWuExXeAwRKagrh
7HKqKCA1WkGV306FNdW5so52i+KejtGr2w+HnrJ2UIwrsTb0HTIqC/XjJg2cepuSTyiIgHmdtUY0
PBM5+lpxGUFrSCGWjJ79Rl/gpodh5CJcVSjbi9Dihkq1M/kt82JPeZRXuH85+hTiOSd9TEo0O/I7
iC0p+XZp4snQNWUr9jzMZKvwB+Xj1z4apPAM+wE3juaA+5o5lzzDkjkRb0qev/WlutiLFJHLdcPH
YktzWMk98TudLIMZjbKrSwGDunuOqs1i6QS6q2uRwu8hVTpr3CvsDPjerXEt5q637VmfQd2v9Yt2
lqQiiKuj2miCjG62tDbl9GQbwZHX0FAxLL6EQoLvzjskBrv2DjsOU65I1dx+NI8vrzlq/7nVHLZ4
Hx7Annq0GSjmsi9KSEps0pMDBc03WUbOelu2AUR1hqUZdCN/2gYpw85rib1wFoCl+7hcMmZwfavi
oemWjL//8F9kAokhCuWaoG276HujvW5rorUfeGMCJilQje50/EBKUu14Bz8ajEltVO+cECRe8yta
LM4z+6mDbSa/gyGpNnzO6DcDsFiD4oJU0mqF9MoMQloKejs1sCMlLNk2wPpnBmK1fg+EP0aV0WXJ
0Va8yC+YV1hv5TV3BmZ3JZxP71sWPrL8rogrIfqv9ucCPGcsaitBTiyn6ezukoNeYeow35X4Q6zK
cBSKw7F03zt41LX+uUdiQ2/76fkY8ZQL+f6wLtBTw6w9uy4hSAGPRsXCmztRJ244wwyiJ1KNjrHv
yMq+v1oErupP+D+5w/tYn97Kl1UZgK4CncAyiWmjPmMBBbEf5dvglkRSmk/TNmoohcX5f39tHtiV
InUtnNB1eQSIoCnK+RepegOmSEH3Rund0bDGrYPHOTiouubrrTcLIFecECUD/JZi22wDJFUhwHmc
/H6+6I/+2ThLBkPbsSeZc9Ic4kGqFBc0gEaVYzPS+wk65xXkSqMpf0rOiOZFm2cJx4EbnFtNyjza
41IP1Yxj+ox6AiH0G/81Rkzm6noz1dxGsaGCCgwKpSSs8Pe+gXs64sW5wnBh/uPDLd2BRPW5Up2w
pKLjTzQu+Jrd2Y3JT3SviCUlRnUVthl3/GocYnF64CK5/FKUNLO03/CGhNGctDZ3y71U7qevg5uj
j0+mrIqnF9vjOUvPxztel6c6kdI5QQB/dl7pD9Lp8mHKgVE9JJGzwZ+h7GGn6BMPFgrQV9QCSf8R
fPTXyrHx1KDu1L5wGnHZP/l10UwYUitntqJJ3eMJ5P92Uczl3XM8WePAkqLmYDG+Qe1p+xM9/igT
yLWgv2rpIIsOMoGaRcgblWbuNGIdv3uf2PPOjFCHL716H/1mVJaMtNIKGTlMHhTiApddm7/8AR8P
p46FfK+695qFKqt+0LeAe8tFL5oVdftjPtecZF4w3EG9zXMVQqsBwuYQgwadWXVEKjx4qmahmJAo
LWfbGupnGoGCp7ztJ3EmhNU2pfABvEh/QFANsI3ac7E3RDsFFmcb99OowdJPkNU4CV/PddBjzFL7
2mZJG4WfHlXBs9I46f46vkWaarzTtKBw9I3qpIe9NnNRGe27Hmnpfz0a2a8B+vinDhSFkPO1igJm
PAvwKrV3O/y7sxAMEXDvrio+fULKYpO+s1/hJzT6T6ptxCcVpnKx++F4ihIRGqHQrtVBj6t8kzDW
/3h/JbXFn/iXh4YJlH11+PGWqPX3df9BWaUlJxuPvXPyuzrtJ1wGJbw9pFNdnFiJs3fK828Pxmjy
cKTNG9gbjCTMvK6O9/ivQGC/MtsJNGngr9Dlxy9Wxv5WMtSxYp4iLbBPgqV2Pk/Z/MP/ikhUXRuP
xgQHRvpf8B2DBcVgkd0er/EYU3j0BW7mNWM7Lf699aNZxQijjrsJu3ybeInBeUQbk1EyTFj1Uom0
lfyf0fTy3ymDuPcVtBXSTJDa/LlA/3GC7qGPltf4pryVh/7C6U2Bmv98Q7s3ZlRjV9f3zg7vpazx
TUe7E/dZ+W0IBvq8AhhrkNRsupa+cOKxdZqZx9m+1FY48g+SffZzFDfhK49f/mBYR5f9UhcAG1+S
l574ad4AT/FqZbcLU/onA33f02pX0btSwUfNWUeCuRHP2bBDZqL5QL0424R8VP8BEYoyeinOCzYj
RueIdgc+q1SljF9FV/rRiRg8gFwko1VLVBWsXv8FNaJJ3b+ltRR/8zPx8TwrA5synIZRi8mmGLw6
INKJTFGFXteYwImLvAmdq7ZICVJfJzajuZObvB0sklZ5JOJN1rTs2CxiFMBebIAsXD1XJgSeXA6j
jN3FHQXLawKTKB2ABGL4TAviXuqYTd12qkA92ARJLBwT0sn/bDqHFHZNrdysEzGTff1jHLnj88Io
VLC0WsM4EqJhWPAFvvfIFOgeasUOKDNjLL8vTbshnVF/n7ZD1J9Kdwp37ZkuLs9L46Rdi37Y95NW
8MbpdJtDI3ktYDJiS+Wk4ZRO/6zhMKeEEuEb/Mdsz3NWBmKFfpLUKG+Pskf8tPzfALMsZUV/mm41
hap/JXEyGPtNl7Tmw5nAfQE4XQkfq3Lpok1DEOp5tOE+uJJom57Zq8N24/6NhR0NrCCzx9r/D5ub
Sfb6Qw4gMwnjuvi1hXey2ngcsDCx2Ljw9gMfFZPxstCYHBD3FT3pRzQw5e9QkUh63/4ZwRGBJs7H
hAquIfBkSgqpvyPvOuqY+vrUNK+elehiRLHADNCHfWLv9IWGDfH8/+ZhirUTNpmzilx934GXkWI+
HMaEEr8TdDp2mQzaFAHrNYeAZwFTZdnVSVdWcV+doYX1K4VAx4KqPYeSe2sekqRjrOr01JgjKkoj
/1z4uLeCjs4uyd5tmza+MMS1fQ5+1JvLSnFTCnwyz8afNdAA0+8hHcimxulZEILSxR4aDzFvcKxD
RVp1R6+Qn9cJb++hzcYUvLkcJFv9kIuGwBglwhaP/lS8h0771uuDiu48JIWlYURsuj6dMsuYgUEE
CVdamgNTShKrfo0f5O+EfBAkT64kBg9QtIMWnFZUYz5fUJ2thI2jyOJ/EcMkLTmbHiPrOS/hYFPo
9Rtk9xbVaEZjr5u36oGICCkfK4KrSdJ/lgsJUnYJV6WmvNjuHwZYsKA6VeBF6CG6KjBoj8nMq9jX
xlsgDwJOYYk9d+MHFXkhnvx5AGsfGnLaMcPeW0gCjJiJP/7NcUWXwR9x1LJxmbrzEVnisriNyzDa
1THzOZRu06VuvvkVsvlw0tkm8DkFIbq9g4UNTLI6O5BryL+rXaCetrFBp0cDZGKoxNls94hYJMIl
rwawBaw0QVRrN8+m2PG/8P4c2pvJkOmQ4bgtseSIZ9RnrNNEMbCqNtLW69XkUMdbLxoLriNAreaJ
KWP4YjfnfeCcVK242Y7pok5/QvVj9e5hGNvU+hkVNvRdSXosx2g9iDMBkusKfVkroCDwaejblm/r
ngkVpiEV8UrkpVUag7bZW0XOzsiu9cx0IejHbpfSHZZBgdR00JCDP5gH1vb7TuE/8VQa1F/2VVVH
rk9gTtoFE6FswXA/Y5HhSu1mBCMC2SORVi6U16toG4uVht+U+j/ZXU5syZ6b4ucdPdFT6td1NU6z
zLiq0UOokQ42MG08JZUn49Whzo19IyIGjBv+6hn2TTOyIZ66QdpCXXyNxv8r8KST1OP+DKhYuUvU
0WmlE+N3KkETGZGFXEHHv6aMiOmHewT0HypFZJkPfDyUm+o6dzr34ngI1Y/7AHG0NLiiGg6VL56u
S5HuE+cPPGCtvDLpC8gBiB3e10EeAlq/zZG4jkrO4p3gzFczBpUrzz1r1zM4JN+PmNQcsG61swhQ
8oRPSg5yPUCDu29bR80SXGaFnjlq8TyG54nqJZO2mzcfGTe1u8Lb749+aV5aJ9IOTK88KfwKOaLL
euUvFCvWHlvOAsR/q5ghK3BLPUGCrYNlx+HIic5ebzd37p0GAPDw+Ofd4NkSVqqjHhu/RGK27GQp
/yX/KvsgjNG7ACG9TjklSpd0MCd9LSFd3a6VDvtYDPiaZLd8Wxv4b4akS9j0Wk8Zs1n2qUWZmbU1
W6E6gZWJ03DyIE4mf+W8194b8qoXCC/JeAIlEcorHpooAeHSrib1Jpb24UcQHzYCe6s33cBo163c
fRIZJeFs4yymrlyUGUGfKndxeOVLvtJlSHQbf9a4fBBtm3JmWPer3hZe2zq2v+jINKqpLuWuq0In
LlvaomENL7Q4gSQJmOTTAls3MVDqGpVmz4h57/0w5au+0XCtROOkpHuwYHoVsy68zqKUehBk5O5C
sjBwu3/XHrI6p9Fvo1M7NGC1nbZQC++vIawxbIaFG0jS6bDcwiV7EgVVD0eAXpk6aaEn9IjdDt1O
g9M1AXKaGv+y2Y1kdAPpxPKPMhK/OG4C76W2O4GyPBIz5G/UPRnzyZjVpDqI9uWibd6V2XkRgm4C
nrcc9nPQDAPcWoJMNwq1n9ybRYuqxYRY16nu6EbZhTs7DizGQxaMzmOrVtwacejfznGS9q/DNWMP
G5pNLfyCBnJy6DVdzdkd81p8cL+RgxBmudi2ft9UHVq8sIlBFN6CTVwUs0zWmeW43eAH1UPE2u0T
OA8g6xVX9HtIoXAanxVu773WtzyREPVFYH3O6K83ROVSin0XG0KwN8Bh5zbCfv3P2hCLrtwOEeez
u9Cu1QYFNKtYwyVhhtasEYLyITZelCNj0RHohWLEQAgfY1IBoRYixSGoF5f65FpoXnFHVSsXrPEA
h5/dlkgtdjbzYZ2WOwU/2hoHfAwV0kbGhgdzMN/PYg+UnvYHFMzpIULttBDxIR2eZsLvBHq4oHVv
0bWm5BgrrGc+qjCHJ05HV3simkQVK/FsSfbbBiHiCEfxGeLttqymTMo25IgUvUSN9vYiV7hazSWx
BtVFWfxmV2LcREMoNZ28vmj4x26oznA2ZUk0y/O7+rAK3+R52MIyQ/seOFCeAvzMBbzsD02xEx9s
R+4PDKLWqxQzhtMZAiglpuZN+KDqLgOGW4e+K6JZMOFYFAKBXkj+tMrUEIr2QxAnZ81zoInzR+Y2
mKGnne6HdBbmjnGFyKTygdwBRvx1JCn/RFIPwsaRXGD7K0Y8J7eqauaOEeT6Qnss26gWt2dLeRK7
KBed5Ly5luBAH37Pk0lAyeLyLHtcxrpkAkRsPHOSxbxb6FTpeUIBFUO3fHaROv90fp44D7f3E3wu
jIqBJ5ZMSaN7w0sN/XpNPDpSHkjeVSgVzOD7fKQBdYIFgZy0kBwmDfvA1f/s9Qqo93tCX8Sfpifv
4wr8gvBXQ542qybhoK2TnMrLAXOn6Gn4Dei6e8jADbeES3FmqLZNohq3lHrzGwFOfEO6WT2VLFEf
XJLg+l2OKTGXFgVkTlCNcNw2Vma0H4DGdzSPh+AyX3SlU9ideIzU1VQoghcD1z/F6fdok9q2gWAS
LUQZaXZJ3XKzYC3d38qnvP6DArkIp6gIqIdwn+9pkcfCf5hKJ9bHrQaN6ZOS+4CfzCmZ2zju24dW
9j+e/XuY8L2hxYt/AnhsPLC0QA5vRpD8UAWF0W4BYWBG+ZWR9rWMQwflbuOnSKRzGlvQfQ0V5fJG
Dt7I1v6wfyel5+EzJenGhaq+idXPJqg46fVsWVi6qFe0DCcNK9Ioo40QtSjMaTz+RL0nUfe1SyD2
GeUlL+bczPgEEiL+0CDctaUs73SkS5BpVFkYNoicj1kvFdz+bz5kojZ8/ezFk8aM8AGrE6lmdWX9
PaVvTBJQ2WPPx3S83TgomGv/OV2zC5HFNt3g9qWzBrM4DrDvpyOYPNLXMv2bqEFz8m/YAQlgK0ez
muTfCLmJ+uV1XHrmbYuviTp3GjWchGDvpSpJBP1n1WETz13wnmO+M/OhX6mEn7Rk+oCkUQrtJZbo
vgoZE3jtwakXgd9VNAU7ca/h4RKuEudfJQhiSA/Z0EZilu8aP57ynPHbBoGpemIFIAj+GKXgHdgB
JgYpIG7A5eDPkbcKbD3/+brpCFCBx/YoS3spkDgxyruZHfrL1FHNjGx2Ci5BcMohQU8hAogOMIKE
/GHTVJQC8OskxDcOAnREYajPsUKyxkul5K1ogiE01Fx3r8AqPmZOUfVkjr0p8lMWxhqzpxF60ZQ7
FUbgHwXjeukas5D2xHkM/jWtYHjKKdwIRgFFDURM00fYTJOamaVOkGZl49wWRtu4B9aS2ZHlx//z
i1zvhpqo4j8FVwj+jE/jqPs2Zw8IWT6eAQkWafYEsIFwiHG/Lr/F2DSQ79LDyAsZLkqOOEYhOdDs
6mLVEOSyvHKvvn+GqtpH6dL10/57133xKuxqvaRzkZLCTknaKAzDQyGVjzxvAeOlaLyyJ+81wcsw
2Zs3jIgO/pwS2MVXkhIBrcc6eYoniDtJInz1TzeYdQInwy2orBeKbb5rCIUlNhMZz5NYeHz539+F
XUbgDrzOAHX7H9aui9wiP9zrWC49Bi09WBLYpzzRCeOdiCx8/B0PvN4KEQ9PKlqHVu5G9i6ZxRhC
wuPWE+VSsgIVDRBavdvCQ/FrGwv7dDSvJe5GYzCaMQUvOLc09Xlu/dsC7Vn+wr8ZGziiZKuKTCQD
sviVuvUqdtlEUJbou1TYtubbH+2n9gb/5Q+USth8bxasGUTri91toHZ6ztFU0krnQLRrQt3oyTO0
x082u56TE1OI9Xto7UFJ1R/GK5+twhKGq8eWF+Wi45AY9xhbjxBsg1tdxjg3rL+gWkdoZ4qpHu9E
uaQfUrsdZXcGDAkVJVmnb+CNgamsSh3tH/1a2tbGlMCZ/IKORxLG7EctJhj/pUKm7xSe+XAWJ9oL
CGJ+Or6FdU5njNodFk1dd46LmjeaNYKMUuoCnGjtWxmJxbJ4Ll9MlVfsV4LzGRNZrWWJ2tpBK7zL
dBQ4WiB3M383NRG9fLH2inXUrZwygaR/a2kqM7BKyNGFXpO5oehnBcgiSm3yvT2/aT1oBWS3YJVq
PSLpBOuZfU/TJLxUPaOU46F8FqK19TF+CVY4QVhyzbUStjqisHloV+zu4p+H9w15ybaoe8IDGh/E
l75YvtftUCtsR/XNOWpfWe2+1rpoTXxRaGFtbQgxI+vUb95u5/6x2hOUoUwiEEGotCJPjuH0JuNW
EGeNMu3stm02IvAf6/hzA8xVtPhNvTQ3f0gEqVof5mCvRh2kWAURMEPKxFu9xybXjcxP2j74Tvl6
vRex2jcy545xUsJO5fjJYq6V8TAt/u77bWTp4boZCtWLkmkBFIf+vJSqYm43gE5r1gHKYTfJJyDr
TJAI5g++xVBndQd5CM79SxX7hHz46MjrlJ3Vevpfz13xs5BvX85vwsyzXjgRgo037go/Okj3Jog9
1BwcamZdF6BLzU/49dEGJkr/dle4U9gV5TuKUS0DqNSEgTrOgF1WWwD/tlCBjLqEVm69PzK8WODR
avwIQXNTsye6Y4/4iCSVLy82lCf1FCHOd3jB1p/fkPT3TK5kLgekvR+AJdqnWKXbF4I0iTaLDVHV
4ORd8Ikay5SVqg8oudBGNP0ecydkjLAncKqxT65+dJpWLla9AMZzhvA0JqqbNyDD8FTN1JScVUuQ
gsoc4TWCcZIfc6uIreGn1pd8v4eZqcfkL4QoSTdfdsExKVF1eq21SB/xwrqivJv95oE6djs4ykLj
D+xJ6cNjw8BtTbUfw3R/GGhJ7q6WqRfKGrn3C2CwOOCyxDx9slLbWfBVMw2KvJbFLda7XCzI1e4A
CLyzcyTcJJ3jLufMM8uCetJiEiwr4Df7Bb5sArRW5nTs/VrhARjL7du3b9QZh3PVE315D8KEu2U1
fXwyTMkpyw0njiteyfR7t88RDuIxPlRUlDb/AuZYTIPXg850cgzN6Ac8V0UuwWiEW63qmDK7BVqE
K+0ESmkd6EIe9ZLa0Kp1P3j/Dlr4RFQw2aZNx0EJyzisoc23IkvZ0+EpNaat4GbcaBZWSi+HTRcW
62j7hHCn1KPZrgx2Mjx0qr9E9A70CD8NwlwG1QhODpwDCLx7/pw2zOw21dwFV9U94+2yRQ2ofzNW
YdX7n0HjrH8cW5csYp7mfNRi23P2lamUniE3GpNU3RvgZKaK8p/fmhdJ4OafYzNhoMmE35Yulai8
4Jpv3xYvuZq5SFfncwpt4zM8gGvosUIqMOsZbok1fa7dGlV6GWE02Dn68HQU+OgZMd6cTDkXXZNZ
2HJsi7bBFBnLO9i5pizE4W46l+DfXhRU1Gf4PkRo2TUfUGYB+y1ARqU70Jc/ni2jgQQ4ML76RAj4
3WzGs/YBGrVFaWVvKjVxxlJsgQH534DZ3Tiyer8IX8MjvQ+zK3xOaY5oJreiVnN9pMLw32AQg7RQ
GFcMTk2j4bfnHVlGzWkbV0mhp05+ILsk9P0Kgsmo2RJkgMFAHVvTt8Sou3L4ixdsQNv5fTaPvwf/
fE9LRbIgr0ahL6FFlfq+6uTTm6lyoQZqdgFFus6kq1lrGIyQhMmS+zD7xvZyBdWaay9AEGXJExki
NLVfYGw9VdrGCHqzWBx9ziq4WvoS7I7xtq+oBVR1+3BVcO1pLpsewr4h8lVkkEbbqJt3Dx2PpNz5
fMVKTNRbqDi2c3DaU/ih0UH/BXl5F3t4ilpQzXJM0OEnaLziBvhm6gYnTPKGclJK3AsCwbdWJrio
5R61RjDgnqelB5C8+Ri8agxmp0Blrzx4ofk+c+iYjggvQofreHq/z5Ou1qjdwk9pntBJ2LbowzxN
8jz6iC394AOt7FLkekxls12lGhyewAqr9JKDOtUY3eYtHj3LAc3BMWNzPuHMb9ZkCjvPsM62irZR
kMZlBY3B4CdON3POCcdva+asx0seXNIVuWWeVMWRjOs/KHpZOaxsa2y6aqZoPcpoCJHNnba2Zps2
DrvnSibtbmdfGkLmIp/XCxVss7hZUD29+5yL3yljjN203Le1DLuMnjyUYbIXpmBjtnJyJOuKnQ/I
NHPtWlWqhT/KBjUn/b5Ix/zGXMR5aZ3CUphyvFIE1Zqp3+vAKrzbjsidelRfnAM3BG9Ok3PVI2s/
rr5lczw5ialR11qEvsMYt+BKt7Isb431iPAKQYCc4z0PGUBtkOMkudgsjECpiGhaCBh5TqN0tBce
qtx104EKNI8kzkYrdBYlr5UDyX7Y6cCRFhNg7xlKoMuz9ArcoKtJg91zXsP2gtQ5jAtkz4Ak3WN+
WAs/si9CUHx28Ksi2TSOKgyRmy1vmgplv3DyH08jWNjd28c9meCjZtAD3nla6t5mhB4lgb9AoB36
oHU6R6b4DAPACC9OcHmq8hahleUSYqsf0ylEapxTx+5zfbxGGpTvO9caZHyBJqTy6KUtrLNhg7sM
uosIWAOlEfh4wIfSw7NH3QNcMufO2LhttY+Jxr9N2KfeVp45OVNqcEkG7w+4ydJpSGjtNnmRmlJN
BlJs0iSuwPMFAxsAYsRSlXb5UacYXtfDzb8sUYIPChaFtY+1MowaCHm83s76CbtJrijV9H8RP7B1
D0zgi4OxqLd4TPdxMJVF/dszY1j+6GgMbMvNAjgPAWEqnRvxHcYKGZHVZo6+O+BNb76WNYb53Jap
+M1o6yrkWIvxj8GxrXNBKigNg+LMNtfp9h+E3MDbbe3jt/a3AV5MkanVXw2Fam0V0O3W1WYcPPmi
MeVk0MMI5tPyjMlpLSesK5+rZcUJP6WXwGIzNY3YUFd2qXNd0cU9Ga5nbs6/rU7Vlv+61Mb96PGs
PCj7Z8y+b+v00T0c3eDzKS+n4oCE7RMHVkotaQncjOSzlijK88CaKq4c4Nlqc5gTMP6QmlGdnNx7
0zZtLjB7sO3qlCLJ5OU5PTb3lgKQpt+N9RuQ9jKz73l/7iiWodWe0+vuWiyzzqq5bMC6pzEt8KTR
vcEEpdoI6Lo2vpM66ne0Zaev/O1yx+f3Qnen8TNvuVcUi0vt750puaPLT2oOleaOC0973SeDYLeG
MqrqgeRtDV3Fuqd/NKVhb4BGCii38oRctXbObcXc1TzVrvyqa6uEpbuB7LmLEzbdHXuVyAMHd6cI
L+nW2kzmSh+HBla4Q0eumzTJwttz6KJLDvjb5g2TmPJSYTSR8TsvfVbBK5tnRkWGUP142ih8rQPo
q//Hg36oHoJtNS+3iaV45mWZWaM5jCE2X1CjJom7jPw0KsITQ7403eLNIEi/wJmo2CYedxXjGWKT
+4YFtSMKQM15CAy8q0yrJaYQr1V4mRKW69DVDjsN3XbN4uhxj8luTWPIDNxixt0IW6FhqEJrXL/P
IxWpFJGYgwEc/95NRxaTituuWx2fVw+Afcs9v6eOfjY1It7i9qaeBXnaXrPWiti2uW+jSr0/lzRj
NLOKWVtFEtqKjbR+Zaxyc6WqMn9732N3ulVr1Ayf//WbnuCWu6T7lzWgme9QGZs0Rr+J3CsXZln+
oZlmKsMK0MqfNy5QsXvKbtOpg2leHZhgFIfKXyfwP+3CidVEO3IlarMOTCzk4f0l4TcwK0uZal/f
nD0muIZHAW/3cb1sAT6R9TVLUzKdVAKfet6iO47YwWg+xm131gY86AiTNfxR/Gn4mZ5/7VEOsnqJ
8KEXT2vBtZqM7gtkM0JynEliIchPtSWVafHn1JbQD0lfs3KFgIEuE6O21yEszYfCyDrw/QFLRJQP
azgy+Z5Ki7UTlmt1g3UkJGkEuqrsdJbcx9pXXNt7nfWqFtxlng98Zc8jqoSZOZTqO8VkGIgbnkXu
3XxuvOGH20vmjwumPpToxAdTZT8DEXrnazb9abrPWaJg6ExHUj5CD9Vdhqe7kz7qu3LOXn/4mpFu
PuM39Z+uRxaXFm9dyL6w3vH8/dyh+lYt/GPz4xTH4XrMgkomdT9OUzOqCh8+vUsgOVYmWULu5c6i
XHrcusgbiZCAtmrERosIZdpPgZpHToDj36Tai8Gs67W9POEp2jJmI/ZVi3rATxNdVg6TsnU+PuxV
XidNhUIeiTU2EtBhTXQiprNzWvOaC20UB9qpl1fH9rQPu9wRF8jzrX9NkgxMnp+hNl9wdSDETzo+
69clhkAbzuIZhk14db7qFW1Is9ps9ggLMCtKD3qaHRjK7aUfBaGvytYOKfYMLy2Z4FcJ32N99fqT
ZS2ZQNrzLSfILgtp3ZCWbr4HDOFSSUHm1SH/RK7+uLurQwlXEA1q648I04pmDEeAuN9UKArzhgwh
tyCPJtxLu4B/7qWLSpd/BRMr9VgcPiKMVTSiK1PL8Lye0Hd3VB+++hJVjZ6DXVXufoqAjCnakDR6
QBZjegQ/dOTw2qzQEoa9bAr+ZzqdSjMddX3ykXGkex6I8lWvm/k0Kn3JNwKIs0greFMiRdXpLA+i
DpZnxiRs9Cjc8tla7n13wZoRZaQnr1rE54cXL6VVlomxHw0ndje1J4/XwX+4tedfiooE5DERNcW3
TsrNiiBqeZZpy56OkmA93cKCYuZBNZ5tEgg15DW55B2hdK2p7nhGYuowzPtVaSj6kvQ+ga3lOzL2
xHvS2v37ZLvPCBeaQZ8xBWdZBTrjdEwxqzD0LqwMduz5z/xl+AOXQCDbVDs2fTml/uVoj5zIrezg
o1lWz1I9yGnrXqycLRV/DXH8K5RTkmastblDfutmoHT77r4rjSymDFs3M/QHAckPBakdf6eoVHnG
iC6QG/veEQGyI52vc0I9RJOy5dIger7z7qS0acCvedRY/lFBVTKJfzk5fT6+Lfal1Jf1kjOis16b
JwfH2/WIfrZ5bHhZRqEdmdMyirI+06/jnincb/6L8eERxpgVqEg6Hw02l2WNa2KyERcAqiH0UyYl
xNxo2bbJVLhT/gniXqaSXfZTezHrrO3nZ5RQL2LBTA4ePlnbXSUCs8DT0yq20asqIX+e6Juis66P
xHJg+79yjvoibX9BNp8Oc6OtZqRfNAbE1npQN5AhJsa+25aJezopxbm2c1/cKYUjXQt1Dd/oHOrS
csPrRba3kn6RI4Znk+bZXI0Yfo3+gbpaPLmx7a9jXbli31RMTqyP8AB4+8/drS3wTc5eyQ+QvRmS
9wyVrLu4XJHEniM8chY0VvDOiDDnmF7UzkdT0qlEsDUCNSPSzR8tRkoDGcNgNIIQB5hlFGAtQU6a
1B2HpVGCRSJZi+wOqGOVaf+N6ujQ9xNuulZ25p+Hvn/3YpeOjRmSRw8Uk5zmuAHVULe6b+6ZtjEd
G+NoIzBdwszdzYsXU0LYX9gHOHknpm2VpbKgqT+iAeY3AlLTdUCPslrfcRXDLUi2bQSHwsY8Gyze
6MUCih0rQUK8DUotJDgk+LtGCV+sAMC5czW56/4B6oWiIj5riJKKMOpSn2XXQhcWmx/INedMwa/a
PHbcIv6ARnfgDeuCnxj3/UqEoUPo3mb5PaGsg3sVVTHDTWocVZ4dPQVcCjbJ1VpPe/0TGfGcl0Y6
BiRAzsxefjf30FY/ciflHWrE+3DlQ7UJDMgGVkAJ1R0pailT60Jwgr5q26d+8CxRG9+ajXF3HiH/
ivmJ95Z+0waDhYOJKCnGaCSafJ6gU0kWFAqjD00mZExJDsiTiNEU6yOSuKt49oc/jeTjjQ0UFWrW
jbDmRdTSzvgW74P2JyAClg3fWVPyHeLKecCqZtYVCCst3myPpEQgWDBeIVxjR5hvBukXYJ4ECStq
x2spWN7zlxIpGrEh6oC0DCdoejvCy4IyGkFOplycGy5M39G+O4UHwUSGJucnDQtHbN6v7FFwgODd
gp/o/njo5hAp0MXXw92vGGnbSCD6JTqOT3k2WrbB5KWpjW+2Ik//8tqNKcX23gKvM3n9cBvjxgSr
gXdHotuRNwbocaNCKxwaROle3Cfd2i/IMZfMOe4hzjHWmxhhYOuh6CyOLpLYForr6xNedXxR6c8l
5CF4sy9lWUXbM/nzJ/FaNZCF5RyaaPT14qKvxnkHQbMW+SZpJwdgawOkzUMRPpuuYhGh6gC6Jmil
sAL4IXva8Ggk9/Qf1Z5EdOFhylY9MCVBaVj6+ShBa7UZ9b5lX1hxWSuzvjC1uff/ZmHLMW1FSIAq
q+J+4ZhkN3Cv13Gjy9X45emBALWcbHbe6thkWU4lpwk0ufp+/au3rTs7JnA8wToxM1wD/mqOI3Xe
tzoogq2zrlw7CqcHDxGUq5FR2a8Tkf1vuuuJuU6CpXNnkdsybbR9bAf3tSLQMJ1Y9OUO73iK3tPQ
q8BXCJY6WnuBg0N96g1bopldhldY/A5Pvxxddz0/ISPxZsbKxJSWWm9OwfyNpiQHYp3pPonSAd9D
Na2+WZCdVX2lhhLFH6p7OUnIJV4DkI1jo5sdbCV6EC9Xgeb1MVrr72/lk7omzvLJkZFzCoYN2NdO
xCl3zq+g2mveHCu2qusz5fryh+X3EI6Yn1fIzHrwySgO47uTAAVFW7d6kBaOwL0Mcucc+er59qIR
8UHfOnwOHGZe24YtX39k757sETiH1+4UyOAZxhoBcwTcBz2pazP6z+uIE/HCrT2gfKn7+v7uH4E4
+TeRA9+mvpB8xn45/gV8XdfcgFulfb9J4hiDSGudt9bdTB/dEynK+04DZymrpbMJZmn5pgAyzwLk
EET639MdmE7uVNyEE7gdt5mSg4kY4N0GFTdLR4muw77BRZyTIecRC/Gru57tmMqwhVztZ/qvzRrE
OUmu1o6CTmVpuKX80wxx6QZU8W6rWc7cJ88zZDk7Rn0KcjuRijk/6gC+dN11hxs17H1/2WS0So+H
rE7C8nqQ3uc3RfSk8e//xQtIzipgdwsv5EHGgdX+nrHBZfv/BRUzCi1znIBsXFxToc9RevqKCKkQ
kEVnrUvSmBXtPjUK4agk+jGnpRWrUhgXlalw07MJyAVwIT0cFtQIOYxyT6FRTfav/zKpaRYzanpE
qxYA7chJFui6jiiCPodDSnAUiDlJr+ygEetmOLNCm6wF5J4v1bC7Skvv+H2lJNROkpHXGRifUKeZ
3wWeu84I2T0xrbMFsU/6KEOOkX7n21D/raoJ5NiluLCbawctlVzXf9wL8XoF3O4XHaH9Q0j0LJiw
EBru6GNVtCVhsDE0tL/KDvkHl3Qfeu1J8em4aEj44vT23TLFlIladfrdfGPsvoUnq1ranwqcucWz
rrfbk4VAO/PjshYkIlHpYgoLCKhzOVmB3mFQapvLst7PVQtsKqfbwhMaZvItiNL63e9HGtwt39m/
gR3okxCUxSTdnymglnw9pYfmXjpspqtUX5x6R4Sm+q2SIyrn2+Y4r2vK6vWHaoUKNKJsBZwrX3bE
BCDrB+Zrn7OBFwjMg6PwdFVij3VQAsBuAJz9KgBSiwXrfeGuHOmIUo1vQ8uVCxYMhvjGgENkexNo
R92I13pul49Lb9XrpPl7BQSrW/rwgI10WD7kUhQFLjD3S9cPrvLRRdhJ9zwFUm7wjsjJtGXG/oeg
oSBDIe6zNe29BC+NKMNH+uJx103H761azklA4+kjjfV3kzWgRj9EOjmshrP8p4SZF1G/wPPb5rIQ
3gKPo9hOvf5gQG3+cMEnoljRl+hNLTEYoS4u8IYMYEa6zI+j5UnBrm42XWXcjP8kTM57jvZz66sM
yiDzYm63amnl4wqmdaC0L8iWB+VkzpZt3fhHoH97xPiQbwDZBvMlrYltklfRKwMf6Hm2alE899XY
CmwUyubmAfM+RldxnZ+e1u5r+lwU/dXNu0b9FgcRX8+a4+F6rRjofNlLYIlFpUfUS0pQVsfy0EtC
N657IRzVT8boKojHz7LkmEIc10Ovdes/c6u+w77Z+Az717dk82u6IvSMR5lNxQvvbCQCVftWaFnh
ZARMOFTqB1XOSsy9a/dDoc23avzEs0AuQ61iyjlD8alZotr0leEavXCr2iAmrgJNYfVdukbl71l4
rcOtAFU3Is4pc56ys7slk9DWz2u2h/h5xQCPn380uwfAOPNqQJImLfvGAteElNKaeTAPdf1+zsWr
wD7HD4LGDBpql6y8Yyq3XH44DNTOlFPwsPkhF8eyhjCBmkmDL/yHxoF8NzW9oeRJFq51aUWSclLE
9hH+P5XC+LXmZke0w+AD09DWUIw0hAtnX2Pn7EN4UqOKuRHI/HY+iBvnqPFgDkYdXj5I4Cl5HrTf
2nkC/nin1d6xXjU/bCCTtPwMDworqlRhg4cUhqGmZ4l4mSSDIZcQuQvb0WCXM51jPo9C1L60pAwk
yrzgi8DWGg/iNnXBqVb6oolbXOAfYUCwr0I6uYBFBYXGbrscmHlyjtlvJdLvT8tLOyLkYvkEKRur
B/eTDgJdczgaSfpjiQ8/bDC/ceLC9yXgCSdBPUZWn4mxW3Gucy9rTVmgAu78fCBK3w1JrhLGwbgg
V6jcANg2Ovr4UHbt5PGBUXw0CrnQx2Gk5g/1PHQhPJeDg4bvOG7ZRifFeCSyjY/9yQhNjK1n7Hl0
rtX8CPSNiTMixZSGLx6XOpczhqxRUk3tuCidf8hrsMjuFLC0XruP9w9P8wBcxRKOdJTIX7Lc8P3K
j3a97G6GJkewd4YFgaMNEXASFMKZUJxXlc4d8gDU8u89b7G4YGA0q1AbS8FtZmUojVJjPS2VoKNV
Wkbl4zSjkGTSeDqrQbbJu6yDZx0+LNe/jbQ3Y2dJieuuZKY4KUof4VmkoLXRmP7qO4wYb5GLjFHg
eOnYC9jqGsrZb30O7WX5twv6rbKyTljmsZifxroNGeD5V5XhKg00PfV1FZhBxeU4LX06t3R2oex0
Khg06nrPKz2OecQvhgl/u42885NDhhKg6jX8jsxwYk3hXAk3uoMUpihUWbt8Vu7DG/oQ+0GwnCP0
MciI5udqrvn6ykzykwMMs9vjvG+mcdZ7JCW4f/ngqkgJHVoLrhOLyxXE4xrZus/nvL5WmIwKrwsB
pQSY6Ryc/m0BUy0McZD0QcwxZ4IvRnKyXK9nSguSWxkGQoFiEcVdWa26aWDkAGP1adfntfXgVDl0
UA3q3gd1AGN+Mgd2Gj/xp8cPdMPu/rHrXUXYCdBW4bAdjByGMq2OVUBtR8KHSO5dxCuiTTGyl1+x
qaNAZSiYQl2nMAeu5Tvy92iMGJHOzQxCLUe48Wi6UErCfHcjBJz3+ydroeeAW1t7OwD3LPwuzVD7
yoeKSWQTDMDmxz2OXqnFbRl9zEY8Yl+4VYOZZ+H2cKlnvei3xiarlm4HtvB7gDw0wk1NYdYMZ5Bf
dt1BRo93pqzpZSESJkACUOMr46UkJrVNmMWTWX64bYKgaPN4g8+pGDqZDq7XG8wIc5LKx81YS+t7
1o/sYJ07UInLgDiUZ4h8vipp6SOd3k7U7CQXbUk7/gqExtwfHtJhgRHrQMrIER6AfEnE3VBUGgoI
Y015T7ww569r92Q3wyoKUNjVoZrLCNvu/pwZuQRtDAqs+zvGkHBXNNI9SD0fsH55md08NTduKRIq
I3pHNg+SoOuh+W5y9qmhUaoZrn1tTxsjkOyLFBfhAiG/mmF1tsC9OGQ5Nx3uv3zIsLvrf1+9k8/E
J2RefbISzzcm4Ig+UlVkEGq+SxPJXDgmzZU7pP57bWRoLveNB9Dw+bxUps3dDYoEk8+l6+qv6png
b3H+i/eJKR+nnLpcY+cS1FSencQmIRo6gf39EmDBouDkrnR0XHN+pd7GI+62Jpe7kQpUSGMK+wzQ
B5qFQA5dKTlOVzJGna5H2Ovn542Vi4ZImZh3JBlo9qUIxFC0fePS1WjOAH62100yrYrFycOMYee0
6T+zJNh4zfqcMwfDmmXR0MhonwPc50/Vqobp1KdGHSA93fJYelFYAKBtGMDw8E4eBZXnomuHXfae
ozy2d4cHtfat0x2tpSIi3Z3rFeXLSkuVLWJrZXWq1v509nQVuqWYeQUIwbTsQJ4tWYKd/2F0X3q1
pRSswulHvO0MKfUPKGuraoU0lzn68LLMgsk5LuwZunljICK73XJzvOZzMlNCBzTfw5SzfvnKYpX2
zOOHVptH12i0jRkjI9rnkfWhNH675eq/E/A+yF7MiU00U/+GCeOICBH9Cx/bNK8K9ZxOIcUh7UpW
plZPH5333Jbap8I23bNyMgUWebDt56I5fNoTVr+7hHYEiEs5VfIB50YXmrtbkX+qQHnav0IKbtO1
70SfAtnH8M/H+j5LYkB7/F2PeD50BonOGCg5OEr5kW+O4YvuwvM2BQ6ReZ8LjdouhVmXxnS0psdN
LKt+8OB0hv+ZzMQtcG3HL+OvUyrOBuI3d70buS2JQjs1l7UQmWv3fpbW2nEY69aYmR+IEyICUdDx
/B6alFNWUZg3y/fe153EQ4BuhapozS8N7tRWNAlHgl9TJp9Y4Y/ZQ/S/29ANxixxK5yIulDsnVGn
7Fpyzq5fDOLrvRqLJMfrzGqUf2d0cotL1F2g9jzXZRsfQiNAOVhVl8PSaYTdL670NFjBLwYBw/ob
dWvGEyZu14+A1iqUjwnn81HAGm1Rbdf5KFISEih9H9ohZPjpt42tycmtnyp3C82B2nbwYdpswiDs
f/F7wl/FhNMM3CJKBahsALGWOcjLjULCkOIwfdIxXLEa4AwwuSgdLPWK/CHojVNVK0WN3sh0iJyt
vJh/Hj9R16AUoZYMX1S+QbnNN5CS68SBpesRxtQFE7cUVw8979/es4IaWimwB8E5ZFVhSioSOgi1
TE9eaVviwhu569dTci34HnZAAauLJ1KA1fkUkhsuSno53rqqrn4fUMoEGXDK9eQL1xpxFptDpvEV
O2XldFoh3Fw0FKyayuGJd2UZwkBOGiZI8mWFe7AIQKO7awX8a3N1MMf3EoicVRJCnFlZ7q4xgIbr
9WilNYe2cUj2KFwuVonNpdoxix6JQW106XS2WyeCfVTQ91+95DG1nW7O+uzqTZSwsGfIMsrtBpfS
PXxd8lFel11csWMfduK/D6Hwg90Q+SOCN/uxDWTR80UdHazbjFD6aDuYsuTE8AuDIyBaow0VnLNU
besmiEFGA7QmPaEXGiMajgFCdjVSevWa13KyTxg4y/wSA1ZbcK//G7IIaUt6lTzt7Ogyz1evDr3o
BwfxS2NwTfSPtXh22IXK1aHTBf1AeYwkIoTSoVF/CKdpXzcoTDRWs7AVAyZuAJpTySb7LRgr4jUC
uyk5VLLppp2m2qAOVofACDeX0snCHV8C27FHbcd7OnL2r1IplndBXdjjM3FS6qk82c3wF0CE0qoY
eLcc73wbfkvcgHvesC0ljfFjvFS64cV6aOY8wa9snDg7XDB5jw3MLr30glCvy0V+Z8aHcszXQ77o
TM4pxyCCy99JcePoRcoL+ljIAZ3KSQoWZ0LuFgD/STBRuoLNldKKbLkIcOW+zTssraBK9R5k2ceP
Us3/9/083Bp1cIRdQvwyhjdvRt9vo3y3e+US1RigXgp0am3VlcJwCmBoD+4lqL2jcFIz1oq4o9u9
38kM1AsoahUUrBepkbmFsrjqnzQDwl7hqvjZp9PKeo5SfeF5UsKPOYCEJbGMDosb77QcKHD6mF3q
Qv8g9aNFTW9NvMiSGxA9UrkJ4iyrWY5tVblO2EcmZHIBk64KP+ibZ7BL8l5qI99kB/FJs9MCIPCk
mTyh41JmapoJLKSN7IG5cC1iHYTJq/163LgCd/G+PMOsbWro1L8A+OgQniL4sZDukE3/u+i/7Cbj
bMaS+QJrepTU9sdDSvfV9fRgmGvV5PTDLZ33qPeXt7F8Qzgz66g6glDdaMT7VADCnCRCIA8nypD3
eQMMiX0a6L+LJcXcZJRzmXGVkOp9l6oW0giDh/mZW4qjLpf/jqKH32dx74/JZP4JTid2VEDmBdOR
3xzJMI18C66jZlVvdXFznQ4DhBPec5n4O1IoOZYXxVjiRlT3z+5wzXJQLYTCjoDCB5Wn0Bv8076Q
4Rdk9IfM+ztUPE+MDQUMhAWk+ZXftH6JOl33x4FjGEwXqfIx/IAnMK83aXvlvEm39dyyw+hRFPEy
Hy3yAIV0CiJs0kz+AaTFKacWZeGOy87H21KTL0wdgvLiM+GEynBfrpppJ45cl7N/G9lRXn6rkPCw
JzrSZF6D5ObAkUsW9ik6tftOcsY+ic6yjNOR11f0VyO446lE+lRFtz4lhKE7WiXlotuBIsr1Y/WM
vWcGyeS1Aqy8TeRGYeQfNkfgDne+UJjEAOzbNd8MlwyUefpgsKf8Ie3svdKnBtj36tm7lPS4RstX
LLILKQ9n8bJBYhQDEfzt21wBIYqXdru1NhBFRmU8VaejkSY3s6bEI4PJrF6Fc7K4tle1dIWt8rrc
y1AB0zWAwyomF6fdtw8hlxIO6bCYBXtEnIWJjt8onWfZDdCvt4SsJbdoYyI9qlncmgUnEMLT2tyf
VzPV6YNw6y1XBeR36VzHUo46vNTYufhXjHtN566YdlnW3tO5Qkl9TeBLjBH1D/iVemYIWTPInMTz
WreRFkZWk+1l1bwkZgFY+S+9wh2/RNYDXWhN6gzvAxB1tSmfoXezgcuos5TeJGDLWjezLCM3wPsi
TFsj1wa5/0Oj8zGWnJBJt87kIvzSeh56ZstJB+mIRVhSgMVlqLZcTc96KJ3QPYP9/BEbZtb54mxP
CkDkbhkguIB4ZKUTGaYZFt0vSl95FN71D26FvutNKfRkcAbp31RJW7jcTR9Ja+sejKPCSMW7GuBO
arXgyPHxYjp0ewljAOZ9PH1j2dOGP/htf5pDHVoWsLLnkSAsQw0FWlbc66Dog9pltdcCzvll7GD7
TQzTO1QRvZHqsGwK7w/FeAmZH+yQgiZ52C6tGIk8HKbnXIUQpka7vZ2LwgY29mVK9jz2ccKrTTaK
SpeMq/LuUcwfnA/0aVe96DJlTcWj/q4ArFPZh4mNmnzIhnPVcsbwMK44AuHvs9vvcOAuI50zkqtP
CUQpGsuxXs0u1XqX4KMNKP1+7dOHCMk8/fI8YJm9lwUXb0AGcGXufaQdU6qltnO1AcuhBQgL21g7
oAFUpm9NBMQ29ChJdyN3gu48/IBoG5L9ek1vGh/oH96OkiVdInYfCAVtiQaVVOvpyr0pmZqPU44+
nIFEISs1oEwdaHTkwfnkGNL35QE8GYBwwF2U6IcfgBkG1gD0s/CImnxgEw3uPt+zpwW07ljraI+y
EhIQI2YYU8Tgxdxc8ZSv+AwDzVkAe3drMkOJE+VW8AlcqpWSlUqC5wPWPAI3E0oEX9O/sWQ7ILtq
wxqmScQELk3L7w1ApYhYz+WSa7lbM4kPb/ToyGqRmcXTkZHUVhXFue9ozbxx1m7Y4qQ6vJbikdki
5L39X9jYNcOHJpmEnfWwxNf8+Z4WfnvvqPnw9+qFDVg0fosYSYWWXoc1EACt+SuSU9gY2i3/V4/e
CLg5XNseVqeE4ZGVH5cO6z8N5zxuSmCYPEODuheXf7BWGGVJNal4cUS8dM3cvbq+1nfhQVV/LdOB
7YGTyZrA7QDLkhHbb9144OLHHWhPXeiZRvlEjUbJVayK3Zi2vsJqpbvqQw34sDKIiU6W/hMwENxw
AFTCxPRmWMeFi+7etBIDk7xGGxNhNP9NKSpguK6iwkYegVwF3Z7md+oxbZ0ZkcpVcUQmn9zAgKIy
fYoF/J9xuQuaBhoYPLgdQaVtXby+U+5wylfYWmf1BXLgFgerQf4Z2dlquktuyb3LYnQGUfmkGpjL
K2fisSWG5o/X3C79ZBvQYYuEK302ogEXxHjL6sHbj8scEPsER3jnXyLyMyoN9yOt/eWbEKQ2FQkT
1LF/SfgzlIp/0/+XKbDHdR/RcUfrpDgdVh/ezVmFg8NTiKFDfK6KGHmEqKjpGmSsN8GT0sNHUNhT
3DamkNCyC1gH9I34yetsZqUQzSx6+G3w1qridMZD17ojaFJK9Slg2MtbauA6kccwzmFs0Fth79z0
yfqEX4FvTTKgQPw8v1SyIVwTGQvY9Nig5rMuOu6BZYPGz8hZgT8AOLJUjdkbLutFCZJK4hnp8Tw4
Rfy+IfJ/8qEQQUFKDN8AQydCLOM4js2OAvCOBk8wjQtdFWmVq00SlWvuhXxaY55FLmUwyrzV/gEk
31OYaF0DBYhmx4ysduEMgI0DHCH26FbUm8bwFPcWgvLsId0dAUhF0y80MZDaqHS4+2nYV02E4x7W
hgvKnG7h7JFQ6RcSGANrTRkp7cMQqSDcH295douBp3aaXCg/KK2cLR2g+2pq4NYy+5jQyA6wdTnl
16gVR2id3hOIWyNXrsiE993CwxXeEBUTHD3V9gwklcnKZE/qtp3RiC1SiUSqpD/29BPAbytSTFBy
9A5S8RshiD9laVtKiG6VvDREdgBBeUqV9ldRwp9WUQqkaiZa29mGjScarP1CcewXGiqXQRucI3cG
4ymH3+GexC+4HR2lEV+8HnFMeeJvbW0iTif5HP0d2AqApv6mZBGN9U0SaNIW4dlo9F4sDVbT3Eil
LzPvV94usPu8YMrP67uAAUyE8ttcqacWU5Hdm0+/OrzNzfW0RDxBc1EIwySA5USsa9wBRV9pomnH
LEvR/mLEkPVrQ7VjoHl7SI/WHERBdFWUKS+3nI9UXZuBBEh20xJgYjUOKCl6jSriawjYGK6k+OtH
byCOnXfUm4mkmg+KwPlmm+o8TYc/BZ17fydEcreTAYVrN+nDWgjeSBVSptaIF0+Hx7nif+rl2qi2
6V/eSem0TSgMu7q/3WD4strrt+7FLWAQP0LA5nsv7QtFs3SpPjpTVyx5qJtBZYsWbXCoNN+dLPBq
7409FQVsJfbl/bj0JdhE4Q5zIwvjPeeX7cG0aBn3d68bWmOTD6ecaul6rgYp94NFBfwl7jLXjT7L
Zyj4bRo8qNcPKz+BcXgNDUJeu2R25+4lvxeVNgF9jMf38epBct0oABizSWJhXBjkKRecEp9Wy++p
oM/wOSV/9zgm/OCXtaiEACAJjM8ZYNVOiFJs3LUCe84jcdJL74DEmYi9whJTub4ZjlWcO+KDE2VW
1SgEjok4enjPnzWltq0QxsZbaSEMcLOBR6c1ONitoKH9cGwlV7wuQudh8KJmdtuaHs9neVybR9j2
WXf0WuR8UK4S70OflqTVhTOSeAIczQ/v5pi+InO8PJN7hC3CZovtI5XPN82iBeNIbBnZFFjMj67V
kAMy1zomwwQ1C7M8rpsQ4TcqUZMsm/0j37wTdtoBYqWmpVUmGmT1tZJyJjmpVUQw2UZ+FvJ3DQ/g
Khss7l8Q6LbmFueECvhn3D3OSe/cbpqPj/7066dzVLkXzFaKJSUFkKTy1GOGfURJl95xhjmYwcfZ
KdPPGfGxLSeU//HBEOutLmNa5np/FXIeXAd/f+40BP8sxc4lQgUT3KewLXI37pkIGrlYKUGqScK3
mO90WwKEcLtWI0QbSfKjKD3sRlpKZ4mum3ngu66G9jE1p9hn0glC2hAJeK9SNLcqSK8uDjPQ6jIp
6a3bwTP7RY1GopSPhyCebhJNiEaLay4VvkETtHT6ytwSqtUsj+Ieq2FeGu2D8EUSc9x/GHCJnuqp
wlaC78XD4vQcJ9gTUkuowwyvoPASNQYnUNxoLCIMqs2IxyFjkOL5h6Fhpjl+vD5V3zZYTY+UWYG9
WE9PNLIrdI4R19R3UJVeHPJgKNlqFl2M8z9PkOAVjvNvop6OGFRHBxo3g3AB2hIDZVhbeWWnL027
Pfr8HaX6xQGQvQbPpxa7hr3o/UgYhPERzo6Z6anwaB0Ti7HxXnMBf/tgRo1xygUUPsgBT18rNn/i
xjBe1y44whwWNZR9kUO9LNJonpWsoS3zml0QRlKchKMTKpAGcGe4nlFDNok6mkjSVUqnRtyvuDsh
8OHQ2MNfF0DZ5VWRW2pJATddqZ8IWY/W8blaptjAJUtPNneI0VKlM0s80Jvypl4b/HQNqvWzEYWP
vake0ZL0UL4GRdglMM+Vyn5hihPSHNQnHRRg9WVtscDEr038prMYdlW1Ll/O4ct8Z4sKYqF7JMPC
Uu5gAgmVKU4sXxJHIv5znXt7SWeupZxJZ2Qw9uTwvOmJ8G2cBqglll7NkSWg286iFfcnfa1wPUxm
96VLMFhImtAiREFzS1z/BBghjr5Oz465XdZzcZQVJ6h8AamauIR2K6KPG8B3jf6KqyslhqF0A43W
6Z4VacIUOE9G9hfLwnuV+gkbhiHaFQzhuEZXvI70ZijAXrq2xUsZ2X/dXtsNHxdeJKg8nIzPDB4P
TmbKv5mgFXAZCOR1zJySYq9PoEkzO8d0X+t1euoaRU5554FLcw/PZf7zx93aSrX8OdoKyn66Hcbp
qC75FnkADYh/KhIRamf3kA+3OGH4RXl1cUopmf/gYlMu26e0Tgh8WNgDyNbxMhohR9O9qvBfSTV0
op+DQMFvp7UY5Cyo2mknKg8ESNHtbwzK5lcwqqere3JcLhW3k/7+Io+9H0dhxMamM8Z5pJMAeONg
sOFivswccpOAuPCji5Brnzt+m/Go1mNHn3ClyfcO+ySBjRfXule8DqCH2O0MYTbF8axLzgOD1+Fu
RVASKA7ScWmfTVZuPatGa3Hn7bCoViByIjxjCx2sgFoEBOnkhFTT/HkiGLSgIatni4bsL1rZnW4J
8WdWKMwIAJSOkaAq5lkLSb9acAnNQU9pARtMMEvh7M7jiXrqapBlryxo0xkR6IPdOXb+MZkoCmvZ
fHtX3rA66Hl0ilxuCoUkr9qSk/wICg/zUh+JqTbfu8ydK67kIL9eyywBsKroYaQXzPXRI85EQJF1
vZmYskOAD6YObcUqrb/kl0GaVVqznYTgONo127RCsGK/GdjQQEJwEUxmCVHJMoNEe35QUt2sCadX
XcSA/+1yIn9jjb3v9eBjoheLOAtg5CXYaFnKDRRfts6MPEhTXQTjg0cTjqw4mXudj4qcxSZ/7Csc
pQbiHOpfnCfGeEibsQN/pNe/XduC0E21hMdIYAr+Zw3REdCfYGqhU8gIPwuZap4QxQn3EAUguB0s
2w0M9SPPvdHhgG71/IhWhiRI4y730xbr41IKuIAofGbIAjmJwwtXIxutqurJjtToLuEMVJidrBhd
9lDjoPfH/AKnprHGCSO2z0uEzyqGlxWMK6tFOJt/hAAItpbCJM2NaNve0O8qkO+KWGiZQi/+x2Hf
3X1T5Yg94w2BYGv9Stzsavo6PYDqkzh8tk9cz/FkcaH1HkYTyfFeeRP2K9TggLteKRTiFaDq/LyO
jVGYF4JyaISiTlM6GTlcI1uMVn7w6yJeCOGlFwtRYR0Vkp4rVwS7PQAyjffIiBnF93k8JBYOMvx1
5KJlId39zxHdtz0w2K++fhkBa6l7VIz9WNl4tVSNYbm0g6X9gt0ZD83H6NEIMPVhccFke8brwCl0
/VHDJicLvqtBP4TAW6nEOBAVUFMgj3pfm7SOUvaUBdVpqn4h5JdhraKqeJ5lYqjfHQ7vFmLqRBT8
LHMhp0aOKw6Neg9iI3OxQsCWSw4UGZWxZr2aacrq3I1CRE6jacNk2V+yTu+oS02vycnmwQyrIYsG
3lY02uWcyKmd5NAuFrOkXZSz+pyjgBjH4b79BM06WQbTen/m6PI8Cl7pcAm3DxJCRutV7rmBj/xA
FcWKzb6XrLxnd3EbQp++mgTS+tkMzsEYORI0A8bIZ58bycf5+812+p5shHoxotVbCqErmzZQabzf
rN9clBz0tlx8QSRkYqR/dwRsr9c+WRfeT1AaVkbRbiTzmCm5JbArqb0fxXWtUAgsFo8ab6X+O7Jc
grKKMN3L+/Gd1DdYXyTIm8Mm4EI5GAy9TISULIlD15dLbE4/3Th4Dtc81b7JI1iJW5i1wYKPzj8h
7X08hH595Ake8kxPL8E5SCUdvVveV7XrlVgngo+8OpX7haJ8DjngA4+FuoMtawumEOewHY5DRR3R
9dcERkZx4vCne1o9LHpkqQi8/jNDN86s8FvUAgfzr4sDTz8eTafKMamIV/YYUNOJxCOWc8QxdpRd
SiyV+nwYoHwWIIQ/2/F88gGPKSl3+nEKjq52H6vKmBNOIj9SNMMfx2Lg6hByhc0q5p3F6YCoUB5x
LT4O7unBmzoiMYjn8N8wXqrtTwlBHaj2o/dmSM2rjhxkD8g6zLlLOyn2lL8AxPkiLwcPNnfE2dGT
zNsS0YdBDcrS4yQogQDqdcIdeaAN2UT+7ThCaaex11fGo/UB1iiV/s8kyqqdkgM8F9adgJ0SO4uU
YT2P2ZTwm5yDfVDIiW2JsVpQurxiN8zCAuZkBhv6p7Rg7CgMHv0m4Q/zGcSxZdqk0J1/IRzn39Bq
+cGS8vruOlTsQss8e2F8ZvQyTfSvL933YNeQRmkcRauLjVRgBC6F27vwv3vs7wLSZFlNYisKtrt/
xdzvBreT7+7Rum2g1uRtvjgUbQMlbYlT6vBFvb+gbqB7oCCIUk6qJb2I53Kj/7pofoAsMbUwJZxo
iyQ8l2ciiG3UORfHN6lvqo1TCOlcJSmnCQh/YBzNwhrBg2NEmCTEI2upx6T/tmNb+BNPb/edaPWR
HZbr7g7YfBPHoC2bbjx7+kUS2pU7Huxe1xo5GUN8ELsAfjnOB66JAQuW13InF7uuUoo4keW924kH
dKBfujbMdM82XrqN4ZkD2KZmgWW92lrFRwo8TP4mk/mF3/rwWVEUHknPJk8V4Knt1KSH7KFIXxYe
kjaWVwRnHyTSoJdhABARyrbot7LmWnUVMcm8nEhaA1COFx/2XEoOzzpApfjd7vVW/rrcS7kgnL1Z
PcbtZZhGLo7eNvRRxYlmV36EUUez730SpW0mSK/zMgznsUqIRc/gMuJ9NWCnGrfgRbkF+VRAZY8Z
oP0OK51MdqJ/mpa9CJdlQC2ZP/gOWnQToZqhi58kULsMkA1GcOBJ5V1CTG8+F4LGni6k/DFB2EYN
M0Br3TKVktsEyudIwoNSHulm66FvBQ3QyUxviMTSCvm6gRZ22tMWmidzLY4Ipdeo6Rn5pJqZIw4p
urbc7kk3tNzIQAQGEuVspfmwU0ssx2RRMx4AFzRvpKtDyLJ5WULMMviGhsTNgFWldubtSQSl1et2
xVKf826NDxbVoJsedMTrIK0JvrD69GP5OJ36wmE1MEOhMmnFxcRgyedZZ3ETch1UPDsxlZpzha5n
3LUP1Imy4ILLFRKnEX7AoBwKclEXQ4/bw5Nx7GDPGFhOqZ2oTJdLT9e2j6EO6a3DMD7h9N/r8JER
kPqGkBZBINZ8O7kBkMuwE84UwlpV3kxFk99Egj03X0RteaBsmWdUbuFbUc4pmWb2ZjCfkbGqzmvl
wTY7oLSgrP15ml2JQd7NSVkpn3Yo6GlCL6NEyrSvMlQ0QsBxMhUrjrgqhRbc16Kz4emSSvbiuZJx
gQd0u8WPwsn5RkgY2vFNUgG4tmbY0RTCk9RYoiTvNQfG1jmc1K28bnVhn0NxQX6nZEXltpRdGbCr
jllZw3g6fQIZsrK4UiiDrrSwvcKNFFggr/AibyVs5jcJXL2FXu6koZTD6HY2ze4Orb9curS3lanj
964eks6bKNCv+h9EvDZrEBspa71q4LzLNx4QIXCkO/Yc8fZ0HjV0Eg5miwpJxp5D8JRdp4auqM2o
ibMFpo0gBtz36JiuxBbOKmitEFMxGo1ecGTA4M0p8cT1YTb2S1KUPaFr9kUATMbbXUvIwy2l5NZe
jpQajxRfKSVqIyUSJZdX0BNLU32prG84WPTMqeojkLyxHGWPyTlnPoP/UbznUwcI3EDdLfb5p6AT
92y/rW7nLEpCdJUNZrzZcKpb2AGVDWPx1lBBCnX4vB9ShdF38aTo0kSOE5BWZDzTa13hnRGOl9Uo
/hbd89vpcANNrnIpanCEZz1S+Ja6mFlPTpFkhijcbKFzCQqBc+K4uKdIWmmImhBhQ+F3mDm8FxuJ
lwshwIxv0TEpVmiAqlUFNZQ2kVdXGQ+Yr3kUEEedimVmGcHXMsutU4MrbY4G/SXldZN9k6zHsXlf
dQSIcbwKWi0YWK/FaU4YnVZbALFNVJ74ei+qCExVUGhRRZy66oqXl2Pc6Q7AVTFCK3iedup5VIko
8Lj6Ue/gQ+lY261HQv379MC0boiU58okY32tdvsfu2U+RUbodSK3TEpRf2CONfkjYXscW9IIIq9A
UAKv2RWpVcdAqe6pnYlk5cnSp2+tnz8PDHfRw+1CNT27As6kRhutDZ9lK3QDs+QqsFOHL0e45USZ
GqKyL1dOfmZQyX5GsfgeuuXQutRIXVSIcqMXs34VKiVay7DBGfaGtPImUCFLPyVcHxPY4hTvePcA
saH3ioM/Ibi0NZbo2LgX08p7xALxkaZyTqso1R3DI9tfWvrKe8Opznz6IYDlr9Ucd6cCp8wTLmhL
83vKo+BBZ0aZltzXca0SiL0tSnsgdDKuuKZQoCwcBbbNiJque7IWQ9ycMt6Y4b0J3Nq1tZ6dyCBS
5dWxefzW715VzSguxWMEaMAuZy0Vz5wF50t4+3FpZgpIlzNdxplJ0+StFFfoX4MvCtMheDTS325T
9jHx0Ama+62MWRWsk8v1s1M1EOEslM+ctLxPBGrIY/cfoWIY8WMxptTjHW5V7qVQOOeJo2WO3kJP
FVTZrfny+iW4cz1fdYyp9mpY3EZuTIsrGsRrrHp2OWKCiggrCKwp0jtUU1Rx3f0UbST08y+QJ3gs
JjuN/OnBnBIjN0mhljOmC+X7Q5CKWcpspxtXFnt+dmsptRTm9+wV7qHKKNGO1AH/CrdzqU1m/PyR
cPINI5riXfWDcFdRN+WdKN4ygrmSnGaUIOCM7E/b8R2Nb4dd0CcODFF60X1WkBy5/kgqlT4sxma7
F8VMCIiHpUoCVJnF1yuQZGT8eC3B9o+BnoCvuwUwL7J1qRkz3pAEwwUOrimB+AwQRKRIMkhpUygD
0Zv0pnFlwSMdrtMyqx53CdFpuj46PblFToxNCIw20h6QeNMdl8sHQ+rY+OPP9KePj4M7Maykam0o
JQmOeduEpLlOE0Z9Fk14+mL4JzrnEMjkCf8Nf4kZQfbK/5nDiGXEU0CHABnB7bf2FwDUIxHYQlrx
jTXKHUFuJA5o5rJ+dixT6rlFw2zeWXCxpWTO8/r7lTQ7nPfZanI+DkgD4LWbXLse4asbbRqTIAOj
H835ju2DzO9VnX6ZI47KEyVY+moDVVujtWYokcE2nz8kRiGwMtV9LCGzPrcBF+mZF27FM77Mw3Y/
1aEHXbfE4DMjLffUSIZqVjgu//EazZCqU4vt/V+n/6BMiumNRNA8BKcqekc2mgKrseW/ibCg/y/y
w6//3mygXLTvSxLyYFO+lVXDkkEgLTp6BRBK9MaJRRh9SSjFPu/Flgt3zkBj7E2upxBOSXhRLO78
XhCtiG9Rg7iq8iksdfjFrTJl4jr1wOwwpoXlIec6cjmrHGt/50qLelsalxdNgpXHvgxd3YKmedfP
XqbE3tzag0qc237TC2wwPG61wfhkeXYbjJL+DPSzn2Xp4YwHaLVRz87HH+xxrQUSBaWhT1WEFDgZ
oj7TAirjKsa35rdVnjf5UN2Js4LBl5aCwPon0JC0HfwIotzex9W9MG+lBQr5hEdg1RCy6rMwqvOi
IemkH5sQWGZpR7nS0shGPC3Y5I60puOnayWcj+8XdgPS7pHmgRBSeaEXAUA1NccLNy/evnKD/Xd/
gKZ6MT9zMxnfBKEXq/yw8EGMJFQ/2gWzY14xC2sVjQBLqYUv59eG3nigwnxHQyxKvcKmXoPqvl6r
D4izkQkZL3kA5ldWlUTIDrHsGlH1YMjpir3kPELNHqiD3UsJETLkm8wTggTeY63IvT1om3HnpptZ
AVgNnA+s7l+82Ee7suBmn/X1LazcyD9IE4kDAQkVeZNwwzqyIIrEON+MStWSkGNhbr7EdT55F0nl
+hKHPkra09q6C9kr8C5enqcPXA/KiNsvABDU4tM30SYR/cZeFvyPgHSO0zUq66e+gvUOZz5MuL+N
bUlMxOIoeHk93UG8lKq6tJfSROMcSw83Z1gd5ePI6iDw1EQra9UhohQ1VM3pCobGqNA361KlzxWO
sZ71J9J6fi8qPoF47foE+97ogZh+PuMg+OVLDJKffDASahk5yTQEY8ryb1Bmh4/gmXdx8FUkO+Mn
KGIPoARNubiDtu5GuePWEs0/NYwm6Ql0jBn4qgVmY5MkviaTC7V+0plrlZYBpLos9kX/+eBlvJxj
MWSSjx2RA+KH6WKovwMLoLJy7pGdx9iFbn9Rr4ZuL9dXtHe1WkD56c8A5J9tfBu+hTb4DRQFiNSt
8WcHF9H757lytYagt5T+TvQd62gCOQLrzbT8t8JhhyiKfsSYXY5C26bBbM3TPMjOs8SMfIaAg7CI
xLP61t5mF/1ec3G8GPbt1qIjW8QpkAWyy7QNE72x8D8D9VRTQazgotfZTC90+sTcABFGYxjAwZ6I
i7iRKr3i0vvOOO0a+JDkw+yTm/j43mpWeX99YhVZr1aFmWmknAXN2HA57Mh+InXaSOuE3tbY9XPT
54bwpu3NrUctHMU0hDx+hN0CLJKh57DDbB0d2FCqfl26aS0yzJ9E1qZiQwVJzZ0NTKxSUTfgiGnD
Z2UYwVAK62fS5tZhSLHQQTsxdXkoSnj3DN5vPFfU9T9AyDcMZwOQndBDfr9E0175eJwN9wKdR186
XWCs52VT8wC/80shc0b/wWZlx85TShsydRnmf3tvLXm0hz7X1ifbzrRm8XrAO699o0u3jdata5Mz
M4Vi8F4sKEmqFmuD53l0AXKwoPG+Rs00uI/jbV+taIz14VhzHy5C2m6885jQ1LCNggVIrwgC+eG1
97MwpbU/nVI/pwn+eLnMfQRz6ognKEXaT9Y9TfhokRVgW8eG7yZAgY44ICEMHZVmlQm80K9X4rkT
FQVI78Pk80wvasXyWZBJYjYbvX2wyI9xsfA7cbUt/8rGmu60yhgUn6MkWGjAUlw06VN3jT4aBGyM
aTLTQ+mFY6PdDd+wL9Fuf+D4P4GaTVf1ivZGT6d0bQcdj/W1vryzrjnWCVeYMiKCua3/pjfsJGRM
mS+TAQS1ucJKPaPRXX/SG0qsTq15v+8KNg3f6XQg1mxJ/iWSODTvNc3XSIEc+LEGr12Ik67D7c5I
WL/9CRfoRw8locH1Kco+9+LZIJpmnaopbpb9/a13BqOXy0SQ3e27x88mVBfD3udcEM/3T6N5gFCD
WCPBIxHibrU7q+pIkYqjm98YYjKFIsJhtY97zu8HaOAJP2h4GVtUY5Dw3QG3V83306X3Ok15dP3a
0YNmlA72LOKO2T88BEb7ETWfwf0RV2Koj1hVLl7qMGJ2ommsiWb9r4g4quE322ZwmV0fH9L1jpBl
S+9MAExL1MEEB6A/OnPkflstMa36ycXc8k9nzfXnDYWL5MN5+8Kwj42I0DicLNdXMc3vrleCeto0
9JSjlWf2dF4TdE2wcpLLrgX3HwQAT1/SlPCnnx7tYfVJBKQEEoarJ3UfFFfgjn9JIM8WPqC8P71G
VNGIxLMf1EYzFnPqIiOsLd6CC1bj3gyCrriNq6G6ubkNZXSRImnddXfbGw/XN/Zf0/7AidxCbWBM
vtEXEoaiTYt+3H0xU/BgzV9kbxgpkFd5GCqVzVYqJM4hVX3uqVuTmby69C/D5hhV44O/GCWud5D/
7F/KhFNP9dwV19n4PfAGGZuHMsHryuqcn451dCcO9DBFHYZb2wihCuJxfrz7UCpAq0ztYfl52J1n
FtK/jxDaA6WjsEOGl2wxawZoE8f956qRA1dWO/cPmjouCp3ku/6wEg19SJGkdcPN1zP/r/+ZSFtE
l3PThUJupb9QM3b9X4bI8LRRALdRr6RnAKMeMi87zRXrrJIdApYwW0GP1f2gP3L0Sar5jYbg/OrE
RiAq/cmR17gxQw7L66hxp/8PXXIcxlqygAICeoh41lxk67hNWRAK+SpNP2HcG+/UwmURAAISv24+
bLDzs7xdr2ipGDtJU/D7h7OMa6ga+WRofCkIUODHnQQcUG0dlF1zsoNe5J/Qzn3px7/esJhDj+vO
m5roxs5UamqYxdPbonUaxkTJ02yKQ6rAkbTS+Wk8W+NMUbhZHktB1NUabnjIrA1gywyg+DeS/kJh
xyPVOJczoydST4kWln/L9MWuIDC7wxCzjv2gXz9HzSI812B4cw6ooE9NS7BJa8y5SngQciniC75G
O0HWg1JZ6uioVWfy/nyIofbgdflqXcr8i3aQtuxYJuY4hlhGMeW2765Patk6I9pEXcYl+Vh7OiIu
GmEICuTPbvQLx4LmTUWMX8OY0XmWNDjfoNmzA7K/wreoyh06EmMhTdYkpNPLugwfMeEDaCLrbqBk
97jeZB8cFMZBzrOUCcvXF4mk8/JgRV4CZ1uldi+LVYFUbY/HmSmyb0kPdn1IQ9CLk74ipM11b1po
qBb6kAumsGMQ4ZKd0uTKKHSumkV3RpnEdQAqL6E+Ao1ZEK/WzRO1NttzZ65gop6fczUqe3O/2PgS
Bw3Dk+VmrC6F/FITX969pRYki6CNcEmzVtWFWyibmJslsWT7igGBVX1SxqMvGzzC5amQoIs8Q2HC
tIOX/wKLhvw0yeiVMaXUBteulOzibAwoNRfFwvoiqykTT69/aAKj1xocQF7donJuuhIzcGu73AId
j6XershhWJxcZwDCBN5ec+ysZUBK7JrcxlyN3ScX+wPkv8poUK9OnHQTpf4e55OUCdMBYjk/ku8n
hMChhWNipRC13iAK+rc/Ms54/f9bl11Y2alkkyMHPWGUmVWFPSJAlS0ZWj4KecmgGeze5fBRqihB
n/Wo61vz6ZOVbhiLIKR5xiOj0mQUrPL05T2ue4qAvllGHc55qZ1K2Iz7TXdasmC3Hd7zoG5L1oVR
G0Bgq/PGcqPQfXRBsgG6FQKzb2K0QPHg7oWCQYwfsHQJC2mqSfPFRK9B93OVFKoBk066i+ewzCCV
rqwgucGv3RhpL/TjEMOM6WCSlHekpiWlGXb1Ldo3EmYd/ZT/UtcQFZYMVsNkgG52a7CZ90uO/ZOz
JlJ3u9J/ySQjspgMekFRpELA5N0q0kUKPudR+Chj08XORgkyn3AmTDixaHUG+hoSpe1yWNT8omqV
VTXzktBrIUfFTDMMj9KFQipU0aRFNzkCfie37HKH5VKLzA+6Yjw/C6zREC7oAwTXpHplyKtoQvPN
RoydhUrZASkjg/VwzF7oO6o4lyQFCjC6R2uJ9Hsvd0zOKO/UD6QFLpBV1CPX3EN0/9WRpg0y8Uit
9UZAOPaveXx4bAsiDDdlI70GpT8ZJ155d1N0FXrtN7OtaVQiypl1fvau8/6CUOKbvfWkunrN1XGd
nWokCzEt1J16HFziXbZoGp9nFy7XDmEZ0i6ami87R960y223K3ueA4Z+n1jfSxD96qVNIUTVQWZe
NYkiyGzURvLQIYQOvnsx0EGT0LIvDjzl3lsgN3kNPSzsXqZcjYTuhMQapvjPwQpnQha0y8SyQeFh
2KcGJpkRVZAXSi/MAZIBSThAPRrghuCwTRi51hDV47+ArTQiXIn9aEpwMptE3BF4RgM+roHsIUhg
tph9wxk0vQ0suKsjKqiAREZ+vJI9iHMXYpbOEZArf+VmDtdzg6tZ2Yy7g+VwbD1VQ/LtlR5R2Emr
Tce7acTKsfSEUS9m/YPhrZ/ojqVgwWMZYUBf3fSBBS1OTEl/a2Ksga0Tzw8r3zcF/wGb6imsJ19D
YoBuvvvVIxlpN6f9x77xEEfvtLN2V78T0+SjzpMEsXPm5sql0WEut9mbVmOJB7hpnexmgh1hDu0A
FPbzB1OmHdmw270LKdr2EA2Iauz9qLp59C//qW0OgAqWJRfzvtQPkKWbS4bKVcMo0tC6gHb5EYM+
2gQGTMvwjkygRABnlb07mKz2VZ1+c7s4VEobVpBZaGbeIMwQ9KCOOsIGIhdNVunO+vgq3zYZbcPQ
1w6npFcVR8dFNUkQURJXOiruHVs12BmGw3fVOdhA5H2bvxpwpLWIChVIh0bJS+zwXE/xb/RtXKD/
NAhJmGviPzwqZTqHHL1qnhf+iOqAUSrOFi3chaiVdh1I++Wje/9fXzfWax7oPjWu6WsXOQbuUwj1
MuL5OBCErSXMF93eTMRsXP4gcNHNxlNynDOtxYnu+6vp2dn/219UIOVdwCdESFa2P5WmUuAO7jKU
fTbZkfYQAeO6vsuNewik74T8cf4/aBrjL0Ir9gE0y0Deu0firf1eyfFOIzDJHIDoA/vPRjKokVv9
bumu8A35MLeNm6QVDlSVQx8MZWPSwX2PHmrHX3/vNKPOnfkVIWzJuVJ4y0j2erXq9tr4jo+SJBlf
Nd+55buHBuEnOuAvIzNhwQi9s621KkRE4Pn9L3HYjitFroL9j/3LcMUScuuP5G+FB+7lsldjJMGr
0R0LgkO5WxYMpndNmYH8lcvdeeOzi5bD/oYQLLOk7GUzQYRC/bE/cHJ4TPl8yxEyn7KDKKLcSOOj
F2MEE0O06SadQO7f/6xaPPBPKPjsaos/Y/Tx9HYzqg079IJRK2lhAAdcQfbd2RAl/7gU0vq+pB3U
JsJcZvYn32REC1byZM59MfDXjvlEDMuwcIX74S8SP15pJCkbXO/sFnCUgEQXBua9YVUGOEQ9lhQ8
CLBRPYkzLeTBbz0H0uht5BSQFfuQ6sd5yB1piWoOQZNh3i2p6ZE8p6m60p5Gl88bEDbPjAJPHIVJ
I6lrACAnRwTGtgGNnZN4QWbvTgyueyzgzV+lzHVGf21FMGvNXi7jEwfypfjMOPUlSzNrlmIJFgjE
bD53acO2sVuFpTkS5VMuLVtH3X150sGsqqyvI8f24c6hgVf+8/sTCmD/DMn7oNapeo/WFsFwoQqL
l3EB2+x+ETFVyfOKxvTDoPAfOMNIDklmJiZ7y1dcOG6l/L4bK66o0s5KG8zWQzlrZdelfKJ4MskS
KKgNstWR77kOmX+UIpe1U+7D6C9WiUsb5xkM3hA3nx/OKKDaD0QIU4toAljKZpPI1/ziyPzR3e65
iGmVBBbBuHZJn2HHplqGAqO7c8IfTcNqjxRmnLhO/GSml9djZ6C/muYNuBU046eiyWNaH2wiAfiK
5fcmpMFhIfJBAiIc69/N6kzIwufkOlKHps4rlEzoDX0Hsvg2+Caa4U85qohJfKgd/r5Tz/6k+xYc
4qW4qQEf1YQprTmf+BRr64WT3fc4nysshGRt9WpvvtomnZ/5A1S5k4lH47q7SJQRy/WeMvhuK3xs
wdHpmScIUq2pZO45BFoY/dPOXtfEPvix/nDdI6w81HqyFcRE3s+S+2LomDdMik7ChXtcMPEFJJAj
Uba7EJ371v/hYfZMu13K9a4nAfS0ry0UhlDJkEeQabuOwDUP+oNAxE1CkBN5ebXmcAC9Nxzi0/oP
FdsHW7iehtO7PkXDVJKNuzvUBU9gyjbq+JH/8YUvTCdG6De7N11xhz0X++aEO7Nq2HYh00r3Q+lS
yxZ6UrAuzKBZ6iLMkFks/bMqEdDiRr0zBmKXp6kTTNk+ctqD0GZ43IqvYz0anLXSN+FBe+wRzYpe
R9crQqz+hDXQ5G29eZh48vqH26g6BHDPUnlB0YDMx3jBOhaC9aDeDg3uqvU55nk4+iqHa3Uu+2cK
KiWQGXlP1mSDjtxKwvvgR2XFKnN0iCBu29JBgElwSsqDpMA/rQwcvnLbDPPeqGQkks5qvRUrONki
g0jTW5HEWwdwXClElRGxeNfA8lOFtnkS62c/e2uk5hDKei2MvD0nDMc23ldN4JZ79rzcf5g3ovB7
TRMheVhii+zkoJzLNn4XnxPm248sqk699iqhu6VzUD/Tjh6oGLBW+0m/HI6xBfC+1T5+QsJRV2no
k9tVoaY4XmO3cJC3OWtqmmhCQ5yKAgLtHj6dZyBYqB7AbCEtzE1arx+dI3jMCF4r8u7rUGtzHnCW
p39BBpI1+9C4x8gZzEJ8uqJ95073nZaBO9cBBh+9NrT862oBO97QbjRfJYE1DWW9+iBaE2B/RcyN
kD2JquSe58qFwbBMkA+8IrN639sNU6oB4gjLJvjnosu8yd1meTey3ProQNH4jhkOdoe/OdzuHRkH
Cy5MGgjg/TeuRrc3XRCK87NYAtLzfOzV9EXknD21tFAkIUMjrI2nwHGHXb7MPdQgvAQcebDjrZSC
9f7mbRJ+Z8hPn6Nlp2IFMJR3m7jrwZ9H397Ey4yxQXtUwjAqK7CbLCNLvQLHJEn2Eu69Aj8+x30f
FaCp6Eucco4hC8MI238X4ddPMDnhY/8aLNaBAIm+vGKj35tD5HcYaJ3fmCshnN+h3tE9ckeZzKEI
R5vdUsS1NPzoRiffnb2leM/BrtNRskpFSIBnbJ1TgPNEjQOW8G2EB3A0Skje05VRPkdnwz3RRXga
KGL69kRBruKjmZiOLjnrSbO+Yt3K/ZAxox4Qj/r4Au/nRDYOguHBVe1fPU7/UVQv8ePrMfZxs8+Z
UpWcNMHckcLsiolCdNEAWr+sJyJuTh7uDWHdYsrIUqiuGmITC0kpX/w9WZAnXWJ5agfg4w6WzCBt
VCMvqVEMPXWyIaI/DtfadRF29N/c/ggjHuaf/PaBDdmUnn1qTl4KRXh0byw5OZjqVjCZ255zOUQl
bugrPqEWhAI92q3/cxbMwJtDgEO7gsS4n70Zecg05GHEBdKxviJD/3rkKd7XVIM9B9VfVWPzPP4Q
29XXA3PmPGbenMrigxXX4XhYKBuPIRY5CZcuqi4BKb1NRHmJt4WQT+MRVY0L/HanxEA2Pf46lpCz
NVL+9Nas9pNTjn3ifUUJ+A3XXReJHRClHh01ESd/J8E5Er32x0hRCUkyTiuCTcA9FtXm/YZjrMbe
oRtkITIXyiQtreUHY+HqMBYh5U50Fy4evjY3lVI7lt4tF+79NdShvLDNMepKmiiIQhVHu/SIkhuy
AJ8RNQmf10Hsiz40xzF+fepoi18stbukSaoERg3V0pRG5p0bcNYq22Ld9RpI8akUedDMlwyCeYqh
p9vHNhZmvx1VrNAkrnFxi3WyRvTASqH8q1kdihmeA7K+jAvtTUB5LP3d6Jt0ofbpTCLSWUIhrylb
0p+t+ap5rwz/y+doikfMzfhBZxZjfi4i96gJYJWjbyt0z+pmxtq++j9zjbFaW14ylN42N3MPOGTy
tt7qAitn1Xn46/a1BDkf9x1JGq6CoQgWl+hDPh0zUYR8onR30evYrzlwELUmkdVlyBkCj7DdRBtJ
JJN+Y/ODh8ep24piZQj/DOlFncw5/z+lMKK5syN4y8Jb701dX3yyNd7q1gHVcIS2gGcYc5jA3yeC
zd7BWT/UpwXnwxjVvWdq6QrTvSZGvW0azdccm0RHZ5h1Kq+zxKWuPzzmj6fJaQTLOyU8Wrigx7sn
3spSEMCe27sNV9aKw/tqWuhRgpvtUs8XaZxjp84SnVdtyz6F0fYhkEXcOHLY4msFYtq2cQyaylq6
685DCTbIJ8HHPjtB351npuNtc9P8l1lIWInr0TTUZ7FkISdtmNTszAFhY0fF+J53R0zsLQ86W0QW
/jEBhwlTxwkbz6fCo+RVyP2IYySDA+vupo4mTETLcKRB8xD8ddtcsNZ6zjsXm/bX55Ts6uOl+jXX
LUhlwb29FWjdXoFqHUO5zxcSiv6OgvG6n/U4mRJ5NaP/swxqbGtGJbo85I1O7uQ0QhsSgvq4l0RY
+gmMQ/nLlP68xq9VzTPI5CJdvFA46OG07nq90Fws0fwApXWIZw3EHIdbXAlx2d07YpwZ71BLXdHr
d1ZUtHLplBvuwkcQvKFjfkcY+s30P7LCrk64ynfm3yuNq9QINbshdPq9wTJ7R62Y2U3qBUQn9zCw
x4vdZvTuSZTF0CA685EqNuVoJsKh3u3x8MIvYV6xZXaIPW81c6cupAEuMAsldnGRVEwtpi1LVq6t
EZML5NxNYsOtihvQQx0WiX6I+EpAwdFazHMifhyUNtbUzL5jIHi1XuZwYyFprCzQYVsbBWjBbleG
iDN6m91qLqkGz98SPcFDiRgJKD9hJiBOjay6sa1Hl+/o3ORKT9J9R4xcIJ5Xh9P9BMlneqzE4stb
U3cyxWttRc/7cjaeRPSDATSMeGqLOBM0XN5hBxgVMXhiE3KT93yF/QIt4MfrE9JLfjxRKwwVHEFR
0XW/Z26XEq46hph+jZc1oxm1Kai8kebHvVsBxaztwLGRaFpYdaNZ8MejsijWEvsf32zjGZJ0ud+C
Qrf2Qq9tgh32bRrkaRbTEg75vI6wrp6vVG1EkACXAiP6ecV3gJz74QiJMY+s+mxAoxEqMgJLcLnl
nX1KmFZr9AyPJ/DBV6uvRBzSxCQJqqy819YJHIL+5xfaaRgWJtVxg544DTbXFrxbFbMndtOPaUYq
UefXvedV+btCtU7kCwIJ7QosP0es0t7ht+89dGJ4xKylOU7pvO3iDvejC3HRUrVaT6IiGa6XrAUz
4sLvfHpggoH6N89CVX/9IupaXdKnNIMd9zTg4h9KMvo2XOA+CxmJKLJ6PmVTpCv14mUnx+uDWJHt
UEOYa0o0xaVBeT4/uTDw7UGn48Ip0l4ILA7zkhVjcsA+qS+7vOSIyttVnMxwdpCC82maNgVWG+G1
+hKk0ylzKUZIwxM4FRGxBBwHND7ihKimoZgI3CuvXnv9hAPDZENOpypDDvI8K6Ebm9/Lsld44RUM
7lRf9XenVUpsy5kfD/4N65MEpNax3GNgrDeD2/vvlcWbq6K2S41+MK9J6vzDMJqU68P5Twf3gDjH
iY/V+u1sPqRQ40FwMx/qasT6ztBe5fL/PZHdd+KEC9wdzXp9sZhZgZ8OqO29Fos+KaOObakXpUU8
7isRp2HWHTcU2AbgIYQ3ONFyYMCDDxzrb+BT3KsEhr5PGSuPKULtGEK+3pUx2s3VWnrQ3b/sg48q
vWRhETKqFYcs6E5bYYGQwRRZZZbkNnLqQD7w2sosrupDQlkkFcY7loEAdL1rD0CPKGzAsgCVs6EG
LPhGvopPoTE4xlEJn00dy1gW3QmJDjKtb6stUFnV7tYbhfCwHWjbnvJPFc/dpj2JUjLnK2hhF8Dr
YIOHu8oPhFhBnA4L90MuFU1DVVEUDMzfcsOC8oQGxji9QTRUL27Qq0is4iwrt2je6WO025qHsOhz
yM3AiZ/7BuDIMxyUIWC4sJlgMWiAVPXZfxerfeR6bJVWyYIdaQLzERMXv/Fr/4OY+OnUM3ap0Vi8
MxpDSszAEyi0maSChYxgCg/yP1qV99g/JSCRM3nU6BycqltnDzh427wvZ/FmfXv09x1KoZfJlfGw
OZw/AEyXFPiVJPsNDFB7SRe5P1wtz2jA1WiHzvxCQJiUh79GHql7a+6RcJccXMLIt8fxEaAXSCU3
S3YCYshS5mauj3/P0LfG8q7JJ+bMm07exrDhjzCr3FJ3C4CAmujIdkk1pxNlTaphqB7v45Q5p2Ua
Z451PXiuIkFkLn/eiOexExveJzRHEe1u1gxQWLgMNPFUc+r3TMSW0JJXMp7cXN0Q6uiQMqm1dFTp
4xi4nyoOAhQoaWU+OccdmKrdg+d6nWvfNGE4WqzpoWrAr8gyDRLk73w4Qz2d2IZJ2h1WwyeHWK19
xXI7ragWc//P8f86mV3HOarZxfp4R9j+vrBgiYuLiS05ljx8m3KUoPqX9kYjOKQmXkZY46/rChuG
1Q4flhlg4GAgZt7dpabBJItY3jfG8VCdZZ4R0kcQcWDmYdXMfV24UDW5/PzgHaLSMNrwfwlibzUr
SBZP5Ib+GYSTNUOAkFxxRYrGxRupaMV3PU75UBZtapTDfiCAcbAGCQSJv7BUEfbgTGzvw+deGu1C
JrtCdQA71YWgs49C2lHyM/l0LnsvD6li+5jgznMSC9wqyBEEbs/zrfn4038fpZrxiWsn352ICpql
zeTEbVXklghTHkNGaYM6c5cw3P2sP95EzK5cyAoMDTYDnB/eVSEW99zseqUvJkqjulNeeBLcNnzW
BcPdkEgTTmunCKHo2aFiAoIhA+JELchHR+3T5iICERPRV1/OdzLVfqN+TQne2CQ6blHJY4HPvb05
5BQc80BfmFg+Yg2ZouqUOTHsNXmG2pvRADY+hUjJzIEal7w8AGJF26upM4qcG8UT6C7uLwRPSHx0
OK08YHCZHRaM0EDI3e8Hh2vgSzLJnwqbDm7ncO4gYjPqhM/2C8RQMcD5WOgc6AnBc8obnSTK9vKP
GfowFOiGZnN/BFNRGrpg31R85vUi5kUgHaZL4KzrvGJeU9vMiFPele7kOyAW6UMM2JQ0Zc2RLu9/
QXbNw3xndViZ45NohmvX8Y/rFk9zaGpb6ThxEKp4p0aDEMgo2rgR6bHzQsiPP/mrvuw4pAjmR8bQ
6vwuCkA+XJLfLzhQ1k2Vx6I+wyIm1wr+fr7lbU4jsf+J/QGYxVMMk+0rwHs5fdr7ynBPMqi4oIIR
yDt8fWZhKUcn5S8qavbV0Gd7TTek7ag+l3F7+0uXmUs2RD89boPmyX74L0p+OBFywBYewnlytJl2
cXXFYgvsE8QCVnHBPBT5mpLTFqlsMwUAxpMg9pfQ+YM41FJgdGw2JzbWFzuym+VzSPqhdJ5qxvKS
e6cD+wlV4F381xkLiFvO+tKYmcrUtFrf/lWF3vshEpCpohuL0LzlR3A6klEUOSxbDEm9CDKejuMc
15S6Fyc6KlncR0wj/rVqI66q3af4/N9Pjncyer1VxYg28YTC426F3V9tFUiGdh5MiTF7pN/wKMrf
Iq8+BSArXqPGXmlPWN89h1dUmTbbDh4Iu3ggNZ9IQBOoOQzwQxEfki81at4hIcL1QVT1ld3i3zPh
VSr3IDH1kxULOICO/GUkR1OIJEuTFmv67lQeJku1E3BcS6buVrttbsEcHLjVJQBhYwr8pg3E0i0I
GpETY5QfUFM7v+dJQKitOoEnKQkMkALS9BEJUGtVhc5QKoeHY4lldon7gK72lIC4AQtyc4drIK+n
DQywOPlKULfaOGCTe9bZXV3pHd/gXo4DoGp2ioGqwBNLgze4Hdj+GLqssCkG+hHXLwhsgDRovqTl
5hJ40R/HHhqxuHuKey6daUqVKiNxBm/yZQZyNKnUKkgNK3DyC1Ld7QWaoaOhXMgSKIoHG8bvx8uK
p52fVjOTw4WVzpfgi3T9X83a4i00wHP1iRw2mEh87s8NOWphkzxb0PeNR2hvr1TB/wWExNhP2cIg
A9N/HzPW9tT5k0wjcpj/RQaml2lgjkO/HW+pqejoCC+22Zden3WKOOG4bBk5HDEe2Wq2j+H/Zwi4
PV+8V1KfW2XtaKLVmsV+rYYQt7OLsB0ZQ6mWeQBeftpl35LYzXf16yuWnJM2IM2hsodiSu9W3Rnx
Nqj8iU/X6r2njffKb68uEUkGxPyYlR000nZ1qWAveg7+yMq30FuMlV6hdbjkPFv7QTy+5oUzd6um
KjTRVvi4KrY3f9cRZInjjEb3Wh+joVm71FPTooocEKhHgcanKP0nCmYbGugzUVcfem+dAwa0lk3x
iRoCCzy1/1FBrNJzhD5whkRC8H8KEfpZW0kfV9XQ3YF6Xt7pzi2T4SwKAnt3qVpvtHH/QmD2CLUl
o+q3X9Wxl2SkAd7rdvwDaBMoT3D6VlVrW2epPRb2WGFVfeQ6IMiWfEgRArXwIorVZql2yVYCQnRN
smo8LtK27bpldfyNZZiGDRhnaSLYsbn5uiWnDtPbTfLoz1Hxa0o5qxTmrI4qgTY05HTMI8ixhkXl
1oepBUjtEliw6e130Ng1vkS58SJv+PgWjd1LQWi7Q24Yiw+hDCyLsr51WQNASHtNSFaP2NA8PGS+
Fh9W6KVoUyYqoqvu9FUnsVfd0JpT3PWQNDYWM+7AAeDK/1kM5aSMRLbuqIeaE4zBqEY0ZqGjLeHA
oox54i0HpLmKetLg9fbB1vhGBBfCpEt2LzaMkBKfxVYPeXq8Tu8Q4bxsgGB5sLPetlDIlcYLAQ5g
3iAX38CZl5Wz3mJYSJsiLaxs79FKbausdhXxdewrLygfL3Hc0VjcpGwatiYUqsbhuBicynUq+Rsk
mKmBDMxU5Ke7xW2omoaQtQmv75jmp7Rb2PCXzBtUgM4vZ28CLzuQj9+V81/MU2K/Tq5+9XYHcG4g
BDp63H/A4j0JBPOwIfXDqM5MfLX0zF3ffCV7HS9UZPJ1RyNLyrnWqAxlOplSmOPMl2ys3KDv+Yom
jVCCASkPlIYyOw8eFZiTaSoWR53QwVIYDx88fgZg+AcNpgi7h+1FUZo0AWcDPgsELOGpYQrsmlFt
pysYj12SnkrqQ16zHPQWjCgDSdkLlzCGKH8IzD8iVYoJflZoLwl4SvPcY1ziYsKEM9IpCqIG6hNG
pZUPhEbLQcwSBODKe89wCvF2yMvT3VSvsm59zPfwKYES5tYNjwK+CseZelCY5qsyEg4KGcfUJaop
9OKcMeblIbJKp6oFXVbft4MyjSzmvpcRiTZUookp6XI9bk4HJIT07T5VmHkqDvSC1BqmAdPOGERX
HswFi01fsnIK+dYIrwPIksEIfc0Voych7ttM24mHlu+4wTwROo0g6TAmsNHBsLbQ/r/Fh68aybR3
p0ZZYoCGGm5S1KCKnkvNPS6SNBhJ1tmEH4NyE4PeeFCRLrsH6FcCtk/xNpWv4J4HPGuW9nHGDW8v
cT6LfRPCtzPE4bQurjOzwwID0YKG7h5Q3pW5tcR5mX3IVQDOYc1bgumg+9PsDcbrBY5JO78CEmbo
yJoKBDBf2SxEnsr+wCoC4Z9HBgWhKtjLkMJHOSRC5zlH7GRaGw63ynAeaZIXyL2UaGOcCXFzPOGc
Ge6xqYI2YOqV4biO40d8SrLfP8KxDGpXNdIKm3wt1I74tcamR12VetXsT8YYZvJsx78WkoYjJ8ag
aHlKYyQfs8A6wZ+LEP5rXI1n6os/vhvyYMz7uo1qUPXVcCHU21Ms6ijNbUGwnN39ZjdDCuF4fpSb
3shN97AnNsIDTF5mOxvWbj8T2VMTz+LeVuS6ntWz85SObLt7v0whzaZOuv+CXrdJpvvjFELrqZ5T
7N44//DWMMXR1lVJChjvyYSh0gwZo1M2GAF2QBhFvvSxBVw95j60S+6E5vP2cRZ3GrbxCrGQrQdl
dSGsB0E/li5TGMHu8xPfP6B2J+pYq6z2Lyw5P+F++LZ9cSLmT1LY/dAvSnvrg5Gc6iIvozC9pXPo
te01pOAKx7jA9rjpy6gDJTe3BKz1bZ4/EwLnTUvINPZEnOeDuEwHZKrtFj6WF5QuhyOT2/kxVZTx
d0qOlyL8eAXnRhxF/2hqzcwjK4FaK02k8LbAs97r0RcGnGNQ4tg8ID96CcqqBLuU4NXE7HiNxvh/
YBlBKa62I3zRm4zPNS+K2Cezhuy3kUm/NMs/dWHQRLETZXAoO1eNLVIxbwcuVfUCjd4WXsJxpf8P
FPUD7RqsvikXR03/rF7EKRw95h5fw3W7Rk6wKArk0gVK9M+7MP9ShGKC/LT+ZJ/4Uo+jzVH81O/r
NS68OL4H3wJor/jRVS5VA4NEJ1vjc8f2pCvptKFJ5UfcdvLwJ5Efnkhj00451z/aVkIBc8KieSoG
amXsfjmlAp+bdQXxe9X/m3jIJMRdnoUG1xD3LEwwGfZkuVTyVc28t/CVFBzsvXRfGYWspw11tglQ
+VWlHVm+ZzK1h3acdFthNTR7EaPO4DG57LRMoM583j28nogNswQGwufwyh/RyDCwbl5lyiCyohg9
DwmgN7o7OBIee2QshWhPgSymlJBAbCCDqYr3DOGwBcHvwULFPI0WwwkGkYTJrKVM6XveBHh0XSXD
BNRCoP6fONGlApkLgSKt6D0C4ZfLcKsmfGja4ny6W9/rY7QhcvTYRIIoHseInfiWBkTtjCmwsuXg
AglN02PIFcQz5F/O0GrmV5HzFTQkHJ5TAjG/QivrGACrz/1IRnSqq6Of0Rhhclx1aJgtzggXFTn+
tfxuZLLQ5/Ut/rEt8Lr2lHnla0/pGhpYTNDAY1NNNe+6zVUGO2tuqkG2vZu7T5D/TFxvFjfMKX8x
eNZT65AbDqZnMlY/aTegoKQy4+FohiO75Pi1EhOioLdZoAMnsc4Y0ebbpRedpWBJk2++H4R1AOgC
TeJ2QT8TNdsnpL/GSEiaxxzl7nOCHJwijlqhI+kw7cC1QCDR8jG7i/Up4JNXe7j2jcIcQnSqGnvX
coHbYAi9krP11oJtGBFnWmx9+R6aPp9l6SbTNauNV33GKjnStHzqJPS6/AqmV7zWg9gQURb40hcs
MiZAvZCZi/CWuC7sa8ZeGbcLTWcr4AB3MoAxPxiphIAKoKvvJ804x8ca4/CadhNjQlvz2jloc5nJ
YFSKw8WdjXW2VLpirpqQjBiyO8fLz+LgSjTWaA5geEq54HHIej9Ui+EEYTS2g52Z5rX16H9KUUqf
ozhqzTcpAt4CYWAJdlFe8w4FF3tWzutbWIBTjpRcdhxDjBrOI/3Y+SmiZEJ5moVGbU41gJyZ27we
nn1HocZYVzuA4dRAUMrL+49xG11lwFmcRSktNPS74a3hl0JNYQ57UWazBcP9x/FPxDGuFcxmnSvx
gzjo74kl3VCEX7hsss4ey/M/Kj+4L6bHe+bRA3WOC0GRgCD6wox3Euo70Wyy1aa5K8MxWMXPG0Gm
tCO9iNykSBzKaKCtLrI3U9QA+aJP2hU0Zq+5jKliqineDuSGJawoqlSmL3VhvMKhcrOjpi4NIGog
ic5+zWSOXNm+XnfwLUirynohTy/jm7Cv48wvUoN1WplqqjOGuaAfOO/PMx8o81i0V0W73ZjlKpiz
3mkiHxqtbvAetkxWbonqeYeWctBDWr9JOc3fFTtqVGCGY5GrUC3LxSiJcDYg/S/KbP4ig2we2DAW
wpdYV1gGNUq1KqbR91GGCnKi9clvqQ8zlJLv6JAXPtkpm0XxjT71gTBZjI9J3zOYdnnvF9m20n96
F4puAGGJT5aRw8yORfgAXfVK/TPvfo0wHeCrL7mZfkF6bZTeAWpQtXd/+uNlBAmA/nNGFNpg+2ic
t46Cd8sK/wt0WurR63hF1ZY1GMPtc02gJ8DHarPAU65s/Q+flS26SoRsbSr8uw2iQ5xKygwDFusp
LWQer+KjtyGmmLhmVH3H0qERwTBitY1eeLKDGQttS64gpmT+geOwtMKvX9SAhD5HBkZXlN9xMNKb
G4FO1Yibjpf2bwz04Jz34xHIKrOt4unCirMMgx4770Kp0IVi0ToQtQ9jIQ/uKlq8fRnSCPKyRwOP
ZbI0Lv8MaCwnk0oZoZGSJn5YvUMEsJO81I5IqdXyk7WzwI1o9zSknvv/BRCXUjQ/7hsdWFHreHDS
3tm+2JgziFQWeKLI/7/qGDrawUaWOYAZfn0O1nBvMAikKcPq7AnjxUyVQcHl+cvgd61Ggsobf5ra
FXyJfh9FASw/jiXu+XWqYu3n/RDQ1370KTHa1U22n0u/YHuccMTjGRoYE33D8f8jdLP78x/OEz/r
RSRFr0UqwbXvM4lzQYbbL+SwoYeBRohM/uh9YNOq3eKveWpEY2QVWLEf8jUEy/hsInPOWOFfqAj0
rFnXeEm9Xr+gN3oALaI5z6nixHj13Zc5DeT9rU8DWzfia4zogsgoIid0JQHUaRPzPOlvoLMBxsRq
oahqeFfl8nqvo7/ZmizmlFDHbnm5TZmejW1arOHGAxCmdDhgoOQNq8HHw49y3BlgMhaGoRY5G6L1
ExVWSC8LeAqC34BiTHf31A3GJc8u9enwUiVNyessVHJQycroM/if/PXqPkRDjY0J2comh7+y8NPG
VdSUwdthE1ioi91jscwe6tRQgQQJMvLb+6U4vXspXYLFon6d0j1J5ImAqcxZCCyEK5CijpyD7O7r
sbDXaPBO8yX56P8cNcwktiUW9SRsFLnlrWX2EBVU32pjkD2MEQgWiSVB4ywssh16tw9xk+/7/bIF
/IjZXwUSmRCEZMeMoK/VYA8/Do13oDm2FpcvI4ysyovD2fLd0lUg/AfejdEuUz1/lQBWAcmSxLeD
IBfdMPARiqxeO6CKh40YAuRZqsztqedHo0AA60Bj6hOA4G1FpypdnMvTQ/ZAjgKRu6XfzaSb3241
ojtTEFgbnVBvAxmLLnsEF7P3RxI2fQCB/gHwnwX7LWtr35xHja29iMv2x0keZeX1hO00j1FoLxfN
rQ1NEfFrh4h4ZbXzuX9liV/hEg96j5S5lOSM9rVULpDYaxVyAR8wp/C7+i3t7GrbyoDZsfKG2XfI
NaCmKcGP67Rq/K/5m62arEXIpZeuxTdekNAl85+bYrHXLbxwhISEEKMDuBazlW72Hw6YH1Dwa2oE
26bAP4sRcLnF0+64/wykkGmK23SKMV0kv9f2T53sEvnFUHWBnZacLzOH59/vsrM9qOWOojXAWKof
U9ZetK1jg2BvSpc8gYZQ63LRffCMs2nAqlOv6PuTS0d1Ap7jNKsTuoIKxbexubmiyDTu9HN5W+sK
TInqwc6U1t7pTWfZvVtj4k61hrmkbVJyQqrFJgwBJUrs3arbwGWNY6hNmpIRfLQ2HDvc9LWCc+6C
uQjwS2LnFRxUbi1IlmqUSzA/+2RlxryrHfq88+4MmGGdToTb7JUHgP56Lol3eKVWYvAuE+EWg+sg
WLWCNuxJ/oZvpmVLeWnES8CgBhQVvbKU/EUQ1e7ShYH4b10KZeoiL5zbEEbc+VdPjwSVu91RyD/Y
50zh+p4lrTTRZ4jVqzpV7Q+DhusVAJITi5XW5Lw5TR8YzF8/GTsMC6j+CON1qRpxweSjVXdG37Rl
hfEgpWSUfr3IyRVu93ybqJTfsLzUOCt/FwQpqxKkANnTx6sUbb5UrvUlMvqPxcnsb67QYg4dnWR1
qy1sYZVRFPLIqVuX2ygZLe+zW4kJx81XSSoSHeyoAALBXSWdCkOm+zajl48AM7W78EVeJl6CIZi1
Va18YWVY74WSHLEQOQT0aV/rmZjuCp3ywo0t1lKz6JyG4RpE2JC1yyFtWJXKQFLD7rd8HMT4xnqy
w+n4kQIMOEZA8kGkz1+HJgh1jZadGjpsJJCf3JcAylC/e7PGItnaCY3RGew/ijvD2reGZwzOSRIs
+m7CnfuP87oRn9KaMCbtx3HMnuRALHvk+CHLJ3JZPvkUeK6whXFa9Mt8y8qtxGeyv6K63Km6D/BC
iXIW2zawvEs9jjzDZQ0Tvob22Sqb2+j4zt70QKURriPLYo8Hqa8aVs7DM081UVyBYawW1LnX9NRG
130ncHby7t4tiFNcsGDVpG9gEUExXWcCqb39/TVwQzaUNQFnrO7zmQ8OTwkj1YXw7eK/ac67GRDx
ps5KtgmRs3dzsInnnOrR2j548FA3PZKYSQgZ2hJWSk9XafnyRqj606HOYGvkeZOjKa764KytFg7Q
9eC+wqFOdVdYDMcVVZOHUkMvGhI8A5s0oEp3K1Wnankd6rYsgc8Ldpgnar4XrBUcUHNKWIWAby2B
mzol5uCeAEtyOZUpNglP5IiITO2YPZbWNJ4JSx2AUGYcT9lRw2heGSSKDZVTsQH27FzOYD8Nl6cb
nrsPUpbRywfM5yKQsABVuQ6Gie9Z5b0LjUqYEUiEOyIQcZ7uEY52sLCumVIvnmH1Ysd6gwYDoprq
sJlvu3MKpVSWl1Ri9Bgv2DdfuGLsN2umyzk7s224ehcJ8SKmjlqbn7J4c5bADVmf8KtWKTrcTR5T
OYOIhfVxa3172hyQ06q30CHZYbZvN8jRKyNu9ySmA0hmp2FubWlj8TMm/uVMLeez4K+ijhaCgMwc
Ieg7XjDSF/ljXHFAbHlKnqCfMzy0nz7D5ueg/MeZxYLAP9fhd9e1FW1fC6NwM4q/OJEQvGghOKwy
HrGw6YDiwubi6Le7Y6jO0gR0ohQvnsBZdnN9QjMlh/NMenpooQ57bZmaEbIo7VZJCvZANODJSR9M
GGdhwpc9iBEccf1THfRTN4a6dJLtm3lXodwmB5u8yH+z+hOCsELgztN5acxFdDY4Zi6vJ6ltSMUA
kQKKDylNSAZ+3QWsikXzUrcew08ZSJBZqRE9DUKLRF0CTBKwEM0C1A08YCsWEYKyUJ2YeUEeOCII
bBMFK96UXQXeY92b4aJhXzDLFnG6aYYIp8LfL0JBuw37iTOC5BJPcporjXs9zGKjKMOjk1R6lrxB
iIzCivVILLO9hVbPVmZXHXhnH29dLed61sh3KaTmWNjtSMtd2KzQcEVk4FlzY2ms+k0++qRrYRxJ
S9oTSe2RDEVMpeIW6YkUThV8ecpIdwpDM9F75HZZj1FexdgHmDQBm1pcoHnPFVAFUq6huq5TYD8L
U8mYI5KUmZb6gEf70AWHUkzXXefGQDi8hZnCA2d9Vgr2ZFNXgRZL/5HellocOgwfj1RpEffp5qyO
uBdYWYn0eEHHLbZUC4xnVxfdMu141eKO49594UMf04YOAuhH8+rrzLuvx0LwowatJ0LP6c5qO4XF
E5RuInSCmsDASIzIVAa7nlKAhh+NbqV3sM4Dyga4b8a7pibbbd+kMTXIJb6SvZKxSx68GyeXGVrS
63y/iJG8HhesqeRT9PuO+S1MDPqYnFav1rUNv3WdC0aMs4Flj4Y+GZFHc5XH+oVlwD+0lXpEX5P+
/jkOSMThrAm4j0QmgdrDTi53UbnEqMlc+9//WELVNmbfC40HTTM8GjW5qWLK4YMm+U8I5NaLdG/4
WuvPVNzTvVTnN1Rjv/Tay072/C7+XVUtUJEOu4tw+Qt9pZNnb08oXiJmQiRpVGdWV23rvGPLfdB4
pn6qO6ohPOGpnP3Wt4GGUjaaiEMZ7VMpsQE1Hx+0ROo4lOtsqUFDJPiXFpb+RkkM6bfT7cr4Qsee
C+sLKjFrdTzJWkeID/na8CoNLP2VaIcPxae48r0fdKFePkoWRB2FTvANhniixIX41iFkG28yJ39B
mB/SNSt8rrS25/heLVtQcZzk6OdZdaQDNbfo6ktEdsTHhEf270KiC2GDiLH8WCF7ozGym/yAq/xe
TaNbDZpJhF/Yp7uI58joLip9zaceoOFf4SyIxqFN1c9a54OlHRc9gdhibJPpNIZX/dyujxVDfNGM
cOfqvlvQUBSv9XlZvNuMCpQY/Cgn+CkXuMnT7ETLGTwHYhQlcmXeoOEITb8OPzKEJYvPvqYcZC6a
uvLejQl0X67ES8+NEBq4Lo0IkebmPIpJ+evmYVw8o9aSFL9hJkqlj3AkMQIOFZvaiFuEohMk9ACB
idQUiaCFmCLD6ZzHafx2r8boxAaSo5jk1MxHBb7O7s9wUzJybRyKAmH/0bWRETCkVTZQ8xXIGV8l
+Wcn671wjJWRDZ1QB/X5+FS3WAJcLYDgZzCbhLfq3tRwOoxHryxlESanEIab1p7Tp1v6IEl7bgsJ
p2bmKCEBosmPAhJCwm6AxbkVy2SZvgvZwLwlasgzvo0/PGIVaaGZYRdEIdGvcIafNXT7oN/FCa6c
lUjP7DMEov6We1MwWetPExlZcKUf66cGZDRXBe1qCw6t39vjxx60A+7+mjJtJMg9/9Gf9vrQSAZM
Y6yW2Va2TFLkoHgMiDJPXGxX3e3jyzpQlBfkJlgO9GE1b9n+JrgRpUWitDkvmyfZR/Hpw2mPx4Ub
lV2fcVWWHS2nR2zIggmNbwcLCb1hJnUIOLjREbj0vmMQqhuFOfL4DdKwI4/iEDRTjeTT9XSvrDKH
+kza0NUEVtGvRmehpARk0B72kGFJe9PfFMU7byjANSTexB640DXDoayXnZza6HcjH5co0/nicA44
wHWjlNF+5EoAYEcCFgeShklu1o1fqtZ8yTa/Yfn/3VPQXkGfMXPmHKrkJ3E9CULVqBfMfuiIaK2M
Nv7e01DSQ4CoLAGIW9yotyuVe0O/cZ0aUJqvhXsQSUNH9+FZypGMc7uD8HmtBPHflQ0t3x0Yx3A1
0/zG50iJ+oDREkIB13OFG+XpyNAKPVHByvE49ff/gi76LUrpdiF64R3zRVlve2av4ltZut+c7rwS
w7ksI1jZx2TuO8QuLAhqdXVtgmTakKe1Y1VfqC2A48VWKWGALRPCEqLb0qNk3jMQsInvF2Qg9CVF
FquS88HGMD1Szk9u2KayBma1MQMupoXxc53XTAZLL5pZbiwyKw+u7Nh7/Yi/xlU2fYh+HsfX/BoA
GFTSAQXfh/tJ+i7V8ESeQEp28cnWUsU8zT9qVzhRTsskxM/0pK4HOgRelivVi62/mOEG7HCymEET
pLyQNEsgPNQdJ2bZxQJbqxj/JE1CJ3+zIbP+mrg0bYP59zn1g41bGvj6ouNGitvO9mXG+O+JkT6T
aty3hF/grZxz/WKIoUyXTyGBZrROmPnUhJ6N0QwyT/uauZiUQXy3G893dWfUQADwk3vZcCQN4OfZ
Qx2Rp31BFPx0x6/3aawmEW4LUseqkr7H0Xwp0mW5TkXVYTlKZxySoADkvzWSwPNYwHfd9upA3Jik
usynQYYGxZFCIWYKhqVqsqSQyGA0lbK/L+IUZ1mS9tM4vhVAUdRfoMU931BL/J/J7DIdNwpNZLav
v5Cj2+lGYlToXjnzCWI76bD4HsP+iurRF0VUR9/L39DqvmzRZPIIF+i2mW4M5G8XqHrweUGmDoy6
xq4u4jWs8dINhOxTlVBKD4OKiYhBjJHBzD0MyFoerv4JG01ftClBi27aajVHaiCHlx+CAAN+AGnX
tEz7AGgtq6pdGeIW42wDWnCMBRKz4gaZH45OtmDdMVz8lYO8WS/hwdXu5m12E2OM7LwgDL3H9IXP
3n1Tg44HKA0rxkdV4kbDT4oU3wAuPMKzTE77MzYLeeRbjF1nG2YKNJfTonIBQQC06XONavV1wr/n
jXbkY3VQ+Czc8wyWZYlTafMKF0lSXo0BxW8wWGBkb6jPV2mRFUGjQYHN09IfpovK8wFeEm20fWKZ
5+5OiaDp5Ohr2VB3UmnF2+DpEZB6mkvUadsLx13UpIqHJUuoA6KjoMr3gncDLKZ6M5MCvIyGJntf
l5BEzdZCJBejoJpAF5ClbAOkqAm0N3h33xR0NbzPHFpaalLvaboGgl235evbXszznGqOtctBqXJI
6Z+hJ6L6UonlCQRmiaS41tpxlvCcqleLrGS7UVQMUqhl0csZWJdVmCboKCgavx3GTxN6N2lmFMux
AOa1SPI+89QY/ErBlNtC/HxwEryrKQ0VfLaF9j3mdJUol5rfRUgVHJsywUxiMsIdprpaaQSFBFbT
GuAy4FL5p8IALzxKO5GRQ0bK/AbGm2GTjp0TeWU/X2TWPhMksDe7AIij9/VqG8J/Sv618FuHOWUn
8LUXy3eU4/MqLf2xfmnvWYjyC3Zt2EAili/9u0f4bnNPHxIy1zCKewP+MMPptKnMIxqwfWpmksPR
zjen4jPzKtFEj9CRyvFdhdq+lQb8O+PArrAREUaFTNzcmOmCb4CBiyfaWdY1u7hzoz08PswzRO3w
xX4udPZMGQmdizaPIcJt/lWd/HTyceNv0Ex14uR0GueYVJbty3C++guu6M0T4pWFtAhVNXqoTlAz
ORFHrLbDZrxf96o2OzyluhFgDN5Boz9He+p5vrwRt1qgLfvWQfTAYJFpBKGpun23xusWOc6YL+ae
0oJfxM+C7QsC/HZ6FBTDChyElTmz6MGt7D3VwZf9Nsmvv/ulAMVmeyuzU3BImNAfIvNsMJ1SYH+J
GuoYu6Xe/CFouFhlMkaqRXIhsABKICr9OY10I4ssJGC553Rn/ogZi0z1zgCoEgw25Z1qrCKdmOq4
GaBAp6bLydTV2EVtJX4c3V20vCuKT+p7R40gJ6JchSEI9+jAJhM7opL/wjPMX51Meq3OXVnu6j5C
CRY70GAi9aDs25RncohInrueC1+DjIHIDkxl69aycUD11xlnWOK/k2Asve8nJGWgZo1NZwJ+mNU2
udPyuZtSf4Nmlv5q7b1s2SfDB+KqrD1WG/IIj8FV1KuiX75iouPrlrzALMSl4kqHFYUd1pEDAah0
Nvc7SCJW/GV48+WANV7qcc0ED0lk77T/mUHXOkuNYOpIniyP+Y7YGdescc/9v7EtSBx1OVlWQU7+
nWBdlr/Dvahnb2A1kwyC96dC0HnzCHegS2RkJnWSQA/T9VFumBPsIkEWz6k4/a0ewhPD36Yj2Sn1
oSFLcqvo3VTETtUhJkrFcOAiIPC5SJFGIeIEo6PzBk1NgO/2+wdp1ySZqBGHtPbY61wXOAI4lXUF
bSUs7xehxVgl/jwJEvm4j4X6jPRGbQcExjeUPBFxtZynsN2LheON5J+IWeILBy2pEzk68Sc6TyE3
X9wH/vxBcOAhTZydnyEoAkZUkjp95S4s2NLwTshMvK9WVWdlLknai4j8xkhnH4pgtU4EFDIx49rI
rieDuUZEDhN4/IIbX9/O2zHPTNWS+RmR+yaUyJ7Om9TewZSGQeRkNJWSgctl3GNi7/TU284gdkTt
h/f9g2SehVwy5peEwLCHUtH8A/vFIdi7Y+6Y6dz6tRhXDIPCpcUuoGeJ5BesMVWNcmxZMG3pDWx8
pFvnP2JuHpObykvn2/tyd9ra6qn1pvrUIRy7q7+hRq4BfEUqIDWl34iTeRw8781B2y6tH8NuTkPA
zV+BqHA7gfQZbxy6YAsLSTKGrIVw443De7PWHBV/rnOhvbzZd+Zn1pW5WFrGwSsq0Mlmj8N/XiE5
BOXt17bq3xRoayfFFrgDUAhYljBH4MblLZHOcu60bwHhZNtKE6smg8AcFGZ11pighN2PwCtBx80D
s5encUPWBv0JpOnmPCdF/DMAQXkZEoKpMTr8N0TfagN3G8tkQNMmzrmYcceqP0yWp/orq5Z7H+3C
aBqDWFQmgdwYClh1nm0IX+bMoB5q9Hwd17bUeRblh3Jv48xsuIuUEZ/dxzr7SsPzLlxO8y1V89gu
Vu2BCTefrFXkPTt5YweGLFZsMvfFe/TpmMpK6+N2kni//GqfLOM2s0zlyGRrddouJW4cQ5wZCKKE
mDDmlu/lqiNO4Gi5q6TRO2FroLdfB2jgIQBtSEygV3NvbG8BYgA7PPBGsW/gu2Rw1x3T5e+NVzyT
UvGmaxU8MBJhijte7YomgR/5JB1X9exwkjxk7DDRl1zG8kPcbCx5relbbBD2zuPHVm3JJN0JCe+d
nYXcV2HP13eMKX4+I9Xyu2CcPaSDcAxJL0kpoCbT7uaA/QvnvhTiShQ+F29QwhFH9fn/j61kLQFb
WQT6ln8N2N3/KunKYkyJX+rxiFIIIRvbh6DqpB/k3W8byZMdmhkmDwzayivbEQWHsflu6cCZ5NHS
VkwS5ibCMIyySC09BvHSy0SVrrz4k5vZpcTrpcXIbKI7HyvxC6wtSbPTbV4c5a02XHReU88Gl0Fx
YBhfJzpyNAR3oITz8LYS3i1tOnnyeMkaDvRvKtpWb2Xr7VPl4kro7oFTFQC/sZvu4trLgoxfpyY7
7UqqkibErJ6efjJnIzX/ueGgFCpwj4+AdLIYBW4ANxB56WjbFXc+iZl7UFW85O4q8Imt6aN1oHo5
ZnHe3WUto3ghb00XJ0cNgEURAbr37ny7DBtrlrzuqvPMm4YEm99hQd0PXujxD7urUIaE+PzpNxU6
ghnygzxxKSyoWh6Y6l1dIs++htou10iyd1ke81gRqFXx39M4vRIhJtq6OzuzfTU+yeXsI3lzjYlu
vXwwsccIBNTs/eRWOcaLEg6ZJjDsPC9KVYmgifzLlxLexKJ2xKtVl4YfFk3p99YYPxG7+16jODmc
kwxXjqDUloVIidcKRm6tetxLr0zIggN1jxxeflaQNPe4Bu2D7qX7svvMc7NRXJqUFSJpaFQEBcCe
gR+KYNRKZ97jPtLR/SR1UEQz2ki2DIkCyhv42Wo9lpOSiPz3oRIWtejIz7MWuZ2ZDzABcNoWvngc
mG0La5PgS8lcgbWrKCnJR4LzqoY6tb7eM4WUws1QaghY0ICFIaF8vLoABh92UmZCf2hT83h9/P87
F90fdSEGX5NJXsWI1d2zpq3wTZoddeX9qKiuc0oqRaeTVIpojNfHP8+iJJaKPjTIhJEaKokX6HHZ
6H0Eb7QbONUBC1b+51Dfhby0u1xFXve1Fr++92Fq2mdvQI2Z1V94teNMWuglAhFeF0efC1NVS4no
vpxEIP0csjSMoPZepJIW2FEcqNy58LX/mh9PR6y8UotiPFP+Hgx+wPh8DFbDAA30NFKNlg28Vv6E
l9Sk4wzqSZ+sh+Z8Tm6d3ntDWqM37VH3x1tJ3xTxIdnxLufcXybiglZRng0BkFa5b0VsAapzwqaM
kPmGG01sjYUByyMiThnEdvrKxm9CfBVpG/kuf2WV17SuvE4tqU4/bmVdI2JngLUSvABdcNt0HyQS
0VyWKXSeVuq1ipJympZN9cMlaA0hTcRLMWue6I2tib8nUbAY8GA2pMHcZHwZHnQQ22Xo2jWx92wm
nXdsAqxKk9sLgh15bOwiEOwenQjIksbb12b1FmD1c4CUKxDI63u7nGIN/QHeccJyeVFWfl/PUdBs
GFLca1WutCbKJBZIEwsxcV8HbivZP1RaH8zaRT1tuAOzfDsOQc+GsHEDuBPZiZebfVIYt0NuDlEz
KoXaSO8t1hWJxgtKrxftvhc3T6ouTYjFb36KhhocYGW/+fWvSZQ5xLMpwabCOpNQrxl9Bnxphs7U
TVO6CoKPEQgH5J9JB+OIqe1pzvkhyavRZFEhhnddhUxjOSjU+YgOPbdO0jeYUxYzzcUKwOZCsXHu
uAiZmixSxiNwKqoH48JWbu+XVPQvSBEREoDModZlvHKQdquiAc6dRlBmefhKqJrs964I6EgFOsxj
RtoVeQdcg8mEuN1sm5Ec9NEpCBtJR+Xrv31lyrj7bzgu5gL6RGgHidh3yeHkTTtehol8/0ZTdmyd
lzGf8FRCe23bi6PZuJu8pr69DrkWjRq4JcI3xKybPJ8p/7iko/h/W25RpOJ5PepEmPwkII2N/dd6
yJhLId+acpiaUt6jWySRc0xUXroIj3/lS0n1OLsf4FKPv/l4NJsTl3VoAHBHnzrKPVk3VEHg0EID
VWQiWa+CwS9clgABlW74pd5L99i2vlur82Lv+vkp9U2lpIMWEVrH5sZdI+k/mbaHToe94ACuKQCZ
WRPJWMgW/sxsleM7Kdn3ar+Q1fmmQ6T/xNHNZ2R8Dys6D/fBuW1z0rW5Qp+JJdKw9IbpfqLp2BLF
mm7YdeovhhKsX2sq+2j+q6tXpDXUnvGlLxTNxkIF8WHwWnK5G/xmz/A3ghfYF0zyrIL/QxHILTVe
MzVir/4V0uBPa4Ivz72bbGB+K4iIDK0B9yzQCqnxe1J3PzuA0OCt2AmhffIyhsoSudJ16AxBYR09
GdBioutMLVU07XjK6JBLdB6fSu8kunjwZ3UuQBJIKoLCKzCthl35n8//HlTsdDQUjWGv/8ph8sED
9FtEwMLykYwibWygeuUL4JKPW7orMYGJ8rM6xd+BH3RX0cGrkhgzG9BNs5Rt9NQfn6wKq+mdaUqN
pIOBvosAqqi1umFboYAGAXktCFo+fPJThJ5CJjJTBbNWeMngFCrLw/5ukrfANhaMIMdCEIgs3KFl
wdVfwGQEm1B+DQq0lFXS9Ejj0yDm5KHlWo71wAC1bH8G9Nh0CGqy2IkgDZRSSNhA9XFJcUp2Zckd
YtepdX9YGWLcyxdTdkdb+pj/wYdaxxaVNMmB4C1AE/nXwI2ps/23rF1v9czXErYKQEOxpiH3Zr4R
C8KiuPUlGVHvZPDLhXkGv4qxgK+X1u6oOb5a2DCyGLvP7YuO4My622E8oDe+SzzjvdnhkLuMPE6Z
sZFhq5ovJxsvK3mgDY9HRXXy/i31TIPkn0DUZv5wNBnr+6EellqgE5L53sTuJ3Zn90cigw7T0DTY
L7+CAsFPPqKW2OjsNUvqciYInJ+VAq0OTaRZ9VdZ/Ejq3XCBQiYMfY3Ad/c3cZxZ7kATt/P+I7y7
ohGdqr1hoZQMJNQEE/X5zdE+YaMxtTwFQCBxUuR8yiGZweXso64Le27PW1NNlpsZa8ewaB5Q1Bag
xavF/Ur+CiV+kS4KGwOb9Ubi0r4VZBEpPOFGCo+slqLgPJVgw9cVo1dMA4LZUnAwLCbPY9dgvmZo
GgurVS9Q1iamg/9U3gCdDIk8xgUMwq/tcrLCw/Fl6AmqL7clUkeEIxPwt8//ZGXIEb+DNKwmO1eM
UO1Nc6X2y3GGZbzCWvkGPyTqRKTUqvq11zXfu1LvvrMP1MkxUxwBTV0bj710z+HlLbE2VLtZvtmn
jtPhboYNdLR500iXjZ1HNtV+Mwk2J4tGOpX6zoEEmxTjQQsnTQfLsLxSZeDr9B/WLs87OfHxPK4+
Ldt8yfP/9N0FEHo6y3tATdd3gSxqlGgKtUNTE7aLdspV+YIpdIEdqw6QGKm51xaqZYDhr5mUKKFz
BR6Gt4dZHEJGjdwibpO/bbCWnTMX2c7cORsML1/NYLo/KH+teu8ltPTRbuzW+ozpZ8DtFXfvyI58
IWYZbigalwARsRPfsGG/2TI4zV+VqjzjVthFGydmjH+rJQX4t+E9xtclxEdZJqZxG1D/N0VxW68C
tm0Onpd8niBPHl4nOFAOjANP87lBfYcHcw5EamhzIRM7KcpaICNo+s2vAURyLY8xcVFq6lNs2E8k
6UbJ/PvLzUntNko0RhYb7JRIIJeCQg7ZQru8+cEbNVD7cprTEBrYQ1n42hmVqPDVb/aELmwCD7kB
+W2qi61V4NvdyATCoAR+Cr7jsxMVkFX+St0mWZfAdzEFWOUIuSZ+ztvg4IPPxJQ0u3w3cgXfPoTc
AuCQBSTIAMvUIvnua5MlFEf2M90jbDcSd6YxFaVd7rEaVGQqZdbduSpxn2wgCNDBcw+GhxztJwy2
Yu5guoiBnksF946lbBHXvT9lP8LkX0DBecXT1HMNhW9Tin8P+EkgpqEwINh92lecrCS7wEomX9KM
cyZcBDEUJH5RSoEsoXcHM2Yin9pitUQkR8ctgalSRSRypKL6sHzUOF7vKRLdlNBhFLia/UK24pci
TZtC2b31Q8Dp8JVQYoTaZbM6d1xnIxeDsDu6tmNW6EvQljRzMz51kbCkCw45xv0Zq792bktKKFil
DaEMEuelPMpAMhsBTWDASMCixXgdu9YBoxLpQe8X3wDxa6mLk8DXlZpMpHB5lhQ8yeYkRSa/VbFo
ceLBU8ckaU4gT4yR7V7YHspNZJCY7ObIBNOXbnpQ3qPS40GBStj2efqrNj9wcfyn1CrUfeS68CQl
au0HifIj6W7XV5vpq2YuleZTqfF05Zuw2Yc3Cwf2qQtOlGV7bbIJpbNqN6cmDEz9dXnfDoMDyGdf
x+YSyCIzF/fSFhiGSbev3rTOfTqdmYtcA5eBCbt9y5nRU34B5kjxnL3nN02BU9ZewJknM20pwn4H
m18IvsIL7ue6mUceATcfw1Lkhs94PSk91bgzMRZh4mZloaf30abQMOEtixk1aFvHk6ZzOqhqgrjU
SAomTmY/bsnpmfSHC7Pwhb1ekGvfGRIQgnyI+LOEjquS91ltiwjpzxLKRhlYjkQc8E97uX3SkFiQ
gJkfiSkt0Hjn0K3+C8bRLtMU4TgkqJ/92dNH/2A5XLZ52X/vQOVGvCqKD6CpMqsiD6MmMe291D6h
Xw5Mxc2oITYelXvTO7rlEhWiBF7Vof4z0i0IbfIpwBFvBSnmUg4Us8nbCZvNqUlTujoWAHhBq6KU
aKGZlR4Wry4jM74Orcm+Mb95X/e6CC2XxrDbT+jlKC56hqTMTRa1c2MMUUbC9SGArtfc1Cc5ylO6
px8TquZMAT4E8Ajf855HmgPPHNF5j8nXDaaPdkXPUfoHQPZzwdZc/i8R1PnwKet3dXHYYK4UHeR8
7SpMo6Fef9kY8XmAow+MbyZrNLtGTzPi/rlUMax0/KnARdDwoWA808E4krPz6KfQfSKrSmXhMdUf
ksx/inWvdkVmZmMV0QyfI42JgOOAP06grLVm44ur1cNA2NZ2x5PoDq6QLgIBjOAsOf5djI5JepbU
2MGEkZ8lFhLvaKjYhIvh9WUSXkQgkDXjgSnX2v/Upy69UaF9anE3xqFg45vCwV5/+F0QvfnWlbAj
ABfHMlAdjM2D9Fk0BYsziFdTr7oLy5B56/DHhucWf6aB9hCDZIKD3b3tOuf9ONXZ0JzK04JJbjD1
OC2KESuv9OpKMpgxge64UY9OWrlGDgdPL907IRaOwBqFcxhsWJvce6SjkjxuMJZKTG02k4MnYOQA
qpzFcHSeTrxPHQFcw2wN4qat6PsqbBY6jX4/zjT91hC6floUVBm1FDQXE10+yvOcOWB4HHt5eTw7
CZxjzXncJZ5cw1VTD2U29NA+dbPLtg2dXFXq1Yqe7KE4yFjJDefwDqk1xIBtCn1Scg3FHS1k0bNY
kdt2j/6JZep6Bdy4zoJ5TBPm/wriMoXGTIhwp0vvAVJ0U+2IsO/4kFW62s0/JQy3mKoXhV89nCuw
/hAhPkepqX+uDSW1mvVfrSYNqTTvOeJlMG3NISmP2LPt/8Lc2QCyoZPV2VI7wSx6JhjCPJcYU6gN
q+G8MiuSLY+PI4UYq2i59tAl9fzabwCmxdzrluDb6g1+wmgpA93Od08W8U9F25hxptmc6cy5jF4u
5E4MLobO4wFNxlPJ5wcqYtw6fnfd+tIo+I4FSbwXhrs9kP4pL/J7Vn7uoA2fc0oLPDHJaAvAPxWd
F3SCgj4eOVcwO+whRy2ipVwc4jsp0X2YKKmYXzTGIkuu35g4P+QTXik03hgtjtFpkKuGsxa+djDi
DoFSMlDBlkYlWHgRLy2IMdggedLgnlMHzdYDDfYf6J2E0zRzzWyJLRnCLr4B6gtCy/gVbpcdQyQZ
8W3mw1rdxm7aLjAcEl6RXuWE4lPgMp/mIf+uxT/5aoAG4eBDxPpkM/jiiAawbPiIvUkgZI4HRhvq
COzJ0uteE0W+AyWNaL5sYz6f6c/9Bc0fTHc4k8GBZ6E3RTp866vcDuzJp7ctyXe/+GHpBA4CUYWf
axBNyV1X9l7iGPpK0mJ5VQUkqU2A4XJ7p8SlTmxd3Tx+HFBPINXfAIF7SaYRUsgmcPws3IYaCT9F
Tlfmz72pKsA9Cg7ikN27VozKSxz04hs+7POL0ew3wtrQ7jhOn87awPcFhkpWDBMEleHaBOUNAm5O
jtqkuEvjHMMEA4gAA65GDjHDS0JirrHvR7V2czKDpTB4zRa1JHps9aOlJAR0v5uTrydUdAjGUDVV
NNyVfl5ZPN65WeeRbyq998ZJs1PYiC16DINN95ZEoPYD6naEJJduCV3ZCBcXOm36Oi3ClkbUII4T
ZX8GOvqny/fx5JMgFuFMmzL8kiT8SM3M3tMSnpvjhsiBwHJFVx5Zfe2cIAkF/mwHVoEYor9c+dmH
Lm96AaNeO8lWwAXYjRat38mWgD6qDl1/GyLOgBbeA+gWttr9wlsiiuSPi7LxRbQ0k1iDWir9Z//3
VJMJsTgDFPBUW+yzi889BHR2JRBVRgoYL3YTJtW9bESAA4SYMmnfVuhHYVjCU3Aj9hQQTH3j9E0G
CfC1WifGwk14Ssc8H1NyvQBXHUUQH6aYFzYDTHtFteGI9weIcSPnXJt6BT3lf97VLLQZS9H/btix
+piZIue4WJEQ7VyYtfo6GF2hLUFoM0gCphcOYCTjNdUBJPQnGreyrq9O9Iavtgc+xCyVEzZf4GWv
dWFXtLMCvL0w5sXGI/XOvFr+BNxU/YhUvfNyfL0b6AfjCi4OCx5uLITnPmtdvroz1ZvmkJiS+GpS
D/4PZmDK6pQ/e5q3xl/Or5rHkgu1fT9dj9iXpPKbA2ZYMqMtfqSg2IvFjaKiZEMyV26TITjbMkjP
hW8XVj1UjHH2aSf9jE92aDg0H3yK7U2mlyB8vtnHXvQXXZoCOLUgBKlQLYzBuEWYLQF5zZ9I6xdD
7OqexK84fZxwedmebJi9qAI0Oh+PFuJVAsbW2OrPz0YTHdiGXyJRcozfcu6peI2uDyT3R+L07OOi
L7br8XtBx9VQKSiLlNgZ28IsyE7Yi/SrPV08xp5sSTS9rjsmqEO6x5Q1FsRsrLOv7QCQN8K/Aghl
PB8jLVZqGxg/MSnl8xlxmMypgnYFY8/uqXcEReiY7deeH42xeRKQCqPDLQdCcsNUD02eZjgLHnYA
AKWJgNVlcRehnfbi9tAcJ0UBpIwwfJFkArqA84ptiwm8x3D03n1iI7HLMVOm/QOKDTMBnfOguBWA
5M1y36HtS3qjnyARmaL7D5nmZRyyi1mqJHnHOcYsgQH2uzwHf/LqR5tC2FVMffy2Un6xdVBOdP0d
ksHz/guGQhSTN+cqGRe68zK1wJ6SRUiNJJ4Fi2mkThVfp71+sL7yjS469CDRF8CUwKRflD6NyH9u
lI654dhYlaRuRq/1uIfccT3SHJKe1EqnHP7bk9Zd1JAX55Gksx30FhENKhR13riZ09sV3vgJOKws
cXeA5exv6ZVoMIx3Y6ls5vuoF7vAHt3RPlSYJ8KUTeMbJjXdCfdX0pwkINzMHt4jtsJ0jlJj50a0
8BpsRJTNvvuCcjTbS76whjJ51g1fFIWA+7KAslTfBi/G5YI7D8fTgB32FtkBhTyYUNnM+KpEptrd
2w6oJKB0QG7hoFal2tDpB0pZ1Ox0cMUJn14C0oG35CXKaZdL30wPIO/un/OAUY7MuY9l63SEseBV
u9gqGh2/NU317XG8FluTOBpaUxyXzoL/bsjHZ1HVnxT8M6TtpGzSkBsocb8H/2aF7B91QVHBix/E
CMuIlomDjCXiKljCtUVs6YCvY2zzSJG7+SC6F8P6+cdsh/UD03zs+CcyyLSbRoPcmqNgs/1F3T1i
Has2OND7TQ8nNf50e2WqR2QQ3mtU0p2LXpQshL0tXbTqeO+6UtMPnEPL3eRyYM8aRSXqwOOwyiQH
2lPRuPyctKp/IpNB+pZ6uF70ML6qJzHua/MMoNAxyyqayQPljhnyhX9x+CdmcKedPfXX/zXMxs2E
Sy0y/lSXq2zH78xv2IXJcHm+QOSMj3M0TJYODh2QwdAoJXIOdPt+jSSj+jmQPICtn1gdVDEH/oYa
IPuo6fC9Jjs9qggeMOCPFPgzr/PRCgdbH6WzbyAEigGLkkiHyGgoAgWI7UOBXsfbru5FjFPQbOR4
SvqzKiXcBfVnqdxPVm2IZCgc/+uvc09m6vliHaBjyrIPIrkihRs7yDHe3OXkJ6pNL0zhPlfBzREB
ilGhatDWGnDqf0Hx/4xgw58KtiGFVvd/qMXIUKLLW+Bf2U5iMAN/SrYcfnaklzjXtwVoy+KDMqYj
PEwf9df2cWTl8uGk/Zn/adP1j5DHwsL3dR506dVSPDBrABABJ1JJsDeeyozHX0gGajdpHGc8USGM
P5rFWH0u0G7lkWd305ftJi0GGvSzubAFmWXFuDSnVUXwC/o0AhJLHPya0/ZSPW6xdnzP3qQLZLtM
xI3u0zhDR4SlQ+8Lh5Iil8P1vFZPbgvhx+CvTH7vShpXItexnKDGQ7ChhJ0RGW5H9RrUFXqdkDlH
AuUOnDGni5canvevQMYO4nX1a4Bob9kQUTsAr5aBDCXY0bMUfElYWrHM9ZSGdN5nMPZWwLnS5FyG
Ft+E6bfRi2N63pnGoKUYrO/Lzw0E/XBgtAckLSC3ed+4e5oB4gI9h2uLR2GdI7STmrRwDu13YxZZ
vQiMcPftGt8WWRDYxdTVYOZt+XaiKxwyTz03l0Y0QqETwlbsPnwfPShnHhMhZoCQXDwn7tY8lci4
CVtECRFL3YvGebpp02D+sirKU9F8CPKVcSuKEWySDXD9ZGsZjQOJTBBYySfk4ERZL7/p2XE7TQxR
WMMfJa8ohwqgPkNm5z4IMS/OunkHwLJac+oq/U7GVXKatFJlGPIAWpSh1eMqPqo62MH19fxyT9KZ
bxVZ1DnWuGgF5qZ47Re+Kw1nB0h/tZxpzD4RgzBfX7sqsWAXx5Cx+HTf2T3MZxsZSGb6hphcLx9n
MED9AWrAHCMrQlvLU7br9Szvm3vJoMWA/75Vs7L9vJKjFSupzb7Aa11QvVNOmkIVAXZHvb3ySAYE
6dMkv31B/lGl1TmsiHI3N0qh4jJB9YAtekS3sbMGqPy4IvZU682+I8j1DmyQmJZBJ6YvYXq8Xg6o
DWHghvxc6+hbaWeJCkcrcWGZaXPqWDsFhg+AZTbehoLIlVBHDEGXk4k23oXpGg+U6xjeIuBXzwIb
XWermCyW8OEZWrejtrvSiDWWv2izzr9wyvBAxHlQ/aHaUFFkLviI7RY3LGPsSoJIDUvWi961jmx9
+sQG99nxhvUeF5nizzj0PaQ63p81KGtXgfKdYsGmcPk+GInzRXmraEo70PRELwP8OwWVgmrMqigC
aKPJAzA7f6N7uTMnTlG6dQZFtJ3lH7u4b2JxbKNClg765y9SoKCOu6oWW1BdVtgB76y3yMX4J95+
KawK/ZBJ8IQQrC5TC+aY9rYreOIxWXrCSe29HQjVjQhC9ylXPFZfDVo15Ut1GTliDR7WlZSO2Ryu
DRC6dVfIPAMxQhsc9C/TrOfjZQD4gqvh7Sw/LatM7hqXm5EzrjEiv59kmz7i45yXKD9RK4TIdlmH
p0iEWVzXiNrMirS0PTIayp7x+w13iqHLKw/fCfMko/WhHW5YDp4Z011JETlcExCgmR6ON265+Fyt
NWQx4na32XVx8FdCPoQeUwNdks8WUm38osyIcR44lel0nmoZqNTH7p11fWX+RCg/xPD1eTCYxqPK
FOaH1SYiLSownyoWObjxqz3n0c9lRplboxDI+xinSHBn4RJn09JmIQYV61oPySjlZtJ0wpAwfkKf
SM0ve9qIz+hgNzldR/75BVa9i6ciVG9hftuEUEgZrEoK4Xq0n7l1Mx66X1SFP88FcgvKAoVHbuCU
om0cYwh+MLKCxB/WcQWI1gGbJnDj5kQDKk+LqPwPCSmrGgb21f0oxsl+XYKFWyNsX0uC1vYohyjY
qDTeR3h0FGdEtFRF/HL42ZPv+HIdJFMxuURmjUzxai5Rcy1tOeTNoU6r+qHPSQzdzdSKh9Mq9Etd
CaIj4FBvTYPFlxoSD8zmZyTGeUv5WEXLFeMGgUUhut6Ha5YlRX8F2nQuIW4x3aEPAgsUFkYeayLH
0qUURMq1WrsiVZUiHdr6V9M/UlcmyLXDPR6eWHKWFT2oKjkdjwoEgyPbx3Hsrmo+I3WjHsI3NSQx
WNkjruWDUJOWruMB8seGI5yq0iNjDRYwz1v/SjDxiEpVNprssUGZCGTa6IYCvKH6tYjG33bpcEKj
HZZNdwFs0HIhee7TIyxGit0jk7QffjzoT5anVN7ong9/rqvSRavHMK7qzK684okOT5fcM7GJ5nYE
SK5oyx0azeKhGGgsjoEO6kSqKpm2ngxwr++ae8WWKbxNQRQCrTQE9u6wteZ/xs8JspgSg9BUtVC5
cQZKWpsU2HcQuZwecb0C1bHPQTPIqz/xlo06CMNyBqiDgr8ov6ZV8bLj3962YkMppIgqKcssR3Nr
d7IkNlzMLyTkUAJRIa4i6BCTyrbNp31nEyckqMWIdypa7Dg2zqjhq3kh4+lDOS3OmDKgnEJrVbNW
jmwy5yblhKt/pSm2s0j0x7zHV7JT7QvH9Vb2z4/sCwHPBE24jTJ/zlpZO/8XuzhvPFICeu47MD5D
l65Mn31C2jL5zDgLCLgmle4xU1MdZABnIbtCYgc+xCInQkoTvrQAcJ9yaWRsaVqFDaZwvvTG09Tq
cwk6shHf5B+NluklRYWxmN6H3xm64x+iomp+Uw6q7OlxDOgeUoJmlDtqKqTXOVab3kM3C2KpktC2
Nc06uU0PmybdFmIGj1pPCkw+YCfpGbRlEJIb19huTiEtNRyNCA4xp6XZ7A71GlwTbQ/4SLzn2pBl
zmlw6I9GzeDwV0FOz7/hD4jpkNysl46Du4XGyHnub0DDcyQQkl1bhYmV6Z47Ys9JY/6ghfTkWWv1
U3I7izOs8c/A0jxLPPQJVxRy80PcKzBdfUkAOq9OHeelTUu1mDrEyCU8FPZzAlK4GmcF4vOfiG/+
cUFi4j0D1pF6ECzuuq6208dZDPkA+dkqOfIXBNXnIdUVeCXQ9eswqQMDPDDUrYntA4qauY098NFX
kSYz4F2rB1c46D/YS2a+FJwVH4xhsMaRrCUbdM7/mV8e8k2+4Ml8rOJUOtJfiMWjI7lqSC3Gojm3
W94pqgFIQ0cB2h6K/eVtlah5mCLxyuW/Gzw8thJahGxCraS5cZumVVo7joXSYm9hBU3mH2KFS2zD
r3/AOIfwvtVNIQN17EFY/e4xfNlI4zcBpVleRJRhTuC/V22doCiwhb9cu8TCeOo6vEwXQkHKjZtQ
JKzvI5zA2u7n6pijUNjfzPvLtKRlFcbBIqpbCumM8NXgxW1Zzosj8MDFhFcfPYnsYjePwXbaXgk4
1QCyiL4LzCvga7T22AjCiyUyojW5JJfWqMW+X//AK/la9PhbnzDV4rWA80fSKwODrdpPzgWmeFVC
7M0h0qUC2GlNvWbw/BEMEUFDXlQcDXFTV9lTLDLTUN/RfkE4H9cMAV/r+wvfI7WiwjnEGrvxvlGs
gGpH688+0K9i0xBlB+bUeR8slNWLVNoPAAhvTWXTFDv51dtWZ5/jGie1AaBZvM86/IErzMhLIEoI
hsZvrMi3AgMXWt7DKKoPaS55R5rGFESGDO3NMzhT1edtyj3An8ej9LQnjRkHooTRhXjYfWgF8ZUI
SiN//C8/p9PZfMgoJzy63SZ9KQ99q4teFQYF7KFJxhI3E9YMSzBMB5U5ObY+Tdcf/d7WqMiX2m72
qMJ8ekjPn9ebwAbIT7EjjmqRo9RQ2VuyTCXzUVjABQGDUErv2bEY8KCQ3vBzcgKiO+Xqnyw2QHUI
P6qwCBxtzUpw0r1ETF8O8jEFRJW73DIQaWqm3o6Y64u4VDHkL9KQfxoaacHX2vuqlL1Q0FF5Ds8s
O+kcph1I5dPgr2EROnyWu3b1oUNg5l8WGMrzIa9cYQqej25m+JLn5IYOaiLpHenj3ta/4rqSWBeW
MqqSdprs5OgRFsI1dP9CEPT6mjOWXTENJMuIbFGJxwCKHeXELiTe/9xWnXb5UqunksdWBQpI+zXD
QEWWJDHtcXujA+WY/eLji0g0270f3oi6IbzcSyoC/7r8wJOnGO9nips9+a2vXZgKaeo+YIiif92F
AnWJVhTlsKb4cRX1hEapNjpZv8gi0fSDhS2UQTfDf+PTSLm2rDa0qQgFjogycPRVYAVtuGH4RP7k
tD55tzAw/WLuAcszgG34HAhFNok1uTCA8Ggl0rAp12lrGP3AXhEgsbyvilTm8xBqTlb5pGfNiYyh
aABTMjOQdo81RljO2eDW1+FxTWqidrwaMrbVwPxiBjCmxKs7awc8kmi9IqtQmBBMFasSMwEjHrNU
0s1MjC/cx0kxCRmWe4h0zcZ9YeeHDgEAU5JGCZp3uZ9d9Ixj02dXMLxN11To/vZf6lHHGa+UwTuw
LVm1014AIcmYya/shesOMsHEhDRIff/6NJS9EjmeV298MWeUXlY3xq21cNmmi3aV93qa9kATfuis
7RCB45/F+QAVcqC+d0kdaN7sc3Fo7CUB7Sap9E7cvkxQxIKYv32r1M5hXpoOKSiqHEu0kgdYK6LJ
I0kwPZqwfiCNKEtC9GPhQv6b91sf9QkECL597IWTHt82z7GuhnF1uIicbI+4SzOM0kXkGxGnd+8/
N2HpNvme/zMAUX84KwIfaB/ItkQdHBWBdWIFdentSGVuRZKp9FaoAt9zmfj7IKoagQQ568aPSo9L
GBtaufdjfaIK4HrrPbARTBkVrB5Zm8eDLwN+5HmPVaR1GT6oPpLexdNlvPgF7QQteQpI+orAXG5z
a6Reu8NGrXJEtgnC6YeLUrF3zyw/ZTYiaPQIB5myb6VR3tFSxQeDFjoRrYO/KvaWpjHH7raW4rc2
0Sf+QfYnh3fGB1JLG0PmKNJNq72B3+Je6ZL2y/h9f26IXF0pYrWcg1EUgRvHiZ11kp9GoRgrBAqp
83ehlj4TWUydcEcXW8QJrZOJBinyfqYrXaOhAevpIbAlQj2svPBheJTId1hv2OW55O0UeSvcgc9K
Z6xtP3RG4hIBBxq00nyDcq+B3MIMqC5aSzVF40LnXBnJvAhHTMUeRltwPNGwgXwYgnHUz82Bzkkc
+PmblI8la02g5DZXKnglZ9danbShrFuowvQk+rK+HO7kMzPXrDbtP8TCVSQsAvqeF1wCzrH9viGx
9K/IwBCrtyLqZl1h+w1WFQVxc8MyMjaYBkh0Cx77DaeZ3FuzxvD5M3syx2xnFlzh88/W+MLqi32u
sUvC3P9zKRXpRUTmvrFUgXbo9rgmpW34w5Las219haCpqephApv8f2730HZBnsOSQ7x2X8ZR9QDe
9zUPfUWS3/OEHlWu82YPT544TsbaKr6e2xKsdmeqtRluX8h15HJzeR9v3BMtimEzbb2Mnm15h/AW
AbUIZ/C6mc6UcfMlRVQQewNK2vuBy3XSUUC+oC2jA4gdIwfLB8L5BIpVeRuq32i2UGzCixMwEnsj
nL/sPC9FK4A0BUbBc84aKCRR2jlA8uOsF/1EGdxDzwg3csEgrVXrogzScXvcW5mIpU5pGhA8UcN3
W/LwnWbT/LnOig22tq4LfG1ZylByFtIBwCml8yMglzZ+mvFNflkZswaffGxnRNFpk+E9/9rckx5z
pT8lOi8GA5MJX5jU0KOh5g9rFpGBlS7J9b29t0yPz8JczHj2exUF4kfCprBhquS3XrjoHXU+zT2z
BNdr6zAhSfrMw0WjLncuPzj3mWjJtkLj1WEQ0b/54akXOUwWZwoTntzTRwMkUk9ubbpQndyLFJLC
dP74SyuUHoWslJt3q3TvkrZF8CNNCrd+I0Zs2VKVkxXHgI8gTdPpsjKm9UOqPa3ItXvydkNy8hiA
WxCn7kQ5drSgNH22HMBuj76ex8Jfxh8YWQOc+0JstWIPv2nmmFE33vLp9vofgUmQvc/txTImRqxJ
cQQUBMb9FkprdKHvPeMgJAV7I1MtN38DtJuh+3dNAzeNd84YqojIjnADQnzT/nhlGPDT9eiExFRa
nnkB7TZ62f0CMEczL59XbqYBMK7ggD6MPgN3dvLcsiqiGZ37K3yZFN7XyiLXgIqxMDMx6LWCvPH+
EWk/XgYwDiSvTU7oCZAl9xCIon+6jxdXGs4CSKv/RW6gO7W9KbGGnI6scjPm+sLamdD0oE/53F5K
sCwdJCt/6LAyau6IHQAPdYVz3+EtYzS/qwsFRJuBzUUyrMcNMhGO2ySkavlHv4NdosAg/EcOlYaR
xSq+jWc7M/Gri+t5uk5xqXv7v0cpKYP0WX1L+S1YPLmAFiflBRr4UZG3DHtvjdLe4w80DLHV1bwX
F2zDdctCrg9q5jdKbJkQI5X73Nl1UM0Bz9ecdXQs8UTb3Wge0qUwz5lQjfrRCXdWQLgXzo85u+Br
/5k1yb4R7T7wFyibSAMwjB/X+dK4zqHt1601YdE3sPW1fcec+ntChePtDaLcVgRBnSNkdP6Fx4Fr
4CwnK/1s/rGzQxZrfNc3PqSdHClhpH8IYvrvm/KHaUtVsIGrlAD3+0K41Aq7aC+bFxLBqcW0bkgD
9lcUuQ06Xk+cQ6b9OyVrz/+WwseUOkbVK6rokHSTHT96XhVCTP2qsyQS2YohOrwZYkzECBDqAJK3
Jk648Qg5Nh0L6pj0WYZi3EBILtoa+fPdPqaFv1QoREApN4Hq16EdHGK2kr9u0FPRdHNSqdTi5+6r
IJ5gN2P4Odh9H+utmOghgiyERkBLynf5cLdSz55IZqiB8eZ1Bs/8cQM2rUjkEPypAUnUT4YxqK1P
h++HzAUB991FldyP+dCIuyOAMA2uOhrmi9DcTWyBJ4LUeWbsPQU7ASLm5CyFEOv7U/PWFgmUnbRV
WRoq4+9Pe9jnKn4iYPElbr8CF4dzMFni3raS5EGk4hz+jPu07rpn4eidN0fGwC9zSof8ViNU64P3
iYFquYPeVSAUwGJsBqeHFiZSvWbDGMq9FcslGR9RnnU2is40G5iboYx1nEZJTj3N9CU1Tk1Lq5Ii
8MMhPSSbGclqaiRW+sWs5FNI+Rz0XmqXlxuyuPK4sZS9Jr9EIsx9RmS1svvvF/s61GR6K5SnlK68
E/RkcHqfOf/g0MOFdU1pU0W0bhk4tmKimoJFWBoBYdNz1JIfrS5OJNJ6A+Igb4w3UeRSae2rEdBz
81y08umwMJcgyv0w4KEZteDZ8uZfehTQz8wiKkTojUeUpG+0GGbJw4CNSHIwwukPiwYPB3uj3eDw
IV4q+3dujWWAC7Mwug19XaBh1Oacq4uMK/L1KNmxoxeERKqCaBQDsIv7C8Wn8MVMYBaJNNBY8XOg
pB12DrWBuhWflRqUhkyMHQUNXT2s2pafcMc8pKj3+Am5+lSqaFNE319wsBoZc/vvkJSio3j4rzcb
FpgAKgi0SWGWSRSFYK0gcYM8U7MLUQI7gup3xxVAnzrY292g3g2l/W4fqOBGsAHmdz8F35WboMuX
PluLQX4WwRE3F9LKE13yxGkZAhGLwO5wiMi79d/gsbrnk/+hDGHKxzK3a/368QsKUZOMg9O9htIo
Yrg9LupCtG6C/zGkT26KiL1L64MnToaSCbfOOFhZ3hogJpFoJ6ZX2tfeLg1FM9Lwx5ppW1Sy34aU
B1fQGe7SWAPxhrGwfqzZkq4f2Ny89sVrOwvI9QTcuDezFqXCmBKkROtverrSVqy0MbpGM1JLbB1T
hSwXDvkwnlXMQqluajbM3seMg41ITF4MrjmDTE3SvwFESCILUadLS6ld9Fmh2H6BXxMKuwOqGfqM
kg2U6jtpx35b6viVwohIRn5Ud4jENqxPfI/paRXswljwHelSaT1gGk0HrFMCYITjCytl+wKkfupj
krWo98SmY72PbE5QgsgtspDDdgNQDL/0G2N7taNqn/8JcW1pr3aODwpFnq4oRiFhxUWq7JYI9WDl
4ri2WdjgjdWqGokwmPp99mZVAGyvnrN/ARTtZ3G+tMHsp8NAEj7L791woaS7BU1Wwlx84xe7Ro9C
MnjtYqcS9XrnVu+YS84mbqs2Gd7gkbOItVlwvg6qdWo/x8bZMDNsARJNpnSnGIUA/t+3NZhRCsEo
udQ4tTG6xXmP9cjSCsnSYvAIwho3pF+cN9gRXYu3dn/vGwhlGsAhjDOhaZNR+g10c2JI4uG75JZC
7yXuq44MFXX/AmhRPwe015VDo4zFeT9w2urd9mdKFNHGGU2zqv4kK3dF1huAsiwbB8DX5Be0pBVk
m6Oh2vY2jvs4IOl6he90ypaEDNADP4ccQobJ8zv0IM6rl7HwbTRTnB8M4KWMpd9w5NbZixGfAaAU
2QPZGtgPFd6Qw8k63CrRgxkHFStHFD8v2aDpQwq3tc/fC4R8oCBR9KxoLRED6xSPLMyDMYNVP7eD
IyP301PSK49tZLPU0atdNKDfYXyQN6Qw4ciz6Fyz692zrk5WZKefusr0f8fTFAVNu+qFSzu/q68f
JywiBNikM2SFisnrh5wF9G8x9tIi5psb5drKgXu/fyjXlm9iQrqsjaUsTRuI4kV2oh5AAWT25pb8
cvQ7lZkd0M+KUtKfZ6mQFe7ZJI8MLk7wl3OJsCPNdm8jkEvgj+mjX8wCam0s5jK157kOyOJ9BFmw
Dlu9Kq5dz3nrmjS9B9DJmgWByX2inLrb51WvXtm5qbkwtDYQV5A4oG1F4HU1VKfKhoXvaEzh1+3t
X9mM2MCANeqBejLqpoCvARFEtHP8yMXM79G/sZIXsdf/Iz05aWnDYMJw+Yj9IlsbJQ0rQt62YX6P
sU7WP4Wdo6QogzW6DyvN8Dpzfen0PSaue6nRphZIXFOFevcURohUsTSKhRoRCuSN1Bik8U4PSaqK
fVxcN0y5qTElCor2KVCL0+QekCSRugYk2AOGrYozRb6CX2lkL/o9C4Gwgb0Zy0w+Wc/rLCvR5Yf3
zRlH9Vd7uoifqWxw8ZlqnXIRTd1OOdrlI9wDeG9UY/fiaSoej+BkTk+a7cMvQDakSZ8ZHqpepw6D
BTKO22KJFeh6n5vgf26RpXXkuqvUqs7iMZYvy74MgjXMfOqSE96Ysnq+7lNRZaFukuii+LFUseoT
MRTmz9ef7IdawC/aY+JbLCMBu+hQdUrFJymqnjDnx7JTVhYvgJHntZnr8AckXRjo0HqUdWdAaV5G
w0D/Jj7B0cWhzQyxW2y/PiBQteTljquQjFvaF2tcXWQ3Aq6PFRUv5D3maAvyi08hLol8GRShbKEH
e5PRX60z3tzy0tbn8j7J0huUL7JIY6udTqdgHECZNDsj/sH1HcK73iJYwJq3qgZJYU19GTMul188
h3V/s3CyJLpZx3U3Joqx8iKyW20D600r56CGVB/ti61owpxMTqICkL8Ceq8Wa4AkkMpzj7TKff5b
26pJ1Khc7+Kgi8MWFrrZh4Sh7zNqG7qlPRk9qBZUa6V9GV4CPbfeIywIga/tkcITmOVmaPWC02MO
pupgsidgkuZwtB7bsmKBd6Mb1uU9tL2Knjjk5A0SjUDMuvQIGvhetdlm7tnhPGZZPqEAT1u5TLG2
1idUU2AA2dVmGMJNBDWTfK6jBlT4dRbgYYr4qAhV+8vcpv48dYA5kjWQMI/ELiJ0rl+v/Kq/aOdM
EDFhAOHgKg6uynK8LD0eZ1rI3KtQfiBqmXW0qg5E1XHTyr1potm60makQq6eeBpSRtXq0uBeAgEm
RXtsB9ZMkBPcRyUWF9dzLthFxjVlxUIFk0kC9Sg7Q0Jvz9MtAk6O85nZ+4z/cdaO5Jgwc+zgqzGS
z/bM4G3iMYmBsQLtvjjZ+hO/j1MnlcDG+OMxe8MKMOzh4TzKc//NfWFt2/vQjCEw+tgb0HrAlYQL
ZuDUXVi/A+nR5H83J7XVS5e2FhhVgbSBl5kiocVGD1fO0GNAbA7deQnuGpGq7TZdkEv/nOV/J+C1
9/NEC178B4UENXxUsRQLpAIwnfjayenOdYc3nFnsx55/7mJqfnVUB9F+Varqjj628sXhOfJCwAdt
2W9RJAD/xO8vfbWWVizuAyAj69xIIkqSmRoIL0NZ7aVYLPZAPg15vjHdCd2eOQyG/jioQox6AgAc
6Bk9KeyBLDeHwxpylvO6msC/GZhqxk0omSD1qv7Zsii61tLbE8zRGML0v0KZvsS4nYc5U/2h+P0e
5lakUHyqx4LssZjJilG9cl2t1mTpeAGK3x5+ZA3z3ieJ/ATiuNA/FjWqEloN1LhF1KFLSfmCv342
JG5Ss/Unb9ehY+K0dyTnRQIzDF7twvRpTgcDMhYmG8CO6cOp2w4jNjr76oJOvORUqe/MbgbDbf5E
/oMN2Vmr2xB6yLj9WsV7xXnyDbRfZNPUsWqfLsrxSGpwLte5LtdSpHnCLg+ssEU1hkFWcm4wUHMZ
R3E18wUKJJUmEQ3bJOy7u+9nOoeYFBL2lMeoMBnYh+mo96pUklASne3Ms0fYzzSPF1MS8twQFGuS
ndOgS2GsXVFfCCjueUg/mEmQHLq4sNhfBtOl30IvfbUFxyH1BolKKvPGp++Pg15+4DYCcG/xZNqX
LM9C0xLQWAzQxzpcMGy8s1QWr+CkIB00cwiSkKdDFPoN6rjSkI5UFe069fmyCZJv9kienqnPb2mo
hYisDRk26OXwy+6RuLtBkRPJ76UnweGSU8sQR1pVInX68fCpygur1A6uNSZJtjPHh/beeu1MSniw
2eY4MtClstPsiwo3c8Q7UHKkMlshyhhVnpVM8aGKTkCfFfRyQXSvfVoQF+aDlvEVwno1PwMMXy3Y
Gxsuxydqy+yAu4BiBZILhLc0uNr+CGmkYQEVcWsVRSqlnOb8HinhV0/zsbJ/1eC7Br0HE0MrkY+5
p0lTKM1vOcZY1fE4ZyoiJ7jkwWCc0EjaHznxg/XK+02wwwXQW1xqKIRvdQqUQ/R8WMVmZS8ErXTo
M3num/7oGGKeBaRq1ZBDuJDMu4zNmron7KdnNkarLLeAyKjXFCGbARIgqAlm0ZVG1SHgK23PnM2O
r0UWiu3bKwwQY0+2ULcO1ob2wVlGnJRiTxZ89a0ILfWqqySjaM9uyx0b8awD9nXBEnrF1y3clOoN
SRZBrDv9IGje2mh/De7ERDwclgTwLx/j/hT4vQShKB8uXqaROtZggG2YAwdbmKbaQel+6Ix+7UiC
c2fHhDqUC+7/cMIBvXKkt2MNbZNyAg3Ax+diYCrGl0Vm75MY1+8w3khtGWKeNr+xJ1uLOwZl3FHh
VL+c4lxGI+bGdtc4smpELcg5t1Szt03NB51OS1K7qUNUUjz/LOZj8DR9uXWtnQ+sR3KIlJOoPih7
Fzoy7yBA+4AbNkjqFV9/lb2e7NOjEKrmREoKrA0RxCa5vcVrD9AcPlSgJWKQ3mHhSYWnUTokjqdA
cOB0cdLJMqX+p8PE+hY+Eh7dPQinaGFcFJNv/OMl68TB8GbHWxZEZ34MOgbPyXbdAjkf0Df3Cfdb
E7EjH5k0PLtnHO72wMvad9mxzzTVnUBStp7mNpVN6pZ7tNzG5E0eaQSjlTXm06kzk9m2+1JZKvu0
nHwNMK0K7uSy/QWpCrhJI6avvQrJRuJ9K5ECBdzofl3WE70lqflYLyRBDmOQQ8FSLPzUe7TGKggx
ElHARz+bFCcjvu2fOFNrTw6Hlbf72/dzb7OxiTcn9EuGKuYMpopJwDcjitAWWn9QfQ+k79cgSA5i
74+fAPQvONl6PvTOxGHPc6TFmwpLrIKpeG86R2hj+gRebK7M0Ks4IG2JE3hoyUZoZ7OdswHg/FYV
wX9+3febeTbxFQCCzkMIivmqAjnHhk+M88cWZLM+VezGZy4qsxbt4aXyDkYcjtM+HCBbck6sqUw2
pJFxa5UAbibcvr/oMuRbpkqeP+5/5N6U2EvHWXDyyzPsnauh/wYq7TR9IZI01rXhA5xZbgViQvEg
UCDyAZ9EXc6V7fZJGW7LGnVyUms7KAVGGFbYbw1LXWB0E4bBZS237tC8y5xuxD6reS6y31Cwk2fg
q5VugvyZ5rNxsTZcxSjmix5A5ULAuTc1zTXNatWrIdj71M5CBcyWxbn3cvmF55VF+rVF3/VVwzMz
VmgrE6L3szUk25rRGM0Mpt/CKsiQCUG7vDE5sKV031K+yVyAZ4kCAdfisMrj6coi+SN9gpOtm4Dj
D6yRgDeYIYu6IpQquZLyD4p2szuqBbFT1wfjPa4vUbv6+dAdKfhvQ92zMZXjvk/74xLCWAGLbsij
ag1E+YEU8j+LMyx4J8eVTwUzSYJGJR03bYThu+z9kHRjYN7HMB56ELCgiQ5a00dnMNetDYDPBKJ3
ri5jNMo3a7dYYvq1w7nJwQSZC1cm00KPeWAGHGmi+DeTSSPwW+oWIxxA8iGDJ53wFGNIwdaYUVQs
bx42Rbpn//4o7+pGFBQK7wk4KDTgVs3oNoM6ij6BtWwFqVrgNVvDcFXI1a56wxlZnozXWhpteFX8
tHZVLcZEY/o+IwcZ/n8/xgoHuKwp6PUXNE8kjZdcChzhpBFshlr1gLFfYC2+gN+1fCW/v8gJYaG/
qPzq0H5aIta3bfhglME8sBSz0lKn6RoulozI5LFwZdrQo421zDIdR6xU568LHzitf6/K3bjN0UIu
gOJtwmAPI/y670shfdCTkpK+IDKu8as8yvvdQaqcFaXAfhvCtutVEeqJBE3PDQYd3A3Vq89wWiES
Q388nnTupJdJ7PbjSI+pH/USSy2DScxTAY5xqKLos/buxIlvzeCJXfD/cH/415RJ2fc22nlYlb8S
zLrbiNSJ4iJkEk1Yil18/kWz0vI2WHqHwSqmYVLrDz98DVcAGmdGWXjrC3o+ZvapqJ0FdmrckYAs
qMuwvB+ntL7F/Sm+WE0dk0e2s0LFe5J9x9AeF0qwTIvz95tkXkL50PBLA0O5R3CWEHRR0xt3jfVs
f698EMJrjxlg61sED4/lqvgq0hVIHSKbjS42DyoVYe09zJRcleCDJtR08tXt3ZPrNEukvR3D5kAU
wL6A15L9NzklWvGFhYpGhdvaFBdj5JED9KsE91hlpleYuHPahKLi0v3LSsbFRIseqtID4/rjeMzt
p+qvFyEpQD6bxcX+oAFVpn4LHW9j9X5wrGP1EU2gw4fzVvtelJL/fba6f3hVG2s+ZRX/XSAz17f/
PnDWEc5QtsT+HDnjH0sKtxOR0+shS3cLj0Bl5DeTQ9eByNyKKGPalzGCH8pAkmmPW7Bmy2QF1Sc8
8MN7PQYa720bpEaCDejFEAkjZitRuvuLliIJr8hGI6NejnJtxjEll7pOgkEH6jOb2I49WDWOQ8LP
1hdHqPdQb5xGNRSPoW5JX1FgtS1Br0Nk8dqqvws/GZRP8CzteKypRc2wpSpgsXp4wPiEHB8mmQb3
5YcozKw2063s+cqB+TrK4SgDPMFzfU2fEmzehOI73Ot4GJ0HeRz77Bd3ptHI7Xztvu6EpVuhuNAo
461cF8kw1frbVGKqki6nTQfp+cPjj2+CMLOg7C/bh9LQAEENMQB265vCVK/iqEjznN0/7+XLiURk
Ck+rsYe7fAchJQ4kJ21ksBbTvuY6MgSH5Cmoq2kxLtyYtoTU3Uxgxux8N08uHacVZXZRw07afniW
HXGG5pfGeOKVv0Wd0HqLBo9IckKcJkfZAYuxK5iD8bW5QyoqEvdmD4nHgNOfTweeiN0LBAh6jcn9
g6EdH7tBb/bMAT42kWMBTf7nIY3/JJMWORXTgt2nHlVg18F4EIENaS/dy54ywziu3c53rRK5iVXC
pIQtJzC09c89brErdJqTukvLgOH7b4MSH4kUzq6tuJjdQN3M/Xf0judAKCaSf1Gk4UvecUfPb9hy
BysTIySTULgi/s6418WG0UImzAceujx9AH1SSjmJu8pbBtdfVTwxT1dNKg0hl8Aal4MUj87McI5g
xBGUDN4S1nDq4goyHAIur2wb3EdGmw64+Ckmy9Q75cdM4uWWz4fbVT1RZ2GCl7GB8HTqBZ7nBXPm
Oq9jnu+cWgTPQ3PrX9ywxwxc5Ziy3IoTGsJYxCBMgXOOcQ5kkpTo5c9BS0s1r/oAB3ZEx0QfulWh
Xl7nHswuZZTVhfqAAEaALdTTxlJzAmihwBvciAH+Tyawi+zI9FnwyA2uXrEe7tl/szjagRsRejaH
AIBP/8rDt9NQ4VGQ8iWfWuUOIcWwqjfnwXpoOtWcKY+pIf3u+PsqPJq/Vxt9CyFBx1umfbXGnfH5
7UYxzKvkq9DKmkXTP561n5m/yjj4re2HIW1bt1Ah6F7HGejSMrdm3jcTZ65luMgS9lUJ76fSIxuA
dHsNeqLEkJKSQ+IE0cjxpqwkdwkyf2j4+BDdpFXF/YDPtPU7K+vrP2E4uSzOBL5yeIkLvnoOUx0S
JGshZWzncITxzuDMFHsL0APpnkOcZZYn+K79W038Q1D4T80rB9N/NjF+wgpgscdw/8n5jOQzuKCm
0tvdwC9FjWBNzk60VsMIkeKasHMduwPV2Lg+CVjCGfVYEAJFDVSbhyyxhWyDYH6VMsue6I/38lYa
qU8pzFm2oHml4FDUV3pKZz9MlITUzeP+La7dB/UxbJMKIqdtVwVRlIsGiVizjrbn4qLsLYJ8G5nz
vGcc680HBD8U4uFjnSZaIOMNswvzL/UFKUGvuvpRYBw6JVcXxw9CROsA6eloBORxucyXJn1UyLn0
9O4YOVYrj3t4aV7oKvhqOXsAhlUr0C2ylurleOb2sZGl3E3KSguVRZ0bO5ESbK4/nrMSU8yjCZ6G
Qf+S+XuUTEzdmY5CioCL3A0MNBFWL3GLQrQo31SZEUn2JJ9tqlIqXB+EGpFqkz3A5XZsDcSTs+Uy
uD/4LkFKglZVYHTszLzHofm8LGxjdLkQBj9oKhGFkY9HP83NlqCSsPymrWaG6ENyJLmRJ8JVZHTq
fcrNwAu01FFXcD3t3C0kXwadQ9ZB/qyulYiObN7sNdPmnP2vKT830wW1APQTUDoKEp6DVq1+D0eG
2tqSSKbgMdA3Lk6n32fDojPvyM235yJsCMetypkbwrsnjk+IiVLpJK4bTWZqmT0GV9QWLbIkNflw
IZI42XIDE0iyAg1LXWyJ3caab139rH+2YW2wKyYGQZDLQ52V8LTDkh4tPca616ka7ZhIAKuJanWi
tMbjdo1FcnuMyu9gkeCcJrsHhr9NZ/H/2l28JCS61GpSjNJ1Oa4dRjtd1sDNDxcTdwk9M5J1skWS
PsuDQDfLIb6S316BA/Ko0Eucclq3tSwUczcKuwrGb2Bx0sWc9JaYaknjFXmhOxCWVSEE0We1gfFE
hoSnokpkMOB6Hl188Fmh1YfgTrODc4lNEN9MI6fO1rFMLpQ7T9ymAZsVOWpgaTz3Viuu3exIGFds
AkzYlUmlu/PW+76sfzlVuE009NnlUj/f7Uw7Pcqi1/6cYGyZ0oXjRxSCbBUf2byjOADeEIu5ncUq
Nx4NBt4h0DoWxw9wJXZybgmc/xBRruiTR3OPd1QpVjY7E2+iWfRiczTcGa48kcwNRIzCOGpzVmNK
FvSLMdrI/HTeN6c+UWg85m8+Npq1oXh4D061g9oyDy/USbUtxDoiHlnYSlkvHWQfgG5N4UytaYIG
LQhpdRTCoZwNJBdzg6YlibDNVF2OXf/BD1dgu0FOv90xkfTtjZ+XX9Q+zJdzpip78AJu/68ArSfI
twRmCrAUcVVBStIABDx2OYX3S8tysj0TTulx6rg7asoFgyNVDSvWMIU9vrDoN9kv9nTwROTV1FJW
Ia2MG+LqFmPY/5+hCJ5MAgp/CdbdiTKRUSy4zl49eIbi8Uyl4RKUNQbXBTznu0d/ujxFf3keOqbw
Qbugi0sQzGm08RsJnmd6QwqZfwXViz98IZsONuAdUdJmGtt+wzux0Na9xk/4n1bSndd611P2/h0k
LT+SsZ1kQTe/Rv5nc4c8q0gjU8MhCsiXdlWuWoR2hXwMIKaGbDMqAUtCz79gGQvYjNEkMeM8hViX
ezqjAO6HsuDozdUZ88HifaPYzCVeJsLy8aogX15OsW5TH/l5NFJa690r7NufWSIwiy/r8W0zQIO6
ui48pWDQbSR1uBXzFn07OByhZFd0zEgryTZckmVQ1Rm4lvBHFvpMFpZqwap153xKqqwhJGF2bb5g
ovtF5x02n48yL5e/5FnKNX9Fj9zwtY1U5nUbzF3zRm1DAy/nuLhBGllm6T74k1Bpog65gA5xe7E2
WWvkWcQPBq+sOI7CCOwrNbe5WlvF68PHhDb7q8+9xJ1pCUn8KGabJI/Cz6QvWoaI6zYsNFp6FHr8
OIDs10EoFZAoUZ7pS1f5BbUwTEO29JmWK33dW/OccaclkBqYtqD1Bmx6qbT9jsT/HtxSb6ytk55r
RceZylAQTx4hNveXMBl6/u6qRrfkkJvfSs6cw7FmCPodP1DSz9IvIOVnUEda/D86mu6KddJ9D727
EGCoRH7sAAaSVET2tWCC/zJzZelD0242GHrhV3zyz0Txwk2H2XLuv8mAu1mDCUQkPuaCGmdLUt5k
t5giKcrmVl5Rds0Ib6aZD2AUXtisjnI67x6YO2JP2w9szrFy+TACH2UcPSHkzDqpArWMa8QzC4Gr
RC3Zsg5JmUmQ6poAxJZUuorQDI5T90m7BZIpq5bKbL8cjCLwD4KhjJdPd5vevwOA38wYNYR13vxU
h2WBckrukfQHiET/xyHatWNOamfCDMe0OHoiUpgOFp68UPo/KmspRGqm0BJ6r5Svkp+SOBb6txaK
A/DkmFMBdKOXUL5OP589JfAq/yV2OYOJz+sbwXqVFJ3TYNriwwJ1GandUlZ8gR90dZrwpFFxuox/
BaC1g5ucIp9uzjxqlDi+E/gDGxsDbueklmfNZgo4mWjv7rJn3TOhWAT56xIalYuqQW3Doq2TQCNr
iDP/J8U3fpKscjggYKMzZOOktF8bpmuZWc284On1al7dNsEStLGtAaefy3H5WyvQVLWN4Soe64G7
RffeVc3S7AeIZGIJ4U/8WSSUiL7BzL2OjNpiN3M3UfJ/MROXP50pTECHs8MBtrQ31J5Mc9MKGmkR
PBya12jrNjCaGDAg+ZVmVxAd83RQamqK8eGvn6OyvbMm04APuXLP9v5bi9mZp3xZfE2eyiZlaQi2
8hWqVoSqsknl5GsM7unLIFLtVKl1AlExteVJ8PUnpffaVyr9vwL1eDks0xqoWkzT1OErG8K6w1GI
/Z6UgdNUm9nezIIuwBu8DDyCOB7vv+8d46QP8jTqrZSa5GZdqM70qzy5EPAz/4u7me9jl3vgr9zd
icDqeh6jnIsXlLvbbhu7wp3V6/T0h9gLCwE+x3/ZHXHnnkuus271QpV99yq5yRefNSGb7S3bgEl2
IUiTp7Ej86bTKdzYhFlufHVlHqJu9V4nOstNaddk/JyXaUSeXJk/jWrUgt/1c7HnpUw7syUYbm/G
hyHYeTKYW0A7eflRqq4u4lb4XB7VB9z7AMTd/+iq//kkTCM3ApCVu1+dPvbazVn/cQ0yoVN99zdE
+GETvis915EC1vapv5O5PAs4VF6d5H2i5DjQAmw8Lj+up7DF4hV+y2EYIeiOr685AhbwkRkMPV9f
53Fht4xJpqj1rh1KWbI28M2eXBX3R5lHksYDEAZsUgMKuNFLUAgI76+zHLiRtQmqsWWSs3C0Jy2/
A7PbCWAV8k4WIWfm3qfP8+1BQnpmIUZ+c79VDKbe+WNllHq+XX8Vn2gSl0ZkqWu6CvMmyDRvKXly
Q9xshVXKSDYNMsW7vIfaAyHCdq1lvhOf9yEiVix0w9ioRrMDxuhErNU6XVWC9gjmEMfclsvl8iG/
Sh7y6yybs7grwQkCvekkN/k465gOndS28CWd6lo8NCA/HZpTLsR5a86bejmtt0RfEh/nJ6ywcmH9
HyPdnPWMisneUYW8vygpvFG7Zb+I7nxCGCAfwj6rrtrIhPaCJ4u2sEq+YpmWF36vmUe6NkoYnT1C
f5gfCjRmwz/CzSlREdqwUmZHYA32h8weeRAHpgABGk0wkrQCjgFkacskJeDSy9RebvBS0yVsKtQc
RR3fOF+VHNBydAnbTGbETYjoQhggTv3x/UQH4GKKhVR6ZGEmrw6MxLa7rOWUQWNkqYifWC7fengR
tvAjmy5SyTy2AIltAaXxy3N3rrGH4FcOnPRl2bRr6CXGSdZm1TboVs0v8gEE5VPM0qoR/Pjebzwt
l3AxXSjHFVUFVk8ONe7lDSdoj0UL1qFjjJQWS55FhPBvNEWS4GG/X9F0V3R7WhJuDvSWG2ZGS+NT
oHnFySXUTiOQ4ZOVTHrddogd7z9R0V2Z3jYF+FIzlrYY54B2XFt0/DezptxxVJQnqKkergSOD5uj
vHfcR2pjfPkGCkYKx5CvE0zpW1wGNB8YGKEXRohaxV/Cozx+UiH4o/kyjmcyas2sbbN6qGoEBuvo
KWxMrzhkwo+lJBiB/OKWImhX9FGccR4oSHRQAmRQnruScDDgyjik4GqOB6ZhlgFJ69KwTAN2/A2n
B5bQxR+r0Og9vEtBfos+nSPmLRwyqqcTD/Suz6X3oP+yrkB2htNnmX7qKvz8bfBPFKfekNZ2H20a
mpmT56S9KuFqtTotlb0+FP7LbTNWdBeDm5IRukBsFmVCo8/JSYIektAB/CNuUCL44n6kXEE8p/sx
/hBjQ9nXxFvxXJfIyOaSUQDA2Rp0r0RiFEKo/EPCRrFqCcTyymq5aGy5oEavc0gEVJrBiG7jy+uu
Tdv1qhEkXSmE3U2WKqfGZiRP+rVdJwIDuadTvVIQ+ZgZhvE4FqbOOQJR/8OaGkm5QJDGk8TUK1Hx
U2tDJDQ1gq1s+6P/pJyBvlIcVYzdkab0QPUnx6B776Ud3caAsiNyieqbHFzD0sYrqE56NBbFnW/C
4MtKZ+QEfGi5jmna8YYYfePdPkSDl/APsWVsUUllp4q+TOtiiTFDxcx+grQUyp/5D5ycD6BIwtu7
AeeqGTe9vjbFc9NSDNz7V673wFpDk8sq9U9r35GRWDvm60FyCHWVgm9dzkIS0TbLnGYY7yzLOD2Q
JqzU2t1KVts7zE2O1zu71D3mx2vCu27XTO94nG5WqePZxeHf1UR+jeQr3xGXYl6L1xtITMp3w/Ja
hUDilJ1YDRau4OMxIKK+NL0y38m2w5Vt8dIxwmcvvoqpvkJbyMPaFxS6BHdaf/+g3w18LO1jDQYi
ox1T1PWgL3GRWt3gadj/7cBLb+A+t2B3aeLB2vXBNUArflxNm6KnPJ8k/G7GpiZSE9Bx7NGCsenC
G84yN9su7OVcsLlg0txiFzRqQ0CdtPNsHtOWyfd8I7DsaLPQe+uZN12QqXDhBUPaiSWAdWSccY58
Zg3EmDXgGxDzo1mxuplIUffUVnyNgRjrqH37Hp52hocxezlokKEsgT/kk8+Jo9+lN8gtB87rxYRM
VcjKiBlil9M9HSs22ARpI+fGteUT67RJtQDCJA7wJvJFpYvADRf19+E/POOl/A0QOL4MusHDyCTF
gDz2CCn1YKSOdbG5nVkuYAmYDhFzw9RMzKRRa71TILTWIGdG0E/4GdcvsKe2X5tMuKIdNBt13QH2
hzxhxjZq3/SSXcvLfEHvjpBp6Q9jtZdlmPc/Ohxd1NK9oYZeSEvVegywCQoofpjBcxDxWLIDcibw
E/tqEdmhnqRQExg2ge6aV2U7uSv6lbAGBOwSMWu6cqdgl+XWONIcBCmI+gqZcpaOsLxKLwbBwiWA
N0BbDLesYXexaYhiM1GMwDgmFLEwqjcs/fwdL10T6iJ+/v9Lm5C/6LFMOTMaBi4PUEmvnqKECl0g
5+OoLos+aDCJ4aoC8SxwoaQzrmhFKb+9geutcapKrpV34my2dSgHx/O2Ut2WBb9R4Dt34aTkjwRD
EC/OTVMnW4Bo09PcU8kzNJgu0GjRslEEH4Nuci+7mVrsNriSczKQRUtyrxv7wVAbHBCYTrNdfsRg
DiR57d5cSHE5JKzu913kJ4IDfBy8PdJLUrHpi/NjqjGTC238VZVsxse0Ea3oh61NF0IgQayBNp7Q
55yc5MR2sIy3/X6uibli4qSWz8aspxhyYnYmfwn8MEAtZ+foZZzvTdGtYrMUNHjMBvdpIrPze5lR
3vTdZu0385nbajyIVb1flt5e8Emr3UNhu4UW9YK19ACp7LNcuM1W14873fu9pfP5UT/je6YypGuI
7iyA1uw2TJO9gCwdMoP4NxFOd1IMY/VqNRHIdWrj+RawxFun/pCTHTP8oxvDStfD9V4Hegx0baeO
rYcP9XTuZaCW+M9kzFTliAHAewlzyKn9XbvafSy9GsncvLfF9qlQ2ceRoo8W9P3nnY490Bnm+smW
OO8GCTqAsL8xVeYrSotWhWWLNWaO0m69QrL9TDdOzF9Sj7txDhpYTe4tb+o2r7vnTJYj/T+To/Tb
LcFESOANQ9JwRqs9UU9ypwCzKlu+Vy6szZrX0uy01YlPSHz45rGYyk/BVWOYoSfIvGMtpiTq3mII
ykoY8EB1KE8CE1BED4Iz4IUbprYYEvelaOeVMA5KTOhFXA27DxI8QzYndc+1ZqYhEiFJvHu/mJmr
icEQ76W/1yDDQWkb9876p0/40RzaK/Ujfgbe8zwAb4H7MmwOltzp0Acepbbft0elMrAye+wyr7r/
Z3sGQ2jjo6wCeCTKQtCc60AxoxLHAiunxF2PYUqRTk8A0McqLhjbBiTcQZItFnJ6G76DoB1V/YhY
h2tdwzX18+y6i5rokSp1qJ95BScCz5AjgZQmtKDGJFnt3xj2J0xl/zQInDj/BDQ9e0hwUWrmhR87
Ih/NW3KNo7i44+4TGfclcVd49SDr7mumcpvRzVedNvi27tOuNVxA2lDYqC1xFiIL/x4yC3EXkhHe
iYdjNu4W19LgZsRIdM7jxHRPtPYNCf1B+zfLVk3PpdDoUBz/DdJjJsUq4hgNSIb1cGgyKFNfjOqw
8IMnedBrHO2USq+vnzSvkBen6rcpvnWRra57inwhNJE6T0LJy0IdX/E1zBXw+phu/9Bzxpo17hn7
eeMATXGPFFHHtLI35HCYHALBZSDHaFwOsGNGNj/bmwZoyBXb3qQ23Hsl/vWZsRNrJIKG0Nm2G+1s
evjufTErtzbmDDOLh2umXIPjqmiJxp9w7qyQub0+6QoMEwwSnlaekx2tLR4h5d2HA9upSmmQJtMZ
UM1UEI/CYASN9I75zWUgWk06Gf6UBla/V+5UgvIDpk8/8QkOKYzseJOJoI7NiLfMPvnCTiihGaYg
z5iUv3VJqxEPlbdN3DshsfAPmzHRoCOI1WUABxnICb227JFyr8Vx0xS+cxadTiNNRNvhZ1QjNlKF
jV6QsrFXkE8UZ0DOxSZ9wVvSpTdPs13rPRmGjttljetMTSks87bTxXKgW8aFTk8LlGjU0MtCrzB7
R889lFNssj/gfvdtt2vQBntHVUSNnpSUu/4Hd81vejeMeb8DmDWw+xeMNBTqaPv2uQ175rG1sWIl
VLUVKvcqYDCa2Jf2BuJBoPkpQmUg1L/DT0fsGikJI6BbdhqcA9lXZ7eOcCzfYG7dgPoomIMOetc0
MPzNhQHcCkx3kvte0Xa1Ks4WINFoPGs+eRt3MNOB7WYd9MaQPqCJrByoEh0OfqPKUm6xzG+0XZxz
xyXtveAVOWzZVtbSVECZycLU7nEHQqi+hvImcu2E16ROM9RRJ+KJQ3J4Rauc9+L7Sd/WDPef92e/
LebqNK+HrkYsYTsOZtRp9tH5BPpooX+0DvJWT5iBoZTGqmDo8rNibqMi/l6iRmbNUiCz+2Bs/WhV
LZxw1RCcQxD1jZHfY594TWBbnjgyNHb4YRXlGlnPr4CZffw3X/z03eahTUBuQ6yE+8qZ8Zmxh/Cr
Y2zhXPCh0BQtnhMu54L6w/ZDTVYoXqKoEUzGeKKsQRtkbVaPSxXgMSNyw/3QgBBcEixue6LccX7+
QEazW+8Q37o2fV44Kg/0qsaX6EZQ2PjMcBj7MHFkpiTYcG5utZO+ER2vwjQUeo6RHj9O05SOYecJ
0YIcwtY8bBkxL764mTVDFFt+HDHcQmYbY3xXBK3hkHxYe7ABCjWKBr43cGF+14A4+4D1JCWYFa/a
O7/OGTkSgHzlOnM88TJ29WFd+J+M73oi0R4nG95hO6+05ABnxawH3mxjDxwcCMuMzJ9Cxgj6wFl6
fwME2Y2T8it6LMGHkBHaVNFM8NyRwvFidqqIFXXfAgd52N2THZJ7WRzwSqubmIKM14nwwQDNfgog
aNs+tNTWz99Ap5hI3kU8fJ+NGe/Pk/Pr3El9QA0/4zoIbgbGsnW32wIJkhksTRpbGzy5iSIfGfMg
r7MTzuI2LR6MEqHe4iEWtYSQEaZ6SNw6R/KpkJW/mxx6gHKh6ZDkeN6tH8do1Oh3IjKVi5kVM1JX
jjGN1S7nhocxQaFebdpqWvJZgDNWijpUGkLtG3DrdrM0noU82ipjlwLcNyKLnpSObJybtwg5pJhS
nQ5mOaOZkn7Ma+vy9LF0ehia9rjmSUQ02tGi8XkWYuZUR4wCd4ML271fAwGhxe4JESPvljJbLNLe
EPBEuRH5hqbQoO/NaDyYvEU6J3qWCoLX9FfhS0Ojd1bDulKKNfFwfp6HTC8jAU8fZ56hqYmwb80F
rDB6odUKapLwtDjpQDOkYUCrf29xI/x0wYerhd+cApW1uWwQ0TsMo4lCWjpe3q2pDiH8zpvO3VIi
0udOHGBAVDNlFtibydotxDt2WdGCyQt1P5wYZz7HxxsKVk2zMmB3Hh1pkT2vtXm6Y/Jf712a0bXh
l01ZmS6xYEqXOJMaYnIi2SGrM4XgbmHtAQe9w7Dq00i7lxUy/4iu1lBoHwop4q+PYCN1OZ2YvZM3
PnCEf0cBCwFdtCH4WOt4XZD94UmRLMi+z6KT0105Op1OI1EsSZxsZhymp893iex4mfyFfrSD31fQ
mFSJmdDJ1wNln9+nm03NuRCEEyDvJz0nwYhrPwjxxiQQwM04/W2uGf5oc21ZXvMK/EQky6nreZnZ
23gbSFTQronvtCR/UvaXKioQlFcbeCLx0CAzU4J5CwS0grOhCf1KfMqDOHDGY8IJP177hdcGct1p
v3eZ/dvFLBZnf/iYDBY+jHksrgRo0hRUtq8Q0DZgbi+/6H/EPh/Q9dvhHKr4gi7OEKVM61DRiYz9
Vk2NWHD5iyM9syKe0pxuuf6i0u4h89AM1cd/HWwajrmmY1ss1LaqeqDr14OrbHw0MlLk6xhrKQFn
v9/vkNg1kzAcz3sKYPfqAVKYk7h/rdMN/9s9pE4UUGG3NPCVGRfY7D+C1R6dJTAvczfWnntutK7U
x7IFh3xAOzEg8TlIQGiH2OsFMNKlxpH/y5b/3NxSr3HZbpwYDQ3MniARuF6vBnutoCEdqnyCfxiE
HqusibAua1m5+ge7cC9VLUXpsLbAY9C1zpMIC684/LvEvhPZtzX85feCAzfsWHAfXdPV0tV5f8nN
YwZkRHtquWEIWxf3y65HWtnpui/H69Ui2bxg8OOv64+gawhaSekptE2HU8ylORpt/LnCVVxx+OyT
iiRQfR9SzjCpN3ihk2lH62qSGTUMBAW/CIoZkwGatuS9G4/d15gaRmo+FMjCsBOP6fVE/3FGsUc/
8zRtCN7JypGs2mtPgpUVTTF9Hn6CBmpe7oxH39pE5LpCcB+YLWUXapL+xZdYw0T/hwM6vCWR+xdc
AE4zo2SBd5ctRAbVbkdraBOcusanyUxns+AzFQGLx+Rly/F2GHvdeb3vyg6odrX6DWGwe3158s5d
EstxKScnXPKs4bZ8AsXrAiwYpXH5J5OGmw068f7b9Wo0Sk/2d+ACkAMISswjNnFenRWPK4Tg+0QM
GrJm80dr5tww4WGsxAgG0hafiaFwVc9q+PYc05P/lW7Fy7JC6+PkLfmar0cIZzhmHybMm+txH4Zo
Odoj4IyfijSkdVual59dqfBenqX40PQeZxvR6FHHPaZGb58jvHcC9sBALA6XECX8PvTlLB+Mzqea
UXyVt0NEWftTKebOn+baFpPnLZVy2WyAbUOf4IenyvmIAdG/jiObpiLGclp7A/tRzoJkfCjfYD+f
Et04q4Npu8QGxY18lyMNY+Yf+ESksKiIJsSgQwzY20FCEjsWV3RPBlnEexiRDsUp7t0NuAUXL/6J
xt37HX01Jo1M/zmN996SDJhI+NVQUd9eY0/r8txUvgZIOYbCVDH7h0ymbCnB28hXoZKjIqVcXfS+
w09eHurBixUtOeo1wMmzTp0ZecEmyPztVNTt41fmRxTWstGnhEMRZ66GtJCzuKwqzzDS6heSy65v
DitpCT2W/QKz0X7+jzbJmDNF+g0bUVAI/9SrQxKvsmI3M/+yB51kgIQweDvGbtR6eNDF7XzOkavR
XHNb8AtZb2/eRHywxJfhLSge2LDguSjDA+sZEI3u+BgDUJknxSmibeFRXYHhzemXJog9Uv2hQnBt
s5GjAzvCXZBfDDSCOjvYBoGUTYQqVOOsIsXuB8NUdGSxD4RpNFmteJPfm9y/i8hUc5eVOXrnz/Ut
kbG6vZ85roaRXvQoIvswzVa5Hvhe3A5mKQJRHPQv05WwpkrPN4oKC1+GmFsbVhfHYA8Ht133LgnZ
0b16U2nCRKR5GUK+BCwJOGeaoW94v78tLdFcd+i7Xs1KTz48o5SnXHFHtBZKa+yAyg6YNAkJSpda
cxOKLbICm51mseB1PTrNNAPUurnfJhMS3pwkTdIxVX6BJiNOG5wy6kPorB/6d1cPvVQwqM5dDrkw
tU8fZ+p1tHen3t+qXJfj7mC84zkK0JQ+P+YQnoMNoOiv1T55h9DsRXVs0I+eqTgNMhgaxvnhmgHg
zttjQBr58H6J7qjtPQ5x+flsLfzaTUxjZXi2Jum1cL4UdEc4ZwJs9tGIcE7StFq+5qGTN4BQrEgw
+fCJLMLqFTKpMe9Gcs7Bkl1dbh9o+np/9CN+PslNGCCZL5ytBz25quHZ3hr45F7cqjDLpBKTcXg0
j2hWScrib0Ya7xUTfBrFKxqJsmFmnVIptOTxiMT5v0vYBYTHblECZh/VsSLMKGnrXbG9vH7MEs93
GfDjORUBQqEqmQ01iW3sIv9lu4cr+D3qjI7lQiUJYkZJr9wv6JKdStuProGE5Q+M0LhUzY9cLQ+3
GvvKdKwiRyXGGDrI6g38CBaOWKdxCHztkklxQdVBEoxJpzO7DrYCkkVOhGHuvEaAno9yxevVtDQ0
Q6Sngnd8Mm1K6Vb28n9GjGRqjhdt8Zb/qVQg9vhy0bkESoRw0wlZaROF1GsZBOebplTD1PFo4lqg
T89M61XwgOaOjDynZOFz/RFgceZbMAGFuEmYALvBJMcj74My24D7q9T86/wJ2+JvPsHZg8DmZQie
kqWCPCmk0rL3A2k5vSFy/yVsG/zAeDb/zZBhNdAINngHsV0S/eDu+H6Z4uPE2OR9xKad0Of5bsXM
Wil6JQyvQn0ZAxXrGmU73gnCmHaN7lcL9V/QtVzJfSe0wY/tPyrVByTNB5fW5dHQnb9161SLsLlR
oBPfVGWXdgyGvZXl4a58hicfE5FppSLVBzHIR9ZfyguZfZmv2bpdeHPvZ/R4WxNQocwAWFMJiiPA
Dm9s9xRkvj6EXw+fXFSGgGPflRVXbkXaUprt5KKP4AqGI/PUiGcQTD4rSxGQAjjP8ROWWqictK1R
fevCX+VpWsgoypBCJkpYwSPjxiSUWKSvDmR/VobLjAqtJ9qujsVLCMEvJ7ql1jQ/ylK2fpySlra4
Pvo1g3HdRDiSxFPhMgMzcsG6bbSrvpvFZ7bg/G31vuOkTx8jMy+zMbWvgjZ+VJOyEJW553pKY5U9
LAvqa5FLmU1OtN1Eektad/63RgK8iRXvRc/AQcYegu5utlRl0z8uaq1wRuRtAxSEtob8sMNia87e
N/D+BichgybX/60Z7288dH9QfjNX6T9DtYhu+08fc1kLOl4yCukRPM/81g/64pP+wfrX3nnIDVpR
9r7FF2I7VD03s/8+E1Sk0SCTFbhYK4O/sCcp7G3anrfSC6jvuewmYoB+92PTI9ojpP+Pl7vRf3Eb
XGT/QgO5bM5Oz8j6xjSse6lla2b1C1sDBQoOBGoX8rKUVmsSzhm82GfPCTCT7k+kf4f46x7KbK8D
1Pm/cRF8jcPJhfRBwRocLI1X2xqmFQElv05xnr8Q7A2jQS4SQUpX/5Rg9NylJ3w5/1EoRQTSE7Ij
WKvIqAYhEOVN+WLzye9X1obN9+kWMyz8kLKggiXTc1Az7SKflHbUshkS9V8go5QNAYrFojwQ6cRw
nWsUUQGhFx3n+2Cq+xuxJ3NtRf5R9SavqZKaEt3qgJdszcLxtv4MQx45pDDPz/hSYRgQtMwwEcnV
Di7SvutQbVKuqL2qnXJ9ATwCQPzL7oC2F69cMG8Omhp0vC6438S3A6Rn72MwBtZhXB+BfC/dD0OM
8EJaVp8mbz5cIvv47mBxgIFcXGb5+lgADWuuCUIUXhWQMxjVQWbJ0DImsBxXznBF85Xx7GAJyP0e
r35E1I8B0b1dh5Wy8bjERLym7JMbm1cSJV5VAi0607bckBTqlUuAmx5bCNS+KZEjBTMJPLKz0FqB
bf722Dol0XDZ+6UKa/Rr1b3U9dc/G7tcznH5seu+KH/lROKE4lRtv+IT8rCTiGe1RIEhcpwZRIWU
2RsXZ++C2Yl9894v1XrpXIzYEVmdJ5ROf3nnB4cNukgAedcJtr9lLDO1XKj+0R4LnV0T+cd+jsHR
KLGSX5GNvP3mnAZt9ZjrYJ0XW4jV5/21pxdKPjbg9dkkZF2dC+4lhtDVcCsMYZkShYBANttJhWqy
OBofDi580M6La/W8J+Zdd+B6dKHL20kQW51h+Hl+y9CsRnU1CpzpRXGkdxb+O64D2ItviBcZ2O7h
CIAci6XnKgtzxkE3ptQZEhaVZxRGUlUUwOP9+s58A2CtLb8II89C3EeotXzBO3xTLfqKADU3yd4J
zmuvJbShAXINBrS8+8tTCXOP9IYXmGvWRH1+B8SYVCnAm98n0NMOr5Amf5qgme6MbMtDCDa0HMI/
WTx7N5GCT3rd0D3s95canJ2Z5uwKox/xhFCyER1rN/I2p3gq9mDhs3Q/Z6PKZ4LN0cMygjZzg1vR
YLV17HZykUAZpA2Qcc1gxO5zheKldcamuRT61iuhF6ImyGQ/90ItT3PVeTDmbUWNd+gEBJ8ZXsBP
2I9WFu1f39zFsFkcF5SZGGg/+qg3SQecDLdv0GAWTdo4rpBpuetOvRMx/GnhoynjLD+P0kJxNNwh
aJ7d0hA0+3ZMhGvhone04ejSE6Cd6lXNliyviQyrY2MhC1KdjdGwuhWuoWlKcTvU24xbUJOkAlyH
Ms3LxLuXrK36aWzmoWuCec0xho8Z109qnXRLzkXi2dKJ65DH19VPbvAI9PO9ANmbN7OzGprQXHK6
lby3BXECiOCitnZD9QjWRnN7XIm8SpdOQy52odYBp7DazorGZJXC/iT/oBVXUJqTOgogLai4FjaE
lbbPNDPlozUhQzMDV+oxtelBUYGmCJJIQuZlAg2BRuscc3EZop6GpFTjzMWi/bZon0L9kLNp3rgf
yhTgikDxVqoxw+J3H3N7PvHD8TvP2sxyMcMF5fuVJmoJFj9sJgHo7w4tlDlkGAPoXYHqF6QqXOhk
U3slMJcHI3C9EVDnWcIIM0aHA8t142hGAg1/ZJ2j/4h9/xKIqrINYeIpplfzsQsDc7v2l+krex8u
7rgir75KVoHvmT410ERYVuXXoeQivQqKOqDwABTFOPsgxgXAqOOoe4HP9VPtOezNendB+yFYjNG5
OBCBxCL4fSS7c6JwL3dk3N7mxuxo820iCM7EG06lyVHUVU+cQ6lxUiKLbd3/IOgh95+PBNAbGPR3
xw6bHLIV5Nfiwmb6jVYNvyNTUFZLctPRrgtCwpNyK6kDmb3jRJlYK5BOaqVTbuaWjUcephczNgCE
E4lEDdD/ILZINvZxXlKuxdT0UGoP9107hTh8gos+u5Q471Ko/bwsVRrSEXxC7imgO1QxEe1RsS+V
ocdPieqv6bvjLz+OD06AqDH3wdwOYxGyQGBEJlDrcV3SVfTqmkPGWI4EawrxQYK4hSSgrntqpC4T
iKy90VCJ3IUg+HUqMn1D1hOiS1A0mSBkIa9vRpWLg8p09yruNGHj6jpNPI9IeUjlDAyT/iJZYRvZ
bGNyhOgGOg7arvxP9HrXlplzick0xjyfKd0pURnMvxo4R2yRdwHymMgmNgwze/NjmhlQS5y11suB
/StyXifd5f8uWLqNqxiy+CoUoTAENmsu+pfqkCRSs03olbqTKh2A76+YPwgB95msvuJg3HBcRxgE
N1CgmXvwoN/8vr38qKbXG7GXOLfDOTs36/c3FVQYi3RYo44iKm5BzImtuDbKORY4lMWdBse5E03D
SKU6XHdwQQEzvuIYiQ7Kqy9kBXPKMHdd9p6yJDxPicxYNJ5ik0gGPR/xQ2WpL2MKWeSuFJ2uLvdA
/go1fySBTAExlZKRl/xb2PKPumhnAJS93Q97lfcNMGglSrXfO7NN+dFzejIyoosHSI+jQ2BkBF5K
9Wn+r+ODvI0xAlZ/+NBK9OHxpmBJaSU3QP/rPxQHuaUxDYclRV06iLTUgWEpc2awNC6/BPYbuJy9
BtUQx587b79/UtK3a5rU+h1IiT5IDgemrn9Hr5gpMGjjJrzRoXlPJSDgsojtTlN3/vLg16THs/fK
eQfHgcu+mnpQL6cuyhmB/fCCgQwhduiUNlmSJUesP/S7h+CshsgsA/MfZP5NfljyME5Wpy1uNGSS
HEsxN2AbbK9Lhu6we9g48qW6YzO1O7t+G0UgEnkhJkpPl5ruYFYXTHwcVLzRrOfd9vwI9MzUblww
Zu0NJ+uYMxZGQfF3PP1cpNdFFUzxpuP4bCH7Pps+lTR+lhOb91aK4Nd+/SwYy/KdxwTlI1W+9Adx
chQjuJatbJpLzq4wVubw4egR9Uy25f+RX6wMuk5fLikfW6g8cCc5owvIsi2cdgP6jVhegeTJk8Zp
UYxbhpYY6jIcZyfRhlUMH3qzYy7DaENEAlbS9WNrio9zPCCXULT9gcAPN+Xc9Biv6T7hLltbEvx/
f0W3estLGiUZKV/J8H9phPQquPbsF7m8doUwUbQLSCOb9hUm8TkM43zi1DHm5vqPIOi3zl3oTQBS
QNa7DodhBcZcW0BdC2zauT56KCM9x7R41KsMDaF+iCDjAKiGX1MWuBO3UdJRK2LZY4GX7xtwV3zc
hERcDcjh9YUCVnkreMV7XJkd3q+4qICxId82dj4tHb5xcf/5DT+FNiA1FenWr3AuyzbCzXQl/Vex
uU/anV8ZbcXq8h7ud6OxB/7I3DziBKoa6CnaZbuE9eeq0ti0v5021Vxr7UPNavcoHlsHVDRzNMVv
qXUDgi9U720Z3u0GEuJymyaodcfzFbN4/QyVwIlNqHEn7g160IEscf6PiV9xQcVXgGiMK6omGqxm
MiAMDBKjZ3exhwkCB8GOFBlUlXzRuaFcpnCpMWfAVtyJ5XhfEvowoVvkpucsZXWx/xv/ABQ8W7uz
eIrdbq3edfOHWyHeqedJhwaQj4/XGZuXbmoV9UgLSQOGnxelBib9i7wTbrVn2ILTmfYnFTskWZQ2
1unPr3oOlQhR80JHhci9FzMqdAZbs8DWvpxkJspIos2WTBoH9B4bBorEB77useMXrQeJVphA1U6v
nsrFb1gU7lTYB6aV6K/ZOoswTwC0Ch6TZRJ4GzShiP9XCcm3bo2oZh2t9CfpinNXlvl/B/aR39qa
IDoYAOdnwECNIWn30oBgJEvDdECErmaAsHZtMVPRZv2FLz07/47Qp5O+wlEwGHfd+UoZZEp8Rjuf
tDGmmhzdP7ekd1dgh8RFev5Rnr3bYfVFQ9WS679Dy+cMCqatqAlDhJlXcKTqMkBBmJcNVG/P0eg0
6cQ/KutTPZQA0BSfyk3ULV9VjyVOeyBgiDV5KNuNz8+NSC7QmJK0+hENJizuWZY2r8NK69ilGgLR
W6luJK+WvmMIWo3379qzVpdMrKQoh+gm61bk4qAFGuyVp/vhOkBs7JZj2OI9qtHdMVX7EeXELJ1s
5lQxh+VAMSt0zQTKFkr+FHvuCfNQaj2ILbVDhLvPShWcV4YBsy691jTiHHCkn+vOX4OpWjJiutLJ
c9031ANNHi1EF2ujm6Sw4Rf8tWk9+hkIQwYbTxh4ECtTFEv42l8VCYQeyYMDOR8AydW4jJ7iw0Xp
FVy5RRFjoyfH1N/xLchfahxgM5WIS+Q6BOuUyMhGG8sHzbw/nYo2l7YPoy7Qgn7/kXVUyZz6iEcO
fjoEyWV8qRAGgLfee5f5hpH59JN2P/ycjsRW3CkJtiYHSBt/MWx8MQO5cCpjJgVNkTwFLju9z14u
4+HsViGhZRKo6WwTBViq+6AGreSKaWI/5UzEInt3g2c8LjDBEwn8cPmgXOZdBtfwIeUZ6tcO2A7N
2sq1O1RAx2ffaJ1LaBmzAvcywQn74brMNV+PDbD37sx2fnYSP9Wmb51Fo2B4h+Ljk/A84TezL5kx
+EbGrOjix9j8P0SeXu/CSCNqCVkMpiBuPDQSVzO4xaBZ+Z3/1xDTkHS6SAr6kTHlyuFk6Rcyj4v5
d92yW8L4rzRwW1nv55t2vr092g/ZOtHVIKvov4Lcba2lXLhxHL2oCAlmrFWXfkMBNUfQOyziX4Yu
P8XS0SAP04ITlwcoqLZ8MphPxcUkHG+egkNNvE3VDB24ZyIDVUM2wYrIl1c757SSzsRZ06ZZlTY7
koOszP0AneDb77Q3Wo31Q2vFnwFCamXOxrNbBt0kdkG6o9jeH33Gj9OoGPjvtOVvfFRXjGPYeSBg
FY9RJhtqqclv5pR3cN17DJS8Y7PHf8YwLltzhAHcE0FYCzWat62iAQPr549k3LvbD9+yfNh6OI3o
3OAi49bqag/4/mxS94mxJeWNgak8DEOinLqNINgpNmjGsMIV6cFpGeBJTc8IpT9SjHcEidtfrC7l
lUASXxZ1gganwceGWu5ogicphAzzJjHTrkfrNUfIyWup4UaTWabjAUuP5ECsM3546voi0+ljGoYG
KZlo+i/ChvUkSa5hv7MFvJvpfNuKd5JUB4v+5SJgKQfQq2SMM1Frf/bssCbMZVMjZ5a9f1UpaqeR
ryBTWfeM9ldClSKtZL7yHUOC7lZLyuBQ9Jws5H0lotrqD58ef+WU/EJ5UJK/VuqZO6iWflpdgqAS
l4wX9ibReC75rkCXWDvenD72ouGDFCaKyyhE6C/xQYxtEK74GyF2o/7DS1OaMLMn5InYJuhuTlLQ
bHg0oAHp0te/MbDsI21wjCACagyQCIdgYkGF47Hr5AJbUwyuWrKgDczlyrNbXkX1uuoA+wGUoTrT
anEk7WT7vKa6HIh7+7lQeuvs6+COHG/i7Jingxhg0mZfXYX1ofnds6DTiOX5nkpTURziY5O55NY7
aDibTgsXyhCgoKwj+BOsXPQcB5ppdxBsmxK54VW/z7yJcr6xHfQkEC30pBXgi6pBXuTk7P7DA73S
yhIGjpDTKTacfIW722U+9VD7dgFQvUQVgXaXfgc9exvOVcUILGTEkSyg7ZSKFt2dvdWak8Sq//AH
lRGK4FOQTAex2ZJEL49HzUj0SdTGOqrmMVdS3EStE8g/TcpLQLpwun2musPlmC9n75o6m/2waEb6
2eGqqlevekJF6dWI1OP+QWAIkc51u5ne72lXfXr9Y9WlKkW2f9nH3WIwsf+drD7uw/m/vAsAGOjG
00Mv0gfbBADIGOKaHdgGwelQp76LJdGF0/nb7CZ/Iyc7OBfGFZjdOzdiNQS8PhjblTOvapCCYT3m
8EO4dtYw7PKIU0B4xOWbvzlsmoIWl4cfB6S5NOa0eBdM2TO4mIkRIxaUjhgjEnGpePjykEjETKeR
1gcKTptBlr0Z6OxZv0TctuYPLcR+jFqNfoDevuNwq9N+nqPq/Ok6/kUNpjIYJi1Kb7eyXMC8nRGZ
05h/7SsJVG1FRnqX/qBS0f99slBMNLrkNnBFK58iW297dgdBdVrLgAmWh6sMrJhUWdIRDGDPL0hP
NfOrdp63IqQ5BM69tLSkoED/JcgfwxLFFzeY+o3UZ4nrb2pf6hNjYwDwe0RFzzzJ61iwx2G5KosU
5BvlgNtN6Ob3TxxqiSjFeFWoy8S92Ol5PAOCcFwrrNHehrW15MulmjjvmVNSl59faRMuJmFcTBxa
bulyRqN66PHx+clHxO8AU1YARQEYeKvncMevw7Amp6i2TXjr/m/r+6+NsEqqVZNoTADdvACd5lHo
Uqo3nwhYxPpuJjDncAJCsXNEYxiN0B8EMMkXaQXbt4SktPLpi8UsA39sJvS+InlLH5krfMbwYCtO
/I9AS2/z9heKj8BtBIsA8xjRBRHLrXbPvw1/OiTuZhS5yvDk8J2ivG4PswYe7wgfhSM1kUDwXhkd
Zfqt06XCx54z37Vysomv00MqC0UGN0lOD0ZdSkwtL+sVjDW2rfFMU0om+tyblc++dyg9U4aeHGiS
KSWDE3T9L24eRBegsP6YNFlV8C1zc6WTy8aYpg58+dHSyWXIzgNwtKPJEBZ16QSMDK3wFwoWbfYy
9v+SGb2RrYZ70s8uy36u3urlFQE+FTCgCK3RSAj0nMd/8i93Nbt7+PoACEkFWciMwplbk5WhPQG0
qn50Tfmrz5s540a+rb5SqmyytDcOEuPqXQBXLyBv9nZJBDgNxSHFNWi0yhuY3Y4rBrCh7fVRYWjQ
u+YdyRYFdemLSIfwUsWS4FnMRswiTqr8I2ZhnwDEI/ZWYUzHR+OirnpjW5ADxsZory9LGqPtDBYt
qDeg4nVbpfKhGqQYu9m1tmYp62/ESZ1Xvr++akV0AlNkVJhF1WHS8GTvCvW3w+QwbYkAp0pcfhkw
lEL9eUqOocbIxJloYA5VrWDa+d5Ho888phHKj1KcsWOYNEU9fqOGLtiSRozBunlucHWo0ZE22Sb5
HbgdIa3yaOKW09cmV2Sjv6VkIyDNvPRy4OOv2HSHzSSnh5O32or26iDcpm6RL54uci+L/vL6LyUW
KGzhl+/jFlvS8IxBUD8cDE9ZCctJWIFrC3qEeuryn0Eg+HxjySaVA0Y8u+uIvD4/gDDFolhQIpdn
yVrlDnFpmRaQ266vZsqMyATqbLungCI2AEDDb3SSn9R0YJBlAvrHAkipBW0VYR51gUaHvaYwOJGJ
EXno1UnRs4cEAdumGlRWSyCMZH4Qi8/O0p23WR9hP1h/VF7tYZcYMNixR3gNfvBBL56lYyITZBJL
rlrL9AXJPdQXwf8rrDsnimkhDBYUTKYQ7GHOnyJTeOGB+1++LWvI2TaGo9u6QUgAykFRuYa88RLI
DPIrvwuqYbY+LP95jSzahXf6icwmX7fnuCmGCIp29Z7v69z5rp2xr64f6AXS6vKoT5i2aamsJq2H
TuVEsetUkzsf0ElxOMPq7LW9VoUPBnXtoAoIgLu7xv73ceuw5LiTP5r2xryomCjDt9fplK7WRENQ
XWnUda29r88M+82zdUOHwwfKfDPlJiykL3v1lsS/DOyfaovPdiR2q8CSNefmP49CEpNwixxXXcVX
Jlt+Pl3s6jI2uH+kZdI/Aax/JI/e/byCMCeB/SzaRlxO5JicdmnpCLVHhtrhUgDjoKnLr9S42eit
ltEF8QIaIOSGTiKgtOdCMEdHdGK26i8I18Oz6Sm7OkyzvJPsr1Jp/5MPdku3fFsXkJzswKUBFCt0
KQkhD+GLtyrDQu9XEAconiXSFeyjg037SGhFKBZQ6xW/GS2aP6KG0kegeZEaorsSG0JtTogoAhjW
1A7pngLuD0puCumbHiDAvgqzSoVHinQlj5laF7W1E5dhnc4sjcZlS8dxLSBRHwE72O6iczVPOlwj
XurxFq5a5edK5q2nMXmf3e25sc2ekROQMJkBw9eMzO7dMTruxbEU84phPmzKTstCpUaiQ9Ab2lfI
7DqirEwlKo6yW39WfaHlu99zBSU9EaQOc1ZLJtKZwhm8/bd0oXnmGnyzRL0HzDHanlHCghEryZF9
7RSnYjcvyRW0jMcX6fqjmJtIAP4YgKu861C+RqTmd5ivax9mpalVGYjXyQzWamaZrlNbwJTr4ltc
I0CZnKTBJzKJQHxaRUEZdjx2L5PKQIecnlNQ1fiOqL6B9RJxdqYqlj8LSG8Y4HbNRrxLrgwswt3X
ezesbRBFWGlfxHYb7vj4BIw7uGv+CUbVtGkdz8hBdi82btM/w9EvY3boj5INq5agS8pSXCMY6y/p
Euq8fU8cb1uJteJe/YqYLdYk5zJR2r8Drk6t/VfB6EP22Ha2qMe0T/mp4uJG+2xyACaNGWXX/Miy
SksRbNY3VqMMtlfuCruGZ0vAO+eflQ9B7IjRuxyO0M1BOeL5XajjQR8lMv/Bn+5rrPDkxFv1Ddmr
ovxIm0+aITsvurKC9GYwERD0jxEk6IU2W1QWUvOVcG2keJZnoTz8v1GHOGxDJ1t+GWr0MCfkELre
LPAKF1J/ckHUo48KOtTAOVYWbVTtcCgO7wwthx8YvGwulVHJXcyF/sMfH1E6S/+NRaSkxhoEjnKX
a6VstAuMqvrjS7RIlpWCjO4DVLUwptvAZvQ37CtdgTZ6cgkn97UP4lM/jNFtSCT0YFlng+sXufLT
cymlHFJOarM/B7hF+hkKiSoLZmSz4nYcJvbt/D98ygVOG5nJqO9m+n6ViiNqvPcgKuTeh1k25gZO
pqjmfmxEUsAc4nHuyLOXYoMfjnCdlyM/efuYAzUZmVsaQf+YiCJoExU9lysh7c8RgloQ+U3nMyUG
ELBJk0ZezBZOV5l0utISJmzLVFtWub1OuoepUh1yp72kJ7UsGXNjCLezX6mk/IqUQ8WznlWozQBM
3lIyS97czd59XzB/9RFfoSdS1K3sguLCZH9b3ymFvrnAZomBiCJKBbIheBJPraNI0kkpxkj2Qqds
snADwkaRME0qvnZXwzJgNGfbynjD0w/NgkjMa6ZKdYVtH/jujrd4BtmEZoZHTw8w0uYR4qKTEuzA
RczJykY3WW7aA53AVrKa2n/cVCzTQiDIvXlROpYgW7oTxjd04Jh9HQVkQsOk0SFMB6RoI2ArZcuh
XsQRkj+45z5S+ylBdRxRJNTu55pIumyqnGNug7baLylAMXv8tCotwo8s4DFKFn6916U17NuzLLb+
PJk2hbhXhDhgLqKwCVvMdFHbx8mQ2Ioy3ekP08DyjSDHLHS8ISVSb+7gwwc5rUjDAsznMR6wpuE3
fTSwczufcuZaaCTDXVoPWk/a4fUDna8WlE6631VJE8wQp246lwRDgSwIjuj8Xjik2DfRMlqOJS7K
FtIIdo/gaW4wwySvGwhOc8PwNTCjkNGx/tJGeuzq8dazrXAnoCI6G/74FgV8HhN+hvGM6OAuojd+
bK9PRiEpb3k8en6PeCtCPncKBQLSnsvurPPTiNrXa/MLM+QKEcq6iCh5/2jciOmt1imKMLWFdv9U
lW1ptUI3wBeej2VvnwKajbf2cAeJZGb8yeYUGUYOGttjBdwJgQvlEwyWESS8RSAFa2mhASFukj6u
F2nOsh1RSkiBzh3leljlJjeADZhPU7jHgLzpEOYfhOlvVHM88EWIs196lcoPrnpzyVynyriXmZSE
bENKA98mk+8/wdbBqirMbGS/UGv0wTxk6R9LUycb6E88nUyIFG9iU4cTLVXz52KaF3BZlK2E1sRo
1Dp12uFikKMeN3nc5ogul3OZd6JERrfyGH+4oGPQ1dm8iz2P3wFS25aDNJurGOQGPedVUKVEIhwF
yiQN5XHc5HHBafNeyWjRstwFPPot+fp9tD47Bc4EbtrBvNTO1KnkbiKpJmGZS+lf9vTezUP5nW/I
7N7dWBzdHH0krMtcuA7TX5yA6PRyqmfQWa+QIb+3XoyE0LY3EYAajunozs8bCxP051l4tjq2m422
BDU/vok7EcCJQFaEHjxp6HqnoR3A7elPp3bJvGmcIBtqc8iTrzxy2m/NJewSzYKQtsKyXHRb2dE/
bdEIM3Ofa7nPaRqiqUdX1tMcuDvhRFri8wW3Uowkg1LT7RGZDuCU7ZvjEVIm8Dua/HG2Ej4TucnO
/xR02gHEO86U/+BtfOx7c1UVDTnB3AvHkPz+3GiwaWL56PL6FIqXc2CW+HJdsfNiB9gI6TV/j7jp
dGLa0dLNEXV/xs2TBVx57UtSV2NkZgJsEPw+r3pumyA0eO8s3gxU/rj6ioiHmWbflnpKIMaq4YnC
ewKgPxN8l8ClpbdRpC4Hf6Cw4pD6qiW6PhJfGfvKxcwMjlBlCh5cTOtpU99M/uujyA2iLV7bs6+y
159vMhVb1OTJmcyZP4VdM7Fpto5HSHmWy14K9F7bQ6kVPHuMDeb9kFwNiBnZzqjWDYRp7FtM6In5
cFZWOL3C8X1ARf5YgGKJxNkAgRez4eSmSaYcj+9EJYUpe6FDTng8lpdj/V8eG+oz4YOdNjNSbM3c
86e7CiO1sOy41NevN58yx5as9bE2Vnnl2LB/PVPKYOsIbg5I2taiZlSR41yZSlLjrHxDGncYcWoS
1/wCxqpk8+9ic4KseY4dpDOi2qzw46vmPixb2d1yEi91u9h3F6pZwjqtkFxg8vo9YsMl4nHapYpd
Dl8VfqSPYOHQJa2glrpXrliSGUGVb043CzmPMV8D7WN4oNtC8h+o2G30W7OG6QnGOTcuuwmRM6vT
KENjRBxg5ZFIsOYftXelcVKCu10HZCqRY2/USy7UJoetiVeeSYkuPqV+/xCfF9XMfZOnJ7WYvUAN
J+DYdt/py2D59W/nqcgofc5XLBrJgSNCrbQs7Wsi49xCgyOc5Wv2Yu6vQfSFnazbVMwur4IVBDt2
F90fdIxBPD6P1eAWikCkaXKdk2GLlXdmPQPkxayxgv5hprLl0ZCloKFMKZQqw2bXXrsfbeuxvSLw
WL/tit/X2KCWpqcnTjltQEued5XnYGGToppgb5stdjZbBYTCJtEkGE5k8EeD4KkJb6IrQgkSGDpk
gbyET/3lgRLmcfhqeUCHM/E+a2vbbokZOUqx4MsEIfm1COThIToWlKwIl0O+dXdeHYZzXUvqRf7B
tkoqGm0KFZNnC20t+sbkMtcbsrhr2wzxs66ofPHrWwf5hQgBjZuiNxZW+PTtbgcp7KH33/ZO9xZv
sOL1j7t2+kn1p5Ix0ODVuTjU+Po+7j7swrakwLBUDFwQNllungaIISw26fzZH5WhWbtoMgRDQ4zo
zqYETiw3tuov9J/F4dExQlgnzY+iJJSTRKmoi8F1oFE+aKoQowyUQpbPuPIs8pyY0ICvaR4oOsn9
ZmgK1GojZga0lOtix1Jx5TIwRsniySePOHHWvNXwS14Ec68FqOQaWL1QVDPEkhvEqpoMcbZbeR2C
SnkSGcF1n/3S0EkDuTbWwKf7c/ceq5bJxT0ZDIWO6nKDu793NjJRr3n17Hi4RKxdr4bIGnc0jkEb
iF6Pn/ztO9z/OmINmuOx8I8R8EeUvnx1z6eoG3RhjGHO3tqlMOzM3FiazExmhqOSxk2IGXIbuhVv
mNr3Vq1ipQuxQz3r+3uPRNaU8jA0JmwXj3i8kTViF0mGJC7f0b23yisfM8f94+FsxJponb/So/Ld
J7Q9AvloPwKhsqUiSUT56HzoYUDdnBE+mDhgNa+prWaDUecCZDOfmkmR89I3t7/V7Ei4YJ2HTDwy
dII5+XAKHLqAOYPskGpaNJDxeuFBgX1c2MLgzbhcwGEJnGFKKCGlzvFyKzriAcFdjhRaRJ38iPOK
hXhWe/QuM8Zps6Zgo8UZRnd/Sk2JsDtQdx/DKy9XwBoPzXt3LvRBGXM/8krU8LiAAd/reCNSvnFH
uGosscwmo9IKvOAlnNRBijThCJ3iK4TzmFVBlRFA5uBbscjw5zUUpQy/c6PHFeHSbihYWTJf8B4C
1binGyturjG/K87jAeO2WgMSbiqi/bG6bi4NrMk39NZNyUUmsxep3IRgveA37C0waUHeUrYFMNPr
ekIT7uREoqErlfZhr0r7LCx6wN+313+96vS9c3R/4BdyR6TlBHu6yEQvsDo/1UpeNfOPjZ5SC4db
CnSu+YZ7bGzGtd88SlfgvOWmjlv0ZvAr+cm4y3Mr6E5anBWkAwl3YMxusn/whNzBsLfWNn8Jwz4r
6kK3PgWIyNQoDg77FX1Nhc9khSEK3SXaKrfzsGGgiqEhzh7fyFuPNujF590YRF/7RuSaZe3DxrG+
bcmMJ5hBFZ1PWy/eenwce7avZR8unPlv0q8dXa7ZweVbCxzZpsyLts5kkbN/kjCU1K1xWeqQ7Cxd
uFMkgYoDObPCLZybz6Q94cvJ6/yHhDjSDfM2LpjetXDRaxQjOlDpGk+HLN35Tk5atXfgjqXhQgi1
t4ax60x4ntmdacFwCvLQKgRrnOUXWlc9k7hZlo3B3rJkUzfeHYQKZnJ4N958Tjt+/RLff4pUrewh
k+3ms9+dwC1VxbLrroZauvWVKa8y9pvuLQFMlqMaE1PweYaOGMy6myA3/vIhbG/0CUR90V0GkrdG
zJ4Gthn7EuXsPOgcSaGXQy/RdI9ZXh61FeqFfZ/rJA8beMxDz9ZqZPmB0yNn76lEhQzQ4p9bdaMe
wYzJSmTzzGtV9HX2ILMZaSh70DWBJYgaCVckXlEIvPP61nNCUZDrN7HrzrH4me7NufJ8sp7tlACg
J/vLEP3E2l2bh0FvDaR/1w6MJXg4H4pR5lXUbrahHQNjtfHZWpUvXfOySP3uTuJK7SQmtusUGGGq
jm9B6JgJU4Fe43C997puMcTIzVr2tOToN7NICQGKrajBy5CLr9IJum5jVAPma6xLyipdoCiA6uj7
/OeCVf20a3VVVpQ6SRa7SjMzJTEaLfL3gtRuj8SJADDrYvdOawkSNf6l3VCQbpmNdCOQ4Q9UwL7a
EKOYXpzv3DOfbc8honsgp+iJT/FI8zU1wV+GuWEraS0mJBH70dGbW1Jr9qRh4aE7KRXTBHazeRef
SMtmURHHHc2GCBhuXVA04/3Fkih6YQnwttyElQqj88wyWVevR+/6/65T5vc5F5I9xjGJVa8AuIaJ
6oBLYyKXPtEJpalvsH467CGpyT1gR7REWLIamAoH2a4g64125SWk9E392BWxsguBwHRDAHt0oJET
Oa0AnrA+aA8GakasX4qTd87Zj/ypPiY5XD4gWLPfjeWagHAdDUi1Hgr4+2NKMS3/i/Kl55WbrWd9
oGxP0eQWuyrz1kkl9x0QQb+yeBF0x07uS5hIju6PwWDBnK2X+sGTkQPIuqjQ7k1GBbPeYLLbrhaK
biee+Dtd0AZcgStLv9t3/h6+BFMsP9cfmnfQkbi/ThEFpgzauEhp+atPR43X+d4sGEURRp5aTjOC
amn+vJBNzRUNGCjyMsyzYy1iNF4dRNkvsgVBa1YAzgy9MVHlY6yup2ZgMidPjYZHZoWTxSulDOEl
hsG3Sx7shJhSyeiK3M0wFbRnOp90zMj7aAk4qwr9AFUmolMPgkJLPK6jrvh9VKMvdfrNhhHbVYrC
fwHmg4KP48PPYT81D4kid4ZMRdgO/GqdRzEPBMs4805gvPe562iVfPfdP0Zr7keyPUN3gFyCLBES
60LdsF0lLu9YFa4GH4aTZPLfc+rdb7eJfIIc6noY2RsK/M2RRwX43mU6UjhJTy2AkeyulkYr+fsz
B+FaRzHtWxt2KCwHyOs26u2oqouS0zztaWe5vlkm4xgMsLv+kK8d4/va5kaf4Qphcf6bkyDt+uru
4T2sa0+3VDkpPMp5AJ5DXVu5gx065+OwMzklNqGBqA4dO6XfUgvlQGauhUyqZVeEH+DI09vZ4yD7
oHGAdOj3xQUiZBzI0GGz3vPnu2zaBxzpipG/iAAhKuLCViBieaAxBD6Xvbbgyq+KZ8MZtfhPDFyl
6V4LIM0sF7YAzNPJBUGVl6kzs8yrYKnZ6hILDe53TbGvAMB0XdDHfLU/rPOKoNLCKX9H1lqY7MfZ
he/bCmjxP/kgcZ6/FDODo0DYsMkWF7CUxUI74TUowyFPlM6nbp26Qkl8cMNJccdjAxcSbMyDGNeY
+P8LcC71LxBF5JsqWXgVK+r8tmm0mhP2lgLKHaHQlnfQcQrqGxcxznIjPZHMDy7pp46ceza2zsff
Lw8OkydJAGthgPx+esxIJGcJsxbvSDFC+Ez1RGeAmmZ6qZf2QDF3I74eusawYW9YbD2nDJJlUdA/
77xzHmU9CiJoDrCWYFFxhHok6PTss6eXIviTPjzRII4ATHh8e8pj4PsPCSBQDSUJS8dZ+STQK2W0
+6wu1CRLHIp0UCkj6VOfAeyLgPiXtyPHqVMINoDsmof0tX87Q7ZuIbX0CbvB0X+NxUV/Mj6yK/Pv
UIaXLvZCDbe2vViAreetqn9/UqtapwG1F2LMfi/FVEGQKjApuqJu0MASmyz2UiKXsvOhriLINbY7
+9+p+c/9ipkiWhRWsgEnpLHSg9FIidhEo0Vp+bVvArNYnwo/YcPsUXYi8aQ1k/RrQfNWYXUn9uih
8+zhbb9WCTxBrOZcCULrL6/MFw3cE9w5mwPPKExZhI5d8EnWSnNrofp+eGmKxjQvMvJA90DCtVvK
hUF4CLQeoaWYTzKjapl4GjBCEGoTC0o8vcnJY4x4Vk//B8AHLz4tPeERtXlG1mzu3tXcIobrqU6C
E4Gu+13tfEOezqE9TAmxFcUJcMNuIF9VYKdCPldX9RguR/C/G20LLxhBErj3O3jYqzW7s3Qry8v3
HS4nU9x0K6a7mlO/3dXW2929Jr/8MwHttHG6zw6adtiby1OX8/7QgpF3BOA+/HWOH43L+c25f0+I
C0bOTCwPPAxTnEZ6tBzzWqrXZxLG7S90Hab3zTCbBand14vp8Edg3SsRa8Zr/W35L+Ul6wLxylAH
vwdTuToQSjKXq+gHK6xINE7a/yXlPcaa5NGNQHKPJPzv/Bi+zF/bQJF1XuQ/41e1WRVLZnTs78sR
Q76x077z7EyVCEiWz2R9+ytHlrC1KrEMDUCx4zus2/ViEB2pNJ1euyCYH1yuKkUG7LBTQARL+CtS
ITRKzIrOp2pnd7KaHhxyAlsCO9FlFX+ZxjvyRIHf38OB+9UhKGI5nUTBKcPBcQ/YEdCJtOfQvZI+
b3RA5I4wRz3TgMPL1kJxqL7MpiNAAE9z875imbJSoxJAnrWA8e5DMhZxlWGEiydS049v0Glh8P2F
u2aTzeuJpOgyaGsnMeq/UjIV/hEroSm8YlYetJ9kKVl1VO2EvdmMcvuFGU4wpHCTVtiY7wHnJ479
oI4QjzaEJ0zvGp+CTSnPtCmC4E9fPaLcCF7srNNsQRi61Mg3oqCosIDmRN66QSwE1uidjEJcckE2
W2HK9JoLl9OoFnzXprHSH6gvmEJbSqPjwtFTSKptb9y4LzgVve4VF6WVukBsKBmmLasZEV18XZM+
otfhGuo2K8wPeiDvVGGfC6pAwde7tNs30RqnfrSON6X0TP47qcrb9omCq6jaPO6kpkVbZRXcNdYE
l5mXa6I8BcqnSZPJl/VHEzpDbqXG0nOoL6d0ZLA8vc7N6mX2h4hSfP+X0IcwYa1Sq1U9jUV7T3B8
VJKEw5jPfxx/ZQldCkkJZx9ws1RUaI1nybQnQERV8sIy8WYuDy4l9FGiVBdzcAzmp+4Fiuk28+u5
tKtWChEmTIV8DMBOVSR8ZrBucLVPoAbNKvBznmvzFzOxhL8T58Tld8zP8RRVAN/uzwKOO8vEuPn7
FU9x5iFDXdEQ4V5VZMRHFl7/0k3F7iMwcjtKoN8R2yeJ/X7wwvsYwKSr7b/N2Yu2mLfKbjK5NbnU
++GTXIuHmEuJH+eVEXMsOrAtxqPtltivbwocRbnGkZERMnT+yfdfGIUmRgKTDe2YqoBvnVLbtePq
sNVFCvKCfykgiaciP/u882RYRzD28ZI9lYWtsyGVaVqc9uRyrwwMWgS/g0xFs5dtU7Zmkdy+L0Bp
UbfAi/6JDhuZmJLEEXfm7N0dgL1emily/cZzafvzyxUp/l9iIdjo7X4xbQTyTsZ4D9euaTXtsgDr
NIFA+u5E+p/1sXrz2LJfMy09l9p73i9ajiNyqbpbHRSzPAYeoVs5d+adITPXyMI+YEEBIMvDn++E
i7w4L9j5noyYBwZLX5pweRWVk78ehsPxfZtu4GWRAxJvjezgs590xZrFEKNPZRLJV6FII50Qe1tk
9NC+Pbg7dp3FXb00OfPXE8EUNNoVjQqsCGRJFzOKSJ30ysZxfwhei0r97+cc7ZyXExc7EVd/k8AQ
c3E3GbPP+nMhub8tDZVf8PtFSnQiPHvf/kettzBP7lx6Mpr8d5/wHNULQhsyn4iQI3TKx4qioyMq
ughwBXq8grFXaXi+c2WNeLPsZYgcBIBOVlyW1q24JATC4B5PaZr+9+MyTkVSzS1Rf8Vtx6N66isK
j4Wp3pE0i00lURC71KDaec30vyUTfDXHbPTL/D6TvFAi57DCQhguMJWlMQwC5+8mAC8d0yK5Yj5/
72MRngHiziXu9NpFYioTWNZOfrwBAYfwSCKivy5claKtbf23mijOUbIeaEHlYBlhhvvZ9qtoQzHC
g+/SPQAWWNlFzYBad8FZi1OxjAyNKSpxE6rh8iyBpPYT0CXWWJQKLwRSIpUnFd6+HKvljlsPyMk6
+LXSi7Xp0m4hcauEMtEqxLshJ/agceCiJF1Bp+nhQ49HZiYr2Rts/bBs6eg3EM/ZcoyDVn7RjhNl
tHt/HCbK5ogz6K+xj/5IYnP1SvQM2AklGlutsNhHaSJc55xSobztxmaeFvg3fiUy9kmEf3KXYXHK
cCJVhxGmGH9Q2CGeyDhQg46klI9/agvxg2PyjXKBikVq3dMoEy+42tNKLB/ueATuUIPkrl1OuO5J
NJTEFJ+2dy+A+aHRVoVL8FAg4beDgtTYzyf+qC17XZ8Sm6oZMWorQGgxhYo0Q9zy5AjeDYpWU+nW
c5QA0tFAQV9cvpMbrAWChCmGVPFEGRAdB9Ro3ZTxJnMwpO0W5WlmlssAMxoDfEhgprLPXoOdlykS
J6DD78nWcs5wmtGGH3CJEuhPfyX3QTFE3RJX5TA9H8i0E2qA9Cz0rlGUxs63V5cgncKZ3rrInWn/
2zzy/awweNCDzOlYGIsYvfryq7tlZjoyXGGLz4nipsbOoFJK30kHGZ7IDk7WYurV+lyEPv9bcuJs
8e7MZKu65fIl8ilsTBJu/GW+OXfP4qQ8jM5U46aY0ktNhvOIL5reCoXijQdI0oKrUYmoskq+HXGu
ZgGK+cqzh8G0/xUYbSq9pwc/Qi9nCm7m6PvG+cL8MFNPMIBUJcGoq4D+wSwJ9C8qXu3Fovhv/PZH
64ZYnbtmRnrrHGUBuSBRI/kzj7pyUVCgNYenBn42E+o3O0r8HwdqR+tL5p4dHCh57K+hwSMP2wzP
JUfftnGvdAuSmknn3TYoM574jHGj3355K4NPzBepni3ZjLTS7aljShzsX8caRm3dRcXXCnTp6mG9
/eN+JZMZkTvlfflh7KFKIBGMipIIZ11E0+GGd84km/lq/li18vPPReqLm692n5cNZS9Jh8xlLYqn
wGAs4H7ouHfzuIszXNe5b/AUUyvrw8LLoO5AnvtfO82c/2odBIK30P1sqf2unsBk6OllvfZC1R1F
fadZZndg5MBumf+QDRXk/viOSgUjb1slv0DKabfhtQRnJRDKNXsCzjsljIDy9/zPO4a0KkHLEj+R
oFeGlVuQpD84XDYpZ51IV/19zyKGKORLXnqsSZrx2kktXeBXe4LEs/mJdLvnd5TKUjYQf8nlrguX
d/FySg2MdGTj1lNTrjDfMNo7bb99KHb3oW2chafMoMcRZVZ2rXtwuM5xQ5Ea0cFAoHQ/3+jCL7ef
Kxyi+8V3tRCdBs3RfZfMgtaFUkPsmkWl1HOPePZGm6wXaq+BrmpJC+Dre80YXcnOsZUibeTudn0C
pUAj1FfE5+6yv/uGarp5arQNPFNynTOI95MAZY+cGsIoj2GJN37xJfo9esmpfPgGSygWEsfrEXmZ
TiDCNlzQB7p4z0cOscMTeLwLBiuENdcHECH/Y2MEvWMz8pnYEU2ZdboQfbIgU7lK2/Jx3H6FnicF
LbTI1yI6GJcFrlN5zqgQ4CpXBVsLUd5R4Vrhxr9jiGdfINX1nfp1/E7dLuOuTPZp3LSWJFQmcfh2
tJrG9etVxjTw//HTfIbENKf/q9rX7L5BI0TJPWm7YRUjc/pw3SU1EPszeAf6P4F8PlC4HtDCHPIU
Dxof2JaDbIkmyvjDa9KJesuQpzN3IKSyZ8AvEHeb48CihD6tg/SYkm7iYZSkmyttzbJ9OKp4CTtQ
b2zm3sNgqaeDHpi/QwykdFNA5kRyAnaTuUAOTTSTa/vJHHwt9UXW5Dt3qtjC4GKdqu8a5ZJk4T1n
3b2GykxzhfSamGLtLmrb23+/ZIu2CkHKafXMafg1NyEOSOnAmkdb7GPF71xaDMDl02ed55lNQ6Ma
NXXWxZGQaq6tTahLE3rVcuQmNtaAtLe6N4VJISGK9xL2otedJ3G5dyPEOr/XyNHIcEvSQ6Rusrvd
+s87nOEQhlQFgWFAgGJ+kNQ2g0xFgvOBY7QLh28lJjSo1wwQ6jimhO3dOJTCsEhY/mfPsCAcgLAU
mXpihQcQMmrCeX1Fs2L6u0Yol+sLsrGxQBBxU8GHvvfJla4FTp1gHb6GQI9dNkG6+DosGkWNLcL3
oGUWiV9SfsUhB0ftYZQEcHPJeDXAF1esWkAahXO58fGJQGiporH3A38nT9lIMHQmlMJbrvNSnxEJ
kyTXO/kD9hpabBf1Sb5aSAd1GPVzVPmuM5j3Nks4z36aJIiLoMpDpe8KwprtUcmShk/GVVGxPtTP
1A/5KRZT85K4qoLasUOk+7kO7LCXXf/QFbWHPHxlPFw6Vi/BJfxOO+a3qKlRiW0XSI/f8eFrk/8p
4j1PsPg7XTbcrSmkp2RAdxC4OnVSPA+R6R77pH+PbBUajwCAnM5w99/EClhvM5R8C0wR2QBYc9PT
+jtyvhLgWHIeQkgkJbX6CyFkUr7mg4BhxMHoA8tcaZVWoU+mPaHnZa2pSXCj5tmRa5OB/ah6WXRM
n6vu5ptIXsvmiQ1w1ELGCS2dtsrVmHrltFV1ew/scSwIE80RUDCy8qVAz7HwmXMuMdcbl0dgzWzQ
fiZJLzTi31qR9fsbNWgN3d4Km7aj0tM5pmTwDrP8CHvQ8hm9PJ4ZTX+9dinvWZ9ESycgVWixwdl5
1aroLKxqoKnfsJziQKWVY92lG7jQxIk4znUmANCBNkRxA5H5QaFDYzL8ZyT2XHTA/Ly/bKQHWgtB
mdLDcA6hz0LxMFlPCExW+IVadqqluNUTmmWu/ORbdR8X65xr9jX3fgYr1Iq2okZXhCn9gHVAG38P
k204tz3XAnTutNqbwaOdC0ummeSbNFGevOniibTtKtHKA8PFVAXcfEvVYcLqaeYmsAp9IHIoLdeN
o8NyIJyRpPsbKPu37GgPdkS20WBo4/doObZL3MQ9L+r6+IQbEOQtuYsRM9nmWnf7oKVzydIPWFov
tZKr3EJNgSEyORDTuq7tlz8oWHbwTMLPbsZF1B75wTUcEMVsiMAHMuDI4jY1r1Rm87SGMXehbdnm
gziQqthzlathre7jpwMse1J5BjRCDzyiOo4oFgDk6aZZVmD/rRwsWZGTTLd1iHRZzdNe9IronLIV
YU0d21WRlBwPTQRky6cre76a0WZPkgFGE8FDfYqDo6x9GqghKQWPJE77evI0RGABioBhj3HKizeo
I4inYBVewIZjlCgh3RJ4v4UPq9UGc3gDfEKW23+HU2bEjK51vEXUaqLDaFylcy5a+CP8otPbDJpz
ibUP5YsVLFSp/UQsOgVjmZ5sxto1vDULP/kjZMqGISx0vUDVCn9Kzo70k8y64SxEOLTnejBgnpr4
ZBiH9WTJWgexg9O/ymTPDDKVIXZg7evdTN4E8yHfg+Q/kkiYNbDGoCUGT4q35bkNNd1cY2Jcj5De
GDH1pULyv7/U+f3nJOR8G0hXeCfpi2JczoeQvCerxbMW1QuCedNfhFUV9AfOfzWpPuLyh2te8pvL
gB6ZlwjHL/JLudTf62A/L5Idiz/CM5LFyuaCndOFt/ehXFMv3pyvUUD2MTQufk2r04QukjuC8PDJ
g+i8S3ANMTXpClbCm0u0xE2KieOiHKPgDDcQcuJUm5Se+gphSkO5Y/1MlYws8zv+MdbkR/LS/R1r
YKqnHUJph2R+1PtYsM/3I5YH2zQwOKwFB/CyzQx/fMTGvtJaElzT3Vc82w9tLS0zlsHwxh9tvvqY
zn8Dziv6R6nWeJ1YsTrC3bbDO1+iPIkeEkdwzqU7VOQEzEPbnNho9xKmQIkmV538q/8Mp1x44q6k
rqzTTBiGSDd8+I+NNjXHNw6bWsXociDDAZ8ZZevdHZzbr9oiIJkD0+HgxrTSoyrk48pZ34j6kjlc
haHuzUh/+QZsntjnj2fkEaiJZNtOYc0BUxs205r5hk1BXA9AsmuYK5fXKf1fkNpShg5HNDDHjBai
lxdIou9SVbijDpWbHId5NjyxPRC8fgGsQ81x5ASmR7BX1ru3HaVjyW+iZz9T6gcmXyB3zkmAVmPz
eRyzexqbSshoaPeDvHGPkPdxKFzLhim1yJaNj9RjFmhnmjSR8fRGcEr9GDovvXEq4ctZBiLwVw6q
i5kW6XF2aarIcfTkyIKMEdgwgXo5gBJuHQ9wARqHsrovhQQbqdLLaOZiAzBoT5x3ZHJo/2Sk8BfX
2aJU4vVJ8ELDPZfpWUpZN824n9FpnpyOOOnSnKmzYpCQLijAthdL0FT8+AQBT7M7q9ScEh3hq9iT
kPMUkmsCZKwwO+PtjsEpcCAlnG6wxnYUL/qaIVTOKQRcTVu1RCS7iEiiiaQsHBlyZcCXbCKADWWu
Ht1Oz4UZKcDuPEXtghlWslN6TWt/HyID+E0EFWGOV/Wezo5Jxi7OgkIV7BmZstvol0apHZLVRcbM
pezZglm8tera9TJHKmVMUernLhZZ3ZSBwf8ogrtApFDDv2+2BucOeSubturAtV6NwGJxzuTHIvrN
ZJFlMeXZsfa7h8yqiIub9xFHm9IY+dUvDR05BywtavZ4rkdZomsaEjA9XSJRgsMNxg/9KvOwKnWK
kfjF1kkVS5M9xVzE2D5JOG2KOy/R086fkzx9+kGByLpNLnDWMRTfA9webRoJUnSnDQnsY1aZq6Bs
AnvLApuhT8/cnLOXQmoGLlG6QG7L4xP2caayjfdnk5MRaMKWZcssZU9MN1EJhhy7FCmQVVNJMbGR
QZ0IAjhUY6WBpOklh4dIrO5h8tZZVIqkox7UzefKF5eaFq3mcJBEXnoBTleC7v/9RxZl4ZRw1aWe
9h0Fz0holVExltQp7zv/+uaBYoj9eLCRlvL+Ctfs2tPfPzv4UuFy7r7cEx57agUfnKIgBfj4tUa8
PdtboNJqVGnjSnSu8A9+x+n0o9riFR250MwCClPWimKlr/9U+HPWuGFT0GK3rCuvbRlB8v/UQew+
2zU74UhmUb1nnnAX3E1DuutFXfZck3hy0gIAKFn1hSsHFTaqgfhjOqMYMVicWvE1MScwQ+YLFGPu
k1mnoVBhK5RhX9QqAzdLidEL3BsiSfCfUMxMEVFbhtwpmfT8rs4L4W5+xvYargqVpvugdbB3FgF7
XVcDUQzBlu20kPFn9jp8J1YPlSIDxUnvCDW1VcHhSrt5MNkLU903GWbUX4CoDRC7WQG9GQ9xtyzv
yqhFQ92la2N/Yo6J4SN4wHvQ6bO9GCB980AR4UfXy1w6HOjU2Ir6yAO4UEm7JemDA2h8lrYmxjh4
Lzhds4js0CAyhR34I9rIt31dHoGDd/4RBMaaHoFPqrrXAl7cOsWPhqKyIn3pyaX6OjfTrxgc/9Em
TKSBeh7OekkLTj3Y+SUVnNRp8l/l1h2+0yNfiChfmWwjDO4jMGAUKgcVG44oTFlYIW1f2Sr/Smoc
8M40kU8MSSoN/VZLm+RliLJhX8tudxFYT/RPNKdlRZK6Z2VB1Ud7EYfRTvQyyD6ASQ0APUwQlVt8
H3UP/TCFSphg+yWdJZZxNY+/hK26BQV2iRtdSJJ4OqB47Of0ItfWJ4+wX/3qxz0wTHxUVGcdG+1Z
risxZK6TUf5aiyVb7kBCTyM8Cr2XknVf+yIIdT3OpiM2IEfODhaZwR3ZOuP1Hfd7izQnCIwcEGIu
CuYggSOSKgfA9Lqjl8eJaUXByLlsMxexPcDhKemv5sp58zbsYzDDvr3nxo9159y7FM1TMRwRp3KW
HVpU72tO8jbXWKl3tNQM8Qqk8xsrOp4Ebsh5wHo6VCWU9aUowdl2Ww6kSXkOBSHyEgyw471OnS7L
H4PHrx6BLQQbaxKm4CFAYCrny9cCRWHWiR3UPg5ATxhpdarFToH98PiSKJKVymfAyqm4hsBXcf9h
3lZOTG+gDDF1rw0774XoTpdj4Op8bczMmVHxg4/Rs7kVysPHl3Z8sLeRabgYzZTCpoSrKS7YNw+y
RRiCHs7Pm3SEHtyBHrE7KUZHIs3ifvjy+a4AJR99PmK1d3lLA+MuuWa4avRVyb+MvYyhpeM1i4Bw
uu0Pb4d6/Jqw7kSP9QnDkU2BNgJMyoBVYxUgLNN5btGjYjhw8bfCTeaLNcnXKiO+PaUM/BPV6BLI
b+Lv6q0sPcZ3C9oF2z5uY1D2c/fEL6wpEvqRT1SB4aFzoo+l5sOI4y0lx5Sy6lPL76FRs5YG0SWt
D0/fTQErXxUpZPyyljC+hPCH70bvRvbocSEPHlsoLWhzP8ebon6ezDSEa5uS8L8LUxbg9EcnuL3E
poNTDQNzyOisaaw9Wb2INBNaKLhx5kFPyq6bFR2OEBliKHuDclqnZw3q5r6hyEkuv+hJji4D8az8
lTnvaQYvWdko61T5mSvMbc6w091p/Q1VMtVA6NZEn8GQ4ONZJYgIFuDhzo28nmDWvimVA9fdlEkD
JA+XcIZBWg9/8IPEdCQUbkblKoqZiMUha7TeuVEtIn4z1+I3JvdVWJmB2yQ3bKifRXwp9xNNffBc
sIQbUnXY1yhx/xY6vhDdWyxLb+aWkgdruRmmB5LHt3UM19WmVn0ionvHZ7+0DuiZXbF5blJ4ifBB
M42RyhP+EXzbJ2YD5o3hi4Bo1vZLH94qp6a8DKYzrR7tgeHlD8+KmTh6D2RUOWsx7uosxyn9f23k
C+kW8Ve7cQ9VI/bNMQ6/zZCqEWXiZK04XXSG8WNO2QpSRJrKFcW29f1gsaLQOEoWNBMtmSuf1/DM
EFrfaTRYFXqgHy6vtBJqSM2UPYeGXqBDpirzqDX6BrBOTq9Lzo6qmxRO720JVUqtOsKyyMp/5COE
cLnaQnZIUbWrwP7VCDhtop3S80wl50ET1bskuhboAOB8wySgQCPalwcGIWKA3qT/fi8NDO2sHuL5
0unnts4u8gxSjtHB6OYQV7tuzfXkdeHEaQffrwNK3FWIQfGzlfy0xxv1Q3Pw9zgmnv3lS+5N4qII
DxYk6qS8d+EfZISTM8m0lpDl/GX69jLWg4co3TJprRJM/ntNlzS5KfrYrwSN1z6CU03Fi8WYhbki
daBIaPp7rbrWzf3Vy6RzZyy0VD+pGtUelsBFMmYEUG4jJpCB/hMnRB/LTKWpIP7TwGcuiV3tVwRH
fV4Zvy6IZvsUAQCgS98vTza+ZXYNCCdo15OYE2poo6M9Jbk2BUVuK7mi87cdFBCx1QYSPbMQRKlq
0Sdi9rZ8wHJHNDr1St3I/+winQD8DqT3CNL/RaNKksCzOt2IDdMSywDlajfwuYzqvK/5RMFa9i2n
nXAKOgCpMGZwIBjKNDHf4CBRNxjTdKIGaI0QdqC9dnzUUx+yGkndltFh23vTxJKLWfWyrKnAUNFC
4/Bl4P5BJnS7kyCb8qfoG0n4SUe2D5J+Lbgy/u53U6FZTY3FQOkWDrxOJB2V9k++bXmJIE6V/3cf
OxP5B6ngcpjTbZCPvqbFUROyK5Vg1hG/yBhjWNnpF6YYcAYlAnpJJKeyexGh2m3sxDpBzhAYJ3eS
KBEvMTlNXXotmQZMaALJNl7QwFVqcoJWldHS1HkFIzIdjgL69t6fPkzViaLBlubh/3BO/NOPtBMH
RdODRzB+PrYZ+pr0MIs6UH5E3dGXxcFMcuAyd9M5L6X97FSJ+RaQ9sOIXeTJZlv5nvjOa9EaZB2Y
/ufWgimWYAJqxs0JvzwEoWkXua8HC/KsxbOWuXVQtkCkH39hswJMlsr25ZrWR81ftiqF/XvfA1jo
CP7abRDJ/IzfpciVBLHzAkCbLBg8tK5UsbEhnH5pzaEX6tZV6ySyXNnCWfE5sFvH1jxBJCeoLMD4
UZrpyZ++SalM1R1MDm11NsDvRmeujVPGiR/CwtwEtUh4UFbTLuFF2kNW+0ADtO+RzCILc2Of60CL
0OhJCLkAkipmmMcfgI4IprSXVZRrTH7JZx3nI5vNqRV9Vbz7o6KW7pcWx5C63H6X5y6sLPxJfUxW
Xr34CxCGyvzXLuqCrg6+R3C/KXCSq7Xex4qoMWkX8x49UP+2ZLx7Hhila3RTls3NJolylXghNlFM
HPIPI8+HLlRU/nli3DIva4A8HsVa7iYMxza5XpeSVo7ZjO3Qtiq+XDY/19obOKAQgrNNHogd47UK
87s+MaaS8VEsW14jD4xE4R61f1/kDWo4yHnsPZevLxr4hotYpLQgK5YV8Bb/MdF9Xfcb4RyYuEu/
GWq2NCI0+DO3tCIexhOvpQND9XmZwtzl1tWE4BWlmLu9PE/AMUAtHjpVarxVTYPbhV5Doo0pfvpi
z/9uqMNJL6UTPJSapjbq/0wR/y4YuQcICE1qPhaabxs3tnd1tLVl6tCfntqJlJKzPukj7cAzTcXN
E2DHpdFL8zqk2LdlteSe04ZLD9eCl1fmwaCe0KaZ3aG6jeITe9rXy0bOtVN3DcEGNIa7bFpmmtOY
q1C2rAOEAOlCaKZAVUYhfY5wDliCt8rRDct5rv0h0gUkyM0or/nNTjbrN2+EjqeR4zV5xPe4dpp+
0jvItE7R8ouS2uxN10AxHpHsOR35sb7eghohY35Vtu7aGBsMVCSctnOEozSzE3netT7GGwx39LXg
KSTE5tGxFiK6OWUpSirKESyU8/EcVubCB0KHrn+TjyEN7FOu5fG9FlyVyyLpgRLrvN5JK0cF84z2
d5QVm2c5e6Gr12kW6v9Wup+/lVohEh7iYSZCNF8KxyUFf4eR5ev5jXLyFx4e7LZT2a90u6750/uU
P5kO3V2a2JwPusOZJw1Ksi04DF81m9OR0DF76C7VaBCoIVv8rT6gymAfJRxbsZF2UdXu6VfHeDsB
s/g0wcjpnhWk2JIuoYOQlfudgN7k6ukqHPfLKgcIFBAXu8mgCGdtgkyJ1cP4TELGuQCsRPCSH2Wo
fSXFYzoN/K/dcxXuVrqT1sLXRexX5A0xmd+O24QnG+FnIEOqTXbzDuzsxYToUUM0qTmwWwnpy2Th
9JdXe5AZNq2ah+84l+LVKzj+oROnKL2SZ017raZJ9KQ2GibDJdglBpBK4IbUcqGqFUENfEMiqtJz
6No7gW5SUePgyScGWmfs76q4o84NTyNfeez4yuAA+lD8wT3YGfr3WboFaw73jc/IQJq/CtWSQtCt
keQUPFXEkwin5zKKZeDhu5CuGue9JbiVqT2B2laxLTexgyfVpA912r+2erdZsyThcbhh3fIF4dFf
IB50YIdqBQHQ0CE5vrQMJJPHFtOeYoJ9ihSkyBAOcZJwdQFrFrzKGAxzkV7U4yX/HGUTve4nnHTd
eUOoBJrMgDVUVuzAUjZ1GfnngJTZ40DUUDLSGMuGAInPQX4JX47jz/4+1YGkb8iNmxG8FD5ntm9x
Td7DkwBKO4XY7sdwM729l/OkAmHgGqqXnN0CRjTJlEzWc/rqbZc/mhMhnsfI4tnIJQh0N3tmArQ2
Q4yAF4wkanVYgCheiythCLp+qsjfVo8Fyk2ZQ2QYb+lR+wEuhWbTz1xNenTPc4pxTodJb9z3nda1
54CWLERg7odBK/8wize/3oBmk9kiQgvhwjHsx/nvAdR61Q0OZPGbWkbWzlZZaUTaHIMIOttlTHXb
OigX799h+BaYQ0z6ZtZhXmxDFCbm4yeU0unj6vxvkVm+uMO8NvAuaWoAf9ucp9Qw1L4KbS5SEL23
ebU7u7gXCdT5aPrbu5zbfsX8lM9JutKqeHA4Nob78sYtby6n4sPOhlnqUyo3ffA0FWYnTfnkzAY6
wd3lWkJ3i6C82e71vJN1UP4Hea7jDDw+NUhe1GEqjRkfmCfllNDFiiuEgJqqGSGLBc8tPsLQdmeM
8+CAZpSv1veBZQtfgktxaWcieMPm7zhpWaHlQ3IX80nT6B5WjIhovx2IgxNesE/6HRfpN/g4L/DJ
/4ZmCdq1AhvpE9A50XiWz+nUbYLsXwpCaaSoFZpthIDBIrl1FY5ieDtE47ujwQNuW4cGwGBF/2H1
ktwOZ/e5UaYM6KgjjZM1JBUIc2jsKLX+6tlSxXFzIdemW+aARaT1bS7D+75HerLtwxnIgFekIMPP
S3SyIv8h49AyqLrYtJU4XXnIy5Xj5h2YjRZXAbsEVug8rwvf8BGCRCaDJO6f18joHnx5RCo87vD4
rtPOtp4P0XETHHL+RDbU0tM/LqhKd2yAP9c7iX2CQmT1axBnjd/DbJA9LVTFDjJ09y//uOkCPPH3
BM8Q53BikWoqYKe8M6aZsuEry358K2lcDzPBqRTtqs1XLchiG1Fnyeykqu55BX1fwqdoG7jfEp8f
MdPCYWv8TckBUoyKO7Q19jFohhxgtQmrHjPEmQ9MnHE4Uju5Xq5qOTJQSIPsoIH+SvOtg0t6691b
O9xtW2GBNvGZC2L7DD3Dd0gZH4RpTJwG6S65ypFceB2nMK8ShHEp+Li8CfysV/LoCkzva+B+V4wr
6RMJhuHx4Xt5Vn91pM/o5aGCbVnMfqUe3mdLgor9lOUeHNLAjOuioQHefygSu+6zq3h0TTcV9Xi/
NOvpDXE+lL0zA/wjPZ150KfkrBFBoPHIEtmvAUraXfRq170lJS5xLwjbOkzln94003pYnhf8Lq/N
L4t2HsJV3tFpOWGifP3mH8pNbfi9cbEqmONNQdle7wCPH0rPJBy4CbNF3+bVcux9MNKbOx2G+ff+
efsTFFp5SXXWxGV2U/lL0o2KHUaeJBG4uCArGXmIk5bAB/yhVj8dLwevWhROaToPIOKmy7YLOvkx
BxJWnLN7BYDOuFFxwBdovjvH+QvHDz3ZeGPWSae1/hXAOYobv5rjyCGr/WGcGMcZsyyM5cPrEAo/
hoOQ7KQcn8f2s/M5vVIPUkdPrHvB+r1tD+WIiwmZCvSJitX2nWQRXIVvMCRMsEBrkHYy32ooO4OA
1sRGYrhe+Crl+z9aoCcAKubQiGE+1Jm06zJr7rujOwIgRgnESKPPQ9i1hi12MSaqY2ydx70e0blI
rvilQKaJ1ODdaMWmRG63RJzvSl8Pc+Lg//mrlc4UjmWgc8JdXzGAbMtILbmgqOwypqf2rtCPep03
pP9TziK43Jj2zg0Qs12GRsludsbO9HQLdpWu1qIkL7tgWZgY6D73WmoKEV05lKEAmia4k6IfolcI
Xwtl9AKA2m0nVWT2GbXTYDw22LutUaN3v+0ftRlHNxdz2V0R4I+e6hJFtqb/g0rvyRcKxealqfLa
a6dW+LmkwOA8btpDlPOZfSsJ8JR3Dipbe9TgU8QWSFdX1JP+BhlMbpjhIsDHUA+4GWPUPkDX6xR9
RSC7+/VjNu3zi8zxmg+KIaL/3gb2pJ8DR/TIaO3VB3V5j2ET6rb89aTb23gGUI7tKaCJkSO187SS
41lYynjn1YtW8S4B3L6kqCwW1DjfW/vIhCX/XsDX76HP20+2E1IEsTa/sudPfwW0duvMhNsPYaES
YtvTMXBwCaZSg44QWoWWQmcV1VNsZqDjUP7BBZjdL7HAma7+wS57zfA+aqSWt7574mLXFg6xoKHe
ia+ccZAk6e9YMyAxiBh3XYPL1ri5672gmKpRlGFUEYmL5mesgwOQhqr9kvrPgI5hS2IcXkxPHMEx
6TFGQzcxOAOKNUyG3yCouNPb6y72y43uuI5/APm08AL0gYYSG3hKw+4DXh2kKc1E4mm9biqxrXZY
Sme2rrPBNpNiEgHa7kgGHi+GgsK4re9+azXMNEi5nuFLKh5Nb4e8yJM7C0eBWNzt/O04DL9WWqfZ
7pYILxJBNS3LwwWofAfYV1XhphKxaPZ31t/MrnOZB0nQbQw9Xlem6xBI6+WY/TX7QJy3tBxivbaj
2RNa+ruz6u84YEcIisixGuDiMBLnyFcGfrSCIKUERHMbvpase3+Oh8eh7LKamZf6QKdvY3hp80aJ
vyVDyWiVuj6ypZs5L/QJjcH4YKYoDJrK3Bs2zYnJCvUYDh5GXOjNse9mzZwIolWqg7O+SruJCXGg
PygJtP3+rCsLwSW4FGz0sEaKoAy369jNFiogzaOpo7ZfVgOkBfBwcxevi8ZX4+sl6tpxEaJqmLyG
iOgh5YtdqFz2c79knMWhW9Uzdb3TvOAmaXdv9hIjJ3Nvah9YoBhmYqAXYlOu0YUs2i5MzQDdxbE6
YgG1XVh55yZqJSTGY6Hxi4rpgeVToU/akNM7tnEVAmznMoZqRtaYeiaqDcqJMI8Hfg9Tn410kJF4
lsRvqj2zjnwQsToq8N4SZr1l9NDesFuK7M9j6kTbcDJy93owq78PHl+hAqWNsHS6bCs1cbuaT1ld
eT+6VT9+W5ogCJdiP6FRyHSIMyWKn+WEnRjM03RtXy1Ljy5ippwOZPmXzvZUIBFDnk1QqvAuvCir
lbGGdRpuJub2gNhkMDbK2nRPHWKYgphgMOMoQsuVDVQ9orBbCSAeZNcDYMCTjr8ZVNAGAtoQxEUi
UBmaecQgKPZH7Rpjy/JLa0LIiSHP7TFEHwk57OXcsZfoQsMjtHqdCLxbV8uFKbzl65lrQu76hpSi
h5iJYOEcBZCr8bZUqYCxPwdl560e5C2CJ78s+ioDYNLWPQWKyu+4UKQ/DF5h7Q2QwCHV0q9E45gb
N9mh3xNfuaPpzL46U2HY9I/8k5IKzbjLGnHnV2TLKdHTY+ueAiutCedMGZPu9hD1TQN6YTcoo/AB
KK2hMsjAG6YYp6mbZC35vgEHrCkmxcxl47Wx86MR+pccLo4I6yHKFB6CkLsIDqRWD0A4x7eyZ566
ZfBivE8IiKfj6TYoZjlXtf634srtBewMYcefduFgH8oCp+Yx1U8k2z2wD2O+LISLRe9y850LCI86
gwtonRbO7kmbBdkDvLa6GK3AKdTU7fCrg8YZu3WuyTpD5xpwJWL9E+AYm2sL0s6QGZFR0bqZ0/vL
Qg37F6X0fEgMxcVlGt+vcVEisUiGOdX+bbIRuwk3QstFkPPoioEAWTHR8jcHUr7yt0XdEZi5zm4V
FY7ETzjBJ99jmWVJmZcrL0PTF3zIQZHJFtY6HVxaaKjMoRhsjfzwSZZVILd9J+t0QSmPTdYtt8on
ykSUvGq+4HymH+E+HZXGRkCA5I0APQXkjuU7e8gmR3QQR0T6lZriBT/I5eDLjN4DpB6xYuSXO2N0
o7zjZ1DxQXSYomwGQXCDDKEGoYiU61Kx+m1DIPo8DAT5IEDwIEPOBk20OYbFr8WjtLL0rMNfs1OW
f1qU2MXdAwlc1p9mAStqjqxtu3qb4WQugL8M41PyIrw/BbA+fWAyynqFoAFOc3n8q/Bw276N5H5J
TpdzDp6SrcSJdfBwIhQbzEuRID2GbZAabH94F5u5BSlVTypzwbICwpOLxnXWvWnxOUMBbkDKjMKj
/SqpZUcL6RCCmcH2uNzVdYR9jYVA89ZWfXkQPSZAgq3vrhPYiDdQizo4dkl0fXgPi4Qc0RCD9mv4
2JOVb1xADYbjIizrmPv23hU2OcXDFzX5Guztd2BAS9JDMOWuel/lol2ZrHzx0PJkVnJDiKRlL1ca
lqY3QWy1nd2humyJyC+5pdQ/pPnQTw2+YAHYM5Jl2V5ecUVrkFgJKCEfdj7lanBqtL+UlqYderWE
Hr7WLnXW6yfpCl2ule5qug0IccH2EuITtzSn2HJ2qR7lVR2Ty9U8cVtGeo+vNq3qzOZwYxbF3v2K
YagcTOF8DlkAAjBrRF7Pyxt0O/2tAJniJXImyfwZhWOCtb1TcLLC7YI/1xzUnDXlbbDOnNL3awgn
ZHJ0kJ//ep+VBGUo1Hm+u5rtwfnWDNzQTta3IrVfAD2mU1EhriE+N1d0TVSvjKiQWCWe1ejvrKkZ
mdfckXRrd97DOYFfCwt2x9YRhsi7ikq0e6apj+tC/niJHCDo+4gJ3x9t3N8MLUnyKf5RfXfAXp11
UeQ30NrtngDQ9R9AU9hoMkkMABu0OMaVtcEBFbSGE6cq1arpDvEKgacEk7pXzmc+KN/TZR+2c8/H
JS2H1GlndGQjPzBFQyy2xZF8L+RL77navsKt8wyiZdQx4GDPTXc/cVmRC2bFnM67Ik2iSJS0q6HG
X+GYquUE+kFg5KmpRBCJnUVEjiEyhgWSO+Ar/ml9jAp6tcmwrpFpBPLBEsKYqOyL3ttXmqPijbOh
oN54586WyO3lydL2wa8t/wB9Jg+4mqAD1ZTD9m9Ex2Ph+NdVfbjkYBWoVKycu6G3sasZrabWMoQY
6gIjequ7MlCqXJqUgrQs7hvj5X0FpIrT0jlhAaLKdla3RCP7tkzPFfeTu2d41aly94LgLeFanLwa
oJwY0EFX9Az5IMwyBGo5o5iY3C14vvgAWRrg2EkcF7274A00+9A0Yv8vBTASmzRSVITzUrYxyb2L
m86MjFSzD1vxPXDuM3/D7R1VuSUTgTDHJ6YzgIenTnmKBipuLc+qAaH3zVFDQF2h2jb9FuZERtYM
+pobgILL8UoZmos04l5d/7QeV/GXU3SG4WZadqaiKI3xufV9aKfalakLbiHilDtUgzLK50uSzZiE
LjfN75gNCMQDdbInzGKhfs0E4x2Kx1jo0dbgG6SKbcII5hD3AuYG3jDmEY3vaDWfS9G7D9g0pYrA
G1vJ+e8y+AulaAqsUpjastr7T0dcAKxMZCXe6r27v/s15XGrlSETPJENn+eNzUPQ11nM8zU2NLL/
557o3PwWoEfS3fHJf4W3G6KKx23ubei/fKrZvA4q5d/gqZwRwl0zTh9EuzkDbPEdpe6Q5Ourpe4x
bXHr05EKtRZsUmkhAdq64hdmnu9iZrWUVNSaFpknS1URB+JP0Tye945sBFYvZ+hmjwGXIzfgY159
c7whFtqv8oSIx+xmeSxc0ypChr4r2zHGf7dGrcfcn3r6uUc4O7/03f4IQQwz+V1VzE4mgdwwCsif
lGaNko6S9VzDprO1C88Ex/grS2FbtpAb99C8XgRGXPgQJwD/Kd4+klOc43eX/IRATZ9QB8ahCZVn
yV7QEdTUJI5p3KQVOvcYvTarfQznu3GIAazzIM9x5MgZ00mvzcf9Upz8q17sTeSFU0nCRF2144IE
qJ13D/ieRyJ4K+orYudbN9nkbqbBiZw27GKU7O8qawyEjFKMDpdLF6BNdgTkMUnVoaKtJdeouHmC
R1ryIpnQgzWZVe+A1jrZOFtfUANUdfc+y2NVy9SN/mzYxgrIDawgQbiHcKS/y4VcDtA/syosr+ZR
p/o956riYsr7j5VDnOFJUb6HeIjPfzQ35tQy60snQF5/XLy4hj6IuwoxTN/d+nOEeblbBCLAh7XV
WYnkEVwK8GvlLKrxbwUxNwYl8w9z1N0e8P0Ta3S9ww1fTmUeL31W18KiAEX2GM8dQXDexn8fZkaj
ubrL1TmiTk7+zrhWcUXV8t2Lwnn11JtiR7lXdl0g+ePddSLbANUoRLCFWFzq8fp+LmPlyUuYqn+/
rWoASC80vKpwgON/r+ra/px1We5eVSrFh0ItAPrZdkQLWwCbdgx7EvnN0qtm04AT644fpomdwE7F
09ZWrX5+Z9vnKYZIgZVKi9dHgC9Uf3JbXUGToM66j998kAHKM9ebKLYQOtvowh6IWg2IPYiRcYZx
8ekNR0la5wi30XRmtGypxQRtOihRCL98Q1IIntbvJxbYqciQtgoHXbazoUOk4zI2hKY5jGOFO78j
ujRwROBAWSHgunFzRhXbHQpo05+Y9marV4sepPcl7LAavIBfG6geJ1qg/ug9wVIgLKr++N+TGh+Y
3S/SI8U2X3VnUyFTookKMDoNSoDkRBwIUn7qxpSa6QGjIn7hsjRWREKRhy22ZYzFDlI9iOfnFcAY
Xfi/dH7Gg2GZzbEslad1EU+Z+oaYrXjk18LgBTMhmk9mZmdRVVc81AnRUas5KHsEWSUA90Tp+ozi
1OZEdyB4V/UPNAUaWlRck0Fy1egKpysQ2DnJPiXvRp1k/5hMV+Mw/0hfh7PZ+dBPeZpIhOUgTWml
RCHc+BQkp2BqqYBBLV6q763oqWnnfddz8pA3K7WNn6UXH7yT+aqqSwFgAhMDVJt3Vk2D1klHOB65
xmczhL8EKRBD+4VodOhbVMZ8EWQAaXIfLDv1KyCnBhYZpv445ZkoK1fDVD0jC+dxvIxr9w0RKP91
xoKOsG8aCOPjZjGkIIrUVo8CUPTa0ie7hHCrNLGf35MU+r/P6q5a46r0/DGC5SoEv3Ix16pbT+zr
um3dWGDfBpvSCQLM+CjbCSzIJP6rHLYY3qULiMohHsQPWiXSeSzKcvfRXg64lZbn6h5XnmPGuSSa
FENNe4p5iB672M2E5J7+82TA78Z0DqrFjmFOxpnE+AwQVlDGzeocTB3WC606DYNZNeEwr3K5E8bj
9TE/5MWi4vmDh9cnO73/VT3DiH/Ifx+G2cFR+i/+WIEPuRJ9ZyoBqDXRHbgOsr0bos1h33Pkc65B
9NdPWWILnrmaLvtdrxDuRcT6VxRlO/ptWGJKeUjatA3lTYXqMQFFQsUIFvPbgrKv+Sk3Y6x5F/NN
Sjckc9te5uUNUlNO8VdJFoGi45suRJ1bUnl7462cAYY+/zIpEegeMtu8/7vMrePwF+RC058sEST9
XlUHMgJOXO49hS6KTKXpGzBEa/ydfBPvHPp+7tpskZ2fKN4voM0icESsbggJtWkEPPwD4fTslBOb
02uZcLTkRQO4pwvOzRxTos9M15CAGy5fLMgRI83EgLQDeNl2A8aetRK1FdBhAraLCWd3bXz1zwOs
aZIIZQ4iH9WpneRzfx4CEtoSqWOhAzvqjxPUxObATUmQkW2jhd01VBolg22EGEkaF52zLyQWbIP1
SGlU02dAGxwQrHjSOWV+gb+43xMjUwxP6SaaZoVtpd5euO+ElxrAFZx1faZHv48h1ojlcF3UFVlK
Ly+HKcfRrsuHns9r79HkHdwUTPFHpDr0XzxTAwHgKhGTXtUN01PNCVwy4Kq10/gApWQz/8SaoYnh
a+wgK7Sq3K6QNrbXoOQN0q6LxMvRiAiGjlThDvStykb6TO18KIrFU8VeFcfU6JFhiNWFHr09LYCE
C3DOXOUNWPlCunGi7gPl1xWHdfeJ8OZbhkpU6TTpJPSodPoHgFGk0cJN6A37LfNfLakrMV99RbBB
dNL5Opei9mSg8RqZKg9WfRaCivRb2sAhtFM7Pvx/jAZ2qqiPP86hIseKjcM8NuKXpVFivD+omRVq
+X4bwvVlqfryA8Xoui323QQzbDp7gVh4g53YjfVYrjstJOQBTTrSljTMJyADFWd4rsngmhjeq206
BWKWnEvvFdMIJBLNeXXo2es1klGJD+B71bpVt1pgXb/L17zpmt6SZlCZ9mIJaVZ9TuKztvp24Amh
tG6BWYNQMhLCgNHWwPa13Dh/Glks09eXuJH+VlfCoJa8GHos6L4WL9mpmEVViGEh29a/zRLQEhnV
5iP3rOrQ4bzzvUUthGoAsIcFQsn9XuvepeAtzsszen4pv49zA29W4+6jgRh+07gR8yvlDo9zYhnJ
aGhfE8IYOrnscf8HiKdNtx0fSIF0edOY/i59h7f6srRpK6PCo5ELOgV0judl3I3+phGgue88wf27
MsTm2+X7neXbaE63QnqGqepYrtMobMEJUbLyTbTMjyOBeqBiRLGMepzFVRQ3xH1Emk4sjSKGTDmt
r7T4F6Ce2Ud8npkwpRRi9iEVG6MtPZ7yUt+ujPJocdM/Ol0jJw1e0xfl91pVVxGVBS5rYv/aRefW
uM/KLoOGprsfkstePK+vLnohq9qVI6HheUTWRxSgYH+x89d6OYaXvDn12KygUn3d4TVPIXZiFR1e
wBJzmMTjHEkAWy4qMuB3a9uQ2GiTI7TVzDUhDmKzYiufUA6mAWbJvNxx2JqJiDM2JlyZiGeY/INH
gZXQIr1Ky8WdB2RD8TZHGSp4KWgAu5yoqjAn1CaAizk08g+bf+9AlsRavbzGkxwpZeQARdSnqmJK
3SPUnPLwEIdiaxlPkB4URlrPQc0X7YpJMNXbDSOv1MVhdVDWo+yexAA4fvplsS6K2YGvMjkyYON4
sPOzl74IF7gbkI2n7VPJWRls4cqPxy9wp5Z45+05K+7BzwELP/w2gM+oAWuipxTEOXktjjgzqTE2
fxHAkQfdqWLWtkn8KcRaWRxPAzeMvBMllUM4kjl2qFp/9Tc6X31eFiRt8D9+9ma+jReDK+OpV/98
IKaCL7SMGKrIJ/9LOmWKQkox7TaY6LohmGOx3rBOYGuVvI7j5Ty6I5oH3p2nN2eRI+X95DgUWOJq
gnhySuhAQIteYA4ehppcYCbtJxTkjsT81AoIzWD4YrU49MuTZIG8uVgoZV7Hki0W4FsOQdY46qcF
3iECq5rffEJRfyVX3Bd3UfxS7lBSMV/kRBEPu1CcBfnO+CbE1S/9wBy51mGIbYEewv9Ngi+TLo/F
K9Qqjk4oTzKEpUQhQDRCQyplEhIPruM8bJcKD/Bjw0fE0pNVvIW6MhVSKnMDp/Gj99U0r42Q9eYE
+6xDJExMnnFT+bv3YJ/Xj3RaAYuEMlSf8i55aSlOhTQirHAIUvZdZfu+1ulQE/4c2kyZCVhsBUQj
mmg+DU/WvfodnjZtQUoB5s3IwemQ6JcYfLrqemtckpnnXxCXN/z6QL9Jip9CZlAOiarFQeXqduxm
vxOUkLCw3WOYw8f5cFp0IivywCKUfzw5S4smWrycCMDhlXZORkoiyX2SaghIphDTkiMReSTm7tUj
kQNF12cofs7Ss2uSSloNeyeHK00ve/Hru9Baun/Bo624yn3B3I5TqjJBAIz8MLnj1FssNf/o9Ljr
5URSV1zL4x+MX4UihfUBHqyuVhVG9PDW3kxXHEdM1HkKSHb+dYyLrdz38InRBxdslLuQjjrTSLAp
0h3C4JYHBSmtmghCikvtkIj3anR55SHUUzRaHmiFAVBkR+gk8lSlHlCNnBHfdaRHY76hEYqagsgm
SG2E7cJ5mKFTRDL7VEbKIG1Tvwc5Q2Uuk2zOxCRbFptrYAblB726nNnseVQFNX7xe7D+7Jszx2AQ
HASBI+OwNiKpJg9Uk40WSLbzWdQh7jJrVPHjumKq1UiIZm/t+KjviCz7d1NFSS9zzW0lo4NpFWax
qTFaMhSmNWJbWdJMcbEqE2HSqRrH3rjZOhr/N33pDRTZPPlTw/bB+dunipoL5fkjLNoGpX2MvJDM
ZqJ38w8tQpwovV+QtmRJrY04xcReBO3GZIryUvEEDUSe1EQvByJkI7ZjuhU1/0vtgZ1xCxtVs8jB
ejIiN+vK2RHjXo+vuAnYZdc99CaVd0dJOKY3qgJiwwe+5aEr9W6vksLRYQotYxI+jli+plovSc+p
YKnD925u3bLyxbX8gwNHQi00Nzn+CBw0V+zQzeKZbbvHgg4UIOQS0UP+nBV4BpCbZ/l0GmrodF6p
vyhLJcZhl+4A9wwBddQW/YDiJpVGVO4St7ac1dP2fB4xRiZMGeo8USw8sQ67nV9xmA0JB4FtLt5O
H+Ml/YsxAeKXTG/GmMVgueQiDrTNkEnCFNkVasVYYB/HqD2/PGZzbK0Lfqj+iFK9h5XA87rczLWw
ai6xy1D+KFG9Kt1NzxRGvfgQfgyHuFnKDnQd+KlfOpwp3oKgXWxpXzlhl+RvMpzwPkWux0qgCnOz
XuyzcjhQb3/Bbt61Mzsh2ipruVEj3Tg5LDwK5SZOMZTtm8OVBxZw4cEaDvVX1tXpeaRhNgnwu1Ql
F/XJvtz8ymip9SpWbMXfJFm3YLhVcuKheYK0iXqzNJnewYinRpOK2SQeVQlQqd6ddi9oa6hQsyh2
hjl2QaYjBi5MZ4r5+BQlsZ/dy6h70uF6o/VenBFCsUhMUCyZ6opWHUcV+24y3+zd2yXMbCt6r2Um
vOj4r7a5011pP6lzgkVORyQwpM9OEC/fMOYa3b2IwKMdM43ibPvj7uzRAdK71MpCJi6aRcwNdTSL
us7jQLlwB5ALm4btNuTNlUVGU9xaYK5Dcbh9lV3XfVtH5qZCB6lNmsWxEIExv+JzuazDcZxqtrM+
QSl1ghM1eMdHv7k0x3zCq3aFb6zlmI7xk8Su7vsUfFs9Cn2O8jFfZPTizci+ZYAMzGJEzKw4nJK3
ou1Mzit0H7eFPeR3NvINfMg6i7UCkL/UXhLJY2/hI3v+f5Ayx2ZxkdbEqYDf/8p1rbbja48CVfOC
vNpDfguBvntU7OMP4YA5ri13hHDlmyBkwow9qioVCs3c4bjTYRpdX+rEXfpKZJFPSFA7531fsYbX
3i6+jJkfTCMTBvsA7kP+7jMMPZpLFTzRmRzTQwLGERAljvcBQ8cIDwY1N+eN4cM+pk8agMuSXUa9
SO29rSpJdMLbm9OWleNLUZHbY0lnoszVcMqxiEETRmQd82sjENqAVImeh1psMHfAKLx11uRHXfwL
emKUT2NCrBPPZCTRZhyqWPb542GDUs8J9JgkmDijAUFzpqujn+QwARw6VZUZ76owXkEP0uiV2rTM
/Vi/RPVeWsybbyFgcsVYBMBYBg14DLwyAiNX2cxQ6XF0aWYtXDfHp30z3FYkRQGzN+6I0HHkzv5s
uOI5l0Egwl/JX9FbvBh1qCmh28Bm+pIql9XPc1dZ3aRMDFReq+HlOFv3ibYIA/lif4U4iEdM+xWt
CKzAkRwnhwOnx6v60UA5w3pg0OUN70B0nVVaHEQEqU/LnAsdlNfV+cqPMgToJg+r1FWfww83Op/+
er3k+ACkdnrXoBQSCKsgFTvUJztUil97CT8dYn1+9BPT0/bnJ9hvRgslEkfFEBkMceLOI6MK8oqn
7sDeNNyP0leuJVQkjgQ1vFaUM2rMnKTP77C+DsPFsEbMTUctxd4Lk+Qhqv+8JdXbyc3Vsi0DXrtB
qIyI5V0pm6S755oc27xbCPRF1m60aCqoIuiRLtMl76zAh2Z2cY0xUnR1wP794McFd48+C1M4S6Z1
X+xUaBMm2jT2zzpBjAcz5q7k+CK0iI5v9FZDCV3WnLk7UrQrg2FFGoADb7gaHXlvnbSgXNN28v/g
d9zoeuoB9hLTTbtZ9yacnZT1LebB4ThJJqcSCYWUKIuX7cCD5wDoL0JSeybh3tYFbfcY+abPJppT
qkTI2M0j4O236eSRK8azcXK2Lv8f4ZOrimjhP0SYKVv4rBMScc+F7wZi2+l3QkGf1fq//fEdiScj
4ItsuG88Hp/NktyMaKa7mrCLwLZylkwGnl0Nt9lwr7Hxrdqr/X7HkOpOjgDRjggQa4RVhNG1mLbQ
42I3QbLIY4cISDX58saKOdgHftLi379EGF0xUkD8RHXXAn6NK6PJtDjEv1AP5vXCEs9SBbLIC5HD
u14MCoOpdy5UI0dsqkylS+WbrrZovPHZsObsUg2cNKxRxo9Z6+9WLYqPc698hsMTY6tb6F/dsfo1
VHyxZGu+rMwGl+1jKF9yAnrHNjpzu/9wJAtLXe0sFEQ2GsZzaSOpzLdsFJmfIqPZPyW5aW/B+GZ+
kqnZ8+eckTsr8U2tpsuW1rOyRtGyXZazY1K57YNoXlRe4OxEi0LuwcMbs0LLBBtQNThFMLdqEsXr
pVq+q1kVIZi4dSSOAG5mV3X10qCpzgEx2kmDLpcYyCQWqy2mL7HQZ4Q4IGY58We3jiBglnycqUSv
W5vZkjTdWgiM4lR+Fx1lXmPF6P6nJqgbDYU9wScBfRYRJIZBSVzRh8m3RcpL8PV2fCNG6kjQggdw
DkFT0Zicayb1/Y4+1lVtiyCzBA5EL1wwrTX+XOttBiSUI5Tpwh1D2wyMdN++tQsAhRASjlPGk7Oz
sVj+o2sKV3uIUrf6sYbWgqCDPBYFXDJFrHMCPehfD6fPUvWuIofSEpisgJkEae+8kKqEHnC6shsW
lumXPIV66iMkh82yyBcpWHZiKlMVJnGnd7lElAy4J4B4Xv+XrgN+Qatr9AxlSAAtyilaPh4j1cGv
67VQU6WQDi9q+lE9iM63oTMexf6BlOynSITvzNqw5DeklRnkDiwO5SzRY8AiLLkMZRYy/DZnJ+uk
GWOTGSI+GWrcf1DTCW0fCo1jQpJ4yr9G2P+d/1rOMGeY1z/O9dkZsnIGUaVe9s8eV0whUjy5BiHh
1yq/wff0Q5wT3w3R0z6cNwvH5WXtZ9x8bLYoJw2M0cnYhVSwEMw7krOGJc0W2sDSbRiHHaCyIRVL
vQfp6wqI1T2ssWUeCBKQgtjoGJMvpo79lb4HuNijPWY+/j4djriSA03Z7HRpYyTvQIaXkh0DUqKh
pQOX6qR08j2kczk8t4ZGSs3RknCGBy4GR4raknsuwmcXcdIMr1j+tMlxDFoOIokMAzgxh4qTUgwp
TMdMomaaJOFhEUjRGI3LCgxubbrHe2TeVRFchj6m4pRxhVV82UJXzcvvnvsLFGIRzWhmzGGTxs64
xNsn6g0rTmvJBrjs8Gj+hAkjN+V7Ro8hqfzQcGogqsLLgyQzQdtmdLr6o3t9Og57VumlYT4FKgrm
FRZJrlExCu3jcCbGDKT0X+nt/JohgJAX6qUet/eRgxcVdJAkrXjC1X+XTe2riOZlDCSiMBJNSjgX
ScWaYmGyqrOPPYjiHU4dfZrcRSiN0cbH+ypTEEs8QeiGlE4NTkObBBXm2bLbBocUkl97x9Sor2hO
l7/4S3WmIS4VZ1EXJxeWARAAHHe9bg6x5ZuRV6vvQLhqgPdg8OQUUA9evwocoHZj/uAwxim22YPB
a+YEP4+2ZeUzEsT7RKW/NocbNGBicNWsLk4tYIN4cDGJk3VC7ZzceMcMQtAKg+yqeUU5EAV8kQsc
LaOVNHj/dDLtJ3OUXkL6Kd0gS43Tj0JroZ3V25F/LsTzP/7Ri/s6t8BoWM5D3I2a4zFy7nL8GaF2
FktMy2h2QlwUAUs87KvFnvlcHT5Ex/xoKZGmn1PMIkoAIk26wXVxP2Ecrh+C+dp5BX0/8rUlHjNS
67Tty9BMtgru75mYC9jBunpegMZs1newXPC3l8p78hKc2HQEzkBamTCaUPLuvKPlXpbrxzaez0oN
3JH9g75t4fIc4U9t6L5uIWj3ldljbUYPDXii+FjEN1e+lzJdfm2frIrWlVvfUqHQU0xNtHoW7lHT
SNWzMWquTnscqGQ3sC5yuB/YdhkANumk8/Bc/dreGE3VAfnbzDWDIWKl4+nVxmCbpvrWDLSquywv
L2FnPP71ds5K19RlImGIvqZxAW3VPu8sySHepqesRp2wjZ3cllGFWGhbUqT9ZLMQpxI4OVL+2UIn
8sh5V3A0+O8uJj07emWeiAbInPXjC+gaHR9N5CE1zitUtC6mo4Hdxu16F6OiOENnYoKeJtpITWMr
RlQFgDVbstlWgbhH2L6E/9K2l8Utzm03VZUJujI+aSpkLl7hjWz0HI+uXmq4Vj9NU96uPp/NPJx4
SleprmL/l6H3xL/P6pdysU9A3rHYZiC7xEjp0AWzz/Z/7HbHzTir2Oh4dXtfGWASqQ1HQp/gn+x5
epgEM/FPwQ0B3IVxV4VaQD1WrHG0vxbiJVBaA+rId3XmqGySNhC3Jgzj9HFziLPgDKyyOWO3k177
UYA5ljb/4L/sSt1+zeCDcCJj/vJ4I6sn0Hxvu4lQRFXQACwCPzHsQJg8+/4zhE+DOl3hlO8U2gC9
vW6BEoeZIxM/rovyhBKI8A1FALFaSPZQ+p0TPDuPZ2fjOME8MFjqmosyqrjE0kPLQaqytSQQa+yY
DsWf/FtDEWjIA/g+v4UciXUmChPTLKqXCYUnDDShvqkesTEGIieLaIGVTIqgld3E5mByIAuHzZ4x
r/6t/Qwjr9L83QeKFd3jGiAQd5ZowNbWh7ogY2xa3/yo70fwYBypcyt2QCG8Qpl1vwo48kLfYz+L
CbCxOjFz4wb+LAdHAbdXanVko/9C//iitr3gP1jk2BasxidMkUyAuq01yh5RNN4j+Qxanhdz1mWk
V5+doL83j5wt1Q44mlLOUsUk74hMwcFYdRWZ+pFvqT/xtPnb8gFBMcJkCadnKf+dzF3vqUUoUOnm
tNIHdrp6ONZ1RuGyjdjxE9MhS/GQ5ussRit02sTVejqm/pAT7C8Bn0C5yMzn16VsDk/obe+Am2rz
BxO4DB39/r8Zj1IkIKnnted8UmdFVxHZXFh+BEVwTuC7PUdHZIb41HebtDdNFW8/Usi31Lfja1FD
B1oE8ZAhpZN9W8rUhdNaCuIKylNgjSeNe2ZhNntW1FzSWqpUKS4gpbcoOeQ1YoY8IxsHKXDRqrx4
839fehe+HTT37qTyXudnmzPKWc3bocSajaMSIEotkNn1OzbC/EUIyK4Bpmn9tFTiJrPbTQglgyBk
06+3JmPnIwlNDj1CuamA22H3SeDd1VfoGCPD2Vgph2iODNmCaKyFzzviq/B+fhpNi8WxTSCEhDfF
k24Q2AqYN9NdjtKPTQ5nnAMnBrlzIbI3VfmK2rFQQYmAuDkONv0WXgCKdt2FhvQjLOLhus8izWIZ
MN3FX0Ts8EOPc94o46MzMKkrEND+a09kutjagFD3g+VHblFEZT1MHEHLw1kGwqq5tKCkfyKe6ukT
nZvsb/ZgvimuewwcnVZs82a7OTR/li97Tk8qm6+eaCCaaGEKQOvIrOnJer279d4XsQDLpcdhey7u
w049zRUQBDM0GPFi1f5OrntEreFEnpZ2Bb6f8KbQd8cobm3nZmzZjC2d4M/IR8tn+jYxSI8/fJNe
p3as/Sv+f8OufhTx3F3XpPk4FXSueK5BJHe5+QQg1WuC3M31919F+LKdMSDGJ8pmqEm0o9QkxHEs
XjGMIcfngfkIy7wdxtagd5erI7h6+7bLOByKpUlrb5A/J3ZbZlVfkABImOSHdogc7unFsh1tuTEV
o8BsqQFmutBDe0wWOJKp70z3VOP6wrbXSDvmViKXphys9//YC8v811g04KMOFihiJTAuswhfojJ7
JYYMRz4vF81YedO/0xltMUGnM7hukVvyegUsskelXIzZNvLJbIo9lB4yKXmc95BWweJ1usOjHQUh
YoPDJsAEOJhzL44tBDOIcRJTuAl2c/lQqJxAviDUGuVsqWSRSM7VTZioyyGRi7qEcyJSj0eL+yTr
ACi9AfmdBPAtMO83wWZNQJRvyc2TmRXiV0oR7FnURTR/xa8k7ITMFcJ+SZbspB+gKIFg2wdK5o4V
sPK2B3EAHy76fTmk4o8ZQNl8HyGhJBP/e70hCLUpHYaGnh3oANfh+/glukKRTINUcBTNurBoljFe
34k4VMCMf40CEdNIigWGtoEyxQczifLMMnSDco/I4D5Jb+fnhIZtRCpS1+Q9AP6vendSr80QT7nx
XuvwF2fVSXQlK3n5AiXNDBJ3urRfgUPuSHrN+A5ypY2muAN2lj/f7cS079lnR3aE/8yNqiNSg7DW
ICWV7RaS9HxkIDF5jJxgTHar8D9T6kDBMDgKy7ym0BLYVABp2qh5fTQLtlFf9EruHqUPGGyAjOBN
8HAKJ7RK5dnEuizYgI/KhiaD8Rr3YW8j+P/wLLUETroo8hvHMRtght0ZgUhLjTFiNbhRTxErkRUy
voIbvW+XL9ncIPfGD/bw+/rFYiCsvaYRfjsVG/1Sm/xy8nJHg0d1RiDF6qNP15XW+19eUwt5jqII
/Lk72fEXmJJPW/wKiy7sGjweBA5VU9NR5CRKkoF4vt4ajkc6pFr1Yx6wSegEiGKn9No1DFAG89XG
u+RpT3TSXjyEaSWQj5KZHfyrfsnuBGVuoYfX9MtVflkDa9CHLcClJP7rLt/8aZosuSt+cWDFJm7O
ZeRvGwMnZry1IZ68Ofz1HlfhCZfxdOGfSiox/wXrwUcFlB6ZmmbJa7s1+cqfTtIFOnfKf4WVHBHY
cimJuOWFD7x6kIuY7aDaMax+0DLvaWuwvyO6h0AlryeMVYj1+5iwN+x8dosu/DqtiXdLAi0LRI5z
gR/R23BgTeqpgdxxL2+kgqIEV3CKyRMR7sXAPizglMTJgRcKBz2ZI/hvsnR6gGDSRZCZqERnAp0w
nnclebHH0QR247dHG5JMl8Rx2oOqbh+B9ANud+5ge+GTl9j1AP7nnb4QQGI+8n1RWxbVzVfL83EK
Jq+RnPOgygdZE+ZfbZ6vRCT2XOUsO+iTHEhGVjBSmq2gV0vJ1OZsifdFO0/jIhU0AMv+Y7AG8C04
+NdKVMIS/0k11d3VDFg35D0Dbm1TS6Q+p9hJ8XfpRSgteFIUuv54jlpRv195hkFK+XqP2khmxMl3
xUPm/piDBA9GV4Ibu5NfEXFSc38A7X1nx2YvA9595A+mWii01uowlXRsuMkz4QRFJEfs1Kls/BYl
KrNlCWUFuJ0JTsJwBixnMCfvVu0NEnWh1qedqzdzeKI6Pwx9iUAMMyGCCBlzLv6ey1hYHGfwjcV8
LynCFpK58EBWS2aW2xZBJZXe0MZrZFXiLCrW8hAiK58N1CYSS7HMkmk7rspVZt9E5Z/NqULd0B81
K1ySidUoQVZ+45hdtidVOqOZoAZHNJW9FiVpP4n0nqmzhTLnu8OHtLNpX9Mp6MhuAqXPlAoQrBJC
RDLtmHcdUQ8TbeUBoMkkAQ3vzS6rZAt12uMZOq5N2GEzQ/bOsbuEXcspHnXb7koDJGAFI1dsGV/g
o+qIV3Rwc1vou5OKuPyOUZQdzXxdslg39/wRjD425H2tGIp5+6oHC48esJkBovktdABTiSZYyUxj
E8uRbNvQjR9v+O3au+PsjtnSmnekBZnDzWz+QbH00KM4ilghOlbuMHHqQkrdn5AxV2uOh4RXLR96
krQKxRfVlLYum0y6DojS198jg3A7M1itvqUn5szbdPbvfHOiI3tiYZ3v9EgUlB8liFJlsCqMg7Rg
XrXQMp1cvOWTaPzeJFoiHralDTFJulGhS7/48dl1jue6KPViNXO32RYwr9bctRn0yWp6z8IH9jZA
kZYwA09x4Ddf7hpDSisKbllT7O553A5+KT89RAs7XhV0nyfmKLuT79CPGnwyO/rAYz3kS8WjdlKq
0YbiaOVCoyL4chjSjbt5TwULiO5ADS4xXyDw5mWkoQYF2fwQd4tb4AqF1TMsGZxAkoBBiNNPlUXh
xAzDNazJeofn1Jis9/DlA9zXG2wSv+1uKKS8gSx6Yk1aT8wfJnURXxHwA8YVbir3/W7tnNRk7xht
f81b14BFZKwM9mkWlNPei30BpvFtHCcmhvI17ei1ru1SO9/R+TbvYG8r9itE9+tbuXgIMVz1gl7e
YDjo327+fiw4z25IGXMivsqNV/RogN9QWBegUU1ryjdx5KgoKqsJmgVt13I0LQjY2Szcx5xfuD6z
HI06famgu/sYT/5NtvqwTgUAqvdjeWyU9M5MmeTIK92eEtpMdc4VgmtWpkKhvYfPM1PtoVd5/y8k
vNnEdOmNkMlPrDplHGG4c+b5z0f72r9Zre7qav193flPmQ4bXJxzDWHZ1tbuNyGa0N5WPjkGUZsy
mx/+WB2MhE1rrfUKn7SOtu2QcMdf24gsBG5x4hblFSxFcqTSMgPFmnOuOXuJHYDfj8n7HFgD4+XP
Ky4B1oBCjr5wpel1H39SpBEcwHVB5nJ2ApQeQoljFjGs7e29EAdh5+UpK+RQqh+ru0EtS2JsPc7q
99ovjUQAagdy7rZVJmu4pg655fNS6Gk7x5cW6x803gIrOhoQstdNrrsxPEAF/PW+KLGkXU401NiL
1P5JF0PqVPEs16NH9TfsLDbo9omxdzrJnTigpKpb6/YKYmisVZamT1sRtZCWqn5UsGzHYkwdPqJh
CfzGxKMKsa/OJfQESJj2Y5BuoWT7e/jIKkOS9C4ayD5QsuliVEVYj9cqtI6AJWWo8pxIxnqLIixk
E226azMIqJWnejm91gum0Tnd1Tvi4j8OtKr2dZqVn1Jmvz12A1/1qzQH6xyrqxTQRtu+L/TwmIY6
76ICiyxCdWyLm7lFYmYjcJyvsfmp3WHbDTFNs7Cc7NCBavu77G05xfE1TUJooui426dP0ng6XOuQ
693O2NFhL5ggau4CyTq4KUftuP6mnEuuKeH9Cw7FUhm1omWlLzFAWYLrRqG0BeLd4EfediqTgE2T
OFkI+m4Ag6ysN4HqYwcVxezUlaGdcSp4BPoKAdbhElsi9W205Q7PdXx1TndHVqltkzNURuAove2D
TOuTUnpgxQ8UhYNcbVAJFGg5pHbCr0cQUtI1TSSVUvBZk/QkcIuMo6d3SRb6Apvb/j4ZI2Ox9Net
Jk8yZgZQLmjmKBp+JfKGq8OjHxGgC2GyffvLRcozJreMGJjGfSVitJyBe8if3eTDoeZfKnjDibMy
U1jV6YxTspWuRJLC/tFq/wy1UFCY8sDgxfKY9zv7GwAjY5XEMFJC7A4+B9zFKpZZ+dK1TlnbQ5PR
SqwlczrKPumIYyC0sI3opjrzudv//MTh2NhikW2Z8195J8e3pCEwzFmjdkRbwABQTW56kVTTmgaE
djmk5GI0uDfSkFsb1baZtMBtdCuiTT0SylSKlnTVZqIOZAr8d9he38svyhNZ144lkKcARdP9h9Jg
0MbCS6Yp3bpPFm5wTJJuamBa6aLglGOxBUq3m6y+oHrnc0aKskfRG2oqz9dAaeWbnjhq48GxRZV4
U2QECh0AXknf6SSeJA9tSpHhd9Dot8ic6RvKAi0vaj9ohahBL68erI9DSCGG4JJTjFE94/xy7HOJ
rC4RIjX7r7+LPqZocuuFzUoBaL3MEodyaXm4SzA9eYnUqEHNv9BbaB9uwsrOidbUqiAzC6E+vyEy
Ex2E0wEJxnUNVFjxobLJsyByohlcjY8W89RKoweFrQzIs505+AbMS2nvKfJU1ml+EUQZVkZe3UoK
aPrcN5Voi+KdZV21Hs0Hwmi7/6KSO79NTwvtpzXNlJjY7H05/7RHbUp5Ro+7prn2MBD9qOZTbD+T
ZKpW/72uL4B5FttIO/ECSPROLRKEpLcDECsT9pJtqZxyJjDXQglOgybIn6Ano4Jr2oEnDDkLQB/1
yLA8y70jJcTcL+ldiTlldgQK5rQwRgpp45e9WQe72dwc93PgPQ2UQSMhr43zzzov6VzORiYJLENf
ndnyzZZKpZKKuTZ5HIGE6gEDAGkkkh1o0h9XAVlaeb4Cus6FK3EXW0E/newBp1bW8fATe9V9Tkii
q9xX3eQZl8L1I8tIoBPioQd9bJhG1bmgmZtZZlTxMqls3KAviWc6uvAv+nyevQ6YcblGapUn6aMS
nm6xmxcRirgh+MUO0Qjl3reMGwjgOESBPhInTr5ob5Zb+ellmWXM6J3NsWT9YEPHincCfGAUzybp
M620kvPmf+JxasxDv05v7HrEYskv6pA5CaqmV4VXw1dx
`pragma protect end_protected
