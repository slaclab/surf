-------------------------------------------------------------------------------
-- File       : Code7b8bPkg.vhd
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2013-05-02
-- Last update: 2017-04-25
-------------------------------------------------------------------------------
-- Description: 7B8B Package File
-------------------------------------------------------------------------------
-- This file is part of 'SLAC Firmware Standard Library'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'SLAC Firmware Standard Library', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

use work.StdRtlPkg.all;

package Code7b8bPkg is

   --Exp
   constant CODE_8B_C : slv8Array(0 to 127) := (
      "01011000",                       -- 0
      "00011001",                       -- 1
      "00011010",                       -- 2
      "00100011",                       -- 3
      "01100100",                       -- 4
      "10000101",                       -- 5
      "10000110",                       -- 6
      "10000111",                       -- 7
      "01101000",                       -- 8
      "10001001",                       -- 9
      "01001010",                       -- 10
      "10001011",                       -- 11
      "01001100",                       -- 12
      "10001101",                       -- 13
      "10001110",                       -- 14
      "11000111",                       -- 15
      "00010011",                       -- 16
      "10010001",                       -- 17
      "10010010",                       -- 18
      "10010011",                       -- 19
      "10010100",                       -- 20
      "10010101",                       -- 21
      "10010110",                       -- 22
      "00010111",                       -- 23
      "10011000",                       -- 24
      "10011001",                       -- 25
      "10011010",                       -- 26
      "00011011",                       -- 27
      "10011100",                       -- 28
      "00011101",                       -- 29
      "00011110",                       -- 30
      "00011100",                       -- 31
      "00100101",                       -- 32
      "10100001",                       -- 33
      "00100110",                       -- 34
      "10100011",                       -- 35
      "10100100",                       -- 36
      "10100101",                       -- 37
      "10100110",                       -- 38
      "00100111",                       -- 39
      "00101001",                       -- 40
      "10101001",                       -- 41
      "10101010",                       -- 42
      "00101011",                       -- 43
      "10101100",                       -- 44
      "00101101",                       -- 45
      "00101110",                       -- 46
      "00101010",                       -- 47
      "00110010",                       -- 48
      "10110001",                       -- 49
      "10110010",                       -- 50
      "00110011",                       -- 51
      "10110100",                       -- 52
      "00110101",                       -- 53
      "00110110",                       -- 54
      "00110111",                       -- 55
      "10111000",                       -- 56
      "00111001",                       -- 57
      "00111010",                       -- 58
      "00111011",                       -- 59
      "00111100",                       -- 60
      "10111101",                       -- 61
      "00110100",                       -- 62
      "10111011",                       -- 63
      "01010100",                       -- 64
      "11000001",                       -- 65
      "11000010",                       -- 66
      "11000011",                       -- 67
      "01000001",                       -- 68
      "11000101",                       -- 69
      "11000110",                       -- 70
      "01000111",                       -- 71
      "01001001",                       -- 72
      "11001001",                       -- 73
      "11001010",                       -- 74
      "01001011",                       -- 75
      "11001100",                       -- 76
      "01001101",                       -- 77
      "01001110",                       -- 78
      "01000101",                       -- 79
      "01000011",                       -- 80
      "11010001",                       -- 81
      "11010010",                       -- 82
      "01010011",                       -- 83
      "11010100",                       -- 84
      "01010101",                       -- 85
      "01010110",                       -- 86
      "01010111",                       -- 87
      "11011000",                       -- 88
      "01011001",                       -- 89
      "01011010",                       -- 90
      "11010011",                       -- 91
      "01011100",                       -- 92
      "01011101",                       -- 93
      "11001110",                       -- 94
      "11011110",                       -- 95
      "01100010",                       -- 96
      "11100001",                       -- 97
      "11100010",                       -- 98
      "01100011",                       -- 99
      "11100100",                       -- 100
      "01100101",                       -- 101
      "01100110",                       -- 102
      "11100111",                       -- 103
      "11101000",                       -- 104
      "01101001",                       -- 105
      "01101010",                       -- 106
      "11101011",                       -- 107
      "01101100",                       -- 108
      "11101001",                       -- 109
      "11101010",                       -- 110
      "11101101",                       -- 111
      "00100100",                       -- 112
      "01110001",                       -- 113
      "01110010",                       -- 114
      "01010001",                       -- 115
      "01110100",                       -- 116
      "01110101",                       -- 117
      "01010010",                       -- 118
      "01110111",                       -- 119
      "01111000",                       -- 120
      "01100001",                       -- 121
      "01111011",                       -- 122
      "01110011",                       -- 123
      "01111100",                       -- 124
      "01111101",                       -- 125
      "01111110",                       -- 126
      "11101110");                      -- 127

--    constant CODE_8B_C : Slv8Array(0 to 127) := (
--       "00011010", "11110001", "10101110", "00100011", "00001101", "00010101",
--       "00100110", "10000111", "00010011", "00100101", "00101001", "10001011",
--       "00101100", "10001101", "10001110", "00001111", "00101010", "00110001",
--       "00110010", "10010011", "00110100", "10010101", "10010110", "00010111",
--       "01000101", "10011001", "10011010", "10011011", "10011100", "00011101",
--       "00011110", "00011001", "01000111", "01100001", "01001001", "10100011",
--       "01001010", "10100101", "10100110", "00100111", "01011000", "10101001",
--       "10101010", "10101011", "10101100", "10101101", "00101110", "00101111",
--       "01001100", "10110001", "10110010", "00110011", "10110100", "00110101",
--       "00110110", "00110111", "10111000", "00111001", "00111010", "00111011",
--       "00111100", "00111101", "00111110", "00011011", "01000100", "00011100",
--       "01100010", "11000011", "00100100", "11000101", "11000110", "11000111",
--       "01101000", "11001001", "11001010", "01001011", "11001100", "01001101",
--       "01001110", "01001111", "01110000", "11010001", "11010010", "01010011",
--       "11010100", "01010101", "01010110", "01010111", "11011000", "01011001",
--       "01011010", "01011011", "01011100", "01011101", "01011110", "00101011",
--       "00101101", "11100001", "11100010", "01100011", "11100100", "01100101",
--       "01100110", "01100111", "11101000", "01101001", "01101010", "01101011",
--       "01101100", "01101101", "01101110", "01000011", "11110000", "01110001",
--       "01110010", "01110011", "01110100", "01110101", "01110110", "01110111",
--       "01111000", "01111001", "01111010", "01111011", "01111100", "10111101",
--       "11110100", "11101001");
   

end package Code7b8bPkg;

