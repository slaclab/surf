`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
MvH1+ext0W/9Gayularhe2zvdFDkB3VRF5NrA2mCAadeWWhR8/Zd8j419ypmyHVmY9DBjIG76z9w
zEuHRVfJ7Q==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
OiR9k2g6wPZAriX/bBytrxdgko1kSCAbGNTq5O1LkvJ7uS5js8cdcxvqtGS56w3jLnjgNoFVSsXs
QFOrF0IcDepvltesU7t/u+RbtporZxINnRZZeXM+I8osW44IiK8BFWkE6ybFgGDuG9Xq0PfTF3NF
Wz5TDi6YX6BDfBPI1E4=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
j44dDJpPIRMl7/1Ic1Af8fDaw4DdXA92MMSTVik/jQVxjTxy487hOdu3GK87nyCpBmNwztfHGDbD
TVJ/nkaYIs9wBfClxorUgenNjscZ+S67GCL24li/r8INvXXXc+F+HyK2+O0qm/FtzJtbSY8Gc6vP
dWmQr3MgDMHd14NtwKI=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Lia1J8liJNcDaSn5jpXIyPC9iTTpZyezvyfxIx3S5Gw7+IX3oSNWaUXa58F9Syw5YLrrFirADtrl
5IgBe8bpsXsf+skFpWO0Dft+cIxRkuxv38jhOYP4FuXEsq00lJmbl4E8hdG4qw9Dv9wkQGEbGy1B
2ME9bEgAr1Rm4lXDz6UyFDSKrF8CDesAtNUAaO1jBj97iN+AbnmCfRuQ4tbrKnBiTe8KoLjn5xiH
lnjCTs8MRHhTHaXapfvU9SMzR7AB72kV+QfOQ03fmWmdQJrt1fbdkAmUFicuZnn+YBKBlGXqRKPI
2Rdml8c7K5c7lsGgpu2DFe/+4KSRQ+iqDI6QKw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
I3j8XINxcyMnvwvw+5eoUv16lgfNprr6kpzTKWljkJjcGuwS1Uno9TFu7I0+54dXnXjD2Zkrs+On
1cCM1Z703dfvnAgEtPvJxKIcTHpWf/uDHvGEMpqjZL/7xusuLdD0WT0D3JqktVLftOq7kloB0inK
c8yrftk0g7u+dTVONcVjAlS+k6t0mgNuTAIpwYO7jDRMwImowq1ca92bwJiOpEEq6uK+dKl/fZue
dBJces4S7utetZTx9iez2n6g3FvDQ2FcXdR6eFYQfkDCnB89lJQ5zQCYaah2bqpa3z3/xwpqbzBR
KYfFISxdgoM7n+cUkvmJYLXefY6N815rYfBTjA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rdMteE4bQ7bs3fvZa2ez95qF2REE7/5oLG5IkDbnT5zGv7RJDeZ2jgWAJDIfQbgqutq4zjuLCsl9
uACwCPXT5Iq0ZXfiSnHXzsicuXyFyTlZWun2iNACNhotKK3M7RWXFb/Mlye2SPcuXfRs5bVemCIa
h4CYt4o0XW4Jdw6kYvxK+rtaJCn9qUtoV94nxTcuEnGGz4KmLfKPzvfesl6PMLY56gLzzuAGpfi0
2gjdT/S9B90OkqmnDORaIcKzArypNrXVQS6h0WmBI98rpjd1P9oi0K8M8biPYPudyNV+qy4hRPav
/EB+T7bLaxLfSGc+/AUd7uaN3L6Le9JqtiSUrw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15104)
`pragma protect data_block
uBs9wu98ujKeFiGYHGE1n5TTSj1VIpEkqez7DF6OtwKUdZpflvZ0ntuHkpL51SKqFn/bUJQobQIC
8aQfPK+fE6h0/2S4BmLQ80zt5TESb350BX0eNqrlLp+YIXxEJeY2PlKb3+WrY+hElzIuW0Ov9F/u
cs4rep40PmEzRQZodV8xRDrWhTuFAff0irA5gTFH1Fu+MQC24NPp+FyeJIVEGIEX802rSrARRAw2
EIQtgEtN9+dwzVcx6EmQ859PpUZJYaJYwLD5HaeJDamdyqCgwO3SAXEXjtTFbEVi0LTYwUglcYhh
u9ZWluCwu63mRyw0GkP9ZibrsFX3LEDPzeXorgCQvnYiX4m8tSV9d/jxx7DnG8xTgTlsPeZWLe0b
qbLQ1ay7zQSBTf89X93QC4m7+Z2OVQvHoPwdNoGE8OPfNwy2bfEBu4d/rCA0eJM4O0nknfxKK6b8
m4KHRP//khfFiO1tDRhNsmbgLy4flleAfMhDhdqTNWm3lgcAX6v4s9QKMwEcfrpR9ZlqDvnxS44x
4t8wiBgIJ/2Y5Fi7JmPUELyzyvsslo+mQXvS3JASoXh/lJ1U2yBZCc6wHJke4yVyuniqCYiJjaOZ
JjQvlYw52q6XsmlWBdPhMKUi/HFrJhjqiV5LpP+3uRyzJrf0S4H0W57ji5p+7YqVafHWKMZaj2Ex
0XV0iqcB0lhB4vzEDaqynCY8k8VkKjdlTAgGeTtb82jAoXHOwP2SDzFYmRF3RTv1jjGeVCqnRiwH
7npOrDNOGTpHT+Gvp26npSjMqe/arth8hiWwSIrseNZA2hvzQWiPC5v+meouOVX1y21gCCNer5fT
RzN86InUkR64UwHoQ4WplUafoemikosbqS3V2qftzUwQysShkDIUiZ1T3XVsV2IdMmWiMJ4Hh9Np
bT9HlgxphzKNYeoULT+tUAS76q1iKGJCahFspraE4T0A8XGbvtOAI8PcDpXEjrMXtGyvZrSjrLIp
p6p3TiPwpT3xcTbWoXUyDt1PW5F40EYzRlZgHyA7RWgKNA4TASJB2C/S2uaxpzdgGqKEsmWkWCGc
R96LOxzzr+2nzMNmPVCXsK/7UU2lX/VEgoSosmmV4PFztJw1JdWV0ZWco2g258Bqgf4XkR4f4jKS
dgt9TQbVT+vkFPeJCAhjHHR7r5LikyN4HxRY+jPdrmq1MOo1ZNEh8L66Vx+kOaFjb0t6T0ifplsk
Q7eYQj41VNHk89o4KVDbLhlmFnRPoyWZEG9yYXKIk5T0Y0etVFpZQOTx5yxCT6jUq8IkXnrNe9fe
DfqxdlsYJKzLwsGU48mUWkZBQr1C4/rX3Z4Re4kmB4X14J3bz6Ju7DzfJoiSVeYv775Mh37prouP
mFpGHwDNpzSu+wG/kJbd2wMuqvx6ttXqiWdD+AQ8nfsZ5j4LJO0y+6yUvmWNtrulr5GkgS8o8cpB
05SfJnXLjRVwLfBhZ1dwDEXzT+J1ZFKwk4vjk1kPP/v6P66d5byyiDZ2EAwcE65bK4BozQBy4Z72
9bj387VTj/auA081Vyi3acc0GWgcVpV8TuFEuDyYL7MIGVOuyCXT+ouHCecyYjX9IkcO/8SZjCWj
sTx6wMWMcYFQ4AnEPzooJk9pCWeaMHddWOwyxZqdZYxgIiBnlNqgic+/oR06wVnfaZttKqsHrkDs
Oi0+ynai2j4IfOC6Vu++Uu9Ej3x7P82q9QOglNRZB5egco/nxSNlxy94EwO94R6RWt9t8ZIoXMya
+tPLvNLJaLDA3Buzs4wGtOs9BjNzUwXloz738LpcmBHmeOBPHOx9NYd2ZRREm9e+LaGCxkZztYL8
o74AoOb9vFCZqMrOdnPaxl8c72bbKWnOWD3OXThrFHxzMvkWsjghjMIn3sDTquFwh4dlX5UW03qS
MB+/Y5PBP/fwV2/Woo7+lal8b1cyRDUWPHmj+UX8eW7nlucUF+a/n2NWBxY9mWRLOiNB5dwrYnJq
LZ/5+Y9PakGAfBwpoJwtXl8YTWheAsTk+5xSTR9UA4jeDTqyc2cZnsAZwEP4P9hJHA7WbQWDe7AE
sqJsoQDQAImu+xkyDxNXceIfE0LKb0TuBTtB/PPBLF8LDSNOCsQHyFMIdMry5KKtqB07tyi6hFm7
8DDoPN0WK3P9RvYi67+cqf6JavOaBoYISBvJlqZMOPaDqU218jSxBQbJ9lYaqCGy0Wlvg1ItSM0C
VZci4kuzVOwtwMRyEyBmrqy53X70+V0T3+naXpbbpDv+cRNI/rZb7m43AfTJa/lcZq7qL7FkaPCx
i+mYVeslo0txBkygnT0aZkr6iaaL7UIc17fg5V6ylV/PmTwn8yxZIZCVTfWuhOqpX/vYYmVqdrbO
LYQ80SUW0q7+S4LCLgMc9M2aylQlsetIEyfbC79fcS6YkoPkcbh50HFJmGL0TGY4MbodZRvgLUEn
BGQKYhRMCHq7ju4YT9ScGgXhA2EkHLAafkiRW1CWHmDgEnYzByvTSslZRQwrh5M8+olSicqurwAP
waavw0rVBQ0ZGFwdX6Cl56yHo3gtuJY6/hkpgv4MwGdPJAjB8mxdIML1dvi4GjIv3LYvAaAAufBd
WJlRQchUnjIUaezuQKjZZ2ExqXr6tur1nfRdyQJRxkKi8ntckxJHLu+m2aq9mx/2Xgp+OTexmzeI
or/hh9I7OPx0LXYJiCXwCAZcWvcRiApBdXU4PJ8lljs2F/khFXi2eYtL4capH295q9ogrECrB0qW
QLHRFBo3fTMZTKDZAb429w5LzjT8eDuGQHdUthXT3D7VZWmrzQEZ1cvqSvXwzpa+VVo9akSjf2kY
5fSQBm/BYdqYV7oDVfqqr07pyjSWal6o5kXC5J6kKyHg7yGz+i72gxA05cCK2xteeAKcYbTMtQ3j
VEKIbQ2Lb9Glp8+eV2wSa5N0jowKCnjJiAnygODDEwUQvndvZkfFds9e9Te5OBauJdIi6I+xK88a
BNbpNxeBWiLmzXMeaOohIzJd0DcKUv3Mh+iwUePHlWJvJ/NpkMMgojtH5PykXb4SqPjFUzzZyndY
7J5ilBggcGUWfE+NMomy6IAkjCaOeced7tQD0IDXd8EveVN49q+CzzIUhvlqyYoNYN74tVBdUHoJ
fBfY1MhSCpoVZCVCNOjs39ZwNe71wH5QYwr4PKr4jX3g3nthYqpzc76DKPCVVzTNGpL+VxVpS29e
o0B+c35yKUitXmZLUN/EZWd956OKmfXeTCnrOBQTP0qpbi11680xcvjfxDcKJnVE4zG8GmpaeBOj
+RW3PQF+8BtW+17xHqa+p0Vo3HYeKBMdBKYHxQbc4FZRzSpjwAZ2TyRExwtJF6dicO91ZUEGnrdA
FNc+1QeWXJFwdc3bQ8SJwBZ8fQHi6ihMCZ3/eipjgOqu5qDsyWm2zJ+0AcoR93+nd78Lb5LgKTv5
hbCUZzpwIAFKNJnjwNjkZ7vt0qSjfXokH0g+dQsGpiv2GS337wplHOa5qL5E69Gc0ZHbQdsWmwry
A9XHYwYexyEh21cbtmc6zSuYBZUnx+Jor4A7sdGxhcesY0EmVPzsDOikythi6uuxEllo1yYnwkPn
UgAAyj9LGg63jLgBR3q05tq4lr2TDgcNDI007XbDaLoMqN/yUxv9DMosqimfhfk3poXclabrR7Jc
RppZe5+416SNA4S+M7v57/XAdN+6njwuCwxF9mWbd7Sdbq7urZ6t1tbOgagqKyvACYzBsE6XbIMc
MAcK1TqS+5TEgm6PP2rm+IW3jz229u1AtupGqX77ULmeL1NFb7tTwdZFPI40rWX8is8qe5KScwBe
V1krIoeRxblS7GAs/Rh8ssRhTVf5ocT2yVDwmHYjFzeo+N15WBFMNAQUwGGhUg30/uKtuJ3XrJy5
g/wJeogH2o3Knqj8k/MJJDe5FJzV9XDjQw15DCKLHOl4j3KtpaMWu8uSK9Cmkan6v+N+5IC3UFaZ
DekvAmA3KWWVSgWB5UNTp7yK3lp+83JNIFbz+pwoVUZRuXwRLN74BRNzPAZWbOB7qSVAMlhk+x3q
TdkmUrR72BPBSCMHNNeBPul2CGjvGwhbNlJNiV342C9OfpjTP4ueYGTPnW+5ArUqWfLHum7GZYIl
y881Whhae0fIPlyIRM7mJrDPTt6VB5pi6h9oDrRhKTkFFr+P6mISOsAA1OyJe3meldG/UMwPLoQ+
GwHhG7uSR9stU5lN7u6r4IjJWqF8csQ7D8GvGvyO3FL7SVyj1c/H4MC7YzWjGMbaobznFe8BMGto
g59ZDH/jpr6b3A0vcOYxwHqx3cj8D5v5dFFWSqBjF83LHX07BrpKGEofYBivzmD0aURtliAC4Skn
InO7g1Uid0L4q9Vj/REiZbRTyMlo++m9OVATtNfI0WM1lhSTMa3/HmEH8TlO8HsnFMbu+y/+1pd0
8f0EjRs3QjwuDoZ6CUVCxWQ0GXtUc/3K2PLatAxwHDAObmQfXXx1++0P3bggkxQVd/42QTAbUhjE
wLMD4ETE1o2/oo7q6bvpQmhkv8SlnMjTSTCWqRFIKPE4pF2emCVSOxoLeN7edRMZxevMCvJ1sNyV
CZbB0MppldksAzZ5puvtwPu61DKv948CvQQLglAwCEpzogm5J6mD9XA0Dxocv04biDbfiVimighO
S/QpPAIFN+r5PgY9v7/S91uZcfHVTmI1Mkea1dj+KFhsG0R45qWcENzhDObKC3hVvR2Zp3e2o9Pf
16JEWJAbrSFXHTX3/D9hAoghuERttqPvWehoeVAxs8TnVJlD66OuVFfjupEFF4giY+sG+Vmj6PDN
+h+ok6hZuHoam8nPDnEtasursrsDr6lrXrTpu7MDKBWLMktJt6521zVLULRCg6hAkIQaDLX372kO
N9uQvsr2k70DmEIbugufPki/CP0B5/7aWn7i6oCJpgH/HsuGncpRTkSkYYPE1/oEDNhwsnQ02Gqs
Xro3xH7Y0OtBWAcA7GvB9A3c6I1IKjnCg6K71pnsXYeYVZuti2AduBfOh0aJ1gXmRE6t6N0HwvcR
R2K6eV2uRwYn0GHh64hPolB2a0JCoNRO+0x/ZXrFDAp7MX08KoTwtxFV3+YnYc6QHWv/YTzGh0LM
ZnEJSiT1P9Vllg3S855XpR2fbY/36+XDkCFrhe6FcZu5pHpxaAFOlinD1LLIvc4g56kzWVeVLQWs
z0Ihu2fZY3Tz1n3kJuGjckdztX+RLQWkL3PN0SuurKI8Kev/JBquQUuAXXSLSJ9gQUDTieFHmG1u
KX0zsK5a0BS++++a3jrc7UklA7HjH9ImGGxDqWAWaFPySnIX9Si24/gEp2PapbzNF9QY+Hcea/9G
+B9cryOf7xqlUOjtW74Zl2wpYeM+6dlhxYFmDlkbzCDNm6l01WVZ2vxKuW2q0Z6vJCUSdEgbRLl5
xF4fmMSO868aw8WNWDQZEvWFaAJmqlAIhqIM4N1FnhiyHl9SWUFkL98T5Bh9se9CV/w1aVOzPBcS
AcRVuRYrnUQ4o48t4jBKE1jAm/gQNHPExrtrdCZBeLfXl8jt2ZMmHk12xdh1LKgYaWwg9+Sz4jRI
AVF6erdyl/xxFRYibZVhwyHjcG5eKkDAU906bUonxCozbjZYJOqhwMx20zlATNZ22D6vOAsydsdx
jAkNIkyssATUfxypHtJohXknivOG5y7nNi7YzvHvCh+iARUyVMvuBRo/kgw4SXmYDvwkmyPO6W6r
SglBYUR/V8qYau8rw694fYyGQ1nNfTBj1fa5VCPlklakguAXOT7yS7zVyag+EUq03SVjR6pA5bxv
mRN4Kd5EclGUWEFPQLNKDeCzQkRHIW/zQ2rSRddrkQooNZWp0vHYaMUf0RJQ+cWd4It+I1DZJVid
GbGrUQXXrn2/DC71Oj0TbZ9VjF1mqtB7uuXPSiZISLwrD5/tkHZOa0gsa4RjZhddpvv9eiLm+0F4
QhbKxwMug7ggwFKtx1qj5y8vR6cT2bntYN7jn420l1MbRgZBrywsaS/3GIt7Qzrh52flb69ifbju
ZYxf6OrzHfb5mOPoVztpbHepWJlVGsu6ni4SXZpMljIRQAF5o6s1RXtqa4sJCN9taylZDS5osNTa
gLcFEhq9mIMQU0GPCVqGaSCMIq5oGJIqX5CSoru90xWPlzH8LDxXXS5MZ/qtoQrZQCb2GkUy1uUY
a5Kup3wmX1U9sLtY5jdmxyVGV41kljR0z1CH+PAjuMSzb4mjXQQqEPjbupKG2komAMzw64YnUqfR
YujatTAJsRTuGTHxDUZPT4ss9aDx0IHD5ogJWPKpxJtIHvKDr5Rz/bzpIOfRlu9AXZf5x9JsvL1f
59lCb3avRgCmf14EQgYpkhDncxiRbQRFEFPLkIPfilWX45xiET1/dYtM73DsgEsh2hzJ5tI91GV3
giyRDOu0O2mcW7aM7CD+RLb1/6fFBwHHXbLFJwJ8R0EL9ZQNYlz3Rmwf4jOCUlfuJ2ax+QQWzpgx
3VT903tt7DqyL5PipGxJ2qvwEcbOOEvt7VNtNObsQpVcMpRZzVVvl8Arjc/iwPCtD4An4gDz8zwk
DTCeplsirf/WApZo4jjHWtcL3IEIMsmhCrNuiGKD8JyprYhlasniexqJNQS6aGGNx585ChAc4CNp
Edqp9hzwbGUUW8+yY+Z4I7k9q/WqOdb7ZkuPaYUGIAAqjUypUoa7MX4bXXTE7IPv7zH8goF4siO8
G9EiNyXzD1l4+jd9GUQVe0TpDO/1NqJGyy3N3Wa31thj9SrgBx44aGUTGx1T928Y2ZaRJXa+dr4p
BTiXP2sp0/3RFDtZ59r0tizTko8y1F7Q19y+edwjfd5y5c7K6C58UObkg8vRgzTAilQwmgsZr2Kq
Jn4sQp39gexDgrGzXx8G/QPRdUl1wEOf5LZ2pDICCIzsuJVw78l2YpKkEzCWSOessUBvV4CF6oDk
5nGxDdNfdnAMFvRlmsMcztO0z4943raOPI+epUJRrNN5EeI7G3uoaEWcmPliue6ARc3Tp5dAkMPs
iWokaJeLWvkNg+Gh0OuluOsu07tya0jhsfIAGBsa3uIL+OW4sUZCsL8ho7ATiX6VC9SldLW1dpAO
sUDshYKjVxeNjQ6tEH/iOAjT7UzGpoQVVNigmwAsMmQv09DL4r2qL5yDj3b5qM1/9j/avbTionVU
8GNxF4NFfY1cTioafmW1NE1GgvpN+5EecIw3fYJP82dmm0NxFbUAKRR3bRoWOoNMUEzcGPKVTGHp
NVV/NJibkocmqz/FSen4VmtOQkH5hQmvjYUVBdqJzZx6/84VnRU9FU7AZKY+5rQuTHd5UZ4YaT5y
k62kP2E9IQNBC22d6m20JVsmqWi8FgkJnBrw4pGH6DvGJWgsB1hOAzYf1nQ5uFpyf7rrl0jmNa30
fxq7UpVwXlnvEf9Q0HDHKgpf+fWJ1i4uQVtWIrFmskwHG3wMsR0o0CS6bE27BbzVRf6YzMqVui92
gVQGMxbOcbP1w91F2FLK4EqF3UOtqrWG/6JlqeLxC0hfj0h3IlgY/bD86+vYpKIN9a2AWqfZ+lJ0
PVwurpKe9OSTFvQY9yATyJ6rG3hs+T1O01Uull3HCUnx9K6f4m8sIMAqvOGYts1kmQuGK+m8P9El
sJgNpTtoyZSfGg6kLHkojsaZa5VskgnEtek1X0LGvADSFnARCloasdyBnEmSubzutWV1i/Y+1sBI
3UFu2neptZaszMFqKnepHTQMyIel48HJNLY17zQVyYQStw8txBIfWuuXsz7nap2sCFmF2Zm/5fTy
Uoh5lshFwMb0ypDwB5XndmGKPpZQI1mmSm4RdplskvwQ4r85gMRnoeSi8l4ZkaqSQLo06z1ehLRd
tQhZVA7sU5/ZtOeuSYflAN5zpntoQaF/t0LchzfQCL1XyjUfmUg4tyOdOx19UI0pDD3qubtvKw/A
Vk+lzIru7+zvQCcmWdMuvWYaFq5BeBboHpivLgYeyBwIQQjEmaXLHrxSPaFpgph3eCSgo3jxJKlx
SQ6BUTrT3rkfAmcwvso3INnud78bYXCRry9MDjwlogGnFB7zD3Pba5Ev2pBiK67euLFUilZypU3+
TW4+ypTBuNKWAvX2uAn1LUtnDvU6qADZcmaM8torHVysctnqg+e9hsh426PlmsQBIjfAagj3MUzx
Zdj6pggdYG6pmHJ/axPDI/AUE/k1blS0w0tr5bLdAJUeAgCy+O9UgC01vx+hyYIeAbnY5gc38h7e
e2NP4E0OHLD8BmVNWLjx/4PT+VKj2EQDcuRqgjMvgVvC1zyPCYpymfMAxdl3ju69eFzKsUxSWaQT
L4TeEAgUzm4Z2QBeCFCicwexQkHmj4dv8nbH08N3kafLyFJ896MizbI9xXhUjThskzo+JaeFvm7J
6r00WKu572nvwQKBrWsbHx7qeyh8/t4FAsPUV+ackmVn1KYhExtVArxvWIQJNZ01ju//dZX0+VSB
AsJWI9MibhI2BXioQxBim7MEepHvMHqN1ekIYBqftJtnfw0WCSNBFhNJNWn+0DqZwS+5jWr5trjt
iXL+VoGOqz3gBSlSQfqsC0Rn0coieMKYdtNjYsLr/UH4C4T4BSDI54cvPL+7T5zTwOqJB/rCiybz
OkaDrT+mtgQkWP60nLGTcxIS3ZQj076FZs2bODPhwcykB/UJM0+patKB8t++H+WGaXMRP8oHeHeR
QWbRPCKU5XoW4HLJC2RBMK3LQA8a+M5N9Vr+5MZ6zn+VCkboVow08Lfdqro/UjbhYbmK2Qq2xQs4
KSVp6vq8gxYAW4B9nm4tGZHmDOyHYnL9VeGoxQyFvBV24ae1DbKc6W92/CZj6wHNMXsRwrkvjJBt
HxPguPA8cglUcBsWMCJ4GpmnWExdeuRS7sTselgDF847wFEj47GuNASMXYebTitBAKWqu+HxdbZM
/ldBUPGg2XsteEJHlnhVJviagzz9imBvnMfV3JikNaSAJvEL8iU0IBkS9f0fGhRzJU3ckxTA1+vP
BUKeaZ5lhgR+OSLZsyWjp4umtouqc8lplAw1gZnPeVEx3K4vUValVlD7vsCN3xzUctoNxgysGw2k
M54IiYsYaOpgQzLagjaWfQOaJqAgftHuRZ4HuHAXm4quzVH9u/6DcE41jqIWxtEnAmLzFETvT8n5
HWly/MunZD7J5qGNIEr8kLe4RKXCO/04dVF4PCOhpi86OTyyMjJNd5tbHV7vB/DpdYQPpsyLUh5c
Fdwhyq16k0HTQUDXjxJhHiH6yuF75DTp4/8CYAK+R5ail4TKFcvDuTuKvWYxr/9MHQQBoF0bWlkW
a8ZO69So+cICIZBaY2fVE/jzDtIiRjg+3cHj4iyQWF0LFBNudNSKuktFGZQd+4ywu9qkiegM704k
HgqMj2nHvFuXi0t+BQn0aoO64RyFRPZogGV2ozl0qZltdm3jolYRxwkzmebQEQJtrknV55h0wFmR
dxibcbAjwgaRnTQgsgPuJ8DrJwfxZjuCFCj4Z3Pk+X5G0sWuK+61hqQr44ISbGWbqrNklWCHlikr
M8R8o2S6LmSmMYniKM38KfbpQjVr5cwh9YH/nCbRDnAAhICH3FHLjS7YZXWoZd4YXKH/+prtHbXK
RUo5YHQpsySkszjOKVZGe6y3i9+YeLWP8s3AOxIoWWDtY9ggQry4Axsn0dgqTSDeQqLVn3fMP9vs
YV4oQ60ZCWsegHMv8NyY3kO3HNLqkS391+CmX5YX6lTDSL0RX/jQWsFqfuyac+3hf3/bu9Cpxje4
nlj16BtTOUgT8Ban+6yyKjyGpJWiTXq2XOTHXj8kLyeqPtClOytEmKdcukEjYe528FUaX8YK0meU
HQC/hmkLyxIH8NwW7lLDIGXLvQyGirTai4R+lxsbomEACs/obwTdlBP8uoOiCBN9oKzC47irNTKE
x+1L+ekOKkwl5nRV+LoJR8xchNBs+dcYWJ2BmdxIgsbDSPAUdQXjXaiE9NClvrkAs7q9kGBkAqwD
PlvJ+GI3lA6dDgU+vG7Fm0hJvwpmIg3BHarLyNw+Kkha8Ii+VZ9Lm9Rq1OEMaR5kpHbTok8Svu0D
eMiomlD7CVL0Kb15Q6ixcQqfzfD0H42bzZevcxD4nNczmEhhFDv+O8NfqrLUq9YkOgdfOJJYSQIY
OIWHBjiUeNvjnxHZVfBWk8E8FaTMoi0PRcnAMa9YQ3RTlJVOqnEjMRANQI7BOhgug6+IfFe9ZKpr
q/h2wJii6ECKV0Z6s+JOdRUlaTtGvfKsh4p7vEub5VBXowQGfuc+KiT4Sp9jgJhMPyGfligocQza
RhH4pxhhuRFD4u4p9kUkOSI+VfHo0McqZGs7880wAGDiPBmM1F199aJ9Ff02jvn9PtspSITSk2yi
Y+hNinYxV+atqAevo/i1a9Jy1EJ5PsRgB97QAu2lLUv9OdyVLxxxBjYi7ZECz6UYD4jcx+X0FhAb
KUJc4rYwLpR98Z987Jm5ZNcz5C4icnHNYES8W1wTsJRYlApbE9ES7o2yxHD43KRWr7e+y/x49ME/
MBd1DXlOY61XhMpezNfkE+iblcxIiERC268e/9m8MzAY67Wz8eV3oxUOLM4avYN2aJkBk3mxQTSn
6NpBbwTHiIHagpLiDnt5cACYOktS6/SELJVOUqfJfdLPYuTT3XuckNqHdOjFbK/iOapwpsMpYOVI
PxHxwfBG/EFkPJTuldlbJi2UyYm83qIH9ABK9b+gJgKgm9A+v2iFjREsoi6QBpBnBR06bNOuDO2P
R+H9997rSDPo4tkfUiSoY6eYc8Zvugh9jSOyK1JyuJmgtSyn5AnhmrN8TgqoLZz49JgFZtfGQa7t
RGWCVNBWJ1GeSo8cClRz/d4ry57FmrJHlBf4D7X51IUzA4VPKf0NGw90OroWmxSEvO/UdSHXrSb8
rNMFjal9NrOaA2NdJyUb/UaMGskOAm8PmdAgNar3aOMzbuzLlJ6ZWDnXyp0ta/PNt/ZqTsBTnXMb
u0djo5a2r3mfyTFCZ64Bcx4cx92zKTHpuypnLPNPJCbeD4nH4FDqf8mnyoGK0E0XX0l1xm6vvY9f
3bTRTlpPNygBvpFuWCbtxYfVYu76Ho1tomu5LImn2CHUM/P/IlPhgeHHkxxBhzSd7ISCBVPUPawk
2gpDBAHLvBlPDhURoH5lyVO/cUHof0o3avgnV9DvvMPS23PKFrcxx24Up8TkfMI7+0lIUasvx0er
qEupVkP2sZbsPpENtlsrbD9p8AsENh5LHpMtcNIIVsllw/MvugrmIHcJrhnCRtZGk2fDB33MTBQp
bkKFg/CIjqxS4XDgE2zgrGId1I6L5xu+sWNlPjHEY7+UmQxmA3Yz1mxbxXN7EXWzIIJdPi8pZPGE
DFn8l+1YX+7XTlTwr42tkBpggfvEoG3+PiWy96NJ53ab3P0e2u66wMOilMou7bwo0hCTgsYNPZ4o
UT8KcNzOT1OZXoztvzpNlsV6Cs1szY9tD5JN2Z6Wye6L07PCAJcwEHTdFvM8HmhV/ItP9wBuSYJF
JGio74XkqY3np6EaqE/6Sig01D/GIMYB/x1MdHbtyNJO+O87IuR1SRPCtCM+wRRFXPxsy3ny50WQ
25SQZfPGbqwx5UDmY650vcWWl/EylVZwhG8J9axZbAKGx+keHmS7nkZfDYSOjvd1rkARiApF98Hd
Ofa5NwULOXeddtUNtOeOHvyPR4jzmVfCD7dJiQrgB1iJmZnHHrXuBIqHHcxSkQB2cbaTwQMVrDag
MlZ0JB9FAoGHixuNITKI/nKWboS7RyweaCOeMCd2WycwRNVWTIXMSQhmIStJS9bRg4JjsNVA5QxP
Oe4/cX9RY3Co5gKz535W6IF8GQkyVE3QdVgMIQYt3XFl331AxWo4x8tDpZ06WTrweZaHV+ebx5Qk
RyR9s7vEmhh3RCWlEzy7viSDjvJIJxJSYMkMriKcjMSb8zescK6ld06o8GO9l5jfIuO0duhL0SJs
i+TC6bmaUSKGPXxU4C5HBoSSuYMCMy49PaDeN/Ajt4d4RrIcSEsv8Ox+m9JSraEdkdbShm+9lnLn
HFAY+fxPRwUOQc4x2R8ISrVsSWNf1BE30TmfIzQR3n+zMGdsOgTWqD6ICN08YHcDuGuLb2PO29YW
MaVDMoUli2GSuimVnIgZ9ZxqelVdiCi7lWbtwVnSEZuNbOHwuNb2m9KBWKRzTfs0zxd+rcmjAemy
CHiza1nKjTvydkRRuYnJtYSi5eAd/iwwOL+ikAODQfX6jdl6YGDfKf8ubNYVp0d7pEwhBfjyyht9
xHIJ4Kt5R9WRKZQFDatvGSjnCzKlF0JGxepzh1e/CEfO0gpU6LsUFV9Yr15O+OKr2/vQSOsN7071
Q1I2rYcxG7BzkchgMQxYkw90miQYzxGldlhnMPMZyE4y6+0GH/zfufmTCrvO4BGBKs7MumFLLXdr
E8kER+fOgjd4ICOP44qwWvt4hZxQCUrxyHCx0mYkSTma9E4d2yn0vxqwngWKvH0kbodSPEHQfNsF
2nqeoLudMiDOTWNTIzWDrDgdJF5iXOHMDEA4Fjx04rArc4z8JLFLZj6H8Bd2YTs4T6RdZQFPNc/M
3IzpE03VdFdjmSg/Gc4+NQEqnuBlDjdzp7zdalkUAGswHIe0zeV5onObhC5dvL3o9VM+WH9ioFnL
pbEWSlgNS7yVFzoMnX6o645XhOfUQH8Ld28q+BhkNPYtiKh1kW88yNDNeuojWzUbLVdwjEpZc6y4
LpKfaY0178Dx45TOIKTt3WYIFYRFv5rTnY+dWlWRdBol1D5qia/e/aoA1/As8LwDgo4ZcJ5DVFIj
C8mO8XlIKqlMGfrBOhFRT7CS8pf64LY5prPmTlUTnTtftQgAGJBc0F8uy5j6ZCz9Y4l2l3RDZT06
Ssc2wvXcn7lZ3/wnmzUjR24EQ8fInX7H1osYr74ifJ5N1ZR0pNMDxSJPDY1jn0fTC+CJ2C8xMibu
gydLdb6ueCIXj/5cWmjm6cCksgoPRkBBpEYySCTVpuQsd7gnKTgdqpBjAbGbnYnxgAZoDDFOWhbr
n9NixltncAm7OPf/78souhJeg3GebezHMnocZuAmNCA5Xi16Hw8gAwsNQKNNQsW2u6m/7hsZY0Jc
PggUt1mdzOz4NObMJ8vXwljRdU8JLqKIZFFtQDg2gq4rlIwQZG3xyfEyhZJl8Cx+OheeR1kVGZ0b
GjdkF7cC+mJkHPDFsOuvUHlf6hDzK+znHS1mBZR8l/MCISlXnhTqmH+KlIHyp/khfCvCTGhD39Qv
rFidkAJmomh2lCgjVUa6E5d7AI1Fq2NNHyP7ZAMeFuvGiq/RoYbaqOSSSD0CBOzw7s4TnzuJXXYN
4LSzcUl1AhUOZNSvY4Mb3J1QEw8ipWMMH3knOQjQbfMo5z/s3GxYZ5EQJrlah2YYRI1Glh74PxB9
yISilmAN5Z+5T82v71a9K2y4qOB2KAaV2Zip2FQMlAnZJlEmLKvJq4C9/TE3cPAJ1GRT0nOKNPbz
BNHeI1ZibTwqoPqyt1CImUgfzV7+n4ul/f2dvNfDGsRyAfncYTWFOtZefQ0JOy1qzbQeWcLcr9dP
qGr0QJMp43/1sRePVqDnCPhMEE4sno9Bya/QRq7XiOJcSw1GgEX18S4Cd6VA8/tq4AjYqoyrKb+A
OaTklOyo+eLp4LNhpy7DRZvgpiRga08y5Ya80siwMpNtBqb+A2p+8OZGkb62aIREPiMRlOCVPBvU
tZ43BX0DEtHBwVAvnEsQAPNFfAicgXVzx/CBTQzG5pa0ZCCN4NZiB0itmmnFW9EpoZ9H3FBHEmjI
WqW9vicQOxusTrrz7WK0QGB+upFvPbBKn6rHmQeulZUKylTP8t1hrz5rKPdlcz1oxSUshrLd36oI
JGfFXeA9wgaIKqJWXyZNg1zEGnlCO3rEFE/2vA4ckKIg8Ak4XdtzQHl9b3/dwAKyAj2zNkD3gQtt
yb/kPgj9MKC1fUzs5JB5u/8dDqtrx5TtOJfEdadtSxHSySA6X+Y7BWYyqi27unKPYje0X2u7uMBu
XNX/XbBr13qGrq27WXxbQPq2SmWMLaRfWeBgG0uvrdGx3QRWnxdK2WZofun9I3ZP3pCzh/vNxMxe
ElnMDbCxVbrzBekn/1Lf7yJsz7zBPLfwcf9k2TP7nUH3oMyrMQrbifhwHtCPFUg1IOcUiffrElEx
lOEZ4TJlvJV/f44z5RCPamqXEzV9N0oDgXLAf+Nimyhw6bb1dmVsCC1k1h7ed30dgxV9HBRrGZTe
wWRMjLyPHfvl/7Hn03ETqj/E1kpYjfXk3n0gIXQ/IwRQ5QkKJM1uTjTTTN+kwDH59bfo2SqP3p2m
kew2ZF8GxUpuutCHqggTOXIZu+1mBzkUH/zGT9iGBSMmYD+S4XgwTrKyDBfh4jBbRPAjVpb/iJjt
odEhwrtjruWRnWBZHwq/UuM6fLHHbW4Aveb37anSNc8H5J8SJEqf+s7QUd7biUMgRD56DyINtSyL
SUnLPQTQ/6UfI8ZrkbbVJ2xcdEDqKxUD8vLNHu+5FD0v5SLxePCnaAQ00SpHdFAgDvUhJI/q9jox
e3KGuplqloUBexpEyl2YsFWzxO4+thzbMVe+HxFuxEaXdwBv2WC1MTtL6ggWrzU4gBEDqrqBrIoJ
u2Iq5MyOQbkngNPl9J4YynGu+sv9fM0XPIEN+6tw4kwDsJManiNN5bSnBudaAD7HsInaHrc6W8xU
cP7AkF38ojbPYnjHEJKJG2NIPJRidoAMP4s9T+qhxTVCNmyAdAMZXabWJry51cjHZCPeEz3tkXbP
5FZRVVJIcrZsKXAUsu51TLYzjIwGUC40IcQxZBSKcOrqM3z6WvV1fmLbcvvgvkoIqzX+aH8tNOxl
DoNbcHZuq8pNkG+XxZYM4eDNopb3ZIMX9G78XmHA5FhE2Ad0ZhHSEs2ZUTFHy/qNWuaqsNTI7o8w
nITBQhrsVvwgfZUC8RpfQeKx7T8699W6UqraEki02/qCJeu+13yY3Isf3RsfjLsDa8nTK22BOV7H
U4z45kKkgIelpTRLeosfmEyzU5NS30GkhUSBESoXARjZn3c3/2wB2e04zDg3xV8v8ZrsvtFI+IiL
9z0wJw/1OTwOCllNYOuBdDyduco2MlF5a+rW0KznEwGcLRxUgYKC3EqaJK+SzxzKtoDSay+jztot
on0ipnajRCcjDk51DsV5Oa/B4FJyzQRgtgQ5D5+i+XFbMDUd1ApiaMzQu1VlWXSNl2CFnLE8ZCQN
/jwMsJMwSR/uGZwTrh0CECKrLCYb3oW/VG/EYCXahURDRt+X1bBmmgncMVJg76LhbQPuMEF2H1G5
La1Vgmoj5sN8hRABGRElO1xBtpZcinwKUUmocrb/iJoESwZcms84gaIEAoATddS3UPZug71BpK7c
s3nLx/U3dEWZS7yGRwS+dhFiAlNiRUNyFBR8GJwlcIJg22+S/ermPMsUh4j+lZ/7jOV8Lr8YGbNK
1JLTWfzFd5VIkBuRBLKZwyWW5xb1azJ4z1mk2VM15FJlzInx+6ZB1kjD7SnE5CRxkI746u+zlwWn
/EJdKCbjVtrYTxVCcLj872WxBoTu0di3HN9RpT8MbA3WXtq/jEUdWlgZ0svywfe8iXFmym8ffKFh
ptUoKprK+3pJMjS+ecQwg0ACG3MxP+G0AgyxGXwoREXgXG/3K5LczrlbcnCC4YGhymqaH1CrqLaz
Ha6Au6BMPPNMsLlHf2g2b4fgP2/rLZeyPlBdjBItyzsrneqFkOQb48XCmrve2vPzewSOXcu2BqU2
1V3UpPJnNV3s3nGtFUYT4MUhSBB2OlG8posQ/G8EKz8S5sbqmP++PfqgcikGbVmXHnpKJpboxYZp
6Gp5CuIp+qgj5yrrhdYrOIhfcKQBjwuM5aUZ8xgEGJHoi8YteHDUcn1gRCd7DjBdm3RU7ArK0pNc
/AU5K0t8DMkdFp5ykICw1V0hsrzYMh2PY7LyCPVbKK0+oADhV7HfsHcC4d0H9S2l9xflvJBn/cBk
ZjnZV6xfkys2VfgQGckPQWvnIK5ah4CuYhMTurOlsi8oKOAB5iKxDj4Li+OcFbvNOEqyaAMc6BWt
LoFZv+Wav3WQomrC35nHEYCHE0Eplfx4P/Uor5gw5BADQcA1YZscOo2aDoceHhYOTznAyjt1xHp3
eN5Un+aohdlMntuEhRQVgXj7v6Lx5NO+grlipS/aalskl2B+kXYhk+J1XPAU10z6YMs6Wtm9vPVB
N6GboF6d+0QVq64TEM4hMqLjexIwSCC4NcL2aXi/ujyJ37MrprURDOnfnOqxvkSjP5VPgpLKX/Y7
AStOR7+47njULZFtuUvnHSPz47f1gD9t7QG5s6IPOp3ZY6eyTJJUFXdYG5GEDm9rN8aCcKxGFRcA
e6fF8vv2ntzivEqENjwhyx86RdifmyXNWXVZRsWKcSUmLNP9PRXqybEjEJzLl77mX1s7GiksJ2in
g566jwbnD5mnTNCEOigGk4cjztGKZcOygf2vw6eKxCTf4T7+Z8ACHuqP2kRZK4CKF6pWeXAfTRbz
qXoNy/LiDjZefLaeMHqGu88QQstTVJXZ7osxp02vuWBY/dQ0168ATAUvTCkBj1f6bZYuAHKT7zJJ
pgoL0gHupIdIkKUCSN7CQxEMG/hGaDNm78DzR9YFFgqGp4R2SdiYgtiekO646v/EWhl846if4pfj
EzWGiJ6ccqC8LyybR6/NOWLs8HdzxDxl9J3oICkTFGUpdwGrGhwI4+pzeQGWmGUmkQbnn7sfGhgl
y90CNJuo/PMBwzeqo9ekxSf4J1wMQ6/kUSW0G5Q1uCsIOKsm4c/hq3iUPMuQ3BZRN1byVEFnyyBA
YLZ3iA1KAHGQL3CNyPHvnq1+Pw4o5wd5dnbL/Yz7awQbdYV9RcD0m1XzkBvCmKppPDLS4n28blxY
fLhOmCUjMV+KP0CpbS0NXzJATZVNq7ndXHYWfYok8wrKFGqLJXaKK6jHC1kJx/0p0XYoBcmtLPOb
y0DRxop8yQ89Syt99qvjvWsjTDF2oMqYeIqIOXRLATSUh5iheH+cTH8Oj9u1lhkbnMnq4o1g4xFI
+u7RNIFe3Qiv8UtcrJ9roUSOVFuhESjqM+A/xOb13OkioJSvDpEJb0VEbh3bPo9xTuxHfhGinWvr
/xww0Bm4RnX2VyjQP7IgK+urdvUbTOXbQuT8XIhrAatdoYjzzuDEjM4z3IEUcAeEHodbRbNCqjRn
2ADouBBgqAEd1FLytdQzoAXSzGaxRa6iR21bsMPLttW7yCp0h9xnndkfQeSwDtjGsvAUW6sMMeaD
V8ffYzJnpa7r3jCAz5ezSflUthOaH8990D7eQi15qABLkLt5bQVDSGiL5aE9/Pq+N21OBk+DV/vC
LNJF6oizOuTOdXHmlIO8V+GgxKiYc+2XSIlDw8+KqXatWxrRTWWfFpkz2M3y2JgwyMSgOWXX45Ug
yU2BiTEs5vXnmrPP4RD7gnKWgyG4NPMnIEgV34vAMrb36BuFKRlEdpR9EzxCUBiE65pYWZmgGzO7
yN7gwInpFiP82l06ciDS/dX6dFSkCW4SPW38TpItZb4fyhC5dz2sDRGuibRUY8vfb9+S91UgIxBT
zET/ZW+SnMlpTy99dcR+8CJ9P1pfvEhk2wmW2Kezukgq4kfvy5+bTSofis6E9IqCxEmvBVnHbk3w
zlHW3yggolYGdhs2lttj/U3Agi2KGxlFnbqYzDtYHal6exay9C6WZl3b19JpSRpMj4qIhYkFcwD8
JUTMlpAcByBWiwaUXFWpCS3bv4/SyrIwu3m1mjKn8/vpQ7q8912MPhlpUC4Kxg7kXdHK+u7cHEEy
Um+53/HJG+20OFQhTPEoERN0kWYNsbxv96+dOgi9xeiPAg3MI5MaB0JOMYlxH0AOzXNxceKgquGR
2G331Z5C+vk55BStVN5s1VsuZYLDqdi8DKhl25iIiURKxGtgLMc+2ayaenwV9KoJrx9GMFsC+KAn
cK6DvqaZqip4+Ozw4yyQhjXRVhnRHaLvORJxGTIBBNUInQVlcXKnEsjBLItOlhtWjmFn5GVVKhTA
HCkI510i2eyS+TjlhK+ptpn+/3cIV75GJyyGOklyhNof/yzhOMp9hzRS2I8epoypcAfgDDXBoK3h
MQ9cVJllSJ9CcfW6dId5QjmbIEuhEksUvMR6pKLQtD/46PYaZgTcdfIkgoChvR5tOv8ziigaku8D
gQ/Y4Xr3P5XvSB301wFMoD0/WHgCt0vQ4Y7zil3Mg8J0piXUl6ts3HfXNGMDQH8U9hKcBjwWZvod
YtcBz63slxp2EmSz6YmwVDJ7ajFm2wi+fWJgbhi7va1OVYlm2IlOLVGwdERRiwPGoXfFLn5TgtEb
3OxTcpCJ+VBjsaKaCnVTL8mc4YndMn5iysV/k6Cl1BjhVT0DsBXYMgtlYUoEV/JdmWzdtu/2Okle
RN0BBnR+HxLpnn0mNvnL9wn2W2gvtyP0v0mkckGQq+2pxNsNSzmYAFys9W9NZYTBtt8cSOS63efJ
hRwQheYJcJU8XfEjpoTR5c524o1Joupzn7F8fU8RCzguMZpc9BNVcrTcmmVdDDIJn6Ia3/pO/XOo
GrRQYn1ER/xm5egy90hrfklZwp0wGn9m6Nlhak2qFxz0Lp5n8tLOFgHPbKZ6hMCodh+DkbW1hq3g
DGYqruu/LAC4jhJZoaBdliJ1Vvu+EtGYZi1bBR5NELodoDrBo5ZZMgxbxBX6yAmfs/sA1bdXzxCl
r/z9V93pEocgfism7gi7Ki2FGw9BahQwvhRC5zrZFN1jvxMypQTlidWTiJ0Bx0/Rr+vY6U2KA+Ut
CE90SZg+24wiiNeW7n+zB9R2Nt2gNSRK0UOpA9hy9XBlowl4bqJzK75aVLhsVA8XZWgswDHFUvNz
OAfJSfy4Ipu0v1eAmrxqMAK0TJumQ5QTOHno3WO1PrZYhXNe/4zb5TTW+7DhMKBkxoz25jUqUlos
6fta2DeKVRwu/SpQ8RENMBvKacda2axXy+y+pgzMRV5ZIQpAbHL6mW4W+22Vnzz0dMPbQv/X9D0g
diJBjBHTHOhnf1tLRkcFHG6Rjras1gHcAeuaNfZTmIufnYfsCXPdalvoYs3dzThlclU8nuCOsiyf
qIEnHSCNGINC02ONDu4TFhK62rklpfhR9mSggPFZzhZHoql3FMxpqz3hgweYI9mgycjDl80Z8OjS
WGVaJPmzbQSk3w3qu+/f+D2ivi4mrj0mdoypV2dkvbOngvE5oLyeQRbI+vy5SiFmtWmK3k+Nt7C0
eDfoo7abJ8dReSoSed3gp12yYrnp3tjK/sKQe+MteFMeMJuJ5xn0qg//ooLqSs+c1xjvV0L/do69
UvDnDPJvXEevVKiqA4OX5gLpVUjJcf0Tc+2RDe2m0d5M2loiKjFMVoEHFP9/40bUXGg69p+5TFlJ
Uw+CiurzxxAwhGJyjd8Ap7DydLgHXUZPs7mr4niuPEK8sWVxQdthGNC0O2I7kKAK1a6W+6VgPOc/
PvtJoYjpgQbqdTyAhWs8nclwsfV8AjMoLpByB1PRPjDmCPVj44V9zpDqPhxpn1ejHJoaN+F4/SA1
BOvnmSD158PYWzsgym+oJ2wFJkx0RU8EZ7NIjTo6LzJgF3ztoNSyZYAcjfv6A5cHveTw2ezzAtM0
SQiDESl2uEG9+/EY3Fibk6mcO2mX353UaCj74EcerS97gQvv2oMgDzFUGl+3zKCQd6oJuWRCm8Z6
fDdYLvQEaXyp+gUDlmHCNfAbei3q6zoKsAC53gPJ/KcqXAjGDil+3zNlg3bEXsDNu93OeJ/Mb292
l8sHXI3mdd3/HEADi9ISYWnNhDua8NLiOvJ6EzUBPxiFMYXBGnI7zim4XUJ/LpbyupmM+4ZSMbaB
49wLTbJ1iy+vDEt4lQycctD6aye5e+cYwfG0uit0weSU6FAthh1gHp32ulQWRjTv4KK0I/+Pq9r7
M5Iu5mtcJ1zUC4UVYJpWZ0X7Ui0Tb5/Gz+qrsbsKBhOB/xe3QsmM2V5nvze+Y/7B8thuvKqUgsYX
AuIYRzwQ2giPSL1n3uyTDWg6lcbzSwqJ0BiDSt6Z2CSFq6ak1nUzV+uzZB5Ze3v3bRr0GMSCfWnm
lzwoW2CY/81Oacg383Vt9rJ1OE2sT50jPcEXzrBt0neiWVmYaWYBCsdgaiE/Vd9XsSbAULOPc+U=
`pragma protect end_protected
