 -------------------------------------------------------------------------------
-- File       : EthCrc32Pkg.vhd
-- Company    : SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------
-- Description: Ethernet CRC32 Ethernet/AAL5 Package File
-- Polynomial: x^32 + x^26 + x^23 + x^22 + x^16 + x^12 + x^11 + x^10 + x^8 + x^7 + x^5 + x^4 + x^2 + x^1 + 1
-------------------------------------------------------------------------------
-- This file is part of 'SLAC Firmware Standard Library'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'SLAC Firmware Standard Library', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

use work.StdRtlPkg.all;

package EthCrc32Pkg is

   function crc32Parallel1Byte (crcCur : slv(31 downto 0); data : slv(7 downto 0)) return slv;
   function crc32Parallel2Byte (crcCur : slv(31 downto 0); data : slv(15 downto 0)) return slv;
   function crc32Parallel3Byte (crcCur : slv(31 downto 0); data : slv(23 downto 0)) return slv;
   function crc32Parallel4Byte (crcCur : slv(31 downto 0); data : slv(31 downto 0)) return slv;
   function crc32Parallel5Byte (crcCur : slv(31 downto 0); data : slv(39 downto 0)) return slv;
   function crc32Parallel6Byte (crcCur : slv(31 downto 0); data : slv(47 downto 0)) return slv;
   function crc32Parallel7Byte (crcCur : slv(31 downto 0); data : slv(55 downto 0)) return slv;
   function crc32Parallel8Byte (crcCur : slv(31 downto 0); data : slv(63 downto 0)) return slv;
   function crc32Parallel9Byte (crcCur : slv(31 downto 0); data : slv(71 downto 0)) return slv;
   function crc32Parallel10Byte (crcCur : slv(31 downto 0); data : slv(79 downto 0)) return slv;
   function crc32Parallel11Byte (crcCur : slv(31 downto 0); data : slv(87 downto 0)) return slv;
   function crc32Parallel12Byte (crcCur : slv(31 downto 0); data : slv(95 downto 0)) return slv;
   function crc32Parallel13Byte (crcCur : slv(31 downto 0); data : slv(103 downto 0)) return slv;
   function crc32Parallel14Byte (crcCur : slv(31 downto 0); data : slv(111 downto 0)) return slv;
   function crc32Parallel15Byte (crcCur : slv(31 downto 0); data : slv(119 downto 0)) return slv;
   function crc32Parallel16Byte (crcCur : slv(31 downto 0); data : slv(127 downto 0)) return slv;

   procedure xorBitMap1Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(7 downto 0));

   procedure xorBitMap2Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(15 downto 0));

   procedure xorBitMap3Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(23 downto 0));

   procedure xorBitMap4Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(31 downto 0));

   procedure xorBitMap5Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(39 downto 0));

   procedure xorBitMap6Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(47 downto 0));

   procedure xorBitMap7Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(55 downto 0));

   procedure xorBitMap8Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(63 downto 0));

   procedure xorBitMap1Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(7 downto 0));

   procedure xorBitMap2Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(15 downto 0));

   procedure xorBitMap3Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(23 downto 0));

   procedure xorBitMap4Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(31 downto 0));

   procedure xorBitMap5Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(39 downto 0));

   procedure xorBitMap6Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(47 downto 0));

   procedure xorBitMap7Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(55 downto 0));

   procedure xorBitMap8Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(63 downto 0));

   procedure xorBitMap9Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(71 downto 0));

   procedure xorBitMap10Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(79 downto 0));

   procedure xorBitMap11Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(87 downto 0));

   procedure xorBitMap12Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(95 downto 0));

   procedure xorBitMap13Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(103 downto 0));

   procedure xorBitMap14Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(111 downto 0));

   procedure xorBitMap15Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(119 downto 0));

   procedure xorBitMap16Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(127 downto 0));

end package EthCrc32Pkg;

package body EthCrc32Pkg is

   function crc32Parallel1Byte (crcCur : slv(31 downto 0); data : slv(7 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor crcCur(24) xor crcCur(30);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor crcCur(24) xor crcCur(25) xor crcCur(30) xor crcCur(31);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor crcCur(0) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor crcCur(1) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor crcCur(2) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(29);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor crcCur(3) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor crcCur(4) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor crcCur(5) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor crcCur(6) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor crcCur(7) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(16) := data(0) xor data(4) xor data(5) xor crcCur(8) xor crcCur(24) xor crcCur(28) xor crcCur(29);
      retVar(17) := data(1) xor data(5) xor data(6) xor crcCur(9) xor crcCur(25) xor crcCur(29) xor crcCur(30);
      retVar(18) := data(2) xor data(6) xor data(7) xor crcCur(10) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(19) := data(3) xor data(7) xor crcCur(11) xor crcCur(27) xor crcCur(31);
      retVar(20) := data(4) xor crcCur(12) xor crcCur(28);
      retVar(21) := data(5) xor crcCur(13) xor crcCur(29);
      retVar(22) := data(0) xor crcCur(14) xor crcCur(24);
      retVar(23) := data(0) xor data(1) xor data(6) xor crcCur(15) xor crcCur(24) xor crcCur(25) xor crcCur(30);
      retVar(24) := data(1) xor data(2) xor data(7) xor crcCur(16) xor crcCur(25) xor crcCur(26) xor crcCur(31);
      retVar(25) := data(2) xor data(3) xor crcCur(17) xor crcCur(26) xor crcCur(27);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor crcCur(18) xor crcCur(24) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor crcCur(19) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(28) := data(2) xor data(5) xor data(6) xor crcCur(20) xor crcCur(26) xor crcCur(29) xor crcCur(30);
      retVar(29) := data(3) xor data(6) xor data(7) xor crcCur(21) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(30) := data(4) xor data(7) xor crcCur(22) xor crcCur(28) xor crcCur(31);
      retVar(31) := data(5) xor crcCur(23) xor crcCur(29);
      return retVar;
   end function;

   function crc32Parallel2Byte (crcCur : slv(31 downto 0); data : slv(15 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor crcCur(16) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(28);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor crcCur(16) xor crcCur(17) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(29) xor crcCur(30);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(26) xor crcCur(29);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(30);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(25) xor crcCur(29) xor crcCur(30);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(25) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(26) xor crcCur(29) xor crcCur(30);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(31);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor crcCur(0) xor crcCur(16) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(28) xor crcCur(29);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor crcCur(1) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(29) xor crcCur(30);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor crcCur(2) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor crcCur(3) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(31);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor crcCur(4) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(28);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor crcCur(5) xor crcCur(21) xor crcCur(25) xor crcCur(26) xor crcCur(29);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor crcCur(6) xor crcCur(16) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor crcCur(7) xor crcCur(16) xor crcCur(17) xor crcCur(22) xor crcCur(25) xor crcCur(29) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor crcCur(8) xor crcCur(17) xor crcCur(18) xor crcCur(23) xor crcCur(26) xor crcCur(30);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor crcCur(9) xor crcCur(18) xor crcCur(19) xor crcCur(24) xor crcCur(27) xor crcCur(31);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor crcCur(10) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(26);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor crcCur(11) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(27);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor crcCur(12) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(28);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor crcCur(13) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(29);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor crcCur(14) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(30);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor crcCur(15) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(31);
      return retVar;
   end function;

   function crc32Parallel3Byte (crcCur : slv(31 downto 0); data : slv(23 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor crcCur(8) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(24);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor crcCur(8) xor crcCur(9) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(25);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(18) xor crcCur(21) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(22) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(23) xor crcCur(24) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(25) xor crcCur(30) xor crcCur(31);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(26) xor crcCur(31);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(27);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(17) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(28);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(29);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(30);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(28) xor crcCur(29);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor crcCur(8) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(20) xor crcCur(21) xor crcCur(25) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(26) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(28) xor crcCur(30);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(29) xor crcCur(31);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor crcCur(13) xor crcCur(17) xor crcCur(18) xor crcCur(21) xor crcCur(25) xor crcCur(26) xor crcCur(30);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor crcCur(8) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor crcCur(8) xor crcCur(9) xor crcCur(14) xor crcCur(17) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor crcCur(0) xor crcCur(9) xor crcCur(10) xor crcCur(15) xor crcCur(18) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor crcCur(1) xor crcCur(10) xor crcCur(11) xor crcCur(16) xor crcCur(19) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor crcCur(2) xor crcCur(8) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(18) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor crcCur(3) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(19) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor crcCur(4) xor crcCur(10) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(20) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor crcCur(5) xor crcCur(11) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(21) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor crcCur(6) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(22) xor crcCur(30) xor crcCur(31);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor crcCur(7) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(23) xor crcCur(31);
      return retVar;
   end function;

   function crc32Parallel4Byte (crcCur : slv(31 downto 0); data : slv(31 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor crcCur(0) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(16) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor crcCur(0) xor crcCur(1) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(24) xor crcCur(27) xor crcCur(28);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(24) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(25) xor crcCur(27) xor crcCur(31);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(10) xor crcCur(13) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(28) xor crcCur(29);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(11) xor crcCur(14) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(29) xor crcCur(30);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(15) xor crcCur(16) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(29);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(17) xor crcCur(22) xor crcCur(23) xor crcCur(28) xor crcCur(31);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(18) xor crcCur(23) xor crcCur(24) xor crcCur(29);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(19) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(9) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(21) xor crcCur(24) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(10) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(25) xor crcCur(28) xor crcCur(31);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(11) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(26) xor crcCur(29);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(27) xor crcCur(30);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor crcCur(0) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(12) xor crcCur(13) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(29) xor crcCur(30);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor crcCur(1) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(28) xor crcCur(31);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(29);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor crcCur(5) xor crcCur(9) xor crcCur(10) xor crcCur(13) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor crcCur(0) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor crcCur(0) xor crcCur(1) xor crcCur(6) xor crcCur(9) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor crcCur(1) xor crcCur(2) xor crcCur(7) xor crcCur(10) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor crcCur(2) xor crcCur(3) xor crcCur(8) xor crcCur(11) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor crcCur(0) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(10) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(31);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor crcCur(1) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(11) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor crcCur(2) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(12) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor crcCur(3) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(13) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(14) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(15) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      return retVar;
   end function;

   function crc32Parallel5Byte (crcCur : slv(31 downto 0); data : slv(39 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(8) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(29);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor crcCur(0) xor crcCur(1) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(16) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(17) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor crcCur(0) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(30) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor crcCur(2) xor crcCur(5) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(20) xor crcCur(21) xor crcCur(29) xor crcCur(31);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor crcCur(0) xor crcCur(3) xor crcCur(6) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(30);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor crcCur(0) xor crcCur(2) xor crcCur(7) xor crcCur(8) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(26) xor crcCur(29) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(9) xor crcCur(14) xor crcCur(15) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(10) xor crcCur(15) xor crcCur(16) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor crcCur(1) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(11) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor crcCur(1) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(25) xor crcCur(28);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor crcCur(1) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(13) xor crcCur(16) xor crcCur(19) xor crcCur(22) xor crcCur(23);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor crcCur(2) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(17) xor crcCur(20) xor crcCur(23) xor crcCur(24);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor crcCur(0) xor crcCur(3) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(18) xor crcCur(21) xor crcCur(24) xor crcCur(25);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(19) xor crcCur(22) xor crcCur(25) xor crcCur(26);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor crcCur(0) xor crcCur(4) xor crcCur(5) xor crcCur(9) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(27) xor crcCur(29);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor crcCur(1) xor crcCur(5) xor crcCur(6) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(28) xor crcCur(30);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(29) xor crcCur(31);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor crcCur(0) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(30);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(31);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor crcCur(1) xor crcCur(2) xor crcCur(5) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(29);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor crcCur(1) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor crcCur(2) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor crcCur(0) xor crcCur(3) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor crcCur(2) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(23) xor crcCur(30) xor crcCur(31);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor crcCur(3) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(24) xor crcCur(31);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor crcCur(0) xor crcCur(4) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(25);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor crcCur(1) xor crcCur(5) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(26);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor crcCur(0) xor crcCur(2) xor crcCur(6) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(27);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(7) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(28);
      return retVar;
   end function;

   function crc32Parallel6Byte (crcCur : slv(31 downto 0); data : slv(47 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor crcCur(0) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(21) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor crcCur(0) xor crcCur(1) xor crcCur(8) xor crcCur(11) xor crcCur(12) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(8) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(28);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(9) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(29);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(12) xor crcCur(13) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor crcCur(0) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(18) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor crcCur(1) xor crcCur(6) xor crcCur(7) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor crcCur(2) xor crcCur(7) xor crcCur(8) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor crcCur(0) xor crcCur(3) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(26);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(17) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor crcCur(1) xor crcCur(2) xor crcCur(5) xor crcCur(8) xor crcCur(11) xor crcCur(14) xor crcCur(15) xor crcCur(25) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(9) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(10) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(27) xor crcCur(28);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor crcCur(0) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(11) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(28) xor crcCur(29);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor crcCur(1) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(19) xor crcCur(21) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor crcCur(2) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(20) xor crcCur(22) xor crcCur(29) xor crcCur(31);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(21) xor crcCur(23) xor crcCur(30);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor crcCur(0) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(22) xor crcCur(24) xor crcCur(31);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor crcCur(0) xor crcCur(1) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(23) xor crcCur(25);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor crcCur(1) xor crcCur(2) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(24) xor crcCur(26);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(31);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(28);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(15) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(31);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(16) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(29);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(17) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(19) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(20) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      return retVar;
   end function;

   function crc32Parallel7Byte (crcCur : slv(31 downto 0); data : slv(55 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(53) xor data(54) xor data(55) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(13) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(53) xor crcCur(0) xor crcCur(3) xor crcCur(4) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor data(51) xor data(52) xor data(53) xor data(55) xor crcCur(0) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(20) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor data(52) xor data(53) xor data(54) xor crcCur(1) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(21) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor data(48) xor data(50) xor crcCur(0) xor crcCur(1) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(53) xor data(54) xor data(55) xor crcCur(0) xor crcCur(4) xor crcCur(5) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(55) xor crcCur(1) xor crcCur(5) xor crcCur(6) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(10) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor data(50) xor data(51) xor data(52) xor data(54) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor data(51) xor data(52) xor data(53) xor data(55) xor crcCur(0) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor data(50) xor data(52) xor data(55) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(26) xor crcCur(28) xor crcCur(31);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(51) xor data(54) xor data(55) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(9) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor crcCur(0) xor crcCur(3) xor crcCur(6) xor crcCur(7) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor crcCur(1) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor crcCur(2) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor data(49) xor data(50) xor data(52) xor data(53) xor data(54) xor data(55) xor crcCur(0) xor crcCur(3) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(20) xor crcCur(21) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor data(48) xor data(51) xor crcCur(0) xor crcCur(2) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(11) xor crcCur(13) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(27);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor data(48) xor data(49) xor data(52) xor crcCur(1) xor crcCur(3) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(12) xor crcCur(14) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(28);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor data(48) xor data(49) xor data(50) xor data(53) xor crcCur(0) xor crcCur(2) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(13) xor crcCur(15) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(29);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor data(49) xor data(50) xor data(51) xor data(54) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(14) xor crcCur(16) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(30);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor data(48) xor data(50) xor data(51) xor data(52) xor data(55) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(15) xor crcCur(17) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor data(49) xor data(51) xor data(52) xor data(53) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(16) xor crcCur(18) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(52) xor data(55) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(28) xor crcCur(31);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(54) xor data(55) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(55) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor data(48) xor data(49) xor data(52) xor data(54) xor data(55) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(7) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor data(48) xor data(49) xor data(50) xor data(53) xor data(55) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(8) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(29) xor crcCur(31);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(54) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(9) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(30);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(55) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor data(48) xor data(51) xor data(52) xor data(53) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(11) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor data(49) xor data(52) xor data(53) xor data(54) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(12) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      return retVar;
   end function;

   function crc32Parallel8Byte (crcCur : slv(31 downto 0); data : slv(63 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(53) xor data(54) xor data(55) xor data(58) xor data(60) xor data(61) xor data(63) xor crcCur(0) xor crcCur(2) xor crcCur(5) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(53) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor data(51) xor data(52) xor data(53) xor data(55) xor data(57) xor data(58) xor data(59) xor crcCur(0) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(12) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor data(52) xor data(53) xor data(54) xor data(56) xor data(58) xor data(59) xor data(60) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(13) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor data(48) xor data(50) xor data(57) xor data(58) xor data(59) xor data(63) xor crcCur(1) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(53) xor data(54) xor data(55) xor data(59) xor data(61) xor data(63) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(55) xor data(56) xor data(60) xor data(62) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(28) xor crcCur(30);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(56) xor data(57) xor data(58) xor data(60) xor crcCur(0) xor crcCur(2) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor data(50) xor data(51) xor data(52) xor data(54) xor data(57) xor data(59) xor data(60) xor data(63) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor data(51) xor data(52) xor data(53) xor data(55) xor data(58) xor data(60) xor data(61) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(26) xor crcCur(28) xor crcCur(29);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor data(50) xor data(52) xor data(55) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(18) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(51) xor data(54) xor data(55) xor data(56) xor data(57) xor data(58) xor data(59) xor crcCur(1) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(63) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor crcCur(0) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor crcCur(0) xor crcCur(1) xor crcCur(11) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor data(49) xor data(50) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(57) xor data(59) xor data(60) xor data(62) xor crcCur(1) xor crcCur(2) xor crcCur(12) xor crcCur(13) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor data(48) xor data(51) xor data(56) xor data(57) xor crcCur(0) xor crcCur(3) xor crcCur(5) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(24) xor crcCur(25);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor data(48) xor data(49) xor data(52) xor data(57) xor data(58) xor crcCur(1) xor crcCur(4) xor crcCur(6) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(25) xor crcCur(26);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor data(48) xor data(49) xor data(50) xor data(53) xor data(58) xor data(59) xor crcCur(0) xor crcCur(2) xor crcCur(5) xor crcCur(7) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(21) xor crcCur(26) xor crcCur(27);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor data(49) xor data(50) xor data(51) xor data(54) xor data(59) xor data(60) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(6) xor crcCur(8) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(27) xor crcCur(28);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor data(48) xor data(50) xor data(51) xor data(52) xor data(55) xor data(60) xor data(61) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(7) xor crcCur(9) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(28) xor crcCur(29);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor data(49) xor data(51) xor data(52) xor data(53) xor data(56) xor data(61) xor data(62) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(8) xor crcCur(10) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(29) xor crcCur(30);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(61) xor data(62) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(20) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(54) xor data(55) xor data(56) xor data(59) xor data(60) xor data(62) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(55) xor data(56) xor data(57) xor data(60) xor data(61) xor data(63) xor crcCur(0) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(56) xor data(57) xor data(58) xor data(61) xor data(62) xor crcCur(1) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(29) xor crcCur(30);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor data(48) xor data(49) xor data(52) xor data(54) xor data(55) xor data(57) xor data(59) xor data(60) xor data(61) xor data(62) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor data(48) xor data(49) xor data(50) xor data(53) xor data(55) xor data(56) xor data(58) xor data(60) xor data(61) xor data(62) xor data(63) xor crcCur(0) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(62) xor data(63) xor crcCur(1) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(63) xor crcCur(2) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor data(48) xor data(51) xor data(52) xor data(53) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor crcCur(0) xor crcCur(3) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor data(49) xor data(52) xor data(53) xor data(54) xor data(57) xor data(59) xor data(60) xor data(62) xor crcCur(1) xor crcCur(4) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      return retVar;
   end function;

   function crc32Parallel9Byte (crcCur : slv(31 downto 0); data : slv(71 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(53) xor data(54) xor data(55) xor data(58) xor data(60) xor data(61) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(53) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(29);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor data(51) xor data(52) xor data(53) xor data(55) xor data(57) xor data(58) xor data(59) xor data(64) xor data(67) xor data(68) xor data(70) xor crcCur(4) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(24) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor data(52) xor data(53) xor data(54) xor data(56) xor data(58) xor data(59) xor data(60) xor data(65) xor data(68) xor data(69) xor data(71) xor crcCur(0) xor crcCur(5) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor data(48) xor data(50) xor data(57) xor data(58) xor data(59) xor data(63) xor data(65) xor data(67) xor data(68) xor data(69) xor data(70) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(53) xor data(54) xor data(55) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(67) xor data(69) xor data(70) xor data(71) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(55) xor data(56) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(56) xor data(57) xor data(58) xor data(60) xor data(68) xor data(69) xor data(71) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor data(50) xor data(51) xor data(52) xor data(54) xor data(57) xor data(59) xor data(60) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor data(51) xor data(52) xor data(53) xor data(55) xor data(58) xor data(60) xor data(61) xor data(64) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(71) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor data(50) xor data(52) xor data(55) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(66) xor data(69) xor data(70) xor data(71) xor crcCur(0) xor crcCur(2) xor crcCur(10) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(26) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(51) xor data(54) xor data(55) xor data(56) xor data(57) xor data(58) xor data(59) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(63) xor data(68) xor data(69) xor data(71) xor crcCur(1) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(64) xor data(69) xor data(70) xor crcCur(2) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(29) xor crcCur(30);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(65) xor data(70) xor data(71) xor crcCur(3) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(30) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor data(49) xor data(50) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(66) xor data(71) xor crcCur(4) xor crcCur(5) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(31);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor data(48) xor data(51) xor data(56) xor data(57) xor data(66) xor data(68) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(11) xor crcCur(16) xor crcCur(17) xor crcCur(26) xor crcCur(28);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor data(48) xor data(49) xor data(52) xor data(57) xor data(58) xor data(67) xor data(69) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(17) xor crcCur(18) xor crcCur(27) xor crcCur(29);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor data(48) xor data(49) xor data(50) xor data(53) xor data(58) xor data(59) xor data(68) xor data(70) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(13) xor crcCur(18) xor crcCur(19) xor crcCur(28) xor crcCur(30);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor data(49) xor data(50) xor data(51) xor data(54) xor data(59) xor data(60) xor data(69) xor data(71) xor crcCur(0) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(19) xor crcCur(20) xor crcCur(29) xor crcCur(31);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor data(48) xor data(50) xor data(51) xor data(52) xor data(55) xor data(60) xor data(61) xor data(70) xor crcCur(1) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(20) xor crcCur(21) xor crcCur(30);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor data(49) xor data(51) xor data(52) xor data(53) xor data(56) xor data(61) xor data(62) xor data(71) xor crcCur(0) xor crcCur(2) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(21) xor crcCur(22) xor crcCur(31);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(61) xor data(62) xor data(65) xor data(66) xor data(67) xor data(68) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(12) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(54) xor data(55) xor data(56) xor data(59) xor data(60) xor data(62) xor data(65) xor data(69) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(25) xor crcCur(29);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(55) xor data(56) xor data(57) xor data(60) xor data(61) xor data(63) xor data(66) xor data(70) xor crcCur(0) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(26) xor crcCur(30);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(56) xor data(57) xor data(58) xor data(61) xor data(62) xor data(64) xor data(67) xor data(71) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(27) xor crcCur(31);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor data(48) xor data(49) xor data(52) xor data(54) xor data(55) xor data(57) xor data(59) xor data(60) xor data(61) xor data(62) xor data(66) xor data(67) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(26) xor crcCur(27);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor data(48) xor data(49) xor data(50) xor data(53) xor data(55) xor data(56) xor data(58) xor data(60) xor data(61) xor data(62) xor data(63) xor data(67) xor data(68) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(27) xor crcCur(28);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(62) xor data(63) xor data(64) xor data(68) xor data(69) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(28) xor crcCur(29);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(70) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(29) xor crcCur(30);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor data(48) xor data(51) xor data(52) xor data(53) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(66) xor data(70) xor data(71) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor data(49) xor data(52) xor data(53) xor data(54) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(67) xor data(71) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      return retVar;
   end function;

   function crc32Parallel10Byte (crcCur : slv(31 downto 0); data : slv(79 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(53) xor data(54) xor data(55) xor data(58) xor data(60) xor data(61) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(72) xor data(73) xor data(79) xor crcCur(0) xor crcCur(2) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(53) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(72) xor data(74) xor data(79) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(21) xor crcCur(24) xor crcCur(26) xor crcCur(31);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor data(51) xor data(52) xor data(53) xor data(55) xor data(57) xor data(58) xor data(59) xor data(64) xor data(67) xor data(68) xor data(70) xor data(72) xor data(75) xor data(79) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(27) xor crcCur(31);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor data(52) xor data(53) xor data(54) xor data(56) xor data(58) xor data(59) xor data(60) xor data(65) xor data(68) xor data(69) xor data(71) xor data(73) xor data(76) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(28);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor data(48) xor data(50) xor data(57) xor data(58) xor data(59) xor data(63) xor data(65) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(74) xor data(77) xor data(79) xor crcCur(0) xor crcCur(2) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(29) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(53) xor data(54) xor data(55) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(67) xor data(69) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(78) xor data(79) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(55) xor data(56) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(76) xor data(79) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(56) xor data(57) xor data(58) xor data(60) xor data(68) xor data(69) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(79) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor data(50) xor data(51) xor data(52) xor data(54) xor data(57) xor data(59) xor data(60) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor data(51) xor data(52) xor data(53) xor data(55) xor data(58) xor data(60) xor data(61) xor data(64) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(71) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor data(50) xor data(52) xor data(55) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(66) xor data(69) xor data(70) xor data(71) xor data(73) xor data(75) xor data(77) xor data(78) xor crcCur(2) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(51) xor data(54) xor data(55) xor data(56) xor data(57) xor data(58) xor data(59) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(73) xor data(74) xor data(76) xor data(78) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(63) xor data(68) xor data(69) xor data(71) xor data(73) xor data(74) xor data(75) xor data(77) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(64) xor data(69) xor data(70) xor data(72) xor data(74) xor data(75) xor data(76) xor data(78) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(65) xor data(70) xor data(71) xor data(73) xor data(75) xor data(76) xor data(77) xor data(79) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor data(49) xor data(50) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(66) xor data(71) xor data(72) xor data(74) xor data(76) xor data(77) xor data(78) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor data(48) xor data(51) xor data(56) xor data(57) xor data(66) xor data(68) xor data(75) xor data(77) xor data(78) xor crcCur(0) xor crcCur(3) xor crcCur(8) xor crcCur(9) xor crcCur(18) xor crcCur(20) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor data(48) xor data(49) xor data(52) xor data(57) xor data(58) xor data(67) xor data(69) xor data(76) xor data(78) xor data(79) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(9) xor crcCur(10) xor crcCur(19) xor crcCur(21) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor data(48) xor data(49) xor data(50) xor data(53) xor data(58) xor data(59) xor data(68) xor data(70) xor data(77) xor data(79) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(5) xor crcCur(10) xor crcCur(11) xor crcCur(20) xor crcCur(22) xor crcCur(29) xor crcCur(31);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor data(49) xor data(50) xor data(51) xor data(54) xor data(59) xor data(60) xor data(69) xor data(71) xor data(78) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(11) xor crcCur(12) xor crcCur(21) xor crcCur(23) xor crcCur(30);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor data(48) xor data(50) xor data(51) xor data(52) xor data(55) xor data(60) xor data(61) xor data(70) xor data(72) xor data(79) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(12) xor crcCur(13) xor crcCur(22) xor crcCur(24) xor crcCur(31);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor data(49) xor data(51) xor data(52) xor data(53) xor data(56) xor data(61) xor data(62) xor data(71) xor data(73) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(13) xor crcCur(14) xor crcCur(23) xor crcCur(25);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(61) xor data(62) xor data(65) xor data(66) xor data(67) xor data(68) xor data(73) xor data(74) xor data(79) xor crcCur(0) xor crcCur(4) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(25) xor crcCur(26) xor crcCur(31);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(54) xor data(55) xor data(56) xor data(59) xor data(60) xor data(62) xor data(65) xor data(69) xor data(72) xor data(73) xor data(74) xor data(75) xor data(79) xor crcCur(1) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(17) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(55) xor data(56) xor data(57) xor data(60) xor data(61) xor data(63) xor data(66) xor data(70) xor data(73) xor data(74) xor data(75) xor data(76) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(56) xor data(57) xor data(58) xor data(61) xor data(62) xor data(64) xor data(67) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(19) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor data(48) xor data(49) xor data(52) xor data(54) xor data(55) xor data(57) xor data(59) xor data(60) xor data(61) xor data(62) xor data(66) xor data(67) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(18) xor crcCur(19) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor data(48) xor data(49) xor data(50) xor data(53) xor data(55) xor data(56) xor data(58) xor data(60) xor data(61) xor data(62) xor data(63) xor data(67) xor data(68) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(19) xor crcCur(20) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(62) xor data(63) xor data(64) xor data(68) xor data(69) xor data(75) xor data(77) xor data(78) xor data(79) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(20) xor crcCur(21) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(70) xor data(76) xor data(78) xor data(79) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor data(48) xor data(51) xor data(52) xor data(53) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(66) xor data(70) xor data(71) xor data(77) xor data(79) xor crcCur(0) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(29) xor crcCur(31);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor data(49) xor data(52) xor data(53) xor data(54) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(67) xor data(71) xor data(72) xor data(78) xor crcCur(1) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(30);
      return retVar;
   end function;

   function crc32Parallel11Byte (crcCur : slv(31 downto 0); data : slv(87 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(53) xor data(54) xor data(55) xor data(58) xor data(60) xor data(61) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(72) xor data(73) xor data(79) xor data(81) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(53) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(72) xor data(74) xor data(79) xor data(80) xor data(81) xor data(86) xor data(87) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(13) xor crcCur(16) xor crcCur(18) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(30) xor crcCur(31);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor data(51) xor data(52) xor data(53) xor data(55) xor data(57) xor data(58) xor data(59) xor data(64) xor data(67) xor data(68) xor data(70) xor data(72) xor data(75) xor data(79) xor data(80) xor data(83) xor data(84) xor data(85) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(8) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor data(52) xor data(53) xor data(54) xor data(56) xor data(58) xor data(59) xor data(60) xor data(65) xor data(68) xor data(69) xor data(71) xor data(73) xor data(76) xor data(80) xor data(81) xor data(84) xor data(85) xor data(86) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor data(48) xor data(50) xor data(57) xor data(58) xor data(59) xor data(63) xor data(65) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(74) xor data(77) xor data(79) xor data(83) xor data(84) xor data(86) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(21) xor crcCur(23) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(53) xor data(54) xor data(55) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(67) xor data(69) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(55) xor data(56) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(76) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor crcCur(0) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(56) xor data(57) xor data(58) xor data(60) xor data(68) xor data(69) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(79) xor data(80) xor data(87) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor data(50) xor data(51) xor data(52) xor data(54) xor data(57) xor data(59) xor data(60) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor data(51) xor data(52) xor data(53) xor data(55) xor data(58) xor data(60) xor data(61) xor data(64) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(71) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(84) xor data(85) xor data(86) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor data(50) xor data(52) xor data(55) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(66) xor data(69) xor data(70) xor data(71) xor data(73) xor data(75) xor data(77) xor data(78) xor data(80) xor data(83) xor data(86) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(10) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(27) xor crcCur(30);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(51) xor data(54) xor data(55) xor data(56) xor data(57) xor data(58) xor data(59) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(73) xor data(74) xor data(76) xor data(78) xor data(82) xor data(83) xor data(85) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(26) xor crcCur(27) xor crcCur(29);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(63) xor data(68) xor data(69) xor data(71) xor data(73) xor data(74) xor data(75) xor data(77) xor data(81) xor data(82) xor data(85) xor data(86) xor data(87) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(25) xor crcCur(26) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(64) xor data(69) xor data(70) xor data(72) xor data(74) xor data(75) xor data(76) xor data(78) xor data(82) xor data(83) xor data(86) xor data(87) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(26) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(65) xor data(70) xor data(71) xor data(73) xor data(75) xor data(76) xor data(77) xor data(79) xor data(83) xor data(84) xor data(87) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor data(49) xor data(50) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(66) xor data(71) xor data(72) xor data(74) xor data(76) xor data(77) xor data(78) xor data(80) xor data(84) xor data(85) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(28) xor crcCur(29);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor data(48) xor data(51) xor data(56) xor data(57) xor data(66) xor data(68) xor data(75) xor data(77) xor data(78) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor crcCur(0) xor crcCur(1) xor crcCur(10) xor crcCur(12) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor data(48) xor data(49) xor data(52) xor data(57) xor data(58) xor data(67) xor data(69) xor data(76) xor data(78) xor data(79) xor data(83) xor data(84) xor data(85) xor data(87) xor crcCur(1) xor crcCur(2) xor crcCur(11) xor crcCur(13) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor data(48) xor data(49) xor data(50) xor data(53) xor data(58) xor data(59) xor data(68) xor data(70) xor data(77) xor data(79) xor data(80) xor data(84) xor data(85) xor data(86) xor crcCur(2) xor crcCur(3) xor crcCur(12) xor crcCur(14) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor data(49) xor data(50) xor data(51) xor data(54) xor data(59) xor data(60) xor data(69) xor data(71) xor data(78) xor data(80) xor data(81) xor data(85) xor data(86) xor data(87) xor crcCur(3) xor crcCur(4) xor crcCur(13) xor crcCur(15) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor data(48) xor data(50) xor data(51) xor data(52) xor data(55) xor data(60) xor data(61) xor data(70) xor data(72) xor data(79) xor data(81) xor data(82) xor data(86) xor data(87) xor crcCur(4) xor crcCur(5) xor crcCur(14) xor crcCur(16) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor data(49) xor data(51) xor data(52) xor data(53) xor data(56) xor data(61) xor data(62) xor data(71) xor data(73) xor data(80) xor data(82) xor data(83) xor data(87) xor crcCur(0) xor crcCur(5) xor crcCur(6) xor crcCur(15) xor crcCur(17) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(61) xor data(62) xor data(65) xor data(66) xor data(67) xor data(68) xor data(73) xor data(74) xor data(79) xor data(82) xor data(85) xor data(87) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(17) xor crcCur(18) xor crcCur(23) xor crcCur(26) xor crcCur(29) xor crcCur(31);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(54) xor data(55) xor data(56) xor data(59) xor data(60) xor data(62) xor data(65) xor data(69) xor data(72) xor data(73) xor data(74) xor data(75) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(85) xor data(86) xor data(87) xor crcCur(0) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(9) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(55) xor data(56) xor data(57) xor data(60) xor data(61) xor data(63) xor data(66) xor data(70) xor data(73) xor data(74) xor data(75) xor data(76) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(86) xor data(87) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(56) xor data(57) xor data(58) xor data(61) xor data(62) xor data(64) xor data(67) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(11) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor data(48) xor data(49) xor data(52) xor data(54) xor data(55) xor data(57) xor data(59) xor data(60) xor data(61) xor data(62) xor data(66) xor data(67) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(81) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(10) xor crcCur(11) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(25);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor data(48) xor data(49) xor data(50) xor data(53) xor data(55) xor data(56) xor data(58) xor data(60) xor data(61) xor data(62) xor data(63) xor data(67) xor data(68) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor crcCur(0) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(11) xor crcCur(12) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(62) xor data(63) xor data(64) xor data(68) xor data(69) xor data(75) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(12) xor crcCur(13) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(70) xor data(76) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor data(48) xor data(51) xor data(52) xor data(53) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(66) xor data(70) xor data(71) xor data(77) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor data(49) xor data(52) xor data(53) xor data(54) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(67) xor data(71) xor data(72) xor data(78) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      return retVar;
   end function;

   function crc32Parallel12Byte (crcCur : slv(31 downto 0); data : slv(95 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(53) xor data(54) xor data(55) xor data(58) xor data(60) xor data(61) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(72) xor data(73) xor data(79) xor data(81) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor data(94) xor data(95) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(30) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(53) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(72) xor data(74) xor data(79) xor data(80) xor data(81) xor data(86) xor data(87) xor data(88) xor data(94) xor crcCur(0) xor crcCur(1) xor crcCur(5) xor crcCur(8) xor crcCur(10) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(30);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor data(51) xor data(52) xor data(53) xor data(55) xor data(57) xor data(58) xor data(59) xor data(64) xor data(67) xor data(68) xor data(70) xor data(72) xor data(75) xor data(79) xor data(80) xor data(83) xor data(84) xor data(85) xor data(88) xor data(89) xor data(94) xor crcCur(0) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(30);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor data(52) xor data(53) xor data(54) xor data(56) xor data(58) xor data(59) xor data(60) xor data(65) xor data(68) xor data(69) xor data(71) xor data(73) xor data(76) xor data(80) xor data(81) xor data(84) xor data(85) xor data(86) xor data(89) xor data(90) xor data(95) xor crcCur(1) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(31);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor data(48) xor data(50) xor data(57) xor data(58) xor data(59) xor data(63) xor data(65) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(74) xor data(77) xor data(79) xor data(83) xor data(84) xor data(86) xor data(90) xor data(91) xor data(94) xor data(95) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(13) xor crcCur(15) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(26) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(53) xor data(54) xor data(55) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(67) xor data(69) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(91) xor data(92) xor data(94) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(55) xor data(56) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(76) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(92) xor data(93) xor data(95) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(56) xor data(57) xor data(58) xor data(60) xor data(68) xor data(69) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(79) xor data(80) xor data(87) xor data(93) xor data(95) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(23) xor crcCur(29) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor data(50) xor data(51) xor data(52) xor data(54) xor data(57) xor data(59) xor data(60) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor data(88) xor data(95) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(31);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor data(51) xor data(52) xor data(53) xor data(55) xor data(58) xor data(60) xor data(61) xor data(64) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(71) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(84) xor data(85) xor data(86) xor data(88) xor data(89) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor data(50) xor data(52) xor data(55) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(66) xor data(69) xor data(70) xor data(71) xor data(73) xor data(75) xor data(77) xor data(78) xor data(80) xor data(83) xor data(86) xor data(89) xor data(90) xor data(94) xor data(95) xor crcCur(2) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(19) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(51) xor data(54) xor data(55) xor data(56) xor data(57) xor data(58) xor data(59) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(73) xor data(74) xor data(76) xor data(78) xor data(82) xor data(83) xor data(85) xor data(90) xor data(91) xor data(94) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(26) xor crcCur(27) xor crcCur(30);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(63) xor data(68) xor data(69) xor data(71) xor data(73) xor data(74) xor data(75) xor data(77) xor data(81) xor data(82) xor data(85) xor data(86) xor data(87) xor data(91) xor data(92) xor data(94) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(17) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(64) xor data(69) xor data(70) xor data(72) xor data(74) xor data(75) xor data(76) xor data(78) xor data(82) xor data(83) xor data(86) xor data(87) xor data(88) xor data(92) xor data(93) xor data(95) xor crcCur(0) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(65) xor data(70) xor data(71) xor data(73) xor data(75) xor data(76) xor data(77) xor data(79) xor data(83) xor data(84) xor data(87) xor data(88) xor data(89) xor data(93) xor data(94) xor crcCur(1) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(29) xor crcCur(30);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor data(49) xor data(50) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(66) xor data(71) xor data(72) xor data(74) xor data(76) xor data(77) xor data(78) xor data(80) xor data(84) xor data(85) xor data(88) xor data(89) xor data(90) xor data(94) xor data(95) xor crcCur(0) xor crcCur(2) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor data(48) xor data(51) xor data(56) xor data(57) xor data(66) xor data(68) xor data(75) xor data(77) xor data(78) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor data(89) xor data(90) xor data(91) xor data(94) xor crcCur(2) xor crcCur(4) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(30);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor data(48) xor data(49) xor data(52) xor data(57) xor data(58) xor data(67) xor data(69) xor data(76) xor data(78) xor data(79) xor data(83) xor data(84) xor data(85) xor data(87) xor data(88) xor data(90) xor data(91) xor data(92) xor data(95) xor crcCur(3) xor crcCur(5) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor data(48) xor data(49) xor data(50) xor data(53) xor data(58) xor data(59) xor data(68) xor data(70) xor data(77) xor data(79) xor data(80) xor data(84) xor data(85) xor data(86) xor data(88) xor data(89) xor data(91) xor data(92) xor data(93) xor crcCur(4) xor crcCur(6) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor data(49) xor data(50) xor data(51) xor data(54) xor data(59) xor data(60) xor data(69) xor data(71) xor data(78) xor data(80) xor data(81) xor data(85) xor data(86) xor data(87) xor data(89) xor data(90) xor data(92) xor data(93) xor data(94) xor crcCur(5) xor crcCur(7) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor data(48) xor data(50) xor data(51) xor data(52) xor data(55) xor data(60) xor data(61) xor data(70) xor data(72) xor data(79) xor data(81) xor data(82) xor data(86) xor data(87) xor data(88) xor data(90) xor data(91) xor data(93) xor data(94) xor data(95) xor crcCur(6) xor crcCur(8) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor data(49) xor data(51) xor data(52) xor data(53) xor data(56) xor data(61) xor data(62) xor data(71) xor data(73) xor data(80) xor data(82) xor data(83) xor data(87) xor data(88) xor data(89) xor data(91) xor data(92) xor data(94) xor data(95) xor crcCur(7) xor crcCur(9) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(61) xor data(62) xor data(65) xor data(66) xor data(67) xor data(68) xor data(73) xor data(74) xor data(79) xor data(82) xor data(85) xor data(87) xor data(88) xor data(89) xor data(90) xor data(92) xor data(93) xor data(94) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(9) xor crcCur(10) xor crcCur(15) xor crcCur(18) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(54) xor data(55) xor data(56) xor data(59) xor data(60) xor data(62) xor data(65) xor data(69) xor data(72) xor data(73) xor data(74) xor data(75) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(85) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(93) xor crcCur(1) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(55) xor data(56) xor data(57) xor data(60) xor data(61) xor data(63) xor data(66) xor data(70) xor data(73) xor data(74) xor data(75) xor data(76) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(94) xor crcCur(2) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(56) xor data(57) xor data(58) xor data(61) xor data(62) xor data(64) xor data(67) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(95) xor crcCur(0) xor crcCur(3) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor data(48) xor data(49) xor data(52) xor data(54) xor data(55) xor data(57) xor data(59) xor data(60) xor data(61) xor data(62) xor data(66) xor data(67) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(81) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(95) xor crcCur(2) xor crcCur(3) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor data(48) xor data(49) xor data(50) xor data(53) xor data(55) xor data(56) xor data(58) xor data(60) xor data(61) xor data(62) xor data(63) xor data(67) xor data(68) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(94) xor crcCur(3) xor crcCur(4) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(62) xor data(63) xor data(64) xor data(68) xor data(69) xor data(75) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(90) xor data(91) xor data(92) xor data(93) xor data(94) xor data(95) xor crcCur(0) xor crcCur(4) xor crcCur(5) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(70) xor data(76) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(91) xor data(92) xor data(93) xor data(94) xor data(95) xor crcCur(0) xor crcCur(1) xor crcCur(5) xor crcCur(6) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor data(48) xor data(51) xor data(52) xor data(53) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(66) xor data(70) xor data(71) xor data(77) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(92) xor data(93) xor data(94) xor data(95) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor data(49) xor data(52) xor data(53) xor data(54) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(67) xor data(71) xor data(72) xor data(78) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(93) xor data(94) xor data(95) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      return retVar;
   end function;

   function crc32Parallel13Byte (crcCur : slv(31 downto 0); data : slv(103 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(53) xor data(54) xor data(55) xor data(58) xor data(60) xor data(61) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(72) xor data(73) xor data(79) xor data(81) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor data(94) xor data(95) xor data(96) xor data(97) xor data(98) xor data(99) xor data(101) xor data(103) xor crcCur(0) xor crcCur(1) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(53) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(72) xor data(74) xor data(79) xor data(80) xor data(81) xor data(86) xor data(87) xor data(88) xor data(94) xor data(100) xor data(101) xor data(102) xor data(103) xor crcCur(0) xor crcCur(2) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(22) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor data(51) xor data(52) xor data(53) xor data(55) xor data(57) xor data(58) xor data(59) xor data(64) xor data(67) xor data(68) xor data(70) xor data(72) xor data(75) xor data(79) xor data(80) xor data(83) xor data(84) xor data(85) xor data(88) xor data(89) xor data(94) xor data(96) xor data(97) xor data(98) xor data(99) xor data(102) xor crcCur(0) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(30);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor data(52) xor data(53) xor data(54) xor data(56) xor data(58) xor data(59) xor data(60) xor data(65) xor data(68) xor data(69) xor data(71) xor data(73) xor data(76) xor data(80) xor data(81) xor data(84) xor data(85) xor data(86) xor data(89) xor data(90) xor data(95) xor data(97) xor data(98) xor data(99) xor data(100) xor data(103) xor crcCur(1) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor data(48) xor data(50) xor data(57) xor data(58) xor data(59) xor data(63) xor data(65) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(74) xor data(77) xor data(79) xor data(83) xor data(84) xor data(86) xor data(90) xor data(91) xor data(94) xor data(95) xor data(97) xor data(100) xor data(103) xor crcCur(1) xor crcCur(2) xor crcCur(5) xor crcCur(7) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(28) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(53) xor data(54) xor data(55) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(67) xor data(69) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(91) xor data(92) xor data(94) xor data(97) xor data(99) xor data(103) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(25) xor crcCur(27) xor crcCur(31);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(55) xor data(56) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(76) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(92) xor data(93) xor data(95) xor data(98) xor data(100) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(26) xor crcCur(28);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(56) xor data(57) xor data(58) xor data(60) xor data(68) xor data(69) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(79) xor data(80) xor data(87) xor data(93) xor data(95) xor data(97) xor data(98) xor data(103) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(15) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor data(50) xor data(51) xor data(52) xor data(54) xor data(57) xor data(59) xor data(60) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor data(88) xor data(95) xor data(97) xor data(101) xor data(103) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(23) xor crcCur(25) xor crcCur(29) xor crcCur(31);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor data(51) xor data(52) xor data(53) xor data(55) xor data(58) xor data(60) xor data(61) xor data(64) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(71) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(84) xor data(85) xor data(86) xor data(88) xor data(89) xor data(96) xor data(98) xor data(102) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(24) xor crcCur(26) xor crcCur(30);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor data(50) xor data(52) xor data(55) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(66) xor data(69) xor data(70) xor data(71) xor data(73) xor data(75) xor data(77) xor data(78) xor data(80) xor data(83) xor data(86) xor data(89) xor data(90) xor data(94) xor data(95) xor data(96) xor data(98) xor data(101) xor crcCur(1) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(11) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(29);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(51) xor data(54) xor data(55) xor data(56) xor data(57) xor data(58) xor data(59) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(73) xor data(74) xor data(76) xor data(78) xor data(82) xor data(83) xor data(85) xor data(90) xor data(91) xor data(94) xor data(98) xor data(101) xor data(102) xor data(103) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(6) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(26) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(63) xor data(68) xor data(69) xor data(71) xor data(73) xor data(74) xor data(75) xor data(77) xor data(81) xor data(82) xor data(85) xor data(86) xor data(87) xor data(91) xor data(92) xor data(94) xor data(96) xor data(97) xor data(98) xor data(101) xor data(102) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(9) xor crcCur(10) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(29) xor crcCur(30);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(64) xor data(69) xor data(70) xor data(72) xor data(74) xor data(75) xor data(76) xor data(78) xor data(82) xor data(83) xor data(86) xor data(87) xor data(88) xor data(92) xor data(93) xor data(95) xor data(97) xor data(98) xor data(99) xor data(102) xor data(103) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(65) xor data(70) xor data(71) xor data(73) xor data(75) xor data(76) xor data(77) xor data(79) xor data(83) xor data(84) xor data(87) xor data(88) xor data(89) xor data(93) xor data(94) xor data(96) xor data(98) xor data(99) xor data(100) xor data(103) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor data(49) xor data(50) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(66) xor data(71) xor data(72) xor data(74) xor data(76) xor data(77) xor data(78) xor data(80) xor data(84) xor data(85) xor data(88) xor data(89) xor data(90) xor data(94) xor data(95) xor data(97) xor data(99) xor data(100) xor data(101) xor crcCur(0) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor data(48) xor data(51) xor data(56) xor data(57) xor data(66) xor data(68) xor data(75) xor data(77) xor data(78) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor data(89) xor data(90) xor data(91) xor data(94) xor data(97) xor data(99) xor data(100) xor data(102) xor data(103) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor data(48) xor data(49) xor data(52) xor data(57) xor data(58) xor data(67) xor data(69) xor data(76) xor data(78) xor data(79) xor data(83) xor data(84) xor data(85) xor data(87) xor data(88) xor data(90) xor data(91) xor data(92) xor data(95) xor data(98) xor data(100) xor data(101) xor data(103) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor data(48) xor data(49) xor data(50) xor data(53) xor data(58) xor data(59) xor data(68) xor data(70) xor data(77) xor data(79) xor data(80) xor data(84) xor data(85) xor data(86) xor data(88) xor data(89) xor data(91) xor data(92) xor data(93) xor data(96) xor data(99) xor data(101) xor data(102) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor data(49) xor data(50) xor data(51) xor data(54) xor data(59) xor data(60) xor data(69) xor data(71) xor data(78) xor data(80) xor data(81) xor data(85) xor data(86) xor data(87) xor data(89) xor data(90) xor data(92) xor data(93) xor data(94) xor data(97) xor data(100) xor data(102) xor data(103) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor data(48) xor data(50) xor data(51) xor data(52) xor data(55) xor data(60) xor data(61) xor data(70) xor data(72) xor data(79) xor data(81) xor data(82) xor data(86) xor data(87) xor data(88) xor data(90) xor data(91) xor data(93) xor data(94) xor data(95) xor data(98) xor data(101) xor data(103) xor crcCur(0) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(26) xor crcCur(29) xor crcCur(31);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor data(49) xor data(51) xor data(52) xor data(53) xor data(56) xor data(61) xor data(62) xor data(71) xor data(73) xor data(80) xor data(82) xor data(83) xor data(87) xor data(88) xor data(89) xor data(91) xor data(92) xor data(94) xor data(95) xor data(96) xor data(99) xor data(102) xor crcCur(1) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(30);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(61) xor data(62) xor data(65) xor data(66) xor data(67) xor data(68) xor data(73) xor data(74) xor data(79) xor data(82) xor data(85) xor data(87) xor data(88) xor data(89) xor data(90) xor data(92) xor data(93) xor data(94) xor data(98) xor data(99) xor data(100) xor data(101) xor crcCur(1) xor crcCur(2) xor crcCur(7) xor crcCur(10) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(54) xor data(55) xor data(56) xor data(59) xor data(60) xor data(62) xor data(65) xor data(69) xor data(72) xor data(73) xor data(74) xor data(75) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(85) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(93) xor data(96) xor data(97) xor data(98) xor data(100) xor data(102) xor data(103) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(55) xor data(56) xor data(57) xor data(60) xor data(61) xor data(63) xor data(66) xor data(70) xor data(73) xor data(74) xor data(75) xor data(76) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(94) xor data(97) xor data(98) xor data(99) xor data(101) xor data(103) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(56) xor data(57) xor data(58) xor data(61) xor data(62) xor data(64) xor data(67) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(95) xor data(98) xor data(99) xor data(100) xor data(102) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor data(48) xor data(49) xor data(52) xor data(54) xor data(55) xor data(57) xor data(59) xor data(60) xor data(61) xor data(62) xor data(66) xor data(67) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(81) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(95) xor data(97) xor data(98) xor data(100) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(28);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor data(48) xor data(49) xor data(50) xor data(53) xor data(55) xor data(56) xor data(58) xor data(60) xor data(61) xor data(62) xor data(63) xor data(67) xor data(68) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(94) xor data(96) xor data(98) xor data(99) xor data(101) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(29);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(62) xor data(63) xor data(64) xor data(68) xor data(69) xor data(75) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(90) xor data(91) xor data(92) xor data(93) xor data(94) xor data(95) xor data(97) xor data(99) xor data(100) xor data(102) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(70) xor data(76) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(91) xor data(92) xor data(93) xor data(94) xor data(95) xor data(96) xor data(98) xor data(100) xor data(101) xor data(103) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor data(48) xor data(51) xor data(52) xor data(53) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(66) xor data(70) xor data(71) xor data(77) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(92) xor data(93) xor data(94) xor data(95) xor data(96) xor data(97) xor data(99) xor data(101) xor data(102) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor data(49) xor data(52) xor data(53) xor data(54) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(67) xor data(71) xor data(72) xor data(78) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(93) xor data(94) xor data(95) xor data(96) xor data(97) xor data(98) xor data(100) xor data(102) xor data(103) xor crcCur(0) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      return retVar;
   end function;

   function crc32Parallel14Byte (crcCur : slv(31 downto 0); data : slv(111 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(53) xor data(54) xor data(55) xor data(58) xor data(60) xor data(61) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(72) xor data(73) xor data(79) xor data(81) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor data(94) xor data(95) xor data(96) xor data(97) xor data(98) xor data(99) xor data(101) xor data(103) xor data(104) xor data(106) xor data(110) xor data(111) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(53) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(72) xor data(74) xor data(79) xor data(80) xor data(81) xor data(86) xor data(87) xor data(88) xor data(94) xor data(100) xor data(101) xor data(102) xor data(103) xor data(105) xor data(106) xor data(107) xor data(110) xor crcCur(0) xor crcCur(1) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(14) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(30);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor data(51) xor data(52) xor data(53) xor data(55) xor data(57) xor data(58) xor data(59) xor data(64) xor data(67) xor data(68) xor data(70) xor data(72) xor data(75) xor data(79) xor data(80) xor data(83) xor data(84) xor data(85) xor data(88) xor data(89) xor data(94) xor data(96) xor data(97) xor data(98) xor data(99) xor data(102) xor data(107) xor data(108) xor data(110) xor crcCur(0) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(27) xor crcCur(28) xor crcCur(30);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor data(52) xor data(53) xor data(54) xor data(56) xor data(58) xor data(59) xor data(60) xor data(65) xor data(68) xor data(69) xor data(71) xor data(73) xor data(76) xor data(80) xor data(81) xor data(84) xor data(85) xor data(86) xor data(89) xor data(90) xor data(95) xor data(97) xor data(98) xor data(99) xor data(100) xor data(103) xor data(108) xor data(109) xor data(111) xor crcCur(0) xor crcCur(1) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor data(48) xor data(50) xor data(57) xor data(58) xor data(59) xor data(63) xor data(65) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(74) xor data(77) xor data(79) xor data(83) xor data(84) xor data(86) xor data(90) xor data(91) xor data(94) xor data(95) xor data(97) xor data(100) xor data(103) xor data(106) xor data(109) xor data(111) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(20) xor crcCur(23) xor crcCur(26) xor crcCur(29) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(53) xor data(54) xor data(55) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(67) xor data(69) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(91) xor data(92) xor data(94) xor data(97) xor data(99) xor data(103) xor data(106) xor data(107) xor data(111) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(17) xor crcCur(19) xor crcCur(23) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(55) xor data(56) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(76) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(92) xor data(93) xor data(95) xor data(98) xor data(100) xor data(104) xor data(107) xor data(108) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(20) xor crcCur(24) xor crcCur(27) xor crcCur(28);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(56) xor data(57) xor data(58) xor data(60) xor data(68) xor data(69) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(79) xor data(80) xor data(87) xor data(93) xor data(95) xor data(97) xor data(98) xor data(103) xor data(104) xor data(105) xor data(106) xor data(108) xor data(109) xor data(110) xor data(111) xor crcCur(0) xor crcCur(7) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor data(50) xor data(51) xor data(52) xor data(54) xor data(57) xor data(59) xor data(60) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor data(88) xor data(95) xor data(97) xor data(101) xor data(103) xor data(105) xor data(107) xor data(109) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(15) xor crcCur(17) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(29);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor data(51) xor data(52) xor data(53) xor data(55) xor data(58) xor data(60) xor data(61) xor data(64) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(71) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(84) xor data(85) xor data(86) xor data(88) xor data(89) xor data(96) xor data(98) xor data(102) xor data(104) xor data(106) xor data(108) xor data(110) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(16) xor crcCur(18) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(28) xor crcCur(30);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor data(50) xor data(52) xor data(55) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(66) xor data(69) xor data(70) xor data(71) xor data(73) xor data(75) xor data(77) xor data(78) xor data(80) xor data(83) xor data(86) xor data(89) xor data(90) xor data(94) xor data(95) xor data(96) xor data(98) xor data(101) xor data(104) xor data(105) xor data(106) xor data(107) xor data(109) xor data(110) xor crcCur(0) xor crcCur(3) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(51) xor data(54) xor data(55) xor data(56) xor data(57) xor data(58) xor data(59) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(73) xor data(74) xor data(76) xor data(78) xor data(82) xor data(83) xor data(85) xor data(90) xor data(91) xor data(94) xor data(98) xor data(101) xor data(102) xor data(103) xor data(104) xor data(105) xor data(107) xor data(108) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(63) xor data(68) xor data(69) xor data(71) xor data(73) xor data(74) xor data(75) xor data(77) xor data(81) xor data(82) xor data(85) xor data(86) xor data(87) xor data(91) xor data(92) xor data(94) xor data(96) xor data(97) xor data(98) xor data(101) xor data(102) xor data(105) xor data(108) xor data(109) xor data(110) xor data(111) xor crcCur(1) xor crcCur(2) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(64) xor data(69) xor data(70) xor data(72) xor data(74) xor data(75) xor data(76) xor data(78) xor data(82) xor data(83) xor data(86) xor data(87) xor data(88) xor data(92) xor data(93) xor data(95) xor data(97) xor data(98) xor data(99) xor data(102) xor data(103) xor data(106) xor data(109) xor data(110) xor data(111) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(26) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(65) xor data(70) xor data(71) xor data(73) xor data(75) xor data(76) xor data(77) xor data(79) xor data(83) xor data(84) xor data(87) xor data(88) xor data(89) xor data(93) xor data(94) xor data(96) xor data(98) xor data(99) xor data(100) xor data(103) xor data(104) xor data(107) xor data(110) xor data(111) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor data(49) xor data(50) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(66) xor data(71) xor data(72) xor data(74) xor data(76) xor data(77) xor data(78) xor data(80) xor data(84) xor data(85) xor data(88) xor data(89) xor data(90) xor data(94) xor data(95) xor data(97) xor data(99) xor data(100) xor data(101) xor data(104) xor data(105) xor data(108) xor data(111) xor crcCur(0) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(31);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor data(48) xor data(51) xor data(56) xor data(57) xor data(66) xor data(68) xor data(75) xor data(77) xor data(78) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor data(89) xor data(90) xor data(91) xor data(94) xor data(97) xor data(99) xor data(100) xor data(102) xor data(103) xor data(104) xor data(105) xor data(109) xor data(110) xor data(111) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor data(48) xor data(49) xor data(52) xor data(57) xor data(58) xor data(67) xor data(69) xor data(76) xor data(78) xor data(79) xor data(83) xor data(84) xor data(85) xor data(87) xor data(88) xor data(90) xor data(91) xor data(92) xor data(95) xor data(98) xor data(100) xor data(101) xor data(103) xor data(104) xor data(105) xor data(106) xor data(110) xor data(111) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(30) xor crcCur(31);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor data(48) xor data(49) xor data(50) xor data(53) xor data(58) xor data(59) xor data(68) xor data(70) xor data(77) xor data(79) xor data(80) xor data(84) xor data(85) xor data(86) xor data(88) xor data(89) xor data(91) xor data(92) xor data(93) xor data(96) xor data(99) xor data(101) xor data(102) xor data(104) xor data(105) xor data(106) xor data(107) xor data(111) xor crcCur(0) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor data(49) xor data(50) xor data(51) xor data(54) xor data(59) xor data(60) xor data(69) xor data(71) xor data(78) xor data(80) xor data(81) xor data(85) xor data(86) xor data(87) xor data(89) xor data(90) xor data(92) xor data(93) xor data(94) xor data(97) xor data(100) xor data(102) xor data(103) xor data(105) xor data(106) xor data(107) xor data(108) xor crcCur(0) xor crcCur(1) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor data(48) xor data(50) xor data(51) xor data(52) xor data(55) xor data(60) xor data(61) xor data(70) xor data(72) xor data(79) xor data(81) xor data(82) xor data(86) xor data(87) xor data(88) xor data(90) xor data(91) xor data(93) xor data(94) xor data(95) xor data(98) xor data(101) xor data(103) xor data(104) xor data(106) xor data(107) xor data(108) xor data(109) xor crcCur(1) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(18) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor data(49) xor data(51) xor data(52) xor data(53) xor data(56) xor data(61) xor data(62) xor data(71) xor data(73) xor data(80) xor data(82) xor data(83) xor data(87) xor data(88) xor data(89) xor data(91) xor data(92) xor data(94) xor data(95) xor data(96) xor data(99) xor data(102) xor data(104) xor data(105) xor data(107) xor data(108) xor data(109) xor data(110) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(61) xor data(62) xor data(65) xor data(66) xor data(67) xor data(68) xor data(73) xor data(74) xor data(79) xor data(82) xor data(85) xor data(87) xor data(88) xor data(89) xor data(90) xor data(92) xor data(93) xor data(94) xor data(98) xor data(99) xor data(100) xor data(101) xor data(104) xor data(105) xor data(108) xor data(109) xor crcCur(2) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(29);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(54) xor data(55) xor data(56) xor data(59) xor data(60) xor data(62) xor data(65) xor data(69) xor data(72) xor data(73) xor data(74) xor data(75) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(85) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(93) xor data(96) xor data(97) xor data(98) xor data(100) xor data(102) xor data(103) xor data(104) xor data(105) xor data(109) xor data(111) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(29) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(55) xor data(56) xor data(57) xor data(60) xor data(61) xor data(63) xor data(66) xor data(70) xor data(73) xor data(74) xor data(75) xor data(76) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(94) xor data(97) xor data(98) xor data(99) xor data(101) xor data(103) xor data(104) xor data(105) xor data(106) xor data(110) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(30);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(56) xor data(57) xor data(58) xor data(61) xor data(62) xor data(64) xor data(67) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(95) xor data(98) xor data(99) xor data(100) xor data(102) xor data(104) xor data(105) xor data(106) xor data(107) xor data(111) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor data(48) xor data(49) xor data(52) xor data(54) xor data(55) xor data(57) xor data(59) xor data(60) xor data(61) xor data(62) xor data(66) xor data(67) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(81) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(95) xor data(97) xor data(98) xor data(100) xor data(104) xor data(105) xor data(107) xor data(108) xor data(110) xor data(111) xor crcCur(1) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor data(48) xor data(49) xor data(50) xor data(53) xor data(55) xor data(56) xor data(58) xor data(60) xor data(61) xor data(62) xor data(63) xor data(67) xor data(68) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(94) xor data(96) xor data(98) xor data(99) xor data(101) xor data(105) xor data(106) xor data(108) xor data(109) xor data(111) xor crcCur(0) xor crcCur(2) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(62) xor data(63) xor data(64) xor data(68) xor data(69) xor data(75) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(90) xor data(91) xor data(92) xor data(93) xor data(94) xor data(95) xor data(97) xor data(99) xor data(100) xor data(102) xor data(106) xor data(107) xor data(109) xor data(110) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(70) xor data(76) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(91) xor data(92) xor data(93) xor data(94) xor data(95) xor data(96) xor data(98) xor data(100) xor data(101) xor data(103) xor data(107) xor data(108) xor data(110) xor data(111) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor data(48) xor data(51) xor data(52) xor data(53) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(66) xor data(70) xor data(71) xor data(77) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(92) xor data(93) xor data(94) xor data(95) xor data(96) xor data(97) xor data(99) xor data(101) xor data(102) xor data(104) xor data(108) xor data(109) xor data(111) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor data(49) xor data(52) xor data(53) xor data(54) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(67) xor data(71) xor data(72) xor data(78) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(93) xor data(94) xor data(95) xor data(96) xor data(97) xor data(98) xor data(100) xor data(102) xor data(103) xor data(105) xor data(109) xor data(110) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(29) xor crcCur(30);
      return retVar;
   end function;

   function crc32Parallel15Byte (crcCur : slv(31 downto 0); data : slv(119 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(53) xor data(54) xor data(55) xor data(58) xor data(60) xor data(61) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(72) xor data(73) xor data(79) xor data(81) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor data(94) xor data(95) xor data(96) xor data(97) xor data(98) xor data(99) xor data(101) xor data(103) xor data(104) xor data(106) xor data(110) xor data(111) xor data(113) xor data(114) xor data(116) xor data(117) xor data(118) xor data(119) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(53) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(72) xor data(74) xor data(79) xor data(80) xor data(81) xor data(86) xor data(87) xor data(88) xor data(94) xor data(100) xor data(101) xor data(102) xor data(103) xor data(105) xor data(106) xor data(107) xor data(110) xor data(112) xor data(113) xor data(115) xor data(116) xor crcCur(0) xor crcCur(6) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor data(51) xor data(52) xor data(53) xor data(55) xor data(57) xor data(58) xor data(59) xor data(64) xor data(67) xor data(68) xor data(70) xor data(72) xor data(75) xor data(79) xor data(80) xor data(83) xor data(84) xor data(85) xor data(88) xor data(89) xor data(94) xor data(96) xor data(97) xor data(98) xor data(99) xor data(102) xor data(107) xor data(108) xor data(110) xor data(118) xor data(119) xor crcCur(0) xor crcCur(1) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(30) xor crcCur(31);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor data(52) xor data(53) xor data(54) xor data(56) xor data(58) xor data(59) xor data(60) xor data(65) xor data(68) xor data(69) xor data(71) xor data(73) xor data(76) xor data(80) xor data(81) xor data(84) xor data(85) xor data(86) xor data(89) xor data(90) xor data(95) xor data(97) xor data(98) xor data(99) xor data(100) xor data(103) xor data(108) xor data(109) xor data(111) xor data(119) xor crcCur(1) xor crcCur(2) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(31);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor data(48) xor data(50) xor data(57) xor data(58) xor data(59) xor data(63) xor data(65) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(74) xor data(77) xor data(79) xor data(83) xor data(84) xor data(86) xor data(90) xor data(91) xor data(94) xor data(95) xor data(97) xor data(100) xor data(103) xor data(106) xor data(109) xor data(111) xor data(112) xor data(113) xor data(114) xor data(116) xor data(117) xor data(118) xor data(119) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(12) xor crcCur(15) xor crcCur(18) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(53) xor data(54) xor data(55) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(67) xor data(69) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(91) xor data(92) xor data(94) xor data(97) xor data(99) xor data(103) xor data(106) xor data(107) xor data(111) xor data(112) xor data(115) xor data(116) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(9) xor crcCur(11) xor crcCur(15) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(28);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(55) xor data(56) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(76) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(92) xor data(93) xor data(95) xor data(98) xor data(100) xor data(104) xor data(107) xor data(108) xor data(112) xor data(113) xor data(116) xor data(117) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(12) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(29);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(56) xor data(57) xor data(58) xor data(60) xor data(68) xor data(69) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(79) xor data(80) xor data(87) xor data(93) xor data(95) xor data(97) xor data(98) xor data(103) xor data(104) xor data(105) xor data(106) xor data(108) xor data(109) xor data(110) xor data(111) xor data(116) xor data(119) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(28) xor crcCur(31);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor data(50) xor data(51) xor data(52) xor data(54) xor data(57) xor data(59) xor data(60) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor data(88) xor data(95) xor data(97) xor data(101) xor data(103) xor data(105) xor data(107) xor data(109) xor data(112) xor data(113) xor data(114) xor data(116) xor data(118) xor data(119) xor crcCur(0) xor crcCur(7) xor crcCur(9) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor data(51) xor data(52) xor data(53) xor data(55) xor data(58) xor data(60) xor data(61) xor data(64) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(71) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(84) xor data(85) xor data(86) xor data(88) xor data(89) xor data(96) xor data(98) xor data(102) xor data(104) xor data(106) xor data(108) xor data(110) xor data(113) xor data(114) xor data(115) xor data(117) xor data(119) xor crcCur(0) xor crcCur(1) xor crcCur(8) xor crcCur(10) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor data(50) xor data(52) xor data(55) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(66) xor data(69) xor data(70) xor data(71) xor data(73) xor data(75) xor data(77) xor data(78) xor data(80) xor data(83) xor data(86) xor data(89) xor data(90) xor data(94) xor data(95) xor data(96) xor data(98) xor data(101) xor data(104) xor data(105) xor data(106) xor data(107) xor data(109) xor data(110) xor data(113) xor data(115) xor data(117) xor data(119) xor crcCur(1) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(25) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(51) xor data(54) xor data(55) xor data(56) xor data(57) xor data(58) xor data(59) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(73) xor data(74) xor data(76) xor data(78) xor data(82) xor data(83) xor data(85) xor data(90) xor data(91) xor data(94) xor data(98) xor data(101) xor data(102) xor data(103) xor data(104) xor data(105) xor data(107) xor data(108) xor data(113) xor data(117) xor data(119) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(10) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(25) xor crcCur(29) xor crcCur(31);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(63) xor data(68) xor data(69) xor data(71) xor data(73) xor data(74) xor data(75) xor data(77) xor data(81) xor data(82) xor data(85) xor data(86) xor data(87) xor data(91) xor data(92) xor data(94) xor data(96) xor data(97) xor data(98) xor data(101) xor data(102) xor data(105) xor data(108) xor data(109) xor data(110) xor data(111) xor data(113) xor data(116) xor data(117) xor data(119) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(64) xor data(69) xor data(70) xor data(72) xor data(74) xor data(75) xor data(76) xor data(78) xor data(82) xor data(83) xor data(86) xor data(87) xor data(88) xor data(92) xor data(93) xor data(95) xor data(97) xor data(98) xor data(99) xor data(102) xor data(103) xor data(106) xor data(109) xor data(110) xor data(111) xor data(112) xor data(114) xor data(117) xor data(118) xor crcCur(0) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(15) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(29) xor crcCur(30);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(65) xor data(70) xor data(71) xor data(73) xor data(75) xor data(76) xor data(77) xor data(79) xor data(83) xor data(84) xor data(87) xor data(88) xor data(89) xor data(93) xor data(94) xor data(96) xor data(98) xor data(99) xor data(100) xor data(103) xor data(104) xor data(107) xor data(110) xor data(111) xor data(112) xor data(113) xor data(115) xor data(118) xor data(119) xor crcCur(0) xor crcCur(1) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor data(49) xor data(50) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(66) xor data(71) xor data(72) xor data(74) xor data(76) xor data(77) xor data(78) xor data(80) xor data(84) xor data(85) xor data(88) xor data(89) xor data(90) xor data(94) xor data(95) xor data(97) xor data(99) xor data(100) xor data(101) xor data(104) xor data(105) xor data(108) xor data(111) xor data(112) xor data(113) xor data(114) xor data(116) xor data(119) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(31);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor data(48) xor data(51) xor data(56) xor data(57) xor data(66) xor data(68) xor data(75) xor data(77) xor data(78) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor data(89) xor data(90) xor data(91) xor data(94) xor data(97) xor data(99) xor data(100) xor data(102) xor data(103) xor data(104) xor data(105) xor data(109) xor data(110) xor data(111) xor data(112) xor data(115) xor data(116) xor data(118) xor data(119) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor data(48) xor data(49) xor data(52) xor data(57) xor data(58) xor data(67) xor data(69) xor data(76) xor data(78) xor data(79) xor data(83) xor data(84) xor data(85) xor data(87) xor data(88) xor data(90) xor data(91) xor data(92) xor data(95) xor data(98) xor data(100) xor data(101) xor data(103) xor data(104) xor data(105) xor data(106) xor data(110) xor data(111) xor data(112) xor data(113) xor data(116) xor data(117) xor data(119) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(29) xor crcCur(31);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor data(48) xor data(49) xor data(50) xor data(53) xor data(58) xor data(59) xor data(68) xor data(70) xor data(77) xor data(79) xor data(80) xor data(84) xor data(85) xor data(86) xor data(88) xor data(89) xor data(91) xor data(92) xor data(93) xor data(96) xor data(99) xor data(101) xor data(102) xor data(104) xor data(105) xor data(106) xor data(107) xor data(111) xor data(112) xor data(113) xor data(114) xor data(117) xor data(118) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(29) xor crcCur(30);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor data(49) xor data(50) xor data(51) xor data(54) xor data(59) xor data(60) xor data(69) xor data(71) xor data(78) xor data(80) xor data(81) xor data(85) xor data(86) xor data(87) xor data(89) xor data(90) xor data(92) xor data(93) xor data(94) xor data(97) xor data(100) xor data(102) xor data(103) xor data(105) xor data(106) xor data(107) xor data(108) xor data(112) xor data(113) xor data(114) xor data(115) xor data(118) xor data(119) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(30) xor crcCur(31);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor data(48) xor data(50) xor data(51) xor data(52) xor data(55) xor data(60) xor data(61) xor data(70) xor data(72) xor data(79) xor data(81) xor data(82) xor data(86) xor data(87) xor data(88) xor data(90) xor data(91) xor data(93) xor data(94) xor data(95) xor data(98) xor data(101) xor data(103) xor data(104) xor data(106) xor data(107) xor data(108) xor data(109) xor data(113) xor data(114) xor data(115) xor data(116) xor data(119) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(10) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor data(49) xor data(51) xor data(52) xor data(53) xor data(56) xor data(61) xor data(62) xor data(71) xor data(73) xor data(80) xor data(82) xor data(83) xor data(87) xor data(88) xor data(89) xor data(91) xor data(92) xor data(94) xor data(95) xor data(96) xor data(99) xor data(102) xor data(104) xor data(105) xor data(107) xor data(108) xor data(109) xor data(110) xor data(114) xor data(115) xor data(116) xor data(117) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(11) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(61) xor data(62) xor data(65) xor data(66) xor data(67) xor data(68) xor data(73) xor data(74) xor data(79) xor data(82) xor data(85) xor data(87) xor data(88) xor data(89) xor data(90) xor data(92) xor data(93) xor data(94) xor data(98) xor data(99) xor data(100) xor data(101) xor data(104) xor data(105) xor data(108) xor data(109) xor data(113) xor data(114) xor data(115) xor data(119) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(54) xor data(55) xor data(56) xor data(59) xor data(60) xor data(62) xor data(65) xor data(69) xor data(72) xor data(73) xor data(74) xor data(75) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(85) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(93) xor data(96) xor data(97) xor data(98) xor data(100) xor data(102) xor data(103) xor data(104) xor data(105) xor data(109) xor data(111) xor data(113) xor data(115) xor data(117) xor data(118) xor data(119) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(21) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(55) xor data(56) xor data(57) xor data(60) xor data(61) xor data(63) xor data(66) xor data(70) xor data(73) xor data(74) xor data(75) xor data(76) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(94) xor data(97) xor data(98) xor data(99) xor data(101) xor data(103) xor data(104) xor data(105) xor data(106) xor data(110) xor data(112) xor data(114) xor data(116) xor data(118) xor data(119) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(24) xor crcCur(26) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(56) xor data(57) xor data(58) xor data(61) xor data(62) xor data(64) xor data(67) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(95) xor data(98) xor data(99) xor data(100) xor data(102) xor data(104) xor data(105) xor data(106) xor data(107) xor data(111) xor data(113) xor data(115) xor data(117) xor data(119) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor data(48) xor data(49) xor data(52) xor data(54) xor data(55) xor data(57) xor data(59) xor data(60) xor data(61) xor data(62) xor data(66) xor data(67) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(81) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(95) xor data(97) xor data(98) xor data(100) xor data(104) xor data(105) xor data(107) xor data(108) xor data(110) xor data(111) xor data(112) xor data(113) xor data(117) xor data(119) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(29) xor crcCur(31);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor data(48) xor data(49) xor data(50) xor data(53) xor data(55) xor data(56) xor data(58) xor data(60) xor data(61) xor data(62) xor data(63) xor data(67) xor data(68) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(94) xor data(96) xor data(98) xor data(99) xor data(101) xor data(105) xor data(106) xor data(108) xor data(109) xor data(111) xor data(112) xor data(113) xor data(114) xor data(118) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(30);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(62) xor data(63) xor data(64) xor data(68) xor data(69) xor data(75) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(90) xor data(91) xor data(92) xor data(93) xor data(94) xor data(95) xor data(97) xor data(99) xor data(100) xor data(102) xor data(106) xor data(107) xor data(109) xor data(110) xor data(112) xor data(113) xor data(114) xor data(115) xor data(119) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(70) xor data(76) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(91) xor data(92) xor data(93) xor data(94) xor data(95) xor data(96) xor data(98) xor data(100) xor data(101) xor data(103) xor data(107) xor data(108) xor data(110) xor data(111) xor data(113) xor data(114) xor data(115) xor data(116) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor data(48) xor data(51) xor data(52) xor data(53) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(66) xor data(70) xor data(71) xor data(77) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(92) xor data(93) xor data(94) xor data(95) xor data(96) xor data(97) xor data(99) xor data(101) xor data(102) xor data(104) xor data(108) xor data(109) xor data(111) xor data(112) xor data(114) xor data(115) xor data(116) xor data(117) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor data(49) xor data(52) xor data(53) xor data(54) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(67) xor data(71) xor data(72) xor data(78) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(93) xor data(94) xor data(95) xor data(96) xor data(97) xor data(98) xor data(100) xor data(102) xor data(103) xor data(105) xor data(109) xor data(110) xor data(112) xor data(113) xor data(115) xor data(116) xor data(117) xor data(118) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      return retVar;
   end function;

   function crc32Parallel16Byte (crcCur : slv(31 downto 0); data : slv(127 downto 0)) return slv is
      variable retVar : slv(31 downto 0) := (others => '0');
   begin
      retVar(0) := data(0) xor data(6) xor data(9) xor data(10) xor data(12) xor data(16) xor data(24) xor data(25) xor data(26) xor data(28) xor data(29) xor data(30) xor data(31) xor data(32) xor data(34) xor data(37) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(53) xor data(54) xor data(55) xor data(58) xor data(60) xor data(61) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(72) xor data(73) xor data(79) xor data(81) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor data(94) xor data(95) xor data(96) xor data(97) xor data(98) xor data(99) xor data(101) xor data(103) xor data(104) xor data(106) xor data(110) xor data(111) xor data(113) xor data(114) xor data(116) xor data(117) xor data(118) xor data(119) xor data(123) xor data(125) xor data(126) xor data(127) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(1) := data(0) xor data(1) xor data(6) xor data(7) xor data(9) xor data(11) xor data(12) xor data(13) xor data(16) xor data(17) xor data(24) xor data(27) xor data(28) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(44) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(53) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(72) xor data(74) xor data(79) xor data(80) xor data(81) xor data(86) xor data(87) xor data(88) xor data(94) xor data(100) xor data(101) xor data(102) xor data(103) xor data(105) xor data(106) xor data(107) xor data(110) xor data(112) xor data(113) xor data(115) xor data(116) xor data(120) xor data(123) xor data(124) xor data(125) xor crcCur(4) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(2) := data(0) xor data(1) xor data(2) xor data(6) xor data(7) xor data(8) xor data(9) xor data(13) xor data(14) xor data(16) xor data(17) xor data(18) xor data(24) xor data(26) xor data(30) xor data(31) xor data(32) xor data(35) xor data(36) xor data(37) xor data(38) xor data(39) xor data(44) xor data(51) xor data(52) xor data(53) xor data(55) xor data(57) xor data(58) xor data(59) xor data(64) xor data(67) xor data(68) xor data(70) xor data(72) xor data(75) xor data(79) xor data(80) xor data(83) xor data(84) xor data(85) xor data(88) xor data(89) xor data(94) xor data(96) xor data(97) xor data(98) xor data(99) xor data(102) xor data(107) xor data(108) xor data(110) xor data(118) xor data(119) xor data(121) xor data(123) xor data(124) xor data(127) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(3) := data(1) xor data(2) xor data(3) xor data(7) xor data(8) xor data(9) xor data(10) xor data(14) xor data(15) xor data(17) xor data(18) xor data(19) xor data(25) xor data(27) xor data(31) xor data(32) xor data(33) xor data(36) xor data(37) xor data(38) xor data(39) xor data(40) xor data(45) xor data(52) xor data(53) xor data(54) xor data(56) xor data(58) xor data(59) xor data(60) xor data(65) xor data(68) xor data(69) xor data(71) xor data(73) xor data(76) xor data(80) xor data(81) xor data(84) xor data(85) xor data(86) xor data(89) xor data(90) xor data(95) xor data(97) xor data(98) xor data(99) xor data(100) xor data(103) xor data(108) xor data(109) xor data(111) xor data(119) xor data(120) xor data(122) xor data(124) xor data(125) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(28) xor crcCur(29);
      retVar(4) := data(0) xor data(2) xor data(3) xor data(4) xor data(6) xor data(8) xor data(11) xor data(12) xor data(15) xor data(18) xor data(19) xor data(20) xor data(24) xor data(25) xor data(29) xor data(30) xor data(31) xor data(33) xor data(38) xor data(39) xor data(40) xor data(41) xor data(44) xor data(45) xor data(46) xor data(47) xor data(48) xor data(50) xor data(57) xor data(58) xor data(59) xor data(63) xor data(65) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(74) xor data(77) xor data(79) xor data(83) xor data(84) xor data(86) xor data(90) xor data(91) xor data(94) xor data(95) xor data(97) xor data(100) xor data(103) xor data(106) xor data(109) xor data(111) xor data(112) xor data(113) xor data(114) xor data(116) xor data(117) xor data(118) xor data(119) xor data(120) xor data(121) xor data(127) xor crcCur(1) xor crcCur(4) xor crcCur(7) xor crcCur(10) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(31);
      retVar(5) := data(0) xor data(1) xor data(3) xor data(4) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(19) xor data(20) xor data(21) xor data(24) xor data(28) xor data(29) xor data(37) xor data(39) xor data(40) xor data(41) xor data(42) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(53) xor data(54) xor data(55) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(67) xor data(69) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(91) xor data(92) xor data(94) xor data(97) xor data(99) xor data(103) xor data(106) xor data(107) xor data(111) xor data(112) xor data(115) xor data(116) xor data(120) xor data(121) xor data(122) xor data(123) xor data(125) xor data(126) xor data(127) xor crcCur(1) xor crcCur(3) xor crcCur(7) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(6) := data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(20) xor data(21) xor data(22) xor data(25) xor data(29) xor data(30) xor data(38) xor data(40) xor data(41) xor data(42) xor data(43) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(55) xor data(56) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(72) xor data(73) xor data(74) xor data(75) xor data(76) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(92) xor data(93) xor data(95) xor data(98) xor data(100) xor data(104) xor data(107) xor data(108) xor data(112) xor data(113) xor data(116) xor data(117) xor data(121) xor data(122) xor data(123) xor data(124) xor data(126) xor data(127) xor crcCur(2) xor crcCur(4) xor crcCur(8) xor crcCur(11) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(7) := data(0) xor data(2) xor data(3) xor data(5) xor data(7) xor data(8) xor data(10) xor data(15) xor data(16) xor data(21) xor data(22) xor data(23) xor data(24) xor data(25) xor data(28) xor data(29) xor data(32) xor data(34) xor data(37) xor data(39) xor data(41) xor data(42) xor data(43) xor data(45) xor data(46) xor data(47) xor data(50) xor data(51) xor data(52) xor data(54) xor data(56) xor data(57) xor data(58) xor data(60) xor data(68) xor data(69) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(79) xor data(80) xor data(87) xor data(93) xor data(95) xor data(97) xor data(98) xor data(103) xor data(104) xor data(105) xor data(106) xor data(108) xor data(109) xor data(110) xor data(111) xor data(116) xor data(119) xor data(122) xor data(124) xor data(126) xor crcCur(1) xor crcCur(2) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(20) xor crcCur(23) xor crcCur(26) xor crcCur(28) xor crcCur(30);
      retVar(8) := data(0) xor data(1) xor data(3) xor data(4) xor data(8) xor data(10) xor data(11) xor data(12) xor data(17) xor data(22) xor data(23) xor data(28) xor data(31) xor data(32) xor data(33) xor data(34) xor data(35) xor data(37) xor data(38) xor data(40) xor data(42) xor data(43) xor data(45) xor data(46) xor data(50) xor data(51) xor data(52) xor data(54) xor data(57) xor data(59) xor data(60) xor data(63) xor data(65) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(83) xor data(84) xor data(85) xor data(87) xor data(88) xor data(95) xor data(97) xor data(101) xor data(103) xor data(105) xor data(107) xor data(109) xor data(112) xor data(113) xor data(114) xor data(116) xor data(118) xor data(119) xor data(120) xor data(126) xor crcCur(1) xor crcCur(5) xor crcCur(7) xor crcCur(9) xor crcCur(11) xor crcCur(13) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(30);
      retVar(9) := data(1) xor data(2) xor data(4) xor data(5) xor data(9) xor data(11) xor data(12) xor data(13) xor data(18) xor data(23) xor data(24) xor data(29) xor data(32) xor data(33) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(41) xor data(43) xor data(44) xor data(46) xor data(47) xor data(51) xor data(52) xor data(53) xor data(55) xor data(58) xor data(60) xor data(61) xor data(64) xor data(66) xor data(67) xor data(68) xor data(69) xor data(70) xor data(71) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(84) xor data(85) xor data(86) xor data(88) xor data(89) xor data(96) xor data(98) xor data(102) xor data(104) xor data(106) xor data(108) xor data(110) xor data(113) xor data(114) xor data(115) xor data(117) xor data(119) xor data(120) xor data(121) xor data(127) xor crcCur(0) xor crcCur(2) xor crcCur(6) xor crcCur(8) xor crcCur(10) xor crcCur(12) xor crcCur(14) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(31);
      retVar(10) := data(0) xor data(2) xor data(3) xor data(5) xor data(9) xor data(13) xor data(14) xor data(16) xor data(19) xor data(26) xor data(28) xor data(29) xor data(31) xor data(32) xor data(33) xor data(35) xor data(36) xor data(39) xor data(40) xor data(42) xor data(50) xor data(52) xor data(55) xor data(56) xor data(58) xor data(59) xor data(60) xor data(62) xor data(63) xor data(66) xor data(69) xor data(70) xor data(71) xor data(73) xor data(75) xor data(77) xor data(78) xor data(80) xor data(83) xor data(86) xor data(89) xor data(90) xor data(94) xor data(95) xor data(96) xor data(98) xor data(101) xor data(104) xor data(105) xor data(106) xor data(107) xor data(109) xor data(110) xor data(113) xor data(115) xor data(117) xor data(119) xor data(120) xor data(121) xor data(122) xor data(123) xor data(125) xor data(126) xor data(127) xor crcCur(0) xor crcCur(2) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      retVar(11) := data(0) xor data(1) xor data(3) xor data(4) xor data(9) xor data(12) xor data(14) xor data(15) xor data(16) xor data(17) xor data(20) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(31) xor data(33) xor data(36) xor data(40) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(50) xor data(51) xor data(54) xor data(55) xor data(56) xor data(57) xor data(58) xor data(59) xor data(64) xor data(65) xor data(66) xor data(68) xor data(70) xor data(71) xor data(73) xor data(74) xor data(76) xor data(78) xor data(82) xor data(83) xor data(85) xor data(90) xor data(91) xor data(94) xor data(98) xor data(101) xor data(102) xor data(103) xor data(104) xor data(105) xor data(107) xor data(108) xor data(113) xor data(117) xor data(119) xor data(120) xor data(121) xor data(122) xor data(124) xor data(125) xor crcCur(2) xor crcCur(5) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(17) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(29);
      retVar(12) := data(0) xor data(1) xor data(2) xor data(4) xor data(5) xor data(6) xor data(9) xor data(12) xor data(13) xor data(15) xor data(17) xor data(18) xor data(21) xor data(24) xor data(27) xor data(30) xor data(31) xor data(41) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(63) xor data(68) xor data(69) xor data(71) xor data(73) xor data(74) xor data(75) xor data(77) xor data(81) xor data(82) xor data(85) xor data(86) xor data(87) xor data(91) xor data(92) xor data(94) xor data(96) xor data(97) xor data(98) xor data(101) xor data(102) xor data(105) xor data(108) xor data(109) xor data(110) xor data(111) xor data(113) xor data(116) xor data(117) xor data(119) xor data(120) xor data(121) xor data(122) xor data(127) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(5) xor crcCur(6) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(31);
      retVar(13) := data(1) xor data(2) xor data(3) xor data(5) xor data(6) xor data(7) xor data(10) xor data(13) xor data(14) xor data(16) xor data(18) xor data(19) xor data(22) xor data(25) xor data(28) xor data(31) xor data(32) xor data(42) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(64) xor data(69) xor data(70) xor data(72) xor data(74) xor data(75) xor data(76) xor data(78) xor data(82) xor data(83) xor data(86) xor data(87) xor data(88) xor data(92) xor data(93) xor data(95) xor data(97) xor data(98) xor data(99) xor data(102) xor data(103) xor data(106) xor data(109) xor data(110) xor data(111) xor data(112) xor data(114) xor data(117) xor data(118) xor data(120) xor data(121) xor data(122) xor data(123) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(6) xor crcCur(7) xor crcCur(10) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27);
      retVar(14) := data(2) xor data(3) xor data(4) xor data(6) xor data(7) xor data(8) xor data(11) xor data(14) xor data(15) xor data(17) xor data(19) xor data(20) xor data(23) xor data(26) xor data(29) xor data(32) xor data(33) xor data(43) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(65) xor data(70) xor data(71) xor data(73) xor data(75) xor data(76) xor data(77) xor data(79) xor data(83) xor data(84) xor data(87) xor data(88) xor data(89) xor data(93) xor data(94) xor data(96) xor data(98) xor data(99) xor data(100) xor data(103) xor data(104) xor data(107) xor data(110) xor data(111) xor data(112) xor data(113) xor data(115) xor data(118) xor data(119) xor data(121) xor data(122) xor data(123) xor data(124) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(7) xor crcCur(8) xor crcCur(11) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(15) := data(3) xor data(4) xor data(5) xor data(7) xor data(8) xor data(9) xor data(12) xor data(15) xor data(16) xor data(18) xor data(20) xor data(21) xor data(24) xor data(27) xor data(30) xor data(33) xor data(34) xor data(44) xor data(45) xor data(49) xor data(50) xor data(52) xor data(53) xor data(54) xor data(55) xor data(56) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(66) xor data(71) xor data(72) xor data(74) xor data(76) xor data(77) xor data(78) xor data(80) xor data(84) xor data(85) xor data(88) xor data(89) xor data(90) xor data(94) xor data(95) xor data(97) xor data(99) xor data(100) xor data(101) xor data(104) xor data(105) xor data(108) xor data(111) xor data(112) xor data(113) xor data(114) xor data(116) xor data(119) xor data(120) xor data(122) xor data(123) xor data(124) xor data(125) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(16) := data(0) xor data(4) xor data(5) xor data(8) xor data(12) xor data(13) xor data(17) xor data(19) xor data(21) xor data(22) xor data(24) xor data(26) xor data(29) xor data(30) xor data(32) xor data(35) xor data(37) xor data(44) xor data(46) xor data(47) xor data(48) xor data(51) xor data(56) xor data(57) xor data(66) xor data(68) xor data(75) xor data(77) xor data(78) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor data(89) xor data(90) xor data(91) xor data(94) xor data(97) xor data(99) xor data(100) xor data(102) xor data(103) xor data(104) xor data(105) xor data(109) xor data(110) xor data(111) xor data(112) xor data(115) xor data(116) xor data(118) xor data(119) xor data(120) xor data(121) xor data(124) xor data(127) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(19) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(28) xor crcCur(31);
      retVar(17) := data(1) xor data(5) xor data(6) xor data(9) xor data(13) xor data(14) xor data(18) xor data(20) xor data(22) xor data(23) xor data(25) xor data(27) xor data(30) xor data(31) xor data(33) xor data(36) xor data(38) xor data(45) xor data(47) xor data(48) xor data(49) xor data(52) xor data(57) xor data(58) xor data(67) xor data(69) xor data(76) xor data(78) xor data(79) xor data(83) xor data(84) xor data(85) xor data(87) xor data(88) xor data(90) xor data(91) xor data(92) xor data(95) xor data(98) xor data(100) xor data(101) xor data(103) xor data(104) xor data(105) xor data(106) xor data(110) xor data(111) xor data(112) xor data(113) xor data(116) xor data(117) xor data(119) xor data(120) xor data(121) xor data(122) xor data(125) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(20) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(29);
      retVar(18) := data(2) xor data(6) xor data(7) xor data(10) xor data(14) xor data(15) xor data(19) xor data(21) xor data(23) xor data(24) xor data(26) xor data(28) xor data(31) xor data(32) xor data(34) xor data(37) xor data(39) xor data(46) xor data(48) xor data(49) xor data(50) xor data(53) xor data(58) xor data(59) xor data(68) xor data(70) xor data(77) xor data(79) xor data(80) xor data(84) xor data(85) xor data(86) xor data(88) xor data(89) xor data(91) xor data(92) xor data(93) xor data(96) xor data(99) xor data(101) xor data(102) xor data(104) xor data(105) xor data(106) xor data(107) xor data(111) xor data(112) xor data(113) xor data(114) xor data(117) xor data(118) xor data(120) xor data(121) xor data(122) xor data(123) xor data(126) xor crcCur(0) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(21) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(30);
      retVar(19) := data(3) xor data(7) xor data(8) xor data(11) xor data(15) xor data(16) xor data(20) xor data(22) xor data(24) xor data(25) xor data(27) xor data(29) xor data(32) xor data(33) xor data(35) xor data(38) xor data(40) xor data(47) xor data(49) xor data(50) xor data(51) xor data(54) xor data(59) xor data(60) xor data(69) xor data(71) xor data(78) xor data(80) xor data(81) xor data(85) xor data(86) xor data(87) xor data(89) xor data(90) xor data(92) xor data(93) xor data(94) xor data(97) xor data(100) xor data(102) xor data(103) xor data(105) xor data(106) xor data(107) xor data(108) xor data(112) xor data(113) xor data(114) xor data(115) xor data(118) xor data(119) xor data(121) xor data(122) xor data(123) xor data(124) xor data(127) xor crcCur(1) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(22) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(31);
      retVar(20) := data(4) xor data(8) xor data(9) xor data(12) xor data(16) xor data(17) xor data(21) xor data(23) xor data(25) xor data(26) xor data(28) xor data(30) xor data(33) xor data(34) xor data(36) xor data(39) xor data(41) xor data(48) xor data(50) xor data(51) xor data(52) xor data(55) xor data(60) xor data(61) xor data(70) xor data(72) xor data(79) xor data(81) xor data(82) xor data(86) xor data(87) xor data(88) xor data(90) xor data(91) xor data(93) xor data(94) xor data(95) xor data(98) xor data(101) xor data(103) xor data(104) xor data(106) xor data(107) xor data(108) xor data(109) xor data(113) xor data(114) xor data(115) xor data(116) xor data(119) xor data(120) xor data(122) xor data(123) xor data(124) xor data(125) xor crcCur(2) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(10) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(21) := data(5) xor data(9) xor data(10) xor data(13) xor data(17) xor data(18) xor data(22) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(37) xor data(40) xor data(42) xor data(49) xor data(51) xor data(52) xor data(53) xor data(56) xor data(61) xor data(62) xor data(71) xor data(73) xor data(80) xor data(82) xor data(83) xor data(87) xor data(88) xor data(89) xor data(91) xor data(92) xor data(94) xor data(95) xor data(96) xor data(99) xor data(102) xor data(104) xor data(105) xor data(107) xor data(108) xor data(109) xor data(110) xor data(114) xor data(115) xor data(116) xor data(117) xor data(120) xor data(121) xor data(123) xor data(124) xor data(125) xor data(126) xor crcCur(0) xor crcCur(3) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(13) xor crcCur(14) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(22) := data(0) xor data(9) xor data(11) xor data(12) xor data(14) xor data(16) xor data(18) xor data(19) xor data(23) xor data(24) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(37) xor data(38) xor data(41) xor data(43) xor data(44) xor data(45) xor data(47) xor data(48) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(61) xor data(62) xor data(65) xor data(66) xor data(67) xor data(68) xor data(73) xor data(74) xor data(79) xor data(82) xor data(85) xor data(87) xor data(88) xor data(89) xor data(90) xor data(92) xor data(93) xor data(94) xor data(98) xor data(99) xor data(100) xor data(101) xor data(104) xor data(105) xor data(108) xor data(109) xor data(113) xor data(114) xor data(115) xor data(119) xor data(121) xor data(122) xor data(123) xor data(124) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(5) xor crcCur(8) xor crcCur(9) xor crcCur(12) xor crcCur(13) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(23) := data(0) xor data(1) xor data(6) xor data(9) xor data(13) xor data(15) xor data(16) xor data(17) xor data(19) xor data(20) xor data(26) xor data(27) xor data(29) xor data(31) xor data(34) xor data(35) xor data(36) xor data(38) xor data(39) xor data(42) xor data(46) xor data(47) xor data(49) xor data(50) xor data(54) xor data(55) xor data(56) xor data(59) xor data(60) xor data(62) xor data(65) xor data(69) xor data(72) xor data(73) xor data(74) xor data(75) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(85) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(93) xor data(96) xor data(97) xor data(98) xor data(100) xor data(102) xor data(103) xor data(104) xor data(105) xor data(109) xor data(111) xor data(113) xor data(115) xor data(117) xor data(118) xor data(119) xor data(120) xor data(122) xor data(124) xor data(126) xor data(127) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(13) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(26) xor crcCur(28) xor crcCur(30) xor crcCur(31);
      retVar(24) := data(1) xor data(2) xor data(7) xor data(10) xor data(14) xor data(16) xor data(17) xor data(18) xor data(20) xor data(21) xor data(27) xor data(28) xor data(30) xor data(32) xor data(35) xor data(36) xor data(37) xor data(39) xor data(40) xor data(43) xor data(47) xor data(48) xor data(50) xor data(51) xor data(55) xor data(56) xor data(57) xor data(60) xor data(61) xor data(63) xor data(66) xor data(70) xor data(73) xor data(74) xor data(75) xor data(76) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(94) xor data(97) xor data(98) xor data(99) xor data(101) xor data(103) xor data(104) xor data(105) xor data(106) xor data(110) xor data(112) xor data(114) xor data(116) xor data(118) xor data(119) xor data(120) xor data(121) xor data(123) xor data(125) xor data(127) xor crcCur(1) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(7) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(14) xor crcCur(16) xor crcCur(18) xor crcCur(20) xor crcCur(22) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(27) xor crcCur(29) xor crcCur(31);
      retVar(25) := data(2) xor data(3) xor data(8) xor data(11) xor data(15) xor data(17) xor data(18) xor data(19) xor data(21) xor data(22) xor data(28) xor data(29) xor data(31) xor data(33) xor data(36) xor data(37) xor data(38) xor data(40) xor data(41) xor data(44) xor data(48) xor data(49) xor data(51) xor data(52) xor data(56) xor data(57) xor data(58) xor data(61) xor data(62) xor data(64) xor data(67) xor data(71) xor data(74) xor data(75) xor data(76) xor data(77) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(87) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(95) xor data(98) xor data(99) xor data(100) xor data(102) xor data(104) xor data(105) xor data(106) xor data(107) xor data(111) xor data(113) xor data(115) xor data(117) xor data(119) xor data(120) xor data(121) xor data(122) xor data(124) xor data(126) xor crcCur(2) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(8) xor crcCur(9) xor crcCur(10) xor crcCur(11) xor crcCur(15) xor crcCur(17) xor crcCur(19) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(28) xor crcCur(30);
      retVar(26) := data(0) xor data(3) xor data(4) xor data(6) xor data(10) xor data(18) xor data(19) xor data(20) xor data(22) xor data(23) xor data(24) xor data(25) xor data(26) xor data(28) xor data(31) xor data(38) xor data(39) xor data(41) xor data(42) xor data(44) xor data(47) xor data(48) xor data(49) xor data(52) xor data(54) xor data(55) xor data(57) xor data(59) xor data(60) xor data(61) xor data(62) xor data(66) xor data(67) xor data(73) xor data(75) xor data(76) xor data(77) xor data(78) xor data(79) xor data(81) xor data(88) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(95) xor data(97) xor data(98) xor data(100) xor data(104) xor data(105) xor data(107) xor data(108) xor data(110) xor data(111) xor data(112) xor data(113) xor data(117) xor data(119) xor data(120) xor data(121) xor data(122) xor data(126) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(8) xor crcCur(9) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(21) xor crcCur(23) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(30);
      retVar(27) := data(1) xor data(4) xor data(5) xor data(7) xor data(11) xor data(19) xor data(20) xor data(21) xor data(23) xor data(24) xor data(25) xor data(26) xor data(27) xor data(29) xor data(32) xor data(39) xor data(40) xor data(42) xor data(43) xor data(45) xor data(48) xor data(49) xor data(50) xor data(53) xor data(55) xor data(56) xor data(58) xor data(60) xor data(61) xor data(62) xor data(63) xor data(67) xor data(68) xor data(74) xor data(76) xor data(77) xor data(78) xor data(79) xor data(80) xor data(82) xor data(89) xor data(90) xor data(91) xor data(92) xor data(93) xor data(94) xor data(96) xor data(98) xor data(99) xor data(101) xor data(105) xor data(106) xor data(108) xor data(109) xor data(111) xor data(112) xor data(113) xor data(114) xor data(118) xor data(120) xor data(121) xor data(122) xor data(123) xor data(127) xor crcCur(0) xor crcCur(2) xor crcCur(3) xor crcCur(5) xor crcCur(9) xor crcCur(10) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(22) xor crcCur(24) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(31);
      retVar(28) := data(2) xor data(5) xor data(6) xor data(8) xor data(12) xor data(20) xor data(21) xor data(22) xor data(24) xor data(25) xor data(26) xor data(27) xor data(28) xor data(30) xor data(33) xor data(40) xor data(41) xor data(43) xor data(44) xor data(46) xor data(49) xor data(50) xor data(51) xor data(54) xor data(56) xor data(57) xor data(59) xor data(61) xor data(62) xor data(63) xor data(64) xor data(68) xor data(69) xor data(75) xor data(77) xor data(78) xor data(79) xor data(80) xor data(81) xor data(83) xor data(90) xor data(91) xor data(92) xor data(93) xor data(94) xor data(95) xor data(97) xor data(99) xor data(100) xor data(102) xor data(106) xor data(107) xor data(109) xor data(110) xor data(112) xor data(113) xor data(114) xor data(115) xor data(119) xor data(121) xor data(122) xor data(123) xor data(124) xor crcCur(1) xor crcCur(3) xor crcCur(4) xor crcCur(6) xor crcCur(10) xor crcCur(11) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(23) xor crcCur(25) xor crcCur(26) xor crcCur(27) xor crcCur(28);
      retVar(29) := data(3) xor data(6) xor data(7) xor data(9) xor data(13) xor data(21) xor data(22) xor data(23) xor data(25) xor data(26) xor data(27) xor data(28) xor data(29) xor data(31) xor data(34) xor data(41) xor data(42) xor data(44) xor data(45) xor data(47) xor data(50) xor data(51) xor data(52) xor data(55) xor data(57) xor data(58) xor data(60) xor data(62) xor data(63) xor data(64) xor data(65) xor data(69) xor data(70) xor data(76) xor data(78) xor data(79) xor data(80) xor data(81) xor data(82) xor data(84) xor data(91) xor data(92) xor data(93) xor data(94) xor data(95) xor data(96) xor data(98) xor data(100) xor data(101) xor data(103) xor data(107) xor data(108) xor data(110) xor data(111) xor data(113) xor data(114) xor data(115) xor data(116) xor data(120) xor data(122) xor data(123) xor data(124) xor data(125) xor crcCur(0) xor crcCur(2) xor crcCur(4) xor crcCur(5) xor crcCur(7) xor crcCur(11) xor crcCur(12) xor crcCur(14) xor crcCur(15) xor crcCur(17) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(24) xor crcCur(26) xor crcCur(27) xor crcCur(28) xor crcCur(29);
      retVar(30) := data(4) xor data(7) xor data(8) xor data(10) xor data(14) xor data(22) xor data(23) xor data(24) xor data(26) xor data(27) xor data(28) xor data(29) xor data(30) xor data(32) xor data(35) xor data(42) xor data(43) xor data(45) xor data(46) xor data(48) xor data(51) xor data(52) xor data(53) xor data(56) xor data(58) xor data(59) xor data(61) xor data(63) xor data(64) xor data(65) xor data(66) xor data(70) xor data(71) xor data(77) xor data(79) xor data(80) xor data(81) xor data(82) xor data(83) xor data(85) xor data(92) xor data(93) xor data(94) xor data(95) xor data(96) xor data(97) xor data(99) xor data(101) xor data(102) xor data(104) xor data(108) xor data(109) xor data(111) xor data(112) xor data(114) xor data(115) xor data(116) xor data(117) xor data(121) xor data(123) xor data(124) xor data(125) xor data(126) xor crcCur(0) xor crcCur(1) xor crcCur(3) xor crcCur(5) xor crcCur(6) xor crcCur(8) xor crcCur(12) xor crcCur(13) xor crcCur(15) xor crcCur(16) xor crcCur(18) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(25) xor crcCur(27) xor crcCur(28) xor crcCur(29) xor crcCur(30);
      retVar(31) := data(5) xor data(8) xor data(9) xor data(11) xor data(15) xor data(23) xor data(24) xor data(25) xor data(27) xor data(28) xor data(29) xor data(30) xor data(31) xor data(33) xor data(36) xor data(43) xor data(44) xor data(46) xor data(47) xor data(49) xor data(52) xor data(53) xor data(54) xor data(57) xor data(59) xor data(60) xor data(62) xor data(64) xor data(65) xor data(66) xor data(67) xor data(71) xor data(72) xor data(78) xor data(80) xor data(81) xor data(82) xor data(83) xor data(84) xor data(86) xor data(93) xor data(94) xor data(95) xor data(96) xor data(97) xor data(98) xor data(100) xor data(102) xor data(103) xor data(105) xor data(109) xor data(110) xor data(112) xor data(113) xor data(115) xor data(116) xor data(117) xor data(118) xor data(122) xor data(124) xor data(125) xor data(126) xor data(127) xor crcCur(0) xor crcCur(1) xor crcCur(2) xor crcCur(4) xor crcCur(6) xor crcCur(7) xor crcCur(9) xor crcCur(13) xor crcCur(14) xor crcCur(16) xor crcCur(17) xor crcCur(19) xor crcCur(20) xor crcCur(21) xor crcCur(22) xor crcCur(26) xor crcCur(28) xor crcCur(29) xor crcCur(30) xor crcCur(31);
      return retVar;
   end function;

   procedure xorBitMap1Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(7 downto 0)) is 
   begin
      xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(88) := previousCrc(24); xorBitMap(0)(94) := previousCrc(30); 
      xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(88) := previousCrc(24); xorBitMap(1)(89) := previousCrc(25); xorBitMap(1)(94) := previousCrc(30); xorBitMap(1)(95) := previousCrc(31); 
      xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(88) := previousCrc(24); xorBitMap(2)(89) := previousCrc(25); xorBitMap(2)(90) := previousCrc(26); xorBitMap(2)(94) := previousCrc(30); xorBitMap(2)(95) := previousCrc(31); 
      xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(89) := previousCrc(25); xorBitMap(3)(90) := previousCrc(26); xorBitMap(3)(91) := previousCrc(27); xorBitMap(3)(95) := previousCrc(31); 
      xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(88) := previousCrc(24); xorBitMap(4)(90) := previousCrc(26); xorBitMap(4)(91) := previousCrc(27); xorBitMap(4)(92) := previousCrc(28); xorBitMap(4)(94) := previousCrc(30); 
      xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(88) := previousCrc(24); xorBitMap(5)(89) := previousCrc(25); xorBitMap(5)(91) := previousCrc(27); xorBitMap(5)(92) := previousCrc(28); xorBitMap(5)(93) := previousCrc(29); xorBitMap(5)(94) := previousCrc(30); xorBitMap(5)(95) := previousCrc(31); 
      xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(89) := previousCrc(25); xorBitMap(6)(90) := previousCrc(26); xorBitMap(6)(92) := previousCrc(28); xorBitMap(6)(93) := previousCrc(29); xorBitMap(6)(94) := previousCrc(30); xorBitMap(6)(95) := previousCrc(31); 
      xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(88) := previousCrc(24); xorBitMap(7)(90) := previousCrc(26); xorBitMap(7)(91) := previousCrc(27); xorBitMap(7)(93) := previousCrc(29); xorBitMap(7)(95) := previousCrc(31); 
      xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(64) := previousCrc(0); xorBitMap(8)(88) := previousCrc(24); xorBitMap(8)(89) := previousCrc(25); xorBitMap(8)(91) := previousCrc(27); xorBitMap(8)(92) := previousCrc(28); 
      xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(65) := previousCrc(1); xorBitMap(9)(89) := previousCrc(25); xorBitMap(9)(90) := previousCrc(26); xorBitMap(9)(92) := previousCrc(28); xorBitMap(9)(93) := previousCrc(29); 
      xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(66) := previousCrc(2); xorBitMap(10)(88) := previousCrc(24); xorBitMap(10)(90) := previousCrc(26); xorBitMap(10)(91) := previousCrc(27); xorBitMap(10)(93) := previousCrc(29); 
      xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(67) := previousCrc(3); xorBitMap(11)(88) := previousCrc(24); xorBitMap(11)(89) := previousCrc(25); xorBitMap(11)(91) := previousCrc(27); xorBitMap(11)(92) := previousCrc(28); 
      xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(68) := previousCrc(4); xorBitMap(12)(88) := previousCrc(24); xorBitMap(12)(89) := previousCrc(25); xorBitMap(12)(90) := previousCrc(26); xorBitMap(12)(92) := previousCrc(28); xorBitMap(12)(93) := previousCrc(29); xorBitMap(12)(94) := previousCrc(30); 
      xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(69) := previousCrc(5); xorBitMap(13)(89) := previousCrc(25); xorBitMap(13)(90) := previousCrc(26); xorBitMap(13)(91) := previousCrc(27); xorBitMap(13)(93) := previousCrc(29); xorBitMap(13)(94) := previousCrc(30); xorBitMap(13)(95) := previousCrc(31); 
      xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(70) := previousCrc(6); xorBitMap(14)(90) := previousCrc(26); xorBitMap(14)(91) := previousCrc(27); xorBitMap(14)(92) := previousCrc(28); xorBitMap(14)(94) := previousCrc(30); xorBitMap(14)(95) := previousCrc(31); 
      xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(71) := previousCrc(7); xorBitMap(15)(91) := previousCrc(27); xorBitMap(15)(92) := previousCrc(28); xorBitMap(15)(93) := previousCrc(29); xorBitMap(15)(95) := previousCrc(31); 
      xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(72) := previousCrc(8); xorBitMap(16)(88) := previousCrc(24); xorBitMap(16)(92) := previousCrc(28); xorBitMap(16)(93) := previousCrc(29); 
      xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(73) := previousCrc(9); xorBitMap(17)(89) := previousCrc(25); xorBitMap(17)(93) := previousCrc(29); xorBitMap(17)(94) := previousCrc(30); 
      xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(74) := previousCrc(10); xorBitMap(18)(90) := previousCrc(26); xorBitMap(18)(94) := previousCrc(30); xorBitMap(18)(95) := previousCrc(31); 
      xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(75) := previousCrc(11); xorBitMap(19)(91) := previousCrc(27); xorBitMap(19)(95) := previousCrc(31); 
      xorBitMap(20)(4) := currentData(4); xorBitMap(20)(76) := previousCrc(12); xorBitMap(20)(92) := previousCrc(28); 
      xorBitMap(21)(5) := currentData(5); xorBitMap(21)(77) := previousCrc(13); xorBitMap(21)(93) := previousCrc(29); 
      xorBitMap(22)(0) := currentData(0); xorBitMap(22)(78) := previousCrc(14); xorBitMap(22)(88) := previousCrc(24); 
      xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(79) := previousCrc(15); xorBitMap(23)(88) := previousCrc(24); xorBitMap(23)(89) := previousCrc(25); xorBitMap(23)(94) := previousCrc(30); 
      xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(80) := previousCrc(16); xorBitMap(24)(89) := previousCrc(25); xorBitMap(24)(90) := previousCrc(26); xorBitMap(24)(95) := previousCrc(31); 
      xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(81) := previousCrc(17); xorBitMap(25)(90) := previousCrc(26); xorBitMap(25)(91) := previousCrc(27); 
      xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(82) := previousCrc(18); xorBitMap(26)(88) := previousCrc(24); xorBitMap(26)(91) := previousCrc(27); xorBitMap(26)(92) := previousCrc(28); xorBitMap(26)(94) := previousCrc(30); 
      xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(83) := previousCrc(19); xorBitMap(27)(89) := previousCrc(25); xorBitMap(27)(92) := previousCrc(28); xorBitMap(27)(93) := previousCrc(29); xorBitMap(27)(95) := previousCrc(31); 
      xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(84) := previousCrc(20); xorBitMap(28)(90) := previousCrc(26); xorBitMap(28)(93) := previousCrc(29); xorBitMap(28)(94) := previousCrc(30); 
      xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(85) := previousCrc(21); xorBitMap(29)(91) := previousCrc(27); xorBitMap(29)(94) := previousCrc(30); xorBitMap(29)(95) := previousCrc(31); 
      xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(86) := previousCrc(22); xorBitMap(30)(92) := previousCrc(28); xorBitMap(30)(95) := previousCrc(31); 
      xorBitMap(31)(5) := currentData(5); xorBitMap(31)(87) := previousCrc(23); xorBitMap(31)(93) := previousCrc(29); 
   end procedure;

   procedure xorBitMap2Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(15 downto 0)) is 
   begin
      xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(80) := previousCrc(16); xorBitMap(0)(86) := previousCrc(22); xorBitMap(0)(89) := previousCrc(25); xorBitMap(0)(90) := previousCrc(26); xorBitMap(0)(92) := previousCrc(28); 
      xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(80) := previousCrc(16); xorBitMap(1)(81) := previousCrc(17); xorBitMap(1)(86) := previousCrc(22); xorBitMap(1)(87) := previousCrc(23); xorBitMap(1)(89) := previousCrc(25); xorBitMap(1)(91) := previousCrc(27); xorBitMap(1)(92) := previousCrc(28); xorBitMap(1)(93) := previousCrc(29); 
      xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(80) := previousCrc(16); xorBitMap(2)(81) := previousCrc(17); xorBitMap(2)(82) := previousCrc(18); xorBitMap(2)(86) := previousCrc(22); xorBitMap(2)(87) := previousCrc(23); xorBitMap(2)(88) := previousCrc(24); xorBitMap(2)(89) := previousCrc(25); xorBitMap(2)(93) := previousCrc(29); xorBitMap(2)(94) := previousCrc(30); 
      xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(81) := previousCrc(17); xorBitMap(3)(82) := previousCrc(18); xorBitMap(3)(83) := previousCrc(19); xorBitMap(3)(87) := previousCrc(23); xorBitMap(3)(88) := previousCrc(24); xorBitMap(3)(89) := previousCrc(25); xorBitMap(3)(90) := previousCrc(26); xorBitMap(3)(94) := previousCrc(30); xorBitMap(3)(95) := previousCrc(31); 
      xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(80) := previousCrc(16); xorBitMap(4)(82) := previousCrc(18); xorBitMap(4)(83) := previousCrc(19); xorBitMap(4)(84) := previousCrc(20); xorBitMap(4)(86) := previousCrc(22); xorBitMap(4)(88) := previousCrc(24); xorBitMap(4)(91) := previousCrc(27); xorBitMap(4)(92) := previousCrc(28); xorBitMap(4)(95) := previousCrc(31); 
      xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(80) := previousCrc(16); xorBitMap(5)(81) := previousCrc(17); xorBitMap(5)(83) := previousCrc(19); xorBitMap(5)(84) := previousCrc(20); xorBitMap(5)(85) := previousCrc(21); xorBitMap(5)(86) := previousCrc(22); xorBitMap(5)(87) := previousCrc(23); xorBitMap(5)(90) := previousCrc(26); xorBitMap(5)(93) := previousCrc(29); 
      xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(81) := previousCrc(17); xorBitMap(6)(82) := previousCrc(18); xorBitMap(6)(84) := previousCrc(20); xorBitMap(6)(85) := previousCrc(21); xorBitMap(6)(86) := previousCrc(22); xorBitMap(6)(87) := previousCrc(23); xorBitMap(6)(88) := previousCrc(24); xorBitMap(6)(91) := previousCrc(27); xorBitMap(6)(94) := previousCrc(30); 
      xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(80) := previousCrc(16); xorBitMap(7)(82) := previousCrc(18); xorBitMap(7)(83) := previousCrc(19); xorBitMap(7)(85) := previousCrc(21); xorBitMap(7)(87) := previousCrc(23); xorBitMap(7)(88) := previousCrc(24); xorBitMap(7)(90) := previousCrc(26); xorBitMap(7)(95) := previousCrc(31); 
      xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(80) := previousCrc(16); xorBitMap(8)(81) := previousCrc(17); xorBitMap(8)(83) := previousCrc(19); xorBitMap(8)(84) := previousCrc(20); xorBitMap(8)(88) := previousCrc(24); xorBitMap(8)(90) := previousCrc(26); xorBitMap(8)(91) := previousCrc(27); xorBitMap(8)(92) := previousCrc(28); 
      xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(81) := previousCrc(17); xorBitMap(9)(82) := previousCrc(18); xorBitMap(9)(84) := previousCrc(20); xorBitMap(9)(85) := previousCrc(21); xorBitMap(9)(89) := previousCrc(25); xorBitMap(9)(91) := previousCrc(27); xorBitMap(9)(92) := previousCrc(28); xorBitMap(9)(93) := previousCrc(29); 
      xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(80) := previousCrc(16); xorBitMap(10)(82) := previousCrc(18); xorBitMap(10)(83) := previousCrc(19); xorBitMap(10)(85) := previousCrc(21); xorBitMap(10)(89) := previousCrc(25); xorBitMap(10)(93) := previousCrc(29); xorBitMap(10)(94) := previousCrc(30); 
      xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(80) := previousCrc(16); xorBitMap(11)(81) := previousCrc(17); xorBitMap(11)(83) := previousCrc(19); xorBitMap(11)(84) := previousCrc(20); xorBitMap(11)(89) := previousCrc(25); xorBitMap(11)(92) := previousCrc(28); xorBitMap(11)(94) := previousCrc(30); xorBitMap(11)(95) := previousCrc(31); 
      xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(80) := previousCrc(16); xorBitMap(12)(81) := previousCrc(17); xorBitMap(12)(82) := previousCrc(18); xorBitMap(12)(84) := previousCrc(20); xorBitMap(12)(85) := previousCrc(21); xorBitMap(12)(86) := previousCrc(22); xorBitMap(12)(89) := previousCrc(25); xorBitMap(12)(92) := previousCrc(28); xorBitMap(12)(93) := previousCrc(29); xorBitMap(12)(95) := previousCrc(31); 
      xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(81) := previousCrc(17); xorBitMap(13)(82) := previousCrc(18); xorBitMap(13)(83) := previousCrc(19); xorBitMap(13)(85) := previousCrc(21); xorBitMap(13)(86) := previousCrc(22); xorBitMap(13)(87) := previousCrc(23); xorBitMap(13)(90) := previousCrc(26); xorBitMap(13)(93) := previousCrc(29); xorBitMap(13)(94) := previousCrc(30); 
      xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(82) := previousCrc(18); xorBitMap(14)(83) := previousCrc(19); xorBitMap(14)(84) := previousCrc(20); xorBitMap(14)(86) := previousCrc(22); xorBitMap(14)(87) := previousCrc(23); xorBitMap(14)(88) := previousCrc(24); xorBitMap(14)(91) := previousCrc(27); xorBitMap(14)(94) := previousCrc(30); xorBitMap(14)(95) := previousCrc(31); 
      xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(83) := previousCrc(19); xorBitMap(15)(84) := previousCrc(20); xorBitMap(15)(85) := previousCrc(21); xorBitMap(15)(87) := previousCrc(23); xorBitMap(15)(88) := previousCrc(24); xorBitMap(15)(89) := previousCrc(25); xorBitMap(15)(92) := previousCrc(28); xorBitMap(15)(95) := previousCrc(31); 
      xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(64) := previousCrc(0); xorBitMap(16)(80) := previousCrc(16); xorBitMap(16)(84) := previousCrc(20); xorBitMap(16)(85) := previousCrc(21); xorBitMap(16)(88) := previousCrc(24); xorBitMap(16)(92) := previousCrc(28); xorBitMap(16)(93) := previousCrc(29); 
      xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(65) := previousCrc(1); xorBitMap(17)(81) := previousCrc(17); xorBitMap(17)(85) := previousCrc(21); xorBitMap(17)(86) := previousCrc(22); xorBitMap(17)(89) := previousCrc(25); xorBitMap(17)(93) := previousCrc(29); xorBitMap(17)(94) := previousCrc(30); 
      xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(66) := previousCrc(2); xorBitMap(18)(82) := previousCrc(18); xorBitMap(18)(86) := previousCrc(22); xorBitMap(18)(87) := previousCrc(23); xorBitMap(18)(90) := previousCrc(26); xorBitMap(18)(94) := previousCrc(30); xorBitMap(18)(95) := previousCrc(31); 
      xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(67) := previousCrc(3); xorBitMap(19)(83) := previousCrc(19); xorBitMap(19)(87) := previousCrc(23); xorBitMap(19)(88) := previousCrc(24); xorBitMap(19)(91) := previousCrc(27); xorBitMap(19)(95) := previousCrc(31); 
      xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(68) := previousCrc(4); xorBitMap(20)(84) := previousCrc(20); xorBitMap(20)(88) := previousCrc(24); xorBitMap(20)(89) := previousCrc(25); xorBitMap(20)(92) := previousCrc(28); 
      xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(69) := previousCrc(5); xorBitMap(21)(85) := previousCrc(21); xorBitMap(21)(89) := previousCrc(25); xorBitMap(21)(90) := previousCrc(26); xorBitMap(21)(93) := previousCrc(29); 
      xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(70) := previousCrc(6); xorBitMap(22)(80) := previousCrc(16); xorBitMap(22)(89) := previousCrc(25); xorBitMap(22)(91) := previousCrc(27); xorBitMap(22)(92) := previousCrc(28); xorBitMap(22)(94) := previousCrc(30); 
      xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(71) := previousCrc(7); xorBitMap(23)(80) := previousCrc(16); xorBitMap(23)(81) := previousCrc(17); xorBitMap(23)(86) := previousCrc(22); xorBitMap(23)(89) := previousCrc(25); xorBitMap(23)(93) := previousCrc(29); xorBitMap(23)(95) := previousCrc(31); 
      xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(72) := previousCrc(8); xorBitMap(24)(81) := previousCrc(17); xorBitMap(24)(82) := previousCrc(18); xorBitMap(24)(87) := previousCrc(23); xorBitMap(24)(90) := previousCrc(26); xorBitMap(24)(94) := previousCrc(30); 
      xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(73) := previousCrc(9); xorBitMap(25)(82) := previousCrc(18); xorBitMap(25)(83) := previousCrc(19); xorBitMap(25)(88) := previousCrc(24); xorBitMap(25)(91) := previousCrc(27); xorBitMap(25)(95) := previousCrc(31); 
      xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(74) := previousCrc(10); xorBitMap(26)(80) := previousCrc(16); xorBitMap(26)(83) := previousCrc(19); xorBitMap(26)(84) := previousCrc(20); xorBitMap(26)(86) := previousCrc(22); xorBitMap(26)(90) := previousCrc(26); 
      xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(75) := previousCrc(11); xorBitMap(27)(81) := previousCrc(17); xorBitMap(27)(84) := previousCrc(20); xorBitMap(27)(85) := previousCrc(21); xorBitMap(27)(87) := previousCrc(23); xorBitMap(27)(91) := previousCrc(27); 
      xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(76) := previousCrc(12); xorBitMap(28)(82) := previousCrc(18); xorBitMap(28)(85) := previousCrc(21); xorBitMap(28)(86) := previousCrc(22); xorBitMap(28)(88) := previousCrc(24); xorBitMap(28)(92) := previousCrc(28); 
      xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(77) := previousCrc(13); xorBitMap(29)(83) := previousCrc(19); xorBitMap(29)(86) := previousCrc(22); xorBitMap(29)(87) := previousCrc(23); xorBitMap(29)(89) := previousCrc(25); xorBitMap(29)(93) := previousCrc(29); 
      xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(78) := previousCrc(14); xorBitMap(30)(84) := previousCrc(20); xorBitMap(30)(87) := previousCrc(23); xorBitMap(30)(88) := previousCrc(24); xorBitMap(30)(90) := previousCrc(26); xorBitMap(30)(94) := previousCrc(30); 
      xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(79) := previousCrc(15); xorBitMap(31)(85) := previousCrc(21); xorBitMap(31)(88) := previousCrc(24); xorBitMap(31)(89) := previousCrc(25); xorBitMap(31)(91) := previousCrc(27); xorBitMap(31)(95) := previousCrc(31); 
   end procedure;

   procedure xorBitMap3Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(23 downto 0)) is 
   begin
      xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(72) := previousCrc(8); xorBitMap(0)(78) := previousCrc(14); xorBitMap(0)(81) := previousCrc(17); xorBitMap(0)(82) := previousCrc(18); xorBitMap(0)(84) := previousCrc(20); xorBitMap(0)(88) := previousCrc(24); 
      xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(72) := previousCrc(8); xorBitMap(1)(73) := previousCrc(9); xorBitMap(1)(78) := previousCrc(14); xorBitMap(1)(79) := previousCrc(15); xorBitMap(1)(81) := previousCrc(17); xorBitMap(1)(83) := previousCrc(19); xorBitMap(1)(84) := previousCrc(20); xorBitMap(1)(85) := previousCrc(21); xorBitMap(1)(88) := previousCrc(24); xorBitMap(1)(89) := previousCrc(25); 
      xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(72) := previousCrc(8); xorBitMap(2)(73) := previousCrc(9); xorBitMap(2)(74) := previousCrc(10); xorBitMap(2)(78) := previousCrc(14); xorBitMap(2)(79) := previousCrc(15); xorBitMap(2)(80) := previousCrc(16); xorBitMap(2)(81) := previousCrc(17); xorBitMap(2)(85) := previousCrc(21); xorBitMap(2)(86) := previousCrc(22); xorBitMap(2)(88) := previousCrc(24); xorBitMap(2)(89) := previousCrc(25); xorBitMap(2)(90) := previousCrc(26); 
      xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(73) := previousCrc(9); xorBitMap(3)(74) := previousCrc(10); xorBitMap(3)(75) := previousCrc(11); xorBitMap(3)(79) := previousCrc(15); xorBitMap(3)(80) := previousCrc(16); xorBitMap(3)(81) := previousCrc(17); xorBitMap(3)(82) := previousCrc(18); xorBitMap(3)(86) := previousCrc(22); xorBitMap(3)(87) := previousCrc(23); xorBitMap(3)(89) := previousCrc(25); xorBitMap(3)(90) := previousCrc(26); xorBitMap(3)(91) := previousCrc(27); 
      xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(72) := previousCrc(8); xorBitMap(4)(74) := previousCrc(10); xorBitMap(4)(75) := previousCrc(11); xorBitMap(4)(76) := previousCrc(12); xorBitMap(4)(78) := previousCrc(14); xorBitMap(4)(80) := previousCrc(16); xorBitMap(4)(83) := previousCrc(19); xorBitMap(4)(84) := previousCrc(20); xorBitMap(4)(87) := previousCrc(23); xorBitMap(4)(90) := previousCrc(26); xorBitMap(4)(91) := previousCrc(27); xorBitMap(4)(92) := previousCrc(28); 
      xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(72) := previousCrc(8); xorBitMap(5)(73) := previousCrc(9); xorBitMap(5)(75) := previousCrc(11); xorBitMap(5)(76) := previousCrc(12); xorBitMap(5)(77) := previousCrc(13); xorBitMap(5)(78) := previousCrc(14); xorBitMap(5)(79) := previousCrc(15); xorBitMap(5)(82) := previousCrc(18); xorBitMap(5)(85) := previousCrc(21); xorBitMap(5)(91) := previousCrc(27); xorBitMap(5)(92) := previousCrc(28); xorBitMap(5)(93) := previousCrc(29); 
      xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(73) := previousCrc(9); xorBitMap(6)(74) := previousCrc(10); xorBitMap(6)(76) := previousCrc(12); xorBitMap(6)(77) := previousCrc(13); xorBitMap(6)(78) := previousCrc(14); xorBitMap(6)(79) := previousCrc(15); xorBitMap(6)(80) := previousCrc(16); xorBitMap(6)(83) := previousCrc(19); xorBitMap(6)(86) := previousCrc(22); xorBitMap(6)(92) := previousCrc(28); xorBitMap(6)(93) := previousCrc(29); xorBitMap(6)(94) := previousCrc(30); 
      xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(72) := previousCrc(8); xorBitMap(7)(74) := previousCrc(10); xorBitMap(7)(75) := previousCrc(11); xorBitMap(7)(77) := previousCrc(13); xorBitMap(7)(79) := previousCrc(15); xorBitMap(7)(80) := previousCrc(16); xorBitMap(7)(82) := previousCrc(18); xorBitMap(7)(87) := previousCrc(23); xorBitMap(7)(88) := previousCrc(24); xorBitMap(7)(93) := previousCrc(29); xorBitMap(7)(94) := previousCrc(30); xorBitMap(7)(95) := previousCrc(31); 
      xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(72) := previousCrc(8); xorBitMap(8)(73) := previousCrc(9); xorBitMap(8)(75) := previousCrc(11); xorBitMap(8)(76) := previousCrc(12); xorBitMap(8)(80) := previousCrc(16); xorBitMap(8)(82) := previousCrc(18); xorBitMap(8)(83) := previousCrc(19); xorBitMap(8)(84) := previousCrc(20); xorBitMap(8)(89) := previousCrc(25); xorBitMap(8)(94) := previousCrc(30); xorBitMap(8)(95) := previousCrc(31); 
      xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(73) := previousCrc(9); xorBitMap(9)(74) := previousCrc(10); xorBitMap(9)(76) := previousCrc(12); xorBitMap(9)(77) := previousCrc(13); xorBitMap(9)(81) := previousCrc(17); xorBitMap(9)(83) := previousCrc(19); xorBitMap(9)(84) := previousCrc(20); xorBitMap(9)(85) := previousCrc(21); xorBitMap(9)(90) := previousCrc(26); xorBitMap(9)(95) := previousCrc(31); 
      xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(72) := previousCrc(8); xorBitMap(10)(74) := previousCrc(10); xorBitMap(10)(75) := previousCrc(11); xorBitMap(10)(77) := previousCrc(13); xorBitMap(10)(81) := previousCrc(17); xorBitMap(10)(85) := previousCrc(21); xorBitMap(10)(86) := previousCrc(22); xorBitMap(10)(88) := previousCrc(24); xorBitMap(10)(91) := previousCrc(27); 
      xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(72) := previousCrc(8); xorBitMap(11)(73) := previousCrc(9); xorBitMap(11)(75) := previousCrc(11); xorBitMap(11)(76) := previousCrc(12); xorBitMap(11)(81) := previousCrc(17); xorBitMap(11)(84) := previousCrc(20); xorBitMap(11)(86) := previousCrc(22); xorBitMap(11)(87) := previousCrc(23); xorBitMap(11)(88) := previousCrc(24); xorBitMap(11)(89) := previousCrc(25); xorBitMap(11)(92) := previousCrc(28); 
      xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(72) := previousCrc(8); xorBitMap(12)(73) := previousCrc(9); xorBitMap(12)(74) := previousCrc(10); xorBitMap(12)(76) := previousCrc(12); xorBitMap(12)(77) := previousCrc(13); xorBitMap(12)(78) := previousCrc(14); xorBitMap(12)(81) := previousCrc(17); xorBitMap(12)(84) := previousCrc(20); xorBitMap(12)(85) := previousCrc(21); xorBitMap(12)(87) := previousCrc(23); xorBitMap(12)(89) := previousCrc(25); xorBitMap(12)(90) := previousCrc(26); xorBitMap(12)(93) := previousCrc(29); 
      xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(73) := previousCrc(9); xorBitMap(13)(74) := previousCrc(10); xorBitMap(13)(75) := previousCrc(11); xorBitMap(13)(77) := previousCrc(13); xorBitMap(13)(78) := previousCrc(14); xorBitMap(13)(79) := previousCrc(15); xorBitMap(13)(82) := previousCrc(18); xorBitMap(13)(85) := previousCrc(21); xorBitMap(13)(86) := previousCrc(22); xorBitMap(13)(88) := previousCrc(24); xorBitMap(13)(90) := previousCrc(26); xorBitMap(13)(91) := previousCrc(27); xorBitMap(13)(94) := previousCrc(30); 
      xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(74) := previousCrc(10); xorBitMap(14)(75) := previousCrc(11); xorBitMap(14)(76) := previousCrc(12); xorBitMap(14)(78) := previousCrc(14); xorBitMap(14)(79) := previousCrc(15); xorBitMap(14)(80) := previousCrc(16); xorBitMap(14)(83) := previousCrc(19); xorBitMap(14)(86) := previousCrc(22); xorBitMap(14)(87) := previousCrc(23); xorBitMap(14)(89) := previousCrc(25); xorBitMap(14)(91) := previousCrc(27); xorBitMap(14)(92) := previousCrc(28); xorBitMap(14)(95) := previousCrc(31); 
      xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(75) := previousCrc(11); xorBitMap(15)(76) := previousCrc(12); xorBitMap(15)(77) := previousCrc(13); xorBitMap(15)(79) := previousCrc(15); xorBitMap(15)(80) := previousCrc(16); xorBitMap(15)(81) := previousCrc(17); xorBitMap(15)(84) := previousCrc(20); xorBitMap(15)(87) := previousCrc(23); xorBitMap(15)(88) := previousCrc(24); xorBitMap(15)(90) := previousCrc(26); xorBitMap(15)(92) := previousCrc(28); xorBitMap(15)(93) := previousCrc(29); 
      xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(72) := previousCrc(8); xorBitMap(16)(76) := previousCrc(12); xorBitMap(16)(77) := previousCrc(13); xorBitMap(16)(80) := previousCrc(16); xorBitMap(16)(84) := previousCrc(20); xorBitMap(16)(85) := previousCrc(21); xorBitMap(16)(89) := previousCrc(25); xorBitMap(16)(91) := previousCrc(27); xorBitMap(16)(93) := previousCrc(29); xorBitMap(16)(94) := previousCrc(30); 
      xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(73) := previousCrc(9); xorBitMap(17)(77) := previousCrc(13); xorBitMap(17)(78) := previousCrc(14); xorBitMap(17)(81) := previousCrc(17); xorBitMap(17)(85) := previousCrc(21); xorBitMap(17)(86) := previousCrc(22); xorBitMap(17)(90) := previousCrc(26); xorBitMap(17)(92) := previousCrc(28); xorBitMap(17)(94) := previousCrc(30); xorBitMap(17)(95) := previousCrc(31); 
      xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(74) := previousCrc(10); xorBitMap(18)(78) := previousCrc(14); xorBitMap(18)(79) := previousCrc(15); xorBitMap(18)(82) := previousCrc(18); xorBitMap(18)(86) := previousCrc(22); xorBitMap(18)(87) := previousCrc(23); xorBitMap(18)(91) := previousCrc(27); xorBitMap(18)(93) := previousCrc(29); xorBitMap(18)(95) := previousCrc(31); 
      xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(75) := previousCrc(11); xorBitMap(19)(79) := previousCrc(15); xorBitMap(19)(80) := previousCrc(16); xorBitMap(19)(83) := previousCrc(19); xorBitMap(19)(87) := previousCrc(23); xorBitMap(19)(88) := previousCrc(24); xorBitMap(19)(92) := previousCrc(28); xorBitMap(19)(94) := previousCrc(30); 
      xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(76) := previousCrc(12); xorBitMap(20)(80) := previousCrc(16); xorBitMap(20)(81) := previousCrc(17); xorBitMap(20)(84) := previousCrc(20); xorBitMap(20)(88) := previousCrc(24); xorBitMap(20)(89) := previousCrc(25); xorBitMap(20)(93) := previousCrc(29); xorBitMap(20)(95) := previousCrc(31); 
      xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(77) := previousCrc(13); xorBitMap(21)(81) := previousCrc(17); xorBitMap(21)(82) := previousCrc(18); xorBitMap(21)(85) := previousCrc(21); xorBitMap(21)(89) := previousCrc(25); xorBitMap(21)(90) := previousCrc(26); xorBitMap(21)(94) := previousCrc(30); 
      xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(72) := previousCrc(8); xorBitMap(22)(81) := previousCrc(17); xorBitMap(22)(83) := previousCrc(19); xorBitMap(22)(84) := previousCrc(20); xorBitMap(22)(86) := previousCrc(22); xorBitMap(22)(88) := previousCrc(24); xorBitMap(22)(90) := previousCrc(26); xorBitMap(22)(91) := previousCrc(27); xorBitMap(22)(95) := previousCrc(31); 
      xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(72) := previousCrc(8); xorBitMap(23)(73) := previousCrc(9); xorBitMap(23)(78) := previousCrc(14); xorBitMap(23)(81) := previousCrc(17); xorBitMap(23)(85) := previousCrc(21); xorBitMap(23)(87) := previousCrc(23); xorBitMap(23)(88) := previousCrc(24); xorBitMap(23)(89) := previousCrc(25); xorBitMap(23)(91) := previousCrc(27); xorBitMap(23)(92) := previousCrc(28); 
      xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(64) := previousCrc(0); xorBitMap(24)(73) := previousCrc(9); xorBitMap(24)(74) := previousCrc(10); xorBitMap(24)(79) := previousCrc(15); xorBitMap(24)(82) := previousCrc(18); xorBitMap(24)(86) := previousCrc(22); xorBitMap(24)(88) := previousCrc(24); xorBitMap(24)(89) := previousCrc(25); xorBitMap(24)(90) := previousCrc(26); xorBitMap(24)(92) := previousCrc(28); xorBitMap(24)(93) := previousCrc(29); 
      xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(65) := previousCrc(1); xorBitMap(25)(74) := previousCrc(10); xorBitMap(25)(75) := previousCrc(11); xorBitMap(25)(80) := previousCrc(16); xorBitMap(25)(83) := previousCrc(19); xorBitMap(25)(87) := previousCrc(23); xorBitMap(25)(89) := previousCrc(25); xorBitMap(25)(90) := previousCrc(26); xorBitMap(25)(91) := previousCrc(27); xorBitMap(25)(93) := previousCrc(29); xorBitMap(25)(94) := previousCrc(30); 
      xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(66) := previousCrc(2); xorBitMap(26)(72) := previousCrc(8); xorBitMap(26)(75) := previousCrc(11); xorBitMap(26)(76) := previousCrc(12); xorBitMap(26)(78) := previousCrc(14); xorBitMap(26)(82) := previousCrc(18); xorBitMap(26)(90) := previousCrc(26); xorBitMap(26)(91) := previousCrc(27); xorBitMap(26)(92) := previousCrc(28); xorBitMap(26)(94) := previousCrc(30); xorBitMap(26)(95) := previousCrc(31); 
      xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(67) := previousCrc(3); xorBitMap(27)(73) := previousCrc(9); xorBitMap(27)(76) := previousCrc(12); xorBitMap(27)(77) := previousCrc(13); xorBitMap(27)(79) := previousCrc(15); xorBitMap(27)(83) := previousCrc(19); xorBitMap(27)(91) := previousCrc(27); xorBitMap(27)(92) := previousCrc(28); xorBitMap(27)(93) := previousCrc(29); xorBitMap(27)(95) := previousCrc(31); 
      xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(68) := previousCrc(4); xorBitMap(28)(74) := previousCrc(10); xorBitMap(28)(77) := previousCrc(13); xorBitMap(28)(78) := previousCrc(14); xorBitMap(28)(80) := previousCrc(16); xorBitMap(28)(84) := previousCrc(20); xorBitMap(28)(92) := previousCrc(28); xorBitMap(28)(93) := previousCrc(29); xorBitMap(28)(94) := previousCrc(30); 
      xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(69) := previousCrc(5); xorBitMap(29)(75) := previousCrc(11); xorBitMap(29)(78) := previousCrc(14); xorBitMap(29)(79) := previousCrc(15); xorBitMap(29)(81) := previousCrc(17); xorBitMap(29)(85) := previousCrc(21); xorBitMap(29)(93) := previousCrc(29); xorBitMap(29)(94) := previousCrc(30); xorBitMap(29)(95) := previousCrc(31); 
      xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(70) := previousCrc(6); xorBitMap(30)(76) := previousCrc(12); xorBitMap(30)(79) := previousCrc(15); xorBitMap(30)(80) := previousCrc(16); xorBitMap(30)(82) := previousCrc(18); xorBitMap(30)(86) := previousCrc(22); xorBitMap(30)(94) := previousCrc(30); xorBitMap(30)(95) := previousCrc(31); 
      xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(71) := previousCrc(7); xorBitMap(31)(77) := previousCrc(13); xorBitMap(31)(80) := previousCrc(16); xorBitMap(31)(81) := previousCrc(17); xorBitMap(31)(83) := previousCrc(19); xorBitMap(31)(87) := previousCrc(23); xorBitMap(31)(95) := previousCrc(31); 
   end procedure;

   procedure xorBitMap4Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(31 downto 0)) is 
   begin
      xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(64) := previousCrc(0); xorBitMap(0)(70) := previousCrc(6); xorBitMap(0)(73) := previousCrc(9); xorBitMap(0)(74) := previousCrc(10); xorBitMap(0)(76) := previousCrc(12); xorBitMap(0)(80) := previousCrc(16); xorBitMap(0)(88) := previousCrc(24); xorBitMap(0)(89) := previousCrc(25); xorBitMap(0)(90) := previousCrc(26); xorBitMap(0)(92) := previousCrc(28); xorBitMap(0)(93) := previousCrc(29); xorBitMap(0)(94) := previousCrc(30); xorBitMap(0)(95) := previousCrc(31); 
      xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(64) := previousCrc(0); xorBitMap(1)(65) := previousCrc(1); xorBitMap(1)(70) := previousCrc(6); xorBitMap(1)(71) := previousCrc(7); xorBitMap(1)(73) := previousCrc(9); xorBitMap(1)(75) := previousCrc(11); xorBitMap(1)(76) := previousCrc(12); xorBitMap(1)(77) := previousCrc(13); xorBitMap(1)(80) := previousCrc(16); xorBitMap(1)(81) := previousCrc(17); xorBitMap(1)(88) := previousCrc(24); xorBitMap(1)(91) := previousCrc(27); xorBitMap(1)(92) := previousCrc(28); 
      xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(64) := previousCrc(0); xorBitMap(2)(65) := previousCrc(1); xorBitMap(2)(66) := previousCrc(2); xorBitMap(2)(70) := previousCrc(6); xorBitMap(2)(71) := previousCrc(7); xorBitMap(2)(72) := previousCrc(8); xorBitMap(2)(73) := previousCrc(9); xorBitMap(2)(77) := previousCrc(13); xorBitMap(2)(78) := previousCrc(14); xorBitMap(2)(80) := previousCrc(16); xorBitMap(2)(81) := previousCrc(17); xorBitMap(2)(82) := previousCrc(18); xorBitMap(2)(88) := previousCrc(24); xorBitMap(2)(90) := previousCrc(26); xorBitMap(2)(94) := previousCrc(30); xorBitMap(2)(95) := previousCrc(31); 
      xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(65) := previousCrc(1); xorBitMap(3)(66) := previousCrc(2); xorBitMap(3)(67) := previousCrc(3); xorBitMap(3)(71) := previousCrc(7); xorBitMap(3)(72) := previousCrc(8); xorBitMap(3)(73) := previousCrc(9); xorBitMap(3)(74) := previousCrc(10); xorBitMap(3)(78) := previousCrc(14); xorBitMap(3)(79) := previousCrc(15); xorBitMap(3)(81) := previousCrc(17); xorBitMap(3)(82) := previousCrc(18); xorBitMap(3)(83) := previousCrc(19); xorBitMap(3)(89) := previousCrc(25); xorBitMap(3)(91) := previousCrc(27); xorBitMap(3)(95) := previousCrc(31); 
      xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(64) := previousCrc(0); xorBitMap(4)(66) := previousCrc(2); xorBitMap(4)(67) := previousCrc(3); xorBitMap(4)(68) := previousCrc(4); xorBitMap(4)(70) := previousCrc(6); xorBitMap(4)(72) := previousCrc(8); xorBitMap(4)(75) := previousCrc(11); xorBitMap(4)(76) := previousCrc(12); xorBitMap(4)(79) := previousCrc(15); xorBitMap(4)(82) := previousCrc(18); xorBitMap(4)(83) := previousCrc(19); xorBitMap(4)(84) := previousCrc(20); xorBitMap(4)(88) := previousCrc(24); xorBitMap(4)(89) := previousCrc(25); xorBitMap(4)(93) := previousCrc(29); xorBitMap(4)(94) := previousCrc(30); xorBitMap(4)(95) := previousCrc(31); 
      xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(64) := previousCrc(0); xorBitMap(5)(65) := previousCrc(1); xorBitMap(5)(67) := previousCrc(3); xorBitMap(5)(68) := previousCrc(4); xorBitMap(5)(69) := previousCrc(5); xorBitMap(5)(70) := previousCrc(6); xorBitMap(5)(71) := previousCrc(7); xorBitMap(5)(74) := previousCrc(10); xorBitMap(5)(77) := previousCrc(13); xorBitMap(5)(83) := previousCrc(19); xorBitMap(5)(84) := previousCrc(20); xorBitMap(5)(85) := previousCrc(21); xorBitMap(5)(88) := previousCrc(24); xorBitMap(5)(92) := previousCrc(28); xorBitMap(5)(93) := previousCrc(29); 
      xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(65) := previousCrc(1); xorBitMap(6)(66) := previousCrc(2); xorBitMap(6)(68) := previousCrc(4); xorBitMap(6)(69) := previousCrc(5); xorBitMap(6)(70) := previousCrc(6); xorBitMap(6)(71) := previousCrc(7); xorBitMap(6)(72) := previousCrc(8); xorBitMap(6)(75) := previousCrc(11); xorBitMap(6)(78) := previousCrc(14); xorBitMap(6)(84) := previousCrc(20); xorBitMap(6)(85) := previousCrc(21); xorBitMap(6)(86) := previousCrc(22); xorBitMap(6)(89) := previousCrc(25); xorBitMap(6)(93) := previousCrc(29); xorBitMap(6)(94) := previousCrc(30); 
      xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(64) := previousCrc(0); xorBitMap(7)(66) := previousCrc(2); xorBitMap(7)(67) := previousCrc(3); xorBitMap(7)(69) := previousCrc(5); xorBitMap(7)(71) := previousCrc(7); xorBitMap(7)(72) := previousCrc(8); xorBitMap(7)(74) := previousCrc(10); xorBitMap(7)(79) := previousCrc(15); xorBitMap(7)(80) := previousCrc(16); xorBitMap(7)(85) := previousCrc(21); xorBitMap(7)(86) := previousCrc(22); xorBitMap(7)(87) := previousCrc(23); xorBitMap(7)(88) := previousCrc(24); xorBitMap(7)(89) := previousCrc(25); xorBitMap(7)(92) := previousCrc(28); xorBitMap(7)(93) := previousCrc(29); 
      xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(64) := previousCrc(0); xorBitMap(8)(65) := previousCrc(1); xorBitMap(8)(67) := previousCrc(3); xorBitMap(8)(68) := previousCrc(4); xorBitMap(8)(72) := previousCrc(8); xorBitMap(8)(74) := previousCrc(10); xorBitMap(8)(75) := previousCrc(11); xorBitMap(8)(76) := previousCrc(12); xorBitMap(8)(81) := previousCrc(17); xorBitMap(8)(86) := previousCrc(22); xorBitMap(8)(87) := previousCrc(23); xorBitMap(8)(92) := previousCrc(28); xorBitMap(8)(95) := previousCrc(31); 
      xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(65) := previousCrc(1); xorBitMap(9)(66) := previousCrc(2); xorBitMap(9)(68) := previousCrc(4); xorBitMap(9)(69) := previousCrc(5); xorBitMap(9)(73) := previousCrc(9); xorBitMap(9)(75) := previousCrc(11); xorBitMap(9)(76) := previousCrc(12); xorBitMap(9)(77) := previousCrc(13); xorBitMap(9)(82) := previousCrc(18); xorBitMap(9)(87) := previousCrc(23); xorBitMap(9)(88) := previousCrc(24); xorBitMap(9)(93) := previousCrc(29); 
      xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(64) := previousCrc(0); xorBitMap(10)(66) := previousCrc(2); xorBitMap(10)(67) := previousCrc(3); xorBitMap(10)(69) := previousCrc(5); xorBitMap(10)(73) := previousCrc(9); xorBitMap(10)(77) := previousCrc(13); xorBitMap(10)(78) := previousCrc(14); xorBitMap(10)(80) := previousCrc(16); xorBitMap(10)(83) := previousCrc(19); xorBitMap(10)(90) := previousCrc(26); xorBitMap(10)(92) := previousCrc(28); xorBitMap(10)(93) := previousCrc(29); xorBitMap(10)(95) := previousCrc(31); 
      xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(64) := previousCrc(0); xorBitMap(11)(65) := previousCrc(1); xorBitMap(11)(67) := previousCrc(3); xorBitMap(11)(68) := previousCrc(4); xorBitMap(11)(73) := previousCrc(9); xorBitMap(11)(76) := previousCrc(12); xorBitMap(11)(78) := previousCrc(14); xorBitMap(11)(79) := previousCrc(15); xorBitMap(11)(80) := previousCrc(16); xorBitMap(11)(81) := previousCrc(17); xorBitMap(11)(84) := previousCrc(20); xorBitMap(11)(88) := previousCrc(24); xorBitMap(11)(89) := previousCrc(25); xorBitMap(11)(90) := previousCrc(26); xorBitMap(11)(91) := previousCrc(27); xorBitMap(11)(92) := previousCrc(28); xorBitMap(11)(95) := previousCrc(31); 
      xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(64) := previousCrc(0); xorBitMap(12)(65) := previousCrc(1); xorBitMap(12)(66) := previousCrc(2); xorBitMap(12)(68) := previousCrc(4); xorBitMap(12)(69) := previousCrc(5); xorBitMap(12)(70) := previousCrc(6); xorBitMap(12)(73) := previousCrc(9); xorBitMap(12)(76) := previousCrc(12); xorBitMap(12)(77) := previousCrc(13); xorBitMap(12)(79) := previousCrc(15); xorBitMap(12)(81) := previousCrc(17); xorBitMap(12)(82) := previousCrc(18); xorBitMap(12)(85) := previousCrc(21); xorBitMap(12)(88) := previousCrc(24); xorBitMap(12)(91) := previousCrc(27); xorBitMap(12)(94) := previousCrc(30); xorBitMap(12)(95) := previousCrc(31); 
      xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(65) := previousCrc(1); xorBitMap(13)(66) := previousCrc(2); xorBitMap(13)(67) := previousCrc(3); xorBitMap(13)(69) := previousCrc(5); xorBitMap(13)(70) := previousCrc(6); xorBitMap(13)(71) := previousCrc(7); xorBitMap(13)(74) := previousCrc(10); xorBitMap(13)(77) := previousCrc(13); xorBitMap(13)(78) := previousCrc(14); xorBitMap(13)(80) := previousCrc(16); xorBitMap(13)(82) := previousCrc(18); xorBitMap(13)(83) := previousCrc(19); xorBitMap(13)(86) := previousCrc(22); xorBitMap(13)(89) := previousCrc(25); xorBitMap(13)(92) := previousCrc(28); xorBitMap(13)(95) := previousCrc(31); 
      xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(66) := previousCrc(2); xorBitMap(14)(67) := previousCrc(3); xorBitMap(14)(68) := previousCrc(4); xorBitMap(14)(70) := previousCrc(6); xorBitMap(14)(71) := previousCrc(7); xorBitMap(14)(72) := previousCrc(8); xorBitMap(14)(75) := previousCrc(11); xorBitMap(14)(78) := previousCrc(14); xorBitMap(14)(79) := previousCrc(15); xorBitMap(14)(81) := previousCrc(17); xorBitMap(14)(83) := previousCrc(19); xorBitMap(14)(84) := previousCrc(20); xorBitMap(14)(87) := previousCrc(23); xorBitMap(14)(90) := previousCrc(26); xorBitMap(14)(93) := previousCrc(29); 
      xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(67) := previousCrc(3); xorBitMap(15)(68) := previousCrc(4); xorBitMap(15)(69) := previousCrc(5); xorBitMap(15)(71) := previousCrc(7); xorBitMap(15)(72) := previousCrc(8); xorBitMap(15)(73) := previousCrc(9); xorBitMap(15)(76) := previousCrc(12); xorBitMap(15)(79) := previousCrc(15); xorBitMap(15)(80) := previousCrc(16); xorBitMap(15)(82) := previousCrc(18); xorBitMap(15)(84) := previousCrc(20); xorBitMap(15)(85) := previousCrc(21); xorBitMap(15)(88) := previousCrc(24); xorBitMap(15)(91) := previousCrc(27); xorBitMap(15)(94) := previousCrc(30); 
      xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(64) := previousCrc(0); xorBitMap(16)(68) := previousCrc(4); xorBitMap(16)(69) := previousCrc(5); xorBitMap(16)(72) := previousCrc(8); xorBitMap(16)(76) := previousCrc(12); xorBitMap(16)(77) := previousCrc(13); xorBitMap(16)(81) := previousCrc(17); xorBitMap(16)(83) := previousCrc(19); xorBitMap(16)(85) := previousCrc(21); xorBitMap(16)(86) := previousCrc(22); xorBitMap(16)(88) := previousCrc(24); xorBitMap(16)(90) := previousCrc(26); xorBitMap(16)(93) := previousCrc(29); xorBitMap(16)(94) := previousCrc(30); 
      xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(65) := previousCrc(1); xorBitMap(17)(69) := previousCrc(5); xorBitMap(17)(70) := previousCrc(6); xorBitMap(17)(73) := previousCrc(9); xorBitMap(17)(77) := previousCrc(13); xorBitMap(17)(78) := previousCrc(14); xorBitMap(17)(82) := previousCrc(18); xorBitMap(17)(84) := previousCrc(20); xorBitMap(17)(86) := previousCrc(22); xorBitMap(17)(87) := previousCrc(23); xorBitMap(17)(89) := previousCrc(25); xorBitMap(17)(91) := previousCrc(27); xorBitMap(17)(94) := previousCrc(30); xorBitMap(17)(95) := previousCrc(31); 
      xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(66) := previousCrc(2); xorBitMap(18)(70) := previousCrc(6); xorBitMap(18)(71) := previousCrc(7); xorBitMap(18)(74) := previousCrc(10); xorBitMap(18)(78) := previousCrc(14); xorBitMap(18)(79) := previousCrc(15); xorBitMap(18)(83) := previousCrc(19); xorBitMap(18)(85) := previousCrc(21); xorBitMap(18)(87) := previousCrc(23); xorBitMap(18)(88) := previousCrc(24); xorBitMap(18)(90) := previousCrc(26); xorBitMap(18)(92) := previousCrc(28); xorBitMap(18)(95) := previousCrc(31); 
      xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(67) := previousCrc(3); xorBitMap(19)(71) := previousCrc(7); xorBitMap(19)(72) := previousCrc(8); xorBitMap(19)(75) := previousCrc(11); xorBitMap(19)(79) := previousCrc(15); xorBitMap(19)(80) := previousCrc(16); xorBitMap(19)(84) := previousCrc(20); xorBitMap(19)(86) := previousCrc(22); xorBitMap(19)(88) := previousCrc(24); xorBitMap(19)(89) := previousCrc(25); xorBitMap(19)(91) := previousCrc(27); xorBitMap(19)(93) := previousCrc(29); 
      xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(68) := previousCrc(4); xorBitMap(20)(72) := previousCrc(8); xorBitMap(20)(73) := previousCrc(9); xorBitMap(20)(76) := previousCrc(12); xorBitMap(20)(80) := previousCrc(16); xorBitMap(20)(81) := previousCrc(17); xorBitMap(20)(85) := previousCrc(21); xorBitMap(20)(87) := previousCrc(23); xorBitMap(20)(89) := previousCrc(25); xorBitMap(20)(90) := previousCrc(26); xorBitMap(20)(92) := previousCrc(28); xorBitMap(20)(94) := previousCrc(30); 
      xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(69) := previousCrc(5); xorBitMap(21)(73) := previousCrc(9); xorBitMap(21)(74) := previousCrc(10); xorBitMap(21)(77) := previousCrc(13); xorBitMap(21)(81) := previousCrc(17); xorBitMap(21)(82) := previousCrc(18); xorBitMap(21)(86) := previousCrc(22); xorBitMap(21)(88) := previousCrc(24); xorBitMap(21)(90) := previousCrc(26); xorBitMap(21)(91) := previousCrc(27); xorBitMap(21)(93) := previousCrc(29); xorBitMap(21)(95) := previousCrc(31); 
      xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(64) := previousCrc(0); xorBitMap(22)(73) := previousCrc(9); xorBitMap(22)(75) := previousCrc(11); xorBitMap(22)(76) := previousCrc(12); xorBitMap(22)(78) := previousCrc(14); xorBitMap(22)(80) := previousCrc(16); xorBitMap(22)(82) := previousCrc(18); xorBitMap(22)(83) := previousCrc(19); xorBitMap(22)(87) := previousCrc(23); xorBitMap(22)(88) := previousCrc(24); xorBitMap(22)(90) := previousCrc(26); xorBitMap(22)(91) := previousCrc(27); xorBitMap(22)(93) := previousCrc(29); xorBitMap(22)(95) := previousCrc(31); 
      xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(64) := previousCrc(0); xorBitMap(23)(65) := previousCrc(1); xorBitMap(23)(70) := previousCrc(6); xorBitMap(23)(73) := previousCrc(9); xorBitMap(23)(77) := previousCrc(13); xorBitMap(23)(79) := previousCrc(15); xorBitMap(23)(80) := previousCrc(16); xorBitMap(23)(81) := previousCrc(17); xorBitMap(23)(83) := previousCrc(19); xorBitMap(23)(84) := previousCrc(20); xorBitMap(23)(90) := previousCrc(26); xorBitMap(23)(91) := previousCrc(27); xorBitMap(23)(93) := previousCrc(29); xorBitMap(23)(95) := previousCrc(31); 
      xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(65) := previousCrc(1); xorBitMap(24)(66) := previousCrc(2); xorBitMap(24)(71) := previousCrc(7); xorBitMap(24)(74) := previousCrc(10); xorBitMap(24)(78) := previousCrc(14); xorBitMap(24)(80) := previousCrc(16); xorBitMap(24)(81) := previousCrc(17); xorBitMap(24)(82) := previousCrc(18); xorBitMap(24)(84) := previousCrc(20); xorBitMap(24)(85) := previousCrc(21); xorBitMap(24)(91) := previousCrc(27); xorBitMap(24)(92) := previousCrc(28); xorBitMap(24)(94) := previousCrc(30); 
      xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(66) := previousCrc(2); xorBitMap(25)(67) := previousCrc(3); xorBitMap(25)(72) := previousCrc(8); xorBitMap(25)(75) := previousCrc(11); xorBitMap(25)(79) := previousCrc(15); xorBitMap(25)(81) := previousCrc(17); xorBitMap(25)(82) := previousCrc(18); xorBitMap(25)(83) := previousCrc(19); xorBitMap(25)(85) := previousCrc(21); xorBitMap(25)(86) := previousCrc(22); xorBitMap(25)(92) := previousCrc(28); xorBitMap(25)(93) := previousCrc(29); xorBitMap(25)(95) := previousCrc(31); 
      xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(64) := previousCrc(0); xorBitMap(26)(67) := previousCrc(3); xorBitMap(26)(68) := previousCrc(4); xorBitMap(26)(70) := previousCrc(6); xorBitMap(26)(74) := previousCrc(10); xorBitMap(26)(82) := previousCrc(18); xorBitMap(26)(83) := previousCrc(19); xorBitMap(26)(84) := previousCrc(20); xorBitMap(26)(86) := previousCrc(22); xorBitMap(26)(87) := previousCrc(23); xorBitMap(26)(88) := previousCrc(24); xorBitMap(26)(89) := previousCrc(25); xorBitMap(26)(90) := previousCrc(26); xorBitMap(26)(92) := previousCrc(28); xorBitMap(26)(95) := previousCrc(31); 
      xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(65) := previousCrc(1); xorBitMap(27)(68) := previousCrc(4); xorBitMap(27)(69) := previousCrc(5); xorBitMap(27)(71) := previousCrc(7); xorBitMap(27)(75) := previousCrc(11); xorBitMap(27)(83) := previousCrc(19); xorBitMap(27)(84) := previousCrc(20); xorBitMap(27)(85) := previousCrc(21); xorBitMap(27)(87) := previousCrc(23); xorBitMap(27)(88) := previousCrc(24); xorBitMap(27)(89) := previousCrc(25); xorBitMap(27)(90) := previousCrc(26); xorBitMap(27)(91) := previousCrc(27); xorBitMap(27)(93) := previousCrc(29); 
      xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(66) := previousCrc(2); xorBitMap(28)(69) := previousCrc(5); xorBitMap(28)(70) := previousCrc(6); xorBitMap(28)(72) := previousCrc(8); xorBitMap(28)(76) := previousCrc(12); xorBitMap(28)(84) := previousCrc(20); xorBitMap(28)(85) := previousCrc(21); xorBitMap(28)(86) := previousCrc(22); xorBitMap(28)(88) := previousCrc(24); xorBitMap(28)(89) := previousCrc(25); xorBitMap(28)(90) := previousCrc(26); xorBitMap(28)(91) := previousCrc(27); xorBitMap(28)(92) := previousCrc(28); xorBitMap(28)(94) := previousCrc(30); 
      xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(67) := previousCrc(3); xorBitMap(29)(70) := previousCrc(6); xorBitMap(29)(71) := previousCrc(7); xorBitMap(29)(73) := previousCrc(9); xorBitMap(29)(77) := previousCrc(13); xorBitMap(29)(85) := previousCrc(21); xorBitMap(29)(86) := previousCrc(22); xorBitMap(29)(87) := previousCrc(23); xorBitMap(29)(89) := previousCrc(25); xorBitMap(29)(90) := previousCrc(26); xorBitMap(29)(91) := previousCrc(27); xorBitMap(29)(92) := previousCrc(28); xorBitMap(29)(93) := previousCrc(29); xorBitMap(29)(95) := previousCrc(31); 
      xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(68) := previousCrc(4); xorBitMap(30)(71) := previousCrc(7); xorBitMap(30)(72) := previousCrc(8); xorBitMap(30)(74) := previousCrc(10); xorBitMap(30)(78) := previousCrc(14); xorBitMap(30)(86) := previousCrc(22); xorBitMap(30)(87) := previousCrc(23); xorBitMap(30)(88) := previousCrc(24); xorBitMap(30)(90) := previousCrc(26); xorBitMap(30)(91) := previousCrc(27); xorBitMap(30)(92) := previousCrc(28); xorBitMap(30)(93) := previousCrc(29); xorBitMap(30)(94) := previousCrc(30); 
      xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(69) := previousCrc(5); xorBitMap(31)(72) := previousCrc(8); xorBitMap(31)(73) := previousCrc(9); xorBitMap(31)(75) := previousCrc(11); xorBitMap(31)(79) := previousCrc(15); xorBitMap(31)(87) := previousCrc(23); xorBitMap(31)(88) := previousCrc(24); xorBitMap(31)(89) := previousCrc(25); xorBitMap(31)(91) := previousCrc(27); xorBitMap(31)(92) := previousCrc(28); xorBitMap(31)(93) := previousCrc(29); xorBitMap(31)(94) := previousCrc(30); xorBitMap(31)(95) := previousCrc(31); 
   end procedure;

   procedure xorBitMap5Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(39 downto 0)) is 
   begin
      xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(65) := previousCrc(1); xorBitMap(0)(66) := previousCrc(2); xorBitMap(0)(68) := previousCrc(4); xorBitMap(0)(72) := previousCrc(8); xorBitMap(0)(80) := previousCrc(16); xorBitMap(0)(81) := previousCrc(17); xorBitMap(0)(82) := previousCrc(18); xorBitMap(0)(84) := previousCrc(20); xorBitMap(0)(85) := previousCrc(21); xorBitMap(0)(86) := previousCrc(22); xorBitMap(0)(87) := previousCrc(23); xorBitMap(0)(88) := previousCrc(24); xorBitMap(0)(90) := previousCrc(26); xorBitMap(0)(93) := previousCrc(29); 
      xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(65) := previousCrc(1); xorBitMap(1)(67) := previousCrc(3); xorBitMap(1)(68) := previousCrc(4); xorBitMap(1)(69) := previousCrc(5); xorBitMap(1)(72) := previousCrc(8); xorBitMap(1)(73) := previousCrc(9); xorBitMap(1)(80) := previousCrc(16); xorBitMap(1)(83) := previousCrc(19); xorBitMap(1)(84) := previousCrc(20); xorBitMap(1)(89) := previousCrc(25); xorBitMap(1)(90) := previousCrc(26); xorBitMap(1)(91) := previousCrc(27); xorBitMap(1)(93) := previousCrc(29); xorBitMap(1)(94) := previousCrc(30); 
      xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(64) := previousCrc(0); xorBitMap(2)(65) := previousCrc(1); xorBitMap(2)(69) := previousCrc(5); xorBitMap(2)(70) := previousCrc(6); xorBitMap(2)(72) := previousCrc(8); xorBitMap(2)(73) := previousCrc(9); xorBitMap(2)(74) := previousCrc(10); xorBitMap(2)(80) := previousCrc(16); xorBitMap(2)(82) := previousCrc(18); xorBitMap(2)(86) := previousCrc(22); xorBitMap(2)(87) := previousCrc(23); xorBitMap(2)(88) := previousCrc(24); xorBitMap(2)(91) := previousCrc(27); xorBitMap(2)(92) := previousCrc(28); xorBitMap(2)(93) := previousCrc(29); xorBitMap(2)(94) := previousCrc(30); xorBitMap(2)(95) := previousCrc(31); 
      xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(64) := previousCrc(0); xorBitMap(3)(65) := previousCrc(1); xorBitMap(3)(66) := previousCrc(2); xorBitMap(3)(70) := previousCrc(6); xorBitMap(3)(71) := previousCrc(7); xorBitMap(3)(73) := previousCrc(9); xorBitMap(3)(74) := previousCrc(10); xorBitMap(3)(75) := previousCrc(11); xorBitMap(3)(81) := previousCrc(17); xorBitMap(3)(83) := previousCrc(19); xorBitMap(3)(87) := previousCrc(23); xorBitMap(3)(88) := previousCrc(24); xorBitMap(3)(89) := previousCrc(25); xorBitMap(3)(92) := previousCrc(28); xorBitMap(3)(93) := previousCrc(29); xorBitMap(3)(94) := previousCrc(30); xorBitMap(3)(95) := previousCrc(31); 
      xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(64) := previousCrc(0); xorBitMap(4)(67) := previousCrc(3); xorBitMap(4)(68) := previousCrc(4); xorBitMap(4)(71) := previousCrc(7); xorBitMap(4)(74) := previousCrc(10); xorBitMap(4)(75) := previousCrc(11); xorBitMap(4)(76) := previousCrc(12); xorBitMap(4)(80) := previousCrc(16); xorBitMap(4)(81) := previousCrc(17); xorBitMap(4)(85) := previousCrc(21); xorBitMap(4)(86) := previousCrc(22); xorBitMap(4)(87) := previousCrc(23); xorBitMap(4)(89) := previousCrc(25); xorBitMap(4)(94) := previousCrc(30); xorBitMap(4)(95) := previousCrc(31); 
      xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(66) := previousCrc(2); xorBitMap(5)(69) := previousCrc(5); xorBitMap(5)(75) := previousCrc(11); xorBitMap(5)(76) := previousCrc(12); xorBitMap(5)(77) := previousCrc(13); xorBitMap(5)(80) := previousCrc(16); xorBitMap(5)(84) := previousCrc(20); xorBitMap(5)(85) := previousCrc(21); xorBitMap(5)(93) := previousCrc(29); xorBitMap(5)(95) := previousCrc(31); 
      xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(64) := previousCrc(0); xorBitMap(6)(67) := previousCrc(3); xorBitMap(6)(70) := previousCrc(6); xorBitMap(6)(76) := previousCrc(12); xorBitMap(6)(77) := previousCrc(13); xorBitMap(6)(78) := previousCrc(14); xorBitMap(6)(81) := previousCrc(17); xorBitMap(6)(85) := previousCrc(21); xorBitMap(6)(86) := previousCrc(22); xorBitMap(6)(94) := previousCrc(30); 
      xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(64) := previousCrc(0); xorBitMap(7)(66) := previousCrc(2); xorBitMap(7)(71) := previousCrc(7); xorBitMap(7)(72) := previousCrc(8); xorBitMap(7)(77) := previousCrc(13); xorBitMap(7)(78) := previousCrc(14); xorBitMap(7)(79) := previousCrc(15); xorBitMap(7)(80) := previousCrc(16); xorBitMap(7)(81) := previousCrc(17); xorBitMap(7)(84) := previousCrc(20); xorBitMap(7)(85) := previousCrc(21); xorBitMap(7)(88) := previousCrc(24); xorBitMap(7)(90) := previousCrc(26); xorBitMap(7)(93) := previousCrc(29); xorBitMap(7)(95) := previousCrc(31); 
      xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(64) := previousCrc(0); xorBitMap(8)(66) := previousCrc(2); xorBitMap(8)(67) := previousCrc(3); xorBitMap(8)(68) := previousCrc(4); xorBitMap(8)(73) := previousCrc(9); xorBitMap(8)(78) := previousCrc(14); xorBitMap(8)(79) := previousCrc(15); xorBitMap(8)(84) := previousCrc(20); xorBitMap(8)(87) := previousCrc(23); xorBitMap(8)(88) := previousCrc(24); xorBitMap(8)(89) := previousCrc(25); xorBitMap(8)(90) := previousCrc(26); xorBitMap(8)(91) := previousCrc(27); xorBitMap(8)(93) := previousCrc(29); xorBitMap(8)(94) := previousCrc(30); 
      xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(65) := previousCrc(1); xorBitMap(9)(67) := previousCrc(3); xorBitMap(9)(68) := previousCrc(4); xorBitMap(9)(69) := previousCrc(5); xorBitMap(9)(74) := previousCrc(10); xorBitMap(9)(79) := previousCrc(15); xorBitMap(9)(80) := previousCrc(16); xorBitMap(9)(85) := previousCrc(21); xorBitMap(9)(88) := previousCrc(24); xorBitMap(9)(89) := previousCrc(25); xorBitMap(9)(90) := previousCrc(26); xorBitMap(9)(91) := previousCrc(27); xorBitMap(9)(92) := previousCrc(28); xorBitMap(9)(94) := previousCrc(30); xorBitMap(9)(95) := previousCrc(31); 
      xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(65) := previousCrc(1); xorBitMap(10)(69) := previousCrc(5); xorBitMap(10)(70) := previousCrc(6); xorBitMap(10)(72) := previousCrc(8); xorBitMap(10)(75) := previousCrc(11); xorBitMap(10)(82) := previousCrc(18); xorBitMap(10)(84) := previousCrc(20); xorBitMap(10)(85) := previousCrc(21); xorBitMap(10)(87) := previousCrc(23); xorBitMap(10)(88) := previousCrc(24); xorBitMap(10)(89) := previousCrc(25); xorBitMap(10)(91) := previousCrc(27); xorBitMap(10)(92) := previousCrc(28); xorBitMap(10)(95) := previousCrc(31); 
      xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(65) := previousCrc(1); xorBitMap(11)(68) := previousCrc(4); xorBitMap(11)(70) := previousCrc(6); xorBitMap(11)(71) := previousCrc(7); xorBitMap(11)(72) := previousCrc(8); xorBitMap(11)(73) := previousCrc(9); xorBitMap(11)(76) := previousCrc(12); xorBitMap(11)(80) := previousCrc(16); xorBitMap(11)(81) := previousCrc(17); xorBitMap(11)(82) := previousCrc(18); xorBitMap(11)(83) := previousCrc(19); xorBitMap(11)(84) := previousCrc(20); xorBitMap(11)(87) := previousCrc(23); xorBitMap(11)(89) := previousCrc(25); xorBitMap(11)(92) := previousCrc(28); 
      xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(65) := previousCrc(1); xorBitMap(12)(68) := previousCrc(4); xorBitMap(12)(69) := previousCrc(5); xorBitMap(12)(71) := previousCrc(7); xorBitMap(12)(73) := previousCrc(9); xorBitMap(12)(74) := previousCrc(10); xorBitMap(12)(77) := previousCrc(13); xorBitMap(12)(80) := previousCrc(16); xorBitMap(12)(83) := previousCrc(19); xorBitMap(12)(86) := previousCrc(22); xorBitMap(12)(87) := previousCrc(23); 
      xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(66) := previousCrc(2); xorBitMap(13)(69) := previousCrc(5); xorBitMap(13)(70) := previousCrc(6); xorBitMap(13)(72) := previousCrc(8); xorBitMap(13)(74) := previousCrc(10); xorBitMap(13)(75) := previousCrc(11); xorBitMap(13)(78) := previousCrc(14); xorBitMap(13)(81) := previousCrc(17); xorBitMap(13)(84) := previousCrc(20); xorBitMap(13)(87) := previousCrc(23); xorBitMap(13)(88) := previousCrc(24); 
      xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(64) := previousCrc(0); xorBitMap(14)(67) := previousCrc(3); xorBitMap(14)(70) := previousCrc(6); xorBitMap(14)(71) := previousCrc(7); xorBitMap(14)(73) := previousCrc(9); xorBitMap(14)(75) := previousCrc(11); xorBitMap(14)(76) := previousCrc(12); xorBitMap(14)(79) := previousCrc(15); xorBitMap(14)(82) := previousCrc(18); xorBitMap(14)(85) := previousCrc(21); xorBitMap(14)(88) := previousCrc(24); xorBitMap(14)(89) := previousCrc(25); 
      xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(64) := previousCrc(0); xorBitMap(15)(65) := previousCrc(1); xorBitMap(15)(68) := previousCrc(4); xorBitMap(15)(71) := previousCrc(7); xorBitMap(15)(72) := previousCrc(8); xorBitMap(15)(74) := previousCrc(10); xorBitMap(15)(76) := previousCrc(12); xorBitMap(15)(77) := previousCrc(13); xorBitMap(15)(80) := previousCrc(16); xorBitMap(15)(83) := previousCrc(19); xorBitMap(15)(86) := previousCrc(22); xorBitMap(15)(89) := previousCrc(25); xorBitMap(15)(90) := previousCrc(26); 
      xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(64) := previousCrc(0); xorBitMap(16)(68) := previousCrc(4); xorBitMap(16)(69) := previousCrc(5); xorBitMap(16)(73) := previousCrc(9); xorBitMap(16)(75) := previousCrc(11); xorBitMap(16)(77) := previousCrc(13); xorBitMap(16)(78) := previousCrc(14); xorBitMap(16)(80) := previousCrc(16); xorBitMap(16)(82) := previousCrc(18); xorBitMap(16)(85) := previousCrc(21); xorBitMap(16)(86) := previousCrc(22); xorBitMap(16)(88) := previousCrc(24); xorBitMap(16)(91) := previousCrc(27); xorBitMap(16)(93) := previousCrc(29); 
      xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(65) := previousCrc(1); xorBitMap(17)(69) := previousCrc(5); xorBitMap(17)(70) := previousCrc(6); xorBitMap(17)(74) := previousCrc(10); xorBitMap(17)(76) := previousCrc(12); xorBitMap(17)(78) := previousCrc(14); xorBitMap(17)(79) := previousCrc(15); xorBitMap(17)(81) := previousCrc(17); xorBitMap(17)(83) := previousCrc(19); xorBitMap(17)(86) := previousCrc(22); xorBitMap(17)(87) := previousCrc(23); xorBitMap(17)(89) := previousCrc(25); xorBitMap(17)(92) := previousCrc(28); xorBitMap(17)(94) := previousCrc(30); 
      xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(66) := previousCrc(2); xorBitMap(18)(70) := previousCrc(6); xorBitMap(18)(71) := previousCrc(7); xorBitMap(18)(75) := previousCrc(11); xorBitMap(18)(77) := previousCrc(13); xorBitMap(18)(79) := previousCrc(15); xorBitMap(18)(80) := previousCrc(16); xorBitMap(18)(82) := previousCrc(18); xorBitMap(18)(84) := previousCrc(20); xorBitMap(18)(87) := previousCrc(23); xorBitMap(18)(88) := previousCrc(24); xorBitMap(18)(90) := previousCrc(26); xorBitMap(18)(93) := previousCrc(29); xorBitMap(18)(95) := previousCrc(31); 
      xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(64) := previousCrc(0); xorBitMap(19)(67) := previousCrc(3); xorBitMap(19)(71) := previousCrc(7); xorBitMap(19)(72) := previousCrc(8); xorBitMap(19)(76) := previousCrc(12); xorBitMap(19)(78) := previousCrc(14); xorBitMap(19)(80) := previousCrc(16); xorBitMap(19)(81) := previousCrc(17); xorBitMap(19)(83) := previousCrc(19); xorBitMap(19)(85) := previousCrc(21); xorBitMap(19)(88) := previousCrc(24); xorBitMap(19)(89) := previousCrc(25); xorBitMap(19)(91) := previousCrc(27); xorBitMap(19)(94) := previousCrc(30); 
      xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(64) := previousCrc(0); xorBitMap(20)(65) := previousCrc(1); xorBitMap(20)(68) := previousCrc(4); xorBitMap(20)(72) := previousCrc(8); xorBitMap(20)(73) := previousCrc(9); xorBitMap(20)(77) := previousCrc(13); xorBitMap(20)(79) := previousCrc(15); xorBitMap(20)(81) := previousCrc(17); xorBitMap(20)(82) := previousCrc(18); xorBitMap(20)(84) := previousCrc(20); xorBitMap(20)(86) := previousCrc(22); xorBitMap(20)(89) := previousCrc(25); xorBitMap(20)(90) := previousCrc(26); xorBitMap(20)(92) := previousCrc(28); xorBitMap(20)(95) := previousCrc(31); 
      xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(65) := previousCrc(1); xorBitMap(21)(66) := previousCrc(2); xorBitMap(21)(69) := previousCrc(5); xorBitMap(21)(73) := previousCrc(9); xorBitMap(21)(74) := previousCrc(10); xorBitMap(21)(78) := previousCrc(14); xorBitMap(21)(80) := previousCrc(16); xorBitMap(21)(82) := previousCrc(18); xorBitMap(21)(83) := previousCrc(19); xorBitMap(21)(85) := previousCrc(21); xorBitMap(21)(87) := previousCrc(23); xorBitMap(21)(90) := previousCrc(26); xorBitMap(21)(91) := previousCrc(27); xorBitMap(21)(93) := previousCrc(29); 
      xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(65) := previousCrc(1); xorBitMap(22)(67) := previousCrc(3); xorBitMap(22)(68) := previousCrc(4); xorBitMap(22)(70) := previousCrc(6); xorBitMap(22)(72) := previousCrc(8); xorBitMap(22)(74) := previousCrc(10); xorBitMap(22)(75) := previousCrc(11); xorBitMap(22)(79) := previousCrc(15); xorBitMap(22)(80) := previousCrc(16); xorBitMap(22)(82) := previousCrc(18); xorBitMap(22)(83) := previousCrc(19); xorBitMap(22)(85) := previousCrc(21); xorBitMap(22)(87) := previousCrc(23); xorBitMap(22)(90) := previousCrc(26); xorBitMap(22)(91) := previousCrc(27); xorBitMap(22)(92) := previousCrc(28); xorBitMap(22)(93) := previousCrc(29); xorBitMap(22)(94) := previousCrc(30); 
      xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(65) := previousCrc(1); xorBitMap(23)(69) := previousCrc(5); xorBitMap(23)(71) := previousCrc(7); xorBitMap(23)(72) := previousCrc(8); xorBitMap(23)(73) := previousCrc(9); xorBitMap(23)(75) := previousCrc(11); xorBitMap(23)(76) := previousCrc(12); xorBitMap(23)(82) := previousCrc(18); xorBitMap(23)(83) := previousCrc(19); xorBitMap(23)(85) := previousCrc(21); xorBitMap(23)(87) := previousCrc(23); xorBitMap(23)(90) := previousCrc(26); xorBitMap(23)(91) := previousCrc(27); xorBitMap(23)(92) := previousCrc(28); xorBitMap(23)(94) := previousCrc(30); xorBitMap(23)(95) := previousCrc(31); 
      xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(66) := previousCrc(2); xorBitMap(24)(70) := previousCrc(6); xorBitMap(24)(72) := previousCrc(8); xorBitMap(24)(73) := previousCrc(9); xorBitMap(24)(74) := previousCrc(10); xorBitMap(24)(76) := previousCrc(12); xorBitMap(24)(77) := previousCrc(13); xorBitMap(24)(83) := previousCrc(19); xorBitMap(24)(84) := previousCrc(20); xorBitMap(24)(86) := previousCrc(22); xorBitMap(24)(88) := previousCrc(24); xorBitMap(24)(91) := previousCrc(27); xorBitMap(24)(92) := previousCrc(28); xorBitMap(24)(93) := previousCrc(29); xorBitMap(24)(95) := previousCrc(31); 
      xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(64) := previousCrc(0); xorBitMap(25)(67) := previousCrc(3); xorBitMap(25)(71) := previousCrc(7); xorBitMap(25)(73) := previousCrc(9); xorBitMap(25)(74) := previousCrc(10); xorBitMap(25)(75) := previousCrc(11); xorBitMap(25)(77) := previousCrc(13); xorBitMap(25)(78) := previousCrc(14); xorBitMap(25)(84) := previousCrc(20); xorBitMap(25)(85) := previousCrc(21); xorBitMap(25)(87) := previousCrc(23); xorBitMap(25)(89) := previousCrc(25); xorBitMap(25)(92) := previousCrc(28); xorBitMap(25)(93) := previousCrc(29); xorBitMap(25)(94) := previousCrc(30); 
      xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(66) := previousCrc(2); xorBitMap(26)(74) := previousCrc(10); xorBitMap(26)(75) := previousCrc(11); xorBitMap(26)(76) := previousCrc(12); xorBitMap(26)(78) := previousCrc(14); xorBitMap(26)(79) := previousCrc(15); xorBitMap(26)(80) := previousCrc(16); xorBitMap(26)(81) := previousCrc(17); xorBitMap(26)(82) := previousCrc(18); xorBitMap(26)(84) := previousCrc(20); xorBitMap(26)(87) := previousCrc(23); xorBitMap(26)(94) := previousCrc(30); xorBitMap(26)(95) := previousCrc(31); 
      xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(67) := previousCrc(3); xorBitMap(27)(75) := previousCrc(11); xorBitMap(27)(76) := previousCrc(12); xorBitMap(27)(77) := previousCrc(13); xorBitMap(27)(79) := previousCrc(15); xorBitMap(27)(80) := previousCrc(16); xorBitMap(27)(81) := previousCrc(17); xorBitMap(27)(82) := previousCrc(18); xorBitMap(27)(83) := previousCrc(19); xorBitMap(27)(85) := previousCrc(21); xorBitMap(27)(88) := previousCrc(24); xorBitMap(27)(95) := previousCrc(31); 
      xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(64) := previousCrc(0); xorBitMap(28)(68) := previousCrc(4); xorBitMap(28)(76) := previousCrc(12); xorBitMap(28)(77) := previousCrc(13); xorBitMap(28)(78) := previousCrc(14); xorBitMap(28)(80) := previousCrc(16); xorBitMap(28)(81) := previousCrc(17); xorBitMap(28)(82) := previousCrc(18); xorBitMap(28)(83) := previousCrc(19); xorBitMap(28)(84) := previousCrc(20); xorBitMap(28)(86) := previousCrc(22); xorBitMap(28)(89) := previousCrc(25); 
      xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(65) := previousCrc(1); xorBitMap(29)(69) := previousCrc(5); xorBitMap(29)(77) := previousCrc(13); xorBitMap(29)(78) := previousCrc(14); xorBitMap(29)(79) := previousCrc(15); xorBitMap(29)(81) := previousCrc(17); xorBitMap(29)(82) := previousCrc(18); xorBitMap(29)(83) := previousCrc(19); xorBitMap(29)(84) := previousCrc(20); xorBitMap(29)(85) := previousCrc(21); xorBitMap(29)(87) := previousCrc(23); xorBitMap(29)(90) := previousCrc(26); 
      xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(64) := previousCrc(0); xorBitMap(30)(66) := previousCrc(2); xorBitMap(30)(70) := previousCrc(6); xorBitMap(30)(78) := previousCrc(14); xorBitMap(30)(79) := previousCrc(15); xorBitMap(30)(80) := previousCrc(16); xorBitMap(30)(82) := previousCrc(18); xorBitMap(30)(83) := previousCrc(19); xorBitMap(30)(84) := previousCrc(20); xorBitMap(30)(85) := previousCrc(21); xorBitMap(30)(86) := previousCrc(22); xorBitMap(30)(88) := previousCrc(24); xorBitMap(30)(91) := previousCrc(27); 
      xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(64) := previousCrc(0); xorBitMap(31)(65) := previousCrc(1); xorBitMap(31)(67) := previousCrc(3); xorBitMap(31)(71) := previousCrc(7); xorBitMap(31)(79) := previousCrc(15); xorBitMap(31)(80) := previousCrc(16); xorBitMap(31)(81) := previousCrc(17); xorBitMap(31)(83) := previousCrc(19); xorBitMap(31)(84) := previousCrc(20); xorBitMap(31)(85) := previousCrc(21); xorBitMap(31)(86) := previousCrc(22); xorBitMap(31)(87) := previousCrc(23); xorBitMap(31)(89) := previousCrc(25); xorBitMap(31)(92) := previousCrc(28); 
   end procedure;

   procedure xorBitMap6Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(47 downto 0)) is 
   begin
      xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(64) := previousCrc(0); xorBitMap(0)(72) := previousCrc(8); xorBitMap(0)(73) := previousCrc(9); xorBitMap(0)(74) := previousCrc(10); xorBitMap(0)(76) := previousCrc(12); xorBitMap(0)(77) := previousCrc(13); xorBitMap(0)(78) := previousCrc(14); xorBitMap(0)(79) := previousCrc(15); xorBitMap(0)(80) := previousCrc(16); xorBitMap(0)(82) := previousCrc(18); xorBitMap(0)(85) := previousCrc(21); xorBitMap(0)(92) := previousCrc(28); xorBitMap(0)(93) := previousCrc(29); xorBitMap(0)(95) := previousCrc(31); 
      xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(64) := previousCrc(0); xorBitMap(1)(65) := previousCrc(1); xorBitMap(1)(72) := previousCrc(8); xorBitMap(1)(75) := previousCrc(11); xorBitMap(1)(76) := previousCrc(12); xorBitMap(1)(81) := previousCrc(17); xorBitMap(1)(82) := previousCrc(18); xorBitMap(1)(83) := previousCrc(19); xorBitMap(1)(85) := previousCrc(21); xorBitMap(1)(86) := previousCrc(22); xorBitMap(1)(92) := previousCrc(28); xorBitMap(1)(94) := previousCrc(30); xorBitMap(1)(95) := previousCrc(31); 
      xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(64) := previousCrc(0); xorBitMap(2)(65) := previousCrc(1); xorBitMap(2)(66) := previousCrc(2); xorBitMap(2)(72) := previousCrc(8); xorBitMap(2)(74) := previousCrc(10); xorBitMap(2)(78) := previousCrc(14); xorBitMap(2)(79) := previousCrc(15); xorBitMap(2)(80) := previousCrc(16); xorBitMap(2)(83) := previousCrc(19); xorBitMap(2)(84) := previousCrc(20); xorBitMap(2)(85) := previousCrc(21); xorBitMap(2)(86) := previousCrc(22); xorBitMap(2)(87) := previousCrc(23); xorBitMap(2)(92) := previousCrc(28); 
      xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(65) := previousCrc(1); xorBitMap(3)(66) := previousCrc(2); xorBitMap(3)(67) := previousCrc(3); xorBitMap(3)(73) := previousCrc(9); xorBitMap(3)(75) := previousCrc(11); xorBitMap(3)(79) := previousCrc(15); xorBitMap(3)(80) := previousCrc(16); xorBitMap(3)(81) := previousCrc(17); xorBitMap(3)(84) := previousCrc(20); xorBitMap(3)(85) := previousCrc(21); xorBitMap(3)(86) := previousCrc(22); xorBitMap(3)(87) := previousCrc(23); xorBitMap(3)(88) := previousCrc(24); xorBitMap(3)(93) := previousCrc(29); 
      xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(66) := previousCrc(2); xorBitMap(4)(67) := previousCrc(3); xorBitMap(4)(68) := previousCrc(4); xorBitMap(4)(72) := previousCrc(8); xorBitMap(4)(73) := previousCrc(9); xorBitMap(4)(77) := previousCrc(13); xorBitMap(4)(78) := previousCrc(14); xorBitMap(4)(79) := previousCrc(15); xorBitMap(4)(81) := previousCrc(17); xorBitMap(4)(86) := previousCrc(22); xorBitMap(4)(87) := previousCrc(23); xorBitMap(4)(88) := previousCrc(24); xorBitMap(4)(89) := previousCrc(25); xorBitMap(4)(92) := previousCrc(28); xorBitMap(4)(93) := previousCrc(29); xorBitMap(4)(94) := previousCrc(30); xorBitMap(4)(95) := previousCrc(31); 
      xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(67) := previousCrc(3); xorBitMap(5)(68) := previousCrc(4); xorBitMap(5)(69) := previousCrc(5); xorBitMap(5)(72) := previousCrc(8); xorBitMap(5)(76) := previousCrc(12); xorBitMap(5)(77) := previousCrc(13); xorBitMap(5)(85) := previousCrc(21); xorBitMap(5)(87) := previousCrc(23); xorBitMap(5)(88) := previousCrc(24); xorBitMap(5)(89) := previousCrc(25); xorBitMap(5)(90) := previousCrc(26); xorBitMap(5)(92) := previousCrc(28); xorBitMap(5)(94) := previousCrc(30); 
      xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(68) := previousCrc(4); xorBitMap(6)(69) := previousCrc(5); xorBitMap(6)(70) := previousCrc(6); xorBitMap(6)(73) := previousCrc(9); xorBitMap(6)(77) := previousCrc(13); xorBitMap(6)(78) := previousCrc(14); xorBitMap(6)(86) := previousCrc(22); xorBitMap(6)(88) := previousCrc(24); xorBitMap(6)(89) := previousCrc(25); xorBitMap(6)(90) := previousCrc(26); xorBitMap(6)(91) := previousCrc(27); xorBitMap(6)(93) := previousCrc(29); xorBitMap(6)(95) := previousCrc(31); 
      xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(64) := previousCrc(0); xorBitMap(7)(69) := previousCrc(5); xorBitMap(7)(70) := previousCrc(6); xorBitMap(7)(71) := previousCrc(7); xorBitMap(7)(72) := previousCrc(8); xorBitMap(7)(73) := previousCrc(9); xorBitMap(7)(76) := previousCrc(12); xorBitMap(7)(77) := previousCrc(13); xorBitMap(7)(80) := previousCrc(16); xorBitMap(7)(82) := previousCrc(18); xorBitMap(7)(85) := previousCrc(21); xorBitMap(7)(87) := previousCrc(23); xorBitMap(7)(89) := previousCrc(25); xorBitMap(7)(90) := previousCrc(26); xorBitMap(7)(91) := previousCrc(27); xorBitMap(7)(93) := previousCrc(29); xorBitMap(7)(94) := previousCrc(30); xorBitMap(7)(95) := previousCrc(31); 
      xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(65) := previousCrc(1); xorBitMap(8)(70) := previousCrc(6); xorBitMap(8)(71) := previousCrc(7); xorBitMap(8)(76) := previousCrc(12); xorBitMap(8)(79) := previousCrc(15); xorBitMap(8)(80) := previousCrc(16); xorBitMap(8)(81) := previousCrc(17); xorBitMap(8)(82) := previousCrc(18); xorBitMap(8)(83) := previousCrc(19); xorBitMap(8)(85) := previousCrc(21); xorBitMap(8)(86) := previousCrc(22); xorBitMap(8)(88) := previousCrc(24); xorBitMap(8)(90) := previousCrc(26); xorBitMap(8)(91) := previousCrc(27); xorBitMap(8)(93) := previousCrc(29); xorBitMap(8)(94) := previousCrc(30); 
      xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(66) := previousCrc(2); xorBitMap(9)(71) := previousCrc(7); xorBitMap(9)(72) := previousCrc(8); xorBitMap(9)(77) := previousCrc(13); xorBitMap(9)(80) := previousCrc(16); xorBitMap(9)(81) := previousCrc(17); xorBitMap(9)(82) := previousCrc(18); xorBitMap(9)(83) := previousCrc(19); xorBitMap(9)(84) := previousCrc(20); xorBitMap(9)(86) := previousCrc(22); xorBitMap(9)(87) := previousCrc(23); xorBitMap(9)(89) := previousCrc(25); xorBitMap(9)(91) := previousCrc(27); xorBitMap(9)(92) := previousCrc(28); xorBitMap(9)(94) := previousCrc(30); xorBitMap(9)(95) := previousCrc(31); 
      xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(64) := previousCrc(0); xorBitMap(10)(67) := previousCrc(3); xorBitMap(10)(74) := previousCrc(10); xorBitMap(10)(76) := previousCrc(12); xorBitMap(10)(77) := previousCrc(13); xorBitMap(10)(79) := previousCrc(15); xorBitMap(10)(80) := previousCrc(16); xorBitMap(10)(81) := previousCrc(17); xorBitMap(10)(83) := previousCrc(19); xorBitMap(10)(84) := previousCrc(20); xorBitMap(10)(87) := previousCrc(23); xorBitMap(10)(88) := previousCrc(24); xorBitMap(10)(90) := previousCrc(26); 
      xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(64) := previousCrc(0); xorBitMap(11)(65) := previousCrc(1); xorBitMap(11)(68) := previousCrc(4); xorBitMap(11)(72) := previousCrc(8); xorBitMap(11)(73) := previousCrc(9); xorBitMap(11)(74) := previousCrc(10); xorBitMap(11)(75) := previousCrc(11); xorBitMap(11)(76) := previousCrc(12); xorBitMap(11)(79) := previousCrc(15); xorBitMap(11)(81) := previousCrc(17); xorBitMap(11)(84) := previousCrc(20); xorBitMap(11)(88) := previousCrc(24); xorBitMap(11)(89) := previousCrc(25); xorBitMap(11)(91) := previousCrc(27); xorBitMap(11)(92) := previousCrc(28); xorBitMap(11)(93) := previousCrc(29); xorBitMap(11)(95) := previousCrc(31); 
      xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(65) := previousCrc(1); xorBitMap(12)(66) := previousCrc(2); xorBitMap(12)(69) := previousCrc(5); xorBitMap(12)(72) := previousCrc(8); xorBitMap(12)(75) := previousCrc(11); xorBitMap(12)(78) := previousCrc(14); xorBitMap(12)(79) := previousCrc(15); xorBitMap(12)(89) := previousCrc(25); xorBitMap(12)(90) := previousCrc(26); xorBitMap(12)(94) := previousCrc(30); xorBitMap(12)(95) := previousCrc(31); 
      xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(64) := previousCrc(0); xorBitMap(13)(66) := previousCrc(2); xorBitMap(13)(67) := previousCrc(3); xorBitMap(13)(70) := previousCrc(6); xorBitMap(13)(73) := previousCrc(9); xorBitMap(13)(76) := previousCrc(12); xorBitMap(13)(79) := previousCrc(15); xorBitMap(13)(80) := previousCrc(16); xorBitMap(13)(90) := previousCrc(26); xorBitMap(13)(91) := previousCrc(27); xorBitMap(13)(95) := previousCrc(31); 
      xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(65) := previousCrc(1); xorBitMap(14)(67) := previousCrc(3); xorBitMap(14)(68) := previousCrc(4); xorBitMap(14)(71) := previousCrc(7); xorBitMap(14)(74) := previousCrc(10); xorBitMap(14)(77) := previousCrc(13); xorBitMap(14)(80) := previousCrc(16); xorBitMap(14)(81) := previousCrc(17); xorBitMap(14)(91) := previousCrc(27); xorBitMap(14)(92) := previousCrc(28); 
      xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(64) := previousCrc(0); xorBitMap(15)(66) := previousCrc(2); xorBitMap(15)(68) := previousCrc(4); xorBitMap(15)(69) := previousCrc(5); xorBitMap(15)(72) := previousCrc(8); xorBitMap(15)(75) := previousCrc(11); xorBitMap(15)(78) := previousCrc(14); xorBitMap(15)(81) := previousCrc(17); xorBitMap(15)(82) := previousCrc(18); xorBitMap(15)(92) := previousCrc(28); xorBitMap(15)(93) := previousCrc(29); 
      xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(65) := previousCrc(1); xorBitMap(16)(67) := previousCrc(3); xorBitMap(16)(69) := previousCrc(5); xorBitMap(16)(70) := previousCrc(6); xorBitMap(16)(72) := previousCrc(8); xorBitMap(16)(74) := previousCrc(10); xorBitMap(16)(77) := previousCrc(13); xorBitMap(16)(78) := previousCrc(14); xorBitMap(16)(80) := previousCrc(16); xorBitMap(16)(83) := previousCrc(19); xorBitMap(16)(85) := previousCrc(21); xorBitMap(16)(92) := previousCrc(28); xorBitMap(16)(94) := previousCrc(30); xorBitMap(16)(95) := previousCrc(31); 
      xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(66) := previousCrc(2); xorBitMap(17)(68) := previousCrc(4); xorBitMap(17)(70) := previousCrc(6); xorBitMap(17)(71) := previousCrc(7); xorBitMap(17)(73) := previousCrc(9); xorBitMap(17)(75) := previousCrc(11); xorBitMap(17)(78) := previousCrc(14); xorBitMap(17)(79) := previousCrc(15); xorBitMap(17)(81) := previousCrc(17); xorBitMap(17)(84) := previousCrc(20); xorBitMap(17)(86) := previousCrc(22); xorBitMap(17)(93) := previousCrc(29); xorBitMap(17)(95) := previousCrc(31); 
      xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(67) := previousCrc(3); xorBitMap(18)(69) := previousCrc(5); xorBitMap(18)(71) := previousCrc(7); xorBitMap(18)(72) := previousCrc(8); xorBitMap(18)(74) := previousCrc(10); xorBitMap(18)(76) := previousCrc(12); xorBitMap(18)(79) := previousCrc(15); xorBitMap(18)(80) := previousCrc(16); xorBitMap(18)(82) := previousCrc(18); xorBitMap(18)(85) := previousCrc(21); xorBitMap(18)(87) := previousCrc(23); xorBitMap(18)(94) := previousCrc(30); 
      xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(64) := previousCrc(0); xorBitMap(19)(68) := previousCrc(4); xorBitMap(19)(70) := previousCrc(6); xorBitMap(19)(72) := previousCrc(8); xorBitMap(19)(73) := previousCrc(9); xorBitMap(19)(75) := previousCrc(11); xorBitMap(19)(77) := previousCrc(13); xorBitMap(19)(80) := previousCrc(16); xorBitMap(19)(81) := previousCrc(17); xorBitMap(19)(83) := previousCrc(19); xorBitMap(19)(86) := previousCrc(22); xorBitMap(19)(88) := previousCrc(24); xorBitMap(19)(95) := previousCrc(31); 
      xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(64) := previousCrc(0); xorBitMap(20)(65) := previousCrc(1); xorBitMap(20)(69) := previousCrc(5); xorBitMap(20)(71) := previousCrc(7); xorBitMap(20)(73) := previousCrc(9); xorBitMap(20)(74) := previousCrc(10); xorBitMap(20)(76) := previousCrc(12); xorBitMap(20)(78) := previousCrc(14); xorBitMap(20)(81) := previousCrc(17); xorBitMap(20)(82) := previousCrc(18); xorBitMap(20)(84) := previousCrc(20); xorBitMap(20)(87) := previousCrc(23); xorBitMap(20)(89) := previousCrc(25); 
      xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(65) := previousCrc(1); xorBitMap(21)(66) := previousCrc(2); xorBitMap(21)(70) := previousCrc(6); xorBitMap(21)(72) := previousCrc(8); xorBitMap(21)(74) := previousCrc(10); xorBitMap(21)(75) := previousCrc(11); xorBitMap(21)(77) := previousCrc(13); xorBitMap(21)(79) := previousCrc(15); xorBitMap(21)(82) := previousCrc(18); xorBitMap(21)(83) := previousCrc(19); xorBitMap(21)(85) := previousCrc(21); xorBitMap(21)(88) := previousCrc(24); xorBitMap(21)(90) := previousCrc(26); 
      xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(64) := previousCrc(0); xorBitMap(22)(66) := previousCrc(2); xorBitMap(22)(67) := previousCrc(3); xorBitMap(22)(71) := previousCrc(7); xorBitMap(22)(72) := previousCrc(8); xorBitMap(22)(74) := previousCrc(10); xorBitMap(22)(75) := previousCrc(11); xorBitMap(22)(77) := previousCrc(13); xorBitMap(22)(79) := previousCrc(15); xorBitMap(22)(82) := previousCrc(18); xorBitMap(22)(83) := previousCrc(19); xorBitMap(22)(84) := previousCrc(20); xorBitMap(22)(85) := previousCrc(21); xorBitMap(22)(86) := previousCrc(22); xorBitMap(22)(89) := previousCrc(25); xorBitMap(22)(91) := previousCrc(27); xorBitMap(22)(92) := previousCrc(28); xorBitMap(22)(93) := previousCrc(29); xorBitMap(22)(95) := previousCrc(31); 
      xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(64) := previousCrc(0); xorBitMap(23)(65) := previousCrc(1); xorBitMap(23)(67) := previousCrc(3); xorBitMap(23)(68) := previousCrc(4); xorBitMap(23)(74) := previousCrc(10); xorBitMap(23)(75) := previousCrc(11); xorBitMap(23)(77) := previousCrc(13); xorBitMap(23)(79) := previousCrc(15); xorBitMap(23)(82) := previousCrc(18); xorBitMap(23)(83) := previousCrc(19); xorBitMap(23)(84) := previousCrc(20); xorBitMap(23)(86) := previousCrc(22); xorBitMap(23)(87) := previousCrc(23); xorBitMap(23)(90) := previousCrc(26); xorBitMap(23)(94) := previousCrc(30); xorBitMap(23)(95) := previousCrc(31); 
      xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(64) := previousCrc(0); xorBitMap(24)(65) := previousCrc(1); xorBitMap(24)(66) := previousCrc(2); xorBitMap(24)(68) := previousCrc(4); xorBitMap(24)(69) := previousCrc(5); xorBitMap(24)(75) := previousCrc(11); xorBitMap(24)(76) := previousCrc(12); xorBitMap(24)(78) := previousCrc(14); xorBitMap(24)(80) := previousCrc(16); xorBitMap(24)(83) := previousCrc(19); xorBitMap(24)(84) := previousCrc(20); xorBitMap(24)(85) := previousCrc(21); xorBitMap(24)(87) := previousCrc(23); xorBitMap(24)(88) := previousCrc(24); xorBitMap(24)(91) := previousCrc(27); xorBitMap(24)(95) := previousCrc(31); 
      xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(65) := previousCrc(1); xorBitMap(25)(66) := previousCrc(2); xorBitMap(25)(67) := previousCrc(3); xorBitMap(25)(69) := previousCrc(5); xorBitMap(25)(70) := previousCrc(6); xorBitMap(25)(76) := previousCrc(12); xorBitMap(25)(77) := previousCrc(13); xorBitMap(25)(79) := previousCrc(15); xorBitMap(25)(81) := previousCrc(17); xorBitMap(25)(84) := previousCrc(20); xorBitMap(25)(85) := previousCrc(21); xorBitMap(25)(86) := previousCrc(22); xorBitMap(25)(88) := previousCrc(24); xorBitMap(25)(89) := previousCrc(25); xorBitMap(25)(92) := previousCrc(28); 
      xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(66) := previousCrc(2); xorBitMap(26)(67) := previousCrc(3); xorBitMap(26)(68) := previousCrc(4); xorBitMap(26)(70) := previousCrc(6); xorBitMap(26)(71) := previousCrc(7); xorBitMap(26)(72) := previousCrc(8); xorBitMap(26)(73) := previousCrc(9); xorBitMap(26)(74) := previousCrc(10); xorBitMap(26)(76) := previousCrc(12); xorBitMap(26)(79) := previousCrc(15); xorBitMap(26)(86) := previousCrc(22); xorBitMap(26)(87) := previousCrc(23); xorBitMap(26)(89) := previousCrc(25); xorBitMap(26)(90) := previousCrc(26); xorBitMap(26)(92) := previousCrc(28); xorBitMap(26)(95) := previousCrc(31); 
      xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(67) := previousCrc(3); xorBitMap(27)(68) := previousCrc(4); xorBitMap(27)(69) := previousCrc(5); xorBitMap(27)(71) := previousCrc(7); xorBitMap(27)(72) := previousCrc(8); xorBitMap(27)(73) := previousCrc(9); xorBitMap(27)(74) := previousCrc(10); xorBitMap(27)(75) := previousCrc(11); xorBitMap(27)(77) := previousCrc(13); xorBitMap(27)(80) := previousCrc(16); xorBitMap(27)(87) := previousCrc(23); xorBitMap(27)(88) := previousCrc(24); xorBitMap(27)(90) := previousCrc(26); xorBitMap(27)(91) := previousCrc(27); xorBitMap(27)(93) := previousCrc(29); 
      xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(68) := previousCrc(4); xorBitMap(28)(69) := previousCrc(5); xorBitMap(28)(70) := previousCrc(6); xorBitMap(28)(72) := previousCrc(8); xorBitMap(28)(73) := previousCrc(9); xorBitMap(28)(74) := previousCrc(10); xorBitMap(28)(75) := previousCrc(11); xorBitMap(28)(76) := previousCrc(12); xorBitMap(28)(78) := previousCrc(14); xorBitMap(28)(81) := previousCrc(17); xorBitMap(28)(88) := previousCrc(24); xorBitMap(28)(89) := previousCrc(25); xorBitMap(28)(91) := previousCrc(27); xorBitMap(28)(92) := previousCrc(28); xorBitMap(28)(94) := previousCrc(30); 
      xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(69) := previousCrc(5); xorBitMap(29)(70) := previousCrc(6); xorBitMap(29)(71) := previousCrc(7); xorBitMap(29)(73) := previousCrc(9); xorBitMap(29)(74) := previousCrc(10); xorBitMap(29)(75) := previousCrc(11); xorBitMap(29)(76) := previousCrc(12); xorBitMap(29)(77) := previousCrc(13); xorBitMap(29)(79) := previousCrc(15); xorBitMap(29)(82) := previousCrc(18); xorBitMap(29)(89) := previousCrc(25); xorBitMap(29)(90) := previousCrc(26); xorBitMap(29)(92) := previousCrc(28); xorBitMap(29)(93) := previousCrc(29); xorBitMap(29)(95) := previousCrc(31); 
      xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(70) := previousCrc(6); xorBitMap(30)(71) := previousCrc(7); xorBitMap(30)(72) := previousCrc(8); xorBitMap(30)(74) := previousCrc(10); xorBitMap(30)(75) := previousCrc(11); xorBitMap(30)(76) := previousCrc(12); xorBitMap(30)(77) := previousCrc(13); xorBitMap(30)(78) := previousCrc(14); xorBitMap(30)(80) := previousCrc(16); xorBitMap(30)(83) := previousCrc(19); xorBitMap(30)(90) := previousCrc(26); xorBitMap(30)(91) := previousCrc(27); xorBitMap(30)(93) := previousCrc(29); xorBitMap(30)(94) := previousCrc(30); 
      xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(71) := previousCrc(7); xorBitMap(31)(72) := previousCrc(8); xorBitMap(31)(73) := previousCrc(9); xorBitMap(31)(75) := previousCrc(11); xorBitMap(31)(76) := previousCrc(12); xorBitMap(31)(77) := previousCrc(13); xorBitMap(31)(78) := previousCrc(14); xorBitMap(31)(79) := previousCrc(15); xorBitMap(31)(81) := previousCrc(17); xorBitMap(31)(84) := previousCrc(20); xorBitMap(31)(91) := previousCrc(27); xorBitMap(31)(92) := previousCrc(28); xorBitMap(31)(94) := previousCrc(30); xorBitMap(31)(95) := previousCrc(31); 
   end procedure;

   procedure xorBitMap7Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(55 downto 0)) is 
   begin
      xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(64) := previousCrc(0); xorBitMap(0)(65) := previousCrc(1); xorBitMap(0)(66) := previousCrc(2); xorBitMap(0)(68) := previousCrc(4); xorBitMap(0)(69) := previousCrc(5); xorBitMap(0)(70) := previousCrc(6); xorBitMap(0)(71) := previousCrc(7); xorBitMap(0)(72) := previousCrc(8); xorBitMap(0)(74) := previousCrc(10); xorBitMap(0)(77) := previousCrc(13); xorBitMap(0)(84) := previousCrc(20); xorBitMap(0)(85) := previousCrc(21); xorBitMap(0)(87) := previousCrc(23); xorBitMap(0)(88) := previousCrc(24); xorBitMap(0)(90) := previousCrc(26); xorBitMap(0)(93) := previousCrc(29); xorBitMap(0)(94) := previousCrc(30); xorBitMap(0)(95) := previousCrc(31); 
      xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(64) := previousCrc(0); xorBitMap(1)(67) := previousCrc(3); xorBitMap(1)(68) := previousCrc(4); xorBitMap(1)(73) := previousCrc(9); xorBitMap(1)(74) := previousCrc(10); xorBitMap(1)(75) := previousCrc(11); xorBitMap(1)(77) := previousCrc(13); xorBitMap(1)(78) := previousCrc(14); xorBitMap(1)(84) := previousCrc(20); xorBitMap(1)(86) := previousCrc(22); xorBitMap(1)(87) := previousCrc(23); xorBitMap(1)(89) := previousCrc(25); xorBitMap(1)(90) := previousCrc(26); xorBitMap(1)(91) := previousCrc(27); xorBitMap(1)(93) := previousCrc(29); 
      xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(64) := previousCrc(0); xorBitMap(2)(66) := previousCrc(2); xorBitMap(2)(70) := previousCrc(6); xorBitMap(2)(71) := previousCrc(7); xorBitMap(2)(72) := previousCrc(8); xorBitMap(2)(75) := previousCrc(11); xorBitMap(2)(76) := previousCrc(12); xorBitMap(2)(77) := previousCrc(13); xorBitMap(2)(78) := previousCrc(14); xorBitMap(2)(79) := previousCrc(15); xorBitMap(2)(84) := previousCrc(20); xorBitMap(2)(91) := previousCrc(27); xorBitMap(2)(92) := previousCrc(28); xorBitMap(2)(93) := previousCrc(29); xorBitMap(2)(95) := previousCrc(31); 
      xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(65) := previousCrc(1); xorBitMap(3)(67) := previousCrc(3); xorBitMap(3)(71) := previousCrc(7); xorBitMap(3)(72) := previousCrc(8); xorBitMap(3)(73) := previousCrc(9); xorBitMap(3)(76) := previousCrc(12); xorBitMap(3)(77) := previousCrc(13); xorBitMap(3)(78) := previousCrc(14); xorBitMap(3)(79) := previousCrc(15); xorBitMap(3)(80) := previousCrc(16); xorBitMap(3)(85) := previousCrc(21); xorBitMap(3)(92) := previousCrc(28); xorBitMap(3)(93) := previousCrc(29); xorBitMap(3)(94) := previousCrc(30); 
      xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(64) := previousCrc(0); xorBitMap(4)(65) := previousCrc(1); xorBitMap(4)(69) := previousCrc(5); xorBitMap(4)(70) := previousCrc(6); xorBitMap(4)(71) := previousCrc(7); xorBitMap(4)(73) := previousCrc(9); xorBitMap(4)(78) := previousCrc(14); xorBitMap(4)(79) := previousCrc(15); xorBitMap(4)(80) := previousCrc(16); xorBitMap(4)(81) := previousCrc(17); xorBitMap(4)(84) := previousCrc(20); xorBitMap(4)(85) := previousCrc(21); xorBitMap(4)(86) := previousCrc(22); xorBitMap(4)(87) := previousCrc(23); xorBitMap(4)(88) := previousCrc(24); xorBitMap(4)(90) := previousCrc(26); 
      xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(64) := previousCrc(0); xorBitMap(5)(68) := previousCrc(4); xorBitMap(5)(69) := previousCrc(5); xorBitMap(5)(77) := previousCrc(13); xorBitMap(5)(79) := previousCrc(15); xorBitMap(5)(80) := previousCrc(16); xorBitMap(5)(81) := previousCrc(17); xorBitMap(5)(82) := previousCrc(18); xorBitMap(5)(84) := previousCrc(20); xorBitMap(5)(86) := previousCrc(22); xorBitMap(5)(89) := previousCrc(25); xorBitMap(5)(90) := previousCrc(26); xorBitMap(5)(91) := previousCrc(27); xorBitMap(5)(93) := previousCrc(29); xorBitMap(5)(94) := previousCrc(30); xorBitMap(5)(95) := previousCrc(31); 
      xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(65) := previousCrc(1); xorBitMap(6)(69) := previousCrc(5); xorBitMap(6)(70) := previousCrc(6); xorBitMap(6)(78) := previousCrc(14); xorBitMap(6)(80) := previousCrc(16); xorBitMap(6)(81) := previousCrc(17); xorBitMap(6)(82) := previousCrc(18); xorBitMap(6)(83) := previousCrc(19); xorBitMap(6)(85) := previousCrc(21); xorBitMap(6)(87) := previousCrc(23); xorBitMap(6)(90) := previousCrc(26); xorBitMap(6)(91) := previousCrc(27); xorBitMap(6)(92) := previousCrc(28); xorBitMap(6)(94) := previousCrc(30); xorBitMap(6)(95) := previousCrc(31); 
      xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(64) := previousCrc(0); xorBitMap(7)(65) := previousCrc(1); xorBitMap(7)(68) := previousCrc(4); xorBitMap(7)(69) := previousCrc(5); xorBitMap(7)(72) := previousCrc(8); xorBitMap(7)(74) := previousCrc(10); xorBitMap(7)(77) := previousCrc(13); xorBitMap(7)(79) := previousCrc(15); xorBitMap(7)(81) := previousCrc(17); xorBitMap(7)(82) := previousCrc(18); xorBitMap(7)(83) := previousCrc(19); xorBitMap(7)(85) := previousCrc(21); xorBitMap(7)(86) := previousCrc(22); xorBitMap(7)(87) := previousCrc(23); xorBitMap(7)(90) := previousCrc(26); xorBitMap(7)(91) := previousCrc(27); xorBitMap(7)(92) := previousCrc(28); xorBitMap(7)(94) := previousCrc(30); 
      xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(68) := previousCrc(4); xorBitMap(8)(71) := previousCrc(7); xorBitMap(8)(72) := previousCrc(8); xorBitMap(8)(73) := previousCrc(9); xorBitMap(8)(74) := previousCrc(10); xorBitMap(8)(75) := previousCrc(11); xorBitMap(8)(77) := previousCrc(13); xorBitMap(8)(78) := previousCrc(14); xorBitMap(8)(80) := previousCrc(16); xorBitMap(8)(82) := previousCrc(18); xorBitMap(8)(83) := previousCrc(19); xorBitMap(8)(85) := previousCrc(21); xorBitMap(8)(86) := previousCrc(22); xorBitMap(8)(90) := previousCrc(26); xorBitMap(8)(91) := previousCrc(27); xorBitMap(8)(92) := previousCrc(28); xorBitMap(8)(94) := previousCrc(30); 
      xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(64) := previousCrc(0); xorBitMap(9)(69) := previousCrc(5); xorBitMap(9)(72) := previousCrc(8); xorBitMap(9)(73) := previousCrc(9); xorBitMap(9)(74) := previousCrc(10); xorBitMap(9)(75) := previousCrc(11); xorBitMap(9)(76) := previousCrc(12); xorBitMap(9)(78) := previousCrc(14); xorBitMap(9)(79) := previousCrc(15); xorBitMap(9)(81) := previousCrc(17); xorBitMap(9)(83) := previousCrc(19); xorBitMap(9)(84) := previousCrc(20); xorBitMap(9)(86) := previousCrc(22); xorBitMap(9)(87) := previousCrc(23); xorBitMap(9)(91) := previousCrc(27); xorBitMap(9)(92) := previousCrc(28); xorBitMap(9)(93) := previousCrc(29); xorBitMap(9)(95) := previousCrc(31); 
      xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(66) := previousCrc(2); xorBitMap(10)(68) := previousCrc(4); xorBitMap(10)(69) := previousCrc(5); xorBitMap(10)(71) := previousCrc(7); xorBitMap(10)(72) := previousCrc(8); xorBitMap(10)(73) := previousCrc(9); xorBitMap(10)(75) := previousCrc(11); xorBitMap(10)(76) := previousCrc(12); xorBitMap(10)(79) := previousCrc(15); xorBitMap(10)(80) := previousCrc(16); xorBitMap(10)(82) := previousCrc(18); xorBitMap(10)(90) := previousCrc(26); xorBitMap(10)(92) := previousCrc(28); xorBitMap(10)(95) := previousCrc(31); 
      xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(64) := previousCrc(0); xorBitMap(11)(65) := previousCrc(1); xorBitMap(11)(66) := previousCrc(2); xorBitMap(11)(67) := previousCrc(3); xorBitMap(11)(68) := previousCrc(4); xorBitMap(11)(71) := previousCrc(7); xorBitMap(11)(73) := previousCrc(9); xorBitMap(11)(76) := previousCrc(12); xorBitMap(11)(80) := previousCrc(16); xorBitMap(11)(81) := previousCrc(17); xorBitMap(11)(83) := previousCrc(19); xorBitMap(11)(84) := previousCrc(20); xorBitMap(11)(85) := previousCrc(21); xorBitMap(11)(87) := previousCrc(23); xorBitMap(11)(88) := previousCrc(24); xorBitMap(11)(90) := previousCrc(26); xorBitMap(11)(91) := previousCrc(27); xorBitMap(11)(94) := previousCrc(30); xorBitMap(11)(95) := previousCrc(31); 
      xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(64) := previousCrc(0); xorBitMap(12)(67) := previousCrc(3); xorBitMap(12)(70) := previousCrc(6); xorBitMap(12)(71) := previousCrc(7); xorBitMap(12)(81) := previousCrc(17); xorBitMap(12)(82) := previousCrc(18); xorBitMap(12)(86) := previousCrc(22); xorBitMap(12)(87) := previousCrc(23); xorBitMap(12)(89) := previousCrc(25); xorBitMap(12)(90) := previousCrc(26); xorBitMap(12)(91) := previousCrc(27); xorBitMap(12)(92) := previousCrc(28); xorBitMap(12)(93) := previousCrc(29); xorBitMap(12)(94) := previousCrc(30); 
      xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(65) := previousCrc(1); xorBitMap(13)(68) := previousCrc(4); xorBitMap(13)(71) := previousCrc(7); xorBitMap(13)(72) := previousCrc(8); xorBitMap(13)(82) := previousCrc(18); xorBitMap(13)(83) := previousCrc(19); xorBitMap(13)(87) := previousCrc(23); xorBitMap(13)(88) := previousCrc(24); xorBitMap(13)(90) := previousCrc(26); xorBitMap(13)(91) := previousCrc(27); xorBitMap(13)(92) := previousCrc(28); xorBitMap(13)(93) := previousCrc(29); xorBitMap(13)(94) := previousCrc(30); xorBitMap(13)(95) := previousCrc(31); 
      xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(66) := previousCrc(2); xorBitMap(14)(69) := previousCrc(5); xorBitMap(14)(72) := previousCrc(8); xorBitMap(14)(73) := previousCrc(9); xorBitMap(14)(83) := previousCrc(19); xorBitMap(14)(84) := previousCrc(20); xorBitMap(14)(88) := previousCrc(24); xorBitMap(14)(89) := previousCrc(25); xorBitMap(14)(91) := previousCrc(27); xorBitMap(14)(92) := previousCrc(28); xorBitMap(14)(93) := previousCrc(29); xorBitMap(14)(94) := previousCrc(30); xorBitMap(14)(95) := previousCrc(31); 
      xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(64) := previousCrc(0); xorBitMap(15)(67) := previousCrc(3); xorBitMap(15)(70) := previousCrc(6); xorBitMap(15)(73) := previousCrc(9); xorBitMap(15)(74) := previousCrc(10); xorBitMap(15)(84) := previousCrc(20); xorBitMap(15)(85) := previousCrc(21); xorBitMap(15)(89) := previousCrc(25); xorBitMap(15)(90) := previousCrc(26); xorBitMap(15)(92) := previousCrc(28); xorBitMap(15)(93) := previousCrc(29); xorBitMap(15)(94) := previousCrc(30); xorBitMap(15)(95) := previousCrc(31); 
      xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(64) := previousCrc(0); xorBitMap(16)(66) := previousCrc(2); xorBitMap(16)(69) := previousCrc(5); xorBitMap(16)(70) := previousCrc(6); xorBitMap(16)(72) := previousCrc(8); xorBitMap(16)(75) := previousCrc(11); xorBitMap(16)(77) := previousCrc(13); xorBitMap(16)(84) := previousCrc(20); xorBitMap(16)(86) := previousCrc(22); xorBitMap(16)(87) := previousCrc(23); xorBitMap(16)(88) := previousCrc(24); xorBitMap(16)(91) := previousCrc(27); 
      xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(65) := previousCrc(1); xorBitMap(17)(67) := previousCrc(3); xorBitMap(17)(70) := previousCrc(6); xorBitMap(17)(71) := previousCrc(7); xorBitMap(17)(73) := previousCrc(9); xorBitMap(17)(76) := previousCrc(12); xorBitMap(17)(78) := previousCrc(14); xorBitMap(17)(85) := previousCrc(21); xorBitMap(17)(87) := previousCrc(23); xorBitMap(17)(88) := previousCrc(24); xorBitMap(17)(89) := previousCrc(25); xorBitMap(17)(92) := previousCrc(28); 
      xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(64) := previousCrc(0); xorBitMap(18)(66) := previousCrc(2); xorBitMap(18)(68) := previousCrc(4); xorBitMap(18)(71) := previousCrc(7); xorBitMap(18)(72) := previousCrc(8); xorBitMap(18)(74) := previousCrc(10); xorBitMap(18)(77) := previousCrc(13); xorBitMap(18)(79) := previousCrc(15); xorBitMap(18)(86) := previousCrc(22); xorBitMap(18)(88) := previousCrc(24); xorBitMap(18)(89) := previousCrc(25); xorBitMap(18)(90) := previousCrc(26); xorBitMap(18)(93) := previousCrc(29); 
      xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(64) := previousCrc(0); xorBitMap(19)(65) := previousCrc(1); xorBitMap(19)(67) := previousCrc(3); xorBitMap(19)(69) := previousCrc(5); xorBitMap(19)(72) := previousCrc(8); xorBitMap(19)(73) := previousCrc(9); xorBitMap(19)(75) := previousCrc(11); xorBitMap(19)(78) := previousCrc(14); xorBitMap(19)(80) := previousCrc(16); xorBitMap(19)(87) := previousCrc(23); xorBitMap(19)(89) := previousCrc(25); xorBitMap(19)(90) := previousCrc(26); xorBitMap(19)(91) := previousCrc(27); xorBitMap(19)(94) := previousCrc(30); 
      xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(65) := previousCrc(1); xorBitMap(20)(66) := previousCrc(2); xorBitMap(20)(68) := previousCrc(4); xorBitMap(20)(70) := previousCrc(6); xorBitMap(20)(73) := previousCrc(9); xorBitMap(20)(74) := previousCrc(10); xorBitMap(20)(76) := previousCrc(12); xorBitMap(20)(79) := previousCrc(15); xorBitMap(20)(81) := previousCrc(17); xorBitMap(20)(88) := previousCrc(24); xorBitMap(20)(90) := previousCrc(26); xorBitMap(20)(91) := previousCrc(27); xorBitMap(20)(92) := previousCrc(28); xorBitMap(20)(95) := previousCrc(31); 
      xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(64) := previousCrc(0); xorBitMap(21)(66) := previousCrc(2); xorBitMap(21)(67) := previousCrc(3); xorBitMap(21)(69) := previousCrc(5); xorBitMap(21)(71) := previousCrc(7); xorBitMap(21)(74) := previousCrc(10); xorBitMap(21)(75) := previousCrc(11); xorBitMap(21)(77) := previousCrc(13); xorBitMap(21)(80) := previousCrc(16); xorBitMap(21)(82) := previousCrc(18); xorBitMap(21)(89) := previousCrc(25); xorBitMap(21)(91) := previousCrc(27); xorBitMap(21)(92) := previousCrc(28); xorBitMap(21)(93) := previousCrc(29); 
      xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(64) := previousCrc(0); xorBitMap(22)(66) := previousCrc(2); xorBitMap(22)(67) := previousCrc(3); xorBitMap(22)(69) := previousCrc(5); xorBitMap(22)(71) := previousCrc(7); xorBitMap(22)(74) := previousCrc(10); xorBitMap(22)(75) := previousCrc(11); xorBitMap(22)(76) := previousCrc(12); xorBitMap(22)(77) := previousCrc(13); xorBitMap(22)(78) := previousCrc(14); xorBitMap(22)(81) := previousCrc(17); xorBitMap(22)(83) := previousCrc(19); xorBitMap(22)(84) := previousCrc(20); xorBitMap(22)(85) := previousCrc(21); xorBitMap(22)(87) := previousCrc(23); xorBitMap(22)(88) := previousCrc(24); xorBitMap(22)(92) := previousCrc(28); xorBitMap(22)(95) := previousCrc(31); 
      xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(66) := previousCrc(2); xorBitMap(23)(67) := previousCrc(3); xorBitMap(23)(69) := previousCrc(5); xorBitMap(23)(71) := previousCrc(7); xorBitMap(23)(74) := previousCrc(10); xorBitMap(23)(75) := previousCrc(11); xorBitMap(23)(76) := previousCrc(12); xorBitMap(23)(78) := previousCrc(14); xorBitMap(23)(79) := previousCrc(15); xorBitMap(23)(82) := previousCrc(18); xorBitMap(23)(86) := previousCrc(22); xorBitMap(23)(87) := previousCrc(23); xorBitMap(23)(89) := previousCrc(25); xorBitMap(23)(90) := previousCrc(26); xorBitMap(23)(94) := previousCrc(30); xorBitMap(23)(95) := previousCrc(31); 
      xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(67) := previousCrc(3); xorBitMap(24)(68) := previousCrc(4); xorBitMap(24)(70) := previousCrc(6); xorBitMap(24)(72) := previousCrc(8); xorBitMap(24)(75) := previousCrc(11); xorBitMap(24)(76) := previousCrc(12); xorBitMap(24)(77) := previousCrc(13); xorBitMap(24)(79) := previousCrc(15); xorBitMap(24)(80) := previousCrc(16); xorBitMap(24)(83) := previousCrc(19); xorBitMap(24)(87) := previousCrc(23); xorBitMap(24)(88) := previousCrc(24); xorBitMap(24)(90) := previousCrc(26); xorBitMap(24)(91) := previousCrc(27); xorBitMap(24)(95) := previousCrc(31); 
      xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(68) := previousCrc(4); xorBitMap(25)(69) := previousCrc(5); xorBitMap(25)(71) := previousCrc(7); xorBitMap(25)(73) := previousCrc(9); xorBitMap(25)(76) := previousCrc(12); xorBitMap(25)(77) := previousCrc(13); xorBitMap(25)(78) := previousCrc(14); xorBitMap(25)(80) := previousCrc(16); xorBitMap(25)(81) := previousCrc(17); xorBitMap(25)(84) := previousCrc(20); xorBitMap(25)(88) := previousCrc(24); xorBitMap(25)(89) := previousCrc(25); xorBitMap(25)(91) := previousCrc(27); xorBitMap(25)(92) := previousCrc(28); 
      xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(64) := previousCrc(0); xorBitMap(26)(65) := previousCrc(1); xorBitMap(26)(66) := previousCrc(2); xorBitMap(26)(68) := previousCrc(4); xorBitMap(26)(71) := previousCrc(7); xorBitMap(26)(78) := previousCrc(14); xorBitMap(26)(79) := previousCrc(15); xorBitMap(26)(81) := previousCrc(17); xorBitMap(26)(82) := previousCrc(18); xorBitMap(26)(84) := previousCrc(20); xorBitMap(26)(87) := previousCrc(23); xorBitMap(26)(88) := previousCrc(24); xorBitMap(26)(89) := previousCrc(25); xorBitMap(26)(92) := previousCrc(28); xorBitMap(26)(94) := previousCrc(30); xorBitMap(26)(95) := previousCrc(31); 
      xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(64) := previousCrc(0); xorBitMap(27)(65) := previousCrc(1); xorBitMap(27)(66) := previousCrc(2); xorBitMap(27)(67) := previousCrc(3); xorBitMap(27)(69) := previousCrc(5); xorBitMap(27)(72) := previousCrc(8); xorBitMap(27)(79) := previousCrc(15); xorBitMap(27)(80) := previousCrc(16); xorBitMap(27)(82) := previousCrc(18); xorBitMap(27)(83) := previousCrc(19); xorBitMap(27)(85) := previousCrc(21); xorBitMap(27)(88) := previousCrc(24); xorBitMap(27)(89) := previousCrc(25); xorBitMap(27)(90) := previousCrc(26); xorBitMap(27)(93) := previousCrc(29); xorBitMap(27)(95) := previousCrc(31); 
      xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(64) := previousCrc(0); xorBitMap(28)(65) := previousCrc(1); xorBitMap(28)(66) := previousCrc(2); xorBitMap(28)(67) := previousCrc(3); xorBitMap(28)(68) := previousCrc(4); xorBitMap(28)(70) := previousCrc(6); xorBitMap(28)(73) := previousCrc(9); xorBitMap(28)(80) := previousCrc(16); xorBitMap(28)(81) := previousCrc(17); xorBitMap(28)(83) := previousCrc(19); xorBitMap(28)(84) := previousCrc(20); xorBitMap(28)(86) := previousCrc(22); xorBitMap(28)(89) := previousCrc(25); xorBitMap(28)(90) := previousCrc(26); xorBitMap(28)(91) := previousCrc(27); xorBitMap(28)(94) := previousCrc(30); 
      xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(65) := previousCrc(1); xorBitMap(29)(66) := previousCrc(2); xorBitMap(29)(67) := previousCrc(3); xorBitMap(29)(68) := previousCrc(4); xorBitMap(29)(69) := previousCrc(5); xorBitMap(29)(71) := previousCrc(7); xorBitMap(29)(74) := previousCrc(10); xorBitMap(29)(81) := previousCrc(17); xorBitMap(29)(82) := previousCrc(18); xorBitMap(29)(84) := previousCrc(20); xorBitMap(29)(85) := previousCrc(21); xorBitMap(29)(87) := previousCrc(23); xorBitMap(29)(90) := previousCrc(26); xorBitMap(29)(91) := previousCrc(27); xorBitMap(29)(92) := previousCrc(28); xorBitMap(29)(95) := previousCrc(31); 
      xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(64) := previousCrc(0); xorBitMap(30)(66) := previousCrc(2); xorBitMap(30)(67) := previousCrc(3); xorBitMap(30)(68) := previousCrc(4); xorBitMap(30)(69) := previousCrc(5); xorBitMap(30)(70) := previousCrc(6); xorBitMap(30)(72) := previousCrc(8); xorBitMap(30)(75) := previousCrc(11); xorBitMap(30)(82) := previousCrc(18); xorBitMap(30)(83) := previousCrc(19); xorBitMap(30)(85) := previousCrc(21); xorBitMap(30)(86) := previousCrc(22); xorBitMap(30)(88) := previousCrc(24); xorBitMap(30)(91) := previousCrc(27); xorBitMap(30)(92) := previousCrc(28); xorBitMap(30)(93) := previousCrc(29); 
      xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(64) := previousCrc(0); xorBitMap(31)(65) := previousCrc(1); xorBitMap(31)(67) := previousCrc(3); xorBitMap(31)(68) := previousCrc(4); xorBitMap(31)(69) := previousCrc(5); xorBitMap(31)(70) := previousCrc(6); xorBitMap(31)(71) := previousCrc(7); xorBitMap(31)(73) := previousCrc(9); xorBitMap(31)(76) := previousCrc(12); xorBitMap(31)(83) := previousCrc(19); xorBitMap(31)(84) := previousCrc(20); xorBitMap(31)(86) := previousCrc(22); xorBitMap(31)(87) := previousCrc(23); xorBitMap(31)(89) := previousCrc(25); xorBitMap(31)(92) := previousCrc(28); xorBitMap(31)(93) := previousCrc(29); xorBitMap(31)(94) := previousCrc(30); 
   end procedure;

   procedure xorBitMap8Byte (
      xorBitMap   : inout Slv96Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(63 downto 0)) is 
   begin
      xorBitMap(0)(63) := currentData(63); xorBitMap(0)(61) := currentData(61); xorBitMap(0)(60) := currentData(60); xorBitMap(0)(58) := currentData(58); xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(64) := previousCrc(0); xorBitMap(0)(66) := previousCrc(2); xorBitMap(0)(69) := previousCrc(5); xorBitMap(0)(76) := previousCrc(12); xorBitMap(0)(77) := previousCrc(13); xorBitMap(0)(79) := previousCrc(15); xorBitMap(0)(80) := previousCrc(16); xorBitMap(0)(82) := previousCrc(18); xorBitMap(0)(85) := previousCrc(21); xorBitMap(0)(86) := previousCrc(22); xorBitMap(0)(87) := previousCrc(23); xorBitMap(0)(90) := previousCrc(26); xorBitMap(0)(92) := previousCrc(28); xorBitMap(0)(93) := previousCrc(29); xorBitMap(0)(95) := previousCrc(31); 
      xorBitMap(1)(63) := currentData(63); xorBitMap(1)(62) := currentData(62); xorBitMap(1)(60) := currentData(60); xorBitMap(1)(59) := currentData(59); xorBitMap(1)(58) := currentData(58); xorBitMap(1)(56) := currentData(56); xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(65) := previousCrc(1); xorBitMap(1)(66) := previousCrc(2); xorBitMap(1)(67) := previousCrc(3); xorBitMap(1)(69) := previousCrc(5); xorBitMap(1)(70) := previousCrc(6); xorBitMap(1)(76) := previousCrc(12); xorBitMap(1)(78) := previousCrc(14); xorBitMap(1)(79) := previousCrc(15); xorBitMap(1)(81) := previousCrc(17); xorBitMap(1)(82) := previousCrc(18); xorBitMap(1)(83) := previousCrc(19); xorBitMap(1)(85) := previousCrc(21); xorBitMap(1)(88) := previousCrc(24); xorBitMap(1)(90) := previousCrc(26); xorBitMap(1)(91) := previousCrc(27); xorBitMap(1)(92) := previousCrc(28); xorBitMap(1)(94) := previousCrc(30); xorBitMap(1)(95) := previousCrc(31); 
      xorBitMap(2)(59) := currentData(59); xorBitMap(2)(58) := currentData(58); xorBitMap(2)(57) := currentData(57); xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(64) := previousCrc(0); xorBitMap(2)(67) := previousCrc(3); xorBitMap(2)(68) := previousCrc(4); xorBitMap(2)(69) := previousCrc(5); xorBitMap(2)(70) := previousCrc(6); xorBitMap(2)(71) := previousCrc(7); xorBitMap(2)(76) := previousCrc(12); xorBitMap(2)(83) := previousCrc(19); xorBitMap(2)(84) := previousCrc(20); xorBitMap(2)(85) := previousCrc(21); xorBitMap(2)(87) := previousCrc(23); xorBitMap(2)(89) := previousCrc(25); xorBitMap(2)(90) := previousCrc(26); xorBitMap(2)(91) := previousCrc(27); 
      xorBitMap(3)(60) := currentData(60); xorBitMap(3)(59) := currentData(59); xorBitMap(3)(58) := currentData(58); xorBitMap(3)(56) := currentData(56); xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(64) := previousCrc(0); xorBitMap(3)(65) := previousCrc(1); xorBitMap(3)(68) := previousCrc(4); xorBitMap(3)(69) := previousCrc(5); xorBitMap(3)(70) := previousCrc(6); xorBitMap(3)(71) := previousCrc(7); xorBitMap(3)(72) := previousCrc(8); xorBitMap(3)(77) := previousCrc(13); xorBitMap(3)(84) := previousCrc(20); xorBitMap(3)(85) := previousCrc(21); xorBitMap(3)(86) := previousCrc(22); xorBitMap(3)(88) := previousCrc(24); xorBitMap(3)(90) := previousCrc(26); xorBitMap(3)(91) := previousCrc(27); xorBitMap(3)(92) := previousCrc(28); 
      xorBitMap(4)(63) := currentData(63); xorBitMap(4)(59) := currentData(59); xorBitMap(4)(58) := currentData(58); xorBitMap(4)(57) := currentData(57); xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(65) := previousCrc(1); xorBitMap(4)(70) := previousCrc(6); xorBitMap(4)(71) := previousCrc(7); xorBitMap(4)(72) := previousCrc(8); xorBitMap(4)(73) := previousCrc(9); xorBitMap(4)(76) := previousCrc(12); xorBitMap(4)(77) := previousCrc(13); xorBitMap(4)(78) := previousCrc(14); xorBitMap(4)(79) := previousCrc(15); xorBitMap(4)(80) := previousCrc(16); xorBitMap(4)(82) := previousCrc(18); xorBitMap(4)(89) := previousCrc(25); xorBitMap(4)(90) := previousCrc(26); xorBitMap(4)(91) := previousCrc(27); xorBitMap(4)(95) := previousCrc(31); 
      xorBitMap(5)(63) := currentData(63); xorBitMap(5)(61) := currentData(61); xorBitMap(5)(59) := currentData(59); xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(69) := previousCrc(5); xorBitMap(5)(71) := previousCrc(7); xorBitMap(5)(72) := previousCrc(8); xorBitMap(5)(73) := previousCrc(9); xorBitMap(5)(74) := previousCrc(10); xorBitMap(5)(76) := previousCrc(12); xorBitMap(5)(78) := previousCrc(14); xorBitMap(5)(81) := previousCrc(17); xorBitMap(5)(82) := previousCrc(18); xorBitMap(5)(83) := previousCrc(19); xorBitMap(5)(85) := previousCrc(21); xorBitMap(5)(86) := previousCrc(22); xorBitMap(5)(87) := previousCrc(23); xorBitMap(5)(91) := previousCrc(27); xorBitMap(5)(93) := previousCrc(29); xorBitMap(5)(95) := previousCrc(31); 
      xorBitMap(6)(62) := currentData(62); xorBitMap(6)(60) := currentData(60); xorBitMap(6)(56) := currentData(56); xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(70) := previousCrc(6); xorBitMap(6)(72) := previousCrc(8); xorBitMap(6)(73) := previousCrc(9); xorBitMap(6)(74) := previousCrc(10); xorBitMap(6)(75) := previousCrc(11); xorBitMap(6)(77) := previousCrc(13); xorBitMap(6)(79) := previousCrc(15); xorBitMap(6)(82) := previousCrc(18); xorBitMap(6)(83) := previousCrc(19); xorBitMap(6)(84) := previousCrc(20); xorBitMap(6)(86) := previousCrc(22); xorBitMap(6)(87) := previousCrc(23); xorBitMap(6)(88) := previousCrc(24); xorBitMap(6)(92) := previousCrc(28); xorBitMap(6)(94) := previousCrc(30); 
      xorBitMap(7)(60) := currentData(60); xorBitMap(7)(58) := currentData(58); xorBitMap(7)(57) := currentData(57); xorBitMap(7)(56) := currentData(56); xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(64) := previousCrc(0); xorBitMap(7)(66) := previousCrc(2); xorBitMap(7)(69) := previousCrc(5); xorBitMap(7)(71) := previousCrc(7); xorBitMap(7)(73) := previousCrc(9); xorBitMap(7)(74) := previousCrc(10); xorBitMap(7)(75) := previousCrc(11); xorBitMap(7)(77) := previousCrc(13); xorBitMap(7)(78) := previousCrc(14); xorBitMap(7)(79) := previousCrc(15); xorBitMap(7)(82) := previousCrc(18); xorBitMap(7)(83) := previousCrc(19); xorBitMap(7)(84) := previousCrc(20); xorBitMap(7)(86) := previousCrc(22); xorBitMap(7)(88) := previousCrc(24); xorBitMap(7)(89) := previousCrc(25); xorBitMap(7)(90) := previousCrc(26); xorBitMap(7)(92) := previousCrc(28); 
      xorBitMap(8)(63) := currentData(63); xorBitMap(8)(60) := currentData(60); xorBitMap(8)(59) := currentData(59); xorBitMap(8)(57) := currentData(57); xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(64) := previousCrc(0); xorBitMap(8)(65) := previousCrc(1); xorBitMap(8)(66) := previousCrc(2); xorBitMap(8)(67) := previousCrc(3); xorBitMap(8)(69) := previousCrc(5); xorBitMap(8)(70) := previousCrc(6); xorBitMap(8)(72) := previousCrc(8); xorBitMap(8)(74) := previousCrc(10); xorBitMap(8)(75) := previousCrc(11); xorBitMap(8)(77) := previousCrc(13); xorBitMap(8)(78) := previousCrc(14); xorBitMap(8)(82) := previousCrc(18); xorBitMap(8)(83) := previousCrc(19); xorBitMap(8)(84) := previousCrc(20); xorBitMap(8)(86) := previousCrc(22); xorBitMap(8)(89) := previousCrc(25); xorBitMap(8)(91) := previousCrc(27); xorBitMap(8)(92) := previousCrc(28); xorBitMap(8)(95) := previousCrc(31); 
      xorBitMap(9)(61) := currentData(61); xorBitMap(9)(60) := currentData(60); xorBitMap(9)(58) := currentData(58); xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(64) := previousCrc(0); xorBitMap(9)(65) := previousCrc(1); xorBitMap(9)(66) := previousCrc(2); xorBitMap(9)(67) := previousCrc(3); xorBitMap(9)(68) := previousCrc(4); xorBitMap(9)(70) := previousCrc(6); xorBitMap(9)(71) := previousCrc(7); xorBitMap(9)(73) := previousCrc(9); xorBitMap(9)(75) := previousCrc(11); xorBitMap(9)(76) := previousCrc(12); xorBitMap(9)(78) := previousCrc(14); xorBitMap(9)(79) := previousCrc(15); xorBitMap(9)(83) := previousCrc(19); xorBitMap(9)(84) := previousCrc(20); xorBitMap(9)(85) := previousCrc(21); xorBitMap(9)(87) := previousCrc(23); xorBitMap(9)(90) := previousCrc(26); xorBitMap(9)(92) := previousCrc(28); xorBitMap(9)(93) := previousCrc(29); 
      xorBitMap(10)(63) := currentData(63); xorBitMap(10)(62) := currentData(62); xorBitMap(10)(60) := currentData(60); xorBitMap(10)(59) := currentData(59); xorBitMap(10)(58) := currentData(58); xorBitMap(10)(56) := currentData(56); xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(64) := previousCrc(0); xorBitMap(10)(65) := previousCrc(1); xorBitMap(10)(67) := previousCrc(3); xorBitMap(10)(68) := previousCrc(4); xorBitMap(10)(71) := previousCrc(7); xorBitMap(10)(72) := previousCrc(8); xorBitMap(10)(74) := previousCrc(10); xorBitMap(10)(82) := previousCrc(18); xorBitMap(10)(84) := previousCrc(20); xorBitMap(10)(87) := previousCrc(23); xorBitMap(10)(88) := previousCrc(24); xorBitMap(10)(90) := previousCrc(26); xorBitMap(10)(91) := previousCrc(27); xorBitMap(10)(92) := previousCrc(28); xorBitMap(10)(94) := previousCrc(30); xorBitMap(10)(95) := previousCrc(31); 
      xorBitMap(11)(59) := currentData(59); xorBitMap(11)(58) := currentData(58); xorBitMap(11)(57) := currentData(57); xorBitMap(11)(56) := currentData(56); xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(65) := previousCrc(1); xorBitMap(11)(68) := previousCrc(4); xorBitMap(11)(72) := previousCrc(8); xorBitMap(11)(73) := previousCrc(9); xorBitMap(11)(75) := previousCrc(11); xorBitMap(11)(76) := previousCrc(12); xorBitMap(11)(77) := previousCrc(13); xorBitMap(11)(79) := previousCrc(15); xorBitMap(11)(80) := previousCrc(16); xorBitMap(11)(82) := previousCrc(18); xorBitMap(11)(83) := previousCrc(19); xorBitMap(11)(86) := previousCrc(22); xorBitMap(11)(87) := previousCrc(23); xorBitMap(11)(88) := previousCrc(24); xorBitMap(11)(89) := previousCrc(25); xorBitMap(11)(90) := previousCrc(26); xorBitMap(11)(91) := previousCrc(27); 
      xorBitMap(12)(63) := currentData(63); xorBitMap(12)(61) := currentData(61); xorBitMap(12)(59) := currentData(59); xorBitMap(12)(57) := currentData(57); xorBitMap(12)(56) := currentData(56); xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(73) := previousCrc(9); xorBitMap(12)(74) := previousCrc(10); xorBitMap(12)(78) := previousCrc(14); xorBitMap(12)(79) := previousCrc(15); xorBitMap(12)(81) := previousCrc(17); xorBitMap(12)(82) := previousCrc(18); xorBitMap(12)(83) := previousCrc(19); xorBitMap(12)(84) := previousCrc(20); xorBitMap(12)(85) := previousCrc(21); xorBitMap(12)(86) := previousCrc(22); xorBitMap(12)(88) := previousCrc(24); xorBitMap(12)(89) := previousCrc(25); xorBitMap(12)(91) := previousCrc(27); xorBitMap(12)(93) := previousCrc(29); xorBitMap(12)(95) := previousCrc(31); 
      xorBitMap(13)(62) := currentData(62); xorBitMap(13)(60) := currentData(60); xorBitMap(13)(58) := currentData(58); xorBitMap(13)(57) := currentData(57); xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(64) := previousCrc(0); xorBitMap(13)(74) := previousCrc(10); xorBitMap(13)(75) := previousCrc(11); xorBitMap(13)(79) := previousCrc(15); xorBitMap(13)(80) := previousCrc(16); xorBitMap(13)(82) := previousCrc(18); xorBitMap(13)(83) := previousCrc(19); xorBitMap(13)(84) := previousCrc(20); xorBitMap(13)(85) := previousCrc(21); xorBitMap(13)(86) := previousCrc(22); xorBitMap(13)(87) := previousCrc(23); xorBitMap(13)(89) := previousCrc(25); xorBitMap(13)(90) := previousCrc(26); xorBitMap(13)(92) := previousCrc(28); xorBitMap(13)(94) := previousCrc(30); 
      xorBitMap(14)(63) := currentData(63); xorBitMap(14)(61) := currentData(61); xorBitMap(14)(59) := currentData(59); xorBitMap(14)(58) := currentData(58); xorBitMap(14)(56) := currentData(56); xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(64) := previousCrc(0); xorBitMap(14)(65) := previousCrc(1); xorBitMap(14)(75) := previousCrc(11); xorBitMap(14)(76) := previousCrc(12); xorBitMap(14)(80) := previousCrc(16); xorBitMap(14)(81) := previousCrc(17); xorBitMap(14)(83) := previousCrc(19); xorBitMap(14)(84) := previousCrc(20); xorBitMap(14)(85) := previousCrc(21); xorBitMap(14)(86) := previousCrc(22); xorBitMap(14)(87) := previousCrc(23); xorBitMap(14)(88) := previousCrc(24); xorBitMap(14)(90) := previousCrc(26); xorBitMap(14)(91) := previousCrc(27); xorBitMap(14)(93) := previousCrc(29); xorBitMap(14)(95) := previousCrc(31); 
      xorBitMap(15)(62) := currentData(62); xorBitMap(15)(60) := currentData(60); xorBitMap(15)(59) := currentData(59); xorBitMap(15)(57) := currentData(57); xorBitMap(15)(56) := currentData(56); xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(65) := previousCrc(1); xorBitMap(15)(66) := previousCrc(2); xorBitMap(15)(76) := previousCrc(12); xorBitMap(15)(77) := previousCrc(13); xorBitMap(15)(81) := previousCrc(17); xorBitMap(15)(82) := previousCrc(18); xorBitMap(15)(84) := previousCrc(20); xorBitMap(15)(85) := previousCrc(21); xorBitMap(15)(86) := previousCrc(22); xorBitMap(15)(87) := previousCrc(23); xorBitMap(15)(88) := previousCrc(24); xorBitMap(15)(89) := previousCrc(25); xorBitMap(15)(91) := previousCrc(27); xorBitMap(15)(92) := previousCrc(28); xorBitMap(15)(94) := previousCrc(30); 
      xorBitMap(16)(57) := currentData(57); xorBitMap(16)(56) := currentData(56); xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(64) := previousCrc(0); xorBitMap(16)(67) := previousCrc(3); xorBitMap(16)(69) := previousCrc(5); xorBitMap(16)(76) := previousCrc(12); xorBitMap(16)(78) := previousCrc(14); xorBitMap(16)(79) := previousCrc(15); xorBitMap(16)(80) := previousCrc(16); xorBitMap(16)(83) := previousCrc(19); xorBitMap(16)(88) := previousCrc(24); xorBitMap(16)(89) := previousCrc(25); 
      xorBitMap(17)(58) := currentData(58); xorBitMap(17)(57) := currentData(57); xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(65) := previousCrc(1); xorBitMap(17)(68) := previousCrc(4); xorBitMap(17)(70) := previousCrc(6); xorBitMap(17)(77) := previousCrc(13); xorBitMap(17)(79) := previousCrc(15); xorBitMap(17)(80) := previousCrc(16); xorBitMap(17)(81) := previousCrc(17); xorBitMap(17)(84) := previousCrc(20); xorBitMap(17)(89) := previousCrc(25); xorBitMap(17)(90) := previousCrc(26); 
      xorBitMap(18)(59) := currentData(59); xorBitMap(18)(58) := currentData(58); xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(64) := previousCrc(0); xorBitMap(18)(66) := previousCrc(2); xorBitMap(18)(69) := previousCrc(5); xorBitMap(18)(71) := previousCrc(7); xorBitMap(18)(78) := previousCrc(14); xorBitMap(18)(80) := previousCrc(16); xorBitMap(18)(81) := previousCrc(17); xorBitMap(18)(82) := previousCrc(18); xorBitMap(18)(85) := previousCrc(21); xorBitMap(18)(90) := previousCrc(26); xorBitMap(18)(91) := previousCrc(27); 
      xorBitMap(19)(60) := currentData(60); xorBitMap(19)(59) := currentData(59); xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(64) := previousCrc(0); xorBitMap(19)(65) := previousCrc(1); xorBitMap(19)(67) := previousCrc(3); xorBitMap(19)(70) := previousCrc(6); xorBitMap(19)(72) := previousCrc(8); xorBitMap(19)(79) := previousCrc(15); xorBitMap(19)(81) := previousCrc(17); xorBitMap(19)(82) := previousCrc(18); xorBitMap(19)(83) := previousCrc(19); xorBitMap(19)(86) := previousCrc(22); xorBitMap(19)(91) := previousCrc(27); xorBitMap(19)(92) := previousCrc(28); 
      xorBitMap(20)(61) := currentData(61); xorBitMap(20)(60) := currentData(60); xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(65) := previousCrc(1); xorBitMap(20)(66) := previousCrc(2); xorBitMap(20)(68) := previousCrc(4); xorBitMap(20)(71) := previousCrc(7); xorBitMap(20)(73) := previousCrc(9); xorBitMap(20)(80) := previousCrc(16); xorBitMap(20)(82) := previousCrc(18); xorBitMap(20)(83) := previousCrc(19); xorBitMap(20)(84) := previousCrc(20); xorBitMap(20)(87) := previousCrc(23); xorBitMap(20)(92) := previousCrc(28); xorBitMap(20)(93) := previousCrc(29); 
      xorBitMap(21)(62) := currentData(62); xorBitMap(21)(61) := currentData(61); xorBitMap(21)(56) := currentData(56); xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(66) := previousCrc(2); xorBitMap(21)(67) := previousCrc(3); xorBitMap(21)(69) := previousCrc(5); xorBitMap(21)(72) := previousCrc(8); xorBitMap(21)(74) := previousCrc(10); xorBitMap(21)(81) := previousCrc(17); xorBitMap(21)(83) := previousCrc(19); xorBitMap(21)(84) := previousCrc(20); xorBitMap(21)(85) := previousCrc(21); xorBitMap(21)(88) := previousCrc(24); xorBitMap(21)(93) := previousCrc(29); xorBitMap(21)(94) := previousCrc(30); 
      xorBitMap(22)(62) := currentData(62); xorBitMap(22)(61) := currentData(61); xorBitMap(22)(60) := currentData(60); xorBitMap(22)(58) := currentData(58); xorBitMap(22)(57) := currentData(57); xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(66) := previousCrc(2); xorBitMap(22)(67) := previousCrc(3); xorBitMap(22)(68) := previousCrc(4); xorBitMap(22)(69) := previousCrc(5); xorBitMap(22)(70) := previousCrc(6); xorBitMap(22)(73) := previousCrc(9); xorBitMap(22)(75) := previousCrc(11); xorBitMap(22)(76) := previousCrc(12); xorBitMap(22)(77) := previousCrc(13); xorBitMap(22)(79) := previousCrc(15); xorBitMap(22)(80) := previousCrc(16); xorBitMap(22)(84) := previousCrc(20); xorBitMap(22)(87) := previousCrc(23); xorBitMap(22)(89) := previousCrc(25); xorBitMap(22)(90) := previousCrc(26); xorBitMap(22)(92) := previousCrc(28); xorBitMap(22)(93) := previousCrc(29); xorBitMap(22)(94) := previousCrc(30); 
      xorBitMap(23)(62) := currentData(62); xorBitMap(23)(60) := currentData(60); xorBitMap(23)(59) := currentData(59); xorBitMap(23)(56) := currentData(56); xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(66) := previousCrc(2); xorBitMap(23)(67) := previousCrc(3); xorBitMap(23)(68) := previousCrc(4); xorBitMap(23)(70) := previousCrc(6); xorBitMap(23)(71) := previousCrc(7); xorBitMap(23)(74) := previousCrc(10); xorBitMap(23)(78) := previousCrc(14); xorBitMap(23)(79) := previousCrc(15); xorBitMap(23)(81) := previousCrc(17); xorBitMap(23)(82) := previousCrc(18); xorBitMap(23)(86) := previousCrc(22); xorBitMap(23)(87) := previousCrc(23); xorBitMap(23)(88) := previousCrc(24); xorBitMap(23)(91) := previousCrc(27); xorBitMap(23)(92) := previousCrc(28); xorBitMap(23)(94) := previousCrc(30); 
      xorBitMap(24)(63) := currentData(63); xorBitMap(24)(61) := currentData(61); xorBitMap(24)(60) := currentData(60); xorBitMap(24)(57) := currentData(57); xorBitMap(24)(56) := currentData(56); xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(64) := previousCrc(0); xorBitMap(24)(67) := previousCrc(3); xorBitMap(24)(68) := previousCrc(4); xorBitMap(24)(69) := previousCrc(5); xorBitMap(24)(71) := previousCrc(7); xorBitMap(24)(72) := previousCrc(8); xorBitMap(24)(75) := previousCrc(11); xorBitMap(24)(79) := previousCrc(15); xorBitMap(24)(80) := previousCrc(16); xorBitMap(24)(82) := previousCrc(18); xorBitMap(24)(83) := previousCrc(19); xorBitMap(24)(87) := previousCrc(23); xorBitMap(24)(88) := previousCrc(24); xorBitMap(24)(89) := previousCrc(25); xorBitMap(24)(92) := previousCrc(28); xorBitMap(24)(93) := previousCrc(29); xorBitMap(24)(95) := previousCrc(31); 
      xorBitMap(25)(62) := currentData(62); xorBitMap(25)(61) := currentData(61); xorBitMap(25)(58) := currentData(58); xorBitMap(25)(57) := currentData(57); xorBitMap(25)(56) := currentData(56); xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(65) := previousCrc(1); xorBitMap(25)(68) := previousCrc(4); xorBitMap(25)(69) := previousCrc(5); xorBitMap(25)(70) := previousCrc(6); xorBitMap(25)(72) := previousCrc(8); xorBitMap(25)(73) := previousCrc(9); xorBitMap(25)(76) := previousCrc(12); xorBitMap(25)(80) := previousCrc(16); xorBitMap(25)(81) := previousCrc(17); xorBitMap(25)(83) := previousCrc(19); xorBitMap(25)(84) := previousCrc(20); xorBitMap(25)(88) := previousCrc(24); xorBitMap(25)(89) := previousCrc(25); xorBitMap(25)(90) := previousCrc(26); xorBitMap(25)(93) := previousCrc(29); xorBitMap(25)(94) := previousCrc(30); 
      xorBitMap(26)(62) := currentData(62); xorBitMap(26)(61) := currentData(61); xorBitMap(26)(60) := currentData(60); xorBitMap(26)(59) := currentData(59); xorBitMap(26)(57) := currentData(57); xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(70) := previousCrc(6); xorBitMap(26)(71) := previousCrc(7); xorBitMap(26)(73) := previousCrc(9); xorBitMap(26)(74) := previousCrc(10); xorBitMap(26)(76) := previousCrc(12); xorBitMap(26)(79) := previousCrc(15); xorBitMap(26)(80) := previousCrc(16); xorBitMap(26)(81) := previousCrc(17); xorBitMap(26)(84) := previousCrc(20); xorBitMap(26)(86) := previousCrc(22); xorBitMap(26)(87) := previousCrc(23); xorBitMap(26)(89) := previousCrc(25); xorBitMap(26)(91) := previousCrc(27); xorBitMap(26)(92) := previousCrc(28); xorBitMap(26)(93) := previousCrc(29); xorBitMap(26)(94) := previousCrc(30); 
      xorBitMap(27)(63) := currentData(63); xorBitMap(27)(62) := currentData(62); xorBitMap(27)(61) := currentData(61); xorBitMap(27)(60) := currentData(60); xorBitMap(27)(58) := currentData(58); xorBitMap(27)(56) := currentData(56); xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(64) := previousCrc(0); xorBitMap(27)(71) := previousCrc(7); xorBitMap(27)(72) := previousCrc(8); xorBitMap(27)(74) := previousCrc(10); xorBitMap(27)(75) := previousCrc(11); xorBitMap(27)(77) := previousCrc(13); xorBitMap(27)(80) := previousCrc(16); xorBitMap(27)(81) := previousCrc(17); xorBitMap(27)(82) := previousCrc(18); xorBitMap(27)(85) := previousCrc(21); xorBitMap(27)(87) := previousCrc(23); xorBitMap(27)(88) := previousCrc(24); xorBitMap(27)(90) := previousCrc(26); xorBitMap(27)(92) := previousCrc(28); xorBitMap(27)(93) := previousCrc(29); xorBitMap(27)(94) := previousCrc(30); xorBitMap(27)(95) := previousCrc(31); 
      xorBitMap(28)(63) := currentData(63); xorBitMap(28)(62) := currentData(62); xorBitMap(28)(61) := currentData(61); xorBitMap(28)(59) := currentData(59); xorBitMap(28)(57) := currentData(57); xorBitMap(28)(56) := currentData(56); xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(65) := previousCrc(1); xorBitMap(28)(72) := previousCrc(8); xorBitMap(28)(73) := previousCrc(9); xorBitMap(28)(75) := previousCrc(11); xorBitMap(28)(76) := previousCrc(12); xorBitMap(28)(78) := previousCrc(14); xorBitMap(28)(81) := previousCrc(17); xorBitMap(28)(82) := previousCrc(18); xorBitMap(28)(83) := previousCrc(19); xorBitMap(28)(86) := previousCrc(22); xorBitMap(28)(88) := previousCrc(24); xorBitMap(28)(89) := previousCrc(25); xorBitMap(28)(91) := previousCrc(27); xorBitMap(28)(93) := previousCrc(29); xorBitMap(28)(94) := previousCrc(30); xorBitMap(28)(95) := previousCrc(31); 
      xorBitMap(29)(63) := currentData(63); xorBitMap(29)(62) := currentData(62); xorBitMap(29)(60) := currentData(60); xorBitMap(29)(58) := currentData(58); xorBitMap(29)(57) := currentData(57); xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(66) := previousCrc(2); xorBitMap(29)(73) := previousCrc(9); xorBitMap(29)(74) := previousCrc(10); xorBitMap(29)(76) := previousCrc(12); xorBitMap(29)(77) := previousCrc(13); xorBitMap(29)(79) := previousCrc(15); xorBitMap(29)(82) := previousCrc(18); xorBitMap(29)(83) := previousCrc(19); xorBitMap(29)(84) := previousCrc(20); xorBitMap(29)(87) := previousCrc(23); xorBitMap(29)(89) := previousCrc(25); xorBitMap(29)(90) := previousCrc(26); xorBitMap(29)(92) := previousCrc(28); xorBitMap(29)(94) := previousCrc(30); xorBitMap(29)(95) := previousCrc(31); 
      xorBitMap(30)(63) := currentData(63); xorBitMap(30)(61) := currentData(61); xorBitMap(30)(59) := currentData(59); xorBitMap(30)(58) := currentData(58); xorBitMap(30)(56) := currentData(56); xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(64) := previousCrc(0); xorBitMap(30)(67) := previousCrc(3); xorBitMap(30)(74) := previousCrc(10); xorBitMap(30)(75) := previousCrc(11); xorBitMap(30)(77) := previousCrc(13); xorBitMap(30)(78) := previousCrc(14); xorBitMap(30)(80) := previousCrc(16); xorBitMap(30)(83) := previousCrc(19); xorBitMap(30)(84) := previousCrc(20); xorBitMap(30)(85) := previousCrc(21); xorBitMap(30)(88) := previousCrc(24); xorBitMap(30)(90) := previousCrc(26); xorBitMap(30)(91) := previousCrc(27); xorBitMap(30)(93) := previousCrc(29); xorBitMap(30)(95) := previousCrc(31); 
      xorBitMap(31)(62) := currentData(62); xorBitMap(31)(60) := currentData(60); xorBitMap(31)(59) := currentData(59); xorBitMap(31)(57) := currentData(57); xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(65) := previousCrc(1); xorBitMap(31)(68) := previousCrc(4); xorBitMap(31)(75) := previousCrc(11); xorBitMap(31)(76) := previousCrc(12); xorBitMap(31)(78) := previousCrc(14); xorBitMap(31)(79) := previousCrc(15); xorBitMap(31)(81) := previousCrc(17); xorBitMap(31)(84) := previousCrc(20); xorBitMap(31)(85) := previousCrc(21); xorBitMap(31)(86) := previousCrc(22); xorBitMap(31)(89) := previousCrc(25); xorBitMap(31)(91) := previousCrc(27); xorBitMap(31)(92) := previousCrc(28); xorBitMap(31)(94) := previousCrc(30); 
   end procedure;

   procedure xorBitMap1Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(7 downto 0)) is 
   begin
      xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(184) := previousCrc(24); xorBitMap(0)(190) := previousCrc(30); 
      xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(184) := previousCrc(24); xorBitMap(1)(185) := previousCrc(25); xorBitMap(1)(190) := previousCrc(30); xorBitMap(1)(191) := previousCrc(31); 
      xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(184) := previousCrc(24); xorBitMap(2)(185) := previousCrc(25); xorBitMap(2)(186) := previousCrc(26); xorBitMap(2)(190) := previousCrc(30); xorBitMap(2)(191) := previousCrc(31); 
      xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(185) := previousCrc(25); xorBitMap(3)(186) := previousCrc(26); xorBitMap(3)(187) := previousCrc(27); xorBitMap(3)(191) := previousCrc(31); 
      xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(184) := previousCrc(24); xorBitMap(4)(186) := previousCrc(26); xorBitMap(4)(187) := previousCrc(27); xorBitMap(4)(188) := previousCrc(28); xorBitMap(4)(190) := previousCrc(30); 
      xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(184) := previousCrc(24); xorBitMap(5)(185) := previousCrc(25); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(188) := previousCrc(28); xorBitMap(5)(189) := previousCrc(29); xorBitMap(5)(190) := previousCrc(30); xorBitMap(5)(191) := previousCrc(31); 
      xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(185) := previousCrc(25); xorBitMap(6)(186) := previousCrc(26); xorBitMap(6)(188) := previousCrc(28); xorBitMap(6)(189) := previousCrc(29); xorBitMap(6)(190) := previousCrc(30); xorBitMap(6)(191) := previousCrc(31); 
      xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(184) := previousCrc(24); xorBitMap(7)(186) := previousCrc(26); xorBitMap(7)(187) := previousCrc(27); xorBitMap(7)(189) := previousCrc(29); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(160) := previousCrc(0); xorBitMap(8)(184) := previousCrc(24); xorBitMap(8)(185) := previousCrc(25); xorBitMap(8)(187) := previousCrc(27); xorBitMap(8)(188) := previousCrc(28); 
      xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(161) := previousCrc(1); xorBitMap(9)(185) := previousCrc(25); xorBitMap(9)(186) := previousCrc(26); xorBitMap(9)(188) := previousCrc(28); xorBitMap(9)(189) := previousCrc(29); 
      xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(162) := previousCrc(2); xorBitMap(10)(184) := previousCrc(24); xorBitMap(10)(186) := previousCrc(26); xorBitMap(10)(187) := previousCrc(27); xorBitMap(10)(189) := previousCrc(29); 
      xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(163) := previousCrc(3); xorBitMap(11)(184) := previousCrc(24); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(187) := previousCrc(27); xorBitMap(11)(188) := previousCrc(28); 
      xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(164) := previousCrc(4); xorBitMap(12)(184) := previousCrc(24); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(186) := previousCrc(26); xorBitMap(12)(188) := previousCrc(28); xorBitMap(12)(189) := previousCrc(29); xorBitMap(12)(190) := previousCrc(30); 
      xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(165) := previousCrc(5); xorBitMap(13)(185) := previousCrc(25); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(187) := previousCrc(27); xorBitMap(13)(189) := previousCrc(29); xorBitMap(13)(190) := previousCrc(30); xorBitMap(13)(191) := previousCrc(31); 
      xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(166) := previousCrc(6); xorBitMap(14)(186) := previousCrc(26); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(188) := previousCrc(28); xorBitMap(14)(190) := previousCrc(30); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(167) := previousCrc(7); xorBitMap(15)(187) := previousCrc(27); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(189) := previousCrc(29); xorBitMap(15)(191) := previousCrc(31); 
      xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(168) := previousCrc(8); xorBitMap(16)(184) := previousCrc(24); xorBitMap(16)(188) := previousCrc(28); xorBitMap(16)(189) := previousCrc(29); 
      xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(169) := previousCrc(9); xorBitMap(17)(185) := previousCrc(25); xorBitMap(17)(189) := previousCrc(29); xorBitMap(17)(190) := previousCrc(30); 
      xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(170) := previousCrc(10); xorBitMap(18)(186) := previousCrc(26); xorBitMap(18)(190) := previousCrc(30); xorBitMap(18)(191) := previousCrc(31); 
      xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(171) := previousCrc(11); xorBitMap(19)(187) := previousCrc(27); xorBitMap(19)(191) := previousCrc(31); 
      xorBitMap(20)(4) := currentData(4); xorBitMap(20)(172) := previousCrc(12); xorBitMap(20)(188) := previousCrc(28); 
      xorBitMap(21)(5) := currentData(5); xorBitMap(21)(173) := previousCrc(13); xorBitMap(21)(189) := previousCrc(29); 
      xorBitMap(22)(0) := currentData(0); xorBitMap(22)(174) := previousCrc(14); xorBitMap(22)(184) := previousCrc(24); 
      xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(175) := previousCrc(15); xorBitMap(23)(184) := previousCrc(24); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(190) := previousCrc(30); 
      xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(176) := previousCrc(16); xorBitMap(24)(185) := previousCrc(25); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(191) := previousCrc(31); 
      xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(177) := previousCrc(17); xorBitMap(25)(186) := previousCrc(26); xorBitMap(25)(187) := previousCrc(27); 
      xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(178) := previousCrc(18); xorBitMap(26)(184) := previousCrc(24); xorBitMap(26)(187) := previousCrc(27); xorBitMap(26)(188) := previousCrc(28); xorBitMap(26)(190) := previousCrc(30); 
      xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(179) := previousCrc(19); xorBitMap(27)(185) := previousCrc(25); xorBitMap(27)(188) := previousCrc(28); xorBitMap(27)(189) := previousCrc(29); xorBitMap(27)(191) := previousCrc(31); 
      xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(180) := previousCrc(20); xorBitMap(28)(186) := previousCrc(26); xorBitMap(28)(189) := previousCrc(29); xorBitMap(28)(190) := previousCrc(30); 
      xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(181) := previousCrc(21); xorBitMap(29)(187) := previousCrc(27); xorBitMap(29)(190) := previousCrc(30); xorBitMap(29)(191) := previousCrc(31); 
      xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(182) := previousCrc(22); xorBitMap(30)(188) := previousCrc(28); xorBitMap(30)(191) := previousCrc(31); 
      xorBitMap(31)(5) := currentData(5); xorBitMap(31)(183) := previousCrc(23); xorBitMap(31)(189) := previousCrc(29); 
   end procedure;

   procedure xorBitMap2Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(15 downto 0)) is 
   begin
      xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(176) := previousCrc(16); xorBitMap(0)(182) := previousCrc(22); xorBitMap(0)(185) := previousCrc(25); xorBitMap(0)(186) := previousCrc(26); xorBitMap(0)(188) := previousCrc(28); 
      xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(176) := previousCrc(16); xorBitMap(1)(177) := previousCrc(17); xorBitMap(1)(182) := previousCrc(22); xorBitMap(1)(183) := previousCrc(23); xorBitMap(1)(185) := previousCrc(25); xorBitMap(1)(187) := previousCrc(27); xorBitMap(1)(188) := previousCrc(28); xorBitMap(1)(189) := previousCrc(29); 
      xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(176) := previousCrc(16); xorBitMap(2)(177) := previousCrc(17); xorBitMap(2)(178) := previousCrc(18); xorBitMap(2)(182) := previousCrc(22); xorBitMap(2)(183) := previousCrc(23); xorBitMap(2)(184) := previousCrc(24); xorBitMap(2)(185) := previousCrc(25); xorBitMap(2)(189) := previousCrc(29); xorBitMap(2)(190) := previousCrc(30); 
      xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(177) := previousCrc(17); xorBitMap(3)(178) := previousCrc(18); xorBitMap(3)(179) := previousCrc(19); xorBitMap(3)(183) := previousCrc(23); xorBitMap(3)(184) := previousCrc(24); xorBitMap(3)(185) := previousCrc(25); xorBitMap(3)(186) := previousCrc(26); xorBitMap(3)(190) := previousCrc(30); xorBitMap(3)(191) := previousCrc(31); 
      xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(176) := previousCrc(16); xorBitMap(4)(178) := previousCrc(18); xorBitMap(4)(179) := previousCrc(19); xorBitMap(4)(180) := previousCrc(20); xorBitMap(4)(182) := previousCrc(22); xorBitMap(4)(184) := previousCrc(24); xorBitMap(4)(187) := previousCrc(27); xorBitMap(4)(188) := previousCrc(28); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(176) := previousCrc(16); xorBitMap(5)(177) := previousCrc(17); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(180) := previousCrc(20); xorBitMap(5)(181) := previousCrc(21); xorBitMap(5)(182) := previousCrc(22); xorBitMap(5)(183) := previousCrc(23); xorBitMap(5)(186) := previousCrc(26); xorBitMap(5)(189) := previousCrc(29); 
      xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(177) := previousCrc(17); xorBitMap(6)(178) := previousCrc(18); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(181) := previousCrc(21); xorBitMap(6)(182) := previousCrc(22); xorBitMap(6)(183) := previousCrc(23); xorBitMap(6)(184) := previousCrc(24); xorBitMap(6)(187) := previousCrc(27); xorBitMap(6)(190) := previousCrc(30); 
      xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(176) := previousCrc(16); xorBitMap(7)(178) := previousCrc(18); xorBitMap(7)(179) := previousCrc(19); xorBitMap(7)(181) := previousCrc(21); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(184) := previousCrc(24); xorBitMap(7)(186) := previousCrc(26); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(176) := previousCrc(16); xorBitMap(8)(177) := previousCrc(17); xorBitMap(8)(179) := previousCrc(19); xorBitMap(8)(180) := previousCrc(20); xorBitMap(8)(184) := previousCrc(24); xorBitMap(8)(186) := previousCrc(26); xorBitMap(8)(187) := previousCrc(27); xorBitMap(8)(188) := previousCrc(28); 
      xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(177) := previousCrc(17); xorBitMap(9)(178) := previousCrc(18); xorBitMap(9)(180) := previousCrc(20); xorBitMap(9)(181) := previousCrc(21); xorBitMap(9)(185) := previousCrc(25); xorBitMap(9)(187) := previousCrc(27); xorBitMap(9)(188) := previousCrc(28); xorBitMap(9)(189) := previousCrc(29); 
      xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(176) := previousCrc(16); xorBitMap(10)(178) := previousCrc(18); xorBitMap(10)(179) := previousCrc(19); xorBitMap(10)(181) := previousCrc(21); xorBitMap(10)(185) := previousCrc(25); xorBitMap(10)(189) := previousCrc(29); xorBitMap(10)(190) := previousCrc(30); 
      xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(176) := previousCrc(16); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(179) := previousCrc(19); xorBitMap(11)(180) := previousCrc(20); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(188) := previousCrc(28); xorBitMap(11)(190) := previousCrc(30); xorBitMap(11)(191) := previousCrc(31); 
      xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(176) := previousCrc(16); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(178) := previousCrc(18); xorBitMap(12)(180) := previousCrc(20); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(182) := previousCrc(22); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(188) := previousCrc(28); xorBitMap(12)(189) := previousCrc(29); xorBitMap(12)(191) := previousCrc(31); 
      xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(177) := previousCrc(17); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(179) := previousCrc(19); xorBitMap(13)(181) := previousCrc(21); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(183) := previousCrc(23); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(189) := previousCrc(29); xorBitMap(13)(190) := previousCrc(30); 
      xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(178) := previousCrc(18); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(180) := previousCrc(20); xorBitMap(14)(182) := previousCrc(22); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(184) := previousCrc(24); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(190) := previousCrc(30); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(179) := previousCrc(19); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(181) := previousCrc(21); xorBitMap(15)(183) := previousCrc(23); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(185) := previousCrc(25); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(191) := previousCrc(31); 
      xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(160) := previousCrc(0); xorBitMap(16)(176) := previousCrc(16); xorBitMap(16)(180) := previousCrc(20); xorBitMap(16)(181) := previousCrc(21); xorBitMap(16)(184) := previousCrc(24); xorBitMap(16)(188) := previousCrc(28); xorBitMap(16)(189) := previousCrc(29); 
      xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(161) := previousCrc(1); xorBitMap(17)(177) := previousCrc(17); xorBitMap(17)(181) := previousCrc(21); xorBitMap(17)(182) := previousCrc(22); xorBitMap(17)(185) := previousCrc(25); xorBitMap(17)(189) := previousCrc(29); xorBitMap(17)(190) := previousCrc(30); 
      xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(162) := previousCrc(2); xorBitMap(18)(178) := previousCrc(18); xorBitMap(18)(182) := previousCrc(22); xorBitMap(18)(183) := previousCrc(23); xorBitMap(18)(186) := previousCrc(26); xorBitMap(18)(190) := previousCrc(30); xorBitMap(18)(191) := previousCrc(31); 
      xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(163) := previousCrc(3); xorBitMap(19)(179) := previousCrc(19); xorBitMap(19)(183) := previousCrc(23); xorBitMap(19)(184) := previousCrc(24); xorBitMap(19)(187) := previousCrc(27); xorBitMap(19)(191) := previousCrc(31); 
      xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(164) := previousCrc(4); xorBitMap(20)(180) := previousCrc(20); xorBitMap(20)(184) := previousCrc(24); xorBitMap(20)(185) := previousCrc(25); xorBitMap(20)(188) := previousCrc(28); 
      xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(165) := previousCrc(5); xorBitMap(21)(181) := previousCrc(21); xorBitMap(21)(185) := previousCrc(25); xorBitMap(21)(186) := previousCrc(26); xorBitMap(21)(189) := previousCrc(29); 
      xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(166) := previousCrc(6); xorBitMap(22)(176) := previousCrc(16); xorBitMap(22)(185) := previousCrc(25); xorBitMap(22)(187) := previousCrc(27); xorBitMap(22)(188) := previousCrc(28); xorBitMap(22)(190) := previousCrc(30); 
      xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(167) := previousCrc(7); xorBitMap(23)(176) := previousCrc(16); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(182) := previousCrc(22); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(189) := previousCrc(29); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(168) := previousCrc(8); xorBitMap(24)(177) := previousCrc(17); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(183) := previousCrc(23); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(190) := previousCrc(30); 
      xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(169) := previousCrc(9); xorBitMap(25)(178) := previousCrc(18); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(184) := previousCrc(24); xorBitMap(25)(187) := previousCrc(27); xorBitMap(25)(191) := previousCrc(31); 
      xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(170) := previousCrc(10); xorBitMap(26)(176) := previousCrc(16); xorBitMap(26)(179) := previousCrc(19); xorBitMap(26)(180) := previousCrc(20); xorBitMap(26)(182) := previousCrc(22); xorBitMap(26)(186) := previousCrc(26); 
      xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(171) := previousCrc(11); xorBitMap(27)(177) := previousCrc(17); xorBitMap(27)(180) := previousCrc(20); xorBitMap(27)(181) := previousCrc(21); xorBitMap(27)(183) := previousCrc(23); xorBitMap(27)(187) := previousCrc(27); 
      xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(172) := previousCrc(12); xorBitMap(28)(178) := previousCrc(18); xorBitMap(28)(181) := previousCrc(21); xorBitMap(28)(182) := previousCrc(22); xorBitMap(28)(184) := previousCrc(24); xorBitMap(28)(188) := previousCrc(28); 
      xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(173) := previousCrc(13); xorBitMap(29)(179) := previousCrc(19); xorBitMap(29)(182) := previousCrc(22); xorBitMap(29)(183) := previousCrc(23); xorBitMap(29)(185) := previousCrc(25); xorBitMap(29)(189) := previousCrc(29); 
      xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(174) := previousCrc(14); xorBitMap(30)(180) := previousCrc(20); xorBitMap(30)(183) := previousCrc(23); xorBitMap(30)(184) := previousCrc(24); xorBitMap(30)(186) := previousCrc(26); xorBitMap(30)(190) := previousCrc(30); 
      xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(175) := previousCrc(15); xorBitMap(31)(181) := previousCrc(21); xorBitMap(31)(184) := previousCrc(24); xorBitMap(31)(185) := previousCrc(25); xorBitMap(31)(187) := previousCrc(27); xorBitMap(31)(191) := previousCrc(31); 
   end procedure;

   procedure xorBitMap3Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(23 downto 0)) is 
   begin
      xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(168) := previousCrc(8); xorBitMap(0)(174) := previousCrc(14); xorBitMap(0)(177) := previousCrc(17); xorBitMap(0)(178) := previousCrc(18); xorBitMap(0)(180) := previousCrc(20); xorBitMap(0)(184) := previousCrc(24); 
      xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(168) := previousCrc(8); xorBitMap(1)(169) := previousCrc(9); xorBitMap(1)(174) := previousCrc(14); xorBitMap(1)(175) := previousCrc(15); xorBitMap(1)(177) := previousCrc(17); xorBitMap(1)(179) := previousCrc(19); xorBitMap(1)(180) := previousCrc(20); xorBitMap(1)(181) := previousCrc(21); xorBitMap(1)(184) := previousCrc(24); xorBitMap(1)(185) := previousCrc(25); 
      xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(168) := previousCrc(8); xorBitMap(2)(169) := previousCrc(9); xorBitMap(2)(170) := previousCrc(10); xorBitMap(2)(174) := previousCrc(14); xorBitMap(2)(175) := previousCrc(15); xorBitMap(2)(176) := previousCrc(16); xorBitMap(2)(177) := previousCrc(17); xorBitMap(2)(181) := previousCrc(21); xorBitMap(2)(182) := previousCrc(22); xorBitMap(2)(184) := previousCrc(24); xorBitMap(2)(185) := previousCrc(25); xorBitMap(2)(186) := previousCrc(26); 
      xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(169) := previousCrc(9); xorBitMap(3)(170) := previousCrc(10); xorBitMap(3)(171) := previousCrc(11); xorBitMap(3)(175) := previousCrc(15); xorBitMap(3)(176) := previousCrc(16); xorBitMap(3)(177) := previousCrc(17); xorBitMap(3)(178) := previousCrc(18); xorBitMap(3)(182) := previousCrc(22); xorBitMap(3)(183) := previousCrc(23); xorBitMap(3)(185) := previousCrc(25); xorBitMap(3)(186) := previousCrc(26); xorBitMap(3)(187) := previousCrc(27); 
      xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(168) := previousCrc(8); xorBitMap(4)(170) := previousCrc(10); xorBitMap(4)(171) := previousCrc(11); xorBitMap(4)(172) := previousCrc(12); xorBitMap(4)(174) := previousCrc(14); xorBitMap(4)(176) := previousCrc(16); xorBitMap(4)(179) := previousCrc(19); xorBitMap(4)(180) := previousCrc(20); xorBitMap(4)(183) := previousCrc(23); xorBitMap(4)(186) := previousCrc(26); xorBitMap(4)(187) := previousCrc(27); xorBitMap(4)(188) := previousCrc(28); 
      xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(168) := previousCrc(8); xorBitMap(5)(169) := previousCrc(9); xorBitMap(5)(171) := previousCrc(11); xorBitMap(5)(172) := previousCrc(12); xorBitMap(5)(173) := previousCrc(13); xorBitMap(5)(174) := previousCrc(14); xorBitMap(5)(175) := previousCrc(15); xorBitMap(5)(178) := previousCrc(18); xorBitMap(5)(181) := previousCrc(21); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(188) := previousCrc(28); xorBitMap(5)(189) := previousCrc(29); 
      xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(169) := previousCrc(9); xorBitMap(6)(170) := previousCrc(10); xorBitMap(6)(172) := previousCrc(12); xorBitMap(6)(173) := previousCrc(13); xorBitMap(6)(174) := previousCrc(14); xorBitMap(6)(175) := previousCrc(15); xorBitMap(6)(176) := previousCrc(16); xorBitMap(6)(179) := previousCrc(19); xorBitMap(6)(182) := previousCrc(22); xorBitMap(6)(188) := previousCrc(28); xorBitMap(6)(189) := previousCrc(29); xorBitMap(6)(190) := previousCrc(30); 
      xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(168) := previousCrc(8); xorBitMap(7)(170) := previousCrc(10); xorBitMap(7)(171) := previousCrc(11); xorBitMap(7)(173) := previousCrc(13); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(176) := previousCrc(16); xorBitMap(7)(178) := previousCrc(18); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(184) := previousCrc(24); xorBitMap(7)(189) := previousCrc(29); xorBitMap(7)(190) := previousCrc(30); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(168) := previousCrc(8); xorBitMap(8)(169) := previousCrc(9); xorBitMap(8)(171) := previousCrc(11); xorBitMap(8)(172) := previousCrc(12); xorBitMap(8)(176) := previousCrc(16); xorBitMap(8)(178) := previousCrc(18); xorBitMap(8)(179) := previousCrc(19); xorBitMap(8)(180) := previousCrc(20); xorBitMap(8)(185) := previousCrc(25); xorBitMap(8)(190) := previousCrc(30); xorBitMap(8)(191) := previousCrc(31); 
      xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(169) := previousCrc(9); xorBitMap(9)(170) := previousCrc(10); xorBitMap(9)(172) := previousCrc(12); xorBitMap(9)(173) := previousCrc(13); xorBitMap(9)(177) := previousCrc(17); xorBitMap(9)(179) := previousCrc(19); xorBitMap(9)(180) := previousCrc(20); xorBitMap(9)(181) := previousCrc(21); xorBitMap(9)(186) := previousCrc(26); xorBitMap(9)(191) := previousCrc(31); 
      xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(168) := previousCrc(8); xorBitMap(10)(170) := previousCrc(10); xorBitMap(10)(171) := previousCrc(11); xorBitMap(10)(173) := previousCrc(13); xorBitMap(10)(177) := previousCrc(17); xorBitMap(10)(181) := previousCrc(21); xorBitMap(10)(182) := previousCrc(22); xorBitMap(10)(184) := previousCrc(24); xorBitMap(10)(187) := previousCrc(27); 
      xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(168) := previousCrc(8); xorBitMap(11)(169) := previousCrc(9); xorBitMap(11)(171) := previousCrc(11); xorBitMap(11)(172) := previousCrc(12); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(180) := previousCrc(20); xorBitMap(11)(182) := previousCrc(22); xorBitMap(11)(183) := previousCrc(23); xorBitMap(11)(184) := previousCrc(24); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(188) := previousCrc(28); 
      xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(168) := previousCrc(8); xorBitMap(12)(169) := previousCrc(9); xorBitMap(12)(170) := previousCrc(10); xorBitMap(12)(172) := previousCrc(12); xorBitMap(12)(173) := previousCrc(13); xorBitMap(12)(174) := previousCrc(14); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(180) := previousCrc(20); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(183) := previousCrc(23); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(186) := previousCrc(26); xorBitMap(12)(189) := previousCrc(29); 
      xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(169) := previousCrc(9); xorBitMap(13)(170) := previousCrc(10); xorBitMap(13)(171) := previousCrc(11); xorBitMap(13)(173) := previousCrc(13); xorBitMap(13)(174) := previousCrc(14); xorBitMap(13)(175) := previousCrc(15); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(181) := previousCrc(21); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(184) := previousCrc(24); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(187) := previousCrc(27); xorBitMap(13)(190) := previousCrc(30); 
      xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(170) := previousCrc(10); xorBitMap(14)(171) := previousCrc(11); xorBitMap(14)(172) := previousCrc(12); xorBitMap(14)(174) := previousCrc(14); xorBitMap(14)(175) := previousCrc(15); xorBitMap(14)(176) := previousCrc(16); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(182) := previousCrc(22); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(185) := previousCrc(25); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(188) := previousCrc(28); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(171) := previousCrc(11); xorBitMap(15)(172) := previousCrc(12); xorBitMap(15)(173) := previousCrc(13); xorBitMap(15)(175) := previousCrc(15); xorBitMap(15)(176) := previousCrc(16); xorBitMap(15)(177) := previousCrc(17); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(183) := previousCrc(23); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(186) := previousCrc(26); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(189) := previousCrc(29); 
      xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(168) := previousCrc(8); xorBitMap(16)(172) := previousCrc(12); xorBitMap(16)(173) := previousCrc(13); xorBitMap(16)(176) := previousCrc(16); xorBitMap(16)(180) := previousCrc(20); xorBitMap(16)(181) := previousCrc(21); xorBitMap(16)(185) := previousCrc(25); xorBitMap(16)(187) := previousCrc(27); xorBitMap(16)(189) := previousCrc(29); xorBitMap(16)(190) := previousCrc(30); 
      xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(169) := previousCrc(9); xorBitMap(17)(173) := previousCrc(13); xorBitMap(17)(174) := previousCrc(14); xorBitMap(17)(177) := previousCrc(17); xorBitMap(17)(181) := previousCrc(21); xorBitMap(17)(182) := previousCrc(22); xorBitMap(17)(186) := previousCrc(26); xorBitMap(17)(188) := previousCrc(28); xorBitMap(17)(190) := previousCrc(30); xorBitMap(17)(191) := previousCrc(31); 
      xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(170) := previousCrc(10); xorBitMap(18)(174) := previousCrc(14); xorBitMap(18)(175) := previousCrc(15); xorBitMap(18)(178) := previousCrc(18); xorBitMap(18)(182) := previousCrc(22); xorBitMap(18)(183) := previousCrc(23); xorBitMap(18)(187) := previousCrc(27); xorBitMap(18)(189) := previousCrc(29); xorBitMap(18)(191) := previousCrc(31); 
      xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(171) := previousCrc(11); xorBitMap(19)(175) := previousCrc(15); xorBitMap(19)(176) := previousCrc(16); xorBitMap(19)(179) := previousCrc(19); xorBitMap(19)(183) := previousCrc(23); xorBitMap(19)(184) := previousCrc(24); xorBitMap(19)(188) := previousCrc(28); xorBitMap(19)(190) := previousCrc(30); 
      xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(172) := previousCrc(12); xorBitMap(20)(176) := previousCrc(16); xorBitMap(20)(177) := previousCrc(17); xorBitMap(20)(180) := previousCrc(20); xorBitMap(20)(184) := previousCrc(24); xorBitMap(20)(185) := previousCrc(25); xorBitMap(20)(189) := previousCrc(29); xorBitMap(20)(191) := previousCrc(31); 
      xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(173) := previousCrc(13); xorBitMap(21)(177) := previousCrc(17); xorBitMap(21)(178) := previousCrc(18); xorBitMap(21)(181) := previousCrc(21); xorBitMap(21)(185) := previousCrc(25); xorBitMap(21)(186) := previousCrc(26); xorBitMap(21)(190) := previousCrc(30); 
      xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(168) := previousCrc(8); xorBitMap(22)(177) := previousCrc(17); xorBitMap(22)(179) := previousCrc(19); xorBitMap(22)(180) := previousCrc(20); xorBitMap(22)(182) := previousCrc(22); xorBitMap(22)(184) := previousCrc(24); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(187) := previousCrc(27); xorBitMap(22)(191) := previousCrc(31); 
      xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(168) := previousCrc(8); xorBitMap(23)(169) := previousCrc(9); xorBitMap(23)(174) := previousCrc(14); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(181) := previousCrc(21); xorBitMap(23)(183) := previousCrc(23); xorBitMap(23)(184) := previousCrc(24); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(187) := previousCrc(27); xorBitMap(23)(188) := previousCrc(28); 
      xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(160) := previousCrc(0); xorBitMap(24)(169) := previousCrc(9); xorBitMap(24)(170) := previousCrc(10); xorBitMap(24)(175) := previousCrc(15); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(182) := previousCrc(22); xorBitMap(24)(184) := previousCrc(24); xorBitMap(24)(185) := previousCrc(25); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(188) := previousCrc(28); xorBitMap(24)(189) := previousCrc(29); 
      xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(161) := previousCrc(1); xorBitMap(25)(170) := previousCrc(10); xorBitMap(25)(171) := previousCrc(11); xorBitMap(25)(176) := previousCrc(16); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(183) := previousCrc(23); xorBitMap(25)(185) := previousCrc(25); xorBitMap(25)(186) := previousCrc(26); xorBitMap(25)(187) := previousCrc(27); xorBitMap(25)(189) := previousCrc(29); xorBitMap(25)(190) := previousCrc(30); 
      xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(162) := previousCrc(2); xorBitMap(26)(168) := previousCrc(8); xorBitMap(26)(171) := previousCrc(11); xorBitMap(26)(172) := previousCrc(12); xorBitMap(26)(174) := previousCrc(14); xorBitMap(26)(178) := previousCrc(18); xorBitMap(26)(186) := previousCrc(26); xorBitMap(26)(187) := previousCrc(27); xorBitMap(26)(188) := previousCrc(28); xorBitMap(26)(190) := previousCrc(30); xorBitMap(26)(191) := previousCrc(31); 
      xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(163) := previousCrc(3); xorBitMap(27)(169) := previousCrc(9); xorBitMap(27)(172) := previousCrc(12); xorBitMap(27)(173) := previousCrc(13); xorBitMap(27)(175) := previousCrc(15); xorBitMap(27)(179) := previousCrc(19); xorBitMap(27)(187) := previousCrc(27); xorBitMap(27)(188) := previousCrc(28); xorBitMap(27)(189) := previousCrc(29); xorBitMap(27)(191) := previousCrc(31); 
      xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(164) := previousCrc(4); xorBitMap(28)(170) := previousCrc(10); xorBitMap(28)(173) := previousCrc(13); xorBitMap(28)(174) := previousCrc(14); xorBitMap(28)(176) := previousCrc(16); xorBitMap(28)(180) := previousCrc(20); xorBitMap(28)(188) := previousCrc(28); xorBitMap(28)(189) := previousCrc(29); xorBitMap(28)(190) := previousCrc(30); 
      xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(165) := previousCrc(5); xorBitMap(29)(171) := previousCrc(11); xorBitMap(29)(174) := previousCrc(14); xorBitMap(29)(175) := previousCrc(15); xorBitMap(29)(177) := previousCrc(17); xorBitMap(29)(181) := previousCrc(21); xorBitMap(29)(189) := previousCrc(29); xorBitMap(29)(190) := previousCrc(30); xorBitMap(29)(191) := previousCrc(31); 
      xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(166) := previousCrc(6); xorBitMap(30)(172) := previousCrc(12); xorBitMap(30)(175) := previousCrc(15); xorBitMap(30)(176) := previousCrc(16); xorBitMap(30)(178) := previousCrc(18); xorBitMap(30)(182) := previousCrc(22); xorBitMap(30)(190) := previousCrc(30); xorBitMap(30)(191) := previousCrc(31); 
      xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(167) := previousCrc(7); xorBitMap(31)(173) := previousCrc(13); xorBitMap(31)(176) := previousCrc(16); xorBitMap(31)(177) := previousCrc(17); xorBitMap(31)(179) := previousCrc(19); xorBitMap(31)(183) := previousCrc(23); xorBitMap(31)(191) := previousCrc(31); 
   end procedure;

   procedure xorBitMap4Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(31 downto 0)) is 
   begin
      xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(160) := previousCrc(0); xorBitMap(0)(166) := previousCrc(6); xorBitMap(0)(169) := previousCrc(9); xorBitMap(0)(170) := previousCrc(10); xorBitMap(0)(172) := previousCrc(12); xorBitMap(0)(176) := previousCrc(16); xorBitMap(0)(184) := previousCrc(24); xorBitMap(0)(185) := previousCrc(25); xorBitMap(0)(186) := previousCrc(26); xorBitMap(0)(188) := previousCrc(28); xorBitMap(0)(189) := previousCrc(29); xorBitMap(0)(190) := previousCrc(30); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(160) := previousCrc(0); xorBitMap(1)(161) := previousCrc(1); xorBitMap(1)(166) := previousCrc(6); xorBitMap(1)(167) := previousCrc(7); xorBitMap(1)(169) := previousCrc(9); xorBitMap(1)(171) := previousCrc(11); xorBitMap(1)(172) := previousCrc(12); xorBitMap(1)(173) := previousCrc(13); xorBitMap(1)(176) := previousCrc(16); xorBitMap(1)(177) := previousCrc(17); xorBitMap(1)(184) := previousCrc(24); xorBitMap(1)(187) := previousCrc(27); xorBitMap(1)(188) := previousCrc(28); 
      xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(160) := previousCrc(0); xorBitMap(2)(161) := previousCrc(1); xorBitMap(2)(162) := previousCrc(2); xorBitMap(2)(166) := previousCrc(6); xorBitMap(2)(167) := previousCrc(7); xorBitMap(2)(168) := previousCrc(8); xorBitMap(2)(169) := previousCrc(9); xorBitMap(2)(173) := previousCrc(13); xorBitMap(2)(174) := previousCrc(14); xorBitMap(2)(176) := previousCrc(16); xorBitMap(2)(177) := previousCrc(17); xorBitMap(2)(178) := previousCrc(18); xorBitMap(2)(184) := previousCrc(24); xorBitMap(2)(186) := previousCrc(26); xorBitMap(2)(190) := previousCrc(30); xorBitMap(2)(191) := previousCrc(31); 
      xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(161) := previousCrc(1); xorBitMap(3)(162) := previousCrc(2); xorBitMap(3)(163) := previousCrc(3); xorBitMap(3)(167) := previousCrc(7); xorBitMap(3)(168) := previousCrc(8); xorBitMap(3)(169) := previousCrc(9); xorBitMap(3)(170) := previousCrc(10); xorBitMap(3)(174) := previousCrc(14); xorBitMap(3)(175) := previousCrc(15); xorBitMap(3)(177) := previousCrc(17); xorBitMap(3)(178) := previousCrc(18); xorBitMap(3)(179) := previousCrc(19); xorBitMap(3)(185) := previousCrc(25); xorBitMap(3)(187) := previousCrc(27); xorBitMap(3)(191) := previousCrc(31); 
      xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(160) := previousCrc(0); xorBitMap(4)(162) := previousCrc(2); xorBitMap(4)(163) := previousCrc(3); xorBitMap(4)(164) := previousCrc(4); xorBitMap(4)(166) := previousCrc(6); xorBitMap(4)(168) := previousCrc(8); xorBitMap(4)(171) := previousCrc(11); xorBitMap(4)(172) := previousCrc(12); xorBitMap(4)(175) := previousCrc(15); xorBitMap(4)(178) := previousCrc(18); xorBitMap(4)(179) := previousCrc(19); xorBitMap(4)(180) := previousCrc(20); xorBitMap(4)(184) := previousCrc(24); xorBitMap(4)(185) := previousCrc(25); xorBitMap(4)(189) := previousCrc(29); xorBitMap(4)(190) := previousCrc(30); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(160) := previousCrc(0); xorBitMap(5)(161) := previousCrc(1); xorBitMap(5)(163) := previousCrc(3); xorBitMap(5)(164) := previousCrc(4); xorBitMap(5)(165) := previousCrc(5); xorBitMap(5)(166) := previousCrc(6); xorBitMap(5)(167) := previousCrc(7); xorBitMap(5)(170) := previousCrc(10); xorBitMap(5)(173) := previousCrc(13); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(180) := previousCrc(20); xorBitMap(5)(181) := previousCrc(21); xorBitMap(5)(184) := previousCrc(24); xorBitMap(5)(188) := previousCrc(28); xorBitMap(5)(189) := previousCrc(29); 
      xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(161) := previousCrc(1); xorBitMap(6)(162) := previousCrc(2); xorBitMap(6)(164) := previousCrc(4); xorBitMap(6)(165) := previousCrc(5); xorBitMap(6)(166) := previousCrc(6); xorBitMap(6)(167) := previousCrc(7); xorBitMap(6)(168) := previousCrc(8); xorBitMap(6)(171) := previousCrc(11); xorBitMap(6)(174) := previousCrc(14); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(181) := previousCrc(21); xorBitMap(6)(182) := previousCrc(22); xorBitMap(6)(185) := previousCrc(25); xorBitMap(6)(189) := previousCrc(29); xorBitMap(6)(190) := previousCrc(30); 
      xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(160) := previousCrc(0); xorBitMap(7)(162) := previousCrc(2); xorBitMap(7)(163) := previousCrc(3); xorBitMap(7)(165) := previousCrc(5); xorBitMap(7)(167) := previousCrc(7); xorBitMap(7)(168) := previousCrc(8); xorBitMap(7)(170) := previousCrc(10); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(176) := previousCrc(16); xorBitMap(7)(181) := previousCrc(21); xorBitMap(7)(182) := previousCrc(22); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(184) := previousCrc(24); xorBitMap(7)(185) := previousCrc(25); xorBitMap(7)(188) := previousCrc(28); xorBitMap(7)(189) := previousCrc(29); 
      xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(160) := previousCrc(0); xorBitMap(8)(161) := previousCrc(1); xorBitMap(8)(163) := previousCrc(3); xorBitMap(8)(164) := previousCrc(4); xorBitMap(8)(168) := previousCrc(8); xorBitMap(8)(170) := previousCrc(10); xorBitMap(8)(171) := previousCrc(11); xorBitMap(8)(172) := previousCrc(12); xorBitMap(8)(177) := previousCrc(17); xorBitMap(8)(182) := previousCrc(22); xorBitMap(8)(183) := previousCrc(23); xorBitMap(8)(188) := previousCrc(28); xorBitMap(8)(191) := previousCrc(31); 
      xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(161) := previousCrc(1); xorBitMap(9)(162) := previousCrc(2); xorBitMap(9)(164) := previousCrc(4); xorBitMap(9)(165) := previousCrc(5); xorBitMap(9)(169) := previousCrc(9); xorBitMap(9)(171) := previousCrc(11); xorBitMap(9)(172) := previousCrc(12); xorBitMap(9)(173) := previousCrc(13); xorBitMap(9)(178) := previousCrc(18); xorBitMap(9)(183) := previousCrc(23); xorBitMap(9)(184) := previousCrc(24); xorBitMap(9)(189) := previousCrc(29); 
      xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(160) := previousCrc(0); xorBitMap(10)(162) := previousCrc(2); xorBitMap(10)(163) := previousCrc(3); xorBitMap(10)(165) := previousCrc(5); xorBitMap(10)(169) := previousCrc(9); xorBitMap(10)(173) := previousCrc(13); xorBitMap(10)(174) := previousCrc(14); xorBitMap(10)(176) := previousCrc(16); xorBitMap(10)(179) := previousCrc(19); xorBitMap(10)(186) := previousCrc(26); xorBitMap(10)(188) := previousCrc(28); xorBitMap(10)(189) := previousCrc(29); xorBitMap(10)(191) := previousCrc(31); 
      xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(160) := previousCrc(0); xorBitMap(11)(161) := previousCrc(1); xorBitMap(11)(163) := previousCrc(3); xorBitMap(11)(164) := previousCrc(4); xorBitMap(11)(169) := previousCrc(9); xorBitMap(11)(172) := previousCrc(12); xorBitMap(11)(174) := previousCrc(14); xorBitMap(11)(175) := previousCrc(15); xorBitMap(11)(176) := previousCrc(16); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(180) := previousCrc(20); xorBitMap(11)(184) := previousCrc(24); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(186) := previousCrc(26); xorBitMap(11)(187) := previousCrc(27); xorBitMap(11)(188) := previousCrc(28); xorBitMap(11)(191) := previousCrc(31); 
      xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(160) := previousCrc(0); xorBitMap(12)(161) := previousCrc(1); xorBitMap(12)(162) := previousCrc(2); xorBitMap(12)(164) := previousCrc(4); xorBitMap(12)(165) := previousCrc(5); xorBitMap(12)(166) := previousCrc(6); xorBitMap(12)(169) := previousCrc(9); xorBitMap(12)(172) := previousCrc(12); xorBitMap(12)(173) := previousCrc(13); xorBitMap(12)(175) := previousCrc(15); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(178) := previousCrc(18); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(184) := previousCrc(24); xorBitMap(12)(187) := previousCrc(27); xorBitMap(12)(190) := previousCrc(30); xorBitMap(12)(191) := previousCrc(31); 
      xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(161) := previousCrc(1); xorBitMap(13)(162) := previousCrc(2); xorBitMap(13)(163) := previousCrc(3); xorBitMap(13)(165) := previousCrc(5); xorBitMap(13)(166) := previousCrc(6); xorBitMap(13)(167) := previousCrc(7); xorBitMap(13)(170) := previousCrc(10); xorBitMap(13)(173) := previousCrc(13); xorBitMap(13)(174) := previousCrc(14); xorBitMap(13)(176) := previousCrc(16); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(179) := previousCrc(19); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(185) := previousCrc(25); xorBitMap(13)(188) := previousCrc(28); xorBitMap(13)(191) := previousCrc(31); 
      xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(162) := previousCrc(2); xorBitMap(14)(163) := previousCrc(3); xorBitMap(14)(164) := previousCrc(4); xorBitMap(14)(166) := previousCrc(6); xorBitMap(14)(167) := previousCrc(7); xorBitMap(14)(168) := previousCrc(8); xorBitMap(14)(171) := previousCrc(11); xorBitMap(14)(174) := previousCrc(14); xorBitMap(14)(175) := previousCrc(15); xorBitMap(14)(177) := previousCrc(17); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(180) := previousCrc(20); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(186) := previousCrc(26); xorBitMap(14)(189) := previousCrc(29); 
      xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(163) := previousCrc(3); xorBitMap(15)(164) := previousCrc(4); xorBitMap(15)(165) := previousCrc(5); xorBitMap(15)(167) := previousCrc(7); xorBitMap(15)(168) := previousCrc(8); xorBitMap(15)(169) := previousCrc(9); xorBitMap(15)(172) := previousCrc(12); xorBitMap(15)(175) := previousCrc(15); xorBitMap(15)(176) := previousCrc(16); xorBitMap(15)(178) := previousCrc(18); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(181) := previousCrc(21); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(187) := previousCrc(27); xorBitMap(15)(190) := previousCrc(30); 
      xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(160) := previousCrc(0); xorBitMap(16)(164) := previousCrc(4); xorBitMap(16)(165) := previousCrc(5); xorBitMap(16)(168) := previousCrc(8); xorBitMap(16)(172) := previousCrc(12); xorBitMap(16)(173) := previousCrc(13); xorBitMap(16)(177) := previousCrc(17); xorBitMap(16)(179) := previousCrc(19); xorBitMap(16)(181) := previousCrc(21); xorBitMap(16)(182) := previousCrc(22); xorBitMap(16)(184) := previousCrc(24); xorBitMap(16)(186) := previousCrc(26); xorBitMap(16)(189) := previousCrc(29); xorBitMap(16)(190) := previousCrc(30); 
      xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(161) := previousCrc(1); xorBitMap(17)(165) := previousCrc(5); xorBitMap(17)(166) := previousCrc(6); xorBitMap(17)(169) := previousCrc(9); xorBitMap(17)(173) := previousCrc(13); xorBitMap(17)(174) := previousCrc(14); xorBitMap(17)(178) := previousCrc(18); xorBitMap(17)(180) := previousCrc(20); xorBitMap(17)(182) := previousCrc(22); xorBitMap(17)(183) := previousCrc(23); xorBitMap(17)(185) := previousCrc(25); xorBitMap(17)(187) := previousCrc(27); xorBitMap(17)(190) := previousCrc(30); xorBitMap(17)(191) := previousCrc(31); 
      xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(162) := previousCrc(2); xorBitMap(18)(166) := previousCrc(6); xorBitMap(18)(167) := previousCrc(7); xorBitMap(18)(170) := previousCrc(10); xorBitMap(18)(174) := previousCrc(14); xorBitMap(18)(175) := previousCrc(15); xorBitMap(18)(179) := previousCrc(19); xorBitMap(18)(181) := previousCrc(21); xorBitMap(18)(183) := previousCrc(23); xorBitMap(18)(184) := previousCrc(24); xorBitMap(18)(186) := previousCrc(26); xorBitMap(18)(188) := previousCrc(28); xorBitMap(18)(191) := previousCrc(31); 
      xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(163) := previousCrc(3); xorBitMap(19)(167) := previousCrc(7); xorBitMap(19)(168) := previousCrc(8); xorBitMap(19)(171) := previousCrc(11); xorBitMap(19)(175) := previousCrc(15); xorBitMap(19)(176) := previousCrc(16); xorBitMap(19)(180) := previousCrc(20); xorBitMap(19)(182) := previousCrc(22); xorBitMap(19)(184) := previousCrc(24); xorBitMap(19)(185) := previousCrc(25); xorBitMap(19)(187) := previousCrc(27); xorBitMap(19)(189) := previousCrc(29); 
      xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(164) := previousCrc(4); xorBitMap(20)(168) := previousCrc(8); xorBitMap(20)(169) := previousCrc(9); xorBitMap(20)(172) := previousCrc(12); xorBitMap(20)(176) := previousCrc(16); xorBitMap(20)(177) := previousCrc(17); xorBitMap(20)(181) := previousCrc(21); xorBitMap(20)(183) := previousCrc(23); xorBitMap(20)(185) := previousCrc(25); xorBitMap(20)(186) := previousCrc(26); xorBitMap(20)(188) := previousCrc(28); xorBitMap(20)(190) := previousCrc(30); 
      xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(165) := previousCrc(5); xorBitMap(21)(169) := previousCrc(9); xorBitMap(21)(170) := previousCrc(10); xorBitMap(21)(173) := previousCrc(13); xorBitMap(21)(177) := previousCrc(17); xorBitMap(21)(178) := previousCrc(18); xorBitMap(21)(182) := previousCrc(22); xorBitMap(21)(184) := previousCrc(24); xorBitMap(21)(186) := previousCrc(26); xorBitMap(21)(187) := previousCrc(27); xorBitMap(21)(189) := previousCrc(29); xorBitMap(21)(191) := previousCrc(31); 
      xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(160) := previousCrc(0); xorBitMap(22)(169) := previousCrc(9); xorBitMap(22)(171) := previousCrc(11); xorBitMap(22)(172) := previousCrc(12); xorBitMap(22)(174) := previousCrc(14); xorBitMap(22)(176) := previousCrc(16); xorBitMap(22)(178) := previousCrc(18); xorBitMap(22)(179) := previousCrc(19); xorBitMap(22)(183) := previousCrc(23); xorBitMap(22)(184) := previousCrc(24); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(187) := previousCrc(27); xorBitMap(22)(189) := previousCrc(29); xorBitMap(22)(191) := previousCrc(31); 
      xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(160) := previousCrc(0); xorBitMap(23)(161) := previousCrc(1); xorBitMap(23)(166) := previousCrc(6); xorBitMap(23)(169) := previousCrc(9); xorBitMap(23)(173) := previousCrc(13); xorBitMap(23)(175) := previousCrc(15); xorBitMap(23)(176) := previousCrc(16); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(179) := previousCrc(19); xorBitMap(23)(180) := previousCrc(20); xorBitMap(23)(186) := previousCrc(26); xorBitMap(23)(187) := previousCrc(27); xorBitMap(23)(189) := previousCrc(29); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(161) := previousCrc(1); xorBitMap(24)(162) := previousCrc(2); xorBitMap(24)(167) := previousCrc(7); xorBitMap(24)(170) := previousCrc(10); xorBitMap(24)(174) := previousCrc(14); xorBitMap(24)(176) := previousCrc(16); xorBitMap(24)(177) := previousCrc(17); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(180) := previousCrc(20); xorBitMap(24)(181) := previousCrc(21); xorBitMap(24)(187) := previousCrc(27); xorBitMap(24)(188) := previousCrc(28); xorBitMap(24)(190) := previousCrc(30); 
      xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(162) := previousCrc(2); xorBitMap(25)(163) := previousCrc(3); xorBitMap(25)(168) := previousCrc(8); xorBitMap(25)(171) := previousCrc(11); xorBitMap(25)(175) := previousCrc(15); xorBitMap(25)(177) := previousCrc(17); xorBitMap(25)(178) := previousCrc(18); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(181) := previousCrc(21); xorBitMap(25)(182) := previousCrc(22); xorBitMap(25)(188) := previousCrc(28); xorBitMap(25)(189) := previousCrc(29); xorBitMap(25)(191) := previousCrc(31); 
      xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(160) := previousCrc(0); xorBitMap(26)(163) := previousCrc(3); xorBitMap(26)(164) := previousCrc(4); xorBitMap(26)(166) := previousCrc(6); xorBitMap(26)(170) := previousCrc(10); xorBitMap(26)(178) := previousCrc(18); xorBitMap(26)(179) := previousCrc(19); xorBitMap(26)(180) := previousCrc(20); xorBitMap(26)(182) := previousCrc(22); xorBitMap(26)(183) := previousCrc(23); xorBitMap(26)(184) := previousCrc(24); xorBitMap(26)(185) := previousCrc(25); xorBitMap(26)(186) := previousCrc(26); xorBitMap(26)(188) := previousCrc(28); xorBitMap(26)(191) := previousCrc(31); 
      xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(161) := previousCrc(1); xorBitMap(27)(164) := previousCrc(4); xorBitMap(27)(165) := previousCrc(5); xorBitMap(27)(167) := previousCrc(7); xorBitMap(27)(171) := previousCrc(11); xorBitMap(27)(179) := previousCrc(19); xorBitMap(27)(180) := previousCrc(20); xorBitMap(27)(181) := previousCrc(21); xorBitMap(27)(183) := previousCrc(23); xorBitMap(27)(184) := previousCrc(24); xorBitMap(27)(185) := previousCrc(25); xorBitMap(27)(186) := previousCrc(26); xorBitMap(27)(187) := previousCrc(27); xorBitMap(27)(189) := previousCrc(29); 
      xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(162) := previousCrc(2); xorBitMap(28)(165) := previousCrc(5); xorBitMap(28)(166) := previousCrc(6); xorBitMap(28)(168) := previousCrc(8); xorBitMap(28)(172) := previousCrc(12); xorBitMap(28)(180) := previousCrc(20); xorBitMap(28)(181) := previousCrc(21); xorBitMap(28)(182) := previousCrc(22); xorBitMap(28)(184) := previousCrc(24); xorBitMap(28)(185) := previousCrc(25); xorBitMap(28)(186) := previousCrc(26); xorBitMap(28)(187) := previousCrc(27); xorBitMap(28)(188) := previousCrc(28); xorBitMap(28)(190) := previousCrc(30); 
      xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(163) := previousCrc(3); xorBitMap(29)(166) := previousCrc(6); xorBitMap(29)(167) := previousCrc(7); xorBitMap(29)(169) := previousCrc(9); xorBitMap(29)(173) := previousCrc(13); xorBitMap(29)(181) := previousCrc(21); xorBitMap(29)(182) := previousCrc(22); xorBitMap(29)(183) := previousCrc(23); xorBitMap(29)(185) := previousCrc(25); xorBitMap(29)(186) := previousCrc(26); xorBitMap(29)(187) := previousCrc(27); xorBitMap(29)(188) := previousCrc(28); xorBitMap(29)(189) := previousCrc(29); xorBitMap(29)(191) := previousCrc(31); 
      xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(164) := previousCrc(4); xorBitMap(30)(167) := previousCrc(7); xorBitMap(30)(168) := previousCrc(8); xorBitMap(30)(170) := previousCrc(10); xorBitMap(30)(174) := previousCrc(14); xorBitMap(30)(182) := previousCrc(22); xorBitMap(30)(183) := previousCrc(23); xorBitMap(30)(184) := previousCrc(24); xorBitMap(30)(186) := previousCrc(26); xorBitMap(30)(187) := previousCrc(27); xorBitMap(30)(188) := previousCrc(28); xorBitMap(30)(189) := previousCrc(29); xorBitMap(30)(190) := previousCrc(30); 
      xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(165) := previousCrc(5); xorBitMap(31)(168) := previousCrc(8); xorBitMap(31)(169) := previousCrc(9); xorBitMap(31)(171) := previousCrc(11); xorBitMap(31)(175) := previousCrc(15); xorBitMap(31)(183) := previousCrc(23); xorBitMap(31)(184) := previousCrc(24); xorBitMap(31)(185) := previousCrc(25); xorBitMap(31)(187) := previousCrc(27); xorBitMap(31)(188) := previousCrc(28); xorBitMap(31)(189) := previousCrc(29); xorBitMap(31)(190) := previousCrc(30); xorBitMap(31)(191) := previousCrc(31); 
   end procedure;

   procedure xorBitMap5Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(39 downto 0)) is 
   begin
      xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(161) := previousCrc(1); xorBitMap(0)(162) := previousCrc(2); xorBitMap(0)(164) := previousCrc(4); xorBitMap(0)(168) := previousCrc(8); xorBitMap(0)(176) := previousCrc(16); xorBitMap(0)(177) := previousCrc(17); xorBitMap(0)(178) := previousCrc(18); xorBitMap(0)(180) := previousCrc(20); xorBitMap(0)(181) := previousCrc(21); xorBitMap(0)(182) := previousCrc(22); xorBitMap(0)(183) := previousCrc(23); xorBitMap(0)(184) := previousCrc(24); xorBitMap(0)(186) := previousCrc(26); xorBitMap(0)(189) := previousCrc(29); 
      xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(161) := previousCrc(1); xorBitMap(1)(163) := previousCrc(3); xorBitMap(1)(164) := previousCrc(4); xorBitMap(1)(165) := previousCrc(5); xorBitMap(1)(168) := previousCrc(8); xorBitMap(1)(169) := previousCrc(9); xorBitMap(1)(176) := previousCrc(16); xorBitMap(1)(179) := previousCrc(19); xorBitMap(1)(180) := previousCrc(20); xorBitMap(1)(185) := previousCrc(25); xorBitMap(1)(186) := previousCrc(26); xorBitMap(1)(187) := previousCrc(27); xorBitMap(1)(189) := previousCrc(29); xorBitMap(1)(190) := previousCrc(30); 
      xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(160) := previousCrc(0); xorBitMap(2)(161) := previousCrc(1); xorBitMap(2)(165) := previousCrc(5); xorBitMap(2)(166) := previousCrc(6); xorBitMap(2)(168) := previousCrc(8); xorBitMap(2)(169) := previousCrc(9); xorBitMap(2)(170) := previousCrc(10); xorBitMap(2)(176) := previousCrc(16); xorBitMap(2)(178) := previousCrc(18); xorBitMap(2)(182) := previousCrc(22); xorBitMap(2)(183) := previousCrc(23); xorBitMap(2)(184) := previousCrc(24); xorBitMap(2)(187) := previousCrc(27); xorBitMap(2)(188) := previousCrc(28); xorBitMap(2)(189) := previousCrc(29); xorBitMap(2)(190) := previousCrc(30); xorBitMap(2)(191) := previousCrc(31); 
      xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(160) := previousCrc(0); xorBitMap(3)(161) := previousCrc(1); xorBitMap(3)(162) := previousCrc(2); xorBitMap(3)(166) := previousCrc(6); xorBitMap(3)(167) := previousCrc(7); xorBitMap(3)(169) := previousCrc(9); xorBitMap(3)(170) := previousCrc(10); xorBitMap(3)(171) := previousCrc(11); xorBitMap(3)(177) := previousCrc(17); xorBitMap(3)(179) := previousCrc(19); xorBitMap(3)(183) := previousCrc(23); xorBitMap(3)(184) := previousCrc(24); xorBitMap(3)(185) := previousCrc(25); xorBitMap(3)(188) := previousCrc(28); xorBitMap(3)(189) := previousCrc(29); xorBitMap(3)(190) := previousCrc(30); xorBitMap(3)(191) := previousCrc(31); 
      xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(160) := previousCrc(0); xorBitMap(4)(163) := previousCrc(3); xorBitMap(4)(164) := previousCrc(4); xorBitMap(4)(167) := previousCrc(7); xorBitMap(4)(170) := previousCrc(10); xorBitMap(4)(171) := previousCrc(11); xorBitMap(4)(172) := previousCrc(12); xorBitMap(4)(176) := previousCrc(16); xorBitMap(4)(177) := previousCrc(17); xorBitMap(4)(181) := previousCrc(21); xorBitMap(4)(182) := previousCrc(22); xorBitMap(4)(183) := previousCrc(23); xorBitMap(4)(185) := previousCrc(25); xorBitMap(4)(190) := previousCrc(30); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(162) := previousCrc(2); xorBitMap(5)(165) := previousCrc(5); xorBitMap(5)(171) := previousCrc(11); xorBitMap(5)(172) := previousCrc(12); xorBitMap(5)(173) := previousCrc(13); xorBitMap(5)(176) := previousCrc(16); xorBitMap(5)(180) := previousCrc(20); xorBitMap(5)(181) := previousCrc(21); xorBitMap(5)(189) := previousCrc(29); xorBitMap(5)(191) := previousCrc(31); 
      xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(160) := previousCrc(0); xorBitMap(6)(163) := previousCrc(3); xorBitMap(6)(166) := previousCrc(6); xorBitMap(6)(172) := previousCrc(12); xorBitMap(6)(173) := previousCrc(13); xorBitMap(6)(174) := previousCrc(14); xorBitMap(6)(177) := previousCrc(17); xorBitMap(6)(181) := previousCrc(21); xorBitMap(6)(182) := previousCrc(22); xorBitMap(6)(190) := previousCrc(30); 
      xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(160) := previousCrc(0); xorBitMap(7)(162) := previousCrc(2); xorBitMap(7)(167) := previousCrc(7); xorBitMap(7)(168) := previousCrc(8); xorBitMap(7)(173) := previousCrc(13); xorBitMap(7)(174) := previousCrc(14); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(176) := previousCrc(16); xorBitMap(7)(177) := previousCrc(17); xorBitMap(7)(180) := previousCrc(20); xorBitMap(7)(181) := previousCrc(21); xorBitMap(7)(184) := previousCrc(24); xorBitMap(7)(186) := previousCrc(26); xorBitMap(7)(189) := previousCrc(29); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(160) := previousCrc(0); xorBitMap(8)(162) := previousCrc(2); xorBitMap(8)(163) := previousCrc(3); xorBitMap(8)(164) := previousCrc(4); xorBitMap(8)(169) := previousCrc(9); xorBitMap(8)(174) := previousCrc(14); xorBitMap(8)(175) := previousCrc(15); xorBitMap(8)(180) := previousCrc(20); xorBitMap(8)(183) := previousCrc(23); xorBitMap(8)(184) := previousCrc(24); xorBitMap(8)(185) := previousCrc(25); xorBitMap(8)(186) := previousCrc(26); xorBitMap(8)(187) := previousCrc(27); xorBitMap(8)(189) := previousCrc(29); xorBitMap(8)(190) := previousCrc(30); 
      xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(161) := previousCrc(1); xorBitMap(9)(163) := previousCrc(3); xorBitMap(9)(164) := previousCrc(4); xorBitMap(9)(165) := previousCrc(5); xorBitMap(9)(170) := previousCrc(10); xorBitMap(9)(175) := previousCrc(15); xorBitMap(9)(176) := previousCrc(16); xorBitMap(9)(181) := previousCrc(21); xorBitMap(9)(184) := previousCrc(24); xorBitMap(9)(185) := previousCrc(25); xorBitMap(9)(186) := previousCrc(26); xorBitMap(9)(187) := previousCrc(27); xorBitMap(9)(188) := previousCrc(28); xorBitMap(9)(190) := previousCrc(30); xorBitMap(9)(191) := previousCrc(31); 
      xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(161) := previousCrc(1); xorBitMap(10)(165) := previousCrc(5); xorBitMap(10)(166) := previousCrc(6); xorBitMap(10)(168) := previousCrc(8); xorBitMap(10)(171) := previousCrc(11); xorBitMap(10)(178) := previousCrc(18); xorBitMap(10)(180) := previousCrc(20); xorBitMap(10)(181) := previousCrc(21); xorBitMap(10)(183) := previousCrc(23); xorBitMap(10)(184) := previousCrc(24); xorBitMap(10)(185) := previousCrc(25); xorBitMap(10)(187) := previousCrc(27); xorBitMap(10)(188) := previousCrc(28); xorBitMap(10)(191) := previousCrc(31); 
      xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(161) := previousCrc(1); xorBitMap(11)(164) := previousCrc(4); xorBitMap(11)(166) := previousCrc(6); xorBitMap(11)(167) := previousCrc(7); xorBitMap(11)(168) := previousCrc(8); xorBitMap(11)(169) := previousCrc(9); xorBitMap(11)(172) := previousCrc(12); xorBitMap(11)(176) := previousCrc(16); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(178) := previousCrc(18); xorBitMap(11)(179) := previousCrc(19); xorBitMap(11)(180) := previousCrc(20); xorBitMap(11)(183) := previousCrc(23); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(188) := previousCrc(28); 
      xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(161) := previousCrc(1); xorBitMap(12)(164) := previousCrc(4); xorBitMap(12)(165) := previousCrc(5); xorBitMap(12)(167) := previousCrc(7); xorBitMap(12)(169) := previousCrc(9); xorBitMap(12)(170) := previousCrc(10); xorBitMap(12)(173) := previousCrc(13); xorBitMap(12)(176) := previousCrc(16); xorBitMap(12)(179) := previousCrc(19); xorBitMap(12)(182) := previousCrc(22); xorBitMap(12)(183) := previousCrc(23); 
      xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(162) := previousCrc(2); xorBitMap(13)(165) := previousCrc(5); xorBitMap(13)(166) := previousCrc(6); xorBitMap(13)(168) := previousCrc(8); xorBitMap(13)(170) := previousCrc(10); xorBitMap(13)(171) := previousCrc(11); xorBitMap(13)(174) := previousCrc(14); xorBitMap(13)(177) := previousCrc(17); xorBitMap(13)(180) := previousCrc(20); xorBitMap(13)(183) := previousCrc(23); xorBitMap(13)(184) := previousCrc(24); 
      xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(160) := previousCrc(0); xorBitMap(14)(163) := previousCrc(3); xorBitMap(14)(166) := previousCrc(6); xorBitMap(14)(167) := previousCrc(7); xorBitMap(14)(169) := previousCrc(9); xorBitMap(14)(171) := previousCrc(11); xorBitMap(14)(172) := previousCrc(12); xorBitMap(14)(175) := previousCrc(15); xorBitMap(14)(178) := previousCrc(18); xorBitMap(14)(181) := previousCrc(21); xorBitMap(14)(184) := previousCrc(24); xorBitMap(14)(185) := previousCrc(25); 
      xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(160) := previousCrc(0); xorBitMap(15)(161) := previousCrc(1); xorBitMap(15)(164) := previousCrc(4); xorBitMap(15)(167) := previousCrc(7); xorBitMap(15)(168) := previousCrc(8); xorBitMap(15)(170) := previousCrc(10); xorBitMap(15)(172) := previousCrc(12); xorBitMap(15)(173) := previousCrc(13); xorBitMap(15)(176) := previousCrc(16); xorBitMap(15)(179) := previousCrc(19); xorBitMap(15)(182) := previousCrc(22); xorBitMap(15)(185) := previousCrc(25); xorBitMap(15)(186) := previousCrc(26); 
      xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(160) := previousCrc(0); xorBitMap(16)(164) := previousCrc(4); xorBitMap(16)(165) := previousCrc(5); xorBitMap(16)(169) := previousCrc(9); xorBitMap(16)(171) := previousCrc(11); xorBitMap(16)(173) := previousCrc(13); xorBitMap(16)(174) := previousCrc(14); xorBitMap(16)(176) := previousCrc(16); xorBitMap(16)(178) := previousCrc(18); xorBitMap(16)(181) := previousCrc(21); xorBitMap(16)(182) := previousCrc(22); xorBitMap(16)(184) := previousCrc(24); xorBitMap(16)(187) := previousCrc(27); xorBitMap(16)(189) := previousCrc(29); 
      xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(161) := previousCrc(1); xorBitMap(17)(165) := previousCrc(5); xorBitMap(17)(166) := previousCrc(6); xorBitMap(17)(170) := previousCrc(10); xorBitMap(17)(172) := previousCrc(12); xorBitMap(17)(174) := previousCrc(14); xorBitMap(17)(175) := previousCrc(15); xorBitMap(17)(177) := previousCrc(17); xorBitMap(17)(179) := previousCrc(19); xorBitMap(17)(182) := previousCrc(22); xorBitMap(17)(183) := previousCrc(23); xorBitMap(17)(185) := previousCrc(25); xorBitMap(17)(188) := previousCrc(28); xorBitMap(17)(190) := previousCrc(30); 
      xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(162) := previousCrc(2); xorBitMap(18)(166) := previousCrc(6); xorBitMap(18)(167) := previousCrc(7); xorBitMap(18)(171) := previousCrc(11); xorBitMap(18)(173) := previousCrc(13); xorBitMap(18)(175) := previousCrc(15); xorBitMap(18)(176) := previousCrc(16); xorBitMap(18)(178) := previousCrc(18); xorBitMap(18)(180) := previousCrc(20); xorBitMap(18)(183) := previousCrc(23); xorBitMap(18)(184) := previousCrc(24); xorBitMap(18)(186) := previousCrc(26); xorBitMap(18)(189) := previousCrc(29); xorBitMap(18)(191) := previousCrc(31); 
      xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(160) := previousCrc(0); xorBitMap(19)(163) := previousCrc(3); xorBitMap(19)(167) := previousCrc(7); xorBitMap(19)(168) := previousCrc(8); xorBitMap(19)(172) := previousCrc(12); xorBitMap(19)(174) := previousCrc(14); xorBitMap(19)(176) := previousCrc(16); xorBitMap(19)(177) := previousCrc(17); xorBitMap(19)(179) := previousCrc(19); xorBitMap(19)(181) := previousCrc(21); xorBitMap(19)(184) := previousCrc(24); xorBitMap(19)(185) := previousCrc(25); xorBitMap(19)(187) := previousCrc(27); xorBitMap(19)(190) := previousCrc(30); 
      xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(160) := previousCrc(0); xorBitMap(20)(161) := previousCrc(1); xorBitMap(20)(164) := previousCrc(4); xorBitMap(20)(168) := previousCrc(8); xorBitMap(20)(169) := previousCrc(9); xorBitMap(20)(173) := previousCrc(13); xorBitMap(20)(175) := previousCrc(15); xorBitMap(20)(177) := previousCrc(17); xorBitMap(20)(178) := previousCrc(18); xorBitMap(20)(180) := previousCrc(20); xorBitMap(20)(182) := previousCrc(22); xorBitMap(20)(185) := previousCrc(25); xorBitMap(20)(186) := previousCrc(26); xorBitMap(20)(188) := previousCrc(28); xorBitMap(20)(191) := previousCrc(31); 
      xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(161) := previousCrc(1); xorBitMap(21)(162) := previousCrc(2); xorBitMap(21)(165) := previousCrc(5); xorBitMap(21)(169) := previousCrc(9); xorBitMap(21)(170) := previousCrc(10); xorBitMap(21)(174) := previousCrc(14); xorBitMap(21)(176) := previousCrc(16); xorBitMap(21)(178) := previousCrc(18); xorBitMap(21)(179) := previousCrc(19); xorBitMap(21)(181) := previousCrc(21); xorBitMap(21)(183) := previousCrc(23); xorBitMap(21)(186) := previousCrc(26); xorBitMap(21)(187) := previousCrc(27); xorBitMap(21)(189) := previousCrc(29); 
      xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(161) := previousCrc(1); xorBitMap(22)(163) := previousCrc(3); xorBitMap(22)(164) := previousCrc(4); xorBitMap(22)(166) := previousCrc(6); xorBitMap(22)(168) := previousCrc(8); xorBitMap(22)(170) := previousCrc(10); xorBitMap(22)(171) := previousCrc(11); xorBitMap(22)(175) := previousCrc(15); xorBitMap(22)(176) := previousCrc(16); xorBitMap(22)(178) := previousCrc(18); xorBitMap(22)(179) := previousCrc(19); xorBitMap(22)(181) := previousCrc(21); xorBitMap(22)(183) := previousCrc(23); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(187) := previousCrc(27); xorBitMap(22)(188) := previousCrc(28); xorBitMap(22)(189) := previousCrc(29); xorBitMap(22)(190) := previousCrc(30); 
      xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(161) := previousCrc(1); xorBitMap(23)(165) := previousCrc(5); xorBitMap(23)(167) := previousCrc(7); xorBitMap(23)(168) := previousCrc(8); xorBitMap(23)(169) := previousCrc(9); xorBitMap(23)(171) := previousCrc(11); xorBitMap(23)(172) := previousCrc(12); xorBitMap(23)(178) := previousCrc(18); xorBitMap(23)(179) := previousCrc(19); xorBitMap(23)(181) := previousCrc(21); xorBitMap(23)(183) := previousCrc(23); xorBitMap(23)(186) := previousCrc(26); xorBitMap(23)(187) := previousCrc(27); xorBitMap(23)(188) := previousCrc(28); xorBitMap(23)(190) := previousCrc(30); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(162) := previousCrc(2); xorBitMap(24)(166) := previousCrc(6); xorBitMap(24)(168) := previousCrc(8); xorBitMap(24)(169) := previousCrc(9); xorBitMap(24)(170) := previousCrc(10); xorBitMap(24)(172) := previousCrc(12); xorBitMap(24)(173) := previousCrc(13); xorBitMap(24)(179) := previousCrc(19); xorBitMap(24)(180) := previousCrc(20); xorBitMap(24)(182) := previousCrc(22); xorBitMap(24)(184) := previousCrc(24); xorBitMap(24)(187) := previousCrc(27); xorBitMap(24)(188) := previousCrc(28); xorBitMap(24)(189) := previousCrc(29); xorBitMap(24)(191) := previousCrc(31); 
      xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(160) := previousCrc(0); xorBitMap(25)(163) := previousCrc(3); xorBitMap(25)(167) := previousCrc(7); xorBitMap(25)(169) := previousCrc(9); xorBitMap(25)(170) := previousCrc(10); xorBitMap(25)(171) := previousCrc(11); xorBitMap(25)(173) := previousCrc(13); xorBitMap(25)(174) := previousCrc(14); xorBitMap(25)(180) := previousCrc(20); xorBitMap(25)(181) := previousCrc(21); xorBitMap(25)(183) := previousCrc(23); xorBitMap(25)(185) := previousCrc(25); xorBitMap(25)(188) := previousCrc(28); xorBitMap(25)(189) := previousCrc(29); xorBitMap(25)(190) := previousCrc(30); 
      xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(162) := previousCrc(2); xorBitMap(26)(170) := previousCrc(10); xorBitMap(26)(171) := previousCrc(11); xorBitMap(26)(172) := previousCrc(12); xorBitMap(26)(174) := previousCrc(14); xorBitMap(26)(175) := previousCrc(15); xorBitMap(26)(176) := previousCrc(16); xorBitMap(26)(177) := previousCrc(17); xorBitMap(26)(178) := previousCrc(18); xorBitMap(26)(180) := previousCrc(20); xorBitMap(26)(183) := previousCrc(23); xorBitMap(26)(190) := previousCrc(30); xorBitMap(26)(191) := previousCrc(31); 
      xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(163) := previousCrc(3); xorBitMap(27)(171) := previousCrc(11); xorBitMap(27)(172) := previousCrc(12); xorBitMap(27)(173) := previousCrc(13); xorBitMap(27)(175) := previousCrc(15); xorBitMap(27)(176) := previousCrc(16); xorBitMap(27)(177) := previousCrc(17); xorBitMap(27)(178) := previousCrc(18); xorBitMap(27)(179) := previousCrc(19); xorBitMap(27)(181) := previousCrc(21); xorBitMap(27)(184) := previousCrc(24); xorBitMap(27)(191) := previousCrc(31); 
      xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(160) := previousCrc(0); xorBitMap(28)(164) := previousCrc(4); xorBitMap(28)(172) := previousCrc(12); xorBitMap(28)(173) := previousCrc(13); xorBitMap(28)(174) := previousCrc(14); xorBitMap(28)(176) := previousCrc(16); xorBitMap(28)(177) := previousCrc(17); xorBitMap(28)(178) := previousCrc(18); xorBitMap(28)(179) := previousCrc(19); xorBitMap(28)(180) := previousCrc(20); xorBitMap(28)(182) := previousCrc(22); xorBitMap(28)(185) := previousCrc(25); 
      xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(161) := previousCrc(1); xorBitMap(29)(165) := previousCrc(5); xorBitMap(29)(173) := previousCrc(13); xorBitMap(29)(174) := previousCrc(14); xorBitMap(29)(175) := previousCrc(15); xorBitMap(29)(177) := previousCrc(17); xorBitMap(29)(178) := previousCrc(18); xorBitMap(29)(179) := previousCrc(19); xorBitMap(29)(180) := previousCrc(20); xorBitMap(29)(181) := previousCrc(21); xorBitMap(29)(183) := previousCrc(23); xorBitMap(29)(186) := previousCrc(26); 
      xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(160) := previousCrc(0); xorBitMap(30)(162) := previousCrc(2); xorBitMap(30)(166) := previousCrc(6); xorBitMap(30)(174) := previousCrc(14); xorBitMap(30)(175) := previousCrc(15); xorBitMap(30)(176) := previousCrc(16); xorBitMap(30)(178) := previousCrc(18); xorBitMap(30)(179) := previousCrc(19); xorBitMap(30)(180) := previousCrc(20); xorBitMap(30)(181) := previousCrc(21); xorBitMap(30)(182) := previousCrc(22); xorBitMap(30)(184) := previousCrc(24); xorBitMap(30)(187) := previousCrc(27); 
      xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(160) := previousCrc(0); xorBitMap(31)(161) := previousCrc(1); xorBitMap(31)(163) := previousCrc(3); xorBitMap(31)(167) := previousCrc(7); xorBitMap(31)(175) := previousCrc(15); xorBitMap(31)(176) := previousCrc(16); xorBitMap(31)(177) := previousCrc(17); xorBitMap(31)(179) := previousCrc(19); xorBitMap(31)(180) := previousCrc(20); xorBitMap(31)(181) := previousCrc(21); xorBitMap(31)(182) := previousCrc(22); xorBitMap(31)(183) := previousCrc(23); xorBitMap(31)(185) := previousCrc(25); xorBitMap(31)(188) := previousCrc(28); 
   end procedure;

   procedure xorBitMap6Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(47 downto 0)) is 
   begin
      xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(160) := previousCrc(0); xorBitMap(0)(168) := previousCrc(8); xorBitMap(0)(169) := previousCrc(9); xorBitMap(0)(170) := previousCrc(10); xorBitMap(0)(172) := previousCrc(12); xorBitMap(0)(173) := previousCrc(13); xorBitMap(0)(174) := previousCrc(14); xorBitMap(0)(175) := previousCrc(15); xorBitMap(0)(176) := previousCrc(16); xorBitMap(0)(178) := previousCrc(18); xorBitMap(0)(181) := previousCrc(21); xorBitMap(0)(188) := previousCrc(28); xorBitMap(0)(189) := previousCrc(29); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(160) := previousCrc(0); xorBitMap(1)(161) := previousCrc(1); xorBitMap(1)(168) := previousCrc(8); xorBitMap(1)(171) := previousCrc(11); xorBitMap(1)(172) := previousCrc(12); xorBitMap(1)(177) := previousCrc(17); xorBitMap(1)(178) := previousCrc(18); xorBitMap(1)(179) := previousCrc(19); xorBitMap(1)(181) := previousCrc(21); xorBitMap(1)(182) := previousCrc(22); xorBitMap(1)(188) := previousCrc(28); xorBitMap(1)(190) := previousCrc(30); xorBitMap(1)(191) := previousCrc(31); 
      xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(160) := previousCrc(0); xorBitMap(2)(161) := previousCrc(1); xorBitMap(2)(162) := previousCrc(2); xorBitMap(2)(168) := previousCrc(8); xorBitMap(2)(170) := previousCrc(10); xorBitMap(2)(174) := previousCrc(14); xorBitMap(2)(175) := previousCrc(15); xorBitMap(2)(176) := previousCrc(16); xorBitMap(2)(179) := previousCrc(19); xorBitMap(2)(180) := previousCrc(20); xorBitMap(2)(181) := previousCrc(21); xorBitMap(2)(182) := previousCrc(22); xorBitMap(2)(183) := previousCrc(23); xorBitMap(2)(188) := previousCrc(28); 
      xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(161) := previousCrc(1); xorBitMap(3)(162) := previousCrc(2); xorBitMap(3)(163) := previousCrc(3); xorBitMap(3)(169) := previousCrc(9); xorBitMap(3)(171) := previousCrc(11); xorBitMap(3)(175) := previousCrc(15); xorBitMap(3)(176) := previousCrc(16); xorBitMap(3)(177) := previousCrc(17); xorBitMap(3)(180) := previousCrc(20); xorBitMap(3)(181) := previousCrc(21); xorBitMap(3)(182) := previousCrc(22); xorBitMap(3)(183) := previousCrc(23); xorBitMap(3)(184) := previousCrc(24); xorBitMap(3)(189) := previousCrc(29); 
      xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(162) := previousCrc(2); xorBitMap(4)(163) := previousCrc(3); xorBitMap(4)(164) := previousCrc(4); xorBitMap(4)(168) := previousCrc(8); xorBitMap(4)(169) := previousCrc(9); xorBitMap(4)(173) := previousCrc(13); xorBitMap(4)(174) := previousCrc(14); xorBitMap(4)(175) := previousCrc(15); xorBitMap(4)(177) := previousCrc(17); xorBitMap(4)(182) := previousCrc(22); xorBitMap(4)(183) := previousCrc(23); xorBitMap(4)(184) := previousCrc(24); xorBitMap(4)(185) := previousCrc(25); xorBitMap(4)(188) := previousCrc(28); xorBitMap(4)(189) := previousCrc(29); xorBitMap(4)(190) := previousCrc(30); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(163) := previousCrc(3); xorBitMap(5)(164) := previousCrc(4); xorBitMap(5)(165) := previousCrc(5); xorBitMap(5)(168) := previousCrc(8); xorBitMap(5)(172) := previousCrc(12); xorBitMap(5)(173) := previousCrc(13); xorBitMap(5)(181) := previousCrc(21); xorBitMap(5)(183) := previousCrc(23); xorBitMap(5)(184) := previousCrc(24); xorBitMap(5)(185) := previousCrc(25); xorBitMap(5)(186) := previousCrc(26); xorBitMap(5)(188) := previousCrc(28); xorBitMap(5)(190) := previousCrc(30); 
      xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(164) := previousCrc(4); xorBitMap(6)(165) := previousCrc(5); xorBitMap(6)(166) := previousCrc(6); xorBitMap(6)(169) := previousCrc(9); xorBitMap(6)(173) := previousCrc(13); xorBitMap(6)(174) := previousCrc(14); xorBitMap(6)(182) := previousCrc(22); xorBitMap(6)(184) := previousCrc(24); xorBitMap(6)(185) := previousCrc(25); xorBitMap(6)(186) := previousCrc(26); xorBitMap(6)(187) := previousCrc(27); xorBitMap(6)(189) := previousCrc(29); xorBitMap(6)(191) := previousCrc(31); 
      xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(160) := previousCrc(0); xorBitMap(7)(165) := previousCrc(5); xorBitMap(7)(166) := previousCrc(6); xorBitMap(7)(167) := previousCrc(7); xorBitMap(7)(168) := previousCrc(8); xorBitMap(7)(169) := previousCrc(9); xorBitMap(7)(172) := previousCrc(12); xorBitMap(7)(173) := previousCrc(13); xorBitMap(7)(176) := previousCrc(16); xorBitMap(7)(178) := previousCrc(18); xorBitMap(7)(181) := previousCrc(21); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(185) := previousCrc(25); xorBitMap(7)(186) := previousCrc(26); xorBitMap(7)(187) := previousCrc(27); xorBitMap(7)(189) := previousCrc(29); xorBitMap(7)(190) := previousCrc(30); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(161) := previousCrc(1); xorBitMap(8)(166) := previousCrc(6); xorBitMap(8)(167) := previousCrc(7); xorBitMap(8)(172) := previousCrc(12); xorBitMap(8)(175) := previousCrc(15); xorBitMap(8)(176) := previousCrc(16); xorBitMap(8)(177) := previousCrc(17); xorBitMap(8)(178) := previousCrc(18); xorBitMap(8)(179) := previousCrc(19); xorBitMap(8)(181) := previousCrc(21); xorBitMap(8)(182) := previousCrc(22); xorBitMap(8)(184) := previousCrc(24); xorBitMap(8)(186) := previousCrc(26); xorBitMap(8)(187) := previousCrc(27); xorBitMap(8)(189) := previousCrc(29); xorBitMap(8)(190) := previousCrc(30); 
      xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(162) := previousCrc(2); xorBitMap(9)(167) := previousCrc(7); xorBitMap(9)(168) := previousCrc(8); xorBitMap(9)(173) := previousCrc(13); xorBitMap(9)(176) := previousCrc(16); xorBitMap(9)(177) := previousCrc(17); xorBitMap(9)(178) := previousCrc(18); xorBitMap(9)(179) := previousCrc(19); xorBitMap(9)(180) := previousCrc(20); xorBitMap(9)(182) := previousCrc(22); xorBitMap(9)(183) := previousCrc(23); xorBitMap(9)(185) := previousCrc(25); xorBitMap(9)(187) := previousCrc(27); xorBitMap(9)(188) := previousCrc(28); xorBitMap(9)(190) := previousCrc(30); xorBitMap(9)(191) := previousCrc(31); 
      xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(160) := previousCrc(0); xorBitMap(10)(163) := previousCrc(3); xorBitMap(10)(170) := previousCrc(10); xorBitMap(10)(172) := previousCrc(12); xorBitMap(10)(173) := previousCrc(13); xorBitMap(10)(175) := previousCrc(15); xorBitMap(10)(176) := previousCrc(16); xorBitMap(10)(177) := previousCrc(17); xorBitMap(10)(179) := previousCrc(19); xorBitMap(10)(180) := previousCrc(20); xorBitMap(10)(183) := previousCrc(23); xorBitMap(10)(184) := previousCrc(24); xorBitMap(10)(186) := previousCrc(26); 
      xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(160) := previousCrc(0); xorBitMap(11)(161) := previousCrc(1); xorBitMap(11)(164) := previousCrc(4); xorBitMap(11)(168) := previousCrc(8); xorBitMap(11)(169) := previousCrc(9); xorBitMap(11)(170) := previousCrc(10); xorBitMap(11)(171) := previousCrc(11); xorBitMap(11)(172) := previousCrc(12); xorBitMap(11)(175) := previousCrc(15); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(180) := previousCrc(20); xorBitMap(11)(184) := previousCrc(24); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(187) := previousCrc(27); xorBitMap(11)(188) := previousCrc(28); xorBitMap(11)(189) := previousCrc(29); xorBitMap(11)(191) := previousCrc(31); 
      xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(161) := previousCrc(1); xorBitMap(12)(162) := previousCrc(2); xorBitMap(12)(165) := previousCrc(5); xorBitMap(12)(168) := previousCrc(8); xorBitMap(12)(171) := previousCrc(11); xorBitMap(12)(174) := previousCrc(14); xorBitMap(12)(175) := previousCrc(15); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(186) := previousCrc(26); xorBitMap(12)(190) := previousCrc(30); xorBitMap(12)(191) := previousCrc(31); 
      xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(160) := previousCrc(0); xorBitMap(13)(162) := previousCrc(2); xorBitMap(13)(163) := previousCrc(3); xorBitMap(13)(166) := previousCrc(6); xorBitMap(13)(169) := previousCrc(9); xorBitMap(13)(172) := previousCrc(12); xorBitMap(13)(175) := previousCrc(15); xorBitMap(13)(176) := previousCrc(16); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(187) := previousCrc(27); xorBitMap(13)(191) := previousCrc(31); 
      xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(161) := previousCrc(1); xorBitMap(14)(163) := previousCrc(3); xorBitMap(14)(164) := previousCrc(4); xorBitMap(14)(167) := previousCrc(7); xorBitMap(14)(170) := previousCrc(10); xorBitMap(14)(173) := previousCrc(13); xorBitMap(14)(176) := previousCrc(16); xorBitMap(14)(177) := previousCrc(17); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(188) := previousCrc(28); 
      xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(160) := previousCrc(0); xorBitMap(15)(162) := previousCrc(2); xorBitMap(15)(164) := previousCrc(4); xorBitMap(15)(165) := previousCrc(5); xorBitMap(15)(168) := previousCrc(8); xorBitMap(15)(171) := previousCrc(11); xorBitMap(15)(174) := previousCrc(14); xorBitMap(15)(177) := previousCrc(17); xorBitMap(15)(178) := previousCrc(18); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(189) := previousCrc(29); 
      xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(161) := previousCrc(1); xorBitMap(16)(163) := previousCrc(3); xorBitMap(16)(165) := previousCrc(5); xorBitMap(16)(166) := previousCrc(6); xorBitMap(16)(168) := previousCrc(8); xorBitMap(16)(170) := previousCrc(10); xorBitMap(16)(173) := previousCrc(13); xorBitMap(16)(174) := previousCrc(14); xorBitMap(16)(176) := previousCrc(16); xorBitMap(16)(179) := previousCrc(19); xorBitMap(16)(181) := previousCrc(21); xorBitMap(16)(188) := previousCrc(28); xorBitMap(16)(190) := previousCrc(30); xorBitMap(16)(191) := previousCrc(31); 
      xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(162) := previousCrc(2); xorBitMap(17)(164) := previousCrc(4); xorBitMap(17)(166) := previousCrc(6); xorBitMap(17)(167) := previousCrc(7); xorBitMap(17)(169) := previousCrc(9); xorBitMap(17)(171) := previousCrc(11); xorBitMap(17)(174) := previousCrc(14); xorBitMap(17)(175) := previousCrc(15); xorBitMap(17)(177) := previousCrc(17); xorBitMap(17)(180) := previousCrc(20); xorBitMap(17)(182) := previousCrc(22); xorBitMap(17)(189) := previousCrc(29); xorBitMap(17)(191) := previousCrc(31); 
      xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(163) := previousCrc(3); xorBitMap(18)(165) := previousCrc(5); xorBitMap(18)(167) := previousCrc(7); xorBitMap(18)(168) := previousCrc(8); xorBitMap(18)(170) := previousCrc(10); xorBitMap(18)(172) := previousCrc(12); xorBitMap(18)(175) := previousCrc(15); xorBitMap(18)(176) := previousCrc(16); xorBitMap(18)(178) := previousCrc(18); xorBitMap(18)(181) := previousCrc(21); xorBitMap(18)(183) := previousCrc(23); xorBitMap(18)(190) := previousCrc(30); 
      xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(160) := previousCrc(0); xorBitMap(19)(164) := previousCrc(4); xorBitMap(19)(166) := previousCrc(6); xorBitMap(19)(168) := previousCrc(8); xorBitMap(19)(169) := previousCrc(9); xorBitMap(19)(171) := previousCrc(11); xorBitMap(19)(173) := previousCrc(13); xorBitMap(19)(176) := previousCrc(16); xorBitMap(19)(177) := previousCrc(17); xorBitMap(19)(179) := previousCrc(19); xorBitMap(19)(182) := previousCrc(22); xorBitMap(19)(184) := previousCrc(24); xorBitMap(19)(191) := previousCrc(31); 
      xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(160) := previousCrc(0); xorBitMap(20)(161) := previousCrc(1); xorBitMap(20)(165) := previousCrc(5); xorBitMap(20)(167) := previousCrc(7); xorBitMap(20)(169) := previousCrc(9); xorBitMap(20)(170) := previousCrc(10); xorBitMap(20)(172) := previousCrc(12); xorBitMap(20)(174) := previousCrc(14); xorBitMap(20)(177) := previousCrc(17); xorBitMap(20)(178) := previousCrc(18); xorBitMap(20)(180) := previousCrc(20); xorBitMap(20)(183) := previousCrc(23); xorBitMap(20)(185) := previousCrc(25); 
      xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(161) := previousCrc(1); xorBitMap(21)(162) := previousCrc(2); xorBitMap(21)(166) := previousCrc(6); xorBitMap(21)(168) := previousCrc(8); xorBitMap(21)(170) := previousCrc(10); xorBitMap(21)(171) := previousCrc(11); xorBitMap(21)(173) := previousCrc(13); xorBitMap(21)(175) := previousCrc(15); xorBitMap(21)(178) := previousCrc(18); xorBitMap(21)(179) := previousCrc(19); xorBitMap(21)(181) := previousCrc(21); xorBitMap(21)(184) := previousCrc(24); xorBitMap(21)(186) := previousCrc(26); 
      xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(160) := previousCrc(0); xorBitMap(22)(162) := previousCrc(2); xorBitMap(22)(163) := previousCrc(3); xorBitMap(22)(167) := previousCrc(7); xorBitMap(22)(168) := previousCrc(8); xorBitMap(22)(170) := previousCrc(10); xorBitMap(22)(171) := previousCrc(11); xorBitMap(22)(173) := previousCrc(13); xorBitMap(22)(175) := previousCrc(15); xorBitMap(22)(178) := previousCrc(18); xorBitMap(22)(179) := previousCrc(19); xorBitMap(22)(180) := previousCrc(20); xorBitMap(22)(181) := previousCrc(21); xorBitMap(22)(182) := previousCrc(22); xorBitMap(22)(185) := previousCrc(25); xorBitMap(22)(187) := previousCrc(27); xorBitMap(22)(188) := previousCrc(28); xorBitMap(22)(189) := previousCrc(29); xorBitMap(22)(191) := previousCrc(31); 
      xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(160) := previousCrc(0); xorBitMap(23)(161) := previousCrc(1); xorBitMap(23)(163) := previousCrc(3); xorBitMap(23)(164) := previousCrc(4); xorBitMap(23)(170) := previousCrc(10); xorBitMap(23)(171) := previousCrc(11); xorBitMap(23)(173) := previousCrc(13); xorBitMap(23)(175) := previousCrc(15); xorBitMap(23)(178) := previousCrc(18); xorBitMap(23)(179) := previousCrc(19); xorBitMap(23)(180) := previousCrc(20); xorBitMap(23)(182) := previousCrc(22); xorBitMap(23)(183) := previousCrc(23); xorBitMap(23)(186) := previousCrc(26); xorBitMap(23)(190) := previousCrc(30); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(160) := previousCrc(0); xorBitMap(24)(161) := previousCrc(1); xorBitMap(24)(162) := previousCrc(2); xorBitMap(24)(164) := previousCrc(4); xorBitMap(24)(165) := previousCrc(5); xorBitMap(24)(171) := previousCrc(11); xorBitMap(24)(172) := previousCrc(12); xorBitMap(24)(174) := previousCrc(14); xorBitMap(24)(176) := previousCrc(16); xorBitMap(24)(179) := previousCrc(19); xorBitMap(24)(180) := previousCrc(20); xorBitMap(24)(181) := previousCrc(21); xorBitMap(24)(183) := previousCrc(23); xorBitMap(24)(184) := previousCrc(24); xorBitMap(24)(187) := previousCrc(27); xorBitMap(24)(191) := previousCrc(31); 
      xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(161) := previousCrc(1); xorBitMap(25)(162) := previousCrc(2); xorBitMap(25)(163) := previousCrc(3); xorBitMap(25)(165) := previousCrc(5); xorBitMap(25)(166) := previousCrc(6); xorBitMap(25)(172) := previousCrc(12); xorBitMap(25)(173) := previousCrc(13); xorBitMap(25)(175) := previousCrc(15); xorBitMap(25)(177) := previousCrc(17); xorBitMap(25)(180) := previousCrc(20); xorBitMap(25)(181) := previousCrc(21); xorBitMap(25)(182) := previousCrc(22); xorBitMap(25)(184) := previousCrc(24); xorBitMap(25)(185) := previousCrc(25); xorBitMap(25)(188) := previousCrc(28); 
      xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(162) := previousCrc(2); xorBitMap(26)(163) := previousCrc(3); xorBitMap(26)(164) := previousCrc(4); xorBitMap(26)(166) := previousCrc(6); xorBitMap(26)(167) := previousCrc(7); xorBitMap(26)(168) := previousCrc(8); xorBitMap(26)(169) := previousCrc(9); xorBitMap(26)(170) := previousCrc(10); xorBitMap(26)(172) := previousCrc(12); xorBitMap(26)(175) := previousCrc(15); xorBitMap(26)(182) := previousCrc(22); xorBitMap(26)(183) := previousCrc(23); xorBitMap(26)(185) := previousCrc(25); xorBitMap(26)(186) := previousCrc(26); xorBitMap(26)(188) := previousCrc(28); xorBitMap(26)(191) := previousCrc(31); 
      xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(163) := previousCrc(3); xorBitMap(27)(164) := previousCrc(4); xorBitMap(27)(165) := previousCrc(5); xorBitMap(27)(167) := previousCrc(7); xorBitMap(27)(168) := previousCrc(8); xorBitMap(27)(169) := previousCrc(9); xorBitMap(27)(170) := previousCrc(10); xorBitMap(27)(171) := previousCrc(11); xorBitMap(27)(173) := previousCrc(13); xorBitMap(27)(176) := previousCrc(16); xorBitMap(27)(183) := previousCrc(23); xorBitMap(27)(184) := previousCrc(24); xorBitMap(27)(186) := previousCrc(26); xorBitMap(27)(187) := previousCrc(27); xorBitMap(27)(189) := previousCrc(29); 
      xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(164) := previousCrc(4); xorBitMap(28)(165) := previousCrc(5); xorBitMap(28)(166) := previousCrc(6); xorBitMap(28)(168) := previousCrc(8); xorBitMap(28)(169) := previousCrc(9); xorBitMap(28)(170) := previousCrc(10); xorBitMap(28)(171) := previousCrc(11); xorBitMap(28)(172) := previousCrc(12); xorBitMap(28)(174) := previousCrc(14); xorBitMap(28)(177) := previousCrc(17); xorBitMap(28)(184) := previousCrc(24); xorBitMap(28)(185) := previousCrc(25); xorBitMap(28)(187) := previousCrc(27); xorBitMap(28)(188) := previousCrc(28); xorBitMap(28)(190) := previousCrc(30); 
      xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(165) := previousCrc(5); xorBitMap(29)(166) := previousCrc(6); xorBitMap(29)(167) := previousCrc(7); xorBitMap(29)(169) := previousCrc(9); xorBitMap(29)(170) := previousCrc(10); xorBitMap(29)(171) := previousCrc(11); xorBitMap(29)(172) := previousCrc(12); xorBitMap(29)(173) := previousCrc(13); xorBitMap(29)(175) := previousCrc(15); xorBitMap(29)(178) := previousCrc(18); xorBitMap(29)(185) := previousCrc(25); xorBitMap(29)(186) := previousCrc(26); xorBitMap(29)(188) := previousCrc(28); xorBitMap(29)(189) := previousCrc(29); xorBitMap(29)(191) := previousCrc(31); 
      xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(166) := previousCrc(6); xorBitMap(30)(167) := previousCrc(7); xorBitMap(30)(168) := previousCrc(8); xorBitMap(30)(170) := previousCrc(10); xorBitMap(30)(171) := previousCrc(11); xorBitMap(30)(172) := previousCrc(12); xorBitMap(30)(173) := previousCrc(13); xorBitMap(30)(174) := previousCrc(14); xorBitMap(30)(176) := previousCrc(16); xorBitMap(30)(179) := previousCrc(19); xorBitMap(30)(186) := previousCrc(26); xorBitMap(30)(187) := previousCrc(27); xorBitMap(30)(189) := previousCrc(29); xorBitMap(30)(190) := previousCrc(30); 
      xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(167) := previousCrc(7); xorBitMap(31)(168) := previousCrc(8); xorBitMap(31)(169) := previousCrc(9); xorBitMap(31)(171) := previousCrc(11); xorBitMap(31)(172) := previousCrc(12); xorBitMap(31)(173) := previousCrc(13); xorBitMap(31)(174) := previousCrc(14); xorBitMap(31)(175) := previousCrc(15); xorBitMap(31)(177) := previousCrc(17); xorBitMap(31)(180) := previousCrc(20); xorBitMap(31)(187) := previousCrc(27); xorBitMap(31)(188) := previousCrc(28); xorBitMap(31)(190) := previousCrc(30); xorBitMap(31)(191) := previousCrc(31); 
   end procedure;

   procedure xorBitMap7Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(55 downto 0)) is 
   begin
      xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(160) := previousCrc(0); xorBitMap(0)(161) := previousCrc(1); xorBitMap(0)(162) := previousCrc(2); xorBitMap(0)(164) := previousCrc(4); xorBitMap(0)(165) := previousCrc(5); xorBitMap(0)(166) := previousCrc(6); xorBitMap(0)(167) := previousCrc(7); xorBitMap(0)(168) := previousCrc(8); xorBitMap(0)(170) := previousCrc(10); xorBitMap(0)(173) := previousCrc(13); xorBitMap(0)(180) := previousCrc(20); xorBitMap(0)(181) := previousCrc(21); xorBitMap(0)(183) := previousCrc(23); xorBitMap(0)(184) := previousCrc(24); xorBitMap(0)(186) := previousCrc(26); xorBitMap(0)(189) := previousCrc(29); xorBitMap(0)(190) := previousCrc(30); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(160) := previousCrc(0); xorBitMap(1)(163) := previousCrc(3); xorBitMap(1)(164) := previousCrc(4); xorBitMap(1)(169) := previousCrc(9); xorBitMap(1)(170) := previousCrc(10); xorBitMap(1)(171) := previousCrc(11); xorBitMap(1)(173) := previousCrc(13); xorBitMap(1)(174) := previousCrc(14); xorBitMap(1)(180) := previousCrc(20); xorBitMap(1)(182) := previousCrc(22); xorBitMap(1)(183) := previousCrc(23); xorBitMap(1)(185) := previousCrc(25); xorBitMap(1)(186) := previousCrc(26); xorBitMap(1)(187) := previousCrc(27); xorBitMap(1)(189) := previousCrc(29); 
      xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(160) := previousCrc(0); xorBitMap(2)(162) := previousCrc(2); xorBitMap(2)(166) := previousCrc(6); xorBitMap(2)(167) := previousCrc(7); xorBitMap(2)(168) := previousCrc(8); xorBitMap(2)(171) := previousCrc(11); xorBitMap(2)(172) := previousCrc(12); xorBitMap(2)(173) := previousCrc(13); xorBitMap(2)(174) := previousCrc(14); xorBitMap(2)(175) := previousCrc(15); xorBitMap(2)(180) := previousCrc(20); xorBitMap(2)(187) := previousCrc(27); xorBitMap(2)(188) := previousCrc(28); xorBitMap(2)(189) := previousCrc(29); xorBitMap(2)(191) := previousCrc(31); 
      xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(161) := previousCrc(1); xorBitMap(3)(163) := previousCrc(3); xorBitMap(3)(167) := previousCrc(7); xorBitMap(3)(168) := previousCrc(8); xorBitMap(3)(169) := previousCrc(9); xorBitMap(3)(172) := previousCrc(12); xorBitMap(3)(173) := previousCrc(13); xorBitMap(3)(174) := previousCrc(14); xorBitMap(3)(175) := previousCrc(15); xorBitMap(3)(176) := previousCrc(16); xorBitMap(3)(181) := previousCrc(21); xorBitMap(3)(188) := previousCrc(28); xorBitMap(3)(189) := previousCrc(29); xorBitMap(3)(190) := previousCrc(30); 
      xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(160) := previousCrc(0); xorBitMap(4)(161) := previousCrc(1); xorBitMap(4)(165) := previousCrc(5); xorBitMap(4)(166) := previousCrc(6); xorBitMap(4)(167) := previousCrc(7); xorBitMap(4)(169) := previousCrc(9); xorBitMap(4)(174) := previousCrc(14); xorBitMap(4)(175) := previousCrc(15); xorBitMap(4)(176) := previousCrc(16); xorBitMap(4)(177) := previousCrc(17); xorBitMap(4)(180) := previousCrc(20); xorBitMap(4)(181) := previousCrc(21); xorBitMap(4)(182) := previousCrc(22); xorBitMap(4)(183) := previousCrc(23); xorBitMap(4)(184) := previousCrc(24); xorBitMap(4)(186) := previousCrc(26); 
      xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(160) := previousCrc(0); xorBitMap(5)(164) := previousCrc(4); xorBitMap(5)(165) := previousCrc(5); xorBitMap(5)(173) := previousCrc(13); xorBitMap(5)(175) := previousCrc(15); xorBitMap(5)(176) := previousCrc(16); xorBitMap(5)(177) := previousCrc(17); xorBitMap(5)(178) := previousCrc(18); xorBitMap(5)(180) := previousCrc(20); xorBitMap(5)(182) := previousCrc(22); xorBitMap(5)(185) := previousCrc(25); xorBitMap(5)(186) := previousCrc(26); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(189) := previousCrc(29); xorBitMap(5)(190) := previousCrc(30); xorBitMap(5)(191) := previousCrc(31); 
      xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(161) := previousCrc(1); xorBitMap(6)(165) := previousCrc(5); xorBitMap(6)(166) := previousCrc(6); xorBitMap(6)(174) := previousCrc(14); xorBitMap(6)(176) := previousCrc(16); xorBitMap(6)(177) := previousCrc(17); xorBitMap(6)(178) := previousCrc(18); xorBitMap(6)(179) := previousCrc(19); xorBitMap(6)(181) := previousCrc(21); xorBitMap(6)(183) := previousCrc(23); xorBitMap(6)(186) := previousCrc(26); xorBitMap(6)(187) := previousCrc(27); xorBitMap(6)(188) := previousCrc(28); xorBitMap(6)(190) := previousCrc(30); xorBitMap(6)(191) := previousCrc(31); 
      xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(160) := previousCrc(0); xorBitMap(7)(161) := previousCrc(1); xorBitMap(7)(164) := previousCrc(4); xorBitMap(7)(165) := previousCrc(5); xorBitMap(7)(168) := previousCrc(8); xorBitMap(7)(170) := previousCrc(10); xorBitMap(7)(173) := previousCrc(13); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(177) := previousCrc(17); xorBitMap(7)(178) := previousCrc(18); xorBitMap(7)(179) := previousCrc(19); xorBitMap(7)(181) := previousCrc(21); xorBitMap(7)(182) := previousCrc(22); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(186) := previousCrc(26); xorBitMap(7)(187) := previousCrc(27); xorBitMap(7)(188) := previousCrc(28); xorBitMap(7)(190) := previousCrc(30); 
      xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(164) := previousCrc(4); xorBitMap(8)(167) := previousCrc(7); xorBitMap(8)(168) := previousCrc(8); xorBitMap(8)(169) := previousCrc(9); xorBitMap(8)(170) := previousCrc(10); xorBitMap(8)(171) := previousCrc(11); xorBitMap(8)(173) := previousCrc(13); xorBitMap(8)(174) := previousCrc(14); xorBitMap(8)(176) := previousCrc(16); xorBitMap(8)(178) := previousCrc(18); xorBitMap(8)(179) := previousCrc(19); xorBitMap(8)(181) := previousCrc(21); xorBitMap(8)(182) := previousCrc(22); xorBitMap(8)(186) := previousCrc(26); xorBitMap(8)(187) := previousCrc(27); xorBitMap(8)(188) := previousCrc(28); xorBitMap(8)(190) := previousCrc(30); 
      xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(160) := previousCrc(0); xorBitMap(9)(165) := previousCrc(5); xorBitMap(9)(168) := previousCrc(8); xorBitMap(9)(169) := previousCrc(9); xorBitMap(9)(170) := previousCrc(10); xorBitMap(9)(171) := previousCrc(11); xorBitMap(9)(172) := previousCrc(12); xorBitMap(9)(174) := previousCrc(14); xorBitMap(9)(175) := previousCrc(15); xorBitMap(9)(177) := previousCrc(17); xorBitMap(9)(179) := previousCrc(19); xorBitMap(9)(180) := previousCrc(20); xorBitMap(9)(182) := previousCrc(22); xorBitMap(9)(183) := previousCrc(23); xorBitMap(9)(187) := previousCrc(27); xorBitMap(9)(188) := previousCrc(28); xorBitMap(9)(189) := previousCrc(29); xorBitMap(9)(191) := previousCrc(31); 
      xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(162) := previousCrc(2); xorBitMap(10)(164) := previousCrc(4); xorBitMap(10)(165) := previousCrc(5); xorBitMap(10)(167) := previousCrc(7); xorBitMap(10)(168) := previousCrc(8); xorBitMap(10)(169) := previousCrc(9); xorBitMap(10)(171) := previousCrc(11); xorBitMap(10)(172) := previousCrc(12); xorBitMap(10)(175) := previousCrc(15); xorBitMap(10)(176) := previousCrc(16); xorBitMap(10)(178) := previousCrc(18); xorBitMap(10)(186) := previousCrc(26); xorBitMap(10)(188) := previousCrc(28); xorBitMap(10)(191) := previousCrc(31); 
      xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(160) := previousCrc(0); xorBitMap(11)(161) := previousCrc(1); xorBitMap(11)(162) := previousCrc(2); xorBitMap(11)(163) := previousCrc(3); xorBitMap(11)(164) := previousCrc(4); xorBitMap(11)(167) := previousCrc(7); xorBitMap(11)(169) := previousCrc(9); xorBitMap(11)(172) := previousCrc(12); xorBitMap(11)(176) := previousCrc(16); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(179) := previousCrc(19); xorBitMap(11)(180) := previousCrc(20); xorBitMap(11)(181) := previousCrc(21); xorBitMap(11)(183) := previousCrc(23); xorBitMap(11)(184) := previousCrc(24); xorBitMap(11)(186) := previousCrc(26); xorBitMap(11)(187) := previousCrc(27); xorBitMap(11)(190) := previousCrc(30); xorBitMap(11)(191) := previousCrc(31); 
      xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(160) := previousCrc(0); xorBitMap(12)(163) := previousCrc(3); xorBitMap(12)(166) := previousCrc(6); xorBitMap(12)(167) := previousCrc(7); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(178) := previousCrc(18); xorBitMap(12)(182) := previousCrc(22); xorBitMap(12)(183) := previousCrc(23); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(186) := previousCrc(26); xorBitMap(12)(187) := previousCrc(27); xorBitMap(12)(188) := previousCrc(28); xorBitMap(12)(189) := previousCrc(29); xorBitMap(12)(190) := previousCrc(30); 
      xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(161) := previousCrc(1); xorBitMap(13)(164) := previousCrc(4); xorBitMap(13)(167) := previousCrc(7); xorBitMap(13)(168) := previousCrc(8); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(179) := previousCrc(19); xorBitMap(13)(183) := previousCrc(23); xorBitMap(13)(184) := previousCrc(24); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(187) := previousCrc(27); xorBitMap(13)(188) := previousCrc(28); xorBitMap(13)(189) := previousCrc(29); xorBitMap(13)(190) := previousCrc(30); xorBitMap(13)(191) := previousCrc(31); 
      xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(162) := previousCrc(2); xorBitMap(14)(165) := previousCrc(5); xorBitMap(14)(168) := previousCrc(8); xorBitMap(14)(169) := previousCrc(9); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(180) := previousCrc(20); xorBitMap(14)(184) := previousCrc(24); xorBitMap(14)(185) := previousCrc(25); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(188) := previousCrc(28); xorBitMap(14)(189) := previousCrc(29); xorBitMap(14)(190) := previousCrc(30); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(160) := previousCrc(0); xorBitMap(15)(163) := previousCrc(3); xorBitMap(15)(166) := previousCrc(6); xorBitMap(15)(169) := previousCrc(9); xorBitMap(15)(170) := previousCrc(10); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(181) := previousCrc(21); xorBitMap(15)(185) := previousCrc(25); xorBitMap(15)(186) := previousCrc(26); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(189) := previousCrc(29); xorBitMap(15)(190) := previousCrc(30); xorBitMap(15)(191) := previousCrc(31); 
      xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(160) := previousCrc(0); xorBitMap(16)(162) := previousCrc(2); xorBitMap(16)(165) := previousCrc(5); xorBitMap(16)(166) := previousCrc(6); xorBitMap(16)(168) := previousCrc(8); xorBitMap(16)(171) := previousCrc(11); xorBitMap(16)(173) := previousCrc(13); xorBitMap(16)(180) := previousCrc(20); xorBitMap(16)(182) := previousCrc(22); xorBitMap(16)(183) := previousCrc(23); xorBitMap(16)(184) := previousCrc(24); xorBitMap(16)(187) := previousCrc(27); 
      xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(161) := previousCrc(1); xorBitMap(17)(163) := previousCrc(3); xorBitMap(17)(166) := previousCrc(6); xorBitMap(17)(167) := previousCrc(7); xorBitMap(17)(169) := previousCrc(9); xorBitMap(17)(172) := previousCrc(12); xorBitMap(17)(174) := previousCrc(14); xorBitMap(17)(181) := previousCrc(21); xorBitMap(17)(183) := previousCrc(23); xorBitMap(17)(184) := previousCrc(24); xorBitMap(17)(185) := previousCrc(25); xorBitMap(17)(188) := previousCrc(28); 
      xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(160) := previousCrc(0); xorBitMap(18)(162) := previousCrc(2); xorBitMap(18)(164) := previousCrc(4); xorBitMap(18)(167) := previousCrc(7); xorBitMap(18)(168) := previousCrc(8); xorBitMap(18)(170) := previousCrc(10); xorBitMap(18)(173) := previousCrc(13); xorBitMap(18)(175) := previousCrc(15); xorBitMap(18)(182) := previousCrc(22); xorBitMap(18)(184) := previousCrc(24); xorBitMap(18)(185) := previousCrc(25); xorBitMap(18)(186) := previousCrc(26); xorBitMap(18)(189) := previousCrc(29); 
      xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(160) := previousCrc(0); xorBitMap(19)(161) := previousCrc(1); xorBitMap(19)(163) := previousCrc(3); xorBitMap(19)(165) := previousCrc(5); xorBitMap(19)(168) := previousCrc(8); xorBitMap(19)(169) := previousCrc(9); xorBitMap(19)(171) := previousCrc(11); xorBitMap(19)(174) := previousCrc(14); xorBitMap(19)(176) := previousCrc(16); xorBitMap(19)(183) := previousCrc(23); xorBitMap(19)(185) := previousCrc(25); xorBitMap(19)(186) := previousCrc(26); xorBitMap(19)(187) := previousCrc(27); xorBitMap(19)(190) := previousCrc(30); 
      xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(161) := previousCrc(1); xorBitMap(20)(162) := previousCrc(2); xorBitMap(20)(164) := previousCrc(4); xorBitMap(20)(166) := previousCrc(6); xorBitMap(20)(169) := previousCrc(9); xorBitMap(20)(170) := previousCrc(10); xorBitMap(20)(172) := previousCrc(12); xorBitMap(20)(175) := previousCrc(15); xorBitMap(20)(177) := previousCrc(17); xorBitMap(20)(184) := previousCrc(24); xorBitMap(20)(186) := previousCrc(26); xorBitMap(20)(187) := previousCrc(27); xorBitMap(20)(188) := previousCrc(28); xorBitMap(20)(191) := previousCrc(31); 
      xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(160) := previousCrc(0); xorBitMap(21)(162) := previousCrc(2); xorBitMap(21)(163) := previousCrc(3); xorBitMap(21)(165) := previousCrc(5); xorBitMap(21)(167) := previousCrc(7); xorBitMap(21)(170) := previousCrc(10); xorBitMap(21)(171) := previousCrc(11); xorBitMap(21)(173) := previousCrc(13); xorBitMap(21)(176) := previousCrc(16); xorBitMap(21)(178) := previousCrc(18); xorBitMap(21)(185) := previousCrc(25); xorBitMap(21)(187) := previousCrc(27); xorBitMap(21)(188) := previousCrc(28); xorBitMap(21)(189) := previousCrc(29); 
      xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(160) := previousCrc(0); xorBitMap(22)(162) := previousCrc(2); xorBitMap(22)(163) := previousCrc(3); xorBitMap(22)(165) := previousCrc(5); xorBitMap(22)(167) := previousCrc(7); xorBitMap(22)(170) := previousCrc(10); xorBitMap(22)(171) := previousCrc(11); xorBitMap(22)(172) := previousCrc(12); xorBitMap(22)(173) := previousCrc(13); xorBitMap(22)(174) := previousCrc(14); xorBitMap(22)(177) := previousCrc(17); xorBitMap(22)(179) := previousCrc(19); xorBitMap(22)(180) := previousCrc(20); xorBitMap(22)(181) := previousCrc(21); xorBitMap(22)(183) := previousCrc(23); xorBitMap(22)(184) := previousCrc(24); xorBitMap(22)(188) := previousCrc(28); xorBitMap(22)(191) := previousCrc(31); 
      xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(162) := previousCrc(2); xorBitMap(23)(163) := previousCrc(3); xorBitMap(23)(165) := previousCrc(5); xorBitMap(23)(167) := previousCrc(7); xorBitMap(23)(170) := previousCrc(10); xorBitMap(23)(171) := previousCrc(11); xorBitMap(23)(172) := previousCrc(12); xorBitMap(23)(174) := previousCrc(14); xorBitMap(23)(175) := previousCrc(15); xorBitMap(23)(178) := previousCrc(18); xorBitMap(23)(182) := previousCrc(22); xorBitMap(23)(183) := previousCrc(23); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(186) := previousCrc(26); xorBitMap(23)(190) := previousCrc(30); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(163) := previousCrc(3); xorBitMap(24)(164) := previousCrc(4); xorBitMap(24)(166) := previousCrc(6); xorBitMap(24)(168) := previousCrc(8); xorBitMap(24)(171) := previousCrc(11); xorBitMap(24)(172) := previousCrc(12); xorBitMap(24)(173) := previousCrc(13); xorBitMap(24)(175) := previousCrc(15); xorBitMap(24)(176) := previousCrc(16); xorBitMap(24)(179) := previousCrc(19); xorBitMap(24)(183) := previousCrc(23); xorBitMap(24)(184) := previousCrc(24); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(187) := previousCrc(27); xorBitMap(24)(191) := previousCrc(31); 
      xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(164) := previousCrc(4); xorBitMap(25)(165) := previousCrc(5); xorBitMap(25)(167) := previousCrc(7); xorBitMap(25)(169) := previousCrc(9); xorBitMap(25)(172) := previousCrc(12); xorBitMap(25)(173) := previousCrc(13); xorBitMap(25)(174) := previousCrc(14); xorBitMap(25)(176) := previousCrc(16); xorBitMap(25)(177) := previousCrc(17); xorBitMap(25)(180) := previousCrc(20); xorBitMap(25)(184) := previousCrc(24); xorBitMap(25)(185) := previousCrc(25); xorBitMap(25)(187) := previousCrc(27); xorBitMap(25)(188) := previousCrc(28); 
      xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(160) := previousCrc(0); xorBitMap(26)(161) := previousCrc(1); xorBitMap(26)(162) := previousCrc(2); xorBitMap(26)(164) := previousCrc(4); xorBitMap(26)(167) := previousCrc(7); xorBitMap(26)(174) := previousCrc(14); xorBitMap(26)(175) := previousCrc(15); xorBitMap(26)(177) := previousCrc(17); xorBitMap(26)(178) := previousCrc(18); xorBitMap(26)(180) := previousCrc(20); xorBitMap(26)(183) := previousCrc(23); xorBitMap(26)(184) := previousCrc(24); xorBitMap(26)(185) := previousCrc(25); xorBitMap(26)(188) := previousCrc(28); xorBitMap(26)(190) := previousCrc(30); xorBitMap(26)(191) := previousCrc(31); 
      xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(160) := previousCrc(0); xorBitMap(27)(161) := previousCrc(1); xorBitMap(27)(162) := previousCrc(2); xorBitMap(27)(163) := previousCrc(3); xorBitMap(27)(165) := previousCrc(5); xorBitMap(27)(168) := previousCrc(8); xorBitMap(27)(175) := previousCrc(15); xorBitMap(27)(176) := previousCrc(16); xorBitMap(27)(178) := previousCrc(18); xorBitMap(27)(179) := previousCrc(19); xorBitMap(27)(181) := previousCrc(21); xorBitMap(27)(184) := previousCrc(24); xorBitMap(27)(185) := previousCrc(25); xorBitMap(27)(186) := previousCrc(26); xorBitMap(27)(189) := previousCrc(29); xorBitMap(27)(191) := previousCrc(31); 
      xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(160) := previousCrc(0); xorBitMap(28)(161) := previousCrc(1); xorBitMap(28)(162) := previousCrc(2); xorBitMap(28)(163) := previousCrc(3); xorBitMap(28)(164) := previousCrc(4); xorBitMap(28)(166) := previousCrc(6); xorBitMap(28)(169) := previousCrc(9); xorBitMap(28)(176) := previousCrc(16); xorBitMap(28)(177) := previousCrc(17); xorBitMap(28)(179) := previousCrc(19); xorBitMap(28)(180) := previousCrc(20); xorBitMap(28)(182) := previousCrc(22); xorBitMap(28)(185) := previousCrc(25); xorBitMap(28)(186) := previousCrc(26); xorBitMap(28)(187) := previousCrc(27); xorBitMap(28)(190) := previousCrc(30); 
      xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(161) := previousCrc(1); xorBitMap(29)(162) := previousCrc(2); xorBitMap(29)(163) := previousCrc(3); xorBitMap(29)(164) := previousCrc(4); xorBitMap(29)(165) := previousCrc(5); xorBitMap(29)(167) := previousCrc(7); xorBitMap(29)(170) := previousCrc(10); xorBitMap(29)(177) := previousCrc(17); xorBitMap(29)(178) := previousCrc(18); xorBitMap(29)(180) := previousCrc(20); xorBitMap(29)(181) := previousCrc(21); xorBitMap(29)(183) := previousCrc(23); xorBitMap(29)(186) := previousCrc(26); xorBitMap(29)(187) := previousCrc(27); xorBitMap(29)(188) := previousCrc(28); xorBitMap(29)(191) := previousCrc(31); 
      xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(160) := previousCrc(0); xorBitMap(30)(162) := previousCrc(2); xorBitMap(30)(163) := previousCrc(3); xorBitMap(30)(164) := previousCrc(4); xorBitMap(30)(165) := previousCrc(5); xorBitMap(30)(166) := previousCrc(6); xorBitMap(30)(168) := previousCrc(8); xorBitMap(30)(171) := previousCrc(11); xorBitMap(30)(178) := previousCrc(18); xorBitMap(30)(179) := previousCrc(19); xorBitMap(30)(181) := previousCrc(21); xorBitMap(30)(182) := previousCrc(22); xorBitMap(30)(184) := previousCrc(24); xorBitMap(30)(187) := previousCrc(27); xorBitMap(30)(188) := previousCrc(28); xorBitMap(30)(189) := previousCrc(29); 
      xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(160) := previousCrc(0); xorBitMap(31)(161) := previousCrc(1); xorBitMap(31)(163) := previousCrc(3); xorBitMap(31)(164) := previousCrc(4); xorBitMap(31)(165) := previousCrc(5); xorBitMap(31)(166) := previousCrc(6); xorBitMap(31)(167) := previousCrc(7); xorBitMap(31)(169) := previousCrc(9); xorBitMap(31)(172) := previousCrc(12); xorBitMap(31)(179) := previousCrc(19); xorBitMap(31)(180) := previousCrc(20); xorBitMap(31)(182) := previousCrc(22); xorBitMap(31)(183) := previousCrc(23); xorBitMap(31)(185) := previousCrc(25); xorBitMap(31)(188) := previousCrc(28); xorBitMap(31)(189) := previousCrc(29); xorBitMap(31)(190) := previousCrc(30); 
   end procedure;

   procedure xorBitMap8Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(63 downto 0)) is 
   begin
      xorBitMap(0)(63) := currentData(63); xorBitMap(0)(61) := currentData(61); xorBitMap(0)(60) := currentData(60); xorBitMap(0)(58) := currentData(58); xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(160) := previousCrc(0); xorBitMap(0)(162) := previousCrc(2); xorBitMap(0)(165) := previousCrc(5); xorBitMap(0)(172) := previousCrc(12); xorBitMap(0)(173) := previousCrc(13); xorBitMap(0)(175) := previousCrc(15); xorBitMap(0)(176) := previousCrc(16); xorBitMap(0)(178) := previousCrc(18); xorBitMap(0)(181) := previousCrc(21); xorBitMap(0)(182) := previousCrc(22); xorBitMap(0)(183) := previousCrc(23); xorBitMap(0)(186) := previousCrc(26); xorBitMap(0)(188) := previousCrc(28); xorBitMap(0)(189) := previousCrc(29); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(63) := currentData(63); xorBitMap(1)(62) := currentData(62); xorBitMap(1)(60) := currentData(60); xorBitMap(1)(59) := currentData(59); xorBitMap(1)(58) := currentData(58); xorBitMap(1)(56) := currentData(56); xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(161) := previousCrc(1); xorBitMap(1)(162) := previousCrc(2); xorBitMap(1)(163) := previousCrc(3); xorBitMap(1)(165) := previousCrc(5); xorBitMap(1)(166) := previousCrc(6); xorBitMap(1)(172) := previousCrc(12); xorBitMap(1)(174) := previousCrc(14); xorBitMap(1)(175) := previousCrc(15); xorBitMap(1)(177) := previousCrc(17); xorBitMap(1)(178) := previousCrc(18); xorBitMap(1)(179) := previousCrc(19); xorBitMap(1)(181) := previousCrc(21); xorBitMap(1)(184) := previousCrc(24); xorBitMap(1)(186) := previousCrc(26); xorBitMap(1)(187) := previousCrc(27); xorBitMap(1)(188) := previousCrc(28); xorBitMap(1)(190) := previousCrc(30); xorBitMap(1)(191) := previousCrc(31); 
      xorBitMap(2)(59) := currentData(59); xorBitMap(2)(58) := currentData(58); xorBitMap(2)(57) := currentData(57); xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(160) := previousCrc(0); xorBitMap(2)(163) := previousCrc(3); xorBitMap(2)(164) := previousCrc(4); xorBitMap(2)(165) := previousCrc(5); xorBitMap(2)(166) := previousCrc(6); xorBitMap(2)(167) := previousCrc(7); xorBitMap(2)(172) := previousCrc(12); xorBitMap(2)(179) := previousCrc(19); xorBitMap(2)(180) := previousCrc(20); xorBitMap(2)(181) := previousCrc(21); xorBitMap(2)(183) := previousCrc(23); xorBitMap(2)(185) := previousCrc(25); xorBitMap(2)(186) := previousCrc(26); xorBitMap(2)(187) := previousCrc(27); 
      xorBitMap(3)(60) := currentData(60); xorBitMap(3)(59) := currentData(59); xorBitMap(3)(58) := currentData(58); xorBitMap(3)(56) := currentData(56); xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(160) := previousCrc(0); xorBitMap(3)(161) := previousCrc(1); xorBitMap(3)(164) := previousCrc(4); xorBitMap(3)(165) := previousCrc(5); xorBitMap(3)(166) := previousCrc(6); xorBitMap(3)(167) := previousCrc(7); xorBitMap(3)(168) := previousCrc(8); xorBitMap(3)(173) := previousCrc(13); xorBitMap(3)(180) := previousCrc(20); xorBitMap(3)(181) := previousCrc(21); xorBitMap(3)(182) := previousCrc(22); xorBitMap(3)(184) := previousCrc(24); xorBitMap(3)(186) := previousCrc(26); xorBitMap(3)(187) := previousCrc(27); xorBitMap(3)(188) := previousCrc(28); 
      xorBitMap(4)(63) := currentData(63); xorBitMap(4)(59) := currentData(59); xorBitMap(4)(58) := currentData(58); xorBitMap(4)(57) := currentData(57); xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(161) := previousCrc(1); xorBitMap(4)(166) := previousCrc(6); xorBitMap(4)(167) := previousCrc(7); xorBitMap(4)(168) := previousCrc(8); xorBitMap(4)(169) := previousCrc(9); xorBitMap(4)(172) := previousCrc(12); xorBitMap(4)(173) := previousCrc(13); xorBitMap(4)(174) := previousCrc(14); xorBitMap(4)(175) := previousCrc(15); xorBitMap(4)(176) := previousCrc(16); xorBitMap(4)(178) := previousCrc(18); xorBitMap(4)(185) := previousCrc(25); xorBitMap(4)(186) := previousCrc(26); xorBitMap(4)(187) := previousCrc(27); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(63) := currentData(63); xorBitMap(5)(61) := currentData(61); xorBitMap(5)(59) := currentData(59); xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(165) := previousCrc(5); xorBitMap(5)(167) := previousCrc(7); xorBitMap(5)(168) := previousCrc(8); xorBitMap(5)(169) := previousCrc(9); xorBitMap(5)(170) := previousCrc(10); xorBitMap(5)(172) := previousCrc(12); xorBitMap(5)(174) := previousCrc(14); xorBitMap(5)(177) := previousCrc(17); xorBitMap(5)(178) := previousCrc(18); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(181) := previousCrc(21); xorBitMap(5)(182) := previousCrc(22); xorBitMap(5)(183) := previousCrc(23); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(189) := previousCrc(29); xorBitMap(5)(191) := previousCrc(31); 
      xorBitMap(6)(62) := currentData(62); xorBitMap(6)(60) := currentData(60); xorBitMap(6)(56) := currentData(56); xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(166) := previousCrc(6); xorBitMap(6)(168) := previousCrc(8); xorBitMap(6)(169) := previousCrc(9); xorBitMap(6)(170) := previousCrc(10); xorBitMap(6)(171) := previousCrc(11); xorBitMap(6)(173) := previousCrc(13); xorBitMap(6)(175) := previousCrc(15); xorBitMap(6)(178) := previousCrc(18); xorBitMap(6)(179) := previousCrc(19); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(182) := previousCrc(22); xorBitMap(6)(183) := previousCrc(23); xorBitMap(6)(184) := previousCrc(24); xorBitMap(6)(188) := previousCrc(28); xorBitMap(6)(190) := previousCrc(30); 
      xorBitMap(7)(60) := currentData(60); xorBitMap(7)(58) := currentData(58); xorBitMap(7)(57) := currentData(57); xorBitMap(7)(56) := currentData(56); xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(160) := previousCrc(0); xorBitMap(7)(162) := previousCrc(2); xorBitMap(7)(165) := previousCrc(5); xorBitMap(7)(167) := previousCrc(7); xorBitMap(7)(169) := previousCrc(9); xorBitMap(7)(170) := previousCrc(10); xorBitMap(7)(171) := previousCrc(11); xorBitMap(7)(173) := previousCrc(13); xorBitMap(7)(174) := previousCrc(14); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(178) := previousCrc(18); xorBitMap(7)(179) := previousCrc(19); xorBitMap(7)(180) := previousCrc(20); xorBitMap(7)(182) := previousCrc(22); xorBitMap(7)(184) := previousCrc(24); xorBitMap(7)(185) := previousCrc(25); xorBitMap(7)(186) := previousCrc(26); xorBitMap(7)(188) := previousCrc(28); 
      xorBitMap(8)(63) := currentData(63); xorBitMap(8)(60) := currentData(60); xorBitMap(8)(59) := currentData(59); xorBitMap(8)(57) := currentData(57); xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(160) := previousCrc(0); xorBitMap(8)(161) := previousCrc(1); xorBitMap(8)(162) := previousCrc(2); xorBitMap(8)(163) := previousCrc(3); xorBitMap(8)(165) := previousCrc(5); xorBitMap(8)(166) := previousCrc(6); xorBitMap(8)(168) := previousCrc(8); xorBitMap(8)(170) := previousCrc(10); xorBitMap(8)(171) := previousCrc(11); xorBitMap(8)(173) := previousCrc(13); xorBitMap(8)(174) := previousCrc(14); xorBitMap(8)(178) := previousCrc(18); xorBitMap(8)(179) := previousCrc(19); xorBitMap(8)(180) := previousCrc(20); xorBitMap(8)(182) := previousCrc(22); xorBitMap(8)(185) := previousCrc(25); xorBitMap(8)(187) := previousCrc(27); xorBitMap(8)(188) := previousCrc(28); xorBitMap(8)(191) := previousCrc(31); 
      xorBitMap(9)(61) := currentData(61); xorBitMap(9)(60) := currentData(60); xorBitMap(9)(58) := currentData(58); xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(160) := previousCrc(0); xorBitMap(9)(161) := previousCrc(1); xorBitMap(9)(162) := previousCrc(2); xorBitMap(9)(163) := previousCrc(3); xorBitMap(9)(164) := previousCrc(4); xorBitMap(9)(166) := previousCrc(6); xorBitMap(9)(167) := previousCrc(7); xorBitMap(9)(169) := previousCrc(9); xorBitMap(9)(171) := previousCrc(11); xorBitMap(9)(172) := previousCrc(12); xorBitMap(9)(174) := previousCrc(14); xorBitMap(9)(175) := previousCrc(15); xorBitMap(9)(179) := previousCrc(19); xorBitMap(9)(180) := previousCrc(20); xorBitMap(9)(181) := previousCrc(21); xorBitMap(9)(183) := previousCrc(23); xorBitMap(9)(186) := previousCrc(26); xorBitMap(9)(188) := previousCrc(28); xorBitMap(9)(189) := previousCrc(29); 
      xorBitMap(10)(63) := currentData(63); xorBitMap(10)(62) := currentData(62); xorBitMap(10)(60) := currentData(60); xorBitMap(10)(59) := currentData(59); xorBitMap(10)(58) := currentData(58); xorBitMap(10)(56) := currentData(56); xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(160) := previousCrc(0); xorBitMap(10)(161) := previousCrc(1); xorBitMap(10)(163) := previousCrc(3); xorBitMap(10)(164) := previousCrc(4); xorBitMap(10)(167) := previousCrc(7); xorBitMap(10)(168) := previousCrc(8); xorBitMap(10)(170) := previousCrc(10); xorBitMap(10)(178) := previousCrc(18); xorBitMap(10)(180) := previousCrc(20); xorBitMap(10)(183) := previousCrc(23); xorBitMap(10)(184) := previousCrc(24); xorBitMap(10)(186) := previousCrc(26); xorBitMap(10)(187) := previousCrc(27); xorBitMap(10)(188) := previousCrc(28); xorBitMap(10)(190) := previousCrc(30); xorBitMap(10)(191) := previousCrc(31); 
      xorBitMap(11)(59) := currentData(59); xorBitMap(11)(58) := currentData(58); xorBitMap(11)(57) := currentData(57); xorBitMap(11)(56) := currentData(56); xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(161) := previousCrc(1); xorBitMap(11)(164) := previousCrc(4); xorBitMap(11)(168) := previousCrc(8); xorBitMap(11)(169) := previousCrc(9); xorBitMap(11)(171) := previousCrc(11); xorBitMap(11)(172) := previousCrc(12); xorBitMap(11)(173) := previousCrc(13); xorBitMap(11)(175) := previousCrc(15); xorBitMap(11)(176) := previousCrc(16); xorBitMap(11)(178) := previousCrc(18); xorBitMap(11)(179) := previousCrc(19); xorBitMap(11)(182) := previousCrc(22); xorBitMap(11)(183) := previousCrc(23); xorBitMap(11)(184) := previousCrc(24); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(186) := previousCrc(26); xorBitMap(11)(187) := previousCrc(27); 
      xorBitMap(12)(63) := currentData(63); xorBitMap(12)(61) := currentData(61); xorBitMap(12)(59) := currentData(59); xorBitMap(12)(57) := currentData(57); xorBitMap(12)(56) := currentData(56); xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(169) := previousCrc(9); xorBitMap(12)(170) := previousCrc(10); xorBitMap(12)(174) := previousCrc(14); xorBitMap(12)(175) := previousCrc(15); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(178) := previousCrc(18); xorBitMap(12)(179) := previousCrc(19); xorBitMap(12)(180) := previousCrc(20); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(182) := previousCrc(22); xorBitMap(12)(184) := previousCrc(24); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(187) := previousCrc(27); xorBitMap(12)(189) := previousCrc(29); xorBitMap(12)(191) := previousCrc(31); 
      xorBitMap(13)(62) := currentData(62); xorBitMap(13)(60) := currentData(60); xorBitMap(13)(58) := currentData(58); xorBitMap(13)(57) := currentData(57); xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(160) := previousCrc(0); xorBitMap(13)(170) := previousCrc(10); xorBitMap(13)(171) := previousCrc(11); xorBitMap(13)(175) := previousCrc(15); xorBitMap(13)(176) := previousCrc(16); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(179) := previousCrc(19); xorBitMap(13)(180) := previousCrc(20); xorBitMap(13)(181) := previousCrc(21); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(183) := previousCrc(23); xorBitMap(13)(185) := previousCrc(25); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(188) := previousCrc(28); xorBitMap(13)(190) := previousCrc(30); 
      xorBitMap(14)(63) := currentData(63); xorBitMap(14)(61) := currentData(61); xorBitMap(14)(59) := currentData(59); xorBitMap(14)(58) := currentData(58); xorBitMap(14)(56) := currentData(56); xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(160) := previousCrc(0); xorBitMap(14)(161) := previousCrc(1); xorBitMap(14)(171) := previousCrc(11); xorBitMap(14)(172) := previousCrc(12); xorBitMap(14)(176) := previousCrc(16); xorBitMap(14)(177) := previousCrc(17); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(180) := previousCrc(20); xorBitMap(14)(181) := previousCrc(21); xorBitMap(14)(182) := previousCrc(22); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(184) := previousCrc(24); xorBitMap(14)(186) := previousCrc(26); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(189) := previousCrc(29); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(62) := currentData(62); xorBitMap(15)(60) := currentData(60); xorBitMap(15)(59) := currentData(59); xorBitMap(15)(57) := currentData(57); xorBitMap(15)(56) := currentData(56); xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(161) := previousCrc(1); xorBitMap(15)(162) := previousCrc(2); xorBitMap(15)(172) := previousCrc(12); xorBitMap(15)(173) := previousCrc(13); xorBitMap(15)(177) := previousCrc(17); xorBitMap(15)(178) := previousCrc(18); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(181) := previousCrc(21); xorBitMap(15)(182) := previousCrc(22); xorBitMap(15)(183) := previousCrc(23); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(185) := previousCrc(25); xorBitMap(15)(187) := previousCrc(27); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(190) := previousCrc(30); 
      xorBitMap(16)(57) := currentData(57); xorBitMap(16)(56) := currentData(56); xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(160) := previousCrc(0); xorBitMap(16)(163) := previousCrc(3); xorBitMap(16)(165) := previousCrc(5); xorBitMap(16)(172) := previousCrc(12); xorBitMap(16)(174) := previousCrc(14); xorBitMap(16)(175) := previousCrc(15); xorBitMap(16)(176) := previousCrc(16); xorBitMap(16)(179) := previousCrc(19); xorBitMap(16)(184) := previousCrc(24); xorBitMap(16)(185) := previousCrc(25); 
      xorBitMap(17)(58) := currentData(58); xorBitMap(17)(57) := currentData(57); xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(161) := previousCrc(1); xorBitMap(17)(164) := previousCrc(4); xorBitMap(17)(166) := previousCrc(6); xorBitMap(17)(173) := previousCrc(13); xorBitMap(17)(175) := previousCrc(15); xorBitMap(17)(176) := previousCrc(16); xorBitMap(17)(177) := previousCrc(17); xorBitMap(17)(180) := previousCrc(20); xorBitMap(17)(185) := previousCrc(25); xorBitMap(17)(186) := previousCrc(26); 
      xorBitMap(18)(59) := currentData(59); xorBitMap(18)(58) := currentData(58); xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(160) := previousCrc(0); xorBitMap(18)(162) := previousCrc(2); xorBitMap(18)(165) := previousCrc(5); xorBitMap(18)(167) := previousCrc(7); xorBitMap(18)(174) := previousCrc(14); xorBitMap(18)(176) := previousCrc(16); xorBitMap(18)(177) := previousCrc(17); xorBitMap(18)(178) := previousCrc(18); xorBitMap(18)(181) := previousCrc(21); xorBitMap(18)(186) := previousCrc(26); xorBitMap(18)(187) := previousCrc(27); 
      xorBitMap(19)(60) := currentData(60); xorBitMap(19)(59) := currentData(59); xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(160) := previousCrc(0); xorBitMap(19)(161) := previousCrc(1); xorBitMap(19)(163) := previousCrc(3); xorBitMap(19)(166) := previousCrc(6); xorBitMap(19)(168) := previousCrc(8); xorBitMap(19)(175) := previousCrc(15); xorBitMap(19)(177) := previousCrc(17); xorBitMap(19)(178) := previousCrc(18); xorBitMap(19)(179) := previousCrc(19); xorBitMap(19)(182) := previousCrc(22); xorBitMap(19)(187) := previousCrc(27); xorBitMap(19)(188) := previousCrc(28); 
      xorBitMap(20)(61) := currentData(61); xorBitMap(20)(60) := currentData(60); xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(161) := previousCrc(1); xorBitMap(20)(162) := previousCrc(2); xorBitMap(20)(164) := previousCrc(4); xorBitMap(20)(167) := previousCrc(7); xorBitMap(20)(169) := previousCrc(9); xorBitMap(20)(176) := previousCrc(16); xorBitMap(20)(178) := previousCrc(18); xorBitMap(20)(179) := previousCrc(19); xorBitMap(20)(180) := previousCrc(20); xorBitMap(20)(183) := previousCrc(23); xorBitMap(20)(188) := previousCrc(28); xorBitMap(20)(189) := previousCrc(29); 
      xorBitMap(21)(62) := currentData(62); xorBitMap(21)(61) := currentData(61); xorBitMap(21)(56) := currentData(56); xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(162) := previousCrc(2); xorBitMap(21)(163) := previousCrc(3); xorBitMap(21)(165) := previousCrc(5); xorBitMap(21)(168) := previousCrc(8); xorBitMap(21)(170) := previousCrc(10); xorBitMap(21)(177) := previousCrc(17); xorBitMap(21)(179) := previousCrc(19); xorBitMap(21)(180) := previousCrc(20); xorBitMap(21)(181) := previousCrc(21); xorBitMap(21)(184) := previousCrc(24); xorBitMap(21)(189) := previousCrc(29); xorBitMap(21)(190) := previousCrc(30); 
      xorBitMap(22)(62) := currentData(62); xorBitMap(22)(61) := currentData(61); xorBitMap(22)(60) := currentData(60); xorBitMap(22)(58) := currentData(58); xorBitMap(22)(57) := currentData(57); xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(162) := previousCrc(2); xorBitMap(22)(163) := previousCrc(3); xorBitMap(22)(164) := previousCrc(4); xorBitMap(22)(165) := previousCrc(5); xorBitMap(22)(166) := previousCrc(6); xorBitMap(22)(169) := previousCrc(9); xorBitMap(22)(171) := previousCrc(11); xorBitMap(22)(172) := previousCrc(12); xorBitMap(22)(173) := previousCrc(13); xorBitMap(22)(175) := previousCrc(15); xorBitMap(22)(176) := previousCrc(16); xorBitMap(22)(180) := previousCrc(20); xorBitMap(22)(183) := previousCrc(23); xorBitMap(22)(185) := previousCrc(25); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(188) := previousCrc(28); xorBitMap(22)(189) := previousCrc(29); xorBitMap(22)(190) := previousCrc(30); 
      xorBitMap(23)(62) := currentData(62); xorBitMap(23)(60) := currentData(60); xorBitMap(23)(59) := currentData(59); xorBitMap(23)(56) := currentData(56); xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(162) := previousCrc(2); xorBitMap(23)(163) := previousCrc(3); xorBitMap(23)(164) := previousCrc(4); xorBitMap(23)(166) := previousCrc(6); xorBitMap(23)(167) := previousCrc(7); xorBitMap(23)(170) := previousCrc(10); xorBitMap(23)(174) := previousCrc(14); xorBitMap(23)(175) := previousCrc(15); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(178) := previousCrc(18); xorBitMap(23)(182) := previousCrc(22); xorBitMap(23)(183) := previousCrc(23); xorBitMap(23)(184) := previousCrc(24); xorBitMap(23)(187) := previousCrc(27); xorBitMap(23)(188) := previousCrc(28); xorBitMap(23)(190) := previousCrc(30); 
      xorBitMap(24)(63) := currentData(63); xorBitMap(24)(61) := currentData(61); xorBitMap(24)(60) := currentData(60); xorBitMap(24)(57) := currentData(57); xorBitMap(24)(56) := currentData(56); xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(160) := previousCrc(0); xorBitMap(24)(163) := previousCrc(3); xorBitMap(24)(164) := previousCrc(4); xorBitMap(24)(165) := previousCrc(5); xorBitMap(24)(167) := previousCrc(7); xorBitMap(24)(168) := previousCrc(8); xorBitMap(24)(171) := previousCrc(11); xorBitMap(24)(175) := previousCrc(15); xorBitMap(24)(176) := previousCrc(16); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(179) := previousCrc(19); xorBitMap(24)(183) := previousCrc(23); xorBitMap(24)(184) := previousCrc(24); xorBitMap(24)(185) := previousCrc(25); xorBitMap(24)(188) := previousCrc(28); xorBitMap(24)(189) := previousCrc(29); xorBitMap(24)(191) := previousCrc(31); 
      xorBitMap(25)(62) := currentData(62); xorBitMap(25)(61) := currentData(61); xorBitMap(25)(58) := currentData(58); xorBitMap(25)(57) := currentData(57); xorBitMap(25)(56) := currentData(56); xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(161) := previousCrc(1); xorBitMap(25)(164) := previousCrc(4); xorBitMap(25)(165) := previousCrc(5); xorBitMap(25)(166) := previousCrc(6); xorBitMap(25)(168) := previousCrc(8); xorBitMap(25)(169) := previousCrc(9); xorBitMap(25)(172) := previousCrc(12); xorBitMap(25)(176) := previousCrc(16); xorBitMap(25)(177) := previousCrc(17); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(180) := previousCrc(20); xorBitMap(25)(184) := previousCrc(24); xorBitMap(25)(185) := previousCrc(25); xorBitMap(25)(186) := previousCrc(26); xorBitMap(25)(189) := previousCrc(29); xorBitMap(25)(190) := previousCrc(30); 
      xorBitMap(26)(62) := currentData(62); xorBitMap(26)(61) := currentData(61); xorBitMap(26)(60) := currentData(60); xorBitMap(26)(59) := currentData(59); xorBitMap(26)(57) := currentData(57); xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(166) := previousCrc(6); xorBitMap(26)(167) := previousCrc(7); xorBitMap(26)(169) := previousCrc(9); xorBitMap(26)(170) := previousCrc(10); xorBitMap(26)(172) := previousCrc(12); xorBitMap(26)(175) := previousCrc(15); xorBitMap(26)(176) := previousCrc(16); xorBitMap(26)(177) := previousCrc(17); xorBitMap(26)(180) := previousCrc(20); xorBitMap(26)(182) := previousCrc(22); xorBitMap(26)(183) := previousCrc(23); xorBitMap(26)(185) := previousCrc(25); xorBitMap(26)(187) := previousCrc(27); xorBitMap(26)(188) := previousCrc(28); xorBitMap(26)(189) := previousCrc(29); xorBitMap(26)(190) := previousCrc(30); 
      xorBitMap(27)(63) := currentData(63); xorBitMap(27)(62) := currentData(62); xorBitMap(27)(61) := currentData(61); xorBitMap(27)(60) := currentData(60); xorBitMap(27)(58) := currentData(58); xorBitMap(27)(56) := currentData(56); xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(160) := previousCrc(0); xorBitMap(27)(167) := previousCrc(7); xorBitMap(27)(168) := previousCrc(8); xorBitMap(27)(170) := previousCrc(10); xorBitMap(27)(171) := previousCrc(11); xorBitMap(27)(173) := previousCrc(13); xorBitMap(27)(176) := previousCrc(16); xorBitMap(27)(177) := previousCrc(17); xorBitMap(27)(178) := previousCrc(18); xorBitMap(27)(181) := previousCrc(21); xorBitMap(27)(183) := previousCrc(23); xorBitMap(27)(184) := previousCrc(24); xorBitMap(27)(186) := previousCrc(26); xorBitMap(27)(188) := previousCrc(28); xorBitMap(27)(189) := previousCrc(29); xorBitMap(27)(190) := previousCrc(30); xorBitMap(27)(191) := previousCrc(31); 
      xorBitMap(28)(63) := currentData(63); xorBitMap(28)(62) := currentData(62); xorBitMap(28)(61) := currentData(61); xorBitMap(28)(59) := currentData(59); xorBitMap(28)(57) := currentData(57); xorBitMap(28)(56) := currentData(56); xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(161) := previousCrc(1); xorBitMap(28)(168) := previousCrc(8); xorBitMap(28)(169) := previousCrc(9); xorBitMap(28)(171) := previousCrc(11); xorBitMap(28)(172) := previousCrc(12); xorBitMap(28)(174) := previousCrc(14); xorBitMap(28)(177) := previousCrc(17); xorBitMap(28)(178) := previousCrc(18); xorBitMap(28)(179) := previousCrc(19); xorBitMap(28)(182) := previousCrc(22); xorBitMap(28)(184) := previousCrc(24); xorBitMap(28)(185) := previousCrc(25); xorBitMap(28)(187) := previousCrc(27); xorBitMap(28)(189) := previousCrc(29); xorBitMap(28)(190) := previousCrc(30); xorBitMap(28)(191) := previousCrc(31); 
      xorBitMap(29)(63) := currentData(63); xorBitMap(29)(62) := currentData(62); xorBitMap(29)(60) := currentData(60); xorBitMap(29)(58) := currentData(58); xorBitMap(29)(57) := currentData(57); xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(162) := previousCrc(2); xorBitMap(29)(169) := previousCrc(9); xorBitMap(29)(170) := previousCrc(10); xorBitMap(29)(172) := previousCrc(12); xorBitMap(29)(173) := previousCrc(13); xorBitMap(29)(175) := previousCrc(15); xorBitMap(29)(178) := previousCrc(18); xorBitMap(29)(179) := previousCrc(19); xorBitMap(29)(180) := previousCrc(20); xorBitMap(29)(183) := previousCrc(23); xorBitMap(29)(185) := previousCrc(25); xorBitMap(29)(186) := previousCrc(26); xorBitMap(29)(188) := previousCrc(28); xorBitMap(29)(190) := previousCrc(30); xorBitMap(29)(191) := previousCrc(31); 
      xorBitMap(30)(63) := currentData(63); xorBitMap(30)(61) := currentData(61); xorBitMap(30)(59) := currentData(59); xorBitMap(30)(58) := currentData(58); xorBitMap(30)(56) := currentData(56); xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(160) := previousCrc(0); xorBitMap(30)(163) := previousCrc(3); xorBitMap(30)(170) := previousCrc(10); xorBitMap(30)(171) := previousCrc(11); xorBitMap(30)(173) := previousCrc(13); xorBitMap(30)(174) := previousCrc(14); xorBitMap(30)(176) := previousCrc(16); xorBitMap(30)(179) := previousCrc(19); xorBitMap(30)(180) := previousCrc(20); xorBitMap(30)(181) := previousCrc(21); xorBitMap(30)(184) := previousCrc(24); xorBitMap(30)(186) := previousCrc(26); xorBitMap(30)(187) := previousCrc(27); xorBitMap(30)(189) := previousCrc(29); xorBitMap(30)(191) := previousCrc(31); 
      xorBitMap(31)(62) := currentData(62); xorBitMap(31)(60) := currentData(60); xorBitMap(31)(59) := currentData(59); xorBitMap(31)(57) := currentData(57); xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(161) := previousCrc(1); xorBitMap(31)(164) := previousCrc(4); xorBitMap(31)(171) := previousCrc(11); xorBitMap(31)(172) := previousCrc(12); xorBitMap(31)(174) := previousCrc(14); xorBitMap(31)(175) := previousCrc(15); xorBitMap(31)(177) := previousCrc(17); xorBitMap(31)(180) := previousCrc(20); xorBitMap(31)(181) := previousCrc(21); xorBitMap(31)(182) := previousCrc(22); xorBitMap(31)(185) := previousCrc(25); xorBitMap(31)(187) := previousCrc(27); xorBitMap(31)(188) := previousCrc(28); xorBitMap(31)(190) := previousCrc(30); 
   end procedure;

   procedure xorBitMap9Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(71 downto 0)) is 
   begin
      xorBitMap(0)(68) := currentData(68); xorBitMap(0)(67) := currentData(67); xorBitMap(0)(66) := currentData(66); xorBitMap(0)(65) := currentData(65); xorBitMap(0)(63) := currentData(63); xorBitMap(0)(61) := currentData(61); xorBitMap(0)(60) := currentData(60); xorBitMap(0)(58) := currentData(58); xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(164) := previousCrc(4); xorBitMap(0)(165) := previousCrc(5); xorBitMap(0)(167) := previousCrc(7); xorBitMap(0)(168) := previousCrc(8); xorBitMap(0)(170) := previousCrc(10); xorBitMap(0)(173) := previousCrc(13); xorBitMap(0)(174) := previousCrc(14); xorBitMap(0)(175) := previousCrc(15); xorBitMap(0)(178) := previousCrc(18); xorBitMap(0)(180) := previousCrc(20); xorBitMap(0)(181) := previousCrc(21); xorBitMap(0)(183) := previousCrc(23); xorBitMap(0)(185) := previousCrc(25); xorBitMap(0)(186) := previousCrc(26); xorBitMap(0)(187) := previousCrc(27); xorBitMap(0)(188) := previousCrc(28); 
      xorBitMap(1)(69) := currentData(69); xorBitMap(1)(65) := currentData(65); xorBitMap(1)(64) := currentData(64); xorBitMap(1)(63) := currentData(63); xorBitMap(1)(62) := currentData(62); xorBitMap(1)(60) := currentData(60); xorBitMap(1)(59) := currentData(59); xorBitMap(1)(58) := currentData(58); xorBitMap(1)(56) := currentData(56); xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(164) := previousCrc(4); xorBitMap(1)(166) := previousCrc(6); xorBitMap(1)(167) := previousCrc(7); xorBitMap(1)(169) := previousCrc(9); xorBitMap(1)(170) := previousCrc(10); xorBitMap(1)(171) := previousCrc(11); xorBitMap(1)(173) := previousCrc(13); xorBitMap(1)(176) := previousCrc(16); xorBitMap(1)(178) := previousCrc(18); xorBitMap(1)(179) := previousCrc(19); xorBitMap(1)(180) := previousCrc(20); xorBitMap(1)(182) := previousCrc(22); xorBitMap(1)(183) := previousCrc(23); xorBitMap(1)(184) := previousCrc(24); xorBitMap(1)(185) := previousCrc(25); xorBitMap(1)(189) := previousCrc(29); 
      xorBitMap(2)(70) := currentData(70); xorBitMap(2)(68) := currentData(68); xorBitMap(2)(67) := currentData(67); xorBitMap(2)(64) := currentData(64); xorBitMap(2)(59) := currentData(59); xorBitMap(2)(58) := currentData(58); xorBitMap(2)(57) := currentData(57); xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(164) := previousCrc(4); xorBitMap(2)(171) := previousCrc(11); xorBitMap(2)(172) := previousCrc(12); xorBitMap(2)(173) := previousCrc(13); xorBitMap(2)(175) := previousCrc(15); xorBitMap(2)(177) := previousCrc(17); xorBitMap(2)(178) := previousCrc(18); xorBitMap(2)(179) := previousCrc(19); xorBitMap(2)(184) := previousCrc(24); xorBitMap(2)(187) := previousCrc(27); xorBitMap(2)(188) := previousCrc(28); xorBitMap(2)(190) := previousCrc(30); 
      xorBitMap(3)(71) := currentData(71); xorBitMap(3)(69) := currentData(69); xorBitMap(3)(68) := currentData(68); xorBitMap(3)(65) := currentData(65); xorBitMap(3)(60) := currentData(60); xorBitMap(3)(59) := currentData(59); xorBitMap(3)(58) := currentData(58); xorBitMap(3)(56) := currentData(56); xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(160) := previousCrc(0); xorBitMap(3)(165) := previousCrc(5); xorBitMap(3)(172) := previousCrc(12); xorBitMap(3)(173) := previousCrc(13); xorBitMap(3)(174) := previousCrc(14); xorBitMap(3)(176) := previousCrc(16); xorBitMap(3)(178) := previousCrc(18); xorBitMap(3)(179) := previousCrc(19); xorBitMap(3)(180) := previousCrc(20); xorBitMap(3)(185) := previousCrc(25); xorBitMap(3)(188) := previousCrc(28); xorBitMap(3)(189) := previousCrc(29); xorBitMap(3)(191) := previousCrc(31); 
      xorBitMap(4)(70) := currentData(70); xorBitMap(4)(69) := currentData(69); xorBitMap(4)(68) := currentData(68); xorBitMap(4)(67) := currentData(67); xorBitMap(4)(65) := currentData(65); xorBitMap(4)(63) := currentData(63); xorBitMap(4)(59) := currentData(59); xorBitMap(4)(58) := currentData(58); xorBitMap(4)(57) := currentData(57); xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(160) := previousCrc(0); xorBitMap(4)(161) := previousCrc(1); xorBitMap(4)(164) := previousCrc(4); xorBitMap(4)(165) := previousCrc(5); xorBitMap(4)(166) := previousCrc(6); xorBitMap(4)(167) := previousCrc(7); xorBitMap(4)(168) := previousCrc(8); xorBitMap(4)(170) := previousCrc(10); xorBitMap(4)(177) := previousCrc(17); xorBitMap(4)(178) := previousCrc(18); xorBitMap(4)(179) := previousCrc(19); xorBitMap(4)(183) := previousCrc(23); xorBitMap(4)(185) := previousCrc(25); xorBitMap(4)(187) := previousCrc(27); xorBitMap(4)(188) := previousCrc(28); xorBitMap(4)(189) := previousCrc(29); xorBitMap(4)(190) := previousCrc(30); 
      xorBitMap(5)(71) := currentData(71); xorBitMap(5)(70) := currentData(70); xorBitMap(5)(69) := currentData(69); xorBitMap(5)(67) := currentData(67); xorBitMap(5)(65) := currentData(65); xorBitMap(5)(64) := currentData(64); xorBitMap(5)(63) := currentData(63); xorBitMap(5)(61) := currentData(61); xorBitMap(5)(59) := currentData(59); xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(160) := previousCrc(0); xorBitMap(5)(161) := previousCrc(1); xorBitMap(5)(162) := previousCrc(2); xorBitMap(5)(164) := previousCrc(4); xorBitMap(5)(166) := previousCrc(6); xorBitMap(5)(169) := previousCrc(9); xorBitMap(5)(170) := previousCrc(10); xorBitMap(5)(171) := previousCrc(11); xorBitMap(5)(173) := previousCrc(13); xorBitMap(5)(174) := previousCrc(14); xorBitMap(5)(175) := previousCrc(15); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(181) := previousCrc(21); xorBitMap(5)(183) := previousCrc(23); xorBitMap(5)(184) := previousCrc(24); xorBitMap(5)(185) := previousCrc(25); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(189) := previousCrc(29); xorBitMap(5)(190) := previousCrc(30); xorBitMap(5)(191) := previousCrc(31); 
      xorBitMap(6)(71) := currentData(71); xorBitMap(6)(70) := currentData(70); xorBitMap(6)(68) := currentData(68); xorBitMap(6)(66) := currentData(66); xorBitMap(6)(65) := currentData(65); xorBitMap(6)(64) := currentData(64); xorBitMap(6)(62) := currentData(62); xorBitMap(6)(60) := currentData(60); xorBitMap(6)(56) := currentData(56); xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(160) := previousCrc(0); xorBitMap(6)(161) := previousCrc(1); xorBitMap(6)(162) := previousCrc(2); xorBitMap(6)(163) := previousCrc(3); xorBitMap(6)(165) := previousCrc(5); xorBitMap(6)(167) := previousCrc(7); xorBitMap(6)(170) := previousCrc(10); xorBitMap(6)(171) := previousCrc(11); xorBitMap(6)(172) := previousCrc(12); xorBitMap(6)(174) := previousCrc(14); xorBitMap(6)(175) := previousCrc(15); xorBitMap(6)(176) := previousCrc(16); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(182) := previousCrc(22); xorBitMap(6)(184) := previousCrc(24); xorBitMap(6)(185) := previousCrc(25); xorBitMap(6)(186) := previousCrc(26); xorBitMap(6)(188) := previousCrc(28); xorBitMap(6)(190) := previousCrc(30); xorBitMap(6)(191) := previousCrc(31); 
      xorBitMap(7)(71) := currentData(71); xorBitMap(7)(69) := currentData(69); xorBitMap(7)(68) := currentData(68); xorBitMap(7)(60) := currentData(60); xorBitMap(7)(58) := currentData(58); xorBitMap(7)(57) := currentData(57); xorBitMap(7)(56) := currentData(56); xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(161) := previousCrc(1); xorBitMap(7)(162) := previousCrc(2); xorBitMap(7)(163) := previousCrc(3); xorBitMap(7)(165) := previousCrc(5); xorBitMap(7)(166) := previousCrc(6); xorBitMap(7)(167) := previousCrc(7); xorBitMap(7)(170) := previousCrc(10); xorBitMap(7)(171) := previousCrc(11); xorBitMap(7)(172) := previousCrc(12); xorBitMap(7)(174) := previousCrc(14); xorBitMap(7)(176) := previousCrc(16); xorBitMap(7)(177) := previousCrc(17); xorBitMap(7)(178) := previousCrc(18); xorBitMap(7)(180) := previousCrc(20); xorBitMap(7)(188) := previousCrc(28); xorBitMap(7)(189) := previousCrc(29); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(70) := currentData(70); xorBitMap(8)(69) := currentData(69); xorBitMap(8)(68) := currentData(68); xorBitMap(8)(67) := currentData(67); xorBitMap(8)(66) := currentData(66); xorBitMap(8)(65) := currentData(65); xorBitMap(8)(63) := currentData(63); xorBitMap(8)(60) := currentData(60); xorBitMap(8)(59) := currentData(59); xorBitMap(8)(57) := currentData(57); xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(160) := previousCrc(0); xorBitMap(8)(162) := previousCrc(2); xorBitMap(8)(163) := previousCrc(3); xorBitMap(8)(165) := previousCrc(5); xorBitMap(8)(166) := previousCrc(6); xorBitMap(8)(170) := previousCrc(10); xorBitMap(8)(171) := previousCrc(11); xorBitMap(8)(172) := previousCrc(12); xorBitMap(8)(174) := previousCrc(14); xorBitMap(8)(177) := previousCrc(17); xorBitMap(8)(179) := previousCrc(19); xorBitMap(8)(180) := previousCrc(20); xorBitMap(8)(183) := previousCrc(23); xorBitMap(8)(185) := previousCrc(25); xorBitMap(8)(186) := previousCrc(26); xorBitMap(8)(187) := previousCrc(27); xorBitMap(8)(188) := previousCrc(28); xorBitMap(8)(189) := previousCrc(29); xorBitMap(8)(190) := previousCrc(30); 
      xorBitMap(9)(71) := currentData(71); xorBitMap(9)(70) := currentData(70); xorBitMap(9)(69) := currentData(69); xorBitMap(9)(68) := currentData(68); xorBitMap(9)(67) := currentData(67); xorBitMap(9)(66) := currentData(66); xorBitMap(9)(64) := currentData(64); xorBitMap(9)(61) := currentData(61); xorBitMap(9)(60) := currentData(60); xorBitMap(9)(58) := currentData(58); xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(161) := previousCrc(1); xorBitMap(9)(163) := previousCrc(3); xorBitMap(9)(164) := previousCrc(4); xorBitMap(9)(166) := previousCrc(6); xorBitMap(9)(167) := previousCrc(7); xorBitMap(9)(171) := previousCrc(11); xorBitMap(9)(172) := previousCrc(12); xorBitMap(9)(173) := previousCrc(13); xorBitMap(9)(175) := previousCrc(15); xorBitMap(9)(178) := previousCrc(18); xorBitMap(9)(180) := previousCrc(20); xorBitMap(9)(181) := previousCrc(21); xorBitMap(9)(184) := previousCrc(24); xorBitMap(9)(186) := previousCrc(26); xorBitMap(9)(187) := previousCrc(27); xorBitMap(9)(188) := previousCrc(28); xorBitMap(9)(189) := previousCrc(29); xorBitMap(9)(190) := previousCrc(30); xorBitMap(9)(191) := previousCrc(31); 
      xorBitMap(10)(71) := currentData(71); xorBitMap(10)(70) := currentData(70); xorBitMap(10)(69) := currentData(69); xorBitMap(10)(66) := currentData(66); xorBitMap(10)(63) := currentData(63); xorBitMap(10)(62) := currentData(62); xorBitMap(10)(60) := currentData(60); xorBitMap(10)(59) := currentData(59); xorBitMap(10)(58) := currentData(58); xorBitMap(10)(56) := currentData(56); xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(160) := previousCrc(0); xorBitMap(10)(162) := previousCrc(2); xorBitMap(10)(170) := previousCrc(10); xorBitMap(10)(172) := previousCrc(12); xorBitMap(10)(175) := previousCrc(15); xorBitMap(10)(176) := previousCrc(16); xorBitMap(10)(178) := previousCrc(18); xorBitMap(10)(179) := previousCrc(19); xorBitMap(10)(180) := previousCrc(20); xorBitMap(10)(182) := previousCrc(22); xorBitMap(10)(183) := previousCrc(23); xorBitMap(10)(186) := previousCrc(26); xorBitMap(10)(189) := previousCrc(29); xorBitMap(10)(190) := previousCrc(30); xorBitMap(10)(191) := previousCrc(31); 
      xorBitMap(11)(71) := currentData(71); xorBitMap(11)(70) := currentData(70); xorBitMap(11)(68) := currentData(68); xorBitMap(11)(66) := currentData(66); xorBitMap(11)(65) := currentData(65); xorBitMap(11)(64) := currentData(64); xorBitMap(11)(59) := currentData(59); xorBitMap(11)(58) := currentData(58); xorBitMap(11)(57) := currentData(57); xorBitMap(11)(56) := currentData(56); xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(160) := previousCrc(0); xorBitMap(11)(161) := previousCrc(1); xorBitMap(11)(163) := previousCrc(3); xorBitMap(11)(164) := previousCrc(4); xorBitMap(11)(165) := previousCrc(5); xorBitMap(11)(167) := previousCrc(7); xorBitMap(11)(168) := previousCrc(8); xorBitMap(11)(170) := previousCrc(10); xorBitMap(11)(171) := previousCrc(11); xorBitMap(11)(174) := previousCrc(14); xorBitMap(11)(175) := previousCrc(15); xorBitMap(11)(176) := previousCrc(16); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(178) := previousCrc(18); xorBitMap(11)(179) := previousCrc(19); xorBitMap(11)(184) := previousCrc(24); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(186) := previousCrc(26); xorBitMap(11)(188) := previousCrc(28); xorBitMap(11)(190) := previousCrc(30); xorBitMap(11)(191) := previousCrc(31); 
      xorBitMap(12)(71) := currentData(71); xorBitMap(12)(69) := currentData(69); xorBitMap(12)(68) := currentData(68); xorBitMap(12)(63) := currentData(63); xorBitMap(12)(61) := currentData(61); xorBitMap(12)(59) := currentData(59); xorBitMap(12)(57) := currentData(57); xorBitMap(12)(56) := currentData(56); xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(161) := previousCrc(1); xorBitMap(12)(162) := previousCrc(2); xorBitMap(12)(166) := previousCrc(6); xorBitMap(12)(167) := previousCrc(7); xorBitMap(12)(169) := previousCrc(9); xorBitMap(12)(170) := previousCrc(10); xorBitMap(12)(171) := previousCrc(11); xorBitMap(12)(172) := previousCrc(12); xorBitMap(12)(173) := previousCrc(13); xorBitMap(12)(174) := previousCrc(14); xorBitMap(12)(176) := previousCrc(16); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(179) := previousCrc(19); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(183) := previousCrc(23); xorBitMap(12)(188) := previousCrc(28); xorBitMap(12)(189) := previousCrc(29); xorBitMap(12)(191) := previousCrc(31); 
      xorBitMap(13)(70) := currentData(70); xorBitMap(13)(69) := currentData(69); xorBitMap(13)(64) := currentData(64); xorBitMap(13)(62) := currentData(62); xorBitMap(13)(60) := currentData(60); xorBitMap(13)(58) := currentData(58); xorBitMap(13)(57) := currentData(57); xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(162) := previousCrc(2); xorBitMap(13)(163) := previousCrc(3); xorBitMap(13)(167) := previousCrc(7); xorBitMap(13)(168) := previousCrc(8); xorBitMap(13)(170) := previousCrc(10); xorBitMap(13)(171) := previousCrc(11); xorBitMap(13)(172) := previousCrc(12); xorBitMap(13)(173) := previousCrc(13); xorBitMap(13)(174) := previousCrc(14); xorBitMap(13)(175) := previousCrc(15); xorBitMap(13)(177) := previousCrc(17); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(180) := previousCrc(20); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(184) := previousCrc(24); xorBitMap(13)(189) := previousCrc(29); xorBitMap(13)(190) := previousCrc(30); 
      xorBitMap(14)(71) := currentData(71); xorBitMap(14)(70) := currentData(70); xorBitMap(14)(65) := currentData(65); xorBitMap(14)(63) := currentData(63); xorBitMap(14)(61) := currentData(61); xorBitMap(14)(59) := currentData(59); xorBitMap(14)(58) := currentData(58); xorBitMap(14)(56) := currentData(56); xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(163) := previousCrc(3); xorBitMap(14)(164) := previousCrc(4); xorBitMap(14)(168) := previousCrc(8); xorBitMap(14)(169) := previousCrc(9); xorBitMap(14)(171) := previousCrc(11); xorBitMap(14)(172) := previousCrc(12); xorBitMap(14)(173) := previousCrc(13); xorBitMap(14)(174) := previousCrc(14); xorBitMap(14)(175) := previousCrc(15); xorBitMap(14)(176) := previousCrc(16); xorBitMap(14)(178) := previousCrc(18); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(181) := previousCrc(21); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(185) := previousCrc(25); xorBitMap(14)(190) := previousCrc(30); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(71) := currentData(71); xorBitMap(15)(66) := currentData(66); xorBitMap(15)(64) := currentData(64); xorBitMap(15)(62) := currentData(62); xorBitMap(15)(60) := currentData(60); xorBitMap(15)(59) := currentData(59); xorBitMap(15)(57) := currentData(57); xorBitMap(15)(56) := currentData(56); xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(164) := previousCrc(4); xorBitMap(15)(165) := previousCrc(5); xorBitMap(15)(169) := previousCrc(9); xorBitMap(15)(170) := previousCrc(10); xorBitMap(15)(172) := previousCrc(12); xorBitMap(15)(173) := previousCrc(13); xorBitMap(15)(174) := previousCrc(14); xorBitMap(15)(175) := previousCrc(15); xorBitMap(15)(176) := previousCrc(16); xorBitMap(15)(177) := previousCrc(17); xorBitMap(15)(179) := previousCrc(19); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(182) := previousCrc(22); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(186) := previousCrc(26); xorBitMap(15)(191) := previousCrc(31); 
      xorBitMap(16)(68) := currentData(68); xorBitMap(16)(66) := currentData(66); xorBitMap(16)(57) := currentData(57); xorBitMap(16)(56) := currentData(56); xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(164) := previousCrc(4); xorBitMap(16)(166) := previousCrc(6); xorBitMap(16)(167) := previousCrc(7); xorBitMap(16)(168) := previousCrc(8); xorBitMap(16)(171) := previousCrc(11); xorBitMap(16)(176) := previousCrc(16); xorBitMap(16)(177) := previousCrc(17); xorBitMap(16)(186) := previousCrc(26); xorBitMap(16)(188) := previousCrc(28); 
      xorBitMap(17)(69) := currentData(69); xorBitMap(17)(67) := currentData(67); xorBitMap(17)(58) := currentData(58); xorBitMap(17)(57) := currentData(57); xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(165) := previousCrc(5); xorBitMap(17)(167) := previousCrc(7); xorBitMap(17)(168) := previousCrc(8); xorBitMap(17)(169) := previousCrc(9); xorBitMap(17)(172) := previousCrc(12); xorBitMap(17)(177) := previousCrc(17); xorBitMap(17)(178) := previousCrc(18); xorBitMap(17)(187) := previousCrc(27); xorBitMap(17)(189) := previousCrc(29); 
      xorBitMap(18)(70) := currentData(70); xorBitMap(18)(68) := currentData(68); xorBitMap(18)(59) := currentData(59); xorBitMap(18)(58) := currentData(58); xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(166) := previousCrc(6); xorBitMap(18)(168) := previousCrc(8); xorBitMap(18)(169) := previousCrc(9); xorBitMap(18)(170) := previousCrc(10); xorBitMap(18)(173) := previousCrc(13); xorBitMap(18)(178) := previousCrc(18); xorBitMap(18)(179) := previousCrc(19); xorBitMap(18)(188) := previousCrc(28); xorBitMap(18)(190) := previousCrc(30); 
      xorBitMap(19)(71) := currentData(71); xorBitMap(19)(69) := currentData(69); xorBitMap(19)(60) := currentData(60); xorBitMap(19)(59) := currentData(59); xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(160) := previousCrc(0); xorBitMap(19)(167) := previousCrc(7); xorBitMap(19)(169) := previousCrc(9); xorBitMap(19)(170) := previousCrc(10); xorBitMap(19)(171) := previousCrc(11); xorBitMap(19)(174) := previousCrc(14); xorBitMap(19)(179) := previousCrc(19); xorBitMap(19)(180) := previousCrc(20); xorBitMap(19)(189) := previousCrc(29); xorBitMap(19)(191) := previousCrc(31); 
      xorBitMap(20)(70) := currentData(70); xorBitMap(20)(61) := currentData(61); xorBitMap(20)(60) := currentData(60); xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(161) := previousCrc(1); xorBitMap(20)(168) := previousCrc(8); xorBitMap(20)(170) := previousCrc(10); xorBitMap(20)(171) := previousCrc(11); xorBitMap(20)(172) := previousCrc(12); xorBitMap(20)(175) := previousCrc(15); xorBitMap(20)(180) := previousCrc(20); xorBitMap(20)(181) := previousCrc(21); xorBitMap(20)(190) := previousCrc(30); 
      xorBitMap(21)(71) := currentData(71); xorBitMap(21)(62) := currentData(62); xorBitMap(21)(61) := currentData(61); xorBitMap(21)(56) := currentData(56); xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(160) := previousCrc(0); xorBitMap(21)(162) := previousCrc(2); xorBitMap(21)(169) := previousCrc(9); xorBitMap(21)(171) := previousCrc(11); xorBitMap(21)(172) := previousCrc(12); xorBitMap(21)(173) := previousCrc(13); xorBitMap(21)(176) := previousCrc(16); xorBitMap(21)(181) := previousCrc(21); xorBitMap(21)(182) := previousCrc(22); xorBitMap(21)(191) := previousCrc(31); 
      xorBitMap(22)(68) := currentData(68); xorBitMap(22)(67) := currentData(67); xorBitMap(22)(66) := currentData(66); xorBitMap(22)(65) := currentData(65); xorBitMap(22)(62) := currentData(62); xorBitMap(22)(61) := currentData(61); xorBitMap(22)(60) := currentData(60); xorBitMap(22)(58) := currentData(58); xorBitMap(22)(57) := currentData(57); xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(161) := previousCrc(1); xorBitMap(22)(163) := previousCrc(3); xorBitMap(22)(164) := previousCrc(4); xorBitMap(22)(165) := previousCrc(5); xorBitMap(22)(167) := previousCrc(7); xorBitMap(22)(168) := previousCrc(8); xorBitMap(22)(172) := previousCrc(12); xorBitMap(22)(175) := previousCrc(15); xorBitMap(22)(177) := previousCrc(17); xorBitMap(22)(178) := previousCrc(18); xorBitMap(22)(180) := previousCrc(20); xorBitMap(22)(181) := previousCrc(21); xorBitMap(22)(182) := previousCrc(22); xorBitMap(22)(185) := previousCrc(25); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(187) := previousCrc(27); xorBitMap(22)(188) := previousCrc(28); 
      xorBitMap(23)(69) := currentData(69); xorBitMap(23)(65) := currentData(65); xorBitMap(23)(62) := currentData(62); xorBitMap(23)(60) := currentData(60); xorBitMap(23)(59) := currentData(59); xorBitMap(23)(56) := currentData(56); xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(162) := previousCrc(2); xorBitMap(23)(166) := previousCrc(6); xorBitMap(23)(167) := previousCrc(7); xorBitMap(23)(169) := previousCrc(9); xorBitMap(23)(170) := previousCrc(10); xorBitMap(23)(174) := previousCrc(14); xorBitMap(23)(175) := previousCrc(15); xorBitMap(23)(176) := previousCrc(16); xorBitMap(23)(179) := previousCrc(19); xorBitMap(23)(180) := previousCrc(20); xorBitMap(23)(182) := previousCrc(22); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(189) := previousCrc(29); 
      xorBitMap(24)(70) := currentData(70); xorBitMap(24)(66) := currentData(66); xorBitMap(24)(63) := currentData(63); xorBitMap(24)(61) := currentData(61); xorBitMap(24)(60) := currentData(60); xorBitMap(24)(57) := currentData(57); xorBitMap(24)(56) := currentData(56); xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(160) := previousCrc(0); xorBitMap(24)(163) := previousCrc(3); xorBitMap(24)(167) := previousCrc(7); xorBitMap(24)(168) := previousCrc(8); xorBitMap(24)(170) := previousCrc(10); xorBitMap(24)(171) := previousCrc(11); xorBitMap(24)(175) := previousCrc(15); xorBitMap(24)(176) := previousCrc(16); xorBitMap(24)(177) := previousCrc(17); xorBitMap(24)(180) := previousCrc(20); xorBitMap(24)(181) := previousCrc(21); xorBitMap(24)(183) := previousCrc(23); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(190) := previousCrc(30); 
      xorBitMap(25)(71) := currentData(71); xorBitMap(25)(67) := currentData(67); xorBitMap(25)(64) := currentData(64); xorBitMap(25)(62) := currentData(62); xorBitMap(25)(61) := currentData(61); xorBitMap(25)(58) := currentData(58); xorBitMap(25)(57) := currentData(57); xorBitMap(25)(56) := currentData(56); xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(160) := previousCrc(0); xorBitMap(25)(161) := previousCrc(1); xorBitMap(25)(164) := previousCrc(4); xorBitMap(25)(168) := previousCrc(8); xorBitMap(25)(169) := previousCrc(9); xorBitMap(25)(171) := previousCrc(11); xorBitMap(25)(172) := previousCrc(12); xorBitMap(25)(176) := previousCrc(16); xorBitMap(25)(177) := previousCrc(17); xorBitMap(25)(178) := previousCrc(18); xorBitMap(25)(181) := previousCrc(21); xorBitMap(25)(182) := previousCrc(22); xorBitMap(25)(184) := previousCrc(24); xorBitMap(25)(187) := previousCrc(27); xorBitMap(25)(191) := previousCrc(31); 
      xorBitMap(26)(67) := currentData(67); xorBitMap(26)(66) := currentData(66); xorBitMap(26)(62) := currentData(62); xorBitMap(26)(61) := currentData(61); xorBitMap(26)(60) := currentData(60); xorBitMap(26)(59) := currentData(59); xorBitMap(26)(57) := currentData(57); xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(161) := previousCrc(1); xorBitMap(26)(162) := previousCrc(2); xorBitMap(26)(164) := previousCrc(4); xorBitMap(26)(167) := previousCrc(7); xorBitMap(26)(168) := previousCrc(8); xorBitMap(26)(169) := previousCrc(9); xorBitMap(26)(172) := previousCrc(12); xorBitMap(26)(174) := previousCrc(14); xorBitMap(26)(175) := previousCrc(15); xorBitMap(26)(177) := previousCrc(17); xorBitMap(26)(179) := previousCrc(19); xorBitMap(26)(180) := previousCrc(20); xorBitMap(26)(181) := previousCrc(21); xorBitMap(26)(182) := previousCrc(22); xorBitMap(26)(186) := previousCrc(26); xorBitMap(26)(187) := previousCrc(27); 
      xorBitMap(27)(68) := currentData(68); xorBitMap(27)(67) := currentData(67); xorBitMap(27)(63) := currentData(63); xorBitMap(27)(62) := currentData(62); xorBitMap(27)(61) := currentData(61); xorBitMap(27)(60) := currentData(60); xorBitMap(27)(58) := currentData(58); xorBitMap(27)(56) := currentData(56); xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(160) := previousCrc(0); xorBitMap(27)(162) := previousCrc(2); xorBitMap(27)(163) := previousCrc(3); xorBitMap(27)(165) := previousCrc(5); xorBitMap(27)(168) := previousCrc(8); xorBitMap(27)(169) := previousCrc(9); xorBitMap(27)(170) := previousCrc(10); xorBitMap(27)(173) := previousCrc(13); xorBitMap(27)(175) := previousCrc(15); xorBitMap(27)(176) := previousCrc(16); xorBitMap(27)(178) := previousCrc(18); xorBitMap(27)(180) := previousCrc(20); xorBitMap(27)(181) := previousCrc(21); xorBitMap(27)(182) := previousCrc(22); xorBitMap(27)(183) := previousCrc(23); xorBitMap(27)(187) := previousCrc(27); xorBitMap(27)(188) := previousCrc(28); 
      xorBitMap(28)(69) := currentData(69); xorBitMap(28)(68) := currentData(68); xorBitMap(28)(64) := currentData(64); xorBitMap(28)(63) := currentData(63); xorBitMap(28)(62) := currentData(62); xorBitMap(28)(61) := currentData(61); xorBitMap(28)(59) := currentData(59); xorBitMap(28)(57) := currentData(57); xorBitMap(28)(56) := currentData(56); xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(160) := previousCrc(0); xorBitMap(28)(161) := previousCrc(1); xorBitMap(28)(163) := previousCrc(3); xorBitMap(28)(164) := previousCrc(4); xorBitMap(28)(166) := previousCrc(6); xorBitMap(28)(169) := previousCrc(9); xorBitMap(28)(170) := previousCrc(10); xorBitMap(28)(171) := previousCrc(11); xorBitMap(28)(174) := previousCrc(14); xorBitMap(28)(176) := previousCrc(16); xorBitMap(28)(177) := previousCrc(17); xorBitMap(28)(179) := previousCrc(19); xorBitMap(28)(181) := previousCrc(21); xorBitMap(28)(182) := previousCrc(22); xorBitMap(28)(183) := previousCrc(23); xorBitMap(28)(184) := previousCrc(24); xorBitMap(28)(188) := previousCrc(28); xorBitMap(28)(189) := previousCrc(29); 
      xorBitMap(29)(70) := currentData(70); xorBitMap(29)(69) := currentData(69); xorBitMap(29)(65) := currentData(65); xorBitMap(29)(64) := currentData(64); xorBitMap(29)(63) := currentData(63); xorBitMap(29)(62) := currentData(62); xorBitMap(29)(60) := currentData(60); xorBitMap(29)(58) := currentData(58); xorBitMap(29)(57) := currentData(57); xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(161) := previousCrc(1); xorBitMap(29)(162) := previousCrc(2); xorBitMap(29)(164) := previousCrc(4); xorBitMap(29)(165) := previousCrc(5); xorBitMap(29)(167) := previousCrc(7); xorBitMap(29)(170) := previousCrc(10); xorBitMap(29)(171) := previousCrc(11); xorBitMap(29)(172) := previousCrc(12); xorBitMap(29)(175) := previousCrc(15); xorBitMap(29)(177) := previousCrc(17); xorBitMap(29)(178) := previousCrc(18); xorBitMap(29)(180) := previousCrc(20); xorBitMap(29)(182) := previousCrc(22); xorBitMap(29)(183) := previousCrc(23); xorBitMap(29)(184) := previousCrc(24); xorBitMap(29)(185) := previousCrc(25); xorBitMap(29)(189) := previousCrc(29); xorBitMap(29)(190) := previousCrc(30); 
      xorBitMap(30)(71) := currentData(71); xorBitMap(30)(70) := currentData(70); xorBitMap(30)(66) := currentData(66); xorBitMap(30)(65) := currentData(65); xorBitMap(30)(64) := currentData(64); xorBitMap(30)(63) := currentData(63); xorBitMap(30)(61) := currentData(61); xorBitMap(30)(59) := currentData(59); xorBitMap(30)(58) := currentData(58); xorBitMap(30)(56) := currentData(56); xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(162) := previousCrc(2); xorBitMap(30)(163) := previousCrc(3); xorBitMap(30)(165) := previousCrc(5); xorBitMap(30)(166) := previousCrc(6); xorBitMap(30)(168) := previousCrc(8); xorBitMap(30)(171) := previousCrc(11); xorBitMap(30)(172) := previousCrc(12); xorBitMap(30)(173) := previousCrc(13); xorBitMap(30)(176) := previousCrc(16); xorBitMap(30)(178) := previousCrc(18); xorBitMap(30)(179) := previousCrc(19); xorBitMap(30)(181) := previousCrc(21); xorBitMap(30)(183) := previousCrc(23); xorBitMap(30)(184) := previousCrc(24); xorBitMap(30)(185) := previousCrc(25); xorBitMap(30)(186) := previousCrc(26); xorBitMap(30)(190) := previousCrc(30); xorBitMap(30)(191) := previousCrc(31); 
      xorBitMap(31)(71) := currentData(71); xorBitMap(31)(67) := currentData(67); xorBitMap(31)(66) := currentData(66); xorBitMap(31)(65) := currentData(65); xorBitMap(31)(64) := currentData(64); xorBitMap(31)(62) := currentData(62); xorBitMap(31)(60) := currentData(60); xorBitMap(31)(59) := currentData(59); xorBitMap(31)(57) := currentData(57); xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(163) := previousCrc(3); xorBitMap(31)(164) := previousCrc(4); xorBitMap(31)(166) := previousCrc(6); xorBitMap(31)(167) := previousCrc(7); xorBitMap(31)(169) := previousCrc(9); xorBitMap(31)(172) := previousCrc(12); xorBitMap(31)(173) := previousCrc(13); xorBitMap(31)(174) := previousCrc(14); xorBitMap(31)(177) := previousCrc(17); xorBitMap(31)(179) := previousCrc(19); xorBitMap(31)(180) := previousCrc(20); xorBitMap(31)(182) := previousCrc(22); xorBitMap(31)(184) := previousCrc(24); xorBitMap(31)(185) := previousCrc(25); xorBitMap(31)(186) := previousCrc(26); xorBitMap(31)(187) := previousCrc(27); xorBitMap(31)(191) := previousCrc(31); 
   end procedure;

   procedure xorBitMap10Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(79 downto 0)) is 
   begin
      xorBitMap(0)(79) := currentData(79); xorBitMap(0)(73) := currentData(73); xorBitMap(0)(72) := currentData(72); xorBitMap(0)(68) := currentData(68); xorBitMap(0)(67) := currentData(67); xorBitMap(0)(66) := currentData(66); xorBitMap(0)(65) := currentData(65); xorBitMap(0)(63) := currentData(63); xorBitMap(0)(61) := currentData(61); xorBitMap(0)(60) := currentData(60); xorBitMap(0)(58) := currentData(58); xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(160) := previousCrc(0); xorBitMap(0)(162) := previousCrc(2); xorBitMap(0)(165) := previousCrc(5); xorBitMap(0)(166) := previousCrc(6); xorBitMap(0)(167) := previousCrc(7); xorBitMap(0)(170) := previousCrc(10); xorBitMap(0)(172) := previousCrc(12); xorBitMap(0)(173) := previousCrc(13); xorBitMap(0)(175) := previousCrc(15); xorBitMap(0)(177) := previousCrc(17); xorBitMap(0)(178) := previousCrc(18); xorBitMap(0)(179) := previousCrc(19); xorBitMap(0)(180) := previousCrc(20); xorBitMap(0)(184) := previousCrc(24); xorBitMap(0)(185) := previousCrc(25); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(79) := currentData(79); xorBitMap(1)(74) := currentData(74); xorBitMap(1)(72) := currentData(72); xorBitMap(1)(69) := currentData(69); xorBitMap(1)(65) := currentData(65); xorBitMap(1)(64) := currentData(64); xorBitMap(1)(63) := currentData(63); xorBitMap(1)(62) := currentData(62); xorBitMap(1)(60) := currentData(60); xorBitMap(1)(59) := currentData(59); xorBitMap(1)(58) := currentData(58); xorBitMap(1)(56) := currentData(56); xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(161) := previousCrc(1); xorBitMap(1)(162) := previousCrc(2); xorBitMap(1)(163) := previousCrc(3); xorBitMap(1)(165) := previousCrc(5); xorBitMap(1)(168) := previousCrc(8); xorBitMap(1)(170) := previousCrc(10); xorBitMap(1)(171) := previousCrc(11); xorBitMap(1)(172) := previousCrc(12); xorBitMap(1)(174) := previousCrc(14); xorBitMap(1)(175) := previousCrc(15); xorBitMap(1)(176) := previousCrc(16); xorBitMap(1)(177) := previousCrc(17); xorBitMap(1)(181) := previousCrc(21); xorBitMap(1)(184) := previousCrc(24); xorBitMap(1)(186) := previousCrc(26); xorBitMap(1)(191) := previousCrc(31); 
      xorBitMap(2)(79) := currentData(79); xorBitMap(2)(75) := currentData(75); xorBitMap(2)(72) := currentData(72); xorBitMap(2)(70) := currentData(70); xorBitMap(2)(68) := currentData(68); xorBitMap(2)(67) := currentData(67); xorBitMap(2)(64) := currentData(64); xorBitMap(2)(59) := currentData(59); xorBitMap(2)(58) := currentData(58); xorBitMap(2)(57) := currentData(57); xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(163) := previousCrc(3); xorBitMap(2)(164) := previousCrc(4); xorBitMap(2)(165) := previousCrc(5); xorBitMap(2)(167) := previousCrc(7); xorBitMap(2)(169) := previousCrc(9); xorBitMap(2)(170) := previousCrc(10); xorBitMap(2)(171) := previousCrc(11); xorBitMap(2)(176) := previousCrc(16); xorBitMap(2)(179) := previousCrc(19); xorBitMap(2)(180) := previousCrc(20); xorBitMap(2)(182) := previousCrc(22); xorBitMap(2)(184) := previousCrc(24); xorBitMap(2)(187) := previousCrc(27); xorBitMap(2)(191) := previousCrc(31); 
      xorBitMap(3)(76) := currentData(76); xorBitMap(3)(73) := currentData(73); xorBitMap(3)(71) := currentData(71); xorBitMap(3)(69) := currentData(69); xorBitMap(3)(68) := currentData(68); xorBitMap(3)(65) := currentData(65); xorBitMap(3)(60) := currentData(60); xorBitMap(3)(59) := currentData(59); xorBitMap(3)(58) := currentData(58); xorBitMap(3)(56) := currentData(56); xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(164) := previousCrc(4); xorBitMap(3)(165) := previousCrc(5); xorBitMap(3)(166) := previousCrc(6); xorBitMap(3)(168) := previousCrc(8); xorBitMap(3)(170) := previousCrc(10); xorBitMap(3)(171) := previousCrc(11); xorBitMap(3)(172) := previousCrc(12); xorBitMap(3)(177) := previousCrc(17); xorBitMap(3)(180) := previousCrc(20); xorBitMap(3)(181) := previousCrc(21); xorBitMap(3)(183) := previousCrc(23); xorBitMap(3)(185) := previousCrc(25); xorBitMap(3)(188) := previousCrc(28); 
      xorBitMap(4)(79) := currentData(79); xorBitMap(4)(77) := currentData(77); xorBitMap(4)(74) := currentData(74); xorBitMap(4)(73) := currentData(73); xorBitMap(4)(70) := currentData(70); xorBitMap(4)(69) := currentData(69); xorBitMap(4)(68) := currentData(68); xorBitMap(4)(67) := currentData(67); xorBitMap(4)(65) := currentData(65); xorBitMap(4)(63) := currentData(63); xorBitMap(4)(59) := currentData(59); xorBitMap(4)(58) := currentData(58); xorBitMap(4)(57) := currentData(57); xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(160) := previousCrc(0); xorBitMap(4)(162) := previousCrc(2); xorBitMap(4)(169) := previousCrc(9); xorBitMap(4)(170) := previousCrc(10); xorBitMap(4)(171) := previousCrc(11); xorBitMap(4)(175) := previousCrc(15); xorBitMap(4)(177) := previousCrc(17); xorBitMap(4)(179) := previousCrc(19); xorBitMap(4)(180) := previousCrc(20); xorBitMap(4)(181) := previousCrc(21); xorBitMap(4)(182) := previousCrc(22); xorBitMap(4)(185) := previousCrc(25); xorBitMap(4)(186) := previousCrc(26); xorBitMap(4)(189) := previousCrc(29); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(79) := currentData(79); xorBitMap(5)(78) := currentData(78); xorBitMap(5)(75) := currentData(75); xorBitMap(5)(74) := currentData(74); xorBitMap(5)(73) := currentData(73); xorBitMap(5)(72) := currentData(72); xorBitMap(5)(71) := currentData(71); xorBitMap(5)(70) := currentData(70); xorBitMap(5)(69) := currentData(69); xorBitMap(5)(67) := currentData(67); xorBitMap(5)(65) := currentData(65); xorBitMap(5)(64) := currentData(64); xorBitMap(5)(63) := currentData(63); xorBitMap(5)(61) := currentData(61); xorBitMap(5)(59) := currentData(59); xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(161) := previousCrc(1); xorBitMap(5)(162) := previousCrc(2); xorBitMap(5)(163) := previousCrc(3); xorBitMap(5)(165) := previousCrc(5); xorBitMap(5)(166) := previousCrc(6); xorBitMap(5)(167) := previousCrc(7); xorBitMap(5)(171) := previousCrc(11); xorBitMap(5)(173) := previousCrc(13); xorBitMap(5)(175) := previousCrc(15); xorBitMap(5)(176) := previousCrc(16); xorBitMap(5)(177) := previousCrc(17); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(181) := previousCrc(21); xorBitMap(5)(182) := previousCrc(22); xorBitMap(5)(183) := previousCrc(23); xorBitMap(5)(184) := previousCrc(24); xorBitMap(5)(185) := previousCrc(25); xorBitMap(5)(186) := previousCrc(26); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(190) := previousCrc(30); xorBitMap(5)(191) := previousCrc(31); 
      xorBitMap(6)(79) := currentData(79); xorBitMap(6)(76) := currentData(76); xorBitMap(6)(75) := currentData(75); xorBitMap(6)(74) := currentData(74); xorBitMap(6)(73) := currentData(73); xorBitMap(6)(72) := currentData(72); xorBitMap(6)(71) := currentData(71); xorBitMap(6)(70) := currentData(70); xorBitMap(6)(68) := currentData(68); xorBitMap(6)(66) := currentData(66); xorBitMap(6)(65) := currentData(65); xorBitMap(6)(64) := currentData(64); xorBitMap(6)(62) := currentData(62); xorBitMap(6)(60) := currentData(60); xorBitMap(6)(56) := currentData(56); xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(162) := previousCrc(2); xorBitMap(6)(163) := previousCrc(3); xorBitMap(6)(164) := previousCrc(4); xorBitMap(6)(166) := previousCrc(6); xorBitMap(6)(167) := previousCrc(7); xorBitMap(6)(168) := previousCrc(8); xorBitMap(6)(172) := previousCrc(12); xorBitMap(6)(174) := previousCrc(14); xorBitMap(6)(176) := previousCrc(16); xorBitMap(6)(177) := previousCrc(17); xorBitMap(6)(178) := previousCrc(18); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(182) := previousCrc(22); xorBitMap(6)(183) := previousCrc(23); xorBitMap(6)(184) := previousCrc(24); xorBitMap(6)(185) := previousCrc(25); xorBitMap(6)(186) := previousCrc(26); xorBitMap(6)(187) := previousCrc(27); xorBitMap(6)(188) := previousCrc(28); xorBitMap(6)(191) := previousCrc(31); 
      xorBitMap(7)(79) := currentData(79); xorBitMap(7)(77) := currentData(77); xorBitMap(7)(76) := currentData(76); xorBitMap(7)(75) := currentData(75); xorBitMap(7)(74) := currentData(74); xorBitMap(7)(71) := currentData(71); xorBitMap(7)(69) := currentData(69); xorBitMap(7)(68) := currentData(68); xorBitMap(7)(60) := currentData(60); xorBitMap(7)(58) := currentData(58); xorBitMap(7)(57) := currentData(57); xorBitMap(7)(56) := currentData(56); xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(162) := previousCrc(2); xorBitMap(7)(163) := previousCrc(3); xorBitMap(7)(164) := previousCrc(4); xorBitMap(7)(166) := previousCrc(6); xorBitMap(7)(168) := previousCrc(8); xorBitMap(7)(169) := previousCrc(9); xorBitMap(7)(170) := previousCrc(10); xorBitMap(7)(172) := previousCrc(12); xorBitMap(7)(180) := previousCrc(20); xorBitMap(7)(181) := previousCrc(21); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(186) := previousCrc(26); xorBitMap(7)(187) := previousCrc(27); xorBitMap(7)(188) := previousCrc(28); xorBitMap(7)(189) := previousCrc(29); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(79) := currentData(79); xorBitMap(8)(78) := currentData(78); xorBitMap(8)(77) := currentData(77); xorBitMap(8)(76) := currentData(76); xorBitMap(8)(75) := currentData(75); xorBitMap(8)(73) := currentData(73); xorBitMap(8)(70) := currentData(70); xorBitMap(8)(69) := currentData(69); xorBitMap(8)(68) := currentData(68); xorBitMap(8)(67) := currentData(67); xorBitMap(8)(66) := currentData(66); xorBitMap(8)(65) := currentData(65); xorBitMap(8)(63) := currentData(63); xorBitMap(8)(60) := currentData(60); xorBitMap(8)(59) := currentData(59); xorBitMap(8)(57) := currentData(57); xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(162) := previousCrc(2); xorBitMap(8)(163) := previousCrc(3); xorBitMap(8)(164) := previousCrc(4); xorBitMap(8)(166) := previousCrc(6); xorBitMap(8)(169) := previousCrc(9); xorBitMap(8)(171) := previousCrc(11); xorBitMap(8)(172) := previousCrc(12); xorBitMap(8)(175) := previousCrc(15); xorBitMap(8)(177) := previousCrc(17); xorBitMap(8)(178) := previousCrc(18); xorBitMap(8)(179) := previousCrc(19); xorBitMap(8)(180) := previousCrc(20); xorBitMap(8)(181) := previousCrc(21); xorBitMap(8)(182) := previousCrc(22); xorBitMap(8)(185) := previousCrc(25); xorBitMap(8)(187) := previousCrc(27); xorBitMap(8)(188) := previousCrc(28); xorBitMap(8)(189) := previousCrc(29); xorBitMap(8)(190) := previousCrc(30); xorBitMap(8)(191) := previousCrc(31); 
      xorBitMap(9)(79) := currentData(79); xorBitMap(9)(78) := currentData(78); xorBitMap(9)(77) := currentData(77); xorBitMap(9)(76) := currentData(76); xorBitMap(9)(74) := currentData(74); xorBitMap(9)(71) := currentData(71); xorBitMap(9)(70) := currentData(70); xorBitMap(9)(69) := currentData(69); xorBitMap(9)(68) := currentData(68); xorBitMap(9)(67) := currentData(67); xorBitMap(9)(66) := currentData(66); xorBitMap(9)(64) := currentData(64); xorBitMap(9)(61) := currentData(61); xorBitMap(9)(60) := currentData(60); xorBitMap(9)(58) := currentData(58); xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(163) := previousCrc(3); xorBitMap(9)(164) := previousCrc(4); xorBitMap(9)(165) := previousCrc(5); xorBitMap(9)(167) := previousCrc(7); xorBitMap(9)(170) := previousCrc(10); xorBitMap(9)(172) := previousCrc(12); xorBitMap(9)(173) := previousCrc(13); xorBitMap(9)(176) := previousCrc(16); xorBitMap(9)(178) := previousCrc(18); xorBitMap(9)(179) := previousCrc(19); xorBitMap(9)(180) := previousCrc(20); xorBitMap(9)(181) := previousCrc(21); xorBitMap(9)(182) := previousCrc(22); xorBitMap(9)(183) := previousCrc(23); xorBitMap(9)(186) := previousCrc(26); xorBitMap(9)(188) := previousCrc(28); xorBitMap(9)(189) := previousCrc(29); xorBitMap(9)(190) := previousCrc(30); xorBitMap(9)(191) := previousCrc(31); 
      xorBitMap(10)(78) := currentData(78); xorBitMap(10)(77) := currentData(77); xorBitMap(10)(75) := currentData(75); xorBitMap(10)(73) := currentData(73); xorBitMap(10)(71) := currentData(71); xorBitMap(10)(70) := currentData(70); xorBitMap(10)(69) := currentData(69); xorBitMap(10)(66) := currentData(66); xorBitMap(10)(63) := currentData(63); xorBitMap(10)(62) := currentData(62); xorBitMap(10)(60) := currentData(60); xorBitMap(10)(59) := currentData(59); xorBitMap(10)(58) := currentData(58); xorBitMap(10)(56) := currentData(56); xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(162) := previousCrc(2); xorBitMap(10)(164) := previousCrc(4); xorBitMap(10)(167) := previousCrc(7); xorBitMap(10)(168) := previousCrc(8); xorBitMap(10)(170) := previousCrc(10); xorBitMap(10)(171) := previousCrc(11); xorBitMap(10)(172) := previousCrc(12); xorBitMap(10)(174) := previousCrc(14); xorBitMap(10)(175) := previousCrc(15); xorBitMap(10)(178) := previousCrc(18); xorBitMap(10)(181) := previousCrc(21); xorBitMap(10)(182) := previousCrc(22); xorBitMap(10)(183) := previousCrc(23); xorBitMap(10)(185) := previousCrc(25); xorBitMap(10)(187) := previousCrc(27); xorBitMap(10)(189) := previousCrc(29); xorBitMap(10)(190) := previousCrc(30); 
      xorBitMap(11)(78) := currentData(78); xorBitMap(11)(76) := currentData(76); xorBitMap(11)(74) := currentData(74); xorBitMap(11)(73) := currentData(73); xorBitMap(11)(71) := currentData(71); xorBitMap(11)(70) := currentData(70); xorBitMap(11)(68) := currentData(68); xorBitMap(11)(66) := currentData(66); xorBitMap(11)(65) := currentData(65); xorBitMap(11)(64) := currentData(64); xorBitMap(11)(59) := currentData(59); xorBitMap(11)(58) := currentData(58); xorBitMap(11)(57) := currentData(57); xorBitMap(11)(56) := currentData(56); xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(160) := previousCrc(0); xorBitMap(11)(162) := previousCrc(2); xorBitMap(11)(163) := previousCrc(3); xorBitMap(11)(166) := previousCrc(6); xorBitMap(11)(167) := previousCrc(7); xorBitMap(11)(168) := previousCrc(8); xorBitMap(11)(169) := previousCrc(9); xorBitMap(11)(170) := previousCrc(10); xorBitMap(11)(171) := previousCrc(11); xorBitMap(11)(176) := previousCrc(16); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(178) := previousCrc(18); xorBitMap(11)(180) := previousCrc(20); xorBitMap(11)(182) := previousCrc(22); xorBitMap(11)(183) := previousCrc(23); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(186) := previousCrc(26); xorBitMap(11)(188) := previousCrc(28); xorBitMap(11)(190) := previousCrc(30); 
      xorBitMap(12)(77) := currentData(77); xorBitMap(12)(75) := currentData(75); xorBitMap(12)(74) := currentData(74); xorBitMap(12)(73) := currentData(73); xorBitMap(12)(71) := currentData(71); xorBitMap(12)(69) := currentData(69); xorBitMap(12)(68) := currentData(68); xorBitMap(12)(63) := currentData(63); xorBitMap(12)(61) := currentData(61); xorBitMap(12)(59) := currentData(59); xorBitMap(12)(57) := currentData(57); xorBitMap(12)(56) := currentData(56); xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(161) := previousCrc(1); xorBitMap(12)(162) := previousCrc(2); xorBitMap(12)(163) := previousCrc(3); xorBitMap(12)(164) := previousCrc(4); xorBitMap(12)(165) := previousCrc(5); xorBitMap(12)(166) := previousCrc(6); xorBitMap(12)(168) := previousCrc(8); xorBitMap(12)(169) := previousCrc(9); xorBitMap(12)(171) := previousCrc(11); xorBitMap(12)(173) := previousCrc(13); xorBitMap(12)(175) := previousCrc(15); xorBitMap(12)(180) := previousCrc(20); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(183) := previousCrc(23); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(186) := previousCrc(26); xorBitMap(12)(187) := previousCrc(27); xorBitMap(12)(189) := previousCrc(29); 
      xorBitMap(13)(78) := currentData(78); xorBitMap(13)(76) := currentData(76); xorBitMap(13)(75) := currentData(75); xorBitMap(13)(74) := currentData(74); xorBitMap(13)(72) := currentData(72); xorBitMap(13)(70) := currentData(70); xorBitMap(13)(69) := currentData(69); xorBitMap(13)(64) := currentData(64); xorBitMap(13)(62) := currentData(62); xorBitMap(13)(60) := currentData(60); xorBitMap(13)(58) := currentData(58); xorBitMap(13)(57) := currentData(57); xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(160) := previousCrc(0); xorBitMap(13)(162) := previousCrc(2); xorBitMap(13)(163) := previousCrc(3); xorBitMap(13)(164) := previousCrc(4); xorBitMap(13)(165) := previousCrc(5); xorBitMap(13)(166) := previousCrc(6); xorBitMap(13)(167) := previousCrc(7); xorBitMap(13)(169) := previousCrc(9); xorBitMap(13)(170) := previousCrc(10); xorBitMap(13)(172) := previousCrc(12); xorBitMap(13)(174) := previousCrc(14); xorBitMap(13)(176) := previousCrc(16); xorBitMap(13)(181) := previousCrc(21); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(184) := previousCrc(24); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(187) := previousCrc(27); xorBitMap(13)(188) := previousCrc(28); xorBitMap(13)(190) := previousCrc(30); 
      xorBitMap(14)(79) := currentData(79); xorBitMap(14)(77) := currentData(77); xorBitMap(14)(76) := currentData(76); xorBitMap(14)(75) := currentData(75); xorBitMap(14)(73) := currentData(73); xorBitMap(14)(71) := currentData(71); xorBitMap(14)(70) := currentData(70); xorBitMap(14)(65) := currentData(65); xorBitMap(14)(63) := currentData(63); xorBitMap(14)(61) := currentData(61); xorBitMap(14)(59) := currentData(59); xorBitMap(14)(58) := currentData(58); xorBitMap(14)(56) := currentData(56); xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(160) := previousCrc(0); xorBitMap(14)(161) := previousCrc(1); xorBitMap(14)(163) := previousCrc(3); xorBitMap(14)(164) := previousCrc(4); xorBitMap(14)(165) := previousCrc(5); xorBitMap(14)(166) := previousCrc(6); xorBitMap(14)(167) := previousCrc(7); xorBitMap(14)(168) := previousCrc(8); xorBitMap(14)(170) := previousCrc(10); xorBitMap(14)(171) := previousCrc(11); xorBitMap(14)(173) := previousCrc(13); xorBitMap(14)(175) := previousCrc(15); xorBitMap(14)(177) := previousCrc(17); xorBitMap(14)(182) := previousCrc(22); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(185) := previousCrc(25); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(188) := previousCrc(28); xorBitMap(14)(189) := previousCrc(29); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(78) := currentData(78); xorBitMap(15)(77) := currentData(77); xorBitMap(15)(76) := currentData(76); xorBitMap(15)(74) := currentData(74); xorBitMap(15)(72) := currentData(72); xorBitMap(15)(71) := currentData(71); xorBitMap(15)(66) := currentData(66); xorBitMap(15)(64) := currentData(64); xorBitMap(15)(62) := currentData(62); xorBitMap(15)(60) := currentData(60); xorBitMap(15)(59) := currentData(59); xorBitMap(15)(57) := currentData(57); xorBitMap(15)(56) := currentData(56); xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(161) := previousCrc(1); xorBitMap(15)(162) := previousCrc(2); xorBitMap(15)(164) := previousCrc(4); xorBitMap(15)(165) := previousCrc(5); xorBitMap(15)(166) := previousCrc(6); xorBitMap(15)(167) := previousCrc(7); xorBitMap(15)(168) := previousCrc(8); xorBitMap(15)(169) := previousCrc(9); xorBitMap(15)(171) := previousCrc(11); xorBitMap(15)(172) := previousCrc(12); xorBitMap(15)(174) := previousCrc(14); xorBitMap(15)(176) := previousCrc(16); xorBitMap(15)(178) := previousCrc(18); xorBitMap(15)(183) := previousCrc(23); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(186) := previousCrc(26); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(189) := previousCrc(29); xorBitMap(15)(190) := previousCrc(30); 
      xorBitMap(16)(78) := currentData(78); xorBitMap(16)(77) := currentData(77); xorBitMap(16)(75) := currentData(75); xorBitMap(16)(68) := currentData(68); xorBitMap(16)(66) := currentData(66); xorBitMap(16)(57) := currentData(57); xorBitMap(16)(56) := currentData(56); xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(160) := previousCrc(0); xorBitMap(16)(163) := previousCrc(3); xorBitMap(16)(168) := previousCrc(8); xorBitMap(16)(169) := previousCrc(9); xorBitMap(16)(178) := previousCrc(18); xorBitMap(16)(180) := previousCrc(20); xorBitMap(16)(187) := previousCrc(27); xorBitMap(16)(189) := previousCrc(29); xorBitMap(16)(190) := previousCrc(30); 
      xorBitMap(17)(79) := currentData(79); xorBitMap(17)(78) := currentData(78); xorBitMap(17)(76) := currentData(76); xorBitMap(17)(69) := currentData(69); xorBitMap(17)(67) := currentData(67); xorBitMap(17)(58) := currentData(58); xorBitMap(17)(57) := currentData(57); xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(160) := previousCrc(0); xorBitMap(17)(161) := previousCrc(1); xorBitMap(17)(164) := previousCrc(4); xorBitMap(17)(169) := previousCrc(9); xorBitMap(17)(170) := previousCrc(10); xorBitMap(17)(179) := previousCrc(19); xorBitMap(17)(181) := previousCrc(21); xorBitMap(17)(188) := previousCrc(28); xorBitMap(17)(190) := previousCrc(30); xorBitMap(17)(191) := previousCrc(31); 
      xorBitMap(18)(79) := currentData(79); xorBitMap(18)(77) := currentData(77); xorBitMap(18)(70) := currentData(70); xorBitMap(18)(68) := currentData(68); xorBitMap(18)(59) := currentData(59); xorBitMap(18)(58) := currentData(58); xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(160) := previousCrc(0); xorBitMap(18)(161) := previousCrc(1); xorBitMap(18)(162) := previousCrc(2); xorBitMap(18)(165) := previousCrc(5); xorBitMap(18)(170) := previousCrc(10); xorBitMap(18)(171) := previousCrc(11); xorBitMap(18)(180) := previousCrc(20); xorBitMap(18)(182) := previousCrc(22); xorBitMap(18)(189) := previousCrc(29); xorBitMap(18)(191) := previousCrc(31); 
      xorBitMap(19)(78) := currentData(78); xorBitMap(19)(71) := currentData(71); xorBitMap(19)(69) := currentData(69); xorBitMap(19)(60) := currentData(60); xorBitMap(19)(59) := currentData(59); xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(161) := previousCrc(1); xorBitMap(19)(162) := previousCrc(2); xorBitMap(19)(163) := previousCrc(3); xorBitMap(19)(166) := previousCrc(6); xorBitMap(19)(171) := previousCrc(11); xorBitMap(19)(172) := previousCrc(12); xorBitMap(19)(181) := previousCrc(21); xorBitMap(19)(183) := previousCrc(23); xorBitMap(19)(190) := previousCrc(30); 
      xorBitMap(20)(79) := currentData(79); xorBitMap(20)(72) := currentData(72); xorBitMap(20)(70) := currentData(70); xorBitMap(20)(61) := currentData(61); xorBitMap(20)(60) := currentData(60); xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(160) := previousCrc(0); xorBitMap(20)(162) := previousCrc(2); xorBitMap(20)(163) := previousCrc(3); xorBitMap(20)(164) := previousCrc(4); xorBitMap(20)(167) := previousCrc(7); xorBitMap(20)(172) := previousCrc(12); xorBitMap(20)(173) := previousCrc(13); xorBitMap(20)(182) := previousCrc(22); xorBitMap(20)(184) := previousCrc(24); xorBitMap(20)(191) := previousCrc(31); 
      xorBitMap(21)(73) := currentData(73); xorBitMap(21)(71) := currentData(71); xorBitMap(21)(62) := currentData(62); xorBitMap(21)(61) := currentData(61); xorBitMap(21)(56) := currentData(56); xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(161) := previousCrc(1); xorBitMap(21)(163) := previousCrc(3); xorBitMap(21)(164) := previousCrc(4); xorBitMap(21)(165) := previousCrc(5); xorBitMap(21)(168) := previousCrc(8); xorBitMap(21)(173) := previousCrc(13); xorBitMap(21)(174) := previousCrc(14); xorBitMap(21)(183) := previousCrc(23); xorBitMap(21)(185) := previousCrc(25); 
      xorBitMap(22)(79) := currentData(79); xorBitMap(22)(74) := currentData(74); xorBitMap(22)(73) := currentData(73); xorBitMap(22)(68) := currentData(68); xorBitMap(22)(67) := currentData(67); xorBitMap(22)(66) := currentData(66); xorBitMap(22)(65) := currentData(65); xorBitMap(22)(62) := currentData(62); xorBitMap(22)(61) := currentData(61); xorBitMap(22)(60) := currentData(60); xorBitMap(22)(58) := currentData(58); xorBitMap(22)(57) := currentData(57); xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(160) := previousCrc(0); xorBitMap(22)(164) := previousCrc(4); xorBitMap(22)(167) := previousCrc(7); xorBitMap(22)(169) := previousCrc(9); xorBitMap(22)(170) := previousCrc(10); xorBitMap(22)(172) := previousCrc(12); xorBitMap(22)(173) := previousCrc(13); xorBitMap(22)(174) := previousCrc(14); xorBitMap(22)(177) := previousCrc(17); xorBitMap(22)(178) := previousCrc(18); xorBitMap(22)(179) := previousCrc(19); xorBitMap(22)(180) := previousCrc(20); xorBitMap(22)(185) := previousCrc(25); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(191) := previousCrc(31); 
      xorBitMap(23)(79) := currentData(79); xorBitMap(23)(75) := currentData(75); xorBitMap(23)(74) := currentData(74); xorBitMap(23)(73) := currentData(73); xorBitMap(23)(72) := currentData(72); xorBitMap(23)(69) := currentData(69); xorBitMap(23)(65) := currentData(65); xorBitMap(23)(62) := currentData(62); xorBitMap(23)(60) := currentData(60); xorBitMap(23)(59) := currentData(59); xorBitMap(23)(56) := currentData(56); xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(161) := previousCrc(1); xorBitMap(23)(162) := previousCrc(2); xorBitMap(23)(166) := previousCrc(6); xorBitMap(23)(167) := previousCrc(7); xorBitMap(23)(168) := previousCrc(8); xorBitMap(23)(171) := previousCrc(11); xorBitMap(23)(172) := previousCrc(12); xorBitMap(23)(174) := previousCrc(14); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(181) := previousCrc(21); xorBitMap(23)(184) := previousCrc(24); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(186) := previousCrc(26); xorBitMap(23)(187) := previousCrc(27); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(76) := currentData(76); xorBitMap(24)(75) := currentData(75); xorBitMap(24)(74) := currentData(74); xorBitMap(24)(73) := currentData(73); xorBitMap(24)(70) := currentData(70); xorBitMap(24)(66) := currentData(66); xorBitMap(24)(63) := currentData(63); xorBitMap(24)(61) := currentData(61); xorBitMap(24)(60) := currentData(60); xorBitMap(24)(57) := currentData(57); xorBitMap(24)(56) := currentData(56); xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(160) := previousCrc(0); xorBitMap(24)(162) := previousCrc(2); xorBitMap(24)(163) := previousCrc(3); xorBitMap(24)(167) := previousCrc(7); xorBitMap(24)(168) := previousCrc(8); xorBitMap(24)(169) := previousCrc(9); xorBitMap(24)(172) := previousCrc(12); xorBitMap(24)(173) := previousCrc(13); xorBitMap(24)(175) := previousCrc(15); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(182) := previousCrc(22); xorBitMap(24)(185) := previousCrc(25); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(187) := previousCrc(27); xorBitMap(24)(188) := previousCrc(28); 
      xorBitMap(25)(77) := currentData(77); xorBitMap(25)(76) := currentData(76); xorBitMap(25)(75) := currentData(75); xorBitMap(25)(74) := currentData(74); xorBitMap(25)(71) := currentData(71); xorBitMap(25)(67) := currentData(67); xorBitMap(25)(64) := currentData(64); xorBitMap(25)(62) := currentData(62); xorBitMap(25)(61) := currentData(61); xorBitMap(25)(58) := currentData(58); xorBitMap(25)(57) := currentData(57); xorBitMap(25)(56) := currentData(56); xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(160) := previousCrc(0); xorBitMap(25)(161) := previousCrc(1); xorBitMap(25)(163) := previousCrc(3); xorBitMap(25)(164) := previousCrc(4); xorBitMap(25)(168) := previousCrc(8); xorBitMap(25)(169) := previousCrc(9); xorBitMap(25)(170) := previousCrc(10); xorBitMap(25)(173) := previousCrc(13); xorBitMap(25)(174) := previousCrc(14); xorBitMap(25)(176) := previousCrc(16); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(183) := previousCrc(23); xorBitMap(25)(186) := previousCrc(26); xorBitMap(25)(187) := previousCrc(27); xorBitMap(25)(188) := previousCrc(28); xorBitMap(25)(189) := previousCrc(29); 
      xorBitMap(26)(79) := currentData(79); xorBitMap(26)(78) := currentData(78); xorBitMap(26)(77) := currentData(77); xorBitMap(26)(76) := currentData(76); xorBitMap(26)(75) := currentData(75); xorBitMap(26)(73) := currentData(73); xorBitMap(26)(67) := currentData(67); xorBitMap(26)(66) := currentData(66); xorBitMap(26)(62) := currentData(62); xorBitMap(26)(61) := currentData(61); xorBitMap(26)(60) := currentData(60); xorBitMap(26)(59) := currentData(59); xorBitMap(26)(57) := currentData(57); xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(160) := previousCrc(0); xorBitMap(26)(161) := previousCrc(1); xorBitMap(26)(164) := previousCrc(4); xorBitMap(26)(166) := previousCrc(6); xorBitMap(26)(167) := previousCrc(7); xorBitMap(26)(169) := previousCrc(9); xorBitMap(26)(171) := previousCrc(11); xorBitMap(26)(172) := previousCrc(12); xorBitMap(26)(173) := previousCrc(13); xorBitMap(26)(174) := previousCrc(14); xorBitMap(26)(178) := previousCrc(18); xorBitMap(26)(179) := previousCrc(19); xorBitMap(26)(185) := previousCrc(25); xorBitMap(26)(187) := previousCrc(27); xorBitMap(26)(188) := previousCrc(28); xorBitMap(26)(189) := previousCrc(29); xorBitMap(26)(190) := previousCrc(30); xorBitMap(26)(191) := previousCrc(31); 
      xorBitMap(27)(79) := currentData(79); xorBitMap(27)(78) := currentData(78); xorBitMap(27)(77) := currentData(77); xorBitMap(27)(76) := currentData(76); xorBitMap(27)(74) := currentData(74); xorBitMap(27)(68) := currentData(68); xorBitMap(27)(67) := currentData(67); xorBitMap(27)(63) := currentData(63); xorBitMap(27)(62) := currentData(62); xorBitMap(27)(61) := currentData(61); xorBitMap(27)(60) := currentData(60); xorBitMap(27)(58) := currentData(58); xorBitMap(27)(56) := currentData(56); xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(160) := previousCrc(0); xorBitMap(27)(161) := previousCrc(1); xorBitMap(27)(162) := previousCrc(2); xorBitMap(27)(165) := previousCrc(5); xorBitMap(27)(167) := previousCrc(7); xorBitMap(27)(168) := previousCrc(8); xorBitMap(27)(170) := previousCrc(10); xorBitMap(27)(172) := previousCrc(12); xorBitMap(27)(173) := previousCrc(13); xorBitMap(27)(174) := previousCrc(14); xorBitMap(27)(175) := previousCrc(15); xorBitMap(27)(179) := previousCrc(19); xorBitMap(27)(180) := previousCrc(20); xorBitMap(27)(186) := previousCrc(26); xorBitMap(27)(188) := previousCrc(28); xorBitMap(27)(189) := previousCrc(29); xorBitMap(27)(190) := previousCrc(30); xorBitMap(27)(191) := previousCrc(31); 
      xorBitMap(28)(79) := currentData(79); xorBitMap(28)(78) := currentData(78); xorBitMap(28)(77) := currentData(77); xorBitMap(28)(75) := currentData(75); xorBitMap(28)(69) := currentData(69); xorBitMap(28)(68) := currentData(68); xorBitMap(28)(64) := currentData(64); xorBitMap(28)(63) := currentData(63); xorBitMap(28)(62) := currentData(62); xorBitMap(28)(61) := currentData(61); xorBitMap(28)(59) := currentData(59); xorBitMap(28)(57) := currentData(57); xorBitMap(28)(56) := currentData(56); xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(161) := previousCrc(1); xorBitMap(28)(162) := previousCrc(2); xorBitMap(28)(163) := previousCrc(3); xorBitMap(28)(166) := previousCrc(6); xorBitMap(28)(168) := previousCrc(8); xorBitMap(28)(169) := previousCrc(9); xorBitMap(28)(171) := previousCrc(11); xorBitMap(28)(173) := previousCrc(13); xorBitMap(28)(174) := previousCrc(14); xorBitMap(28)(175) := previousCrc(15); xorBitMap(28)(176) := previousCrc(16); xorBitMap(28)(180) := previousCrc(20); xorBitMap(28)(181) := previousCrc(21); xorBitMap(28)(187) := previousCrc(27); xorBitMap(28)(189) := previousCrc(29); xorBitMap(28)(190) := previousCrc(30); xorBitMap(28)(191) := previousCrc(31); 
      xorBitMap(29)(79) := currentData(79); xorBitMap(29)(78) := currentData(78); xorBitMap(29)(76) := currentData(76); xorBitMap(29)(70) := currentData(70); xorBitMap(29)(69) := currentData(69); xorBitMap(29)(65) := currentData(65); xorBitMap(29)(64) := currentData(64); xorBitMap(29)(63) := currentData(63); xorBitMap(29)(62) := currentData(62); xorBitMap(29)(60) := currentData(60); xorBitMap(29)(58) := currentData(58); xorBitMap(29)(57) := currentData(57); xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(162) := previousCrc(2); xorBitMap(29)(163) := previousCrc(3); xorBitMap(29)(164) := previousCrc(4); xorBitMap(29)(167) := previousCrc(7); xorBitMap(29)(169) := previousCrc(9); xorBitMap(29)(170) := previousCrc(10); xorBitMap(29)(172) := previousCrc(12); xorBitMap(29)(174) := previousCrc(14); xorBitMap(29)(175) := previousCrc(15); xorBitMap(29)(176) := previousCrc(16); xorBitMap(29)(177) := previousCrc(17); xorBitMap(29)(181) := previousCrc(21); xorBitMap(29)(182) := previousCrc(22); xorBitMap(29)(188) := previousCrc(28); xorBitMap(29)(190) := previousCrc(30); xorBitMap(29)(191) := previousCrc(31); 
      xorBitMap(30)(79) := currentData(79); xorBitMap(30)(77) := currentData(77); xorBitMap(30)(71) := currentData(71); xorBitMap(30)(70) := currentData(70); xorBitMap(30)(66) := currentData(66); xorBitMap(30)(65) := currentData(65); xorBitMap(30)(64) := currentData(64); xorBitMap(30)(63) := currentData(63); xorBitMap(30)(61) := currentData(61); xorBitMap(30)(59) := currentData(59); xorBitMap(30)(58) := currentData(58); xorBitMap(30)(56) := currentData(56); xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(160) := previousCrc(0); xorBitMap(30)(163) := previousCrc(3); xorBitMap(30)(164) := previousCrc(4); xorBitMap(30)(165) := previousCrc(5); xorBitMap(30)(168) := previousCrc(8); xorBitMap(30)(170) := previousCrc(10); xorBitMap(30)(171) := previousCrc(11); xorBitMap(30)(173) := previousCrc(13); xorBitMap(30)(175) := previousCrc(15); xorBitMap(30)(176) := previousCrc(16); xorBitMap(30)(177) := previousCrc(17); xorBitMap(30)(178) := previousCrc(18); xorBitMap(30)(182) := previousCrc(22); xorBitMap(30)(183) := previousCrc(23); xorBitMap(30)(189) := previousCrc(29); xorBitMap(30)(191) := previousCrc(31); 
      xorBitMap(31)(78) := currentData(78); xorBitMap(31)(72) := currentData(72); xorBitMap(31)(71) := currentData(71); xorBitMap(31)(67) := currentData(67); xorBitMap(31)(66) := currentData(66); xorBitMap(31)(65) := currentData(65); xorBitMap(31)(64) := currentData(64); xorBitMap(31)(62) := currentData(62); xorBitMap(31)(60) := currentData(60); xorBitMap(31)(59) := currentData(59); xorBitMap(31)(57) := currentData(57); xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(161) := previousCrc(1); xorBitMap(31)(164) := previousCrc(4); xorBitMap(31)(165) := previousCrc(5); xorBitMap(31)(166) := previousCrc(6); xorBitMap(31)(169) := previousCrc(9); xorBitMap(31)(171) := previousCrc(11); xorBitMap(31)(172) := previousCrc(12); xorBitMap(31)(174) := previousCrc(14); xorBitMap(31)(176) := previousCrc(16); xorBitMap(31)(177) := previousCrc(17); xorBitMap(31)(178) := previousCrc(18); xorBitMap(31)(179) := previousCrc(19); xorBitMap(31)(183) := previousCrc(23); xorBitMap(31)(184) := previousCrc(24); xorBitMap(31)(190) := previousCrc(30); 
   end procedure;

   procedure xorBitMap11Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(87 downto 0)) is 
   begin
      xorBitMap(0)(87) := currentData(87); xorBitMap(0)(85) := currentData(85); xorBitMap(0)(84) := currentData(84); xorBitMap(0)(83) := currentData(83); xorBitMap(0)(82) := currentData(82); xorBitMap(0)(81) := currentData(81); xorBitMap(0)(79) := currentData(79); xorBitMap(0)(73) := currentData(73); xorBitMap(0)(72) := currentData(72); xorBitMap(0)(68) := currentData(68); xorBitMap(0)(67) := currentData(67); xorBitMap(0)(66) := currentData(66); xorBitMap(0)(65) := currentData(65); xorBitMap(0)(63) := currentData(63); xorBitMap(0)(61) := currentData(61); xorBitMap(0)(60) := currentData(60); xorBitMap(0)(58) := currentData(58); xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(162) := previousCrc(2); xorBitMap(0)(164) := previousCrc(4); xorBitMap(0)(165) := previousCrc(5); xorBitMap(0)(167) := previousCrc(7); xorBitMap(0)(169) := previousCrc(9); xorBitMap(0)(170) := previousCrc(10); xorBitMap(0)(171) := previousCrc(11); xorBitMap(0)(172) := previousCrc(12); xorBitMap(0)(176) := previousCrc(16); xorBitMap(0)(177) := previousCrc(17); xorBitMap(0)(183) := previousCrc(23); xorBitMap(0)(185) := previousCrc(25); xorBitMap(0)(186) := previousCrc(26); xorBitMap(0)(187) := previousCrc(27); xorBitMap(0)(188) := previousCrc(28); xorBitMap(0)(189) := previousCrc(29); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(87) := currentData(87); xorBitMap(1)(86) := currentData(86); xorBitMap(1)(81) := currentData(81); xorBitMap(1)(80) := currentData(80); xorBitMap(1)(79) := currentData(79); xorBitMap(1)(74) := currentData(74); xorBitMap(1)(72) := currentData(72); xorBitMap(1)(69) := currentData(69); xorBitMap(1)(65) := currentData(65); xorBitMap(1)(64) := currentData(64); xorBitMap(1)(63) := currentData(63); xorBitMap(1)(62) := currentData(62); xorBitMap(1)(60) := currentData(60); xorBitMap(1)(59) := currentData(59); xorBitMap(1)(58) := currentData(58); xorBitMap(1)(56) := currentData(56); xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(160) := previousCrc(0); xorBitMap(1)(162) := previousCrc(2); xorBitMap(1)(163) := previousCrc(3); xorBitMap(1)(164) := previousCrc(4); xorBitMap(1)(166) := previousCrc(6); xorBitMap(1)(167) := previousCrc(7); xorBitMap(1)(168) := previousCrc(8); xorBitMap(1)(169) := previousCrc(9); xorBitMap(1)(173) := previousCrc(13); xorBitMap(1)(176) := previousCrc(16); xorBitMap(1)(178) := previousCrc(18); xorBitMap(1)(183) := previousCrc(23); xorBitMap(1)(184) := previousCrc(24); xorBitMap(1)(185) := previousCrc(25); xorBitMap(1)(190) := previousCrc(30); xorBitMap(1)(191) := previousCrc(31); 
      xorBitMap(2)(85) := currentData(85); xorBitMap(2)(84) := currentData(84); xorBitMap(2)(83) := currentData(83); xorBitMap(2)(80) := currentData(80); xorBitMap(2)(79) := currentData(79); xorBitMap(2)(75) := currentData(75); xorBitMap(2)(72) := currentData(72); xorBitMap(2)(70) := currentData(70); xorBitMap(2)(68) := currentData(68); xorBitMap(2)(67) := currentData(67); xorBitMap(2)(64) := currentData(64); xorBitMap(2)(59) := currentData(59); xorBitMap(2)(58) := currentData(58); xorBitMap(2)(57) := currentData(57); xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(161) := previousCrc(1); xorBitMap(2)(162) := previousCrc(2); xorBitMap(2)(163) := previousCrc(3); xorBitMap(2)(168) := previousCrc(8); xorBitMap(2)(171) := previousCrc(11); xorBitMap(2)(172) := previousCrc(12); xorBitMap(2)(174) := previousCrc(14); xorBitMap(2)(176) := previousCrc(16); xorBitMap(2)(179) := previousCrc(19); xorBitMap(2)(183) := previousCrc(23); xorBitMap(2)(184) := previousCrc(24); xorBitMap(2)(187) := previousCrc(27); xorBitMap(2)(188) := previousCrc(28); xorBitMap(2)(189) := previousCrc(29); 
      xorBitMap(3)(86) := currentData(86); xorBitMap(3)(85) := currentData(85); xorBitMap(3)(84) := currentData(84); xorBitMap(3)(81) := currentData(81); xorBitMap(3)(80) := currentData(80); xorBitMap(3)(76) := currentData(76); xorBitMap(3)(73) := currentData(73); xorBitMap(3)(71) := currentData(71); xorBitMap(3)(69) := currentData(69); xorBitMap(3)(68) := currentData(68); xorBitMap(3)(65) := currentData(65); xorBitMap(3)(60) := currentData(60); xorBitMap(3)(59) := currentData(59); xorBitMap(3)(58) := currentData(58); xorBitMap(3)(56) := currentData(56); xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(160) := previousCrc(0); xorBitMap(3)(162) := previousCrc(2); xorBitMap(3)(163) := previousCrc(3); xorBitMap(3)(164) := previousCrc(4); xorBitMap(3)(169) := previousCrc(9); xorBitMap(3)(172) := previousCrc(12); xorBitMap(3)(173) := previousCrc(13); xorBitMap(3)(175) := previousCrc(15); xorBitMap(3)(177) := previousCrc(17); xorBitMap(3)(180) := previousCrc(20); xorBitMap(3)(184) := previousCrc(24); xorBitMap(3)(185) := previousCrc(25); xorBitMap(3)(188) := previousCrc(28); xorBitMap(3)(189) := previousCrc(29); xorBitMap(3)(190) := previousCrc(30); 
      xorBitMap(4)(86) := currentData(86); xorBitMap(4)(84) := currentData(84); xorBitMap(4)(83) := currentData(83); xorBitMap(4)(79) := currentData(79); xorBitMap(4)(77) := currentData(77); xorBitMap(4)(74) := currentData(74); xorBitMap(4)(73) := currentData(73); xorBitMap(4)(70) := currentData(70); xorBitMap(4)(69) := currentData(69); xorBitMap(4)(68) := currentData(68); xorBitMap(4)(67) := currentData(67); xorBitMap(4)(65) := currentData(65); xorBitMap(4)(63) := currentData(63); xorBitMap(4)(59) := currentData(59); xorBitMap(4)(58) := currentData(58); xorBitMap(4)(57) := currentData(57); xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(161) := previousCrc(1); xorBitMap(4)(162) := previousCrc(2); xorBitMap(4)(163) := previousCrc(3); xorBitMap(4)(167) := previousCrc(7); xorBitMap(4)(169) := previousCrc(9); xorBitMap(4)(171) := previousCrc(11); xorBitMap(4)(172) := previousCrc(12); xorBitMap(4)(173) := previousCrc(13); xorBitMap(4)(174) := previousCrc(14); xorBitMap(4)(177) := previousCrc(17); xorBitMap(4)(178) := previousCrc(18); xorBitMap(4)(181) := previousCrc(21); xorBitMap(4)(183) := previousCrc(23); xorBitMap(4)(187) := previousCrc(27); xorBitMap(4)(188) := previousCrc(28); xorBitMap(4)(190) := previousCrc(30); 
      xorBitMap(5)(83) := currentData(83); xorBitMap(5)(82) := currentData(82); xorBitMap(5)(81) := currentData(81); xorBitMap(5)(80) := currentData(80); xorBitMap(5)(79) := currentData(79); xorBitMap(5)(78) := currentData(78); xorBitMap(5)(75) := currentData(75); xorBitMap(5)(74) := currentData(74); xorBitMap(5)(73) := currentData(73); xorBitMap(5)(72) := currentData(72); xorBitMap(5)(71) := currentData(71); xorBitMap(5)(70) := currentData(70); xorBitMap(5)(69) := currentData(69); xorBitMap(5)(67) := currentData(67); xorBitMap(5)(65) := currentData(65); xorBitMap(5)(64) := currentData(64); xorBitMap(5)(63) := currentData(63); xorBitMap(5)(61) := currentData(61); xorBitMap(5)(59) := currentData(59); xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(163) := previousCrc(3); xorBitMap(5)(165) := previousCrc(5); xorBitMap(5)(167) := previousCrc(7); xorBitMap(5)(168) := previousCrc(8); xorBitMap(5)(169) := previousCrc(9); xorBitMap(5)(171) := previousCrc(11); xorBitMap(5)(173) := previousCrc(13); xorBitMap(5)(174) := previousCrc(14); xorBitMap(5)(175) := previousCrc(15); xorBitMap(5)(176) := previousCrc(16); xorBitMap(5)(177) := previousCrc(17); xorBitMap(5)(178) := previousCrc(18); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(182) := previousCrc(22); xorBitMap(5)(183) := previousCrc(23); xorBitMap(5)(184) := previousCrc(24); xorBitMap(5)(185) := previousCrc(25); xorBitMap(5)(186) := previousCrc(26); xorBitMap(5)(187) := previousCrc(27); 
      xorBitMap(6)(84) := currentData(84); xorBitMap(6)(83) := currentData(83); xorBitMap(6)(82) := currentData(82); xorBitMap(6)(81) := currentData(81); xorBitMap(6)(80) := currentData(80); xorBitMap(6)(79) := currentData(79); xorBitMap(6)(76) := currentData(76); xorBitMap(6)(75) := currentData(75); xorBitMap(6)(74) := currentData(74); xorBitMap(6)(73) := currentData(73); xorBitMap(6)(72) := currentData(72); xorBitMap(6)(71) := currentData(71); xorBitMap(6)(70) := currentData(70); xorBitMap(6)(68) := currentData(68); xorBitMap(6)(66) := currentData(66); xorBitMap(6)(65) := currentData(65); xorBitMap(6)(64) := currentData(64); xorBitMap(6)(62) := currentData(62); xorBitMap(6)(60) := currentData(60); xorBitMap(6)(56) := currentData(56); xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(160) := previousCrc(0); xorBitMap(6)(164) := previousCrc(4); xorBitMap(6)(166) := previousCrc(6); xorBitMap(6)(168) := previousCrc(8); xorBitMap(6)(169) := previousCrc(9); xorBitMap(6)(170) := previousCrc(10); xorBitMap(6)(172) := previousCrc(12); xorBitMap(6)(174) := previousCrc(14); xorBitMap(6)(175) := previousCrc(15); xorBitMap(6)(176) := previousCrc(16); xorBitMap(6)(177) := previousCrc(17); xorBitMap(6)(178) := previousCrc(18); xorBitMap(6)(179) := previousCrc(19); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(183) := previousCrc(23); xorBitMap(6)(184) := previousCrc(24); xorBitMap(6)(185) := previousCrc(25); xorBitMap(6)(186) := previousCrc(26); xorBitMap(6)(187) := previousCrc(27); xorBitMap(6)(188) := previousCrc(28); 
      xorBitMap(7)(87) := currentData(87); xorBitMap(7)(80) := currentData(80); xorBitMap(7)(79) := currentData(79); xorBitMap(7)(77) := currentData(77); xorBitMap(7)(76) := currentData(76); xorBitMap(7)(75) := currentData(75); xorBitMap(7)(74) := currentData(74); xorBitMap(7)(71) := currentData(71); xorBitMap(7)(69) := currentData(69); xorBitMap(7)(68) := currentData(68); xorBitMap(7)(60) := currentData(60); xorBitMap(7)(58) := currentData(58); xorBitMap(7)(57) := currentData(57); xorBitMap(7)(56) := currentData(56); xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(160) := previousCrc(0); xorBitMap(7)(161) := previousCrc(1); xorBitMap(7)(162) := previousCrc(2); xorBitMap(7)(164) := previousCrc(4); xorBitMap(7)(172) := previousCrc(12); xorBitMap(7)(173) := previousCrc(13); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(178) := previousCrc(18); xorBitMap(7)(179) := previousCrc(19); xorBitMap(7)(180) := previousCrc(20); xorBitMap(7)(181) := previousCrc(21); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(184) := previousCrc(24); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(87) := currentData(87); xorBitMap(8)(85) := currentData(85); xorBitMap(8)(84) := currentData(84); xorBitMap(8)(83) := currentData(83); xorBitMap(8)(82) := currentData(82); xorBitMap(8)(80) := currentData(80); xorBitMap(8)(79) := currentData(79); xorBitMap(8)(78) := currentData(78); xorBitMap(8)(77) := currentData(77); xorBitMap(8)(76) := currentData(76); xorBitMap(8)(75) := currentData(75); xorBitMap(8)(73) := currentData(73); xorBitMap(8)(70) := currentData(70); xorBitMap(8)(69) := currentData(69); xorBitMap(8)(68) := currentData(68); xorBitMap(8)(67) := currentData(67); xorBitMap(8)(66) := currentData(66); xorBitMap(8)(65) := currentData(65); xorBitMap(8)(63) := currentData(63); xorBitMap(8)(60) := currentData(60); xorBitMap(8)(59) := currentData(59); xorBitMap(8)(57) := currentData(57); xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(161) := previousCrc(1); xorBitMap(8)(163) := previousCrc(3); xorBitMap(8)(164) := previousCrc(4); xorBitMap(8)(167) := previousCrc(7); xorBitMap(8)(169) := previousCrc(9); xorBitMap(8)(170) := previousCrc(10); xorBitMap(8)(171) := previousCrc(11); xorBitMap(8)(172) := previousCrc(12); xorBitMap(8)(173) := previousCrc(13); xorBitMap(8)(174) := previousCrc(14); xorBitMap(8)(177) := previousCrc(17); xorBitMap(8)(179) := previousCrc(19); xorBitMap(8)(180) := previousCrc(20); xorBitMap(8)(181) := previousCrc(21); xorBitMap(8)(182) := previousCrc(22); xorBitMap(8)(183) := previousCrc(23); xorBitMap(8)(184) := previousCrc(24); xorBitMap(8)(186) := previousCrc(26); xorBitMap(8)(187) := previousCrc(27); xorBitMap(8)(188) := previousCrc(28); xorBitMap(8)(189) := previousCrc(29); xorBitMap(8)(191) := previousCrc(31); 
      xorBitMap(9)(86) := currentData(86); xorBitMap(9)(85) := currentData(85); xorBitMap(9)(84) := currentData(84); xorBitMap(9)(83) := currentData(83); xorBitMap(9)(81) := currentData(81); xorBitMap(9)(80) := currentData(80); xorBitMap(9)(79) := currentData(79); xorBitMap(9)(78) := currentData(78); xorBitMap(9)(77) := currentData(77); xorBitMap(9)(76) := currentData(76); xorBitMap(9)(74) := currentData(74); xorBitMap(9)(71) := currentData(71); xorBitMap(9)(70) := currentData(70); xorBitMap(9)(69) := currentData(69); xorBitMap(9)(68) := currentData(68); xorBitMap(9)(67) := currentData(67); xorBitMap(9)(66) := currentData(66); xorBitMap(9)(64) := currentData(64); xorBitMap(9)(61) := currentData(61); xorBitMap(9)(60) := currentData(60); xorBitMap(9)(58) := currentData(58); xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(162) := previousCrc(2); xorBitMap(9)(164) := previousCrc(4); xorBitMap(9)(165) := previousCrc(5); xorBitMap(9)(168) := previousCrc(8); xorBitMap(9)(170) := previousCrc(10); xorBitMap(9)(171) := previousCrc(11); xorBitMap(9)(172) := previousCrc(12); xorBitMap(9)(173) := previousCrc(13); xorBitMap(9)(174) := previousCrc(14); xorBitMap(9)(175) := previousCrc(15); xorBitMap(9)(178) := previousCrc(18); xorBitMap(9)(180) := previousCrc(20); xorBitMap(9)(181) := previousCrc(21); xorBitMap(9)(182) := previousCrc(22); xorBitMap(9)(183) := previousCrc(23); xorBitMap(9)(184) := previousCrc(24); xorBitMap(9)(185) := previousCrc(25); xorBitMap(9)(187) := previousCrc(27); xorBitMap(9)(188) := previousCrc(28); xorBitMap(9)(189) := previousCrc(29); xorBitMap(9)(190) := previousCrc(30); 
      xorBitMap(10)(86) := currentData(86); xorBitMap(10)(83) := currentData(83); xorBitMap(10)(80) := currentData(80); xorBitMap(10)(78) := currentData(78); xorBitMap(10)(77) := currentData(77); xorBitMap(10)(75) := currentData(75); xorBitMap(10)(73) := currentData(73); xorBitMap(10)(71) := currentData(71); xorBitMap(10)(70) := currentData(70); xorBitMap(10)(69) := currentData(69); xorBitMap(10)(66) := currentData(66); xorBitMap(10)(63) := currentData(63); xorBitMap(10)(62) := currentData(62); xorBitMap(10)(60) := currentData(60); xorBitMap(10)(59) := currentData(59); xorBitMap(10)(58) := currentData(58); xorBitMap(10)(56) := currentData(56); xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(160) := previousCrc(0); xorBitMap(10)(162) := previousCrc(2); xorBitMap(10)(163) := previousCrc(3); xorBitMap(10)(164) := previousCrc(4); xorBitMap(10)(166) := previousCrc(6); xorBitMap(10)(167) := previousCrc(7); xorBitMap(10)(170) := previousCrc(10); xorBitMap(10)(173) := previousCrc(13); xorBitMap(10)(174) := previousCrc(14); xorBitMap(10)(175) := previousCrc(15); xorBitMap(10)(177) := previousCrc(17); xorBitMap(10)(179) := previousCrc(19); xorBitMap(10)(181) := previousCrc(21); xorBitMap(10)(182) := previousCrc(22); xorBitMap(10)(184) := previousCrc(24); xorBitMap(10)(187) := previousCrc(27); xorBitMap(10)(190) := previousCrc(30); 
      xorBitMap(11)(85) := currentData(85); xorBitMap(11)(83) := currentData(83); xorBitMap(11)(82) := currentData(82); xorBitMap(11)(78) := currentData(78); xorBitMap(11)(76) := currentData(76); xorBitMap(11)(74) := currentData(74); xorBitMap(11)(73) := currentData(73); xorBitMap(11)(71) := currentData(71); xorBitMap(11)(70) := currentData(70); xorBitMap(11)(68) := currentData(68); xorBitMap(11)(66) := currentData(66); xorBitMap(11)(65) := currentData(65); xorBitMap(11)(64) := currentData(64); xorBitMap(11)(59) := currentData(59); xorBitMap(11)(58) := currentData(58); xorBitMap(11)(57) := currentData(57); xorBitMap(11)(56) := currentData(56); xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(160) := previousCrc(0); xorBitMap(11)(161) := previousCrc(1); xorBitMap(11)(162) := previousCrc(2); xorBitMap(11)(163) := previousCrc(3); xorBitMap(11)(168) := previousCrc(8); xorBitMap(11)(169) := previousCrc(9); xorBitMap(11)(170) := previousCrc(10); xorBitMap(11)(172) := previousCrc(12); xorBitMap(11)(174) := previousCrc(14); xorBitMap(11)(175) := previousCrc(15); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(178) := previousCrc(18); xorBitMap(11)(180) := previousCrc(20); xorBitMap(11)(182) := previousCrc(22); xorBitMap(11)(186) := previousCrc(26); xorBitMap(11)(187) := previousCrc(27); xorBitMap(11)(189) := previousCrc(29); 
      xorBitMap(12)(87) := currentData(87); xorBitMap(12)(86) := currentData(86); xorBitMap(12)(85) := currentData(85); xorBitMap(12)(82) := currentData(82); xorBitMap(12)(81) := currentData(81); xorBitMap(12)(77) := currentData(77); xorBitMap(12)(75) := currentData(75); xorBitMap(12)(74) := currentData(74); xorBitMap(12)(73) := currentData(73); xorBitMap(12)(71) := currentData(71); xorBitMap(12)(69) := currentData(69); xorBitMap(12)(68) := currentData(68); xorBitMap(12)(63) := currentData(63); xorBitMap(12)(61) := currentData(61); xorBitMap(12)(59) := currentData(59); xorBitMap(12)(57) := currentData(57); xorBitMap(12)(56) := currentData(56); xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(160) := previousCrc(0); xorBitMap(12)(161) := previousCrc(1); xorBitMap(12)(163) := previousCrc(3); xorBitMap(12)(165) := previousCrc(5); xorBitMap(12)(167) := previousCrc(7); xorBitMap(12)(172) := previousCrc(12); xorBitMap(12)(173) := previousCrc(13); xorBitMap(12)(175) := previousCrc(15); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(178) := previousCrc(18); xorBitMap(12)(179) := previousCrc(19); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(186) := previousCrc(26); xorBitMap(12)(189) := previousCrc(29); xorBitMap(12)(190) := previousCrc(30); xorBitMap(12)(191) := previousCrc(31); 
      xorBitMap(13)(87) := currentData(87); xorBitMap(13)(86) := currentData(86); xorBitMap(13)(83) := currentData(83); xorBitMap(13)(82) := currentData(82); xorBitMap(13)(78) := currentData(78); xorBitMap(13)(76) := currentData(76); xorBitMap(13)(75) := currentData(75); xorBitMap(13)(74) := currentData(74); xorBitMap(13)(72) := currentData(72); xorBitMap(13)(70) := currentData(70); xorBitMap(13)(69) := currentData(69); xorBitMap(13)(64) := currentData(64); xorBitMap(13)(62) := currentData(62); xorBitMap(13)(60) := currentData(60); xorBitMap(13)(58) := currentData(58); xorBitMap(13)(57) := currentData(57); xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(161) := previousCrc(1); xorBitMap(13)(162) := previousCrc(2); xorBitMap(13)(164) := previousCrc(4); xorBitMap(13)(166) := previousCrc(6); xorBitMap(13)(168) := previousCrc(8); xorBitMap(13)(173) := previousCrc(13); xorBitMap(13)(174) := previousCrc(14); xorBitMap(13)(176) := previousCrc(16); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(179) := previousCrc(19); xorBitMap(13)(180) := previousCrc(20); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(187) := previousCrc(27); xorBitMap(13)(190) := previousCrc(30); xorBitMap(13)(191) := previousCrc(31); 
      xorBitMap(14)(87) := currentData(87); xorBitMap(14)(84) := currentData(84); xorBitMap(14)(83) := currentData(83); xorBitMap(14)(79) := currentData(79); xorBitMap(14)(77) := currentData(77); xorBitMap(14)(76) := currentData(76); xorBitMap(14)(75) := currentData(75); xorBitMap(14)(73) := currentData(73); xorBitMap(14)(71) := currentData(71); xorBitMap(14)(70) := currentData(70); xorBitMap(14)(65) := currentData(65); xorBitMap(14)(63) := currentData(63); xorBitMap(14)(61) := currentData(61); xorBitMap(14)(59) := currentData(59); xorBitMap(14)(58) := currentData(58); xorBitMap(14)(56) := currentData(56); xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(160) := previousCrc(0); xorBitMap(14)(162) := previousCrc(2); xorBitMap(14)(163) := previousCrc(3); xorBitMap(14)(165) := previousCrc(5); xorBitMap(14)(167) := previousCrc(7); xorBitMap(14)(169) := previousCrc(9); xorBitMap(14)(174) := previousCrc(14); xorBitMap(14)(175) := previousCrc(15); xorBitMap(14)(177) := previousCrc(17); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(180) := previousCrc(20); xorBitMap(14)(181) := previousCrc(21); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(188) := previousCrc(28); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(85) := currentData(85); xorBitMap(15)(84) := currentData(84); xorBitMap(15)(80) := currentData(80); xorBitMap(15)(78) := currentData(78); xorBitMap(15)(77) := currentData(77); xorBitMap(15)(76) := currentData(76); xorBitMap(15)(74) := currentData(74); xorBitMap(15)(72) := currentData(72); xorBitMap(15)(71) := currentData(71); xorBitMap(15)(66) := currentData(66); xorBitMap(15)(64) := currentData(64); xorBitMap(15)(62) := currentData(62); xorBitMap(15)(60) := currentData(60); xorBitMap(15)(59) := currentData(59); xorBitMap(15)(57) := currentData(57); xorBitMap(15)(56) := currentData(56); xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(160) := previousCrc(0); xorBitMap(15)(161) := previousCrc(1); xorBitMap(15)(163) := previousCrc(3); xorBitMap(15)(164) := previousCrc(4); xorBitMap(15)(166) := previousCrc(6); xorBitMap(15)(168) := previousCrc(8); xorBitMap(15)(170) := previousCrc(10); xorBitMap(15)(175) := previousCrc(15); xorBitMap(15)(176) := previousCrc(16); xorBitMap(15)(178) := previousCrc(18); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(181) := previousCrc(21); xorBitMap(15)(182) := previousCrc(22); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(189) := previousCrc(29); 
      xorBitMap(16)(87) := currentData(87); xorBitMap(16)(86) := currentData(86); xorBitMap(16)(84) := currentData(84); xorBitMap(16)(83) := currentData(83); xorBitMap(16)(82) := currentData(82); xorBitMap(16)(78) := currentData(78); xorBitMap(16)(77) := currentData(77); xorBitMap(16)(75) := currentData(75); xorBitMap(16)(68) := currentData(68); xorBitMap(16)(66) := currentData(66); xorBitMap(16)(57) := currentData(57); xorBitMap(16)(56) := currentData(56); xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(160) := previousCrc(0); xorBitMap(16)(161) := previousCrc(1); xorBitMap(16)(170) := previousCrc(10); xorBitMap(16)(172) := previousCrc(12); xorBitMap(16)(179) := previousCrc(19); xorBitMap(16)(181) := previousCrc(21); xorBitMap(16)(182) := previousCrc(22); xorBitMap(16)(186) := previousCrc(26); xorBitMap(16)(187) := previousCrc(27); xorBitMap(16)(188) := previousCrc(28); xorBitMap(16)(190) := previousCrc(30); xorBitMap(16)(191) := previousCrc(31); 
      xorBitMap(17)(87) := currentData(87); xorBitMap(17)(85) := currentData(85); xorBitMap(17)(84) := currentData(84); xorBitMap(17)(83) := currentData(83); xorBitMap(17)(79) := currentData(79); xorBitMap(17)(78) := currentData(78); xorBitMap(17)(76) := currentData(76); xorBitMap(17)(69) := currentData(69); xorBitMap(17)(67) := currentData(67); xorBitMap(17)(58) := currentData(58); xorBitMap(17)(57) := currentData(57); xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(161) := previousCrc(1); xorBitMap(17)(162) := previousCrc(2); xorBitMap(17)(171) := previousCrc(11); xorBitMap(17)(173) := previousCrc(13); xorBitMap(17)(180) := previousCrc(20); xorBitMap(17)(182) := previousCrc(22); xorBitMap(17)(183) := previousCrc(23); xorBitMap(17)(187) := previousCrc(27); xorBitMap(17)(188) := previousCrc(28); xorBitMap(17)(189) := previousCrc(29); xorBitMap(17)(191) := previousCrc(31); 
      xorBitMap(18)(86) := currentData(86); xorBitMap(18)(85) := currentData(85); xorBitMap(18)(84) := currentData(84); xorBitMap(18)(80) := currentData(80); xorBitMap(18)(79) := currentData(79); xorBitMap(18)(77) := currentData(77); xorBitMap(18)(70) := currentData(70); xorBitMap(18)(68) := currentData(68); xorBitMap(18)(59) := currentData(59); xorBitMap(18)(58) := currentData(58); xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(162) := previousCrc(2); xorBitMap(18)(163) := previousCrc(3); xorBitMap(18)(172) := previousCrc(12); xorBitMap(18)(174) := previousCrc(14); xorBitMap(18)(181) := previousCrc(21); xorBitMap(18)(183) := previousCrc(23); xorBitMap(18)(184) := previousCrc(24); xorBitMap(18)(188) := previousCrc(28); xorBitMap(18)(189) := previousCrc(29); xorBitMap(18)(190) := previousCrc(30); 
      xorBitMap(19)(87) := currentData(87); xorBitMap(19)(86) := currentData(86); xorBitMap(19)(85) := currentData(85); xorBitMap(19)(81) := currentData(81); xorBitMap(19)(80) := currentData(80); xorBitMap(19)(78) := currentData(78); xorBitMap(19)(71) := currentData(71); xorBitMap(19)(69) := currentData(69); xorBitMap(19)(60) := currentData(60); xorBitMap(19)(59) := currentData(59); xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(163) := previousCrc(3); xorBitMap(19)(164) := previousCrc(4); xorBitMap(19)(173) := previousCrc(13); xorBitMap(19)(175) := previousCrc(15); xorBitMap(19)(182) := previousCrc(22); xorBitMap(19)(184) := previousCrc(24); xorBitMap(19)(185) := previousCrc(25); xorBitMap(19)(189) := previousCrc(29); xorBitMap(19)(190) := previousCrc(30); xorBitMap(19)(191) := previousCrc(31); 
      xorBitMap(20)(87) := currentData(87); xorBitMap(20)(86) := currentData(86); xorBitMap(20)(82) := currentData(82); xorBitMap(20)(81) := currentData(81); xorBitMap(20)(79) := currentData(79); xorBitMap(20)(72) := currentData(72); xorBitMap(20)(70) := currentData(70); xorBitMap(20)(61) := currentData(61); xorBitMap(20)(60) := currentData(60); xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(164) := previousCrc(4); xorBitMap(20)(165) := previousCrc(5); xorBitMap(20)(174) := previousCrc(14); xorBitMap(20)(176) := previousCrc(16); xorBitMap(20)(183) := previousCrc(23); xorBitMap(20)(185) := previousCrc(25); xorBitMap(20)(186) := previousCrc(26); xorBitMap(20)(190) := previousCrc(30); xorBitMap(20)(191) := previousCrc(31); 
      xorBitMap(21)(87) := currentData(87); xorBitMap(21)(83) := currentData(83); xorBitMap(21)(82) := currentData(82); xorBitMap(21)(80) := currentData(80); xorBitMap(21)(73) := currentData(73); xorBitMap(21)(71) := currentData(71); xorBitMap(21)(62) := currentData(62); xorBitMap(21)(61) := currentData(61); xorBitMap(21)(56) := currentData(56); xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(160) := previousCrc(0); xorBitMap(21)(165) := previousCrc(5); xorBitMap(21)(166) := previousCrc(6); xorBitMap(21)(175) := previousCrc(15); xorBitMap(21)(177) := previousCrc(17); xorBitMap(21)(184) := previousCrc(24); xorBitMap(21)(186) := previousCrc(26); xorBitMap(21)(187) := previousCrc(27); xorBitMap(21)(191) := previousCrc(31); 
      xorBitMap(22)(87) := currentData(87); xorBitMap(22)(85) := currentData(85); xorBitMap(22)(82) := currentData(82); xorBitMap(22)(79) := currentData(79); xorBitMap(22)(74) := currentData(74); xorBitMap(22)(73) := currentData(73); xorBitMap(22)(68) := currentData(68); xorBitMap(22)(67) := currentData(67); xorBitMap(22)(66) := currentData(66); xorBitMap(22)(65) := currentData(65); xorBitMap(22)(62) := currentData(62); xorBitMap(22)(61) := currentData(61); xorBitMap(22)(60) := currentData(60); xorBitMap(22)(58) := currentData(58); xorBitMap(22)(57) := currentData(57); xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(161) := previousCrc(1); xorBitMap(22)(162) := previousCrc(2); xorBitMap(22)(164) := previousCrc(4); xorBitMap(22)(165) := previousCrc(5); xorBitMap(22)(166) := previousCrc(6); xorBitMap(22)(169) := previousCrc(9); xorBitMap(22)(170) := previousCrc(10); xorBitMap(22)(171) := previousCrc(11); xorBitMap(22)(172) := previousCrc(12); xorBitMap(22)(177) := previousCrc(17); xorBitMap(22)(178) := previousCrc(18); xorBitMap(22)(183) := previousCrc(23); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(189) := previousCrc(29); xorBitMap(22)(191) := previousCrc(31); 
      xorBitMap(23)(87) := currentData(87); xorBitMap(23)(86) := currentData(86); xorBitMap(23)(85) := currentData(85); xorBitMap(23)(84) := currentData(84); xorBitMap(23)(82) := currentData(82); xorBitMap(23)(81) := currentData(81); xorBitMap(23)(80) := currentData(80); xorBitMap(23)(79) := currentData(79); xorBitMap(23)(75) := currentData(75); xorBitMap(23)(74) := currentData(74); xorBitMap(23)(73) := currentData(73); xorBitMap(23)(72) := currentData(72); xorBitMap(23)(69) := currentData(69); xorBitMap(23)(65) := currentData(65); xorBitMap(23)(62) := currentData(62); xorBitMap(23)(60) := currentData(60); xorBitMap(23)(59) := currentData(59); xorBitMap(23)(56) := currentData(56); xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(160) := previousCrc(0); xorBitMap(23)(163) := previousCrc(3); xorBitMap(23)(164) := previousCrc(4); xorBitMap(23)(166) := previousCrc(6); xorBitMap(23)(169) := previousCrc(9); xorBitMap(23)(173) := previousCrc(13); xorBitMap(23)(176) := previousCrc(16); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(178) := previousCrc(18); xorBitMap(23)(179) := previousCrc(19); xorBitMap(23)(183) := previousCrc(23); xorBitMap(23)(184) := previousCrc(24); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(186) := previousCrc(26); xorBitMap(23)(188) := previousCrc(28); xorBitMap(23)(189) := previousCrc(29); xorBitMap(23)(190) := previousCrc(30); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(87) := currentData(87); xorBitMap(24)(86) := currentData(86); xorBitMap(24)(85) := currentData(85); xorBitMap(24)(83) := currentData(83); xorBitMap(24)(82) := currentData(82); xorBitMap(24)(81) := currentData(81); xorBitMap(24)(80) := currentData(80); xorBitMap(24)(76) := currentData(76); xorBitMap(24)(75) := currentData(75); xorBitMap(24)(74) := currentData(74); xorBitMap(24)(73) := currentData(73); xorBitMap(24)(70) := currentData(70); xorBitMap(24)(66) := currentData(66); xorBitMap(24)(63) := currentData(63); xorBitMap(24)(61) := currentData(61); xorBitMap(24)(60) := currentData(60); xorBitMap(24)(57) := currentData(57); xorBitMap(24)(56) := currentData(56); xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(160) := previousCrc(0); xorBitMap(24)(161) := previousCrc(1); xorBitMap(24)(164) := previousCrc(4); xorBitMap(24)(165) := previousCrc(5); xorBitMap(24)(167) := previousCrc(7); xorBitMap(24)(170) := previousCrc(10); xorBitMap(24)(174) := previousCrc(14); xorBitMap(24)(177) := previousCrc(17); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(179) := previousCrc(19); xorBitMap(24)(180) := previousCrc(20); xorBitMap(24)(184) := previousCrc(24); xorBitMap(24)(185) := previousCrc(25); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(187) := previousCrc(27); xorBitMap(24)(189) := previousCrc(29); xorBitMap(24)(190) := previousCrc(30); xorBitMap(24)(191) := previousCrc(31); 
      xorBitMap(25)(87) := currentData(87); xorBitMap(25)(86) := currentData(86); xorBitMap(25)(84) := currentData(84); xorBitMap(25)(83) := currentData(83); xorBitMap(25)(82) := currentData(82); xorBitMap(25)(81) := currentData(81); xorBitMap(25)(77) := currentData(77); xorBitMap(25)(76) := currentData(76); xorBitMap(25)(75) := currentData(75); xorBitMap(25)(74) := currentData(74); xorBitMap(25)(71) := currentData(71); xorBitMap(25)(67) := currentData(67); xorBitMap(25)(64) := currentData(64); xorBitMap(25)(62) := currentData(62); xorBitMap(25)(61) := currentData(61); xorBitMap(25)(58) := currentData(58); xorBitMap(25)(57) := currentData(57); xorBitMap(25)(56) := currentData(56); xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(160) := previousCrc(0); xorBitMap(25)(161) := previousCrc(1); xorBitMap(25)(162) := previousCrc(2); xorBitMap(25)(165) := previousCrc(5); xorBitMap(25)(166) := previousCrc(6); xorBitMap(25)(168) := previousCrc(8); xorBitMap(25)(171) := previousCrc(11); xorBitMap(25)(175) := previousCrc(15); xorBitMap(25)(178) := previousCrc(18); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(180) := previousCrc(20); xorBitMap(25)(181) := previousCrc(21); xorBitMap(25)(185) := previousCrc(25); xorBitMap(25)(186) := previousCrc(26); xorBitMap(25)(187) := previousCrc(27); xorBitMap(25)(188) := previousCrc(28); xorBitMap(25)(190) := previousCrc(30); xorBitMap(25)(191) := previousCrc(31); 
      xorBitMap(26)(81) := currentData(81); xorBitMap(26)(79) := currentData(79); xorBitMap(26)(78) := currentData(78); xorBitMap(26)(77) := currentData(77); xorBitMap(26)(76) := currentData(76); xorBitMap(26)(75) := currentData(75); xorBitMap(26)(73) := currentData(73); xorBitMap(26)(67) := currentData(67); xorBitMap(26)(66) := currentData(66); xorBitMap(26)(62) := currentData(62); xorBitMap(26)(61) := currentData(61); xorBitMap(26)(60) := currentData(60); xorBitMap(26)(59) := currentData(59); xorBitMap(26)(57) := currentData(57); xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(161) := previousCrc(1); xorBitMap(26)(163) := previousCrc(3); xorBitMap(26)(164) := previousCrc(4); xorBitMap(26)(165) := previousCrc(5); xorBitMap(26)(166) := previousCrc(6); xorBitMap(26)(170) := previousCrc(10); xorBitMap(26)(171) := previousCrc(11); xorBitMap(26)(177) := previousCrc(17); xorBitMap(26)(179) := previousCrc(19); xorBitMap(26)(180) := previousCrc(20); xorBitMap(26)(181) := previousCrc(21); xorBitMap(26)(182) := previousCrc(22); xorBitMap(26)(183) := previousCrc(23); xorBitMap(26)(185) := previousCrc(25); 
      xorBitMap(27)(82) := currentData(82); xorBitMap(27)(80) := currentData(80); xorBitMap(27)(79) := currentData(79); xorBitMap(27)(78) := currentData(78); xorBitMap(27)(77) := currentData(77); xorBitMap(27)(76) := currentData(76); xorBitMap(27)(74) := currentData(74); xorBitMap(27)(68) := currentData(68); xorBitMap(27)(67) := currentData(67); xorBitMap(27)(63) := currentData(63); xorBitMap(27)(62) := currentData(62); xorBitMap(27)(61) := currentData(61); xorBitMap(27)(60) := currentData(60); xorBitMap(27)(58) := currentData(58); xorBitMap(27)(56) := currentData(56); xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(160) := previousCrc(0); xorBitMap(27)(162) := previousCrc(2); xorBitMap(27)(164) := previousCrc(4); xorBitMap(27)(165) := previousCrc(5); xorBitMap(27)(166) := previousCrc(6); xorBitMap(27)(167) := previousCrc(7); xorBitMap(27)(171) := previousCrc(11); xorBitMap(27)(172) := previousCrc(12); xorBitMap(27)(178) := previousCrc(18); xorBitMap(27)(180) := previousCrc(20); xorBitMap(27)(181) := previousCrc(21); xorBitMap(27)(182) := previousCrc(22); xorBitMap(27)(183) := previousCrc(23); xorBitMap(27)(184) := previousCrc(24); xorBitMap(27)(186) := previousCrc(26); 
      xorBitMap(28)(83) := currentData(83); xorBitMap(28)(81) := currentData(81); xorBitMap(28)(80) := currentData(80); xorBitMap(28)(79) := currentData(79); xorBitMap(28)(78) := currentData(78); xorBitMap(28)(77) := currentData(77); xorBitMap(28)(75) := currentData(75); xorBitMap(28)(69) := currentData(69); xorBitMap(28)(68) := currentData(68); xorBitMap(28)(64) := currentData(64); xorBitMap(28)(63) := currentData(63); xorBitMap(28)(62) := currentData(62); xorBitMap(28)(61) := currentData(61); xorBitMap(28)(59) := currentData(59); xorBitMap(28)(57) := currentData(57); xorBitMap(28)(56) := currentData(56); xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(160) := previousCrc(0); xorBitMap(28)(161) := previousCrc(1); xorBitMap(28)(163) := previousCrc(3); xorBitMap(28)(165) := previousCrc(5); xorBitMap(28)(166) := previousCrc(6); xorBitMap(28)(167) := previousCrc(7); xorBitMap(28)(168) := previousCrc(8); xorBitMap(28)(172) := previousCrc(12); xorBitMap(28)(173) := previousCrc(13); xorBitMap(28)(179) := previousCrc(19); xorBitMap(28)(181) := previousCrc(21); xorBitMap(28)(182) := previousCrc(22); xorBitMap(28)(183) := previousCrc(23); xorBitMap(28)(184) := previousCrc(24); xorBitMap(28)(185) := previousCrc(25); xorBitMap(28)(187) := previousCrc(27); 
      xorBitMap(29)(84) := currentData(84); xorBitMap(29)(82) := currentData(82); xorBitMap(29)(81) := currentData(81); xorBitMap(29)(80) := currentData(80); xorBitMap(29)(79) := currentData(79); xorBitMap(29)(78) := currentData(78); xorBitMap(29)(76) := currentData(76); xorBitMap(29)(70) := currentData(70); xorBitMap(29)(69) := currentData(69); xorBitMap(29)(65) := currentData(65); xorBitMap(29)(64) := currentData(64); xorBitMap(29)(63) := currentData(63); xorBitMap(29)(62) := currentData(62); xorBitMap(29)(60) := currentData(60); xorBitMap(29)(58) := currentData(58); xorBitMap(29)(57) := currentData(57); xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(161) := previousCrc(1); xorBitMap(29)(162) := previousCrc(2); xorBitMap(29)(164) := previousCrc(4); xorBitMap(29)(166) := previousCrc(6); xorBitMap(29)(167) := previousCrc(7); xorBitMap(29)(168) := previousCrc(8); xorBitMap(29)(169) := previousCrc(9); xorBitMap(29)(173) := previousCrc(13); xorBitMap(29)(174) := previousCrc(14); xorBitMap(29)(180) := previousCrc(20); xorBitMap(29)(182) := previousCrc(22); xorBitMap(29)(183) := previousCrc(23); xorBitMap(29)(184) := previousCrc(24); xorBitMap(29)(185) := previousCrc(25); xorBitMap(29)(186) := previousCrc(26); xorBitMap(29)(188) := previousCrc(28); 
      xorBitMap(30)(85) := currentData(85); xorBitMap(30)(83) := currentData(83); xorBitMap(30)(82) := currentData(82); xorBitMap(30)(81) := currentData(81); xorBitMap(30)(80) := currentData(80); xorBitMap(30)(79) := currentData(79); xorBitMap(30)(77) := currentData(77); xorBitMap(30)(71) := currentData(71); xorBitMap(30)(70) := currentData(70); xorBitMap(30)(66) := currentData(66); xorBitMap(30)(65) := currentData(65); xorBitMap(30)(64) := currentData(64); xorBitMap(30)(63) := currentData(63); xorBitMap(30)(61) := currentData(61); xorBitMap(30)(59) := currentData(59); xorBitMap(30)(58) := currentData(58); xorBitMap(30)(56) := currentData(56); xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(160) := previousCrc(0); xorBitMap(30)(162) := previousCrc(2); xorBitMap(30)(163) := previousCrc(3); xorBitMap(30)(165) := previousCrc(5); xorBitMap(30)(167) := previousCrc(7); xorBitMap(30)(168) := previousCrc(8); xorBitMap(30)(169) := previousCrc(9); xorBitMap(30)(170) := previousCrc(10); xorBitMap(30)(174) := previousCrc(14); xorBitMap(30)(175) := previousCrc(15); xorBitMap(30)(181) := previousCrc(21); xorBitMap(30)(183) := previousCrc(23); xorBitMap(30)(184) := previousCrc(24); xorBitMap(30)(185) := previousCrc(25); xorBitMap(30)(186) := previousCrc(26); xorBitMap(30)(187) := previousCrc(27); xorBitMap(30)(189) := previousCrc(29); 
      xorBitMap(31)(86) := currentData(86); xorBitMap(31)(84) := currentData(84); xorBitMap(31)(83) := currentData(83); xorBitMap(31)(82) := currentData(82); xorBitMap(31)(81) := currentData(81); xorBitMap(31)(80) := currentData(80); xorBitMap(31)(78) := currentData(78); xorBitMap(31)(72) := currentData(72); xorBitMap(31)(71) := currentData(71); xorBitMap(31)(67) := currentData(67); xorBitMap(31)(66) := currentData(66); xorBitMap(31)(65) := currentData(65); xorBitMap(31)(64) := currentData(64); xorBitMap(31)(62) := currentData(62); xorBitMap(31)(60) := currentData(60); xorBitMap(31)(59) := currentData(59); xorBitMap(31)(57) := currentData(57); xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(161) := previousCrc(1); xorBitMap(31)(163) := previousCrc(3); xorBitMap(31)(164) := previousCrc(4); xorBitMap(31)(166) := previousCrc(6); xorBitMap(31)(168) := previousCrc(8); xorBitMap(31)(169) := previousCrc(9); xorBitMap(31)(170) := previousCrc(10); xorBitMap(31)(171) := previousCrc(11); xorBitMap(31)(175) := previousCrc(15); xorBitMap(31)(176) := previousCrc(16); xorBitMap(31)(182) := previousCrc(22); xorBitMap(31)(184) := previousCrc(24); xorBitMap(31)(185) := previousCrc(25); xorBitMap(31)(186) := previousCrc(26); xorBitMap(31)(187) := previousCrc(27); xorBitMap(31)(188) := previousCrc(28); xorBitMap(31)(190) := previousCrc(30); 
   end procedure;

   procedure xorBitMap12Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(95 downto 0)) is 
   begin
      xorBitMap(0)(95) := currentData(95); xorBitMap(0)(94) := currentData(94); xorBitMap(0)(87) := currentData(87); xorBitMap(0)(85) := currentData(85); xorBitMap(0)(84) := currentData(84); xorBitMap(0)(83) := currentData(83); xorBitMap(0)(82) := currentData(82); xorBitMap(0)(81) := currentData(81); xorBitMap(0)(79) := currentData(79); xorBitMap(0)(73) := currentData(73); xorBitMap(0)(72) := currentData(72); xorBitMap(0)(68) := currentData(68); xorBitMap(0)(67) := currentData(67); xorBitMap(0)(66) := currentData(66); xorBitMap(0)(65) := currentData(65); xorBitMap(0)(63) := currentData(63); xorBitMap(0)(61) := currentData(61); xorBitMap(0)(60) := currentData(60); xorBitMap(0)(58) := currentData(58); xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(161) := previousCrc(1); xorBitMap(0)(162) := previousCrc(2); xorBitMap(0)(163) := previousCrc(3); xorBitMap(0)(164) := previousCrc(4); xorBitMap(0)(168) := previousCrc(8); xorBitMap(0)(169) := previousCrc(9); xorBitMap(0)(175) := previousCrc(15); xorBitMap(0)(177) := previousCrc(17); xorBitMap(0)(178) := previousCrc(18); xorBitMap(0)(179) := previousCrc(19); xorBitMap(0)(180) := previousCrc(20); xorBitMap(0)(181) := previousCrc(21); xorBitMap(0)(183) := previousCrc(23); xorBitMap(0)(190) := previousCrc(30); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(94) := currentData(94); xorBitMap(1)(88) := currentData(88); xorBitMap(1)(87) := currentData(87); xorBitMap(1)(86) := currentData(86); xorBitMap(1)(81) := currentData(81); xorBitMap(1)(80) := currentData(80); xorBitMap(1)(79) := currentData(79); xorBitMap(1)(74) := currentData(74); xorBitMap(1)(72) := currentData(72); xorBitMap(1)(69) := currentData(69); xorBitMap(1)(65) := currentData(65); xorBitMap(1)(64) := currentData(64); xorBitMap(1)(63) := currentData(63); xorBitMap(1)(62) := currentData(62); xorBitMap(1)(60) := currentData(60); xorBitMap(1)(59) := currentData(59); xorBitMap(1)(58) := currentData(58); xorBitMap(1)(56) := currentData(56); xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(160) := previousCrc(0); xorBitMap(1)(161) := previousCrc(1); xorBitMap(1)(165) := previousCrc(5); xorBitMap(1)(168) := previousCrc(8); xorBitMap(1)(170) := previousCrc(10); xorBitMap(1)(175) := previousCrc(15); xorBitMap(1)(176) := previousCrc(16); xorBitMap(1)(177) := previousCrc(17); xorBitMap(1)(182) := previousCrc(22); xorBitMap(1)(183) := previousCrc(23); xorBitMap(1)(184) := previousCrc(24); xorBitMap(1)(190) := previousCrc(30); 
      xorBitMap(2)(94) := currentData(94); xorBitMap(2)(89) := currentData(89); xorBitMap(2)(88) := currentData(88); xorBitMap(2)(85) := currentData(85); xorBitMap(2)(84) := currentData(84); xorBitMap(2)(83) := currentData(83); xorBitMap(2)(80) := currentData(80); xorBitMap(2)(79) := currentData(79); xorBitMap(2)(75) := currentData(75); xorBitMap(2)(72) := currentData(72); xorBitMap(2)(70) := currentData(70); xorBitMap(2)(68) := currentData(68); xorBitMap(2)(67) := currentData(67); xorBitMap(2)(64) := currentData(64); xorBitMap(2)(59) := currentData(59); xorBitMap(2)(58) := currentData(58); xorBitMap(2)(57) := currentData(57); xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(160) := previousCrc(0); xorBitMap(2)(163) := previousCrc(3); xorBitMap(2)(164) := previousCrc(4); xorBitMap(2)(166) := previousCrc(6); xorBitMap(2)(168) := previousCrc(8); xorBitMap(2)(171) := previousCrc(11); xorBitMap(2)(175) := previousCrc(15); xorBitMap(2)(176) := previousCrc(16); xorBitMap(2)(179) := previousCrc(19); xorBitMap(2)(180) := previousCrc(20); xorBitMap(2)(181) := previousCrc(21); xorBitMap(2)(184) := previousCrc(24); xorBitMap(2)(185) := previousCrc(25); xorBitMap(2)(190) := previousCrc(30); 
      xorBitMap(3)(95) := currentData(95); xorBitMap(3)(90) := currentData(90); xorBitMap(3)(89) := currentData(89); xorBitMap(3)(86) := currentData(86); xorBitMap(3)(85) := currentData(85); xorBitMap(3)(84) := currentData(84); xorBitMap(3)(81) := currentData(81); xorBitMap(3)(80) := currentData(80); xorBitMap(3)(76) := currentData(76); xorBitMap(3)(73) := currentData(73); xorBitMap(3)(71) := currentData(71); xorBitMap(3)(69) := currentData(69); xorBitMap(3)(68) := currentData(68); xorBitMap(3)(65) := currentData(65); xorBitMap(3)(60) := currentData(60); xorBitMap(3)(59) := currentData(59); xorBitMap(3)(58) := currentData(58); xorBitMap(3)(56) := currentData(56); xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(161) := previousCrc(1); xorBitMap(3)(164) := previousCrc(4); xorBitMap(3)(165) := previousCrc(5); xorBitMap(3)(167) := previousCrc(7); xorBitMap(3)(169) := previousCrc(9); xorBitMap(3)(172) := previousCrc(12); xorBitMap(3)(176) := previousCrc(16); xorBitMap(3)(177) := previousCrc(17); xorBitMap(3)(180) := previousCrc(20); xorBitMap(3)(181) := previousCrc(21); xorBitMap(3)(182) := previousCrc(22); xorBitMap(3)(185) := previousCrc(25); xorBitMap(3)(186) := previousCrc(26); xorBitMap(3)(191) := previousCrc(31); 
      xorBitMap(4)(95) := currentData(95); xorBitMap(4)(94) := currentData(94); xorBitMap(4)(91) := currentData(91); xorBitMap(4)(90) := currentData(90); xorBitMap(4)(86) := currentData(86); xorBitMap(4)(84) := currentData(84); xorBitMap(4)(83) := currentData(83); xorBitMap(4)(79) := currentData(79); xorBitMap(4)(77) := currentData(77); xorBitMap(4)(74) := currentData(74); xorBitMap(4)(73) := currentData(73); xorBitMap(4)(70) := currentData(70); xorBitMap(4)(69) := currentData(69); xorBitMap(4)(68) := currentData(68); xorBitMap(4)(67) := currentData(67); xorBitMap(4)(65) := currentData(65); xorBitMap(4)(63) := currentData(63); xorBitMap(4)(59) := currentData(59); xorBitMap(4)(58) := currentData(58); xorBitMap(4)(57) := currentData(57); xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(161) := previousCrc(1); xorBitMap(4)(163) := previousCrc(3); xorBitMap(4)(164) := previousCrc(4); xorBitMap(4)(165) := previousCrc(5); xorBitMap(4)(166) := previousCrc(6); xorBitMap(4)(169) := previousCrc(9); xorBitMap(4)(170) := previousCrc(10); xorBitMap(4)(173) := previousCrc(13); xorBitMap(4)(175) := previousCrc(15); xorBitMap(4)(179) := previousCrc(19); xorBitMap(4)(180) := previousCrc(20); xorBitMap(4)(182) := previousCrc(22); xorBitMap(4)(186) := previousCrc(26); xorBitMap(4)(187) := previousCrc(27); xorBitMap(4)(190) := previousCrc(30); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(94) := currentData(94); xorBitMap(5)(92) := currentData(92); xorBitMap(5)(91) := currentData(91); xorBitMap(5)(83) := currentData(83); xorBitMap(5)(82) := currentData(82); xorBitMap(5)(81) := currentData(81); xorBitMap(5)(80) := currentData(80); xorBitMap(5)(79) := currentData(79); xorBitMap(5)(78) := currentData(78); xorBitMap(5)(75) := currentData(75); xorBitMap(5)(74) := currentData(74); xorBitMap(5)(73) := currentData(73); xorBitMap(5)(72) := currentData(72); xorBitMap(5)(71) := currentData(71); xorBitMap(5)(70) := currentData(70); xorBitMap(5)(69) := currentData(69); xorBitMap(5)(67) := currentData(67); xorBitMap(5)(65) := currentData(65); xorBitMap(5)(64) := currentData(64); xorBitMap(5)(63) := currentData(63); xorBitMap(5)(61) := currentData(61); xorBitMap(5)(59) := currentData(59); xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(160) := previousCrc(0); xorBitMap(5)(161) := previousCrc(1); xorBitMap(5)(163) := previousCrc(3); xorBitMap(5)(165) := previousCrc(5); xorBitMap(5)(166) := previousCrc(6); xorBitMap(5)(167) := previousCrc(7); xorBitMap(5)(168) := previousCrc(8); xorBitMap(5)(169) := previousCrc(9); xorBitMap(5)(170) := previousCrc(10); xorBitMap(5)(171) := previousCrc(11); xorBitMap(5)(174) := previousCrc(14); xorBitMap(5)(175) := previousCrc(15); xorBitMap(5)(176) := previousCrc(16); xorBitMap(5)(177) := previousCrc(17); xorBitMap(5)(178) := previousCrc(18); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(188) := previousCrc(28); xorBitMap(5)(190) := previousCrc(30); 
      xorBitMap(6)(95) := currentData(95); xorBitMap(6)(93) := currentData(93); xorBitMap(6)(92) := currentData(92); xorBitMap(6)(84) := currentData(84); xorBitMap(6)(83) := currentData(83); xorBitMap(6)(82) := currentData(82); xorBitMap(6)(81) := currentData(81); xorBitMap(6)(80) := currentData(80); xorBitMap(6)(79) := currentData(79); xorBitMap(6)(76) := currentData(76); xorBitMap(6)(75) := currentData(75); xorBitMap(6)(74) := currentData(74); xorBitMap(6)(73) := currentData(73); xorBitMap(6)(72) := currentData(72); xorBitMap(6)(71) := currentData(71); xorBitMap(6)(70) := currentData(70); xorBitMap(6)(68) := currentData(68); xorBitMap(6)(66) := currentData(66); xorBitMap(6)(65) := currentData(65); xorBitMap(6)(64) := currentData(64); xorBitMap(6)(62) := currentData(62); xorBitMap(6)(60) := currentData(60); xorBitMap(6)(56) := currentData(56); xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(160) := previousCrc(0); xorBitMap(6)(161) := previousCrc(1); xorBitMap(6)(162) := previousCrc(2); xorBitMap(6)(164) := previousCrc(4); xorBitMap(6)(166) := previousCrc(6); xorBitMap(6)(167) := previousCrc(7); xorBitMap(6)(168) := previousCrc(8); xorBitMap(6)(169) := previousCrc(9); xorBitMap(6)(170) := previousCrc(10); xorBitMap(6)(171) := previousCrc(11); xorBitMap(6)(172) := previousCrc(12); xorBitMap(6)(175) := previousCrc(15); xorBitMap(6)(176) := previousCrc(16); xorBitMap(6)(177) := previousCrc(17); xorBitMap(6)(178) := previousCrc(18); xorBitMap(6)(179) := previousCrc(19); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(188) := previousCrc(28); xorBitMap(6)(189) := previousCrc(29); xorBitMap(6)(191) := previousCrc(31); 
      xorBitMap(7)(95) := currentData(95); xorBitMap(7)(93) := currentData(93); xorBitMap(7)(87) := currentData(87); xorBitMap(7)(80) := currentData(80); xorBitMap(7)(79) := currentData(79); xorBitMap(7)(77) := currentData(77); xorBitMap(7)(76) := currentData(76); xorBitMap(7)(75) := currentData(75); xorBitMap(7)(74) := currentData(74); xorBitMap(7)(71) := currentData(71); xorBitMap(7)(69) := currentData(69); xorBitMap(7)(68) := currentData(68); xorBitMap(7)(60) := currentData(60); xorBitMap(7)(58) := currentData(58); xorBitMap(7)(57) := currentData(57); xorBitMap(7)(56) := currentData(56); xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(164) := previousCrc(4); xorBitMap(7)(165) := previousCrc(5); xorBitMap(7)(167) := previousCrc(7); xorBitMap(7)(170) := previousCrc(10); xorBitMap(7)(171) := previousCrc(11); xorBitMap(7)(172) := previousCrc(12); xorBitMap(7)(173) := previousCrc(13); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(176) := previousCrc(16); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(189) := previousCrc(29); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(95) := currentData(95); xorBitMap(8)(88) := currentData(88); xorBitMap(8)(87) := currentData(87); xorBitMap(8)(85) := currentData(85); xorBitMap(8)(84) := currentData(84); xorBitMap(8)(83) := currentData(83); xorBitMap(8)(82) := currentData(82); xorBitMap(8)(80) := currentData(80); xorBitMap(8)(79) := currentData(79); xorBitMap(8)(78) := currentData(78); xorBitMap(8)(77) := currentData(77); xorBitMap(8)(76) := currentData(76); xorBitMap(8)(75) := currentData(75); xorBitMap(8)(73) := currentData(73); xorBitMap(8)(70) := currentData(70); xorBitMap(8)(69) := currentData(69); xorBitMap(8)(68) := currentData(68); xorBitMap(8)(67) := currentData(67); xorBitMap(8)(66) := currentData(66); xorBitMap(8)(65) := currentData(65); xorBitMap(8)(63) := currentData(63); xorBitMap(8)(60) := currentData(60); xorBitMap(8)(59) := currentData(59); xorBitMap(8)(57) := currentData(57); xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(161) := previousCrc(1); xorBitMap(8)(162) := previousCrc(2); xorBitMap(8)(163) := previousCrc(3); xorBitMap(8)(164) := previousCrc(4); xorBitMap(8)(165) := previousCrc(5); xorBitMap(8)(166) := previousCrc(6); xorBitMap(8)(169) := previousCrc(9); xorBitMap(8)(171) := previousCrc(11); xorBitMap(8)(172) := previousCrc(12); xorBitMap(8)(173) := previousCrc(13); xorBitMap(8)(174) := previousCrc(14); xorBitMap(8)(175) := previousCrc(15); xorBitMap(8)(176) := previousCrc(16); xorBitMap(8)(178) := previousCrc(18); xorBitMap(8)(179) := previousCrc(19); xorBitMap(8)(180) := previousCrc(20); xorBitMap(8)(181) := previousCrc(21); xorBitMap(8)(183) := previousCrc(23); xorBitMap(8)(184) := previousCrc(24); xorBitMap(8)(191) := previousCrc(31); 
      xorBitMap(9)(89) := currentData(89); xorBitMap(9)(88) := currentData(88); xorBitMap(9)(86) := currentData(86); xorBitMap(9)(85) := currentData(85); xorBitMap(9)(84) := currentData(84); xorBitMap(9)(83) := currentData(83); xorBitMap(9)(81) := currentData(81); xorBitMap(9)(80) := currentData(80); xorBitMap(9)(79) := currentData(79); xorBitMap(9)(78) := currentData(78); xorBitMap(9)(77) := currentData(77); xorBitMap(9)(76) := currentData(76); xorBitMap(9)(74) := currentData(74); xorBitMap(9)(71) := currentData(71); xorBitMap(9)(70) := currentData(70); xorBitMap(9)(69) := currentData(69); xorBitMap(9)(68) := currentData(68); xorBitMap(9)(67) := currentData(67); xorBitMap(9)(66) := currentData(66); xorBitMap(9)(64) := currentData(64); xorBitMap(9)(61) := currentData(61); xorBitMap(9)(60) := currentData(60); xorBitMap(9)(58) := currentData(58); xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(160) := previousCrc(0); xorBitMap(9)(162) := previousCrc(2); xorBitMap(9)(163) := previousCrc(3); xorBitMap(9)(164) := previousCrc(4); xorBitMap(9)(165) := previousCrc(5); xorBitMap(9)(166) := previousCrc(6); xorBitMap(9)(167) := previousCrc(7); xorBitMap(9)(170) := previousCrc(10); xorBitMap(9)(172) := previousCrc(12); xorBitMap(9)(173) := previousCrc(13); xorBitMap(9)(174) := previousCrc(14); xorBitMap(9)(175) := previousCrc(15); xorBitMap(9)(176) := previousCrc(16); xorBitMap(9)(177) := previousCrc(17); xorBitMap(9)(179) := previousCrc(19); xorBitMap(9)(180) := previousCrc(20); xorBitMap(9)(181) := previousCrc(21); xorBitMap(9)(182) := previousCrc(22); xorBitMap(9)(184) := previousCrc(24); xorBitMap(9)(185) := previousCrc(25); 
      xorBitMap(10)(95) := currentData(95); xorBitMap(10)(94) := currentData(94); xorBitMap(10)(90) := currentData(90); xorBitMap(10)(89) := currentData(89); xorBitMap(10)(86) := currentData(86); xorBitMap(10)(83) := currentData(83); xorBitMap(10)(80) := currentData(80); xorBitMap(10)(78) := currentData(78); xorBitMap(10)(77) := currentData(77); xorBitMap(10)(75) := currentData(75); xorBitMap(10)(73) := currentData(73); xorBitMap(10)(71) := currentData(71); xorBitMap(10)(70) := currentData(70); xorBitMap(10)(69) := currentData(69); xorBitMap(10)(66) := currentData(66); xorBitMap(10)(63) := currentData(63); xorBitMap(10)(62) := currentData(62); xorBitMap(10)(60) := currentData(60); xorBitMap(10)(59) := currentData(59); xorBitMap(10)(58) := currentData(58); xorBitMap(10)(56) := currentData(56); xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(162) := previousCrc(2); xorBitMap(10)(165) := previousCrc(5); xorBitMap(10)(166) := previousCrc(6); xorBitMap(10)(167) := previousCrc(7); xorBitMap(10)(169) := previousCrc(9); xorBitMap(10)(171) := previousCrc(11); xorBitMap(10)(173) := previousCrc(13); xorBitMap(10)(174) := previousCrc(14); xorBitMap(10)(176) := previousCrc(16); xorBitMap(10)(179) := previousCrc(19); xorBitMap(10)(182) := previousCrc(22); xorBitMap(10)(185) := previousCrc(25); xorBitMap(10)(186) := previousCrc(26); xorBitMap(10)(190) := previousCrc(30); xorBitMap(10)(191) := previousCrc(31); 
      xorBitMap(11)(94) := currentData(94); xorBitMap(11)(91) := currentData(91); xorBitMap(11)(90) := currentData(90); xorBitMap(11)(85) := currentData(85); xorBitMap(11)(83) := currentData(83); xorBitMap(11)(82) := currentData(82); xorBitMap(11)(78) := currentData(78); xorBitMap(11)(76) := currentData(76); xorBitMap(11)(74) := currentData(74); xorBitMap(11)(73) := currentData(73); xorBitMap(11)(71) := currentData(71); xorBitMap(11)(70) := currentData(70); xorBitMap(11)(68) := currentData(68); xorBitMap(11)(66) := currentData(66); xorBitMap(11)(65) := currentData(65); xorBitMap(11)(64) := currentData(64); xorBitMap(11)(59) := currentData(59); xorBitMap(11)(58) := currentData(58); xorBitMap(11)(57) := currentData(57); xorBitMap(11)(56) := currentData(56); xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(160) := previousCrc(0); xorBitMap(11)(161) := previousCrc(1); xorBitMap(11)(162) := previousCrc(2); xorBitMap(11)(164) := previousCrc(4); xorBitMap(11)(166) := previousCrc(6); xorBitMap(11)(167) := previousCrc(7); xorBitMap(11)(169) := previousCrc(9); xorBitMap(11)(170) := previousCrc(10); xorBitMap(11)(172) := previousCrc(12); xorBitMap(11)(174) := previousCrc(14); xorBitMap(11)(178) := previousCrc(18); xorBitMap(11)(179) := previousCrc(19); xorBitMap(11)(181) := previousCrc(21); xorBitMap(11)(186) := previousCrc(26); xorBitMap(11)(187) := previousCrc(27); xorBitMap(11)(190) := previousCrc(30); 
      xorBitMap(12)(94) := currentData(94); xorBitMap(12)(92) := currentData(92); xorBitMap(12)(91) := currentData(91); xorBitMap(12)(87) := currentData(87); xorBitMap(12)(86) := currentData(86); xorBitMap(12)(85) := currentData(85); xorBitMap(12)(82) := currentData(82); xorBitMap(12)(81) := currentData(81); xorBitMap(12)(77) := currentData(77); xorBitMap(12)(75) := currentData(75); xorBitMap(12)(74) := currentData(74); xorBitMap(12)(73) := currentData(73); xorBitMap(12)(71) := currentData(71); xorBitMap(12)(69) := currentData(69); xorBitMap(12)(68) := currentData(68); xorBitMap(12)(63) := currentData(63); xorBitMap(12)(61) := currentData(61); xorBitMap(12)(59) := currentData(59); xorBitMap(12)(57) := currentData(57); xorBitMap(12)(56) := currentData(56); xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(164) := previousCrc(4); xorBitMap(12)(165) := previousCrc(5); xorBitMap(12)(167) := previousCrc(7); xorBitMap(12)(169) := previousCrc(9); xorBitMap(12)(170) := previousCrc(10); xorBitMap(12)(171) := previousCrc(11); xorBitMap(12)(173) := previousCrc(13); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(178) := previousCrc(18); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(182) := previousCrc(22); xorBitMap(12)(183) := previousCrc(23); xorBitMap(12)(187) := previousCrc(27); xorBitMap(12)(188) := previousCrc(28); xorBitMap(12)(190) := previousCrc(30); 
      xorBitMap(13)(95) := currentData(95); xorBitMap(13)(93) := currentData(93); xorBitMap(13)(92) := currentData(92); xorBitMap(13)(88) := currentData(88); xorBitMap(13)(87) := currentData(87); xorBitMap(13)(86) := currentData(86); xorBitMap(13)(83) := currentData(83); xorBitMap(13)(82) := currentData(82); xorBitMap(13)(78) := currentData(78); xorBitMap(13)(76) := currentData(76); xorBitMap(13)(75) := currentData(75); xorBitMap(13)(74) := currentData(74); xorBitMap(13)(72) := currentData(72); xorBitMap(13)(70) := currentData(70); xorBitMap(13)(69) := currentData(69); xorBitMap(13)(64) := currentData(64); xorBitMap(13)(62) := currentData(62); xorBitMap(13)(60) := currentData(60); xorBitMap(13)(58) := currentData(58); xorBitMap(13)(57) := currentData(57); xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(160) := previousCrc(0); xorBitMap(13)(165) := previousCrc(5); xorBitMap(13)(166) := previousCrc(6); xorBitMap(13)(168) := previousCrc(8); xorBitMap(13)(170) := previousCrc(10); xorBitMap(13)(171) := previousCrc(11); xorBitMap(13)(172) := previousCrc(12); xorBitMap(13)(174) := previousCrc(14); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(179) := previousCrc(19); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(183) := previousCrc(23); xorBitMap(13)(184) := previousCrc(24); xorBitMap(13)(188) := previousCrc(28); xorBitMap(13)(189) := previousCrc(29); xorBitMap(13)(191) := previousCrc(31); 
      xorBitMap(14)(94) := currentData(94); xorBitMap(14)(93) := currentData(93); xorBitMap(14)(89) := currentData(89); xorBitMap(14)(88) := currentData(88); xorBitMap(14)(87) := currentData(87); xorBitMap(14)(84) := currentData(84); xorBitMap(14)(83) := currentData(83); xorBitMap(14)(79) := currentData(79); xorBitMap(14)(77) := currentData(77); xorBitMap(14)(76) := currentData(76); xorBitMap(14)(75) := currentData(75); xorBitMap(14)(73) := currentData(73); xorBitMap(14)(71) := currentData(71); xorBitMap(14)(70) := currentData(70); xorBitMap(14)(65) := currentData(65); xorBitMap(14)(63) := currentData(63); xorBitMap(14)(61) := currentData(61); xorBitMap(14)(59) := currentData(59); xorBitMap(14)(58) := currentData(58); xorBitMap(14)(56) := currentData(56); xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(161) := previousCrc(1); xorBitMap(14)(166) := previousCrc(6); xorBitMap(14)(167) := previousCrc(7); xorBitMap(14)(169) := previousCrc(9); xorBitMap(14)(171) := previousCrc(11); xorBitMap(14)(172) := previousCrc(12); xorBitMap(14)(173) := previousCrc(13); xorBitMap(14)(175) := previousCrc(15); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(180) := previousCrc(20); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(184) := previousCrc(24); xorBitMap(14)(185) := previousCrc(25); xorBitMap(14)(189) := previousCrc(29); xorBitMap(14)(190) := previousCrc(30); 
      xorBitMap(15)(95) := currentData(95); xorBitMap(15)(94) := currentData(94); xorBitMap(15)(90) := currentData(90); xorBitMap(15)(89) := currentData(89); xorBitMap(15)(88) := currentData(88); xorBitMap(15)(85) := currentData(85); xorBitMap(15)(84) := currentData(84); xorBitMap(15)(80) := currentData(80); xorBitMap(15)(78) := currentData(78); xorBitMap(15)(77) := currentData(77); xorBitMap(15)(76) := currentData(76); xorBitMap(15)(74) := currentData(74); xorBitMap(15)(72) := currentData(72); xorBitMap(15)(71) := currentData(71); xorBitMap(15)(66) := currentData(66); xorBitMap(15)(64) := currentData(64); xorBitMap(15)(62) := currentData(62); xorBitMap(15)(60) := currentData(60); xorBitMap(15)(59) := currentData(59); xorBitMap(15)(57) := currentData(57); xorBitMap(15)(56) := currentData(56); xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(160) := previousCrc(0); xorBitMap(15)(162) := previousCrc(2); xorBitMap(15)(167) := previousCrc(7); xorBitMap(15)(168) := previousCrc(8); xorBitMap(15)(170) := previousCrc(10); xorBitMap(15)(172) := previousCrc(12); xorBitMap(15)(173) := previousCrc(13); xorBitMap(15)(174) := previousCrc(14); xorBitMap(15)(176) := previousCrc(16); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(181) := previousCrc(21); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(185) := previousCrc(25); xorBitMap(15)(186) := previousCrc(26); xorBitMap(15)(190) := previousCrc(30); xorBitMap(15)(191) := previousCrc(31); 
      xorBitMap(16)(94) := currentData(94); xorBitMap(16)(91) := currentData(91); xorBitMap(16)(90) := currentData(90); xorBitMap(16)(89) := currentData(89); xorBitMap(16)(87) := currentData(87); xorBitMap(16)(86) := currentData(86); xorBitMap(16)(84) := currentData(84); xorBitMap(16)(83) := currentData(83); xorBitMap(16)(82) := currentData(82); xorBitMap(16)(78) := currentData(78); xorBitMap(16)(77) := currentData(77); xorBitMap(16)(75) := currentData(75); xorBitMap(16)(68) := currentData(68); xorBitMap(16)(66) := currentData(66); xorBitMap(16)(57) := currentData(57); xorBitMap(16)(56) := currentData(56); xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(162) := previousCrc(2); xorBitMap(16)(164) := previousCrc(4); xorBitMap(16)(171) := previousCrc(11); xorBitMap(16)(173) := previousCrc(13); xorBitMap(16)(174) := previousCrc(14); xorBitMap(16)(178) := previousCrc(18); xorBitMap(16)(179) := previousCrc(19); xorBitMap(16)(180) := previousCrc(20); xorBitMap(16)(182) := previousCrc(22); xorBitMap(16)(183) := previousCrc(23); xorBitMap(16)(185) := previousCrc(25); xorBitMap(16)(186) := previousCrc(26); xorBitMap(16)(187) := previousCrc(27); xorBitMap(16)(190) := previousCrc(30); 
      xorBitMap(17)(95) := currentData(95); xorBitMap(17)(92) := currentData(92); xorBitMap(17)(91) := currentData(91); xorBitMap(17)(90) := currentData(90); xorBitMap(17)(88) := currentData(88); xorBitMap(17)(87) := currentData(87); xorBitMap(17)(85) := currentData(85); xorBitMap(17)(84) := currentData(84); xorBitMap(17)(83) := currentData(83); xorBitMap(17)(79) := currentData(79); xorBitMap(17)(78) := currentData(78); xorBitMap(17)(76) := currentData(76); xorBitMap(17)(69) := currentData(69); xorBitMap(17)(67) := currentData(67); xorBitMap(17)(58) := currentData(58); xorBitMap(17)(57) := currentData(57); xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(163) := previousCrc(3); xorBitMap(17)(165) := previousCrc(5); xorBitMap(17)(172) := previousCrc(12); xorBitMap(17)(174) := previousCrc(14); xorBitMap(17)(175) := previousCrc(15); xorBitMap(17)(179) := previousCrc(19); xorBitMap(17)(180) := previousCrc(20); xorBitMap(17)(181) := previousCrc(21); xorBitMap(17)(183) := previousCrc(23); xorBitMap(17)(184) := previousCrc(24); xorBitMap(17)(186) := previousCrc(26); xorBitMap(17)(187) := previousCrc(27); xorBitMap(17)(188) := previousCrc(28); xorBitMap(17)(191) := previousCrc(31); 
      xorBitMap(18)(93) := currentData(93); xorBitMap(18)(92) := currentData(92); xorBitMap(18)(91) := currentData(91); xorBitMap(18)(89) := currentData(89); xorBitMap(18)(88) := currentData(88); xorBitMap(18)(86) := currentData(86); xorBitMap(18)(85) := currentData(85); xorBitMap(18)(84) := currentData(84); xorBitMap(18)(80) := currentData(80); xorBitMap(18)(79) := currentData(79); xorBitMap(18)(77) := currentData(77); xorBitMap(18)(70) := currentData(70); xorBitMap(18)(68) := currentData(68); xorBitMap(18)(59) := currentData(59); xorBitMap(18)(58) := currentData(58); xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(164) := previousCrc(4); xorBitMap(18)(166) := previousCrc(6); xorBitMap(18)(173) := previousCrc(13); xorBitMap(18)(175) := previousCrc(15); xorBitMap(18)(176) := previousCrc(16); xorBitMap(18)(180) := previousCrc(20); xorBitMap(18)(181) := previousCrc(21); xorBitMap(18)(182) := previousCrc(22); xorBitMap(18)(184) := previousCrc(24); xorBitMap(18)(185) := previousCrc(25); xorBitMap(18)(187) := previousCrc(27); xorBitMap(18)(188) := previousCrc(28); xorBitMap(18)(189) := previousCrc(29); 
      xorBitMap(19)(94) := currentData(94); xorBitMap(19)(93) := currentData(93); xorBitMap(19)(92) := currentData(92); xorBitMap(19)(90) := currentData(90); xorBitMap(19)(89) := currentData(89); xorBitMap(19)(87) := currentData(87); xorBitMap(19)(86) := currentData(86); xorBitMap(19)(85) := currentData(85); xorBitMap(19)(81) := currentData(81); xorBitMap(19)(80) := currentData(80); xorBitMap(19)(78) := currentData(78); xorBitMap(19)(71) := currentData(71); xorBitMap(19)(69) := currentData(69); xorBitMap(19)(60) := currentData(60); xorBitMap(19)(59) := currentData(59); xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(165) := previousCrc(5); xorBitMap(19)(167) := previousCrc(7); xorBitMap(19)(174) := previousCrc(14); xorBitMap(19)(176) := previousCrc(16); xorBitMap(19)(177) := previousCrc(17); xorBitMap(19)(181) := previousCrc(21); xorBitMap(19)(182) := previousCrc(22); xorBitMap(19)(183) := previousCrc(23); xorBitMap(19)(185) := previousCrc(25); xorBitMap(19)(186) := previousCrc(26); xorBitMap(19)(188) := previousCrc(28); xorBitMap(19)(189) := previousCrc(29); xorBitMap(19)(190) := previousCrc(30); 
      xorBitMap(20)(95) := currentData(95); xorBitMap(20)(94) := currentData(94); xorBitMap(20)(93) := currentData(93); xorBitMap(20)(91) := currentData(91); xorBitMap(20)(90) := currentData(90); xorBitMap(20)(88) := currentData(88); xorBitMap(20)(87) := currentData(87); xorBitMap(20)(86) := currentData(86); xorBitMap(20)(82) := currentData(82); xorBitMap(20)(81) := currentData(81); xorBitMap(20)(79) := currentData(79); xorBitMap(20)(72) := currentData(72); xorBitMap(20)(70) := currentData(70); xorBitMap(20)(61) := currentData(61); xorBitMap(20)(60) := currentData(60); xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(166) := previousCrc(6); xorBitMap(20)(168) := previousCrc(8); xorBitMap(20)(175) := previousCrc(15); xorBitMap(20)(177) := previousCrc(17); xorBitMap(20)(178) := previousCrc(18); xorBitMap(20)(182) := previousCrc(22); xorBitMap(20)(183) := previousCrc(23); xorBitMap(20)(184) := previousCrc(24); xorBitMap(20)(186) := previousCrc(26); xorBitMap(20)(187) := previousCrc(27); xorBitMap(20)(189) := previousCrc(29); xorBitMap(20)(190) := previousCrc(30); xorBitMap(20)(191) := previousCrc(31); 
      xorBitMap(21)(95) := currentData(95); xorBitMap(21)(94) := currentData(94); xorBitMap(21)(92) := currentData(92); xorBitMap(21)(91) := currentData(91); xorBitMap(21)(89) := currentData(89); xorBitMap(21)(88) := currentData(88); xorBitMap(21)(87) := currentData(87); xorBitMap(21)(83) := currentData(83); xorBitMap(21)(82) := currentData(82); xorBitMap(21)(80) := currentData(80); xorBitMap(21)(73) := currentData(73); xorBitMap(21)(71) := currentData(71); xorBitMap(21)(62) := currentData(62); xorBitMap(21)(61) := currentData(61); xorBitMap(21)(56) := currentData(56); xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(167) := previousCrc(7); xorBitMap(21)(169) := previousCrc(9); xorBitMap(21)(176) := previousCrc(16); xorBitMap(21)(178) := previousCrc(18); xorBitMap(21)(179) := previousCrc(19); xorBitMap(21)(183) := previousCrc(23); xorBitMap(21)(184) := previousCrc(24); xorBitMap(21)(185) := previousCrc(25); xorBitMap(21)(187) := previousCrc(27); xorBitMap(21)(188) := previousCrc(28); xorBitMap(21)(190) := previousCrc(30); xorBitMap(21)(191) := previousCrc(31); 
      xorBitMap(22)(94) := currentData(94); xorBitMap(22)(93) := currentData(93); xorBitMap(22)(92) := currentData(92); xorBitMap(22)(90) := currentData(90); xorBitMap(22)(89) := currentData(89); xorBitMap(22)(88) := currentData(88); xorBitMap(22)(87) := currentData(87); xorBitMap(22)(85) := currentData(85); xorBitMap(22)(82) := currentData(82); xorBitMap(22)(79) := currentData(79); xorBitMap(22)(74) := currentData(74); xorBitMap(22)(73) := currentData(73); xorBitMap(22)(68) := currentData(68); xorBitMap(22)(67) := currentData(67); xorBitMap(22)(66) := currentData(66); xorBitMap(22)(65) := currentData(65); xorBitMap(22)(62) := currentData(62); xorBitMap(22)(61) := currentData(61); xorBitMap(22)(60) := currentData(60); xorBitMap(22)(58) := currentData(58); xorBitMap(22)(57) := currentData(57); xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(161) := previousCrc(1); xorBitMap(22)(162) := previousCrc(2); xorBitMap(22)(163) := previousCrc(3); xorBitMap(22)(164) := previousCrc(4); xorBitMap(22)(169) := previousCrc(9); xorBitMap(22)(170) := previousCrc(10); xorBitMap(22)(175) := previousCrc(15); xorBitMap(22)(178) := previousCrc(18); xorBitMap(22)(181) := previousCrc(21); xorBitMap(22)(183) := previousCrc(23); xorBitMap(22)(184) := previousCrc(24); xorBitMap(22)(185) := previousCrc(25); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(188) := previousCrc(28); xorBitMap(22)(189) := previousCrc(29); xorBitMap(22)(190) := previousCrc(30); 
      xorBitMap(23)(93) := currentData(93); xorBitMap(23)(91) := currentData(91); xorBitMap(23)(90) := currentData(90); xorBitMap(23)(89) := currentData(89); xorBitMap(23)(88) := currentData(88); xorBitMap(23)(87) := currentData(87); xorBitMap(23)(86) := currentData(86); xorBitMap(23)(85) := currentData(85); xorBitMap(23)(84) := currentData(84); xorBitMap(23)(82) := currentData(82); xorBitMap(23)(81) := currentData(81); xorBitMap(23)(80) := currentData(80); xorBitMap(23)(79) := currentData(79); xorBitMap(23)(75) := currentData(75); xorBitMap(23)(74) := currentData(74); xorBitMap(23)(73) := currentData(73); xorBitMap(23)(72) := currentData(72); xorBitMap(23)(69) := currentData(69); xorBitMap(23)(65) := currentData(65); xorBitMap(23)(62) := currentData(62); xorBitMap(23)(60) := currentData(60); xorBitMap(23)(59) := currentData(59); xorBitMap(23)(56) := currentData(56); xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(161) := previousCrc(1); xorBitMap(23)(165) := previousCrc(5); xorBitMap(23)(168) := previousCrc(8); xorBitMap(23)(169) := previousCrc(9); xorBitMap(23)(170) := previousCrc(10); xorBitMap(23)(171) := previousCrc(11); xorBitMap(23)(175) := previousCrc(15); xorBitMap(23)(176) := previousCrc(16); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(178) := previousCrc(18); xorBitMap(23)(180) := previousCrc(20); xorBitMap(23)(181) := previousCrc(21); xorBitMap(23)(182) := previousCrc(22); xorBitMap(23)(183) := previousCrc(23); xorBitMap(23)(184) := previousCrc(24); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(186) := previousCrc(26); xorBitMap(23)(187) := previousCrc(27); xorBitMap(23)(189) := previousCrc(29); 
      xorBitMap(24)(94) := currentData(94); xorBitMap(24)(92) := currentData(92); xorBitMap(24)(91) := currentData(91); xorBitMap(24)(90) := currentData(90); xorBitMap(24)(89) := currentData(89); xorBitMap(24)(88) := currentData(88); xorBitMap(24)(87) := currentData(87); xorBitMap(24)(86) := currentData(86); xorBitMap(24)(85) := currentData(85); xorBitMap(24)(83) := currentData(83); xorBitMap(24)(82) := currentData(82); xorBitMap(24)(81) := currentData(81); xorBitMap(24)(80) := currentData(80); xorBitMap(24)(76) := currentData(76); xorBitMap(24)(75) := currentData(75); xorBitMap(24)(74) := currentData(74); xorBitMap(24)(73) := currentData(73); xorBitMap(24)(70) := currentData(70); xorBitMap(24)(66) := currentData(66); xorBitMap(24)(63) := currentData(63); xorBitMap(24)(61) := currentData(61); xorBitMap(24)(60) := currentData(60); xorBitMap(24)(57) := currentData(57); xorBitMap(24)(56) := currentData(56); xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(162) := previousCrc(2); xorBitMap(24)(166) := previousCrc(6); xorBitMap(24)(169) := previousCrc(9); xorBitMap(24)(170) := previousCrc(10); xorBitMap(24)(171) := previousCrc(11); xorBitMap(24)(172) := previousCrc(12); xorBitMap(24)(176) := previousCrc(16); xorBitMap(24)(177) := previousCrc(17); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(179) := previousCrc(19); xorBitMap(24)(181) := previousCrc(21); xorBitMap(24)(182) := previousCrc(22); xorBitMap(24)(183) := previousCrc(23); xorBitMap(24)(184) := previousCrc(24); xorBitMap(24)(185) := previousCrc(25); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(187) := previousCrc(27); xorBitMap(24)(188) := previousCrc(28); xorBitMap(24)(190) := previousCrc(30); 
      xorBitMap(25)(95) := currentData(95); xorBitMap(25)(93) := currentData(93); xorBitMap(25)(92) := currentData(92); xorBitMap(25)(91) := currentData(91); xorBitMap(25)(90) := currentData(90); xorBitMap(25)(89) := currentData(89); xorBitMap(25)(88) := currentData(88); xorBitMap(25)(87) := currentData(87); xorBitMap(25)(86) := currentData(86); xorBitMap(25)(84) := currentData(84); xorBitMap(25)(83) := currentData(83); xorBitMap(25)(82) := currentData(82); xorBitMap(25)(81) := currentData(81); xorBitMap(25)(77) := currentData(77); xorBitMap(25)(76) := currentData(76); xorBitMap(25)(75) := currentData(75); xorBitMap(25)(74) := currentData(74); xorBitMap(25)(71) := currentData(71); xorBitMap(25)(67) := currentData(67); xorBitMap(25)(64) := currentData(64); xorBitMap(25)(62) := currentData(62); xorBitMap(25)(61) := currentData(61); xorBitMap(25)(58) := currentData(58); xorBitMap(25)(57) := currentData(57); xorBitMap(25)(56) := currentData(56); xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(160) := previousCrc(0); xorBitMap(25)(163) := previousCrc(3); xorBitMap(25)(167) := previousCrc(7); xorBitMap(25)(170) := previousCrc(10); xorBitMap(25)(171) := previousCrc(11); xorBitMap(25)(172) := previousCrc(12); xorBitMap(25)(173) := previousCrc(13); xorBitMap(25)(177) := previousCrc(17); xorBitMap(25)(178) := previousCrc(18); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(180) := previousCrc(20); xorBitMap(25)(182) := previousCrc(22); xorBitMap(25)(183) := previousCrc(23); xorBitMap(25)(184) := previousCrc(24); xorBitMap(25)(185) := previousCrc(25); xorBitMap(25)(186) := previousCrc(26); xorBitMap(25)(187) := previousCrc(27); xorBitMap(25)(188) := previousCrc(28); xorBitMap(25)(189) := previousCrc(29); xorBitMap(25)(191) := previousCrc(31); 
      xorBitMap(26)(95) := currentData(95); xorBitMap(26)(93) := currentData(93); xorBitMap(26)(92) := currentData(92); xorBitMap(26)(91) := currentData(91); xorBitMap(26)(90) := currentData(90); xorBitMap(26)(89) := currentData(89); xorBitMap(26)(88) := currentData(88); xorBitMap(26)(81) := currentData(81); xorBitMap(26)(79) := currentData(79); xorBitMap(26)(78) := currentData(78); xorBitMap(26)(77) := currentData(77); xorBitMap(26)(76) := currentData(76); xorBitMap(26)(75) := currentData(75); xorBitMap(26)(73) := currentData(73); xorBitMap(26)(67) := currentData(67); xorBitMap(26)(66) := currentData(66); xorBitMap(26)(62) := currentData(62); xorBitMap(26)(61) := currentData(61); xorBitMap(26)(60) := currentData(60); xorBitMap(26)(59) := currentData(59); xorBitMap(26)(57) := currentData(57); xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(162) := previousCrc(2); xorBitMap(26)(163) := previousCrc(3); xorBitMap(26)(169) := previousCrc(9); xorBitMap(26)(171) := previousCrc(11); xorBitMap(26)(172) := previousCrc(12); xorBitMap(26)(173) := previousCrc(13); xorBitMap(26)(174) := previousCrc(14); xorBitMap(26)(175) := previousCrc(15); xorBitMap(26)(177) := previousCrc(17); xorBitMap(26)(184) := previousCrc(24); xorBitMap(26)(185) := previousCrc(25); xorBitMap(26)(186) := previousCrc(26); xorBitMap(26)(187) := previousCrc(27); xorBitMap(26)(188) := previousCrc(28); xorBitMap(26)(189) := previousCrc(29); xorBitMap(26)(191) := previousCrc(31); 
      xorBitMap(27)(94) := currentData(94); xorBitMap(27)(93) := currentData(93); xorBitMap(27)(92) := currentData(92); xorBitMap(27)(91) := currentData(91); xorBitMap(27)(90) := currentData(90); xorBitMap(27)(89) := currentData(89); xorBitMap(27)(82) := currentData(82); xorBitMap(27)(80) := currentData(80); xorBitMap(27)(79) := currentData(79); xorBitMap(27)(78) := currentData(78); xorBitMap(27)(77) := currentData(77); xorBitMap(27)(76) := currentData(76); xorBitMap(27)(74) := currentData(74); xorBitMap(27)(68) := currentData(68); xorBitMap(27)(67) := currentData(67); xorBitMap(27)(63) := currentData(63); xorBitMap(27)(62) := currentData(62); xorBitMap(27)(61) := currentData(61); xorBitMap(27)(60) := currentData(60); xorBitMap(27)(58) := currentData(58); xorBitMap(27)(56) := currentData(56); xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(163) := previousCrc(3); xorBitMap(27)(164) := previousCrc(4); xorBitMap(27)(170) := previousCrc(10); xorBitMap(27)(172) := previousCrc(12); xorBitMap(27)(173) := previousCrc(13); xorBitMap(27)(174) := previousCrc(14); xorBitMap(27)(175) := previousCrc(15); xorBitMap(27)(176) := previousCrc(16); xorBitMap(27)(178) := previousCrc(18); xorBitMap(27)(185) := previousCrc(25); xorBitMap(27)(186) := previousCrc(26); xorBitMap(27)(187) := previousCrc(27); xorBitMap(27)(188) := previousCrc(28); xorBitMap(27)(189) := previousCrc(29); xorBitMap(27)(190) := previousCrc(30); 
      xorBitMap(28)(95) := currentData(95); xorBitMap(28)(94) := currentData(94); xorBitMap(28)(93) := currentData(93); xorBitMap(28)(92) := currentData(92); xorBitMap(28)(91) := currentData(91); xorBitMap(28)(90) := currentData(90); xorBitMap(28)(83) := currentData(83); xorBitMap(28)(81) := currentData(81); xorBitMap(28)(80) := currentData(80); xorBitMap(28)(79) := currentData(79); xorBitMap(28)(78) := currentData(78); xorBitMap(28)(77) := currentData(77); xorBitMap(28)(75) := currentData(75); xorBitMap(28)(69) := currentData(69); xorBitMap(28)(68) := currentData(68); xorBitMap(28)(64) := currentData(64); xorBitMap(28)(63) := currentData(63); xorBitMap(28)(62) := currentData(62); xorBitMap(28)(61) := currentData(61); xorBitMap(28)(59) := currentData(59); xorBitMap(28)(57) := currentData(57); xorBitMap(28)(56) := currentData(56); xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(160) := previousCrc(0); xorBitMap(28)(164) := previousCrc(4); xorBitMap(28)(165) := previousCrc(5); xorBitMap(28)(171) := previousCrc(11); xorBitMap(28)(173) := previousCrc(13); xorBitMap(28)(174) := previousCrc(14); xorBitMap(28)(175) := previousCrc(15); xorBitMap(28)(176) := previousCrc(16); xorBitMap(28)(177) := previousCrc(17); xorBitMap(28)(179) := previousCrc(19); xorBitMap(28)(186) := previousCrc(26); xorBitMap(28)(187) := previousCrc(27); xorBitMap(28)(188) := previousCrc(28); xorBitMap(28)(189) := previousCrc(29); xorBitMap(28)(190) := previousCrc(30); xorBitMap(28)(191) := previousCrc(31); 
      xorBitMap(29)(95) := currentData(95); xorBitMap(29)(94) := currentData(94); xorBitMap(29)(93) := currentData(93); xorBitMap(29)(92) := currentData(92); xorBitMap(29)(91) := currentData(91); xorBitMap(29)(84) := currentData(84); xorBitMap(29)(82) := currentData(82); xorBitMap(29)(81) := currentData(81); xorBitMap(29)(80) := currentData(80); xorBitMap(29)(79) := currentData(79); xorBitMap(29)(78) := currentData(78); xorBitMap(29)(76) := currentData(76); xorBitMap(29)(70) := currentData(70); xorBitMap(29)(69) := currentData(69); xorBitMap(29)(65) := currentData(65); xorBitMap(29)(64) := currentData(64); xorBitMap(29)(63) := currentData(63); xorBitMap(29)(62) := currentData(62); xorBitMap(29)(60) := currentData(60); xorBitMap(29)(58) := currentData(58); xorBitMap(29)(57) := currentData(57); xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(160) := previousCrc(0); xorBitMap(29)(161) := previousCrc(1); xorBitMap(29)(165) := previousCrc(5); xorBitMap(29)(166) := previousCrc(6); xorBitMap(29)(172) := previousCrc(12); xorBitMap(29)(174) := previousCrc(14); xorBitMap(29)(175) := previousCrc(15); xorBitMap(29)(176) := previousCrc(16); xorBitMap(29)(177) := previousCrc(17); xorBitMap(29)(178) := previousCrc(18); xorBitMap(29)(180) := previousCrc(20); xorBitMap(29)(187) := previousCrc(27); xorBitMap(29)(188) := previousCrc(28); xorBitMap(29)(189) := previousCrc(29); xorBitMap(29)(190) := previousCrc(30); xorBitMap(29)(191) := previousCrc(31); 
      xorBitMap(30)(95) := currentData(95); xorBitMap(30)(94) := currentData(94); xorBitMap(30)(93) := currentData(93); xorBitMap(30)(92) := currentData(92); xorBitMap(30)(85) := currentData(85); xorBitMap(30)(83) := currentData(83); xorBitMap(30)(82) := currentData(82); xorBitMap(30)(81) := currentData(81); xorBitMap(30)(80) := currentData(80); xorBitMap(30)(79) := currentData(79); xorBitMap(30)(77) := currentData(77); xorBitMap(30)(71) := currentData(71); xorBitMap(30)(70) := currentData(70); xorBitMap(30)(66) := currentData(66); xorBitMap(30)(65) := currentData(65); xorBitMap(30)(64) := currentData(64); xorBitMap(30)(63) := currentData(63); xorBitMap(30)(61) := currentData(61); xorBitMap(30)(59) := currentData(59); xorBitMap(30)(58) := currentData(58); xorBitMap(30)(56) := currentData(56); xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(160) := previousCrc(0); xorBitMap(30)(161) := previousCrc(1); xorBitMap(30)(162) := previousCrc(2); xorBitMap(30)(166) := previousCrc(6); xorBitMap(30)(167) := previousCrc(7); xorBitMap(30)(173) := previousCrc(13); xorBitMap(30)(175) := previousCrc(15); xorBitMap(30)(176) := previousCrc(16); xorBitMap(30)(177) := previousCrc(17); xorBitMap(30)(178) := previousCrc(18); xorBitMap(30)(179) := previousCrc(19); xorBitMap(30)(181) := previousCrc(21); xorBitMap(30)(188) := previousCrc(28); xorBitMap(30)(189) := previousCrc(29); xorBitMap(30)(190) := previousCrc(30); xorBitMap(30)(191) := previousCrc(31); 
      xorBitMap(31)(95) := currentData(95); xorBitMap(31)(94) := currentData(94); xorBitMap(31)(93) := currentData(93); xorBitMap(31)(86) := currentData(86); xorBitMap(31)(84) := currentData(84); xorBitMap(31)(83) := currentData(83); xorBitMap(31)(82) := currentData(82); xorBitMap(31)(81) := currentData(81); xorBitMap(31)(80) := currentData(80); xorBitMap(31)(78) := currentData(78); xorBitMap(31)(72) := currentData(72); xorBitMap(31)(71) := currentData(71); xorBitMap(31)(67) := currentData(67); xorBitMap(31)(66) := currentData(66); xorBitMap(31)(65) := currentData(65); xorBitMap(31)(64) := currentData(64); xorBitMap(31)(62) := currentData(62); xorBitMap(31)(60) := currentData(60); xorBitMap(31)(59) := currentData(59); xorBitMap(31)(57) := currentData(57); xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(160) := previousCrc(0); xorBitMap(31)(161) := previousCrc(1); xorBitMap(31)(162) := previousCrc(2); xorBitMap(31)(163) := previousCrc(3); xorBitMap(31)(167) := previousCrc(7); xorBitMap(31)(168) := previousCrc(8); xorBitMap(31)(174) := previousCrc(14); xorBitMap(31)(176) := previousCrc(16); xorBitMap(31)(177) := previousCrc(17); xorBitMap(31)(178) := previousCrc(18); xorBitMap(31)(179) := previousCrc(19); xorBitMap(31)(180) := previousCrc(20); xorBitMap(31)(182) := previousCrc(22); xorBitMap(31)(189) := previousCrc(29); xorBitMap(31)(190) := previousCrc(30); xorBitMap(31)(191) := previousCrc(31); 
   end procedure;

   procedure xorBitMap13Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(103 downto 0)) is 
   begin
      xorBitMap(0)(103) := currentData(103); xorBitMap(0)(101) := currentData(101); xorBitMap(0)(99) := currentData(99); xorBitMap(0)(98) := currentData(98); xorBitMap(0)(97) := currentData(97); xorBitMap(0)(96) := currentData(96); xorBitMap(0)(95) := currentData(95); xorBitMap(0)(94) := currentData(94); xorBitMap(0)(87) := currentData(87); xorBitMap(0)(85) := currentData(85); xorBitMap(0)(84) := currentData(84); xorBitMap(0)(83) := currentData(83); xorBitMap(0)(82) := currentData(82); xorBitMap(0)(81) := currentData(81); xorBitMap(0)(79) := currentData(79); xorBitMap(0)(73) := currentData(73); xorBitMap(0)(72) := currentData(72); xorBitMap(0)(68) := currentData(68); xorBitMap(0)(67) := currentData(67); xorBitMap(0)(66) := currentData(66); xorBitMap(0)(65) := currentData(65); xorBitMap(0)(63) := currentData(63); xorBitMap(0)(61) := currentData(61); xorBitMap(0)(60) := currentData(60); xorBitMap(0)(58) := currentData(58); xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(160) := previousCrc(0); xorBitMap(0)(161) := previousCrc(1); xorBitMap(0)(167) := previousCrc(7); xorBitMap(0)(169) := previousCrc(9); xorBitMap(0)(170) := previousCrc(10); xorBitMap(0)(171) := previousCrc(11); xorBitMap(0)(172) := previousCrc(12); xorBitMap(0)(173) := previousCrc(13); xorBitMap(0)(175) := previousCrc(15); xorBitMap(0)(182) := previousCrc(22); xorBitMap(0)(183) := previousCrc(23); xorBitMap(0)(184) := previousCrc(24); xorBitMap(0)(185) := previousCrc(25); xorBitMap(0)(186) := previousCrc(26); xorBitMap(0)(187) := previousCrc(27); xorBitMap(0)(189) := previousCrc(29); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(103) := currentData(103); xorBitMap(1)(102) := currentData(102); xorBitMap(1)(101) := currentData(101); xorBitMap(1)(100) := currentData(100); xorBitMap(1)(94) := currentData(94); xorBitMap(1)(88) := currentData(88); xorBitMap(1)(87) := currentData(87); xorBitMap(1)(86) := currentData(86); xorBitMap(1)(81) := currentData(81); xorBitMap(1)(80) := currentData(80); xorBitMap(1)(79) := currentData(79); xorBitMap(1)(74) := currentData(74); xorBitMap(1)(72) := currentData(72); xorBitMap(1)(69) := currentData(69); xorBitMap(1)(65) := currentData(65); xorBitMap(1)(64) := currentData(64); xorBitMap(1)(63) := currentData(63); xorBitMap(1)(62) := currentData(62); xorBitMap(1)(60) := currentData(60); xorBitMap(1)(59) := currentData(59); xorBitMap(1)(58) := currentData(58); xorBitMap(1)(56) := currentData(56); xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(160) := previousCrc(0); xorBitMap(1)(162) := previousCrc(2); xorBitMap(1)(167) := previousCrc(7); xorBitMap(1)(168) := previousCrc(8); xorBitMap(1)(169) := previousCrc(9); xorBitMap(1)(174) := previousCrc(14); xorBitMap(1)(175) := previousCrc(15); xorBitMap(1)(176) := previousCrc(16); xorBitMap(1)(182) := previousCrc(22); xorBitMap(1)(188) := previousCrc(28); xorBitMap(1)(189) := previousCrc(29); xorBitMap(1)(190) := previousCrc(30); xorBitMap(1)(191) := previousCrc(31); 
      xorBitMap(2)(102) := currentData(102); xorBitMap(2)(99) := currentData(99); xorBitMap(2)(98) := currentData(98); xorBitMap(2)(97) := currentData(97); xorBitMap(2)(96) := currentData(96); xorBitMap(2)(94) := currentData(94); xorBitMap(2)(89) := currentData(89); xorBitMap(2)(88) := currentData(88); xorBitMap(2)(85) := currentData(85); xorBitMap(2)(84) := currentData(84); xorBitMap(2)(83) := currentData(83); xorBitMap(2)(80) := currentData(80); xorBitMap(2)(79) := currentData(79); xorBitMap(2)(75) := currentData(75); xorBitMap(2)(72) := currentData(72); xorBitMap(2)(70) := currentData(70); xorBitMap(2)(68) := currentData(68); xorBitMap(2)(67) := currentData(67); xorBitMap(2)(64) := currentData(64); xorBitMap(2)(59) := currentData(59); xorBitMap(2)(58) := currentData(58); xorBitMap(2)(57) := currentData(57); xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(160) := previousCrc(0); xorBitMap(2)(163) := previousCrc(3); xorBitMap(2)(167) := previousCrc(7); xorBitMap(2)(168) := previousCrc(8); xorBitMap(2)(171) := previousCrc(11); xorBitMap(2)(172) := previousCrc(12); xorBitMap(2)(173) := previousCrc(13); xorBitMap(2)(176) := previousCrc(16); xorBitMap(2)(177) := previousCrc(17); xorBitMap(2)(182) := previousCrc(22); xorBitMap(2)(184) := previousCrc(24); xorBitMap(2)(185) := previousCrc(25); xorBitMap(2)(186) := previousCrc(26); xorBitMap(2)(187) := previousCrc(27); xorBitMap(2)(190) := previousCrc(30); 
      xorBitMap(3)(103) := currentData(103); xorBitMap(3)(100) := currentData(100); xorBitMap(3)(99) := currentData(99); xorBitMap(3)(98) := currentData(98); xorBitMap(3)(97) := currentData(97); xorBitMap(3)(95) := currentData(95); xorBitMap(3)(90) := currentData(90); xorBitMap(3)(89) := currentData(89); xorBitMap(3)(86) := currentData(86); xorBitMap(3)(85) := currentData(85); xorBitMap(3)(84) := currentData(84); xorBitMap(3)(81) := currentData(81); xorBitMap(3)(80) := currentData(80); xorBitMap(3)(76) := currentData(76); xorBitMap(3)(73) := currentData(73); xorBitMap(3)(71) := currentData(71); xorBitMap(3)(69) := currentData(69); xorBitMap(3)(68) := currentData(68); xorBitMap(3)(65) := currentData(65); xorBitMap(3)(60) := currentData(60); xorBitMap(3)(59) := currentData(59); xorBitMap(3)(58) := currentData(58); xorBitMap(3)(56) := currentData(56); xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(161) := previousCrc(1); xorBitMap(3)(164) := previousCrc(4); xorBitMap(3)(168) := previousCrc(8); xorBitMap(3)(169) := previousCrc(9); xorBitMap(3)(172) := previousCrc(12); xorBitMap(3)(173) := previousCrc(13); xorBitMap(3)(174) := previousCrc(14); xorBitMap(3)(177) := previousCrc(17); xorBitMap(3)(178) := previousCrc(18); xorBitMap(3)(183) := previousCrc(23); xorBitMap(3)(185) := previousCrc(25); xorBitMap(3)(186) := previousCrc(26); xorBitMap(3)(187) := previousCrc(27); xorBitMap(3)(188) := previousCrc(28); xorBitMap(3)(191) := previousCrc(31); 
      xorBitMap(4)(103) := currentData(103); xorBitMap(4)(100) := currentData(100); xorBitMap(4)(97) := currentData(97); xorBitMap(4)(95) := currentData(95); xorBitMap(4)(94) := currentData(94); xorBitMap(4)(91) := currentData(91); xorBitMap(4)(90) := currentData(90); xorBitMap(4)(86) := currentData(86); xorBitMap(4)(84) := currentData(84); xorBitMap(4)(83) := currentData(83); xorBitMap(4)(79) := currentData(79); xorBitMap(4)(77) := currentData(77); xorBitMap(4)(74) := currentData(74); xorBitMap(4)(73) := currentData(73); xorBitMap(4)(70) := currentData(70); xorBitMap(4)(69) := currentData(69); xorBitMap(4)(68) := currentData(68); xorBitMap(4)(67) := currentData(67); xorBitMap(4)(65) := currentData(65); xorBitMap(4)(63) := currentData(63); xorBitMap(4)(59) := currentData(59); xorBitMap(4)(58) := currentData(58); xorBitMap(4)(57) := currentData(57); xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(161) := previousCrc(1); xorBitMap(4)(162) := previousCrc(2); xorBitMap(4)(165) := previousCrc(5); xorBitMap(4)(167) := previousCrc(7); xorBitMap(4)(171) := previousCrc(11); xorBitMap(4)(172) := previousCrc(12); xorBitMap(4)(174) := previousCrc(14); xorBitMap(4)(178) := previousCrc(18); xorBitMap(4)(179) := previousCrc(19); xorBitMap(4)(182) := previousCrc(22); xorBitMap(4)(183) := previousCrc(23); xorBitMap(4)(185) := previousCrc(25); xorBitMap(4)(188) := previousCrc(28); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(103) := currentData(103); xorBitMap(5)(99) := currentData(99); xorBitMap(5)(97) := currentData(97); xorBitMap(5)(94) := currentData(94); xorBitMap(5)(92) := currentData(92); xorBitMap(5)(91) := currentData(91); xorBitMap(5)(83) := currentData(83); xorBitMap(5)(82) := currentData(82); xorBitMap(5)(81) := currentData(81); xorBitMap(5)(80) := currentData(80); xorBitMap(5)(79) := currentData(79); xorBitMap(5)(78) := currentData(78); xorBitMap(5)(75) := currentData(75); xorBitMap(5)(74) := currentData(74); xorBitMap(5)(73) := currentData(73); xorBitMap(5)(72) := currentData(72); xorBitMap(5)(71) := currentData(71); xorBitMap(5)(70) := currentData(70); xorBitMap(5)(69) := currentData(69); xorBitMap(5)(67) := currentData(67); xorBitMap(5)(65) := currentData(65); xorBitMap(5)(64) := currentData(64); xorBitMap(5)(63) := currentData(63); xorBitMap(5)(61) := currentData(61); xorBitMap(5)(59) := currentData(59); xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(160) := previousCrc(0); xorBitMap(5)(161) := previousCrc(1); xorBitMap(5)(162) := previousCrc(2); xorBitMap(5)(163) := previousCrc(3); xorBitMap(5)(166) := previousCrc(6); xorBitMap(5)(167) := previousCrc(7); xorBitMap(5)(168) := previousCrc(8); xorBitMap(5)(169) := previousCrc(9); xorBitMap(5)(170) := previousCrc(10); xorBitMap(5)(171) := previousCrc(11); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(180) := previousCrc(20); xorBitMap(5)(182) := previousCrc(22); xorBitMap(5)(185) := previousCrc(25); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(191) := previousCrc(31); 
      xorBitMap(6)(100) := currentData(100); xorBitMap(6)(98) := currentData(98); xorBitMap(6)(95) := currentData(95); xorBitMap(6)(93) := currentData(93); xorBitMap(6)(92) := currentData(92); xorBitMap(6)(84) := currentData(84); xorBitMap(6)(83) := currentData(83); xorBitMap(6)(82) := currentData(82); xorBitMap(6)(81) := currentData(81); xorBitMap(6)(80) := currentData(80); xorBitMap(6)(79) := currentData(79); xorBitMap(6)(76) := currentData(76); xorBitMap(6)(75) := currentData(75); xorBitMap(6)(74) := currentData(74); xorBitMap(6)(73) := currentData(73); xorBitMap(6)(72) := currentData(72); xorBitMap(6)(71) := currentData(71); xorBitMap(6)(70) := currentData(70); xorBitMap(6)(68) := currentData(68); xorBitMap(6)(66) := currentData(66); xorBitMap(6)(65) := currentData(65); xorBitMap(6)(64) := currentData(64); xorBitMap(6)(62) := currentData(62); xorBitMap(6)(60) := currentData(60); xorBitMap(6)(56) := currentData(56); xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(160) := previousCrc(0); xorBitMap(6)(161) := previousCrc(1); xorBitMap(6)(162) := previousCrc(2); xorBitMap(6)(163) := previousCrc(3); xorBitMap(6)(164) := previousCrc(4); xorBitMap(6)(167) := previousCrc(7); xorBitMap(6)(168) := previousCrc(8); xorBitMap(6)(169) := previousCrc(9); xorBitMap(6)(170) := previousCrc(10); xorBitMap(6)(171) := previousCrc(11); xorBitMap(6)(172) := previousCrc(12); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(181) := previousCrc(21); xorBitMap(6)(183) := previousCrc(23); xorBitMap(6)(186) := previousCrc(26); xorBitMap(6)(188) := previousCrc(28); 
      xorBitMap(7)(103) := currentData(103); xorBitMap(7)(98) := currentData(98); xorBitMap(7)(97) := currentData(97); xorBitMap(7)(95) := currentData(95); xorBitMap(7)(93) := currentData(93); xorBitMap(7)(87) := currentData(87); xorBitMap(7)(80) := currentData(80); xorBitMap(7)(79) := currentData(79); xorBitMap(7)(77) := currentData(77); xorBitMap(7)(76) := currentData(76); xorBitMap(7)(75) := currentData(75); xorBitMap(7)(74) := currentData(74); xorBitMap(7)(71) := currentData(71); xorBitMap(7)(69) := currentData(69); xorBitMap(7)(68) := currentData(68); xorBitMap(7)(60) := currentData(60); xorBitMap(7)(58) := currentData(58); xorBitMap(7)(57) := currentData(57); xorBitMap(7)(56) := currentData(56); xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(162) := previousCrc(2); xorBitMap(7)(163) := previousCrc(3); xorBitMap(7)(164) := previousCrc(4); xorBitMap(7)(165) := previousCrc(5); xorBitMap(7)(167) := previousCrc(7); xorBitMap(7)(168) := previousCrc(8); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(181) := previousCrc(21); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(185) := previousCrc(25); xorBitMap(7)(186) := previousCrc(26); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(103) := currentData(103); xorBitMap(8)(101) := currentData(101); xorBitMap(8)(97) := currentData(97); xorBitMap(8)(95) := currentData(95); xorBitMap(8)(88) := currentData(88); xorBitMap(8)(87) := currentData(87); xorBitMap(8)(85) := currentData(85); xorBitMap(8)(84) := currentData(84); xorBitMap(8)(83) := currentData(83); xorBitMap(8)(82) := currentData(82); xorBitMap(8)(80) := currentData(80); xorBitMap(8)(79) := currentData(79); xorBitMap(8)(78) := currentData(78); xorBitMap(8)(77) := currentData(77); xorBitMap(8)(76) := currentData(76); xorBitMap(8)(75) := currentData(75); xorBitMap(8)(73) := currentData(73); xorBitMap(8)(70) := currentData(70); xorBitMap(8)(69) := currentData(69); xorBitMap(8)(68) := currentData(68); xorBitMap(8)(67) := currentData(67); xorBitMap(8)(66) := currentData(66); xorBitMap(8)(65) := currentData(65); xorBitMap(8)(63) := currentData(63); xorBitMap(8)(60) := currentData(60); xorBitMap(8)(59) := currentData(59); xorBitMap(8)(57) := currentData(57); xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(161) := previousCrc(1); xorBitMap(8)(163) := previousCrc(3); xorBitMap(8)(164) := previousCrc(4); xorBitMap(8)(165) := previousCrc(5); xorBitMap(8)(166) := previousCrc(6); xorBitMap(8)(167) := previousCrc(7); xorBitMap(8)(168) := previousCrc(8); xorBitMap(8)(170) := previousCrc(10); xorBitMap(8)(171) := previousCrc(11); xorBitMap(8)(172) := previousCrc(12); xorBitMap(8)(173) := previousCrc(13); xorBitMap(8)(175) := previousCrc(15); xorBitMap(8)(176) := previousCrc(16); xorBitMap(8)(183) := previousCrc(23); xorBitMap(8)(185) := previousCrc(25); xorBitMap(8)(189) := previousCrc(29); xorBitMap(8)(191) := previousCrc(31); 
      xorBitMap(9)(102) := currentData(102); xorBitMap(9)(98) := currentData(98); xorBitMap(9)(96) := currentData(96); xorBitMap(9)(89) := currentData(89); xorBitMap(9)(88) := currentData(88); xorBitMap(9)(86) := currentData(86); xorBitMap(9)(85) := currentData(85); xorBitMap(9)(84) := currentData(84); xorBitMap(9)(83) := currentData(83); xorBitMap(9)(81) := currentData(81); xorBitMap(9)(80) := currentData(80); xorBitMap(9)(79) := currentData(79); xorBitMap(9)(78) := currentData(78); xorBitMap(9)(77) := currentData(77); xorBitMap(9)(76) := currentData(76); xorBitMap(9)(74) := currentData(74); xorBitMap(9)(71) := currentData(71); xorBitMap(9)(70) := currentData(70); xorBitMap(9)(69) := currentData(69); xorBitMap(9)(68) := currentData(68); xorBitMap(9)(67) := currentData(67); xorBitMap(9)(66) := currentData(66); xorBitMap(9)(64) := currentData(64); xorBitMap(9)(61) := currentData(61); xorBitMap(9)(60) := currentData(60); xorBitMap(9)(58) := currentData(58); xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(162) := previousCrc(2); xorBitMap(9)(164) := previousCrc(4); xorBitMap(9)(165) := previousCrc(5); xorBitMap(9)(166) := previousCrc(6); xorBitMap(9)(167) := previousCrc(7); xorBitMap(9)(168) := previousCrc(8); xorBitMap(9)(169) := previousCrc(9); xorBitMap(9)(171) := previousCrc(11); xorBitMap(9)(172) := previousCrc(12); xorBitMap(9)(173) := previousCrc(13); xorBitMap(9)(174) := previousCrc(14); xorBitMap(9)(176) := previousCrc(16); xorBitMap(9)(177) := previousCrc(17); xorBitMap(9)(184) := previousCrc(24); xorBitMap(9)(186) := previousCrc(26); xorBitMap(9)(190) := previousCrc(30); 
      xorBitMap(10)(101) := currentData(101); xorBitMap(10)(98) := currentData(98); xorBitMap(10)(96) := currentData(96); xorBitMap(10)(95) := currentData(95); xorBitMap(10)(94) := currentData(94); xorBitMap(10)(90) := currentData(90); xorBitMap(10)(89) := currentData(89); xorBitMap(10)(86) := currentData(86); xorBitMap(10)(83) := currentData(83); xorBitMap(10)(80) := currentData(80); xorBitMap(10)(78) := currentData(78); xorBitMap(10)(77) := currentData(77); xorBitMap(10)(75) := currentData(75); xorBitMap(10)(73) := currentData(73); xorBitMap(10)(71) := currentData(71); xorBitMap(10)(70) := currentData(70); xorBitMap(10)(69) := currentData(69); xorBitMap(10)(66) := currentData(66); xorBitMap(10)(63) := currentData(63); xorBitMap(10)(62) := currentData(62); xorBitMap(10)(60) := currentData(60); xorBitMap(10)(59) := currentData(59); xorBitMap(10)(58) := currentData(58); xorBitMap(10)(56) := currentData(56); xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(161) := previousCrc(1); xorBitMap(10)(163) := previousCrc(3); xorBitMap(10)(165) := previousCrc(5); xorBitMap(10)(166) := previousCrc(6); xorBitMap(10)(168) := previousCrc(8); xorBitMap(10)(171) := previousCrc(11); xorBitMap(10)(174) := previousCrc(14); xorBitMap(10)(177) := previousCrc(17); xorBitMap(10)(178) := previousCrc(18); xorBitMap(10)(182) := previousCrc(22); xorBitMap(10)(183) := previousCrc(23); xorBitMap(10)(184) := previousCrc(24); xorBitMap(10)(186) := previousCrc(26); xorBitMap(10)(189) := previousCrc(29); 
      xorBitMap(11)(103) := currentData(103); xorBitMap(11)(102) := currentData(102); xorBitMap(11)(101) := currentData(101); xorBitMap(11)(98) := currentData(98); xorBitMap(11)(94) := currentData(94); xorBitMap(11)(91) := currentData(91); xorBitMap(11)(90) := currentData(90); xorBitMap(11)(85) := currentData(85); xorBitMap(11)(83) := currentData(83); xorBitMap(11)(82) := currentData(82); xorBitMap(11)(78) := currentData(78); xorBitMap(11)(76) := currentData(76); xorBitMap(11)(74) := currentData(74); xorBitMap(11)(73) := currentData(73); xorBitMap(11)(71) := currentData(71); xorBitMap(11)(70) := currentData(70); xorBitMap(11)(68) := currentData(68); xorBitMap(11)(66) := currentData(66); xorBitMap(11)(65) := currentData(65); xorBitMap(11)(64) := currentData(64); xorBitMap(11)(59) := currentData(59); xorBitMap(11)(58) := currentData(58); xorBitMap(11)(57) := currentData(57); xorBitMap(11)(56) := currentData(56); xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(161) := previousCrc(1); xorBitMap(11)(162) := previousCrc(2); xorBitMap(11)(164) := previousCrc(4); xorBitMap(11)(166) := previousCrc(6); xorBitMap(11)(170) := previousCrc(10); xorBitMap(11)(171) := previousCrc(11); xorBitMap(11)(173) := previousCrc(13); xorBitMap(11)(178) := previousCrc(18); xorBitMap(11)(179) := previousCrc(19); xorBitMap(11)(182) := previousCrc(22); xorBitMap(11)(186) := previousCrc(26); xorBitMap(11)(189) := previousCrc(29); xorBitMap(11)(190) := previousCrc(30); xorBitMap(11)(191) := previousCrc(31); 
      xorBitMap(12)(102) := currentData(102); xorBitMap(12)(101) := currentData(101); xorBitMap(12)(98) := currentData(98); xorBitMap(12)(97) := currentData(97); xorBitMap(12)(96) := currentData(96); xorBitMap(12)(94) := currentData(94); xorBitMap(12)(92) := currentData(92); xorBitMap(12)(91) := currentData(91); xorBitMap(12)(87) := currentData(87); xorBitMap(12)(86) := currentData(86); xorBitMap(12)(85) := currentData(85); xorBitMap(12)(82) := currentData(82); xorBitMap(12)(81) := currentData(81); xorBitMap(12)(77) := currentData(77); xorBitMap(12)(75) := currentData(75); xorBitMap(12)(74) := currentData(74); xorBitMap(12)(73) := currentData(73); xorBitMap(12)(71) := currentData(71); xorBitMap(12)(69) := currentData(69); xorBitMap(12)(68) := currentData(68); xorBitMap(12)(63) := currentData(63); xorBitMap(12)(61) := currentData(61); xorBitMap(12)(59) := currentData(59); xorBitMap(12)(57) := currentData(57); xorBitMap(12)(56) := currentData(56); xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(161) := previousCrc(1); xorBitMap(12)(162) := previousCrc(2); xorBitMap(12)(163) := previousCrc(3); xorBitMap(12)(165) := previousCrc(5); xorBitMap(12)(169) := previousCrc(9); xorBitMap(12)(170) := previousCrc(10); xorBitMap(12)(173) := previousCrc(13); xorBitMap(12)(174) := previousCrc(14); xorBitMap(12)(175) := previousCrc(15); xorBitMap(12)(179) := previousCrc(19); xorBitMap(12)(180) := previousCrc(20); xorBitMap(12)(182) := previousCrc(22); xorBitMap(12)(184) := previousCrc(24); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(186) := previousCrc(26); xorBitMap(12)(189) := previousCrc(29); xorBitMap(12)(190) := previousCrc(30); 
      xorBitMap(13)(103) := currentData(103); xorBitMap(13)(102) := currentData(102); xorBitMap(13)(99) := currentData(99); xorBitMap(13)(98) := currentData(98); xorBitMap(13)(97) := currentData(97); xorBitMap(13)(95) := currentData(95); xorBitMap(13)(93) := currentData(93); xorBitMap(13)(92) := currentData(92); xorBitMap(13)(88) := currentData(88); xorBitMap(13)(87) := currentData(87); xorBitMap(13)(86) := currentData(86); xorBitMap(13)(83) := currentData(83); xorBitMap(13)(82) := currentData(82); xorBitMap(13)(78) := currentData(78); xorBitMap(13)(76) := currentData(76); xorBitMap(13)(75) := currentData(75); xorBitMap(13)(74) := currentData(74); xorBitMap(13)(72) := currentData(72); xorBitMap(13)(70) := currentData(70); xorBitMap(13)(69) := currentData(69); xorBitMap(13)(64) := currentData(64); xorBitMap(13)(62) := currentData(62); xorBitMap(13)(60) := currentData(60); xorBitMap(13)(58) := currentData(58); xorBitMap(13)(57) := currentData(57); xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(160) := previousCrc(0); xorBitMap(13)(162) := previousCrc(2); xorBitMap(13)(163) := previousCrc(3); xorBitMap(13)(164) := previousCrc(4); xorBitMap(13)(166) := previousCrc(6); xorBitMap(13)(170) := previousCrc(10); xorBitMap(13)(171) := previousCrc(11); xorBitMap(13)(174) := previousCrc(14); xorBitMap(13)(175) := previousCrc(15); xorBitMap(13)(176) := previousCrc(16); xorBitMap(13)(180) := previousCrc(20); xorBitMap(13)(181) := previousCrc(21); xorBitMap(13)(183) := previousCrc(23); xorBitMap(13)(185) := previousCrc(25); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(187) := previousCrc(27); xorBitMap(13)(190) := previousCrc(30); xorBitMap(13)(191) := previousCrc(31); 
      xorBitMap(14)(103) := currentData(103); xorBitMap(14)(100) := currentData(100); xorBitMap(14)(99) := currentData(99); xorBitMap(14)(98) := currentData(98); xorBitMap(14)(96) := currentData(96); xorBitMap(14)(94) := currentData(94); xorBitMap(14)(93) := currentData(93); xorBitMap(14)(89) := currentData(89); xorBitMap(14)(88) := currentData(88); xorBitMap(14)(87) := currentData(87); xorBitMap(14)(84) := currentData(84); xorBitMap(14)(83) := currentData(83); xorBitMap(14)(79) := currentData(79); xorBitMap(14)(77) := currentData(77); xorBitMap(14)(76) := currentData(76); xorBitMap(14)(75) := currentData(75); xorBitMap(14)(73) := currentData(73); xorBitMap(14)(71) := currentData(71); xorBitMap(14)(70) := currentData(70); xorBitMap(14)(65) := currentData(65); xorBitMap(14)(63) := currentData(63); xorBitMap(14)(61) := currentData(61); xorBitMap(14)(59) := currentData(59); xorBitMap(14)(58) := currentData(58); xorBitMap(14)(56) := currentData(56); xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(161) := previousCrc(1); xorBitMap(14)(163) := previousCrc(3); xorBitMap(14)(164) := previousCrc(4); xorBitMap(14)(165) := previousCrc(5); xorBitMap(14)(167) := previousCrc(7); xorBitMap(14)(171) := previousCrc(11); xorBitMap(14)(172) := previousCrc(12); xorBitMap(14)(175) := previousCrc(15); xorBitMap(14)(176) := previousCrc(16); xorBitMap(14)(177) := previousCrc(17); xorBitMap(14)(181) := previousCrc(21); xorBitMap(14)(182) := previousCrc(22); xorBitMap(14)(184) := previousCrc(24); xorBitMap(14)(186) := previousCrc(26); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(188) := previousCrc(28); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(101) := currentData(101); xorBitMap(15)(100) := currentData(100); xorBitMap(15)(99) := currentData(99); xorBitMap(15)(97) := currentData(97); xorBitMap(15)(95) := currentData(95); xorBitMap(15)(94) := currentData(94); xorBitMap(15)(90) := currentData(90); xorBitMap(15)(89) := currentData(89); xorBitMap(15)(88) := currentData(88); xorBitMap(15)(85) := currentData(85); xorBitMap(15)(84) := currentData(84); xorBitMap(15)(80) := currentData(80); xorBitMap(15)(78) := currentData(78); xorBitMap(15)(77) := currentData(77); xorBitMap(15)(76) := currentData(76); xorBitMap(15)(74) := currentData(74); xorBitMap(15)(72) := currentData(72); xorBitMap(15)(71) := currentData(71); xorBitMap(15)(66) := currentData(66); xorBitMap(15)(64) := currentData(64); xorBitMap(15)(62) := currentData(62); xorBitMap(15)(60) := currentData(60); xorBitMap(15)(59) := currentData(59); xorBitMap(15)(57) := currentData(57); xorBitMap(15)(56) := currentData(56); xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(160) := previousCrc(0); xorBitMap(15)(162) := previousCrc(2); xorBitMap(15)(164) := previousCrc(4); xorBitMap(15)(165) := previousCrc(5); xorBitMap(15)(166) := previousCrc(6); xorBitMap(15)(168) := previousCrc(8); xorBitMap(15)(172) := previousCrc(12); xorBitMap(15)(173) := previousCrc(13); xorBitMap(15)(176) := previousCrc(16); xorBitMap(15)(177) := previousCrc(17); xorBitMap(15)(178) := previousCrc(18); xorBitMap(15)(182) := previousCrc(22); xorBitMap(15)(183) := previousCrc(23); xorBitMap(15)(185) := previousCrc(25); xorBitMap(15)(187) := previousCrc(27); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(189) := previousCrc(29); 
      xorBitMap(16)(103) := currentData(103); xorBitMap(16)(102) := currentData(102); xorBitMap(16)(100) := currentData(100); xorBitMap(16)(99) := currentData(99); xorBitMap(16)(97) := currentData(97); xorBitMap(16)(94) := currentData(94); xorBitMap(16)(91) := currentData(91); xorBitMap(16)(90) := currentData(90); xorBitMap(16)(89) := currentData(89); xorBitMap(16)(87) := currentData(87); xorBitMap(16)(86) := currentData(86); xorBitMap(16)(84) := currentData(84); xorBitMap(16)(83) := currentData(83); xorBitMap(16)(82) := currentData(82); xorBitMap(16)(78) := currentData(78); xorBitMap(16)(77) := currentData(77); xorBitMap(16)(75) := currentData(75); xorBitMap(16)(68) := currentData(68); xorBitMap(16)(66) := currentData(66); xorBitMap(16)(57) := currentData(57); xorBitMap(16)(56) := currentData(56); xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(163) := previousCrc(3); xorBitMap(16)(165) := previousCrc(5); xorBitMap(16)(166) := previousCrc(6); xorBitMap(16)(170) := previousCrc(10); xorBitMap(16)(171) := previousCrc(11); xorBitMap(16)(172) := previousCrc(12); xorBitMap(16)(174) := previousCrc(14); xorBitMap(16)(175) := previousCrc(15); xorBitMap(16)(177) := previousCrc(17); xorBitMap(16)(178) := previousCrc(18); xorBitMap(16)(179) := previousCrc(19); xorBitMap(16)(182) := previousCrc(22); xorBitMap(16)(185) := previousCrc(25); xorBitMap(16)(187) := previousCrc(27); xorBitMap(16)(188) := previousCrc(28); xorBitMap(16)(190) := previousCrc(30); xorBitMap(16)(191) := previousCrc(31); 
      xorBitMap(17)(103) := currentData(103); xorBitMap(17)(101) := currentData(101); xorBitMap(17)(100) := currentData(100); xorBitMap(17)(98) := currentData(98); xorBitMap(17)(95) := currentData(95); xorBitMap(17)(92) := currentData(92); xorBitMap(17)(91) := currentData(91); xorBitMap(17)(90) := currentData(90); xorBitMap(17)(88) := currentData(88); xorBitMap(17)(87) := currentData(87); xorBitMap(17)(85) := currentData(85); xorBitMap(17)(84) := currentData(84); xorBitMap(17)(83) := currentData(83); xorBitMap(17)(79) := currentData(79); xorBitMap(17)(78) := currentData(78); xorBitMap(17)(76) := currentData(76); xorBitMap(17)(69) := currentData(69); xorBitMap(17)(67) := currentData(67); xorBitMap(17)(58) := currentData(58); xorBitMap(17)(57) := currentData(57); xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(164) := previousCrc(4); xorBitMap(17)(166) := previousCrc(6); xorBitMap(17)(167) := previousCrc(7); xorBitMap(17)(171) := previousCrc(11); xorBitMap(17)(172) := previousCrc(12); xorBitMap(17)(173) := previousCrc(13); xorBitMap(17)(175) := previousCrc(15); xorBitMap(17)(176) := previousCrc(16); xorBitMap(17)(178) := previousCrc(18); xorBitMap(17)(179) := previousCrc(19); xorBitMap(17)(180) := previousCrc(20); xorBitMap(17)(183) := previousCrc(23); xorBitMap(17)(186) := previousCrc(26); xorBitMap(17)(188) := previousCrc(28); xorBitMap(17)(189) := previousCrc(29); xorBitMap(17)(191) := previousCrc(31); 
      xorBitMap(18)(102) := currentData(102); xorBitMap(18)(101) := currentData(101); xorBitMap(18)(99) := currentData(99); xorBitMap(18)(96) := currentData(96); xorBitMap(18)(93) := currentData(93); xorBitMap(18)(92) := currentData(92); xorBitMap(18)(91) := currentData(91); xorBitMap(18)(89) := currentData(89); xorBitMap(18)(88) := currentData(88); xorBitMap(18)(86) := currentData(86); xorBitMap(18)(85) := currentData(85); xorBitMap(18)(84) := currentData(84); xorBitMap(18)(80) := currentData(80); xorBitMap(18)(79) := currentData(79); xorBitMap(18)(77) := currentData(77); xorBitMap(18)(70) := currentData(70); xorBitMap(18)(68) := currentData(68); xorBitMap(18)(59) := currentData(59); xorBitMap(18)(58) := currentData(58); xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(165) := previousCrc(5); xorBitMap(18)(167) := previousCrc(7); xorBitMap(18)(168) := previousCrc(8); xorBitMap(18)(172) := previousCrc(12); xorBitMap(18)(173) := previousCrc(13); xorBitMap(18)(174) := previousCrc(14); xorBitMap(18)(176) := previousCrc(16); xorBitMap(18)(177) := previousCrc(17); xorBitMap(18)(179) := previousCrc(19); xorBitMap(18)(180) := previousCrc(20); xorBitMap(18)(181) := previousCrc(21); xorBitMap(18)(184) := previousCrc(24); xorBitMap(18)(187) := previousCrc(27); xorBitMap(18)(189) := previousCrc(29); xorBitMap(18)(190) := previousCrc(30); 
      xorBitMap(19)(103) := currentData(103); xorBitMap(19)(102) := currentData(102); xorBitMap(19)(100) := currentData(100); xorBitMap(19)(97) := currentData(97); xorBitMap(19)(94) := currentData(94); xorBitMap(19)(93) := currentData(93); xorBitMap(19)(92) := currentData(92); xorBitMap(19)(90) := currentData(90); xorBitMap(19)(89) := currentData(89); xorBitMap(19)(87) := currentData(87); xorBitMap(19)(86) := currentData(86); xorBitMap(19)(85) := currentData(85); xorBitMap(19)(81) := currentData(81); xorBitMap(19)(80) := currentData(80); xorBitMap(19)(78) := currentData(78); xorBitMap(19)(71) := currentData(71); xorBitMap(19)(69) := currentData(69); xorBitMap(19)(60) := currentData(60); xorBitMap(19)(59) := currentData(59); xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(166) := previousCrc(6); xorBitMap(19)(168) := previousCrc(8); xorBitMap(19)(169) := previousCrc(9); xorBitMap(19)(173) := previousCrc(13); xorBitMap(19)(174) := previousCrc(14); xorBitMap(19)(175) := previousCrc(15); xorBitMap(19)(177) := previousCrc(17); xorBitMap(19)(178) := previousCrc(18); xorBitMap(19)(180) := previousCrc(20); xorBitMap(19)(181) := previousCrc(21); xorBitMap(19)(182) := previousCrc(22); xorBitMap(19)(185) := previousCrc(25); xorBitMap(19)(188) := previousCrc(28); xorBitMap(19)(190) := previousCrc(30); xorBitMap(19)(191) := previousCrc(31); 
      xorBitMap(20)(103) := currentData(103); xorBitMap(20)(101) := currentData(101); xorBitMap(20)(98) := currentData(98); xorBitMap(20)(95) := currentData(95); xorBitMap(20)(94) := currentData(94); xorBitMap(20)(93) := currentData(93); xorBitMap(20)(91) := currentData(91); xorBitMap(20)(90) := currentData(90); xorBitMap(20)(88) := currentData(88); xorBitMap(20)(87) := currentData(87); xorBitMap(20)(86) := currentData(86); xorBitMap(20)(82) := currentData(82); xorBitMap(20)(81) := currentData(81); xorBitMap(20)(79) := currentData(79); xorBitMap(20)(72) := currentData(72); xorBitMap(20)(70) := currentData(70); xorBitMap(20)(61) := currentData(61); xorBitMap(20)(60) := currentData(60); xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(160) := previousCrc(0); xorBitMap(20)(167) := previousCrc(7); xorBitMap(20)(169) := previousCrc(9); xorBitMap(20)(170) := previousCrc(10); xorBitMap(20)(174) := previousCrc(14); xorBitMap(20)(175) := previousCrc(15); xorBitMap(20)(176) := previousCrc(16); xorBitMap(20)(178) := previousCrc(18); xorBitMap(20)(179) := previousCrc(19); xorBitMap(20)(181) := previousCrc(21); xorBitMap(20)(182) := previousCrc(22); xorBitMap(20)(183) := previousCrc(23); xorBitMap(20)(186) := previousCrc(26); xorBitMap(20)(189) := previousCrc(29); xorBitMap(20)(191) := previousCrc(31); 
      xorBitMap(21)(102) := currentData(102); xorBitMap(21)(99) := currentData(99); xorBitMap(21)(96) := currentData(96); xorBitMap(21)(95) := currentData(95); xorBitMap(21)(94) := currentData(94); xorBitMap(21)(92) := currentData(92); xorBitMap(21)(91) := currentData(91); xorBitMap(21)(89) := currentData(89); xorBitMap(21)(88) := currentData(88); xorBitMap(21)(87) := currentData(87); xorBitMap(21)(83) := currentData(83); xorBitMap(21)(82) := currentData(82); xorBitMap(21)(80) := currentData(80); xorBitMap(21)(73) := currentData(73); xorBitMap(21)(71) := currentData(71); xorBitMap(21)(62) := currentData(62); xorBitMap(21)(61) := currentData(61); xorBitMap(21)(56) := currentData(56); xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(161) := previousCrc(1); xorBitMap(21)(168) := previousCrc(8); xorBitMap(21)(170) := previousCrc(10); xorBitMap(21)(171) := previousCrc(11); xorBitMap(21)(175) := previousCrc(15); xorBitMap(21)(176) := previousCrc(16); xorBitMap(21)(177) := previousCrc(17); xorBitMap(21)(179) := previousCrc(19); xorBitMap(21)(180) := previousCrc(20); xorBitMap(21)(182) := previousCrc(22); xorBitMap(21)(183) := previousCrc(23); xorBitMap(21)(184) := previousCrc(24); xorBitMap(21)(187) := previousCrc(27); xorBitMap(21)(190) := previousCrc(30); 
      xorBitMap(22)(101) := currentData(101); xorBitMap(22)(100) := currentData(100); xorBitMap(22)(99) := currentData(99); xorBitMap(22)(98) := currentData(98); xorBitMap(22)(94) := currentData(94); xorBitMap(22)(93) := currentData(93); xorBitMap(22)(92) := currentData(92); xorBitMap(22)(90) := currentData(90); xorBitMap(22)(89) := currentData(89); xorBitMap(22)(88) := currentData(88); xorBitMap(22)(87) := currentData(87); xorBitMap(22)(85) := currentData(85); xorBitMap(22)(82) := currentData(82); xorBitMap(22)(79) := currentData(79); xorBitMap(22)(74) := currentData(74); xorBitMap(22)(73) := currentData(73); xorBitMap(22)(68) := currentData(68); xorBitMap(22)(67) := currentData(67); xorBitMap(22)(66) := currentData(66); xorBitMap(22)(65) := currentData(65); xorBitMap(22)(62) := currentData(62); xorBitMap(22)(61) := currentData(61); xorBitMap(22)(60) := currentData(60); xorBitMap(22)(58) := currentData(58); xorBitMap(22)(57) := currentData(57); xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(161) := previousCrc(1); xorBitMap(22)(162) := previousCrc(2); xorBitMap(22)(167) := previousCrc(7); xorBitMap(22)(170) := previousCrc(10); xorBitMap(22)(173) := previousCrc(13); xorBitMap(22)(175) := previousCrc(15); xorBitMap(22)(176) := previousCrc(16); xorBitMap(22)(177) := previousCrc(17); xorBitMap(22)(178) := previousCrc(18); xorBitMap(22)(180) := previousCrc(20); xorBitMap(22)(181) := previousCrc(21); xorBitMap(22)(182) := previousCrc(22); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(187) := previousCrc(27); xorBitMap(22)(188) := previousCrc(28); xorBitMap(22)(189) := previousCrc(29); 
      xorBitMap(23)(103) := currentData(103); xorBitMap(23)(102) := currentData(102); xorBitMap(23)(100) := currentData(100); xorBitMap(23)(98) := currentData(98); xorBitMap(23)(97) := currentData(97); xorBitMap(23)(96) := currentData(96); xorBitMap(23)(93) := currentData(93); xorBitMap(23)(91) := currentData(91); xorBitMap(23)(90) := currentData(90); xorBitMap(23)(89) := currentData(89); xorBitMap(23)(88) := currentData(88); xorBitMap(23)(87) := currentData(87); xorBitMap(23)(86) := currentData(86); xorBitMap(23)(85) := currentData(85); xorBitMap(23)(84) := currentData(84); xorBitMap(23)(82) := currentData(82); xorBitMap(23)(81) := currentData(81); xorBitMap(23)(80) := currentData(80); xorBitMap(23)(79) := currentData(79); xorBitMap(23)(75) := currentData(75); xorBitMap(23)(74) := currentData(74); xorBitMap(23)(73) := currentData(73); xorBitMap(23)(72) := currentData(72); xorBitMap(23)(69) := currentData(69); xorBitMap(23)(65) := currentData(65); xorBitMap(23)(62) := currentData(62); xorBitMap(23)(60) := currentData(60); xorBitMap(23)(59) := currentData(59); xorBitMap(23)(56) := currentData(56); xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(160) := previousCrc(0); xorBitMap(23)(161) := previousCrc(1); xorBitMap(23)(162) := previousCrc(2); xorBitMap(23)(163) := previousCrc(3); xorBitMap(23)(167) := previousCrc(7); xorBitMap(23)(168) := previousCrc(8); xorBitMap(23)(169) := previousCrc(9); xorBitMap(23)(170) := previousCrc(10); xorBitMap(23)(172) := previousCrc(12); xorBitMap(23)(173) := previousCrc(13); xorBitMap(23)(174) := previousCrc(14); xorBitMap(23)(175) := previousCrc(15); xorBitMap(23)(176) := previousCrc(16); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(178) := previousCrc(18); xorBitMap(23)(179) := previousCrc(19); xorBitMap(23)(181) := previousCrc(21); xorBitMap(23)(184) := previousCrc(24); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(186) := previousCrc(26); xorBitMap(23)(188) := previousCrc(28); xorBitMap(23)(190) := previousCrc(30); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(103) := currentData(103); xorBitMap(24)(101) := currentData(101); xorBitMap(24)(99) := currentData(99); xorBitMap(24)(98) := currentData(98); xorBitMap(24)(97) := currentData(97); xorBitMap(24)(94) := currentData(94); xorBitMap(24)(92) := currentData(92); xorBitMap(24)(91) := currentData(91); xorBitMap(24)(90) := currentData(90); xorBitMap(24)(89) := currentData(89); xorBitMap(24)(88) := currentData(88); xorBitMap(24)(87) := currentData(87); xorBitMap(24)(86) := currentData(86); xorBitMap(24)(85) := currentData(85); xorBitMap(24)(83) := currentData(83); xorBitMap(24)(82) := currentData(82); xorBitMap(24)(81) := currentData(81); xorBitMap(24)(80) := currentData(80); xorBitMap(24)(76) := currentData(76); xorBitMap(24)(75) := currentData(75); xorBitMap(24)(74) := currentData(74); xorBitMap(24)(73) := currentData(73); xorBitMap(24)(70) := currentData(70); xorBitMap(24)(66) := currentData(66); xorBitMap(24)(63) := currentData(63); xorBitMap(24)(61) := currentData(61); xorBitMap(24)(60) := currentData(60); xorBitMap(24)(57) := currentData(57); xorBitMap(24)(56) := currentData(56); xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(161) := previousCrc(1); xorBitMap(24)(162) := previousCrc(2); xorBitMap(24)(163) := previousCrc(3); xorBitMap(24)(164) := previousCrc(4); xorBitMap(24)(168) := previousCrc(8); xorBitMap(24)(169) := previousCrc(9); xorBitMap(24)(170) := previousCrc(10); xorBitMap(24)(171) := previousCrc(11); xorBitMap(24)(173) := previousCrc(13); xorBitMap(24)(174) := previousCrc(14); xorBitMap(24)(175) := previousCrc(15); xorBitMap(24)(176) := previousCrc(16); xorBitMap(24)(177) := previousCrc(17); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(179) := previousCrc(19); xorBitMap(24)(180) := previousCrc(20); xorBitMap(24)(182) := previousCrc(22); xorBitMap(24)(185) := previousCrc(25); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(187) := previousCrc(27); xorBitMap(24)(189) := previousCrc(29); xorBitMap(24)(191) := previousCrc(31); 
      xorBitMap(25)(102) := currentData(102); xorBitMap(25)(100) := currentData(100); xorBitMap(25)(99) := currentData(99); xorBitMap(25)(98) := currentData(98); xorBitMap(25)(95) := currentData(95); xorBitMap(25)(93) := currentData(93); xorBitMap(25)(92) := currentData(92); xorBitMap(25)(91) := currentData(91); xorBitMap(25)(90) := currentData(90); xorBitMap(25)(89) := currentData(89); xorBitMap(25)(88) := currentData(88); xorBitMap(25)(87) := currentData(87); xorBitMap(25)(86) := currentData(86); xorBitMap(25)(84) := currentData(84); xorBitMap(25)(83) := currentData(83); xorBitMap(25)(82) := currentData(82); xorBitMap(25)(81) := currentData(81); xorBitMap(25)(77) := currentData(77); xorBitMap(25)(76) := currentData(76); xorBitMap(25)(75) := currentData(75); xorBitMap(25)(74) := currentData(74); xorBitMap(25)(71) := currentData(71); xorBitMap(25)(67) := currentData(67); xorBitMap(25)(64) := currentData(64); xorBitMap(25)(62) := currentData(62); xorBitMap(25)(61) := currentData(61); xorBitMap(25)(58) := currentData(58); xorBitMap(25)(57) := currentData(57); xorBitMap(25)(56) := currentData(56); xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(162) := previousCrc(2); xorBitMap(25)(163) := previousCrc(3); xorBitMap(25)(164) := previousCrc(4); xorBitMap(25)(165) := previousCrc(5); xorBitMap(25)(169) := previousCrc(9); xorBitMap(25)(170) := previousCrc(10); xorBitMap(25)(171) := previousCrc(11); xorBitMap(25)(172) := previousCrc(12); xorBitMap(25)(174) := previousCrc(14); xorBitMap(25)(175) := previousCrc(15); xorBitMap(25)(176) := previousCrc(16); xorBitMap(25)(177) := previousCrc(17); xorBitMap(25)(178) := previousCrc(18); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(180) := previousCrc(20); xorBitMap(25)(181) := previousCrc(21); xorBitMap(25)(183) := previousCrc(23); xorBitMap(25)(186) := previousCrc(26); xorBitMap(25)(187) := previousCrc(27); xorBitMap(25)(188) := previousCrc(28); xorBitMap(25)(190) := previousCrc(30); 
      xorBitMap(26)(100) := currentData(100); xorBitMap(26)(98) := currentData(98); xorBitMap(26)(97) := currentData(97); xorBitMap(26)(95) := currentData(95); xorBitMap(26)(93) := currentData(93); xorBitMap(26)(92) := currentData(92); xorBitMap(26)(91) := currentData(91); xorBitMap(26)(90) := currentData(90); xorBitMap(26)(89) := currentData(89); xorBitMap(26)(88) := currentData(88); xorBitMap(26)(81) := currentData(81); xorBitMap(26)(79) := currentData(79); xorBitMap(26)(78) := currentData(78); xorBitMap(26)(77) := currentData(77); xorBitMap(26)(76) := currentData(76); xorBitMap(26)(75) := currentData(75); xorBitMap(26)(73) := currentData(73); xorBitMap(26)(67) := currentData(67); xorBitMap(26)(66) := currentData(66); xorBitMap(26)(62) := currentData(62); xorBitMap(26)(61) := currentData(61); xorBitMap(26)(60) := currentData(60); xorBitMap(26)(59) := currentData(59); xorBitMap(26)(57) := currentData(57); xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(161) := previousCrc(1); xorBitMap(26)(163) := previousCrc(3); xorBitMap(26)(164) := previousCrc(4); xorBitMap(26)(165) := previousCrc(5); xorBitMap(26)(166) := previousCrc(6); xorBitMap(26)(167) := previousCrc(7); xorBitMap(26)(169) := previousCrc(9); xorBitMap(26)(176) := previousCrc(16); xorBitMap(26)(177) := previousCrc(17); xorBitMap(26)(178) := previousCrc(18); xorBitMap(26)(179) := previousCrc(19); xorBitMap(26)(180) := previousCrc(20); xorBitMap(26)(181) := previousCrc(21); xorBitMap(26)(183) := previousCrc(23); xorBitMap(26)(185) := previousCrc(25); xorBitMap(26)(186) := previousCrc(26); xorBitMap(26)(188) := previousCrc(28); 
      xorBitMap(27)(101) := currentData(101); xorBitMap(27)(99) := currentData(99); xorBitMap(27)(98) := currentData(98); xorBitMap(27)(96) := currentData(96); xorBitMap(27)(94) := currentData(94); xorBitMap(27)(93) := currentData(93); xorBitMap(27)(92) := currentData(92); xorBitMap(27)(91) := currentData(91); xorBitMap(27)(90) := currentData(90); xorBitMap(27)(89) := currentData(89); xorBitMap(27)(82) := currentData(82); xorBitMap(27)(80) := currentData(80); xorBitMap(27)(79) := currentData(79); xorBitMap(27)(78) := currentData(78); xorBitMap(27)(77) := currentData(77); xorBitMap(27)(76) := currentData(76); xorBitMap(27)(74) := currentData(74); xorBitMap(27)(68) := currentData(68); xorBitMap(27)(67) := currentData(67); xorBitMap(27)(63) := currentData(63); xorBitMap(27)(62) := currentData(62); xorBitMap(27)(61) := currentData(61); xorBitMap(27)(60) := currentData(60); xorBitMap(27)(58) := currentData(58); xorBitMap(27)(56) := currentData(56); xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(162) := previousCrc(2); xorBitMap(27)(164) := previousCrc(4); xorBitMap(27)(165) := previousCrc(5); xorBitMap(27)(166) := previousCrc(6); xorBitMap(27)(167) := previousCrc(7); xorBitMap(27)(168) := previousCrc(8); xorBitMap(27)(170) := previousCrc(10); xorBitMap(27)(177) := previousCrc(17); xorBitMap(27)(178) := previousCrc(18); xorBitMap(27)(179) := previousCrc(19); xorBitMap(27)(180) := previousCrc(20); xorBitMap(27)(181) := previousCrc(21); xorBitMap(27)(182) := previousCrc(22); xorBitMap(27)(184) := previousCrc(24); xorBitMap(27)(186) := previousCrc(26); xorBitMap(27)(187) := previousCrc(27); xorBitMap(27)(189) := previousCrc(29); 
      xorBitMap(28)(102) := currentData(102); xorBitMap(28)(100) := currentData(100); xorBitMap(28)(99) := currentData(99); xorBitMap(28)(97) := currentData(97); xorBitMap(28)(95) := currentData(95); xorBitMap(28)(94) := currentData(94); xorBitMap(28)(93) := currentData(93); xorBitMap(28)(92) := currentData(92); xorBitMap(28)(91) := currentData(91); xorBitMap(28)(90) := currentData(90); xorBitMap(28)(83) := currentData(83); xorBitMap(28)(81) := currentData(81); xorBitMap(28)(80) := currentData(80); xorBitMap(28)(79) := currentData(79); xorBitMap(28)(78) := currentData(78); xorBitMap(28)(77) := currentData(77); xorBitMap(28)(75) := currentData(75); xorBitMap(28)(69) := currentData(69); xorBitMap(28)(68) := currentData(68); xorBitMap(28)(64) := currentData(64); xorBitMap(28)(63) := currentData(63); xorBitMap(28)(62) := currentData(62); xorBitMap(28)(61) := currentData(61); xorBitMap(28)(59) := currentData(59); xorBitMap(28)(57) := currentData(57); xorBitMap(28)(56) := currentData(56); xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(163) := previousCrc(3); xorBitMap(28)(165) := previousCrc(5); xorBitMap(28)(166) := previousCrc(6); xorBitMap(28)(167) := previousCrc(7); xorBitMap(28)(168) := previousCrc(8); xorBitMap(28)(169) := previousCrc(9); xorBitMap(28)(171) := previousCrc(11); xorBitMap(28)(178) := previousCrc(18); xorBitMap(28)(179) := previousCrc(19); xorBitMap(28)(180) := previousCrc(20); xorBitMap(28)(181) := previousCrc(21); xorBitMap(28)(182) := previousCrc(22); xorBitMap(28)(183) := previousCrc(23); xorBitMap(28)(185) := previousCrc(25); xorBitMap(28)(187) := previousCrc(27); xorBitMap(28)(188) := previousCrc(28); xorBitMap(28)(190) := previousCrc(30); 
      xorBitMap(29)(103) := currentData(103); xorBitMap(29)(101) := currentData(101); xorBitMap(29)(100) := currentData(100); xorBitMap(29)(98) := currentData(98); xorBitMap(29)(96) := currentData(96); xorBitMap(29)(95) := currentData(95); xorBitMap(29)(94) := currentData(94); xorBitMap(29)(93) := currentData(93); xorBitMap(29)(92) := currentData(92); xorBitMap(29)(91) := currentData(91); xorBitMap(29)(84) := currentData(84); xorBitMap(29)(82) := currentData(82); xorBitMap(29)(81) := currentData(81); xorBitMap(29)(80) := currentData(80); xorBitMap(29)(79) := currentData(79); xorBitMap(29)(78) := currentData(78); xorBitMap(29)(76) := currentData(76); xorBitMap(29)(70) := currentData(70); xorBitMap(29)(69) := currentData(69); xorBitMap(29)(65) := currentData(65); xorBitMap(29)(64) := currentData(64); xorBitMap(29)(63) := currentData(63); xorBitMap(29)(62) := currentData(62); xorBitMap(29)(60) := currentData(60); xorBitMap(29)(58) := currentData(58); xorBitMap(29)(57) := currentData(57); xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(164) := previousCrc(4); xorBitMap(29)(166) := previousCrc(6); xorBitMap(29)(167) := previousCrc(7); xorBitMap(29)(168) := previousCrc(8); xorBitMap(29)(169) := previousCrc(9); xorBitMap(29)(170) := previousCrc(10); xorBitMap(29)(172) := previousCrc(12); xorBitMap(29)(179) := previousCrc(19); xorBitMap(29)(180) := previousCrc(20); xorBitMap(29)(181) := previousCrc(21); xorBitMap(29)(182) := previousCrc(22); xorBitMap(29)(183) := previousCrc(23); xorBitMap(29)(184) := previousCrc(24); xorBitMap(29)(186) := previousCrc(26); xorBitMap(29)(188) := previousCrc(28); xorBitMap(29)(189) := previousCrc(29); xorBitMap(29)(191) := previousCrc(31); 
      xorBitMap(30)(102) := currentData(102); xorBitMap(30)(101) := currentData(101); xorBitMap(30)(99) := currentData(99); xorBitMap(30)(97) := currentData(97); xorBitMap(30)(96) := currentData(96); xorBitMap(30)(95) := currentData(95); xorBitMap(30)(94) := currentData(94); xorBitMap(30)(93) := currentData(93); xorBitMap(30)(92) := currentData(92); xorBitMap(30)(85) := currentData(85); xorBitMap(30)(83) := currentData(83); xorBitMap(30)(82) := currentData(82); xorBitMap(30)(81) := currentData(81); xorBitMap(30)(80) := currentData(80); xorBitMap(30)(79) := currentData(79); xorBitMap(30)(77) := currentData(77); xorBitMap(30)(71) := currentData(71); xorBitMap(30)(70) := currentData(70); xorBitMap(30)(66) := currentData(66); xorBitMap(30)(65) := currentData(65); xorBitMap(30)(64) := currentData(64); xorBitMap(30)(63) := currentData(63); xorBitMap(30)(61) := currentData(61); xorBitMap(30)(59) := currentData(59); xorBitMap(30)(58) := currentData(58); xorBitMap(30)(56) := currentData(56); xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(165) := previousCrc(5); xorBitMap(30)(167) := previousCrc(7); xorBitMap(30)(168) := previousCrc(8); xorBitMap(30)(169) := previousCrc(9); xorBitMap(30)(170) := previousCrc(10); xorBitMap(30)(171) := previousCrc(11); xorBitMap(30)(173) := previousCrc(13); xorBitMap(30)(180) := previousCrc(20); xorBitMap(30)(181) := previousCrc(21); xorBitMap(30)(182) := previousCrc(22); xorBitMap(30)(183) := previousCrc(23); xorBitMap(30)(184) := previousCrc(24); xorBitMap(30)(185) := previousCrc(25); xorBitMap(30)(187) := previousCrc(27); xorBitMap(30)(189) := previousCrc(29); xorBitMap(30)(190) := previousCrc(30); 
      xorBitMap(31)(103) := currentData(103); xorBitMap(31)(102) := currentData(102); xorBitMap(31)(100) := currentData(100); xorBitMap(31)(98) := currentData(98); xorBitMap(31)(97) := currentData(97); xorBitMap(31)(96) := currentData(96); xorBitMap(31)(95) := currentData(95); xorBitMap(31)(94) := currentData(94); xorBitMap(31)(93) := currentData(93); xorBitMap(31)(86) := currentData(86); xorBitMap(31)(84) := currentData(84); xorBitMap(31)(83) := currentData(83); xorBitMap(31)(82) := currentData(82); xorBitMap(31)(81) := currentData(81); xorBitMap(31)(80) := currentData(80); xorBitMap(31)(78) := currentData(78); xorBitMap(31)(72) := currentData(72); xorBitMap(31)(71) := currentData(71); xorBitMap(31)(67) := currentData(67); xorBitMap(31)(66) := currentData(66); xorBitMap(31)(65) := currentData(65); xorBitMap(31)(64) := currentData(64); xorBitMap(31)(62) := currentData(62); xorBitMap(31)(60) := currentData(60); xorBitMap(31)(59) := currentData(59); xorBitMap(31)(57) := currentData(57); xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(160) := previousCrc(0); xorBitMap(31)(166) := previousCrc(6); xorBitMap(31)(168) := previousCrc(8); xorBitMap(31)(169) := previousCrc(9); xorBitMap(31)(170) := previousCrc(10); xorBitMap(31)(171) := previousCrc(11); xorBitMap(31)(172) := previousCrc(12); xorBitMap(31)(174) := previousCrc(14); xorBitMap(31)(181) := previousCrc(21); xorBitMap(31)(182) := previousCrc(22); xorBitMap(31)(183) := previousCrc(23); xorBitMap(31)(184) := previousCrc(24); xorBitMap(31)(185) := previousCrc(25); xorBitMap(31)(186) := previousCrc(26); xorBitMap(31)(188) := previousCrc(28); xorBitMap(31)(190) := previousCrc(30); xorBitMap(31)(191) := previousCrc(31); 
   end procedure;

   procedure xorBitMap14Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(111 downto 0)) is 
   begin
      xorBitMap(0)(111) := currentData(111); xorBitMap(0)(110) := currentData(110); xorBitMap(0)(106) := currentData(106); xorBitMap(0)(104) := currentData(104); xorBitMap(0)(103) := currentData(103); xorBitMap(0)(101) := currentData(101); xorBitMap(0)(99) := currentData(99); xorBitMap(0)(98) := currentData(98); xorBitMap(0)(97) := currentData(97); xorBitMap(0)(96) := currentData(96); xorBitMap(0)(95) := currentData(95); xorBitMap(0)(94) := currentData(94); xorBitMap(0)(87) := currentData(87); xorBitMap(0)(85) := currentData(85); xorBitMap(0)(84) := currentData(84); xorBitMap(0)(83) := currentData(83); xorBitMap(0)(82) := currentData(82); xorBitMap(0)(81) := currentData(81); xorBitMap(0)(79) := currentData(79); xorBitMap(0)(73) := currentData(73); xorBitMap(0)(72) := currentData(72); xorBitMap(0)(68) := currentData(68); xorBitMap(0)(67) := currentData(67); xorBitMap(0)(66) := currentData(66); xorBitMap(0)(65) := currentData(65); xorBitMap(0)(63) := currentData(63); xorBitMap(0)(61) := currentData(61); xorBitMap(0)(60) := currentData(60); xorBitMap(0)(58) := currentData(58); xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(161) := previousCrc(1); xorBitMap(0)(162) := previousCrc(2); xorBitMap(0)(163) := previousCrc(3); xorBitMap(0)(164) := previousCrc(4); xorBitMap(0)(165) := previousCrc(5); xorBitMap(0)(167) := previousCrc(7); xorBitMap(0)(174) := previousCrc(14); xorBitMap(0)(175) := previousCrc(15); xorBitMap(0)(176) := previousCrc(16); xorBitMap(0)(177) := previousCrc(17); xorBitMap(0)(178) := previousCrc(18); xorBitMap(0)(179) := previousCrc(19); xorBitMap(0)(181) := previousCrc(21); xorBitMap(0)(183) := previousCrc(23); xorBitMap(0)(184) := previousCrc(24); xorBitMap(0)(186) := previousCrc(26); xorBitMap(0)(190) := previousCrc(30); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(110) := currentData(110); xorBitMap(1)(107) := currentData(107); xorBitMap(1)(106) := currentData(106); xorBitMap(1)(105) := currentData(105); xorBitMap(1)(103) := currentData(103); xorBitMap(1)(102) := currentData(102); xorBitMap(1)(101) := currentData(101); xorBitMap(1)(100) := currentData(100); xorBitMap(1)(94) := currentData(94); xorBitMap(1)(88) := currentData(88); xorBitMap(1)(87) := currentData(87); xorBitMap(1)(86) := currentData(86); xorBitMap(1)(81) := currentData(81); xorBitMap(1)(80) := currentData(80); xorBitMap(1)(79) := currentData(79); xorBitMap(1)(74) := currentData(74); xorBitMap(1)(72) := currentData(72); xorBitMap(1)(69) := currentData(69); xorBitMap(1)(65) := currentData(65); xorBitMap(1)(64) := currentData(64); xorBitMap(1)(63) := currentData(63); xorBitMap(1)(62) := currentData(62); xorBitMap(1)(60) := currentData(60); xorBitMap(1)(59) := currentData(59); xorBitMap(1)(58) := currentData(58); xorBitMap(1)(56) := currentData(56); xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(160) := previousCrc(0); xorBitMap(1)(161) := previousCrc(1); xorBitMap(1)(166) := previousCrc(6); xorBitMap(1)(167) := previousCrc(7); xorBitMap(1)(168) := previousCrc(8); xorBitMap(1)(174) := previousCrc(14); xorBitMap(1)(180) := previousCrc(20); xorBitMap(1)(181) := previousCrc(21); xorBitMap(1)(182) := previousCrc(22); xorBitMap(1)(183) := previousCrc(23); xorBitMap(1)(185) := previousCrc(25); xorBitMap(1)(186) := previousCrc(26); xorBitMap(1)(187) := previousCrc(27); xorBitMap(1)(190) := previousCrc(30); 
      xorBitMap(2)(110) := currentData(110); xorBitMap(2)(108) := currentData(108); xorBitMap(2)(107) := currentData(107); xorBitMap(2)(102) := currentData(102); xorBitMap(2)(99) := currentData(99); xorBitMap(2)(98) := currentData(98); xorBitMap(2)(97) := currentData(97); xorBitMap(2)(96) := currentData(96); xorBitMap(2)(94) := currentData(94); xorBitMap(2)(89) := currentData(89); xorBitMap(2)(88) := currentData(88); xorBitMap(2)(85) := currentData(85); xorBitMap(2)(84) := currentData(84); xorBitMap(2)(83) := currentData(83); xorBitMap(2)(80) := currentData(80); xorBitMap(2)(79) := currentData(79); xorBitMap(2)(75) := currentData(75); xorBitMap(2)(72) := currentData(72); xorBitMap(2)(70) := currentData(70); xorBitMap(2)(68) := currentData(68); xorBitMap(2)(67) := currentData(67); xorBitMap(2)(64) := currentData(64); xorBitMap(2)(59) := currentData(59); xorBitMap(2)(58) := currentData(58); xorBitMap(2)(57) := currentData(57); xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(160) := previousCrc(0); xorBitMap(2)(163) := previousCrc(3); xorBitMap(2)(164) := previousCrc(4); xorBitMap(2)(165) := previousCrc(5); xorBitMap(2)(168) := previousCrc(8); xorBitMap(2)(169) := previousCrc(9); xorBitMap(2)(174) := previousCrc(14); xorBitMap(2)(176) := previousCrc(16); xorBitMap(2)(177) := previousCrc(17); xorBitMap(2)(178) := previousCrc(18); xorBitMap(2)(179) := previousCrc(19); xorBitMap(2)(182) := previousCrc(22); xorBitMap(2)(187) := previousCrc(27); xorBitMap(2)(188) := previousCrc(28); xorBitMap(2)(190) := previousCrc(30); 
      xorBitMap(3)(111) := currentData(111); xorBitMap(3)(109) := currentData(109); xorBitMap(3)(108) := currentData(108); xorBitMap(3)(103) := currentData(103); xorBitMap(3)(100) := currentData(100); xorBitMap(3)(99) := currentData(99); xorBitMap(3)(98) := currentData(98); xorBitMap(3)(97) := currentData(97); xorBitMap(3)(95) := currentData(95); xorBitMap(3)(90) := currentData(90); xorBitMap(3)(89) := currentData(89); xorBitMap(3)(86) := currentData(86); xorBitMap(3)(85) := currentData(85); xorBitMap(3)(84) := currentData(84); xorBitMap(3)(81) := currentData(81); xorBitMap(3)(80) := currentData(80); xorBitMap(3)(76) := currentData(76); xorBitMap(3)(73) := currentData(73); xorBitMap(3)(71) := currentData(71); xorBitMap(3)(69) := currentData(69); xorBitMap(3)(68) := currentData(68); xorBitMap(3)(65) := currentData(65); xorBitMap(3)(60) := currentData(60); xorBitMap(3)(59) := currentData(59); xorBitMap(3)(58) := currentData(58); xorBitMap(3)(56) := currentData(56); xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(160) := previousCrc(0); xorBitMap(3)(161) := previousCrc(1); xorBitMap(3)(164) := previousCrc(4); xorBitMap(3)(165) := previousCrc(5); xorBitMap(3)(166) := previousCrc(6); xorBitMap(3)(169) := previousCrc(9); xorBitMap(3)(170) := previousCrc(10); xorBitMap(3)(175) := previousCrc(15); xorBitMap(3)(177) := previousCrc(17); xorBitMap(3)(178) := previousCrc(18); xorBitMap(3)(179) := previousCrc(19); xorBitMap(3)(180) := previousCrc(20); xorBitMap(3)(183) := previousCrc(23); xorBitMap(3)(188) := previousCrc(28); xorBitMap(3)(189) := previousCrc(29); xorBitMap(3)(191) := previousCrc(31); 
      xorBitMap(4)(111) := currentData(111); xorBitMap(4)(109) := currentData(109); xorBitMap(4)(106) := currentData(106); xorBitMap(4)(103) := currentData(103); xorBitMap(4)(100) := currentData(100); xorBitMap(4)(97) := currentData(97); xorBitMap(4)(95) := currentData(95); xorBitMap(4)(94) := currentData(94); xorBitMap(4)(91) := currentData(91); xorBitMap(4)(90) := currentData(90); xorBitMap(4)(86) := currentData(86); xorBitMap(4)(84) := currentData(84); xorBitMap(4)(83) := currentData(83); xorBitMap(4)(79) := currentData(79); xorBitMap(4)(77) := currentData(77); xorBitMap(4)(74) := currentData(74); xorBitMap(4)(73) := currentData(73); xorBitMap(4)(70) := currentData(70); xorBitMap(4)(69) := currentData(69); xorBitMap(4)(68) := currentData(68); xorBitMap(4)(67) := currentData(67); xorBitMap(4)(65) := currentData(65); xorBitMap(4)(63) := currentData(63); xorBitMap(4)(59) := currentData(59); xorBitMap(4)(58) := currentData(58); xorBitMap(4)(57) := currentData(57); xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(163) := previousCrc(3); xorBitMap(4)(164) := previousCrc(4); xorBitMap(4)(166) := previousCrc(6); xorBitMap(4)(170) := previousCrc(10); xorBitMap(4)(171) := previousCrc(11); xorBitMap(4)(174) := previousCrc(14); xorBitMap(4)(175) := previousCrc(15); xorBitMap(4)(177) := previousCrc(17); xorBitMap(4)(180) := previousCrc(20); xorBitMap(4)(183) := previousCrc(23); xorBitMap(4)(186) := previousCrc(26); xorBitMap(4)(189) := previousCrc(29); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(111) := currentData(111); xorBitMap(5)(107) := currentData(107); xorBitMap(5)(106) := currentData(106); xorBitMap(5)(103) := currentData(103); xorBitMap(5)(99) := currentData(99); xorBitMap(5)(97) := currentData(97); xorBitMap(5)(94) := currentData(94); xorBitMap(5)(92) := currentData(92); xorBitMap(5)(91) := currentData(91); xorBitMap(5)(83) := currentData(83); xorBitMap(5)(82) := currentData(82); xorBitMap(5)(81) := currentData(81); xorBitMap(5)(80) := currentData(80); xorBitMap(5)(79) := currentData(79); xorBitMap(5)(78) := currentData(78); xorBitMap(5)(75) := currentData(75); xorBitMap(5)(74) := currentData(74); xorBitMap(5)(73) := currentData(73); xorBitMap(5)(72) := currentData(72); xorBitMap(5)(71) := currentData(71); xorBitMap(5)(70) := currentData(70); xorBitMap(5)(69) := currentData(69); xorBitMap(5)(67) := currentData(67); xorBitMap(5)(65) := currentData(65); xorBitMap(5)(64) := currentData(64); xorBitMap(5)(63) := currentData(63); xorBitMap(5)(61) := currentData(61); xorBitMap(5)(59) := currentData(59); xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(160) := previousCrc(0); xorBitMap(5)(161) := previousCrc(1); xorBitMap(5)(162) := previousCrc(2); xorBitMap(5)(163) := previousCrc(3); xorBitMap(5)(171) := previousCrc(11); xorBitMap(5)(172) := previousCrc(12); xorBitMap(5)(174) := previousCrc(14); xorBitMap(5)(177) := previousCrc(17); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(183) := previousCrc(23); xorBitMap(5)(186) := previousCrc(26); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(191) := previousCrc(31); 
      xorBitMap(6)(108) := currentData(108); xorBitMap(6)(107) := currentData(107); xorBitMap(6)(104) := currentData(104); xorBitMap(6)(100) := currentData(100); xorBitMap(6)(98) := currentData(98); xorBitMap(6)(95) := currentData(95); xorBitMap(6)(93) := currentData(93); xorBitMap(6)(92) := currentData(92); xorBitMap(6)(84) := currentData(84); xorBitMap(6)(83) := currentData(83); xorBitMap(6)(82) := currentData(82); xorBitMap(6)(81) := currentData(81); xorBitMap(6)(80) := currentData(80); xorBitMap(6)(79) := currentData(79); xorBitMap(6)(76) := currentData(76); xorBitMap(6)(75) := currentData(75); xorBitMap(6)(74) := currentData(74); xorBitMap(6)(73) := currentData(73); xorBitMap(6)(72) := currentData(72); xorBitMap(6)(71) := currentData(71); xorBitMap(6)(70) := currentData(70); xorBitMap(6)(68) := currentData(68); xorBitMap(6)(66) := currentData(66); xorBitMap(6)(65) := currentData(65); xorBitMap(6)(64) := currentData(64); xorBitMap(6)(62) := currentData(62); xorBitMap(6)(60) := currentData(60); xorBitMap(6)(56) := currentData(56); xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(160) := previousCrc(0); xorBitMap(6)(161) := previousCrc(1); xorBitMap(6)(162) := previousCrc(2); xorBitMap(6)(163) := previousCrc(3); xorBitMap(6)(164) := previousCrc(4); xorBitMap(6)(172) := previousCrc(12); xorBitMap(6)(173) := previousCrc(13); xorBitMap(6)(175) := previousCrc(15); xorBitMap(6)(178) := previousCrc(18); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(184) := previousCrc(24); xorBitMap(6)(187) := previousCrc(27); xorBitMap(6)(188) := previousCrc(28); 
      xorBitMap(7)(111) := currentData(111); xorBitMap(7)(110) := currentData(110); xorBitMap(7)(109) := currentData(109); xorBitMap(7)(108) := currentData(108); xorBitMap(7)(106) := currentData(106); xorBitMap(7)(105) := currentData(105); xorBitMap(7)(104) := currentData(104); xorBitMap(7)(103) := currentData(103); xorBitMap(7)(98) := currentData(98); xorBitMap(7)(97) := currentData(97); xorBitMap(7)(95) := currentData(95); xorBitMap(7)(93) := currentData(93); xorBitMap(7)(87) := currentData(87); xorBitMap(7)(80) := currentData(80); xorBitMap(7)(79) := currentData(79); xorBitMap(7)(77) := currentData(77); xorBitMap(7)(76) := currentData(76); xorBitMap(7)(75) := currentData(75); xorBitMap(7)(74) := currentData(74); xorBitMap(7)(71) := currentData(71); xorBitMap(7)(69) := currentData(69); xorBitMap(7)(68) := currentData(68); xorBitMap(7)(60) := currentData(60); xorBitMap(7)(58) := currentData(58); xorBitMap(7)(57) := currentData(57); xorBitMap(7)(56) := currentData(56); xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(160) := previousCrc(0); xorBitMap(7)(167) := previousCrc(7); xorBitMap(7)(173) := previousCrc(13); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(177) := previousCrc(17); xorBitMap(7)(178) := previousCrc(18); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(184) := previousCrc(24); xorBitMap(7)(185) := previousCrc(25); xorBitMap(7)(186) := previousCrc(26); xorBitMap(7)(188) := previousCrc(28); xorBitMap(7)(189) := previousCrc(29); xorBitMap(7)(190) := previousCrc(30); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(109) := currentData(109); xorBitMap(8)(107) := currentData(107); xorBitMap(8)(105) := currentData(105); xorBitMap(8)(103) := currentData(103); xorBitMap(8)(101) := currentData(101); xorBitMap(8)(97) := currentData(97); xorBitMap(8)(95) := currentData(95); xorBitMap(8)(88) := currentData(88); xorBitMap(8)(87) := currentData(87); xorBitMap(8)(85) := currentData(85); xorBitMap(8)(84) := currentData(84); xorBitMap(8)(83) := currentData(83); xorBitMap(8)(82) := currentData(82); xorBitMap(8)(80) := currentData(80); xorBitMap(8)(79) := currentData(79); xorBitMap(8)(78) := currentData(78); xorBitMap(8)(77) := currentData(77); xorBitMap(8)(76) := currentData(76); xorBitMap(8)(75) := currentData(75); xorBitMap(8)(73) := currentData(73); xorBitMap(8)(70) := currentData(70); xorBitMap(8)(69) := currentData(69); xorBitMap(8)(68) := currentData(68); xorBitMap(8)(67) := currentData(67); xorBitMap(8)(66) := currentData(66); xorBitMap(8)(65) := currentData(65); xorBitMap(8)(63) := currentData(63); xorBitMap(8)(60) := currentData(60); xorBitMap(8)(59) := currentData(59); xorBitMap(8)(57) := currentData(57); xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(160) := previousCrc(0); xorBitMap(8)(162) := previousCrc(2); xorBitMap(8)(163) := previousCrc(3); xorBitMap(8)(164) := previousCrc(4); xorBitMap(8)(165) := previousCrc(5); xorBitMap(8)(167) := previousCrc(7); xorBitMap(8)(168) := previousCrc(8); xorBitMap(8)(175) := previousCrc(15); xorBitMap(8)(177) := previousCrc(17); xorBitMap(8)(181) := previousCrc(21); xorBitMap(8)(183) := previousCrc(23); xorBitMap(8)(185) := previousCrc(25); xorBitMap(8)(187) := previousCrc(27); xorBitMap(8)(189) := previousCrc(29); 
      xorBitMap(9)(110) := currentData(110); xorBitMap(9)(108) := currentData(108); xorBitMap(9)(106) := currentData(106); xorBitMap(9)(104) := currentData(104); xorBitMap(9)(102) := currentData(102); xorBitMap(9)(98) := currentData(98); xorBitMap(9)(96) := currentData(96); xorBitMap(9)(89) := currentData(89); xorBitMap(9)(88) := currentData(88); xorBitMap(9)(86) := currentData(86); xorBitMap(9)(85) := currentData(85); xorBitMap(9)(84) := currentData(84); xorBitMap(9)(83) := currentData(83); xorBitMap(9)(81) := currentData(81); xorBitMap(9)(80) := currentData(80); xorBitMap(9)(79) := currentData(79); xorBitMap(9)(78) := currentData(78); xorBitMap(9)(77) := currentData(77); xorBitMap(9)(76) := currentData(76); xorBitMap(9)(74) := currentData(74); xorBitMap(9)(71) := currentData(71); xorBitMap(9)(70) := currentData(70); xorBitMap(9)(69) := currentData(69); xorBitMap(9)(68) := currentData(68); xorBitMap(9)(67) := currentData(67); xorBitMap(9)(66) := currentData(66); xorBitMap(9)(64) := currentData(64); xorBitMap(9)(61) := currentData(61); xorBitMap(9)(60) := currentData(60); xorBitMap(9)(58) := currentData(58); xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(160) := previousCrc(0); xorBitMap(9)(161) := previousCrc(1); xorBitMap(9)(163) := previousCrc(3); xorBitMap(9)(164) := previousCrc(4); xorBitMap(9)(165) := previousCrc(5); xorBitMap(9)(166) := previousCrc(6); xorBitMap(9)(168) := previousCrc(8); xorBitMap(9)(169) := previousCrc(9); xorBitMap(9)(176) := previousCrc(16); xorBitMap(9)(178) := previousCrc(18); xorBitMap(9)(182) := previousCrc(22); xorBitMap(9)(184) := previousCrc(24); xorBitMap(9)(186) := previousCrc(26); xorBitMap(9)(188) := previousCrc(28); xorBitMap(9)(190) := previousCrc(30); 
      xorBitMap(10)(110) := currentData(110); xorBitMap(10)(109) := currentData(109); xorBitMap(10)(107) := currentData(107); xorBitMap(10)(106) := currentData(106); xorBitMap(10)(105) := currentData(105); xorBitMap(10)(104) := currentData(104); xorBitMap(10)(101) := currentData(101); xorBitMap(10)(98) := currentData(98); xorBitMap(10)(96) := currentData(96); xorBitMap(10)(95) := currentData(95); xorBitMap(10)(94) := currentData(94); xorBitMap(10)(90) := currentData(90); xorBitMap(10)(89) := currentData(89); xorBitMap(10)(86) := currentData(86); xorBitMap(10)(83) := currentData(83); xorBitMap(10)(80) := currentData(80); xorBitMap(10)(78) := currentData(78); xorBitMap(10)(77) := currentData(77); xorBitMap(10)(75) := currentData(75); xorBitMap(10)(73) := currentData(73); xorBitMap(10)(71) := currentData(71); xorBitMap(10)(70) := currentData(70); xorBitMap(10)(69) := currentData(69); xorBitMap(10)(66) := currentData(66); xorBitMap(10)(63) := currentData(63); xorBitMap(10)(62) := currentData(62); xorBitMap(10)(60) := currentData(60); xorBitMap(10)(59) := currentData(59); xorBitMap(10)(58) := currentData(58); xorBitMap(10)(56) := currentData(56); xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(160) := previousCrc(0); xorBitMap(10)(163) := previousCrc(3); xorBitMap(10)(166) := previousCrc(6); xorBitMap(10)(169) := previousCrc(9); xorBitMap(10)(170) := previousCrc(10); xorBitMap(10)(174) := previousCrc(14); xorBitMap(10)(175) := previousCrc(15); xorBitMap(10)(176) := previousCrc(16); xorBitMap(10)(178) := previousCrc(18); xorBitMap(10)(181) := previousCrc(21); xorBitMap(10)(184) := previousCrc(24); xorBitMap(10)(185) := previousCrc(25); xorBitMap(10)(186) := previousCrc(26); xorBitMap(10)(187) := previousCrc(27); xorBitMap(10)(189) := previousCrc(29); xorBitMap(10)(190) := previousCrc(30); 
      xorBitMap(11)(108) := currentData(108); xorBitMap(11)(107) := currentData(107); xorBitMap(11)(105) := currentData(105); xorBitMap(11)(104) := currentData(104); xorBitMap(11)(103) := currentData(103); xorBitMap(11)(102) := currentData(102); xorBitMap(11)(101) := currentData(101); xorBitMap(11)(98) := currentData(98); xorBitMap(11)(94) := currentData(94); xorBitMap(11)(91) := currentData(91); xorBitMap(11)(90) := currentData(90); xorBitMap(11)(85) := currentData(85); xorBitMap(11)(83) := currentData(83); xorBitMap(11)(82) := currentData(82); xorBitMap(11)(78) := currentData(78); xorBitMap(11)(76) := currentData(76); xorBitMap(11)(74) := currentData(74); xorBitMap(11)(73) := currentData(73); xorBitMap(11)(71) := currentData(71); xorBitMap(11)(70) := currentData(70); xorBitMap(11)(68) := currentData(68); xorBitMap(11)(66) := currentData(66); xorBitMap(11)(65) := currentData(65); xorBitMap(11)(64) := currentData(64); xorBitMap(11)(59) := currentData(59); xorBitMap(11)(58) := currentData(58); xorBitMap(11)(57) := currentData(57); xorBitMap(11)(56) := currentData(56); xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(162) := previousCrc(2); xorBitMap(11)(163) := previousCrc(3); xorBitMap(11)(165) := previousCrc(5); xorBitMap(11)(170) := previousCrc(10); xorBitMap(11)(171) := previousCrc(11); xorBitMap(11)(174) := previousCrc(14); xorBitMap(11)(178) := previousCrc(18); xorBitMap(11)(181) := previousCrc(21); xorBitMap(11)(182) := previousCrc(22); xorBitMap(11)(183) := previousCrc(23); xorBitMap(11)(184) := previousCrc(24); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(187) := previousCrc(27); xorBitMap(11)(188) := previousCrc(28); 
      xorBitMap(12)(111) := currentData(111); xorBitMap(12)(110) := currentData(110); xorBitMap(12)(109) := currentData(109); xorBitMap(12)(108) := currentData(108); xorBitMap(12)(105) := currentData(105); xorBitMap(12)(102) := currentData(102); xorBitMap(12)(101) := currentData(101); xorBitMap(12)(98) := currentData(98); xorBitMap(12)(97) := currentData(97); xorBitMap(12)(96) := currentData(96); xorBitMap(12)(94) := currentData(94); xorBitMap(12)(92) := currentData(92); xorBitMap(12)(91) := currentData(91); xorBitMap(12)(87) := currentData(87); xorBitMap(12)(86) := currentData(86); xorBitMap(12)(85) := currentData(85); xorBitMap(12)(82) := currentData(82); xorBitMap(12)(81) := currentData(81); xorBitMap(12)(77) := currentData(77); xorBitMap(12)(75) := currentData(75); xorBitMap(12)(74) := currentData(74); xorBitMap(12)(73) := currentData(73); xorBitMap(12)(71) := currentData(71); xorBitMap(12)(69) := currentData(69); xorBitMap(12)(68) := currentData(68); xorBitMap(12)(63) := currentData(63); xorBitMap(12)(61) := currentData(61); xorBitMap(12)(59) := currentData(59); xorBitMap(12)(57) := currentData(57); xorBitMap(12)(56) := currentData(56); xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(161) := previousCrc(1); xorBitMap(12)(162) := previousCrc(2); xorBitMap(12)(165) := previousCrc(5); xorBitMap(12)(166) := previousCrc(6); xorBitMap(12)(167) := previousCrc(7); xorBitMap(12)(171) := previousCrc(11); xorBitMap(12)(172) := previousCrc(12); xorBitMap(12)(174) := previousCrc(14); xorBitMap(12)(176) := previousCrc(16); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(178) := previousCrc(18); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(182) := previousCrc(22); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(188) := previousCrc(28); xorBitMap(12)(189) := previousCrc(29); xorBitMap(12)(190) := previousCrc(30); xorBitMap(12)(191) := previousCrc(31); 
      xorBitMap(13)(111) := currentData(111); xorBitMap(13)(110) := currentData(110); xorBitMap(13)(109) := currentData(109); xorBitMap(13)(106) := currentData(106); xorBitMap(13)(103) := currentData(103); xorBitMap(13)(102) := currentData(102); xorBitMap(13)(99) := currentData(99); xorBitMap(13)(98) := currentData(98); xorBitMap(13)(97) := currentData(97); xorBitMap(13)(95) := currentData(95); xorBitMap(13)(93) := currentData(93); xorBitMap(13)(92) := currentData(92); xorBitMap(13)(88) := currentData(88); xorBitMap(13)(87) := currentData(87); xorBitMap(13)(86) := currentData(86); xorBitMap(13)(83) := currentData(83); xorBitMap(13)(82) := currentData(82); xorBitMap(13)(78) := currentData(78); xorBitMap(13)(76) := currentData(76); xorBitMap(13)(75) := currentData(75); xorBitMap(13)(74) := currentData(74); xorBitMap(13)(72) := currentData(72); xorBitMap(13)(70) := currentData(70); xorBitMap(13)(69) := currentData(69); xorBitMap(13)(64) := currentData(64); xorBitMap(13)(62) := currentData(62); xorBitMap(13)(60) := currentData(60); xorBitMap(13)(58) := currentData(58); xorBitMap(13)(57) := currentData(57); xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(162) := previousCrc(2); xorBitMap(13)(163) := previousCrc(3); xorBitMap(13)(166) := previousCrc(6); xorBitMap(13)(167) := previousCrc(7); xorBitMap(13)(168) := previousCrc(8); xorBitMap(13)(172) := previousCrc(12); xorBitMap(13)(173) := previousCrc(13); xorBitMap(13)(175) := previousCrc(15); xorBitMap(13)(177) := previousCrc(17); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(179) := previousCrc(19); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(183) := previousCrc(23); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(189) := previousCrc(29); xorBitMap(13)(190) := previousCrc(30); xorBitMap(13)(191) := previousCrc(31); 
      xorBitMap(14)(111) := currentData(111); xorBitMap(14)(110) := currentData(110); xorBitMap(14)(107) := currentData(107); xorBitMap(14)(104) := currentData(104); xorBitMap(14)(103) := currentData(103); xorBitMap(14)(100) := currentData(100); xorBitMap(14)(99) := currentData(99); xorBitMap(14)(98) := currentData(98); xorBitMap(14)(96) := currentData(96); xorBitMap(14)(94) := currentData(94); xorBitMap(14)(93) := currentData(93); xorBitMap(14)(89) := currentData(89); xorBitMap(14)(88) := currentData(88); xorBitMap(14)(87) := currentData(87); xorBitMap(14)(84) := currentData(84); xorBitMap(14)(83) := currentData(83); xorBitMap(14)(79) := currentData(79); xorBitMap(14)(77) := currentData(77); xorBitMap(14)(76) := currentData(76); xorBitMap(14)(75) := currentData(75); xorBitMap(14)(73) := currentData(73); xorBitMap(14)(71) := currentData(71); xorBitMap(14)(70) := currentData(70); xorBitMap(14)(65) := currentData(65); xorBitMap(14)(63) := currentData(63); xorBitMap(14)(61) := currentData(61); xorBitMap(14)(59) := currentData(59); xorBitMap(14)(58) := currentData(58); xorBitMap(14)(56) := currentData(56); xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(163) := previousCrc(3); xorBitMap(14)(164) := previousCrc(4); xorBitMap(14)(167) := previousCrc(7); xorBitMap(14)(168) := previousCrc(8); xorBitMap(14)(169) := previousCrc(9); xorBitMap(14)(173) := previousCrc(13); xorBitMap(14)(174) := previousCrc(14); xorBitMap(14)(176) := previousCrc(16); xorBitMap(14)(178) := previousCrc(18); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(180) := previousCrc(20); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(184) := previousCrc(24); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(190) := previousCrc(30); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(111) := currentData(111); xorBitMap(15)(108) := currentData(108); xorBitMap(15)(105) := currentData(105); xorBitMap(15)(104) := currentData(104); xorBitMap(15)(101) := currentData(101); xorBitMap(15)(100) := currentData(100); xorBitMap(15)(99) := currentData(99); xorBitMap(15)(97) := currentData(97); xorBitMap(15)(95) := currentData(95); xorBitMap(15)(94) := currentData(94); xorBitMap(15)(90) := currentData(90); xorBitMap(15)(89) := currentData(89); xorBitMap(15)(88) := currentData(88); xorBitMap(15)(85) := currentData(85); xorBitMap(15)(84) := currentData(84); xorBitMap(15)(80) := currentData(80); xorBitMap(15)(78) := currentData(78); xorBitMap(15)(77) := currentData(77); xorBitMap(15)(76) := currentData(76); xorBitMap(15)(74) := currentData(74); xorBitMap(15)(72) := currentData(72); xorBitMap(15)(71) := currentData(71); xorBitMap(15)(66) := currentData(66); xorBitMap(15)(64) := currentData(64); xorBitMap(15)(62) := currentData(62); xorBitMap(15)(60) := currentData(60); xorBitMap(15)(59) := currentData(59); xorBitMap(15)(57) := currentData(57); xorBitMap(15)(56) := currentData(56); xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(160) := previousCrc(0); xorBitMap(15)(164) := previousCrc(4); xorBitMap(15)(165) := previousCrc(5); xorBitMap(15)(168) := previousCrc(8); xorBitMap(15)(169) := previousCrc(9); xorBitMap(15)(170) := previousCrc(10); xorBitMap(15)(174) := previousCrc(14); xorBitMap(15)(175) := previousCrc(15); xorBitMap(15)(177) := previousCrc(17); xorBitMap(15)(179) := previousCrc(19); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(181) := previousCrc(21); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(185) := previousCrc(25); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(191) := previousCrc(31); 
      xorBitMap(16)(111) := currentData(111); xorBitMap(16)(110) := currentData(110); xorBitMap(16)(109) := currentData(109); xorBitMap(16)(105) := currentData(105); xorBitMap(16)(104) := currentData(104); xorBitMap(16)(103) := currentData(103); xorBitMap(16)(102) := currentData(102); xorBitMap(16)(100) := currentData(100); xorBitMap(16)(99) := currentData(99); xorBitMap(16)(97) := currentData(97); xorBitMap(16)(94) := currentData(94); xorBitMap(16)(91) := currentData(91); xorBitMap(16)(90) := currentData(90); xorBitMap(16)(89) := currentData(89); xorBitMap(16)(87) := currentData(87); xorBitMap(16)(86) := currentData(86); xorBitMap(16)(84) := currentData(84); xorBitMap(16)(83) := currentData(83); xorBitMap(16)(82) := currentData(82); xorBitMap(16)(78) := currentData(78); xorBitMap(16)(77) := currentData(77); xorBitMap(16)(75) := currentData(75); xorBitMap(16)(68) := currentData(68); xorBitMap(16)(66) := currentData(66); xorBitMap(16)(57) := currentData(57); xorBitMap(16)(56) := currentData(56); xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(162) := previousCrc(2); xorBitMap(16)(163) := previousCrc(3); xorBitMap(16)(164) := previousCrc(4); xorBitMap(16)(166) := previousCrc(6); xorBitMap(16)(167) := previousCrc(7); xorBitMap(16)(169) := previousCrc(9); xorBitMap(16)(170) := previousCrc(10); xorBitMap(16)(171) := previousCrc(11); xorBitMap(16)(174) := previousCrc(14); xorBitMap(16)(177) := previousCrc(17); xorBitMap(16)(179) := previousCrc(19); xorBitMap(16)(180) := previousCrc(20); xorBitMap(16)(182) := previousCrc(22); xorBitMap(16)(183) := previousCrc(23); xorBitMap(16)(184) := previousCrc(24); xorBitMap(16)(185) := previousCrc(25); xorBitMap(16)(189) := previousCrc(29); xorBitMap(16)(190) := previousCrc(30); xorBitMap(16)(191) := previousCrc(31); 
      xorBitMap(17)(111) := currentData(111); xorBitMap(17)(110) := currentData(110); xorBitMap(17)(106) := currentData(106); xorBitMap(17)(105) := currentData(105); xorBitMap(17)(104) := currentData(104); xorBitMap(17)(103) := currentData(103); xorBitMap(17)(101) := currentData(101); xorBitMap(17)(100) := currentData(100); xorBitMap(17)(98) := currentData(98); xorBitMap(17)(95) := currentData(95); xorBitMap(17)(92) := currentData(92); xorBitMap(17)(91) := currentData(91); xorBitMap(17)(90) := currentData(90); xorBitMap(17)(88) := currentData(88); xorBitMap(17)(87) := currentData(87); xorBitMap(17)(85) := currentData(85); xorBitMap(17)(84) := currentData(84); xorBitMap(17)(83) := currentData(83); xorBitMap(17)(79) := currentData(79); xorBitMap(17)(78) := currentData(78); xorBitMap(17)(76) := currentData(76); xorBitMap(17)(69) := currentData(69); xorBitMap(17)(67) := currentData(67); xorBitMap(17)(58) := currentData(58); xorBitMap(17)(57) := currentData(57); xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(163) := previousCrc(3); xorBitMap(17)(164) := previousCrc(4); xorBitMap(17)(165) := previousCrc(5); xorBitMap(17)(167) := previousCrc(7); xorBitMap(17)(168) := previousCrc(8); xorBitMap(17)(170) := previousCrc(10); xorBitMap(17)(171) := previousCrc(11); xorBitMap(17)(172) := previousCrc(12); xorBitMap(17)(175) := previousCrc(15); xorBitMap(17)(178) := previousCrc(18); xorBitMap(17)(180) := previousCrc(20); xorBitMap(17)(181) := previousCrc(21); xorBitMap(17)(183) := previousCrc(23); xorBitMap(17)(184) := previousCrc(24); xorBitMap(17)(185) := previousCrc(25); xorBitMap(17)(186) := previousCrc(26); xorBitMap(17)(190) := previousCrc(30); xorBitMap(17)(191) := previousCrc(31); 
      xorBitMap(18)(111) := currentData(111); xorBitMap(18)(107) := currentData(107); xorBitMap(18)(106) := currentData(106); xorBitMap(18)(105) := currentData(105); xorBitMap(18)(104) := currentData(104); xorBitMap(18)(102) := currentData(102); xorBitMap(18)(101) := currentData(101); xorBitMap(18)(99) := currentData(99); xorBitMap(18)(96) := currentData(96); xorBitMap(18)(93) := currentData(93); xorBitMap(18)(92) := currentData(92); xorBitMap(18)(91) := currentData(91); xorBitMap(18)(89) := currentData(89); xorBitMap(18)(88) := currentData(88); xorBitMap(18)(86) := currentData(86); xorBitMap(18)(85) := currentData(85); xorBitMap(18)(84) := currentData(84); xorBitMap(18)(80) := currentData(80); xorBitMap(18)(79) := currentData(79); xorBitMap(18)(77) := currentData(77); xorBitMap(18)(70) := currentData(70); xorBitMap(18)(68) := currentData(68); xorBitMap(18)(59) := currentData(59); xorBitMap(18)(58) := currentData(58); xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(160) := previousCrc(0); xorBitMap(18)(164) := previousCrc(4); xorBitMap(18)(165) := previousCrc(5); xorBitMap(18)(166) := previousCrc(6); xorBitMap(18)(168) := previousCrc(8); xorBitMap(18)(169) := previousCrc(9); xorBitMap(18)(171) := previousCrc(11); xorBitMap(18)(172) := previousCrc(12); xorBitMap(18)(173) := previousCrc(13); xorBitMap(18)(176) := previousCrc(16); xorBitMap(18)(179) := previousCrc(19); xorBitMap(18)(181) := previousCrc(21); xorBitMap(18)(182) := previousCrc(22); xorBitMap(18)(184) := previousCrc(24); xorBitMap(18)(185) := previousCrc(25); xorBitMap(18)(186) := previousCrc(26); xorBitMap(18)(187) := previousCrc(27); xorBitMap(18)(191) := previousCrc(31); 
      xorBitMap(19)(108) := currentData(108); xorBitMap(19)(107) := currentData(107); xorBitMap(19)(106) := currentData(106); xorBitMap(19)(105) := currentData(105); xorBitMap(19)(103) := currentData(103); xorBitMap(19)(102) := currentData(102); xorBitMap(19)(100) := currentData(100); xorBitMap(19)(97) := currentData(97); xorBitMap(19)(94) := currentData(94); xorBitMap(19)(93) := currentData(93); xorBitMap(19)(92) := currentData(92); xorBitMap(19)(90) := currentData(90); xorBitMap(19)(89) := currentData(89); xorBitMap(19)(87) := currentData(87); xorBitMap(19)(86) := currentData(86); xorBitMap(19)(85) := currentData(85); xorBitMap(19)(81) := currentData(81); xorBitMap(19)(80) := currentData(80); xorBitMap(19)(78) := currentData(78); xorBitMap(19)(71) := currentData(71); xorBitMap(19)(69) := currentData(69); xorBitMap(19)(60) := currentData(60); xorBitMap(19)(59) := currentData(59); xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(160) := previousCrc(0); xorBitMap(19)(161) := previousCrc(1); xorBitMap(19)(165) := previousCrc(5); xorBitMap(19)(166) := previousCrc(6); xorBitMap(19)(167) := previousCrc(7); xorBitMap(19)(169) := previousCrc(9); xorBitMap(19)(170) := previousCrc(10); xorBitMap(19)(172) := previousCrc(12); xorBitMap(19)(173) := previousCrc(13); xorBitMap(19)(174) := previousCrc(14); xorBitMap(19)(177) := previousCrc(17); xorBitMap(19)(180) := previousCrc(20); xorBitMap(19)(182) := previousCrc(22); xorBitMap(19)(183) := previousCrc(23); xorBitMap(19)(185) := previousCrc(25); xorBitMap(19)(186) := previousCrc(26); xorBitMap(19)(187) := previousCrc(27); xorBitMap(19)(188) := previousCrc(28); 
      xorBitMap(20)(109) := currentData(109); xorBitMap(20)(108) := currentData(108); xorBitMap(20)(107) := currentData(107); xorBitMap(20)(106) := currentData(106); xorBitMap(20)(104) := currentData(104); xorBitMap(20)(103) := currentData(103); xorBitMap(20)(101) := currentData(101); xorBitMap(20)(98) := currentData(98); xorBitMap(20)(95) := currentData(95); xorBitMap(20)(94) := currentData(94); xorBitMap(20)(93) := currentData(93); xorBitMap(20)(91) := currentData(91); xorBitMap(20)(90) := currentData(90); xorBitMap(20)(88) := currentData(88); xorBitMap(20)(87) := currentData(87); xorBitMap(20)(86) := currentData(86); xorBitMap(20)(82) := currentData(82); xorBitMap(20)(81) := currentData(81); xorBitMap(20)(79) := currentData(79); xorBitMap(20)(72) := currentData(72); xorBitMap(20)(70) := currentData(70); xorBitMap(20)(61) := currentData(61); xorBitMap(20)(60) := currentData(60); xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(161) := previousCrc(1); xorBitMap(20)(162) := previousCrc(2); xorBitMap(20)(166) := previousCrc(6); xorBitMap(20)(167) := previousCrc(7); xorBitMap(20)(168) := previousCrc(8); xorBitMap(20)(170) := previousCrc(10); xorBitMap(20)(171) := previousCrc(11); xorBitMap(20)(173) := previousCrc(13); xorBitMap(20)(174) := previousCrc(14); xorBitMap(20)(175) := previousCrc(15); xorBitMap(20)(178) := previousCrc(18); xorBitMap(20)(181) := previousCrc(21); xorBitMap(20)(183) := previousCrc(23); xorBitMap(20)(184) := previousCrc(24); xorBitMap(20)(186) := previousCrc(26); xorBitMap(20)(187) := previousCrc(27); xorBitMap(20)(188) := previousCrc(28); xorBitMap(20)(189) := previousCrc(29); 
      xorBitMap(21)(110) := currentData(110); xorBitMap(21)(109) := currentData(109); xorBitMap(21)(108) := currentData(108); xorBitMap(21)(107) := currentData(107); xorBitMap(21)(105) := currentData(105); xorBitMap(21)(104) := currentData(104); xorBitMap(21)(102) := currentData(102); xorBitMap(21)(99) := currentData(99); xorBitMap(21)(96) := currentData(96); xorBitMap(21)(95) := currentData(95); xorBitMap(21)(94) := currentData(94); xorBitMap(21)(92) := currentData(92); xorBitMap(21)(91) := currentData(91); xorBitMap(21)(89) := currentData(89); xorBitMap(21)(88) := currentData(88); xorBitMap(21)(87) := currentData(87); xorBitMap(21)(83) := currentData(83); xorBitMap(21)(82) := currentData(82); xorBitMap(21)(80) := currentData(80); xorBitMap(21)(73) := currentData(73); xorBitMap(21)(71) := currentData(71); xorBitMap(21)(62) := currentData(62); xorBitMap(21)(61) := currentData(61); xorBitMap(21)(56) := currentData(56); xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(160) := previousCrc(0); xorBitMap(21)(162) := previousCrc(2); xorBitMap(21)(163) := previousCrc(3); xorBitMap(21)(167) := previousCrc(7); xorBitMap(21)(168) := previousCrc(8); xorBitMap(21)(169) := previousCrc(9); xorBitMap(21)(171) := previousCrc(11); xorBitMap(21)(172) := previousCrc(12); xorBitMap(21)(174) := previousCrc(14); xorBitMap(21)(175) := previousCrc(15); xorBitMap(21)(176) := previousCrc(16); xorBitMap(21)(179) := previousCrc(19); xorBitMap(21)(182) := previousCrc(22); xorBitMap(21)(184) := previousCrc(24); xorBitMap(21)(185) := previousCrc(25); xorBitMap(21)(187) := previousCrc(27); xorBitMap(21)(188) := previousCrc(28); xorBitMap(21)(189) := previousCrc(29); xorBitMap(21)(190) := previousCrc(30); 
      xorBitMap(22)(109) := currentData(109); xorBitMap(22)(108) := currentData(108); xorBitMap(22)(105) := currentData(105); xorBitMap(22)(104) := currentData(104); xorBitMap(22)(101) := currentData(101); xorBitMap(22)(100) := currentData(100); xorBitMap(22)(99) := currentData(99); xorBitMap(22)(98) := currentData(98); xorBitMap(22)(94) := currentData(94); xorBitMap(22)(93) := currentData(93); xorBitMap(22)(92) := currentData(92); xorBitMap(22)(90) := currentData(90); xorBitMap(22)(89) := currentData(89); xorBitMap(22)(88) := currentData(88); xorBitMap(22)(87) := currentData(87); xorBitMap(22)(85) := currentData(85); xorBitMap(22)(82) := currentData(82); xorBitMap(22)(79) := currentData(79); xorBitMap(22)(74) := currentData(74); xorBitMap(22)(73) := currentData(73); xorBitMap(22)(68) := currentData(68); xorBitMap(22)(67) := currentData(67); xorBitMap(22)(66) := currentData(66); xorBitMap(22)(65) := currentData(65); xorBitMap(22)(62) := currentData(62); xorBitMap(22)(61) := currentData(61); xorBitMap(22)(60) := currentData(60); xorBitMap(22)(58) := currentData(58); xorBitMap(22)(57) := currentData(57); xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(162) := previousCrc(2); xorBitMap(22)(165) := previousCrc(5); xorBitMap(22)(167) := previousCrc(7); xorBitMap(22)(168) := previousCrc(8); xorBitMap(22)(169) := previousCrc(9); xorBitMap(22)(170) := previousCrc(10); xorBitMap(22)(172) := previousCrc(12); xorBitMap(22)(173) := previousCrc(13); xorBitMap(22)(174) := previousCrc(14); xorBitMap(22)(178) := previousCrc(18); xorBitMap(22)(179) := previousCrc(19); xorBitMap(22)(180) := previousCrc(20); xorBitMap(22)(181) := previousCrc(21); xorBitMap(22)(184) := previousCrc(24); xorBitMap(22)(185) := previousCrc(25); xorBitMap(22)(188) := previousCrc(28); xorBitMap(22)(189) := previousCrc(29); 
      xorBitMap(23)(111) := currentData(111); xorBitMap(23)(109) := currentData(109); xorBitMap(23)(105) := currentData(105); xorBitMap(23)(104) := currentData(104); xorBitMap(23)(103) := currentData(103); xorBitMap(23)(102) := currentData(102); xorBitMap(23)(100) := currentData(100); xorBitMap(23)(98) := currentData(98); xorBitMap(23)(97) := currentData(97); xorBitMap(23)(96) := currentData(96); xorBitMap(23)(93) := currentData(93); xorBitMap(23)(91) := currentData(91); xorBitMap(23)(90) := currentData(90); xorBitMap(23)(89) := currentData(89); xorBitMap(23)(88) := currentData(88); xorBitMap(23)(87) := currentData(87); xorBitMap(23)(86) := currentData(86); xorBitMap(23)(85) := currentData(85); xorBitMap(23)(84) := currentData(84); xorBitMap(23)(82) := currentData(82); xorBitMap(23)(81) := currentData(81); xorBitMap(23)(80) := currentData(80); xorBitMap(23)(79) := currentData(79); xorBitMap(23)(75) := currentData(75); xorBitMap(23)(74) := currentData(74); xorBitMap(23)(73) := currentData(73); xorBitMap(23)(72) := currentData(72); xorBitMap(23)(69) := currentData(69); xorBitMap(23)(65) := currentData(65); xorBitMap(23)(62) := currentData(62); xorBitMap(23)(60) := currentData(60); xorBitMap(23)(59) := currentData(59); xorBitMap(23)(56) := currentData(56); xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(160) := previousCrc(0); xorBitMap(23)(161) := previousCrc(1); xorBitMap(23)(162) := previousCrc(2); xorBitMap(23)(164) := previousCrc(4); xorBitMap(23)(165) := previousCrc(5); xorBitMap(23)(166) := previousCrc(6); xorBitMap(23)(167) := previousCrc(7); xorBitMap(23)(168) := previousCrc(8); xorBitMap(23)(169) := previousCrc(9); xorBitMap(23)(170) := previousCrc(10); xorBitMap(23)(171) := previousCrc(11); xorBitMap(23)(173) := previousCrc(13); xorBitMap(23)(176) := previousCrc(16); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(178) := previousCrc(18); xorBitMap(23)(180) := previousCrc(20); xorBitMap(23)(182) := previousCrc(22); xorBitMap(23)(183) := previousCrc(23); xorBitMap(23)(184) := previousCrc(24); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(189) := previousCrc(29); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(110) := currentData(110); xorBitMap(24)(106) := currentData(106); xorBitMap(24)(105) := currentData(105); xorBitMap(24)(104) := currentData(104); xorBitMap(24)(103) := currentData(103); xorBitMap(24)(101) := currentData(101); xorBitMap(24)(99) := currentData(99); xorBitMap(24)(98) := currentData(98); xorBitMap(24)(97) := currentData(97); xorBitMap(24)(94) := currentData(94); xorBitMap(24)(92) := currentData(92); xorBitMap(24)(91) := currentData(91); xorBitMap(24)(90) := currentData(90); xorBitMap(24)(89) := currentData(89); xorBitMap(24)(88) := currentData(88); xorBitMap(24)(87) := currentData(87); xorBitMap(24)(86) := currentData(86); xorBitMap(24)(85) := currentData(85); xorBitMap(24)(83) := currentData(83); xorBitMap(24)(82) := currentData(82); xorBitMap(24)(81) := currentData(81); xorBitMap(24)(80) := currentData(80); xorBitMap(24)(76) := currentData(76); xorBitMap(24)(75) := currentData(75); xorBitMap(24)(74) := currentData(74); xorBitMap(24)(73) := currentData(73); xorBitMap(24)(70) := currentData(70); xorBitMap(24)(66) := currentData(66); xorBitMap(24)(63) := currentData(63); xorBitMap(24)(61) := currentData(61); xorBitMap(24)(60) := currentData(60); xorBitMap(24)(57) := currentData(57); xorBitMap(24)(56) := currentData(56); xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(160) := previousCrc(0); xorBitMap(24)(161) := previousCrc(1); xorBitMap(24)(162) := previousCrc(2); xorBitMap(24)(163) := previousCrc(3); xorBitMap(24)(165) := previousCrc(5); xorBitMap(24)(166) := previousCrc(6); xorBitMap(24)(167) := previousCrc(7); xorBitMap(24)(168) := previousCrc(8); xorBitMap(24)(169) := previousCrc(9); xorBitMap(24)(170) := previousCrc(10); xorBitMap(24)(171) := previousCrc(11); xorBitMap(24)(172) := previousCrc(12); xorBitMap(24)(174) := previousCrc(14); xorBitMap(24)(177) := previousCrc(17); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(179) := previousCrc(19); xorBitMap(24)(181) := previousCrc(21); xorBitMap(24)(183) := previousCrc(23); xorBitMap(24)(184) := previousCrc(24); xorBitMap(24)(185) := previousCrc(25); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(190) := previousCrc(30); 
      xorBitMap(25)(111) := currentData(111); xorBitMap(25)(107) := currentData(107); xorBitMap(25)(106) := currentData(106); xorBitMap(25)(105) := currentData(105); xorBitMap(25)(104) := currentData(104); xorBitMap(25)(102) := currentData(102); xorBitMap(25)(100) := currentData(100); xorBitMap(25)(99) := currentData(99); xorBitMap(25)(98) := currentData(98); xorBitMap(25)(95) := currentData(95); xorBitMap(25)(93) := currentData(93); xorBitMap(25)(92) := currentData(92); xorBitMap(25)(91) := currentData(91); xorBitMap(25)(90) := currentData(90); xorBitMap(25)(89) := currentData(89); xorBitMap(25)(88) := currentData(88); xorBitMap(25)(87) := currentData(87); xorBitMap(25)(86) := currentData(86); xorBitMap(25)(84) := currentData(84); xorBitMap(25)(83) := currentData(83); xorBitMap(25)(82) := currentData(82); xorBitMap(25)(81) := currentData(81); xorBitMap(25)(77) := currentData(77); xorBitMap(25)(76) := currentData(76); xorBitMap(25)(75) := currentData(75); xorBitMap(25)(74) := currentData(74); xorBitMap(25)(71) := currentData(71); xorBitMap(25)(67) := currentData(67); xorBitMap(25)(64) := currentData(64); xorBitMap(25)(62) := currentData(62); xorBitMap(25)(61) := currentData(61); xorBitMap(25)(58) := currentData(58); xorBitMap(25)(57) := currentData(57); xorBitMap(25)(56) := currentData(56); xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(161) := previousCrc(1); xorBitMap(25)(162) := previousCrc(2); xorBitMap(25)(163) := previousCrc(3); xorBitMap(25)(164) := previousCrc(4); xorBitMap(25)(166) := previousCrc(6); xorBitMap(25)(167) := previousCrc(7); xorBitMap(25)(168) := previousCrc(8); xorBitMap(25)(169) := previousCrc(9); xorBitMap(25)(170) := previousCrc(10); xorBitMap(25)(171) := previousCrc(11); xorBitMap(25)(172) := previousCrc(12); xorBitMap(25)(173) := previousCrc(13); xorBitMap(25)(175) := previousCrc(15); xorBitMap(25)(178) := previousCrc(18); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(180) := previousCrc(20); xorBitMap(25)(182) := previousCrc(22); xorBitMap(25)(184) := previousCrc(24); xorBitMap(25)(185) := previousCrc(25); xorBitMap(25)(186) := previousCrc(26); xorBitMap(25)(187) := previousCrc(27); xorBitMap(25)(191) := previousCrc(31); 
      xorBitMap(26)(111) := currentData(111); xorBitMap(26)(110) := currentData(110); xorBitMap(26)(108) := currentData(108); xorBitMap(26)(107) := currentData(107); xorBitMap(26)(105) := currentData(105); xorBitMap(26)(104) := currentData(104); xorBitMap(26)(100) := currentData(100); xorBitMap(26)(98) := currentData(98); xorBitMap(26)(97) := currentData(97); xorBitMap(26)(95) := currentData(95); xorBitMap(26)(93) := currentData(93); xorBitMap(26)(92) := currentData(92); xorBitMap(26)(91) := currentData(91); xorBitMap(26)(90) := currentData(90); xorBitMap(26)(89) := currentData(89); xorBitMap(26)(88) := currentData(88); xorBitMap(26)(81) := currentData(81); xorBitMap(26)(79) := currentData(79); xorBitMap(26)(78) := currentData(78); xorBitMap(26)(77) := currentData(77); xorBitMap(26)(76) := currentData(76); xorBitMap(26)(75) := currentData(75); xorBitMap(26)(73) := currentData(73); xorBitMap(26)(67) := currentData(67); xorBitMap(26)(66) := currentData(66); xorBitMap(26)(62) := currentData(62); xorBitMap(26)(61) := currentData(61); xorBitMap(26)(60) := currentData(60); xorBitMap(26)(59) := currentData(59); xorBitMap(26)(57) := currentData(57); xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(161) := previousCrc(1); xorBitMap(26)(168) := previousCrc(8); xorBitMap(26)(169) := previousCrc(9); xorBitMap(26)(170) := previousCrc(10); xorBitMap(26)(171) := previousCrc(11); xorBitMap(26)(172) := previousCrc(12); xorBitMap(26)(173) := previousCrc(13); xorBitMap(26)(175) := previousCrc(15); xorBitMap(26)(177) := previousCrc(17); xorBitMap(26)(178) := previousCrc(18); xorBitMap(26)(180) := previousCrc(20); xorBitMap(26)(184) := previousCrc(24); xorBitMap(26)(185) := previousCrc(25); xorBitMap(26)(187) := previousCrc(27); xorBitMap(26)(188) := previousCrc(28); xorBitMap(26)(190) := previousCrc(30); xorBitMap(26)(191) := previousCrc(31); 
      xorBitMap(27)(111) := currentData(111); xorBitMap(27)(109) := currentData(109); xorBitMap(27)(108) := currentData(108); xorBitMap(27)(106) := currentData(106); xorBitMap(27)(105) := currentData(105); xorBitMap(27)(101) := currentData(101); xorBitMap(27)(99) := currentData(99); xorBitMap(27)(98) := currentData(98); xorBitMap(27)(96) := currentData(96); xorBitMap(27)(94) := currentData(94); xorBitMap(27)(93) := currentData(93); xorBitMap(27)(92) := currentData(92); xorBitMap(27)(91) := currentData(91); xorBitMap(27)(90) := currentData(90); xorBitMap(27)(89) := currentData(89); xorBitMap(27)(82) := currentData(82); xorBitMap(27)(80) := currentData(80); xorBitMap(27)(79) := currentData(79); xorBitMap(27)(78) := currentData(78); xorBitMap(27)(77) := currentData(77); xorBitMap(27)(76) := currentData(76); xorBitMap(27)(74) := currentData(74); xorBitMap(27)(68) := currentData(68); xorBitMap(27)(67) := currentData(67); xorBitMap(27)(63) := currentData(63); xorBitMap(27)(62) := currentData(62); xorBitMap(27)(61) := currentData(61); xorBitMap(27)(60) := currentData(60); xorBitMap(27)(58) := currentData(58); xorBitMap(27)(56) := currentData(56); xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(160) := previousCrc(0); xorBitMap(27)(162) := previousCrc(2); xorBitMap(27)(169) := previousCrc(9); xorBitMap(27)(170) := previousCrc(10); xorBitMap(27)(171) := previousCrc(11); xorBitMap(27)(172) := previousCrc(12); xorBitMap(27)(173) := previousCrc(13); xorBitMap(27)(174) := previousCrc(14); xorBitMap(27)(176) := previousCrc(16); xorBitMap(27)(178) := previousCrc(18); xorBitMap(27)(179) := previousCrc(19); xorBitMap(27)(181) := previousCrc(21); xorBitMap(27)(185) := previousCrc(25); xorBitMap(27)(186) := previousCrc(26); xorBitMap(27)(188) := previousCrc(28); xorBitMap(27)(189) := previousCrc(29); xorBitMap(27)(191) := previousCrc(31); 
      xorBitMap(28)(110) := currentData(110); xorBitMap(28)(109) := currentData(109); xorBitMap(28)(107) := currentData(107); xorBitMap(28)(106) := currentData(106); xorBitMap(28)(102) := currentData(102); xorBitMap(28)(100) := currentData(100); xorBitMap(28)(99) := currentData(99); xorBitMap(28)(97) := currentData(97); xorBitMap(28)(95) := currentData(95); xorBitMap(28)(94) := currentData(94); xorBitMap(28)(93) := currentData(93); xorBitMap(28)(92) := currentData(92); xorBitMap(28)(91) := currentData(91); xorBitMap(28)(90) := currentData(90); xorBitMap(28)(83) := currentData(83); xorBitMap(28)(81) := currentData(81); xorBitMap(28)(80) := currentData(80); xorBitMap(28)(79) := currentData(79); xorBitMap(28)(78) := currentData(78); xorBitMap(28)(77) := currentData(77); xorBitMap(28)(75) := currentData(75); xorBitMap(28)(69) := currentData(69); xorBitMap(28)(68) := currentData(68); xorBitMap(28)(64) := currentData(64); xorBitMap(28)(63) := currentData(63); xorBitMap(28)(62) := currentData(62); xorBitMap(28)(61) := currentData(61); xorBitMap(28)(59) := currentData(59); xorBitMap(28)(57) := currentData(57); xorBitMap(28)(56) := currentData(56); xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(160) := previousCrc(0); xorBitMap(28)(161) := previousCrc(1); xorBitMap(28)(163) := previousCrc(3); xorBitMap(28)(170) := previousCrc(10); xorBitMap(28)(171) := previousCrc(11); xorBitMap(28)(172) := previousCrc(12); xorBitMap(28)(173) := previousCrc(13); xorBitMap(28)(174) := previousCrc(14); xorBitMap(28)(175) := previousCrc(15); xorBitMap(28)(177) := previousCrc(17); xorBitMap(28)(179) := previousCrc(19); xorBitMap(28)(180) := previousCrc(20); xorBitMap(28)(182) := previousCrc(22); xorBitMap(28)(186) := previousCrc(26); xorBitMap(28)(187) := previousCrc(27); xorBitMap(28)(189) := previousCrc(29); xorBitMap(28)(190) := previousCrc(30); 
      xorBitMap(29)(111) := currentData(111); xorBitMap(29)(110) := currentData(110); xorBitMap(29)(108) := currentData(108); xorBitMap(29)(107) := currentData(107); xorBitMap(29)(103) := currentData(103); xorBitMap(29)(101) := currentData(101); xorBitMap(29)(100) := currentData(100); xorBitMap(29)(98) := currentData(98); xorBitMap(29)(96) := currentData(96); xorBitMap(29)(95) := currentData(95); xorBitMap(29)(94) := currentData(94); xorBitMap(29)(93) := currentData(93); xorBitMap(29)(92) := currentData(92); xorBitMap(29)(91) := currentData(91); xorBitMap(29)(84) := currentData(84); xorBitMap(29)(82) := currentData(82); xorBitMap(29)(81) := currentData(81); xorBitMap(29)(80) := currentData(80); xorBitMap(29)(79) := currentData(79); xorBitMap(29)(78) := currentData(78); xorBitMap(29)(76) := currentData(76); xorBitMap(29)(70) := currentData(70); xorBitMap(29)(69) := currentData(69); xorBitMap(29)(65) := currentData(65); xorBitMap(29)(64) := currentData(64); xorBitMap(29)(63) := currentData(63); xorBitMap(29)(62) := currentData(62); xorBitMap(29)(60) := currentData(60); xorBitMap(29)(58) := currentData(58); xorBitMap(29)(57) := currentData(57); xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(160) := previousCrc(0); xorBitMap(29)(161) := previousCrc(1); xorBitMap(29)(162) := previousCrc(2); xorBitMap(29)(164) := previousCrc(4); xorBitMap(29)(171) := previousCrc(11); xorBitMap(29)(172) := previousCrc(12); xorBitMap(29)(173) := previousCrc(13); xorBitMap(29)(174) := previousCrc(14); xorBitMap(29)(175) := previousCrc(15); xorBitMap(29)(176) := previousCrc(16); xorBitMap(29)(178) := previousCrc(18); xorBitMap(29)(180) := previousCrc(20); xorBitMap(29)(181) := previousCrc(21); xorBitMap(29)(183) := previousCrc(23); xorBitMap(29)(187) := previousCrc(27); xorBitMap(29)(188) := previousCrc(28); xorBitMap(29)(190) := previousCrc(30); xorBitMap(29)(191) := previousCrc(31); 
      xorBitMap(30)(111) := currentData(111); xorBitMap(30)(109) := currentData(109); xorBitMap(30)(108) := currentData(108); xorBitMap(30)(104) := currentData(104); xorBitMap(30)(102) := currentData(102); xorBitMap(30)(101) := currentData(101); xorBitMap(30)(99) := currentData(99); xorBitMap(30)(97) := currentData(97); xorBitMap(30)(96) := currentData(96); xorBitMap(30)(95) := currentData(95); xorBitMap(30)(94) := currentData(94); xorBitMap(30)(93) := currentData(93); xorBitMap(30)(92) := currentData(92); xorBitMap(30)(85) := currentData(85); xorBitMap(30)(83) := currentData(83); xorBitMap(30)(82) := currentData(82); xorBitMap(30)(81) := currentData(81); xorBitMap(30)(80) := currentData(80); xorBitMap(30)(79) := currentData(79); xorBitMap(30)(77) := currentData(77); xorBitMap(30)(71) := currentData(71); xorBitMap(30)(70) := currentData(70); xorBitMap(30)(66) := currentData(66); xorBitMap(30)(65) := currentData(65); xorBitMap(30)(64) := currentData(64); xorBitMap(30)(63) := currentData(63); xorBitMap(30)(61) := currentData(61); xorBitMap(30)(59) := currentData(59); xorBitMap(30)(58) := currentData(58); xorBitMap(30)(56) := currentData(56); xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(160) := previousCrc(0); xorBitMap(30)(161) := previousCrc(1); xorBitMap(30)(162) := previousCrc(2); xorBitMap(30)(163) := previousCrc(3); xorBitMap(30)(165) := previousCrc(5); xorBitMap(30)(172) := previousCrc(12); xorBitMap(30)(173) := previousCrc(13); xorBitMap(30)(174) := previousCrc(14); xorBitMap(30)(175) := previousCrc(15); xorBitMap(30)(176) := previousCrc(16); xorBitMap(30)(177) := previousCrc(17); xorBitMap(30)(179) := previousCrc(19); xorBitMap(30)(181) := previousCrc(21); xorBitMap(30)(182) := previousCrc(22); xorBitMap(30)(184) := previousCrc(24); xorBitMap(30)(188) := previousCrc(28); xorBitMap(30)(189) := previousCrc(29); xorBitMap(30)(191) := previousCrc(31); 
      xorBitMap(31)(110) := currentData(110); xorBitMap(31)(109) := currentData(109); xorBitMap(31)(105) := currentData(105); xorBitMap(31)(103) := currentData(103); xorBitMap(31)(102) := currentData(102); xorBitMap(31)(100) := currentData(100); xorBitMap(31)(98) := currentData(98); xorBitMap(31)(97) := currentData(97); xorBitMap(31)(96) := currentData(96); xorBitMap(31)(95) := currentData(95); xorBitMap(31)(94) := currentData(94); xorBitMap(31)(93) := currentData(93); xorBitMap(31)(86) := currentData(86); xorBitMap(31)(84) := currentData(84); xorBitMap(31)(83) := currentData(83); xorBitMap(31)(82) := currentData(82); xorBitMap(31)(81) := currentData(81); xorBitMap(31)(80) := currentData(80); xorBitMap(31)(78) := currentData(78); xorBitMap(31)(72) := currentData(72); xorBitMap(31)(71) := currentData(71); xorBitMap(31)(67) := currentData(67); xorBitMap(31)(66) := currentData(66); xorBitMap(31)(65) := currentData(65); xorBitMap(31)(64) := currentData(64); xorBitMap(31)(62) := currentData(62); xorBitMap(31)(60) := currentData(60); xorBitMap(31)(59) := currentData(59); xorBitMap(31)(57) := currentData(57); xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(160) := previousCrc(0); xorBitMap(31)(161) := previousCrc(1); xorBitMap(31)(162) := previousCrc(2); xorBitMap(31)(163) := previousCrc(3); xorBitMap(31)(164) := previousCrc(4); xorBitMap(31)(166) := previousCrc(6); xorBitMap(31)(173) := previousCrc(13); xorBitMap(31)(174) := previousCrc(14); xorBitMap(31)(175) := previousCrc(15); xorBitMap(31)(176) := previousCrc(16); xorBitMap(31)(177) := previousCrc(17); xorBitMap(31)(178) := previousCrc(18); xorBitMap(31)(180) := previousCrc(20); xorBitMap(31)(182) := previousCrc(22); xorBitMap(31)(183) := previousCrc(23); xorBitMap(31)(185) := previousCrc(25); xorBitMap(31)(189) := previousCrc(29); xorBitMap(31)(190) := previousCrc(30); 
   end procedure;

   procedure xorBitMap15Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(119 downto 0)) is 
   begin
      xorBitMap(0)(119) := currentData(119); xorBitMap(0)(118) := currentData(118); xorBitMap(0)(117) := currentData(117); xorBitMap(0)(116) := currentData(116); xorBitMap(0)(114) := currentData(114); xorBitMap(0)(113) := currentData(113); xorBitMap(0)(111) := currentData(111); xorBitMap(0)(110) := currentData(110); xorBitMap(0)(106) := currentData(106); xorBitMap(0)(104) := currentData(104); xorBitMap(0)(103) := currentData(103); xorBitMap(0)(101) := currentData(101); xorBitMap(0)(99) := currentData(99); xorBitMap(0)(98) := currentData(98); xorBitMap(0)(97) := currentData(97); xorBitMap(0)(96) := currentData(96); xorBitMap(0)(95) := currentData(95); xorBitMap(0)(94) := currentData(94); xorBitMap(0)(87) := currentData(87); xorBitMap(0)(85) := currentData(85); xorBitMap(0)(84) := currentData(84); xorBitMap(0)(83) := currentData(83); xorBitMap(0)(82) := currentData(82); xorBitMap(0)(81) := currentData(81); xorBitMap(0)(79) := currentData(79); xorBitMap(0)(73) := currentData(73); xorBitMap(0)(72) := currentData(72); xorBitMap(0)(68) := currentData(68); xorBitMap(0)(67) := currentData(67); xorBitMap(0)(66) := currentData(66); xorBitMap(0)(65) := currentData(65); xorBitMap(0)(63) := currentData(63); xorBitMap(0)(61) := currentData(61); xorBitMap(0)(60) := currentData(60); xorBitMap(0)(58) := currentData(58); xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(166) := previousCrc(6); xorBitMap(0)(167) := previousCrc(7); xorBitMap(0)(168) := previousCrc(8); xorBitMap(0)(169) := previousCrc(9); xorBitMap(0)(170) := previousCrc(10); xorBitMap(0)(171) := previousCrc(11); xorBitMap(0)(173) := previousCrc(13); xorBitMap(0)(175) := previousCrc(15); xorBitMap(0)(176) := previousCrc(16); xorBitMap(0)(178) := previousCrc(18); xorBitMap(0)(182) := previousCrc(22); xorBitMap(0)(183) := previousCrc(23); xorBitMap(0)(185) := previousCrc(25); xorBitMap(0)(186) := previousCrc(26); xorBitMap(0)(188) := previousCrc(28); xorBitMap(0)(189) := previousCrc(29); xorBitMap(0)(190) := previousCrc(30); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(116) := currentData(116); xorBitMap(1)(115) := currentData(115); xorBitMap(1)(113) := currentData(113); xorBitMap(1)(112) := currentData(112); xorBitMap(1)(110) := currentData(110); xorBitMap(1)(107) := currentData(107); xorBitMap(1)(106) := currentData(106); xorBitMap(1)(105) := currentData(105); xorBitMap(1)(103) := currentData(103); xorBitMap(1)(102) := currentData(102); xorBitMap(1)(101) := currentData(101); xorBitMap(1)(100) := currentData(100); xorBitMap(1)(94) := currentData(94); xorBitMap(1)(88) := currentData(88); xorBitMap(1)(87) := currentData(87); xorBitMap(1)(86) := currentData(86); xorBitMap(1)(81) := currentData(81); xorBitMap(1)(80) := currentData(80); xorBitMap(1)(79) := currentData(79); xorBitMap(1)(74) := currentData(74); xorBitMap(1)(72) := currentData(72); xorBitMap(1)(69) := currentData(69); xorBitMap(1)(65) := currentData(65); xorBitMap(1)(64) := currentData(64); xorBitMap(1)(63) := currentData(63); xorBitMap(1)(62) := currentData(62); xorBitMap(1)(60) := currentData(60); xorBitMap(1)(59) := currentData(59); xorBitMap(1)(58) := currentData(58); xorBitMap(1)(56) := currentData(56); xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(160) := previousCrc(0); xorBitMap(1)(166) := previousCrc(6); xorBitMap(1)(172) := previousCrc(12); xorBitMap(1)(173) := previousCrc(13); xorBitMap(1)(174) := previousCrc(14); xorBitMap(1)(175) := previousCrc(15); xorBitMap(1)(177) := previousCrc(17); xorBitMap(1)(178) := previousCrc(18); xorBitMap(1)(179) := previousCrc(19); xorBitMap(1)(182) := previousCrc(22); xorBitMap(1)(184) := previousCrc(24); xorBitMap(1)(185) := previousCrc(25); xorBitMap(1)(187) := previousCrc(27); xorBitMap(1)(188) := previousCrc(28); 
      xorBitMap(2)(119) := currentData(119); xorBitMap(2)(118) := currentData(118); xorBitMap(2)(110) := currentData(110); xorBitMap(2)(108) := currentData(108); xorBitMap(2)(107) := currentData(107); xorBitMap(2)(102) := currentData(102); xorBitMap(2)(99) := currentData(99); xorBitMap(2)(98) := currentData(98); xorBitMap(2)(97) := currentData(97); xorBitMap(2)(96) := currentData(96); xorBitMap(2)(94) := currentData(94); xorBitMap(2)(89) := currentData(89); xorBitMap(2)(88) := currentData(88); xorBitMap(2)(85) := currentData(85); xorBitMap(2)(84) := currentData(84); xorBitMap(2)(83) := currentData(83); xorBitMap(2)(80) := currentData(80); xorBitMap(2)(79) := currentData(79); xorBitMap(2)(75) := currentData(75); xorBitMap(2)(72) := currentData(72); xorBitMap(2)(70) := currentData(70); xorBitMap(2)(68) := currentData(68); xorBitMap(2)(67) := currentData(67); xorBitMap(2)(64) := currentData(64); xorBitMap(2)(59) := currentData(59); xorBitMap(2)(58) := currentData(58); xorBitMap(2)(57) := currentData(57); xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(160) := previousCrc(0); xorBitMap(2)(161) := previousCrc(1); xorBitMap(2)(166) := previousCrc(6); xorBitMap(2)(168) := previousCrc(8); xorBitMap(2)(169) := previousCrc(9); xorBitMap(2)(170) := previousCrc(10); xorBitMap(2)(171) := previousCrc(11); xorBitMap(2)(174) := previousCrc(14); xorBitMap(2)(179) := previousCrc(19); xorBitMap(2)(180) := previousCrc(20); xorBitMap(2)(182) := previousCrc(22); xorBitMap(2)(190) := previousCrc(30); xorBitMap(2)(191) := previousCrc(31); 
      xorBitMap(3)(119) := currentData(119); xorBitMap(3)(111) := currentData(111); xorBitMap(3)(109) := currentData(109); xorBitMap(3)(108) := currentData(108); xorBitMap(3)(103) := currentData(103); xorBitMap(3)(100) := currentData(100); xorBitMap(3)(99) := currentData(99); xorBitMap(3)(98) := currentData(98); xorBitMap(3)(97) := currentData(97); xorBitMap(3)(95) := currentData(95); xorBitMap(3)(90) := currentData(90); xorBitMap(3)(89) := currentData(89); xorBitMap(3)(86) := currentData(86); xorBitMap(3)(85) := currentData(85); xorBitMap(3)(84) := currentData(84); xorBitMap(3)(81) := currentData(81); xorBitMap(3)(80) := currentData(80); xorBitMap(3)(76) := currentData(76); xorBitMap(3)(73) := currentData(73); xorBitMap(3)(71) := currentData(71); xorBitMap(3)(69) := currentData(69); xorBitMap(3)(68) := currentData(68); xorBitMap(3)(65) := currentData(65); xorBitMap(3)(60) := currentData(60); xorBitMap(3)(59) := currentData(59); xorBitMap(3)(58) := currentData(58); xorBitMap(3)(56) := currentData(56); xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(161) := previousCrc(1); xorBitMap(3)(162) := previousCrc(2); xorBitMap(3)(167) := previousCrc(7); xorBitMap(3)(169) := previousCrc(9); xorBitMap(3)(170) := previousCrc(10); xorBitMap(3)(171) := previousCrc(11); xorBitMap(3)(172) := previousCrc(12); xorBitMap(3)(175) := previousCrc(15); xorBitMap(3)(180) := previousCrc(20); xorBitMap(3)(181) := previousCrc(21); xorBitMap(3)(183) := previousCrc(23); xorBitMap(3)(191) := previousCrc(31); 
      xorBitMap(4)(119) := currentData(119); xorBitMap(4)(118) := currentData(118); xorBitMap(4)(117) := currentData(117); xorBitMap(4)(116) := currentData(116); xorBitMap(4)(114) := currentData(114); xorBitMap(4)(113) := currentData(113); xorBitMap(4)(112) := currentData(112); xorBitMap(4)(111) := currentData(111); xorBitMap(4)(109) := currentData(109); xorBitMap(4)(106) := currentData(106); xorBitMap(4)(103) := currentData(103); xorBitMap(4)(100) := currentData(100); xorBitMap(4)(97) := currentData(97); xorBitMap(4)(95) := currentData(95); xorBitMap(4)(94) := currentData(94); xorBitMap(4)(91) := currentData(91); xorBitMap(4)(90) := currentData(90); xorBitMap(4)(86) := currentData(86); xorBitMap(4)(84) := currentData(84); xorBitMap(4)(83) := currentData(83); xorBitMap(4)(79) := currentData(79); xorBitMap(4)(77) := currentData(77); xorBitMap(4)(74) := currentData(74); xorBitMap(4)(73) := currentData(73); xorBitMap(4)(70) := currentData(70); xorBitMap(4)(69) := currentData(69); xorBitMap(4)(68) := currentData(68); xorBitMap(4)(67) := currentData(67); xorBitMap(4)(65) := currentData(65); xorBitMap(4)(63) := currentData(63); xorBitMap(4)(59) := currentData(59); xorBitMap(4)(58) := currentData(58); xorBitMap(4)(57) := currentData(57); xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(162) := previousCrc(2); xorBitMap(4)(163) := previousCrc(3); xorBitMap(4)(166) := previousCrc(6); xorBitMap(4)(167) := previousCrc(7); xorBitMap(4)(169) := previousCrc(9); xorBitMap(4)(172) := previousCrc(12); xorBitMap(4)(175) := previousCrc(15); xorBitMap(4)(178) := previousCrc(18); xorBitMap(4)(181) := previousCrc(21); xorBitMap(4)(183) := previousCrc(23); xorBitMap(4)(184) := previousCrc(24); xorBitMap(4)(185) := previousCrc(25); xorBitMap(4)(186) := previousCrc(26); xorBitMap(4)(188) := previousCrc(28); xorBitMap(4)(189) := previousCrc(29); xorBitMap(4)(190) := previousCrc(30); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(116) := currentData(116); xorBitMap(5)(115) := currentData(115); xorBitMap(5)(112) := currentData(112); xorBitMap(5)(111) := currentData(111); xorBitMap(5)(107) := currentData(107); xorBitMap(5)(106) := currentData(106); xorBitMap(5)(103) := currentData(103); xorBitMap(5)(99) := currentData(99); xorBitMap(5)(97) := currentData(97); xorBitMap(5)(94) := currentData(94); xorBitMap(5)(92) := currentData(92); xorBitMap(5)(91) := currentData(91); xorBitMap(5)(83) := currentData(83); xorBitMap(5)(82) := currentData(82); xorBitMap(5)(81) := currentData(81); xorBitMap(5)(80) := currentData(80); xorBitMap(5)(79) := currentData(79); xorBitMap(5)(78) := currentData(78); xorBitMap(5)(75) := currentData(75); xorBitMap(5)(74) := currentData(74); xorBitMap(5)(73) := currentData(73); xorBitMap(5)(72) := currentData(72); xorBitMap(5)(71) := currentData(71); xorBitMap(5)(70) := currentData(70); xorBitMap(5)(69) := currentData(69); xorBitMap(5)(67) := currentData(67); xorBitMap(5)(65) := currentData(65); xorBitMap(5)(64) := currentData(64); xorBitMap(5)(63) := currentData(63); xorBitMap(5)(61) := currentData(61); xorBitMap(5)(59) := currentData(59); xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(163) := previousCrc(3); xorBitMap(5)(164) := previousCrc(4); xorBitMap(5)(166) := previousCrc(6); xorBitMap(5)(169) := previousCrc(9); xorBitMap(5)(171) := previousCrc(11); xorBitMap(5)(175) := previousCrc(15); xorBitMap(5)(178) := previousCrc(18); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(183) := previousCrc(23); xorBitMap(5)(184) := previousCrc(24); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(188) := previousCrc(28); 
      xorBitMap(6)(117) := currentData(117); xorBitMap(6)(116) := currentData(116); xorBitMap(6)(113) := currentData(113); xorBitMap(6)(112) := currentData(112); xorBitMap(6)(108) := currentData(108); xorBitMap(6)(107) := currentData(107); xorBitMap(6)(104) := currentData(104); xorBitMap(6)(100) := currentData(100); xorBitMap(6)(98) := currentData(98); xorBitMap(6)(95) := currentData(95); xorBitMap(6)(93) := currentData(93); xorBitMap(6)(92) := currentData(92); xorBitMap(6)(84) := currentData(84); xorBitMap(6)(83) := currentData(83); xorBitMap(6)(82) := currentData(82); xorBitMap(6)(81) := currentData(81); xorBitMap(6)(80) := currentData(80); xorBitMap(6)(79) := currentData(79); xorBitMap(6)(76) := currentData(76); xorBitMap(6)(75) := currentData(75); xorBitMap(6)(74) := currentData(74); xorBitMap(6)(73) := currentData(73); xorBitMap(6)(72) := currentData(72); xorBitMap(6)(71) := currentData(71); xorBitMap(6)(70) := currentData(70); xorBitMap(6)(68) := currentData(68); xorBitMap(6)(66) := currentData(66); xorBitMap(6)(65) := currentData(65); xorBitMap(6)(64) := currentData(64); xorBitMap(6)(62) := currentData(62); xorBitMap(6)(60) := currentData(60); xorBitMap(6)(56) := currentData(56); xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(164) := previousCrc(4); xorBitMap(6)(165) := previousCrc(5); xorBitMap(6)(167) := previousCrc(7); xorBitMap(6)(170) := previousCrc(10); xorBitMap(6)(172) := previousCrc(12); xorBitMap(6)(176) := previousCrc(16); xorBitMap(6)(179) := previousCrc(19); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(184) := previousCrc(24); xorBitMap(6)(185) := previousCrc(25); xorBitMap(6)(188) := previousCrc(28); xorBitMap(6)(189) := previousCrc(29); 
      xorBitMap(7)(119) := currentData(119); xorBitMap(7)(116) := currentData(116); xorBitMap(7)(111) := currentData(111); xorBitMap(7)(110) := currentData(110); xorBitMap(7)(109) := currentData(109); xorBitMap(7)(108) := currentData(108); xorBitMap(7)(106) := currentData(106); xorBitMap(7)(105) := currentData(105); xorBitMap(7)(104) := currentData(104); xorBitMap(7)(103) := currentData(103); xorBitMap(7)(98) := currentData(98); xorBitMap(7)(97) := currentData(97); xorBitMap(7)(95) := currentData(95); xorBitMap(7)(93) := currentData(93); xorBitMap(7)(87) := currentData(87); xorBitMap(7)(80) := currentData(80); xorBitMap(7)(79) := currentData(79); xorBitMap(7)(77) := currentData(77); xorBitMap(7)(76) := currentData(76); xorBitMap(7)(75) := currentData(75); xorBitMap(7)(74) := currentData(74); xorBitMap(7)(71) := currentData(71); xorBitMap(7)(69) := currentData(69); xorBitMap(7)(68) := currentData(68); xorBitMap(7)(60) := currentData(60); xorBitMap(7)(58) := currentData(58); xorBitMap(7)(57) := currentData(57); xorBitMap(7)(56) := currentData(56); xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(165) := previousCrc(5); xorBitMap(7)(167) := previousCrc(7); xorBitMap(7)(169) := previousCrc(9); xorBitMap(7)(170) := previousCrc(10); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(176) := previousCrc(16); xorBitMap(7)(177) := previousCrc(17); xorBitMap(7)(178) := previousCrc(18); xorBitMap(7)(180) := previousCrc(20); xorBitMap(7)(181) := previousCrc(21); xorBitMap(7)(182) := previousCrc(22); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(188) := previousCrc(28); xorBitMap(7)(191) := previousCrc(31); 
      xorBitMap(8)(119) := currentData(119); xorBitMap(8)(118) := currentData(118); xorBitMap(8)(116) := currentData(116); xorBitMap(8)(114) := currentData(114); xorBitMap(8)(113) := currentData(113); xorBitMap(8)(112) := currentData(112); xorBitMap(8)(109) := currentData(109); xorBitMap(8)(107) := currentData(107); xorBitMap(8)(105) := currentData(105); xorBitMap(8)(103) := currentData(103); xorBitMap(8)(101) := currentData(101); xorBitMap(8)(97) := currentData(97); xorBitMap(8)(95) := currentData(95); xorBitMap(8)(88) := currentData(88); xorBitMap(8)(87) := currentData(87); xorBitMap(8)(85) := currentData(85); xorBitMap(8)(84) := currentData(84); xorBitMap(8)(83) := currentData(83); xorBitMap(8)(82) := currentData(82); xorBitMap(8)(80) := currentData(80); xorBitMap(8)(79) := currentData(79); xorBitMap(8)(78) := currentData(78); xorBitMap(8)(77) := currentData(77); xorBitMap(8)(76) := currentData(76); xorBitMap(8)(75) := currentData(75); xorBitMap(8)(73) := currentData(73); xorBitMap(8)(70) := currentData(70); xorBitMap(8)(69) := currentData(69); xorBitMap(8)(68) := currentData(68); xorBitMap(8)(67) := currentData(67); xorBitMap(8)(66) := currentData(66); xorBitMap(8)(65) := currentData(65); xorBitMap(8)(63) := currentData(63); xorBitMap(8)(60) := currentData(60); xorBitMap(8)(59) := currentData(59); xorBitMap(8)(57) := currentData(57); xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(160) := previousCrc(0); xorBitMap(8)(167) := previousCrc(7); xorBitMap(8)(169) := previousCrc(9); xorBitMap(8)(173) := previousCrc(13); xorBitMap(8)(175) := previousCrc(15); xorBitMap(8)(177) := previousCrc(17); xorBitMap(8)(179) := previousCrc(19); xorBitMap(8)(181) := previousCrc(21); xorBitMap(8)(184) := previousCrc(24); xorBitMap(8)(185) := previousCrc(25); xorBitMap(8)(186) := previousCrc(26); xorBitMap(8)(188) := previousCrc(28); xorBitMap(8)(190) := previousCrc(30); xorBitMap(8)(191) := previousCrc(31); 
      xorBitMap(9)(119) := currentData(119); xorBitMap(9)(117) := currentData(117); xorBitMap(9)(115) := currentData(115); xorBitMap(9)(114) := currentData(114); xorBitMap(9)(113) := currentData(113); xorBitMap(9)(110) := currentData(110); xorBitMap(9)(108) := currentData(108); xorBitMap(9)(106) := currentData(106); xorBitMap(9)(104) := currentData(104); xorBitMap(9)(102) := currentData(102); xorBitMap(9)(98) := currentData(98); xorBitMap(9)(96) := currentData(96); xorBitMap(9)(89) := currentData(89); xorBitMap(9)(88) := currentData(88); xorBitMap(9)(86) := currentData(86); xorBitMap(9)(85) := currentData(85); xorBitMap(9)(84) := currentData(84); xorBitMap(9)(83) := currentData(83); xorBitMap(9)(81) := currentData(81); xorBitMap(9)(80) := currentData(80); xorBitMap(9)(79) := currentData(79); xorBitMap(9)(78) := currentData(78); xorBitMap(9)(77) := currentData(77); xorBitMap(9)(76) := currentData(76); xorBitMap(9)(74) := currentData(74); xorBitMap(9)(71) := currentData(71); xorBitMap(9)(70) := currentData(70); xorBitMap(9)(69) := currentData(69); xorBitMap(9)(68) := currentData(68); xorBitMap(9)(67) := currentData(67); xorBitMap(9)(66) := currentData(66); xorBitMap(9)(64) := currentData(64); xorBitMap(9)(61) := currentData(61); xorBitMap(9)(60) := currentData(60); xorBitMap(9)(58) := currentData(58); xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(160) := previousCrc(0); xorBitMap(9)(161) := previousCrc(1); xorBitMap(9)(168) := previousCrc(8); xorBitMap(9)(170) := previousCrc(10); xorBitMap(9)(174) := previousCrc(14); xorBitMap(9)(176) := previousCrc(16); xorBitMap(9)(178) := previousCrc(18); xorBitMap(9)(180) := previousCrc(20); xorBitMap(9)(182) := previousCrc(22); xorBitMap(9)(185) := previousCrc(25); xorBitMap(9)(186) := previousCrc(26); xorBitMap(9)(187) := previousCrc(27); xorBitMap(9)(189) := previousCrc(29); xorBitMap(9)(191) := previousCrc(31); 
      xorBitMap(10)(119) := currentData(119); xorBitMap(10)(117) := currentData(117); xorBitMap(10)(115) := currentData(115); xorBitMap(10)(113) := currentData(113); xorBitMap(10)(110) := currentData(110); xorBitMap(10)(109) := currentData(109); xorBitMap(10)(107) := currentData(107); xorBitMap(10)(106) := currentData(106); xorBitMap(10)(105) := currentData(105); xorBitMap(10)(104) := currentData(104); xorBitMap(10)(101) := currentData(101); xorBitMap(10)(98) := currentData(98); xorBitMap(10)(96) := currentData(96); xorBitMap(10)(95) := currentData(95); xorBitMap(10)(94) := currentData(94); xorBitMap(10)(90) := currentData(90); xorBitMap(10)(89) := currentData(89); xorBitMap(10)(86) := currentData(86); xorBitMap(10)(83) := currentData(83); xorBitMap(10)(80) := currentData(80); xorBitMap(10)(78) := currentData(78); xorBitMap(10)(77) := currentData(77); xorBitMap(10)(75) := currentData(75); xorBitMap(10)(73) := currentData(73); xorBitMap(10)(71) := currentData(71); xorBitMap(10)(70) := currentData(70); xorBitMap(10)(69) := currentData(69); xorBitMap(10)(66) := currentData(66); xorBitMap(10)(63) := currentData(63); xorBitMap(10)(62) := currentData(62); xorBitMap(10)(60) := currentData(60); xorBitMap(10)(59) := currentData(59); xorBitMap(10)(58) := currentData(58); xorBitMap(10)(56) := currentData(56); xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(161) := previousCrc(1); xorBitMap(10)(162) := previousCrc(2); xorBitMap(10)(166) := previousCrc(6); xorBitMap(10)(167) := previousCrc(7); xorBitMap(10)(168) := previousCrc(8); xorBitMap(10)(170) := previousCrc(10); xorBitMap(10)(173) := previousCrc(13); xorBitMap(10)(176) := previousCrc(16); xorBitMap(10)(177) := previousCrc(17); xorBitMap(10)(178) := previousCrc(18); xorBitMap(10)(179) := previousCrc(19); xorBitMap(10)(181) := previousCrc(21); xorBitMap(10)(182) := previousCrc(22); xorBitMap(10)(185) := previousCrc(25); xorBitMap(10)(187) := previousCrc(27); xorBitMap(10)(189) := previousCrc(29); xorBitMap(10)(191) := previousCrc(31); 
      xorBitMap(11)(119) := currentData(119); xorBitMap(11)(117) := currentData(117); xorBitMap(11)(113) := currentData(113); xorBitMap(11)(108) := currentData(108); xorBitMap(11)(107) := currentData(107); xorBitMap(11)(105) := currentData(105); xorBitMap(11)(104) := currentData(104); xorBitMap(11)(103) := currentData(103); xorBitMap(11)(102) := currentData(102); xorBitMap(11)(101) := currentData(101); xorBitMap(11)(98) := currentData(98); xorBitMap(11)(94) := currentData(94); xorBitMap(11)(91) := currentData(91); xorBitMap(11)(90) := currentData(90); xorBitMap(11)(85) := currentData(85); xorBitMap(11)(83) := currentData(83); xorBitMap(11)(82) := currentData(82); xorBitMap(11)(78) := currentData(78); xorBitMap(11)(76) := currentData(76); xorBitMap(11)(74) := currentData(74); xorBitMap(11)(73) := currentData(73); xorBitMap(11)(71) := currentData(71); xorBitMap(11)(70) := currentData(70); xorBitMap(11)(68) := currentData(68); xorBitMap(11)(66) := currentData(66); xorBitMap(11)(65) := currentData(65); xorBitMap(11)(64) := currentData(64); xorBitMap(11)(59) := currentData(59); xorBitMap(11)(58) := currentData(58); xorBitMap(11)(57) := currentData(57); xorBitMap(11)(56) := currentData(56); xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(162) := previousCrc(2); xorBitMap(11)(163) := previousCrc(3); xorBitMap(11)(166) := previousCrc(6); xorBitMap(11)(170) := previousCrc(10); xorBitMap(11)(173) := previousCrc(13); xorBitMap(11)(174) := previousCrc(14); xorBitMap(11)(175) := previousCrc(15); xorBitMap(11)(176) := previousCrc(16); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(179) := previousCrc(19); xorBitMap(11)(180) := previousCrc(20); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(189) := previousCrc(29); xorBitMap(11)(191) := previousCrc(31); 
      xorBitMap(12)(119) := currentData(119); xorBitMap(12)(117) := currentData(117); xorBitMap(12)(116) := currentData(116); xorBitMap(12)(113) := currentData(113); xorBitMap(12)(111) := currentData(111); xorBitMap(12)(110) := currentData(110); xorBitMap(12)(109) := currentData(109); xorBitMap(12)(108) := currentData(108); xorBitMap(12)(105) := currentData(105); xorBitMap(12)(102) := currentData(102); xorBitMap(12)(101) := currentData(101); xorBitMap(12)(98) := currentData(98); xorBitMap(12)(97) := currentData(97); xorBitMap(12)(96) := currentData(96); xorBitMap(12)(94) := currentData(94); xorBitMap(12)(92) := currentData(92); xorBitMap(12)(91) := currentData(91); xorBitMap(12)(87) := currentData(87); xorBitMap(12)(86) := currentData(86); xorBitMap(12)(85) := currentData(85); xorBitMap(12)(82) := currentData(82); xorBitMap(12)(81) := currentData(81); xorBitMap(12)(77) := currentData(77); xorBitMap(12)(75) := currentData(75); xorBitMap(12)(74) := currentData(74); xorBitMap(12)(73) := currentData(73); xorBitMap(12)(71) := currentData(71); xorBitMap(12)(69) := currentData(69); xorBitMap(12)(68) := currentData(68); xorBitMap(12)(63) := currentData(63); xorBitMap(12)(61) := currentData(61); xorBitMap(12)(59) := currentData(59); xorBitMap(12)(57) := currentData(57); xorBitMap(12)(56) := currentData(56); xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(163) := previousCrc(3); xorBitMap(12)(164) := previousCrc(4); xorBitMap(12)(166) := previousCrc(6); xorBitMap(12)(168) := previousCrc(8); xorBitMap(12)(169) := previousCrc(9); xorBitMap(12)(170) := previousCrc(10); xorBitMap(12)(173) := previousCrc(13); xorBitMap(12)(174) := previousCrc(14); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(180) := previousCrc(20); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(182) := previousCrc(22); xorBitMap(12)(183) := previousCrc(23); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(188) := previousCrc(28); xorBitMap(12)(189) := previousCrc(29); xorBitMap(12)(191) := previousCrc(31); 
      xorBitMap(13)(118) := currentData(118); xorBitMap(13)(117) := currentData(117); xorBitMap(13)(114) := currentData(114); xorBitMap(13)(112) := currentData(112); xorBitMap(13)(111) := currentData(111); xorBitMap(13)(110) := currentData(110); xorBitMap(13)(109) := currentData(109); xorBitMap(13)(106) := currentData(106); xorBitMap(13)(103) := currentData(103); xorBitMap(13)(102) := currentData(102); xorBitMap(13)(99) := currentData(99); xorBitMap(13)(98) := currentData(98); xorBitMap(13)(97) := currentData(97); xorBitMap(13)(95) := currentData(95); xorBitMap(13)(93) := currentData(93); xorBitMap(13)(92) := currentData(92); xorBitMap(13)(88) := currentData(88); xorBitMap(13)(87) := currentData(87); xorBitMap(13)(86) := currentData(86); xorBitMap(13)(83) := currentData(83); xorBitMap(13)(82) := currentData(82); xorBitMap(13)(78) := currentData(78); xorBitMap(13)(76) := currentData(76); xorBitMap(13)(75) := currentData(75); xorBitMap(13)(74) := currentData(74); xorBitMap(13)(72) := currentData(72); xorBitMap(13)(70) := currentData(70); xorBitMap(13)(69) := currentData(69); xorBitMap(13)(64) := currentData(64); xorBitMap(13)(62) := currentData(62); xorBitMap(13)(60) := currentData(60); xorBitMap(13)(58) := currentData(58); xorBitMap(13)(57) := currentData(57); xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(160) := previousCrc(0); xorBitMap(13)(164) := previousCrc(4); xorBitMap(13)(165) := previousCrc(5); xorBitMap(13)(167) := previousCrc(7); xorBitMap(13)(169) := previousCrc(9); xorBitMap(13)(170) := previousCrc(10); xorBitMap(13)(171) := previousCrc(11); xorBitMap(13)(174) := previousCrc(14); xorBitMap(13)(175) := previousCrc(15); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(181) := previousCrc(21); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(183) := previousCrc(23); xorBitMap(13)(184) := previousCrc(24); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(189) := previousCrc(29); xorBitMap(13)(190) := previousCrc(30); 
      xorBitMap(14)(119) := currentData(119); xorBitMap(14)(118) := currentData(118); xorBitMap(14)(115) := currentData(115); xorBitMap(14)(113) := currentData(113); xorBitMap(14)(112) := currentData(112); xorBitMap(14)(111) := currentData(111); xorBitMap(14)(110) := currentData(110); xorBitMap(14)(107) := currentData(107); xorBitMap(14)(104) := currentData(104); xorBitMap(14)(103) := currentData(103); xorBitMap(14)(100) := currentData(100); xorBitMap(14)(99) := currentData(99); xorBitMap(14)(98) := currentData(98); xorBitMap(14)(96) := currentData(96); xorBitMap(14)(94) := currentData(94); xorBitMap(14)(93) := currentData(93); xorBitMap(14)(89) := currentData(89); xorBitMap(14)(88) := currentData(88); xorBitMap(14)(87) := currentData(87); xorBitMap(14)(84) := currentData(84); xorBitMap(14)(83) := currentData(83); xorBitMap(14)(79) := currentData(79); xorBitMap(14)(77) := currentData(77); xorBitMap(14)(76) := currentData(76); xorBitMap(14)(75) := currentData(75); xorBitMap(14)(73) := currentData(73); xorBitMap(14)(71) := currentData(71); xorBitMap(14)(70) := currentData(70); xorBitMap(14)(65) := currentData(65); xorBitMap(14)(63) := currentData(63); xorBitMap(14)(61) := currentData(61); xorBitMap(14)(59) := currentData(59); xorBitMap(14)(58) := currentData(58); xorBitMap(14)(56) := currentData(56); xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(160) := previousCrc(0); xorBitMap(14)(161) := previousCrc(1); xorBitMap(14)(165) := previousCrc(5); xorBitMap(14)(166) := previousCrc(6); xorBitMap(14)(168) := previousCrc(8); xorBitMap(14)(170) := previousCrc(10); xorBitMap(14)(171) := previousCrc(11); xorBitMap(14)(172) := previousCrc(12); xorBitMap(14)(175) := previousCrc(15); xorBitMap(14)(176) := previousCrc(16); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(182) := previousCrc(22); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(184) := previousCrc(24); xorBitMap(14)(185) := previousCrc(25); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(190) := previousCrc(30); xorBitMap(14)(191) := previousCrc(31); 
      xorBitMap(15)(119) := currentData(119); xorBitMap(15)(116) := currentData(116); xorBitMap(15)(114) := currentData(114); xorBitMap(15)(113) := currentData(113); xorBitMap(15)(112) := currentData(112); xorBitMap(15)(111) := currentData(111); xorBitMap(15)(108) := currentData(108); xorBitMap(15)(105) := currentData(105); xorBitMap(15)(104) := currentData(104); xorBitMap(15)(101) := currentData(101); xorBitMap(15)(100) := currentData(100); xorBitMap(15)(99) := currentData(99); xorBitMap(15)(97) := currentData(97); xorBitMap(15)(95) := currentData(95); xorBitMap(15)(94) := currentData(94); xorBitMap(15)(90) := currentData(90); xorBitMap(15)(89) := currentData(89); xorBitMap(15)(88) := currentData(88); xorBitMap(15)(85) := currentData(85); xorBitMap(15)(84) := currentData(84); xorBitMap(15)(80) := currentData(80); xorBitMap(15)(78) := currentData(78); xorBitMap(15)(77) := currentData(77); xorBitMap(15)(76) := currentData(76); xorBitMap(15)(74) := currentData(74); xorBitMap(15)(72) := currentData(72); xorBitMap(15)(71) := currentData(71); xorBitMap(15)(66) := currentData(66); xorBitMap(15)(64) := currentData(64); xorBitMap(15)(62) := currentData(62); xorBitMap(15)(60) := currentData(60); xorBitMap(15)(59) := currentData(59); xorBitMap(15)(57) := currentData(57); xorBitMap(15)(56) := currentData(56); xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(160) := previousCrc(0); xorBitMap(15)(161) := previousCrc(1); xorBitMap(15)(162) := previousCrc(2); xorBitMap(15)(166) := previousCrc(6); xorBitMap(15)(167) := previousCrc(7); xorBitMap(15)(169) := previousCrc(9); xorBitMap(15)(171) := previousCrc(11); xorBitMap(15)(172) := previousCrc(12); xorBitMap(15)(173) := previousCrc(13); xorBitMap(15)(176) := previousCrc(16); xorBitMap(15)(177) := previousCrc(17); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(183) := previousCrc(23); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(185) := previousCrc(25); xorBitMap(15)(186) := previousCrc(26); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(191) := previousCrc(31); 
      xorBitMap(16)(119) := currentData(119); xorBitMap(16)(118) := currentData(118); xorBitMap(16)(116) := currentData(116); xorBitMap(16)(115) := currentData(115); xorBitMap(16)(112) := currentData(112); xorBitMap(16)(111) := currentData(111); xorBitMap(16)(110) := currentData(110); xorBitMap(16)(109) := currentData(109); xorBitMap(16)(105) := currentData(105); xorBitMap(16)(104) := currentData(104); xorBitMap(16)(103) := currentData(103); xorBitMap(16)(102) := currentData(102); xorBitMap(16)(100) := currentData(100); xorBitMap(16)(99) := currentData(99); xorBitMap(16)(97) := currentData(97); xorBitMap(16)(94) := currentData(94); xorBitMap(16)(91) := currentData(91); xorBitMap(16)(90) := currentData(90); xorBitMap(16)(89) := currentData(89); xorBitMap(16)(87) := currentData(87); xorBitMap(16)(86) := currentData(86); xorBitMap(16)(84) := currentData(84); xorBitMap(16)(83) := currentData(83); xorBitMap(16)(82) := currentData(82); xorBitMap(16)(78) := currentData(78); xorBitMap(16)(77) := currentData(77); xorBitMap(16)(75) := currentData(75); xorBitMap(16)(68) := currentData(68); xorBitMap(16)(66) := currentData(66); xorBitMap(16)(57) := currentData(57); xorBitMap(16)(56) := currentData(56); xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(161) := previousCrc(1); xorBitMap(16)(162) := previousCrc(2); xorBitMap(16)(163) := previousCrc(3); xorBitMap(16)(166) := previousCrc(6); xorBitMap(16)(169) := previousCrc(9); xorBitMap(16)(171) := previousCrc(11); xorBitMap(16)(172) := previousCrc(12); xorBitMap(16)(174) := previousCrc(14); xorBitMap(16)(175) := previousCrc(15); xorBitMap(16)(176) := previousCrc(16); xorBitMap(16)(177) := previousCrc(17); xorBitMap(16)(181) := previousCrc(21); xorBitMap(16)(182) := previousCrc(22); xorBitMap(16)(183) := previousCrc(23); xorBitMap(16)(184) := previousCrc(24); xorBitMap(16)(187) := previousCrc(27); xorBitMap(16)(188) := previousCrc(28); xorBitMap(16)(190) := previousCrc(30); xorBitMap(16)(191) := previousCrc(31); 
      xorBitMap(17)(119) := currentData(119); xorBitMap(17)(117) := currentData(117); xorBitMap(17)(116) := currentData(116); xorBitMap(17)(113) := currentData(113); xorBitMap(17)(112) := currentData(112); xorBitMap(17)(111) := currentData(111); xorBitMap(17)(110) := currentData(110); xorBitMap(17)(106) := currentData(106); xorBitMap(17)(105) := currentData(105); xorBitMap(17)(104) := currentData(104); xorBitMap(17)(103) := currentData(103); xorBitMap(17)(101) := currentData(101); xorBitMap(17)(100) := currentData(100); xorBitMap(17)(98) := currentData(98); xorBitMap(17)(95) := currentData(95); xorBitMap(17)(92) := currentData(92); xorBitMap(17)(91) := currentData(91); xorBitMap(17)(90) := currentData(90); xorBitMap(17)(88) := currentData(88); xorBitMap(17)(87) := currentData(87); xorBitMap(17)(85) := currentData(85); xorBitMap(17)(84) := currentData(84); xorBitMap(17)(83) := currentData(83); xorBitMap(17)(79) := currentData(79); xorBitMap(17)(78) := currentData(78); xorBitMap(17)(76) := currentData(76); xorBitMap(17)(69) := currentData(69); xorBitMap(17)(67) := currentData(67); xorBitMap(17)(58) := currentData(58); xorBitMap(17)(57) := currentData(57); xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(160) := previousCrc(0); xorBitMap(17)(162) := previousCrc(2); xorBitMap(17)(163) := previousCrc(3); xorBitMap(17)(164) := previousCrc(4); xorBitMap(17)(167) := previousCrc(7); xorBitMap(17)(170) := previousCrc(10); xorBitMap(17)(172) := previousCrc(12); xorBitMap(17)(173) := previousCrc(13); xorBitMap(17)(175) := previousCrc(15); xorBitMap(17)(176) := previousCrc(16); xorBitMap(17)(177) := previousCrc(17); xorBitMap(17)(178) := previousCrc(18); xorBitMap(17)(182) := previousCrc(22); xorBitMap(17)(183) := previousCrc(23); xorBitMap(17)(184) := previousCrc(24); xorBitMap(17)(185) := previousCrc(25); xorBitMap(17)(188) := previousCrc(28); xorBitMap(17)(189) := previousCrc(29); xorBitMap(17)(191) := previousCrc(31); 
      xorBitMap(18)(118) := currentData(118); xorBitMap(18)(117) := currentData(117); xorBitMap(18)(114) := currentData(114); xorBitMap(18)(113) := currentData(113); xorBitMap(18)(112) := currentData(112); xorBitMap(18)(111) := currentData(111); xorBitMap(18)(107) := currentData(107); xorBitMap(18)(106) := currentData(106); xorBitMap(18)(105) := currentData(105); xorBitMap(18)(104) := currentData(104); xorBitMap(18)(102) := currentData(102); xorBitMap(18)(101) := currentData(101); xorBitMap(18)(99) := currentData(99); xorBitMap(18)(96) := currentData(96); xorBitMap(18)(93) := currentData(93); xorBitMap(18)(92) := currentData(92); xorBitMap(18)(91) := currentData(91); xorBitMap(18)(89) := currentData(89); xorBitMap(18)(88) := currentData(88); xorBitMap(18)(86) := currentData(86); xorBitMap(18)(85) := currentData(85); xorBitMap(18)(84) := currentData(84); xorBitMap(18)(80) := currentData(80); xorBitMap(18)(79) := currentData(79); xorBitMap(18)(77) := currentData(77); xorBitMap(18)(70) := currentData(70); xorBitMap(18)(68) := currentData(68); xorBitMap(18)(59) := currentData(59); xorBitMap(18)(58) := currentData(58); xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(160) := previousCrc(0); xorBitMap(18)(161) := previousCrc(1); xorBitMap(18)(163) := previousCrc(3); xorBitMap(18)(164) := previousCrc(4); xorBitMap(18)(165) := previousCrc(5); xorBitMap(18)(168) := previousCrc(8); xorBitMap(18)(171) := previousCrc(11); xorBitMap(18)(173) := previousCrc(13); xorBitMap(18)(174) := previousCrc(14); xorBitMap(18)(176) := previousCrc(16); xorBitMap(18)(177) := previousCrc(17); xorBitMap(18)(178) := previousCrc(18); xorBitMap(18)(179) := previousCrc(19); xorBitMap(18)(183) := previousCrc(23); xorBitMap(18)(184) := previousCrc(24); xorBitMap(18)(185) := previousCrc(25); xorBitMap(18)(186) := previousCrc(26); xorBitMap(18)(189) := previousCrc(29); xorBitMap(18)(190) := previousCrc(30); 
      xorBitMap(19)(119) := currentData(119); xorBitMap(19)(118) := currentData(118); xorBitMap(19)(115) := currentData(115); xorBitMap(19)(114) := currentData(114); xorBitMap(19)(113) := currentData(113); xorBitMap(19)(112) := currentData(112); xorBitMap(19)(108) := currentData(108); xorBitMap(19)(107) := currentData(107); xorBitMap(19)(106) := currentData(106); xorBitMap(19)(105) := currentData(105); xorBitMap(19)(103) := currentData(103); xorBitMap(19)(102) := currentData(102); xorBitMap(19)(100) := currentData(100); xorBitMap(19)(97) := currentData(97); xorBitMap(19)(94) := currentData(94); xorBitMap(19)(93) := currentData(93); xorBitMap(19)(92) := currentData(92); xorBitMap(19)(90) := currentData(90); xorBitMap(19)(89) := currentData(89); xorBitMap(19)(87) := currentData(87); xorBitMap(19)(86) := currentData(86); xorBitMap(19)(85) := currentData(85); xorBitMap(19)(81) := currentData(81); xorBitMap(19)(80) := currentData(80); xorBitMap(19)(78) := currentData(78); xorBitMap(19)(71) := currentData(71); xorBitMap(19)(69) := currentData(69); xorBitMap(19)(60) := currentData(60); xorBitMap(19)(59) := currentData(59); xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(161) := previousCrc(1); xorBitMap(19)(162) := previousCrc(2); xorBitMap(19)(164) := previousCrc(4); xorBitMap(19)(165) := previousCrc(5); xorBitMap(19)(166) := previousCrc(6); xorBitMap(19)(169) := previousCrc(9); xorBitMap(19)(172) := previousCrc(12); xorBitMap(19)(174) := previousCrc(14); xorBitMap(19)(175) := previousCrc(15); xorBitMap(19)(177) := previousCrc(17); xorBitMap(19)(178) := previousCrc(18); xorBitMap(19)(179) := previousCrc(19); xorBitMap(19)(180) := previousCrc(20); xorBitMap(19)(184) := previousCrc(24); xorBitMap(19)(185) := previousCrc(25); xorBitMap(19)(186) := previousCrc(26); xorBitMap(19)(187) := previousCrc(27); xorBitMap(19)(190) := previousCrc(30); xorBitMap(19)(191) := previousCrc(31); 
      xorBitMap(20)(119) := currentData(119); xorBitMap(20)(116) := currentData(116); xorBitMap(20)(115) := currentData(115); xorBitMap(20)(114) := currentData(114); xorBitMap(20)(113) := currentData(113); xorBitMap(20)(109) := currentData(109); xorBitMap(20)(108) := currentData(108); xorBitMap(20)(107) := currentData(107); xorBitMap(20)(106) := currentData(106); xorBitMap(20)(104) := currentData(104); xorBitMap(20)(103) := currentData(103); xorBitMap(20)(101) := currentData(101); xorBitMap(20)(98) := currentData(98); xorBitMap(20)(95) := currentData(95); xorBitMap(20)(94) := currentData(94); xorBitMap(20)(93) := currentData(93); xorBitMap(20)(91) := currentData(91); xorBitMap(20)(90) := currentData(90); xorBitMap(20)(88) := currentData(88); xorBitMap(20)(87) := currentData(87); xorBitMap(20)(86) := currentData(86); xorBitMap(20)(82) := currentData(82); xorBitMap(20)(81) := currentData(81); xorBitMap(20)(79) := currentData(79); xorBitMap(20)(72) := currentData(72); xorBitMap(20)(70) := currentData(70); xorBitMap(20)(61) := currentData(61); xorBitMap(20)(60) := currentData(60); xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(160) := previousCrc(0); xorBitMap(20)(162) := previousCrc(2); xorBitMap(20)(163) := previousCrc(3); xorBitMap(20)(165) := previousCrc(5); xorBitMap(20)(166) := previousCrc(6); xorBitMap(20)(167) := previousCrc(7); xorBitMap(20)(170) := previousCrc(10); xorBitMap(20)(173) := previousCrc(13); xorBitMap(20)(175) := previousCrc(15); xorBitMap(20)(176) := previousCrc(16); xorBitMap(20)(178) := previousCrc(18); xorBitMap(20)(179) := previousCrc(19); xorBitMap(20)(180) := previousCrc(20); xorBitMap(20)(181) := previousCrc(21); xorBitMap(20)(185) := previousCrc(25); xorBitMap(20)(186) := previousCrc(26); xorBitMap(20)(187) := previousCrc(27); xorBitMap(20)(188) := previousCrc(28); xorBitMap(20)(191) := previousCrc(31); 
      xorBitMap(21)(117) := currentData(117); xorBitMap(21)(116) := currentData(116); xorBitMap(21)(115) := currentData(115); xorBitMap(21)(114) := currentData(114); xorBitMap(21)(110) := currentData(110); xorBitMap(21)(109) := currentData(109); xorBitMap(21)(108) := currentData(108); xorBitMap(21)(107) := currentData(107); xorBitMap(21)(105) := currentData(105); xorBitMap(21)(104) := currentData(104); xorBitMap(21)(102) := currentData(102); xorBitMap(21)(99) := currentData(99); xorBitMap(21)(96) := currentData(96); xorBitMap(21)(95) := currentData(95); xorBitMap(21)(94) := currentData(94); xorBitMap(21)(92) := currentData(92); xorBitMap(21)(91) := currentData(91); xorBitMap(21)(89) := currentData(89); xorBitMap(21)(88) := currentData(88); xorBitMap(21)(87) := currentData(87); xorBitMap(21)(83) := currentData(83); xorBitMap(21)(82) := currentData(82); xorBitMap(21)(80) := currentData(80); xorBitMap(21)(73) := currentData(73); xorBitMap(21)(71) := currentData(71); xorBitMap(21)(62) := currentData(62); xorBitMap(21)(61) := currentData(61); xorBitMap(21)(56) := currentData(56); xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(160) := previousCrc(0); xorBitMap(21)(161) := previousCrc(1); xorBitMap(21)(163) := previousCrc(3); xorBitMap(21)(164) := previousCrc(4); xorBitMap(21)(166) := previousCrc(6); xorBitMap(21)(167) := previousCrc(7); xorBitMap(21)(168) := previousCrc(8); xorBitMap(21)(171) := previousCrc(11); xorBitMap(21)(174) := previousCrc(14); xorBitMap(21)(176) := previousCrc(16); xorBitMap(21)(177) := previousCrc(17); xorBitMap(21)(179) := previousCrc(19); xorBitMap(21)(180) := previousCrc(20); xorBitMap(21)(181) := previousCrc(21); xorBitMap(21)(182) := previousCrc(22); xorBitMap(21)(186) := previousCrc(26); xorBitMap(21)(187) := previousCrc(27); xorBitMap(21)(188) := previousCrc(28); xorBitMap(21)(189) := previousCrc(29); 
      xorBitMap(22)(119) := currentData(119); xorBitMap(22)(115) := currentData(115); xorBitMap(22)(114) := currentData(114); xorBitMap(22)(113) := currentData(113); xorBitMap(22)(109) := currentData(109); xorBitMap(22)(108) := currentData(108); xorBitMap(22)(105) := currentData(105); xorBitMap(22)(104) := currentData(104); xorBitMap(22)(101) := currentData(101); xorBitMap(22)(100) := currentData(100); xorBitMap(22)(99) := currentData(99); xorBitMap(22)(98) := currentData(98); xorBitMap(22)(94) := currentData(94); xorBitMap(22)(93) := currentData(93); xorBitMap(22)(92) := currentData(92); xorBitMap(22)(90) := currentData(90); xorBitMap(22)(89) := currentData(89); xorBitMap(22)(88) := currentData(88); xorBitMap(22)(87) := currentData(87); xorBitMap(22)(85) := currentData(85); xorBitMap(22)(82) := currentData(82); xorBitMap(22)(79) := currentData(79); xorBitMap(22)(74) := currentData(74); xorBitMap(22)(73) := currentData(73); xorBitMap(22)(68) := currentData(68); xorBitMap(22)(67) := currentData(67); xorBitMap(22)(66) := currentData(66); xorBitMap(22)(65) := currentData(65); xorBitMap(22)(62) := currentData(62); xorBitMap(22)(61) := currentData(61); xorBitMap(22)(60) := currentData(60); xorBitMap(22)(58) := currentData(58); xorBitMap(22)(57) := currentData(57); xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(160) := previousCrc(0); xorBitMap(22)(161) := previousCrc(1); xorBitMap(22)(162) := previousCrc(2); xorBitMap(22)(164) := previousCrc(4); xorBitMap(22)(165) := previousCrc(5); xorBitMap(22)(166) := previousCrc(6); xorBitMap(22)(170) := previousCrc(10); xorBitMap(22)(171) := previousCrc(11); xorBitMap(22)(172) := previousCrc(12); xorBitMap(22)(173) := previousCrc(13); xorBitMap(22)(176) := previousCrc(16); xorBitMap(22)(177) := previousCrc(17); xorBitMap(22)(180) := previousCrc(20); xorBitMap(22)(181) := previousCrc(21); xorBitMap(22)(185) := previousCrc(25); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(187) := previousCrc(27); xorBitMap(22)(191) := previousCrc(31); 
      xorBitMap(23)(119) := currentData(119); xorBitMap(23)(118) := currentData(118); xorBitMap(23)(117) := currentData(117); xorBitMap(23)(115) := currentData(115); xorBitMap(23)(113) := currentData(113); xorBitMap(23)(111) := currentData(111); xorBitMap(23)(109) := currentData(109); xorBitMap(23)(105) := currentData(105); xorBitMap(23)(104) := currentData(104); xorBitMap(23)(103) := currentData(103); xorBitMap(23)(102) := currentData(102); xorBitMap(23)(100) := currentData(100); xorBitMap(23)(98) := currentData(98); xorBitMap(23)(97) := currentData(97); xorBitMap(23)(96) := currentData(96); xorBitMap(23)(93) := currentData(93); xorBitMap(23)(91) := currentData(91); xorBitMap(23)(90) := currentData(90); xorBitMap(23)(89) := currentData(89); xorBitMap(23)(88) := currentData(88); xorBitMap(23)(87) := currentData(87); xorBitMap(23)(86) := currentData(86); xorBitMap(23)(85) := currentData(85); xorBitMap(23)(84) := currentData(84); xorBitMap(23)(82) := currentData(82); xorBitMap(23)(81) := currentData(81); xorBitMap(23)(80) := currentData(80); xorBitMap(23)(79) := currentData(79); xorBitMap(23)(75) := currentData(75); xorBitMap(23)(74) := currentData(74); xorBitMap(23)(73) := currentData(73); xorBitMap(23)(72) := currentData(72); xorBitMap(23)(69) := currentData(69); xorBitMap(23)(65) := currentData(65); xorBitMap(23)(62) := currentData(62); xorBitMap(23)(60) := currentData(60); xorBitMap(23)(59) := currentData(59); xorBitMap(23)(56) := currentData(56); xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(160) := previousCrc(0); xorBitMap(23)(161) := previousCrc(1); xorBitMap(23)(162) := previousCrc(2); xorBitMap(23)(163) := previousCrc(3); xorBitMap(23)(165) := previousCrc(5); xorBitMap(23)(168) := previousCrc(8); xorBitMap(23)(169) := previousCrc(9); xorBitMap(23)(170) := previousCrc(10); xorBitMap(23)(172) := previousCrc(12); xorBitMap(23)(174) := previousCrc(14); xorBitMap(23)(175) := previousCrc(15); xorBitMap(23)(176) := previousCrc(16); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(181) := previousCrc(21); xorBitMap(23)(183) := previousCrc(23); xorBitMap(23)(185) := previousCrc(25); xorBitMap(23)(187) := previousCrc(27); xorBitMap(23)(189) := previousCrc(29); xorBitMap(23)(190) := previousCrc(30); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(119) := currentData(119); xorBitMap(24)(118) := currentData(118); xorBitMap(24)(116) := currentData(116); xorBitMap(24)(114) := currentData(114); xorBitMap(24)(112) := currentData(112); xorBitMap(24)(110) := currentData(110); xorBitMap(24)(106) := currentData(106); xorBitMap(24)(105) := currentData(105); xorBitMap(24)(104) := currentData(104); xorBitMap(24)(103) := currentData(103); xorBitMap(24)(101) := currentData(101); xorBitMap(24)(99) := currentData(99); xorBitMap(24)(98) := currentData(98); xorBitMap(24)(97) := currentData(97); xorBitMap(24)(94) := currentData(94); xorBitMap(24)(92) := currentData(92); xorBitMap(24)(91) := currentData(91); xorBitMap(24)(90) := currentData(90); xorBitMap(24)(89) := currentData(89); xorBitMap(24)(88) := currentData(88); xorBitMap(24)(87) := currentData(87); xorBitMap(24)(86) := currentData(86); xorBitMap(24)(85) := currentData(85); xorBitMap(24)(83) := currentData(83); xorBitMap(24)(82) := currentData(82); xorBitMap(24)(81) := currentData(81); xorBitMap(24)(80) := currentData(80); xorBitMap(24)(76) := currentData(76); xorBitMap(24)(75) := currentData(75); xorBitMap(24)(74) := currentData(74); xorBitMap(24)(73) := currentData(73); xorBitMap(24)(70) := currentData(70); xorBitMap(24)(66) := currentData(66); xorBitMap(24)(63) := currentData(63); xorBitMap(24)(61) := currentData(61); xorBitMap(24)(60) := currentData(60); xorBitMap(24)(57) := currentData(57); xorBitMap(24)(56) := currentData(56); xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(160) := previousCrc(0); xorBitMap(24)(161) := previousCrc(1); xorBitMap(24)(162) := previousCrc(2); xorBitMap(24)(163) := previousCrc(3); xorBitMap(24)(164) := previousCrc(4); xorBitMap(24)(166) := previousCrc(6); xorBitMap(24)(169) := previousCrc(9); xorBitMap(24)(170) := previousCrc(10); xorBitMap(24)(171) := previousCrc(11); xorBitMap(24)(173) := previousCrc(13); xorBitMap(24)(175) := previousCrc(15); xorBitMap(24)(176) := previousCrc(16); xorBitMap(24)(177) := previousCrc(17); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(182) := previousCrc(22); xorBitMap(24)(184) := previousCrc(24); xorBitMap(24)(186) := previousCrc(26); xorBitMap(24)(188) := previousCrc(28); xorBitMap(24)(190) := previousCrc(30); xorBitMap(24)(191) := previousCrc(31); 
      xorBitMap(25)(119) := currentData(119); xorBitMap(25)(117) := currentData(117); xorBitMap(25)(115) := currentData(115); xorBitMap(25)(113) := currentData(113); xorBitMap(25)(111) := currentData(111); xorBitMap(25)(107) := currentData(107); xorBitMap(25)(106) := currentData(106); xorBitMap(25)(105) := currentData(105); xorBitMap(25)(104) := currentData(104); xorBitMap(25)(102) := currentData(102); xorBitMap(25)(100) := currentData(100); xorBitMap(25)(99) := currentData(99); xorBitMap(25)(98) := currentData(98); xorBitMap(25)(95) := currentData(95); xorBitMap(25)(93) := currentData(93); xorBitMap(25)(92) := currentData(92); xorBitMap(25)(91) := currentData(91); xorBitMap(25)(90) := currentData(90); xorBitMap(25)(89) := currentData(89); xorBitMap(25)(88) := currentData(88); xorBitMap(25)(87) := currentData(87); xorBitMap(25)(86) := currentData(86); xorBitMap(25)(84) := currentData(84); xorBitMap(25)(83) := currentData(83); xorBitMap(25)(82) := currentData(82); xorBitMap(25)(81) := currentData(81); xorBitMap(25)(77) := currentData(77); xorBitMap(25)(76) := currentData(76); xorBitMap(25)(75) := currentData(75); xorBitMap(25)(74) := currentData(74); xorBitMap(25)(71) := currentData(71); xorBitMap(25)(67) := currentData(67); xorBitMap(25)(64) := currentData(64); xorBitMap(25)(62) := currentData(62); xorBitMap(25)(61) := currentData(61); xorBitMap(25)(58) := currentData(58); xorBitMap(25)(57) := currentData(57); xorBitMap(25)(56) := currentData(56); xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(160) := previousCrc(0); xorBitMap(25)(161) := previousCrc(1); xorBitMap(25)(162) := previousCrc(2); xorBitMap(25)(163) := previousCrc(3); xorBitMap(25)(164) := previousCrc(4); xorBitMap(25)(165) := previousCrc(5); xorBitMap(25)(167) := previousCrc(7); xorBitMap(25)(170) := previousCrc(10); xorBitMap(25)(171) := previousCrc(11); xorBitMap(25)(172) := previousCrc(12); xorBitMap(25)(174) := previousCrc(14); xorBitMap(25)(176) := previousCrc(16); xorBitMap(25)(177) := previousCrc(17); xorBitMap(25)(178) := previousCrc(18); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(183) := previousCrc(23); xorBitMap(25)(185) := previousCrc(25); xorBitMap(25)(187) := previousCrc(27); xorBitMap(25)(189) := previousCrc(29); xorBitMap(25)(191) := previousCrc(31); 
      xorBitMap(26)(119) := currentData(119); xorBitMap(26)(117) := currentData(117); xorBitMap(26)(113) := currentData(113); xorBitMap(26)(112) := currentData(112); xorBitMap(26)(111) := currentData(111); xorBitMap(26)(110) := currentData(110); xorBitMap(26)(108) := currentData(108); xorBitMap(26)(107) := currentData(107); xorBitMap(26)(105) := currentData(105); xorBitMap(26)(104) := currentData(104); xorBitMap(26)(100) := currentData(100); xorBitMap(26)(98) := currentData(98); xorBitMap(26)(97) := currentData(97); xorBitMap(26)(95) := currentData(95); xorBitMap(26)(93) := currentData(93); xorBitMap(26)(92) := currentData(92); xorBitMap(26)(91) := currentData(91); xorBitMap(26)(90) := currentData(90); xorBitMap(26)(89) := currentData(89); xorBitMap(26)(88) := currentData(88); xorBitMap(26)(81) := currentData(81); xorBitMap(26)(79) := currentData(79); xorBitMap(26)(78) := currentData(78); xorBitMap(26)(77) := currentData(77); xorBitMap(26)(76) := currentData(76); xorBitMap(26)(75) := currentData(75); xorBitMap(26)(73) := currentData(73); xorBitMap(26)(67) := currentData(67); xorBitMap(26)(66) := currentData(66); xorBitMap(26)(62) := currentData(62); xorBitMap(26)(61) := currentData(61); xorBitMap(26)(60) := currentData(60); xorBitMap(26)(59) := currentData(59); xorBitMap(26)(57) := currentData(57); xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(160) := previousCrc(0); xorBitMap(26)(161) := previousCrc(1); xorBitMap(26)(162) := previousCrc(2); xorBitMap(26)(163) := previousCrc(3); xorBitMap(26)(164) := previousCrc(4); xorBitMap(26)(165) := previousCrc(5); xorBitMap(26)(167) := previousCrc(7); xorBitMap(26)(169) := previousCrc(9); xorBitMap(26)(170) := previousCrc(10); xorBitMap(26)(172) := previousCrc(12); xorBitMap(26)(176) := previousCrc(16); xorBitMap(26)(177) := previousCrc(17); xorBitMap(26)(179) := previousCrc(19); xorBitMap(26)(180) := previousCrc(20); xorBitMap(26)(182) := previousCrc(22); xorBitMap(26)(183) := previousCrc(23); xorBitMap(26)(184) := previousCrc(24); xorBitMap(26)(185) := previousCrc(25); xorBitMap(26)(189) := previousCrc(29); xorBitMap(26)(191) := previousCrc(31); 
      xorBitMap(27)(118) := currentData(118); xorBitMap(27)(114) := currentData(114); xorBitMap(27)(113) := currentData(113); xorBitMap(27)(112) := currentData(112); xorBitMap(27)(111) := currentData(111); xorBitMap(27)(109) := currentData(109); xorBitMap(27)(108) := currentData(108); xorBitMap(27)(106) := currentData(106); xorBitMap(27)(105) := currentData(105); xorBitMap(27)(101) := currentData(101); xorBitMap(27)(99) := currentData(99); xorBitMap(27)(98) := currentData(98); xorBitMap(27)(96) := currentData(96); xorBitMap(27)(94) := currentData(94); xorBitMap(27)(93) := currentData(93); xorBitMap(27)(92) := currentData(92); xorBitMap(27)(91) := currentData(91); xorBitMap(27)(90) := currentData(90); xorBitMap(27)(89) := currentData(89); xorBitMap(27)(82) := currentData(82); xorBitMap(27)(80) := currentData(80); xorBitMap(27)(79) := currentData(79); xorBitMap(27)(78) := currentData(78); xorBitMap(27)(77) := currentData(77); xorBitMap(27)(76) := currentData(76); xorBitMap(27)(74) := currentData(74); xorBitMap(27)(68) := currentData(68); xorBitMap(27)(67) := currentData(67); xorBitMap(27)(63) := currentData(63); xorBitMap(27)(62) := currentData(62); xorBitMap(27)(61) := currentData(61); xorBitMap(27)(60) := currentData(60); xorBitMap(27)(58) := currentData(58); xorBitMap(27)(56) := currentData(56); xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(161) := previousCrc(1); xorBitMap(27)(162) := previousCrc(2); xorBitMap(27)(163) := previousCrc(3); xorBitMap(27)(164) := previousCrc(4); xorBitMap(27)(165) := previousCrc(5); xorBitMap(27)(166) := previousCrc(6); xorBitMap(27)(168) := previousCrc(8); xorBitMap(27)(170) := previousCrc(10); xorBitMap(27)(171) := previousCrc(11); xorBitMap(27)(173) := previousCrc(13); xorBitMap(27)(177) := previousCrc(17); xorBitMap(27)(178) := previousCrc(18); xorBitMap(27)(180) := previousCrc(20); xorBitMap(27)(181) := previousCrc(21); xorBitMap(27)(183) := previousCrc(23); xorBitMap(27)(184) := previousCrc(24); xorBitMap(27)(185) := previousCrc(25); xorBitMap(27)(186) := previousCrc(26); xorBitMap(27)(190) := previousCrc(30); 
      xorBitMap(28)(119) := currentData(119); xorBitMap(28)(115) := currentData(115); xorBitMap(28)(114) := currentData(114); xorBitMap(28)(113) := currentData(113); xorBitMap(28)(112) := currentData(112); xorBitMap(28)(110) := currentData(110); xorBitMap(28)(109) := currentData(109); xorBitMap(28)(107) := currentData(107); xorBitMap(28)(106) := currentData(106); xorBitMap(28)(102) := currentData(102); xorBitMap(28)(100) := currentData(100); xorBitMap(28)(99) := currentData(99); xorBitMap(28)(97) := currentData(97); xorBitMap(28)(95) := currentData(95); xorBitMap(28)(94) := currentData(94); xorBitMap(28)(93) := currentData(93); xorBitMap(28)(92) := currentData(92); xorBitMap(28)(91) := currentData(91); xorBitMap(28)(90) := currentData(90); xorBitMap(28)(83) := currentData(83); xorBitMap(28)(81) := currentData(81); xorBitMap(28)(80) := currentData(80); xorBitMap(28)(79) := currentData(79); xorBitMap(28)(78) := currentData(78); xorBitMap(28)(77) := currentData(77); xorBitMap(28)(75) := currentData(75); xorBitMap(28)(69) := currentData(69); xorBitMap(28)(68) := currentData(68); xorBitMap(28)(64) := currentData(64); xorBitMap(28)(63) := currentData(63); xorBitMap(28)(62) := currentData(62); xorBitMap(28)(61) := currentData(61); xorBitMap(28)(59) := currentData(59); xorBitMap(28)(57) := currentData(57); xorBitMap(28)(56) := currentData(56); xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(162) := previousCrc(2); xorBitMap(28)(163) := previousCrc(3); xorBitMap(28)(164) := previousCrc(4); xorBitMap(28)(165) := previousCrc(5); xorBitMap(28)(166) := previousCrc(6); xorBitMap(28)(167) := previousCrc(7); xorBitMap(28)(169) := previousCrc(9); xorBitMap(28)(171) := previousCrc(11); xorBitMap(28)(172) := previousCrc(12); xorBitMap(28)(174) := previousCrc(14); xorBitMap(28)(178) := previousCrc(18); xorBitMap(28)(179) := previousCrc(19); xorBitMap(28)(181) := previousCrc(21); xorBitMap(28)(182) := previousCrc(22); xorBitMap(28)(184) := previousCrc(24); xorBitMap(28)(185) := previousCrc(25); xorBitMap(28)(186) := previousCrc(26); xorBitMap(28)(187) := previousCrc(27); xorBitMap(28)(191) := previousCrc(31); 
      xorBitMap(29)(116) := currentData(116); xorBitMap(29)(115) := currentData(115); xorBitMap(29)(114) := currentData(114); xorBitMap(29)(113) := currentData(113); xorBitMap(29)(111) := currentData(111); xorBitMap(29)(110) := currentData(110); xorBitMap(29)(108) := currentData(108); xorBitMap(29)(107) := currentData(107); xorBitMap(29)(103) := currentData(103); xorBitMap(29)(101) := currentData(101); xorBitMap(29)(100) := currentData(100); xorBitMap(29)(98) := currentData(98); xorBitMap(29)(96) := currentData(96); xorBitMap(29)(95) := currentData(95); xorBitMap(29)(94) := currentData(94); xorBitMap(29)(93) := currentData(93); xorBitMap(29)(92) := currentData(92); xorBitMap(29)(91) := currentData(91); xorBitMap(29)(84) := currentData(84); xorBitMap(29)(82) := currentData(82); xorBitMap(29)(81) := currentData(81); xorBitMap(29)(80) := currentData(80); xorBitMap(29)(79) := currentData(79); xorBitMap(29)(78) := currentData(78); xorBitMap(29)(76) := currentData(76); xorBitMap(29)(70) := currentData(70); xorBitMap(29)(69) := currentData(69); xorBitMap(29)(65) := currentData(65); xorBitMap(29)(64) := currentData(64); xorBitMap(29)(63) := currentData(63); xorBitMap(29)(62) := currentData(62); xorBitMap(29)(60) := currentData(60); xorBitMap(29)(58) := currentData(58); xorBitMap(29)(57) := currentData(57); xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(163) := previousCrc(3); xorBitMap(29)(164) := previousCrc(4); xorBitMap(29)(165) := previousCrc(5); xorBitMap(29)(166) := previousCrc(6); xorBitMap(29)(167) := previousCrc(7); xorBitMap(29)(168) := previousCrc(8); xorBitMap(29)(170) := previousCrc(10); xorBitMap(29)(172) := previousCrc(12); xorBitMap(29)(173) := previousCrc(13); xorBitMap(29)(175) := previousCrc(15); xorBitMap(29)(179) := previousCrc(19); xorBitMap(29)(180) := previousCrc(20); xorBitMap(29)(182) := previousCrc(22); xorBitMap(29)(183) := previousCrc(23); xorBitMap(29)(185) := previousCrc(25); xorBitMap(29)(186) := previousCrc(26); xorBitMap(29)(187) := previousCrc(27); xorBitMap(29)(188) := previousCrc(28); 
      xorBitMap(30)(117) := currentData(117); xorBitMap(30)(116) := currentData(116); xorBitMap(30)(115) := currentData(115); xorBitMap(30)(114) := currentData(114); xorBitMap(30)(112) := currentData(112); xorBitMap(30)(111) := currentData(111); xorBitMap(30)(109) := currentData(109); xorBitMap(30)(108) := currentData(108); xorBitMap(30)(104) := currentData(104); xorBitMap(30)(102) := currentData(102); xorBitMap(30)(101) := currentData(101); xorBitMap(30)(99) := currentData(99); xorBitMap(30)(97) := currentData(97); xorBitMap(30)(96) := currentData(96); xorBitMap(30)(95) := currentData(95); xorBitMap(30)(94) := currentData(94); xorBitMap(30)(93) := currentData(93); xorBitMap(30)(92) := currentData(92); xorBitMap(30)(85) := currentData(85); xorBitMap(30)(83) := currentData(83); xorBitMap(30)(82) := currentData(82); xorBitMap(30)(81) := currentData(81); xorBitMap(30)(80) := currentData(80); xorBitMap(30)(79) := currentData(79); xorBitMap(30)(77) := currentData(77); xorBitMap(30)(71) := currentData(71); xorBitMap(30)(70) := currentData(70); xorBitMap(30)(66) := currentData(66); xorBitMap(30)(65) := currentData(65); xorBitMap(30)(64) := currentData(64); xorBitMap(30)(63) := currentData(63); xorBitMap(30)(61) := currentData(61); xorBitMap(30)(59) := currentData(59); xorBitMap(30)(58) := currentData(58); xorBitMap(30)(56) := currentData(56); xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(164) := previousCrc(4); xorBitMap(30)(165) := previousCrc(5); xorBitMap(30)(166) := previousCrc(6); xorBitMap(30)(167) := previousCrc(7); xorBitMap(30)(168) := previousCrc(8); xorBitMap(30)(169) := previousCrc(9); xorBitMap(30)(171) := previousCrc(11); xorBitMap(30)(173) := previousCrc(13); xorBitMap(30)(174) := previousCrc(14); xorBitMap(30)(176) := previousCrc(16); xorBitMap(30)(180) := previousCrc(20); xorBitMap(30)(181) := previousCrc(21); xorBitMap(30)(183) := previousCrc(23); xorBitMap(30)(184) := previousCrc(24); xorBitMap(30)(186) := previousCrc(26); xorBitMap(30)(187) := previousCrc(27); xorBitMap(30)(188) := previousCrc(28); xorBitMap(30)(189) := previousCrc(29); 
      xorBitMap(31)(118) := currentData(118); xorBitMap(31)(117) := currentData(117); xorBitMap(31)(116) := currentData(116); xorBitMap(31)(115) := currentData(115); xorBitMap(31)(113) := currentData(113); xorBitMap(31)(112) := currentData(112); xorBitMap(31)(110) := currentData(110); xorBitMap(31)(109) := currentData(109); xorBitMap(31)(105) := currentData(105); xorBitMap(31)(103) := currentData(103); xorBitMap(31)(102) := currentData(102); xorBitMap(31)(100) := currentData(100); xorBitMap(31)(98) := currentData(98); xorBitMap(31)(97) := currentData(97); xorBitMap(31)(96) := currentData(96); xorBitMap(31)(95) := currentData(95); xorBitMap(31)(94) := currentData(94); xorBitMap(31)(93) := currentData(93); xorBitMap(31)(86) := currentData(86); xorBitMap(31)(84) := currentData(84); xorBitMap(31)(83) := currentData(83); xorBitMap(31)(82) := currentData(82); xorBitMap(31)(81) := currentData(81); xorBitMap(31)(80) := currentData(80); xorBitMap(31)(78) := currentData(78); xorBitMap(31)(72) := currentData(72); xorBitMap(31)(71) := currentData(71); xorBitMap(31)(67) := currentData(67); xorBitMap(31)(66) := currentData(66); xorBitMap(31)(65) := currentData(65); xorBitMap(31)(64) := currentData(64); xorBitMap(31)(62) := currentData(62); xorBitMap(31)(60) := currentData(60); xorBitMap(31)(59) := currentData(59); xorBitMap(31)(57) := currentData(57); xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(165) := previousCrc(5); xorBitMap(31)(166) := previousCrc(6); xorBitMap(31)(167) := previousCrc(7); xorBitMap(31)(168) := previousCrc(8); xorBitMap(31)(169) := previousCrc(9); xorBitMap(31)(170) := previousCrc(10); xorBitMap(31)(172) := previousCrc(12); xorBitMap(31)(174) := previousCrc(14); xorBitMap(31)(175) := previousCrc(15); xorBitMap(31)(177) := previousCrc(17); xorBitMap(31)(181) := previousCrc(21); xorBitMap(31)(182) := previousCrc(22); xorBitMap(31)(184) := previousCrc(24); xorBitMap(31)(185) := previousCrc(25); xorBitMap(31)(187) := previousCrc(27); xorBitMap(31)(188) := previousCrc(28); xorBitMap(31)(189) := previousCrc(29); xorBitMap(31)(190) := previousCrc(30); 
   end procedure;

   procedure xorBitMap16Byte (
      xorBitMap   : inout Slv192Array(31 downto 0);
      previousCrc : in    slv(31 downto 0);
      currentData : in    slv(127 downto 0)) is 
   begin
      xorBitMap(0)(127) := currentData(127); xorBitMap(0)(126) := currentData(126); xorBitMap(0)(125) := currentData(125); xorBitMap(0)(123) := currentData(123); xorBitMap(0)(119) := currentData(119); xorBitMap(0)(118) := currentData(118); xorBitMap(0)(117) := currentData(117); xorBitMap(0)(116) := currentData(116); xorBitMap(0)(114) := currentData(114); xorBitMap(0)(113) := currentData(113); xorBitMap(0)(111) := currentData(111); xorBitMap(0)(110) := currentData(110); xorBitMap(0)(106) := currentData(106); xorBitMap(0)(104) := currentData(104); xorBitMap(0)(103) := currentData(103); xorBitMap(0)(101) := currentData(101); xorBitMap(0)(99) := currentData(99); xorBitMap(0)(98) := currentData(98); xorBitMap(0)(97) := currentData(97); xorBitMap(0)(96) := currentData(96); xorBitMap(0)(95) := currentData(95); xorBitMap(0)(94) := currentData(94); xorBitMap(0)(87) := currentData(87); xorBitMap(0)(85) := currentData(85); xorBitMap(0)(84) := currentData(84); xorBitMap(0)(83) := currentData(83); xorBitMap(0)(82) := currentData(82); xorBitMap(0)(81) := currentData(81); xorBitMap(0)(79) := currentData(79); xorBitMap(0)(73) := currentData(73); xorBitMap(0)(72) := currentData(72); xorBitMap(0)(68) := currentData(68); xorBitMap(0)(67) := currentData(67); xorBitMap(0)(66) := currentData(66); xorBitMap(0)(65) := currentData(65); xorBitMap(0)(63) := currentData(63); xorBitMap(0)(61) := currentData(61); xorBitMap(0)(60) := currentData(60); xorBitMap(0)(58) := currentData(58); xorBitMap(0)(55) := currentData(55); xorBitMap(0)(54) := currentData(54); xorBitMap(0)(53) := currentData(53); xorBitMap(0)(50) := currentData(50); xorBitMap(0)(48) := currentData(48); xorBitMap(0)(47) := currentData(47); xorBitMap(0)(45) := currentData(45); xorBitMap(0)(44) := currentData(44); xorBitMap(0)(37) := currentData(37); xorBitMap(0)(34) := currentData(34); xorBitMap(0)(32) := currentData(32); xorBitMap(0)(31) := currentData(31); xorBitMap(0)(30) := currentData(30); xorBitMap(0)(29) := currentData(29); xorBitMap(0)(28) := currentData(28); xorBitMap(0)(26) := currentData(26); xorBitMap(0)(25) := currentData(25); xorBitMap(0)(24) := currentData(24); xorBitMap(0)(16) := currentData(16); xorBitMap(0)(12) := currentData(12); xorBitMap(0)(10) := currentData(10); xorBitMap(0)(9) := currentData(9); xorBitMap(0)(6) := currentData(6); xorBitMap(0)(0) := currentData(0); xorBitMap(0)(160) := previousCrc(0); xorBitMap(0)(161) := previousCrc(1); xorBitMap(0)(162) := previousCrc(2); xorBitMap(0)(163) := previousCrc(3); xorBitMap(0)(165) := previousCrc(5); xorBitMap(0)(167) := previousCrc(7); xorBitMap(0)(168) := previousCrc(8); xorBitMap(0)(170) := previousCrc(10); xorBitMap(0)(174) := previousCrc(14); xorBitMap(0)(175) := previousCrc(15); xorBitMap(0)(177) := previousCrc(17); xorBitMap(0)(178) := previousCrc(18); xorBitMap(0)(180) := previousCrc(20); xorBitMap(0)(181) := previousCrc(21); xorBitMap(0)(182) := previousCrc(22); xorBitMap(0)(183) := previousCrc(23); xorBitMap(0)(187) := previousCrc(27); xorBitMap(0)(189) := previousCrc(29); xorBitMap(0)(190) := previousCrc(30); xorBitMap(0)(191) := previousCrc(31); 
      xorBitMap(1)(125) := currentData(125); xorBitMap(1)(124) := currentData(124); xorBitMap(1)(123) := currentData(123); xorBitMap(1)(120) := currentData(120); xorBitMap(1)(116) := currentData(116); xorBitMap(1)(115) := currentData(115); xorBitMap(1)(113) := currentData(113); xorBitMap(1)(112) := currentData(112); xorBitMap(1)(110) := currentData(110); xorBitMap(1)(107) := currentData(107); xorBitMap(1)(106) := currentData(106); xorBitMap(1)(105) := currentData(105); xorBitMap(1)(103) := currentData(103); xorBitMap(1)(102) := currentData(102); xorBitMap(1)(101) := currentData(101); xorBitMap(1)(100) := currentData(100); xorBitMap(1)(94) := currentData(94); xorBitMap(1)(88) := currentData(88); xorBitMap(1)(87) := currentData(87); xorBitMap(1)(86) := currentData(86); xorBitMap(1)(81) := currentData(81); xorBitMap(1)(80) := currentData(80); xorBitMap(1)(79) := currentData(79); xorBitMap(1)(74) := currentData(74); xorBitMap(1)(72) := currentData(72); xorBitMap(1)(69) := currentData(69); xorBitMap(1)(65) := currentData(65); xorBitMap(1)(64) := currentData(64); xorBitMap(1)(63) := currentData(63); xorBitMap(1)(62) := currentData(62); xorBitMap(1)(60) := currentData(60); xorBitMap(1)(59) := currentData(59); xorBitMap(1)(58) := currentData(58); xorBitMap(1)(56) := currentData(56); xorBitMap(1)(53) := currentData(53); xorBitMap(1)(51) := currentData(51); xorBitMap(1)(50) := currentData(50); xorBitMap(1)(49) := currentData(49); xorBitMap(1)(47) := currentData(47); xorBitMap(1)(46) := currentData(46); xorBitMap(1)(44) := currentData(44); xorBitMap(1)(38) := currentData(38); xorBitMap(1)(37) := currentData(37); xorBitMap(1)(35) := currentData(35); xorBitMap(1)(34) := currentData(34); xorBitMap(1)(33) := currentData(33); xorBitMap(1)(28) := currentData(28); xorBitMap(1)(27) := currentData(27); xorBitMap(1)(24) := currentData(24); xorBitMap(1)(17) := currentData(17); xorBitMap(1)(16) := currentData(16); xorBitMap(1)(13) := currentData(13); xorBitMap(1)(12) := currentData(12); xorBitMap(1)(11) := currentData(11); xorBitMap(1)(9) := currentData(9); xorBitMap(1)(7) := currentData(7); xorBitMap(1)(6) := currentData(6); xorBitMap(1)(1) := currentData(1); xorBitMap(1)(0) := currentData(0); xorBitMap(1)(164) := previousCrc(4); xorBitMap(1)(165) := previousCrc(5); xorBitMap(1)(166) := previousCrc(6); xorBitMap(1)(167) := previousCrc(7); xorBitMap(1)(169) := previousCrc(9); xorBitMap(1)(170) := previousCrc(10); xorBitMap(1)(171) := previousCrc(11); xorBitMap(1)(174) := previousCrc(14); xorBitMap(1)(176) := previousCrc(16); xorBitMap(1)(177) := previousCrc(17); xorBitMap(1)(179) := previousCrc(19); xorBitMap(1)(180) := previousCrc(20); xorBitMap(1)(184) := previousCrc(24); xorBitMap(1)(187) := previousCrc(27); xorBitMap(1)(188) := previousCrc(28); xorBitMap(1)(189) := previousCrc(29); 
      xorBitMap(2)(127) := currentData(127); xorBitMap(2)(124) := currentData(124); xorBitMap(2)(123) := currentData(123); xorBitMap(2)(121) := currentData(121); xorBitMap(2)(119) := currentData(119); xorBitMap(2)(118) := currentData(118); xorBitMap(2)(110) := currentData(110); xorBitMap(2)(108) := currentData(108); xorBitMap(2)(107) := currentData(107); xorBitMap(2)(102) := currentData(102); xorBitMap(2)(99) := currentData(99); xorBitMap(2)(98) := currentData(98); xorBitMap(2)(97) := currentData(97); xorBitMap(2)(96) := currentData(96); xorBitMap(2)(94) := currentData(94); xorBitMap(2)(89) := currentData(89); xorBitMap(2)(88) := currentData(88); xorBitMap(2)(85) := currentData(85); xorBitMap(2)(84) := currentData(84); xorBitMap(2)(83) := currentData(83); xorBitMap(2)(80) := currentData(80); xorBitMap(2)(79) := currentData(79); xorBitMap(2)(75) := currentData(75); xorBitMap(2)(72) := currentData(72); xorBitMap(2)(70) := currentData(70); xorBitMap(2)(68) := currentData(68); xorBitMap(2)(67) := currentData(67); xorBitMap(2)(64) := currentData(64); xorBitMap(2)(59) := currentData(59); xorBitMap(2)(58) := currentData(58); xorBitMap(2)(57) := currentData(57); xorBitMap(2)(55) := currentData(55); xorBitMap(2)(53) := currentData(53); xorBitMap(2)(52) := currentData(52); xorBitMap(2)(51) := currentData(51); xorBitMap(2)(44) := currentData(44); xorBitMap(2)(39) := currentData(39); xorBitMap(2)(38) := currentData(38); xorBitMap(2)(37) := currentData(37); xorBitMap(2)(36) := currentData(36); xorBitMap(2)(35) := currentData(35); xorBitMap(2)(32) := currentData(32); xorBitMap(2)(31) := currentData(31); xorBitMap(2)(30) := currentData(30); xorBitMap(2)(26) := currentData(26); xorBitMap(2)(24) := currentData(24); xorBitMap(2)(18) := currentData(18); xorBitMap(2)(17) := currentData(17); xorBitMap(2)(16) := currentData(16); xorBitMap(2)(14) := currentData(14); xorBitMap(2)(13) := currentData(13); xorBitMap(2)(9) := currentData(9); xorBitMap(2)(8) := currentData(8); xorBitMap(2)(7) := currentData(7); xorBitMap(2)(6) := currentData(6); xorBitMap(2)(2) := currentData(2); xorBitMap(2)(1) := currentData(1); xorBitMap(2)(0) := currentData(0); xorBitMap(2)(160) := previousCrc(0); xorBitMap(2)(161) := previousCrc(1); xorBitMap(2)(162) := previousCrc(2); xorBitMap(2)(163) := previousCrc(3); xorBitMap(2)(166) := previousCrc(6); xorBitMap(2)(171) := previousCrc(11); xorBitMap(2)(172) := previousCrc(12); xorBitMap(2)(174) := previousCrc(14); xorBitMap(2)(182) := previousCrc(22); xorBitMap(2)(183) := previousCrc(23); xorBitMap(2)(185) := previousCrc(25); xorBitMap(2)(187) := previousCrc(27); xorBitMap(2)(188) := previousCrc(28); xorBitMap(2)(191) := previousCrc(31); 
      xorBitMap(3)(125) := currentData(125); xorBitMap(3)(124) := currentData(124); xorBitMap(3)(122) := currentData(122); xorBitMap(3)(120) := currentData(120); xorBitMap(3)(119) := currentData(119); xorBitMap(3)(111) := currentData(111); xorBitMap(3)(109) := currentData(109); xorBitMap(3)(108) := currentData(108); xorBitMap(3)(103) := currentData(103); xorBitMap(3)(100) := currentData(100); xorBitMap(3)(99) := currentData(99); xorBitMap(3)(98) := currentData(98); xorBitMap(3)(97) := currentData(97); xorBitMap(3)(95) := currentData(95); xorBitMap(3)(90) := currentData(90); xorBitMap(3)(89) := currentData(89); xorBitMap(3)(86) := currentData(86); xorBitMap(3)(85) := currentData(85); xorBitMap(3)(84) := currentData(84); xorBitMap(3)(81) := currentData(81); xorBitMap(3)(80) := currentData(80); xorBitMap(3)(76) := currentData(76); xorBitMap(3)(73) := currentData(73); xorBitMap(3)(71) := currentData(71); xorBitMap(3)(69) := currentData(69); xorBitMap(3)(68) := currentData(68); xorBitMap(3)(65) := currentData(65); xorBitMap(3)(60) := currentData(60); xorBitMap(3)(59) := currentData(59); xorBitMap(3)(58) := currentData(58); xorBitMap(3)(56) := currentData(56); xorBitMap(3)(54) := currentData(54); xorBitMap(3)(53) := currentData(53); xorBitMap(3)(52) := currentData(52); xorBitMap(3)(45) := currentData(45); xorBitMap(3)(40) := currentData(40); xorBitMap(3)(39) := currentData(39); xorBitMap(3)(38) := currentData(38); xorBitMap(3)(37) := currentData(37); xorBitMap(3)(36) := currentData(36); xorBitMap(3)(33) := currentData(33); xorBitMap(3)(32) := currentData(32); xorBitMap(3)(31) := currentData(31); xorBitMap(3)(27) := currentData(27); xorBitMap(3)(25) := currentData(25); xorBitMap(3)(19) := currentData(19); xorBitMap(3)(18) := currentData(18); xorBitMap(3)(17) := currentData(17); xorBitMap(3)(15) := currentData(15); xorBitMap(3)(14) := currentData(14); xorBitMap(3)(10) := currentData(10); xorBitMap(3)(9) := currentData(9); xorBitMap(3)(8) := currentData(8); xorBitMap(3)(7) := currentData(7); xorBitMap(3)(3) := currentData(3); xorBitMap(3)(2) := currentData(2); xorBitMap(3)(1) := currentData(1); xorBitMap(3)(161) := previousCrc(1); xorBitMap(3)(162) := previousCrc(2); xorBitMap(3)(163) := previousCrc(3); xorBitMap(3)(164) := previousCrc(4); xorBitMap(3)(167) := previousCrc(7); xorBitMap(3)(172) := previousCrc(12); xorBitMap(3)(173) := previousCrc(13); xorBitMap(3)(175) := previousCrc(15); xorBitMap(3)(183) := previousCrc(23); xorBitMap(3)(184) := previousCrc(24); xorBitMap(3)(186) := previousCrc(26); xorBitMap(3)(188) := previousCrc(28); xorBitMap(3)(189) := previousCrc(29); 
      xorBitMap(4)(127) := currentData(127); xorBitMap(4)(121) := currentData(121); xorBitMap(4)(120) := currentData(120); xorBitMap(4)(119) := currentData(119); xorBitMap(4)(118) := currentData(118); xorBitMap(4)(117) := currentData(117); xorBitMap(4)(116) := currentData(116); xorBitMap(4)(114) := currentData(114); xorBitMap(4)(113) := currentData(113); xorBitMap(4)(112) := currentData(112); xorBitMap(4)(111) := currentData(111); xorBitMap(4)(109) := currentData(109); xorBitMap(4)(106) := currentData(106); xorBitMap(4)(103) := currentData(103); xorBitMap(4)(100) := currentData(100); xorBitMap(4)(97) := currentData(97); xorBitMap(4)(95) := currentData(95); xorBitMap(4)(94) := currentData(94); xorBitMap(4)(91) := currentData(91); xorBitMap(4)(90) := currentData(90); xorBitMap(4)(86) := currentData(86); xorBitMap(4)(84) := currentData(84); xorBitMap(4)(83) := currentData(83); xorBitMap(4)(79) := currentData(79); xorBitMap(4)(77) := currentData(77); xorBitMap(4)(74) := currentData(74); xorBitMap(4)(73) := currentData(73); xorBitMap(4)(70) := currentData(70); xorBitMap(4)(69) := currentData(69); xorBitMap(4)(68) := currentData(68); xorBitMap(4)(67) := currentData(67); xorBitMap(4)(65) := currentData(65); xorBitMap(4)(63) := currentData(63); xorBitMap(4)(59) := currentData(59); xorBitMap(4)(58) := currentData(58); xorBitMap(4)(57) := currentData(57); xorBitMap(4)(50) := currentData(50); xorBitMap(4)(48) := currentData(48); xorBitMap(4)(47) := currentData(47); xorBitMap(4)(46) := currentData(46); xorBitMap(4)(45) := currentData(45); xorBitMap(4)(44) := currentData(44); xorBitMap(4)(41) := currentData(41); xorBitMap(4)(40) := currentData(40); xorBitMap(4)(39) := currentData(39); xorBitMap(4)(38) := currentData(38); xorBitMap(4)(33) := currentData(33); xorBitMap(4)(31) := currentData(31); xorBitMap(4)(30) := currentData(30); xorBitMap(4)(29) := currentData(29); xorBitMap(4)(25) := currentData(25); xorBitMap(4)(24) := currentData(24); xorBitMap(4)(20) := currentData(20); xorBitMap(4)(19) := currentData(19); xorBitMap(4)(18) := currentData(18); xorBitMap(4)(15) := currentData(15); xorBitMap(4)(12) := currentData(12); xorBitMap(4)(11) := currentData(11); xorBitMap(4)(8) := currentData(8); xorBitMap(4)(6) := currentData(6); xorBitMap(4)(4) := currentData(4); xorBitMap(4)(3) := currentData(3); xorBitMap(4)(2) := currentData(2); xorBitMap(4)(0) := currentData(0); xorBitMap(4)(161) := previousCrc(1); xorBitMap(4)(164) := previousCrc(4); xorBitMap(4)(167) := previousCrc(7); xorBitMap(4)(170) := previousCrc(10); xorBitMap(4)(173) := previousCrc(13); xorBitMap(4)(175) := previousCrc(15); xorBitMap(4)(176) := previousCrc(16); xorBitMap(4)(177) := previousCrc(17); xorBitMap(4)(178) := previousCrc(18); xorBitMap(4)(180) := previousCrc(20); xorBitMap(4)(181) := previousCrc(21); xorBitMap(4)(182) := previousCrc(22); xorBitMap(4)(183) := previousCrc(23); xorBitMap(4)(184) := previousCrc(24); xorBitMap(4)(185) := previousCrc(25); xorBitMap(4)(191) := previousCrc(31); 
      xorBitMap(5)(127) := currentData(127); xorBitMap(5)(126) := currentData(126); xorBitMap(5)(125) := currentData(125); xorBitMap(5)(123) := currentData(123); xorBitMap(5)(122) := currentData(122); xorBitMap(5)(121) := currentData(121); xorBitMap(5)(120) := currentData(120); xorBitMap(5)(116) := currentData(116); xorBitMap(5)(115) := currentData(115); xorBitMap(5)(112) := currentData(112); xorBitMap(5)(111) := currentData(111); xorBitMap(5)(107) := currentData(107); xorBitMap(5)(106) := currentData(106); xorBitMap(5)(103) := currentData(103); xorBitMap(5)(99) := currentData(99); xorBitMap(5)(97) := currentData(97); xorBitMap(5)(94) := currentData(94); xorBitMap(5)(92) := currentData(92); xorBitMap(5)(91) := currentData(91); xorBitMap(5)(83) := currentData(83); xorBitMap(5)(82) := currentData(82); xorBitMap(5)(81) := currentData(81); xorBitMap(5)(80) := currentData(80); xorBitMap(5)(79) := currentData(79); xorBitMap(5)(78) := currentData(78); xorBitMap(5)(75) := currentData(75); xorBitMap(5)(74) := currentData(74); xorBitMap(5)(73) := currentData(73); xorBitMap(5)(72) := currentData(72); xorBitMap(5)(71) := currentData(71); xorBitMap(5)(70) := currentData(70); xorBitMap(5)(69) := currentData(69); xorBitMap(5)(67) := currentData(67); xorBitMap(5)(65) := currentData(65); xorBitMap(5)(64) := currentData(64); xorBitMap(5)(63) := currentData(63); xorBitMap(5)(61) := currentData(61); xorBitMap(5)(59) := currentData(59); xorBitMap(5)(55) := currentData(55); xorBitMap(5)(54) := currentData(54); xorBitMap(5)(53) := currentData(53); xorBitMap(5)(51) := currentData(51); xorBitMap(5)(50) := currentData(50); xorBitMap(5)(49) := currentData(49); xorBitMap(5)(46) := currentData(46); xorBitMap(5)(44) := currentData(44); xorBitMap(5)(42) := currentData(42); xorBitMap(5)(41) := currentData(41); xorBitMap(5)(40) := currentData(40); xorBitMap(5)(39) := currentData(39); xorBitMap(5)(37) := currentData(37); xorBitMap(5)(29) := currentData(29); xorBitMap(5)(28) := currentData(28); xorBitMap(5)(24) := currentData(24); xorBitMap(5)(21) := currentData(21); xorBitMap(5)(20) := currentData(20); xorBitMap(5)(19) := currentData(19); xorBitMap(5)(13) := currentData(13); xorBitMap(5)(10) := currentData(10); xorBitMap(5)(7) := currentData(7); xorBitMap(5)(6) := currentData(6); xorBitMap(5)(5) := currentData(5); xorBitMap(5)(4) := currentData(4); xorBitMap(5)(3) := currentData(3); xorBitMap(5)(1) := currentData(1); xorBitMap(5)(0) := currentData(0); xorBitMap(5)(161) := previousCrc(1); xorBitMap(5)(163) := previousCrc(3); xorBitMap(5)(167) := previousCrc(7); xorBitMap(5)(170) := previousCrc(10); xorBitMap(5)(171) := previousCrc(11); xorBitMap(5)(175) := previousCrc(15); xorBitMap(5)(176) := previousCrc(16); xorBitMap(5)(179) := previousCrc(19); xorBitMap(5)(180) := previousCrc(20); xorBitMap(5)(184) := previousCrc(24); xorBitMap(5)(185) := previousCrc(25); xorBitMap(5)(186) := previousCrc(26); xorBitMap(5)(187) := previousCrc(27); xorBitMap(5)(189) := previousCrc(29); xorBitMap(5)(190) := previousCrc(30); xorBitMap(5)(191) := previousCrc(31); 
      xorBitMap(6)(127) := currentData(127); xorBitMap(6)(126) := currentData(126); xorBitMap(6)(124) := currentData(124); xorBitMap(6)(123) := currentData(123); xorBitMap(6)(122) := currentData(122); xorBitMap(6)(121) := currentData(121); xorBitMap(6)(117) := currentData(117); xorBitMap(6)(116) := currentData(116); xorBitMap(6)(113) := currentData(113); xorBitMap(6)(112) := currentData(112); xorBitMap(6)(108) := currentData(108); xorBitMap(6)(107) := currentData(107); xorBitMap(6)(104) := currentData(104); xorBitMap(6)(100) := currentData(100); xorBitMap(6)(98) := currentData(98); xorBitMap(6)(95) := currentData(95); xorBitMap(6)(93) := currentData(93); xorBitMap(6)(92) := currentData(92); xorBitMap(6)(84) := currentData(84); xorBitMap(6)(83) := currentData(83); xorBitMap(6)(82) := currentData(82); xorBitMap(6)(81) := currentData(81); xorBitMap(6)(80) := currentData(80); xorBitMap(6)(79) := currentData(79); xorBitMap(6)(76) := currentData(76); xorBitMap(6)(75) := currentData(75); xorBitMap(6)(74) := currentData(74); xorBitMap(6)(73) := currentData(73); xorBitMap(6)(72) := currentData(72); xorBitMap(6)(71) := currentData(71); xorBitMap(6)(70) := currentData(70); xorBitMap(6)(68) := currentData(68); xorBitMap(6)(66) := currentData(66); xorBitMap(6)(65) := currentData(65); xorBitMap(6)(64) := currentData(64); xorBitMap(6)(62) := currentData(62); xorBitMap(6)(60) := currentData(60); xorBitMap(6)(56) := currentData(56); xorBitMap(6)(55) := currentData(55); xorBitMap(6)(54) := currentData(54); xorBitMap(6)(52) := currentData(52); xorBitMap(6)(51) := currentData(51); xorBitMap(6)(50) := currentData(50); xorBitMap(6)(47) := currentData(47); xorBitMap(6)(45) := currentData(45); xorBitMap(6)(43) := currentData(43); xorBitMap(6)(42) := currentData(42); xorBitMap(6)(41) := currentData(41); xorBitMap(6)(40) := currentData(40); xorBitMap(6)(38) := currentData(38); xorBitMap(6)(30) := currentData(30); xorBitMap(6)(29) := currentData(29); xorBitMap(6)(25) := currentData(25); xorBitMap(6)(22) := currentData(22); xorBitMap(6)(21) := currentData(21); xorBitMap(6)(20) := currentData(20); xorBitMap(6)(14) := currentData(14); xorBitMap(6)(11) := currentData(11); xorBitMap(6)(8) := currentData(8); xorBitMap(6)(7) := currentData(7); xorBitMap(6)(6) := currentData(6); xorBitMap(6)(5) := currentData(5); xorBitMap(6)(4) := currentData(4); xorBitMap(6)(2) := currentData(2); xorBitMap(6)(1) := currentData(1); xorBitMap(6)(162) := previousCrc(2); xorBitMap(6)(164) := previousCrc(4); xorBitMap(6)(168) := previousCrc(8); xorBitMap(6)(171) := previousCrc(11); xorBitMap(6)(172) := previousCrc(12); xorBitMap(6)(176) := previousCrc(16); xorBitMap(6)(177) := previousCrc(17); xorBitMap(6)(180) := previousCrc(20); xorBitMap(6)(181) := previousCrc(21); xorBitMap(6)(185) := previousCrc(25); xorBitMap(6)(186) := previousCrc(26); xorBitMap(6)(187) := previousCrc(27); xorBitMap(6)(188) := previousCrc(28); xorBitMap(6)(190) := previousCrc(30); xorBitMap(6)(191) := previousCrc(31); 
      xorBitMap(7)(126) := currentData(126); xorBitMap(7)(124) := currentData(124); xorBitMap(7)(122) := currentData(122); xorBitMap(7)(119) := currentData(119); xorBitMap(7)(116) := currentData(116); xorBitMap(7)(111) := currentData(111); xorBitMap(7)(110) := currentData(110); xorBitMap(7)(109) := currentData(109); xorBitMap(7)(108) := currentData(108); xorBitMap(7)(106) := currentData(106); xorBitMap(7)(105) := currentData(105); xorBitMap(7)(104) := currentData(104); xorBitMap(7)(103) := currentData(103); xorBitMap(7)(98) := currentData(98); xorBitMap(7)(97) := currentData(97); xorBitMap(7)(95) := currentData(95); xorBitMap(7)(93) := currentData(93); xorBitMap(7)(87) := currentData(87); xorBitMap(7)(80) := currentData(80); xorBitMap(7)(79) := currentData(79); xorBitMap(7)(77) := currentData(77); xorBitMap(7)(76) := currentData(76); xorBitMap(7)(75) := currentData(75); xorBitMap(7)(74) := currentData(74); xorBitMap(7)(71) := currentData(71); xorBitMap(7)(69) := currentData(69); xorBitMap(7)(68) := currentData(68); xorBitMap(7)(60) := currentData(60); xorBitMap(7)(58) := currentData(58); xorBitMap(7)(57) := currentData(57); xorBitMap(7)(56) := currentData(56); xorBitMap(7)(54) := currentData(54); xorBitMap(7)(52) := currentData(52); xorBitMap(7)(51) := currentData(51); xorBitMap(7)(50) := currentData(50); xorBitMap(7)(47) := currentData(47); xorBitMap(7)(46) := currentData(46); xorBitMap(7)(45) := currentData(45); xorBitMap(7)(43) := currentData(43); xorBitMap(7)(42) := currentData(42); xorBitMap(7)(41) := currentData(41); xorBitMap(7)(39) := currentData(39); xorBitMap(7)(37) := currentData(37); xorBitMap(7)(34) := currentData(34); xorBitMap(7)(32) := currentData(32); xorBitMap(7)(29) := currentData(29); xorBitMap(7)(28) := currentData(28); xorBitMap(7)(25) := currentData(25); xorBitMap(7)(24) := currentData(24); xorBitMap(7)(23) := currentData(23); xorBitMap(7)(22) := currentData(22); xorBitMap(7)(21) := currentData(21); xorBitMap(7)(16) := currentData(16); xorBitMap(7)(15) := currentData(15); xorBitMap(7)(10) := currentData(10); xorBitMap(7)(8) := currentData(8); xorBitMap(7)(7) := currentData(7); xorBitMap(7)(5) := currentData(5); xorBitMap(7)(3) := currentData(3); xorBitMap(7)(2) := currentData(2); xorBitMap(7)(0) := currentData(0); xorBitMap(7)(161) := previousCrc(1); xorBitMap(7)(162) := previousCrc(2); xorBitMap(7)(167) := previousCrc(7); xorBitMap(7)(168) := previousCrc(8); xorBitMap(7)(169) := previousCrc(9); xorBitMap(7)(170) := previousCrc(10); xorBitMap(7)(172) := previousCrc(12); xorBitMap(7)(173) := previousCrc(13); xorBitMap(7)(174) := previousCrc(14); xorBitMap(7)(175) := previousCrc(15); xorBitMap(7)(180) := previousCrc(20); xorBitMap(7)(183) := previousCrc(23); xorBitMap(7)(186) := previousCrc(26); xorBitMap(7)(188) := previousCrc(28); xorBitMap(7)(190) := previousCrc(30); 
      xorBitMap(8)(126) := currentData(126); xorBitMap(8)(120) := currentData(120); xorBitMap(8)(119) := currentData(119); xorBitMap(8)(118) := currentData(118); xorBitMap(8)(116) := currentData(116); xorBitMap(8)(114) := currentData(114); xorBitMap(8)(113) := currentData(113); xorBitMap(8)(112) := currentData(112); xorBitMap(8)(109) := currentData(109); xorBitMap(8)(107) := currentData(107); xorBitMap(8)(105) := currentData(105); xorBitMap(8)(103) := currentData(103); xorBitMap(8)(101) := currentData(101); xorBitMap(8)(97) := currentData(97); xorBitMap(8)(95) := currentData(95); xorBitMap(8)(88) := currentData(88); xorBitMap(8)(87) := currentData(87); xorBitMap(8)(85) := currentData(85); xorBitMap(8)(84) := currentData(84); xorBitMap(8)(83) := currentData(83); xorBitMap(8)(82) := currentData(82); xorBitMap(8)(80) := currentData(80); xorBitMap(8)(79) := currentData(79); xorBitMap(8)(78) := currentData(78); xorBitMap(8)(77) := currentData(77); xorBitMap(8)(76) := currentData(76); xorBitMap(8)(75) := currentData(75); xorBitMap(8)(73) := currentData(73); xorBitMap(8)(70) := currentData(70); xorBitMap(8)(69) := currentData(69); xorBitMap(8)(68) := currentData(68); xorBitMap(8)(67) := currentData(67); xorBitMap(8)(66) := currentData(66); xorBitMap(8)(65) := currentData(65); xorBitMap(8)(63) := currentData(63); xorBitMap(8)(60) := currentData(60); xorBitMap(8)(59) := currentData(59); xorBitMap(8)(57) := currentData(57); xorBitMap(8)(54) := currentData(54); xorBitMap(8)(52) := currentData(52); xorBitMap(8)(51) := currentData(51); xorBitMap(8)(50) := currentData(50); xorBitMap(8)(46) := currentData(46); xorBitMap(8)(45) := currentData(45); xorBitMap(8)(43) := currentData(43); xorBitMap(8)(42) := currentData(42); xorBitMap(8)(40) := currentData(40); xorBitMap(8)(38) := currentData(38); xorBitMap(8)(37) := currentData(37); xorBitMap(8)(35) := currentData(35); xorBitMap(8)(34) := currentData(34); xorBitMap(8)(33) := currentData(33); xorBitMap(8)(32) := currentData(32); xorBitMap(8)(31) := currentData(31); xorBitMap(8)(28) := currentData(28); xorBitMap(8)(23) := currentData(23); xorBitMap(8)(22) := currentData(22); xorBitMap(8)(17) := currentData(17); xorBitMap(8)(12) := currentData(12); xorBitMap(8)(11) := currentData(11); xorBitMap(8)(10) := currentData(10); xorBitMap(8)(8) := currentData(8); xorBitMap(8)(4) := currentData(4); xorBitMap(8)(3) := currentData(3); xorBitMap(8)(1) := currentData(1); xorBitMap(8)(0) := currentData(0); xorBitMap(8)(161) := previousCrc(1); xorBitMap(8)(165) := previousCrc(5); xorBitMap(8)(167) := previousCrc(7); xorBitMap(8)(169) := previousCrc(9); xorBitMap(8)(171) := previousCrc(11); xorBitMap(8)(173) := previousCrc(13); xorBitMap(8)(176) := previousCrc(16); xorBitMap(8)(177) := previousCrc(17); xorBitMap(8)(178) := previousCrc(18); xorBitMap(8)(180) := previousCrc(20); xorBitMap(8)(182) := previousCrc(22); xorBitMap(8)(183) := previousCrc(23); xorBitMap(8)(184) := previousCrc(24); xorBitMap(8)(190) := previousCrc(30); 
      xorBitMap(9)(127) := currentData(127); xorBitMap(9)(121) := currentData(121); xorBitMap(9)(120) := currentData(120); xorBitMap(9)(119) := currentData(119); xorBitMap(9)(117) := currentData(117); xorBitMap(9)(115) := currentData(115); xorBitMap(9)(114) := currentData(114); xorBitMap(9)(113) := currentData(113); xorBitMap(9)(110) := currentData(110); xorBitMap(9)(108) := currentData(108); xorBitMap(9)(106) := currentData(106); xorBitMap(9)(104) := currentData(104); xorBitMap(9)(102) := currentData(102); xorBitMap(9)(98) := currentData(98); xorBitMap(9)(96) := currentData(96); xorBitMap(9)(89) := currentData(89); xorBitMap(9)(88) := currentData(88); xorBitMap(9)(86) := currentData(86); xorBitMap(9)(85) := currentData(85); xorBitMap(9)(84) := currentData(84); xorBitMap(9)(83) := currentData(83); xorBitMap(9)(81) := currentData(81); xorBitMap(9)(80) := currentData(80); xorBitMap(9)(79) := currentData(79); xorBitMap(9)(78) := currentData(78); xorBitMap(9)(77) := currentData(77); xorBitMap(9)(76) := currentData(76); xorBitMap(9)(74) := currentData(74); xorBitMap(9)(71) := currentData(71); xorBitMap(9)(70) := currentData(70); xorBitMap(9)(69) := currentData(69); xorBitMap(9)(68) := currentData(68); xorBitMap(9)(67) := currentData(67); xorBitMap(9)(66) := currentData(66); xorBitMap(9)(64) := currentData(64); xorBitMap(9)(61) := currentData(61); xorBitMap(9)(60) := currentData(60); xorBitMap(9)(58) := currentData(58); xorBitMap(9)(55) := currentData(55); xorBitMap(9)(53) := currentData(53); xorBitMap(9)(52) := currentData(52); xorBitMap(9)(51) := currentData(51); xorBitMap(9)(47) := currentData(47); xorBitMap(9)(46) := currentData(46); xorBitMap(9)(44) := currentData(44); xorBitMap(9)(43) := currentData(43); xorBitMap(9)(41) := currentData(41); xorBitMap(9)(39) := currentData(39); xorBitMap(9)(38) := currentData(38); xorBitMap(9)(36) := currentData(36); xorBitMap(9)(35) := currentData(35); xorBitMap(9)(34) := currentData(34); xorBitMap(9)(33) := currentData(33); xorBitMap(9)(32) := currentData(32); xorBitMap(9)(29) := currentData(29); xorBitMap(9)(24) := currentData(24); xorBitMap(9)(23) := currentData(23); xorBitMap(9)(18) := currentData(18); xorBitMap(9)(13) := currentData(13); xorBitMap(9)(12) := currentData(12); xorBitMap(9)(11) := currentData(11); xorBitMap(9)(9) := currentData(9); xorBitMap(9)(5) := currentData(5); xorBitMap(9)(4) := currentData(4); xorBitMap(9)(2) := currentData(2); xorBitMap(9)(1) := currentData(1); xorBitMap(9)(160) := previousCrc(0); xorBitMap(9)(162) := previousCrc(2); xorBitMap(9)(166) := previousCrc(6); xorBitMap(9)(168) := previousCrc(8); xorBitMap(9)(170) := previousCrc(10); xorBitMap(9)(172) := previousCrc(12); xorBitMap(9)(174) := previousCrc(14); xorBitMap(9)(177) := previousCrc(17); xorBitMap(9)(178) := previousCrc(18); xorBitMap(9)(179) := previousCrc(19); xorBitMap(9)(181) := previousCrc(21); xorBitMap(9)(183) := previousCrc(23); xorBitMap(9)(184) := previousCrc(24); xorBitMap(9)(185) := previousCrc(25); xorBitMap(9)(191) := previousCrc(31); 
      xorBitMap(10)(127) := currentData(127); xorBitMap(10)(126) := currentData(126); xorBitMap(10)(125) := currentData(125); xorBitMap(10)(123) := currentData(123); xorBitMap(10)(122) := currentData(122); xorBitMap(10)(121) := currentData(121); xorBitMap(10)(120) := currentData(120); xorBitMap(10)(119) := currentData(119); xorBitMap(10)(117) := currentData(117); xorBitMap(10)(115) := currentData(115); xorBitMap(10)(113) := currentData(113); xorBitMap(10)(110) := currentData(110); xorBitMap(10)(109) := currentData(109); xorBitMap(10)(107) := currentData(107); xorBitMap(10)(106) := currentData(106); xorBitMap(10)(105) := currentData(105); xorBitMap(10)(104) := currentData(104); xorBitMap(10)(101) := currentData(101); xorBitMap(10)(98) := currentData(98); xorBitMap(10)(96) := currentData(96); xorBitMap(10)(95) := currentData(95); xorBitMap(10)(94) := currentData(94); xorBitMap(10)(90) := currentData(90); xorBitMap(10)(89) := currentData(89); xorBitMap(10)(86) := currentData(86); xorBitMap(10)(83) := currentData(83); xorBitMap(10)(80) := currentData(80); xorBitMap(10)(78) := currentData(78); xorBitMap(10)(77) := currentData(77); xorBitMap(10)(75) := currentData(75); xorBitMap(10)(73) := currentData(73); xorBitMap(10)(71) := currentData(71); xorBitMap(10)(70) := currentData(70); xorBitMap(10)(69) := currentData(69); xorBitMap(10)(66) := currentData(66); xorBitMap(10)(63) := currentData(63); xorBitMap(10)(62) := currentData(62); xorBitMap(10)(60) := currentData(60); xorBitMap(10)(59) := currentData(59); xorBitMap(10)(58) := currentData(58); xorBitMap(10)(56) := currentData(56); xorBitMap(10)(55) := currentData(55); xorBitMap(10)(52) := currentData(52); xorBitMap(10)(50) := currentData(50); xorBitMap(10)(42) := currentData(42); xorBitMap(10)(40) := currentData(40); xorBitMap(10)(39) := currentData(39); xorBitMap(10)(36) := currentData(36); xorBitMap(10)(35) := currentData(35); xorBitMap(10)(33) := currentData(33); xorBitMap(10)(32) := currentData(32); xorBitMap(10)(31) := currentData(31); xorBitMap(10)(29) := currentData(29); xorBitMap(10)(28) := currentData(28); xorBitMap(10)(26) := currentData(26); xorBitMap(10)(19) := currentData(19); xorBitMap(10)(16) := currentData(16); xorBitMap(10)(14) := currentData(14); xorBitMap(10)(13) := currentData(13); xorBitMap(10)(9) := currentData(9); xorBitMap(10)(5) := currentData(5); xorBitMap(10)(3) := currentData(3); xorBitMap(10)(2) := currentData(2); xorBitMap(10)(0) := currentData(0); xorBitMap(10)(160) := previousCrc(0); xorBitMap(10)(162) := previousCrc(2); xorBitMap(10)(165) := previousCrc(5); xorBitMap(10)(168) := previousCrc(8); xorBitMap(10)(169) := previousCrc(9); xorBitMap(10)(170) := previousCrc(10); xorBitMap(10)(171) := previousCrc(11); xorBitMap(10)(173) := previousCrc(13); xorBitMap(10)(174) := previousCrc(14); xorBitMap(10)(177) := previousCrc(17); xorBitMap(10)(179) := previousCrc(19); xorBitMap(10)(181) := previousCrc(21); xorBitMap(10)(183) := previousCrc(23); xorBitMap(10)(184) := previousCrc(24); xorBitMap(10)(185) := previousCrc(25); xorBitMap(10)(186) := previousCrc(26); xorBitMap(10)(187) := previousCrc(27); xorBitMap(10)(189) := previousCrc(29); xorBitMap(10)(190) := previousCrc(30); xorBitMap(10)(191) := previousCrc(31); 
      xorBitMap(11)(125) := currentData(125); xorBitMap(11)(124) := currentData(124); xorBitMap(11)(122) := currentData(122); xorBitMap(11)(121) := currentData(121); xorBitMap(11)(120) := currentData(120); xorBitMap(11)(119) := currentData(119); xorBitMap(11)(117) := currentData(117); xorBitMap(11)(113) := currentData(113); xorBitMap(11)(108) := currentData(108); xorBitMap(11)(107) := currentData(107); xorBitMap(11)(105) := currentData(105); xorBitMap(11)(104) := currentData(104); xorBitMap(11)(103) := currentData(103); xorBitMap(11)(102) := currentData(102); xorBitMap(11)(101) := currentData(101); xorBitMap(11)(98) := currentData(98); xorBitMap(11)(94) := currentData(94); xorBitMap(11)(91) := currentData(91); xorBitMap(11)(90) := currentData(90); xorBitMap(11)(85) := currentData(85); xorBitMap(11)(83) := currentData(83); xorBitMap(11)(82) := currentData(82); xorBitMap(11)(78) := currentData(78); xorBitMap(11)(76) := currentData(76); xorBitMap(11)(74) := currentData(74); xorBitMap(11)(73) := currentData(73); xorBitMap(11)(71) := currentData(71); xorBitMap(11)(70) := currentData(70); xorBitMap(11)(68) := currentData(68); xorBitMap(11)(66) := currentData(66); xorBitMap(11)(65) := currentData(65); xorBitMap(11)(64) := currentData(64); xorBitMap(11)(59) := currentData(59); xorBitMap(11)(58) := currentData(58); xorBitMap(11)(57) := currentData(57); xorBitMap(11)(56) := currentData(56); xorBitMap(11)(55) := currentData(55); xorBitMap(11)(54) := currentData(54); xorBitMap(11)(51) := currentData(51); xorBitMap(11)(50) := currentData(50); xorBitMap(11)(48) := currentData(48); xorBitMap(11)(47) := currentData(47); xorBitMap(11)(45) := currentData(45); xorBitMap(11)(44) := currentData(44); xorBitMap(11)(43) := currentData(43); xorBitMap(11)(41) := currentData(41); xorBitMap(11)(40) := currentData(40); xorBitMap(11)(36) := currentData(36); xorBitMap(11)(33) := currentData(33); xorBitMap(11)(31) := currentData(31); xorBitMap(11)(28) := currentData(28); xorBitMap(11)(27) := currentData(27); xorBitMap(11)(26) := currentData(26); xorBitMap(11)(25) := currentData(25); xorBitMap(11)(24) := currentData(24); xorBitMap(11)(20) := currentData(20); xorBitMap(11)(17) := currentData(17); xorBitMap(11)(16) := currentData(16); xorBitMap(11)(15) := currentData(15); xorBitMap(11)(14) := currentData(14); xorBitMap(11)(12) := currentData(12); xorBitMap(11)(9) := currentData(9); xorBitMap(11)(4) := currentData(4); xorBitMap(11)(3) := currentData(3); xorBitMap(11)(1) := currentData(1); xorBitMap(11)(0) := currentData(0); xorBitMap(11)(162) := previousCrc(2); xorBitMap(11)(165) := previousCrc(5); xorBitMap(11)(166) := previousCrc(6); xorBitMap(11)(167) := previousCrc(7); xorBitMap(11)(168) := previousCrc(8); xorBitMap(11)(169) := previousCrc(9); xorBitMap(11)(171) := previousCrc(11); xorBitMap(11)(172) := previousCrc(12); xorBitMap(11)(177) := previousCrc(17); xorBitMap(11)(181) := previousCrc(21); xorBitMap(11)(183) := previousCrc(23); xorBitMap(11)(184) := previousCrc(24); xorBitMap(11)(185) := previousCrc(25); xorBitMap(11)(186) := previousCrc(26); xorBitMap(11)(188) := previousCrc(28); xorBitMap(11)(189) := previousCrc(29); 
      xorBitMap(12)(127) := currentData(127); xorBitMap(12)(122) := currentData(122); xorBitMap(12)(121) := currentData(121); xorBitMap(12)(120) := currentData(120); xorBitMap(12)(119) := currentData(119); xorBitMap(12)(117) := currentData(117); xorBitMap(12)(116) := currentData(116); xorBitMap(12)(113) := currentData(113); xorBitMap(12)(111) := currentData(111); xorBitMap(12)(110) := currentData(110); xorBitMap(12)(109) := currentData(109); xorBitMap(12)(108) := currentData(108); xorBitMap(12)(105) := currentData(105); xorBitMap(12)(102) := currentData(102); xorBitMap(12)(101) := currentData(101); xorBitMap(12)(98) := currentData(98); xorBitMap(12)(97) := currentData(97); xorBitMap(12)(96) := currentData(96); xorBitMap(12)(94) := currentData(94); xorBitMap(12)(92) := currentData(92); xorBitMap(12)(91) := currentData(91); xorBitMap(12)(87) := currentData(87); xorBitMap(12)(86) := currentData(86); xorBitMap(12)(85) := currentData(85); xorBitMap(12)(82) := currentData(82); xorBitMap(12)(81) := currentData(81); xorBitMap(12)(77) := currentData(77); xorBitMap(12)(75) := currentData(75); xorBitMap(12)(74) := currentData(74); xorBitMap(12)(73) := currentData(73); xorBitMap(12)(71) := currentData(71); xorBitMap(12)(69) := currentData(69); xorBitMap(12)(68) := currentData(68); xorBitMap(12)(63) := currentData(63); xorBitMap(12)(61) := currentData(61); xorBitMap(12)(59) := currentData(59); xorBitMap(12)(57) := currentData(57); xorBitMap(12)(56) := currentData(56); xorBitMap(12)(54) := currentData(54); xorBitMap(12)(53) := currentData(53); xorBitMap(12)(52) := currentData(52); xorBitMap(12)(51) := currentData(51); xorBitMap(12)(50) := currentData(50); xorBitMap(12)(49) := currentData(49); xorBitMap(12)(47) := currentData(47); xorBitMap(12)(46) := currentData(46); xorBitMap(12)(42) := currentData(42); xorBitMap(12)(41) := currentData(41); xorBitMap(12)(31) := currentData(31); xorBitMap(12)(30) := currentData(30); xorBitMap(12)(27) := currentData(27); xorBitMap(12)(24) := currentData(24); xorBitMap(12)(21) := currentData(21); xorBitMap(12)(18) := currentData(18); xorBitMap(12)(17) := currentData(17); xorBitMap(12)(15) := currentData(15); xorBitMap(12)(13) := currentData(13); xorBitMap(12)(12) := currentData(12); xorBitMap(12)(9) := currentData(9); xorBitMap(12)(6) := currentData(6); xorBitMap(12)(5) := currentData(5); xorBitMap(12)(4) := currentData(4); xorBitMap(12)(2) := currentData(2); xorBitMap(12)(1) := currentData(1); xorBitMap(12)(0) := currentData(0); xorBitMap(12)(160) := previousCrc(0); xorBitMap(12)(161) := previousCrc(1); xorBitMap(12)(162) := previousCrc(2); xorBitMap(12)(165) := previousCrc(5); xorBitMap(12)(166) := previousCrc(6); xorBitMap(12)(169) := previousCrc(9); xorBitMap(12)(172) := previousCrc(12); xorBitMap(12)(173) := previousCrc(13); xorBitMap(12)(174) := previousCrc(14); xorBitMap(12)(175) := previousCrc(15); xorBitMap(12)(177) := previousCrc(17); xorBitMap(12)(180) := previousCrc(20); xorBitMap(12)(181) := previousCrc(21); xorBitMap(12)(183) := previousCrc(23); xorBitMap(12)(184) := previousCrc(24); xorBitMap(12)(185) := previousCrc(25); xorBitMap(12)(186) := previousCrc(26); xorBitMap(12)(191) := previousCrc(31); 
      xorBitMap(13)(123) := currentData(123); xorBitMap(13)(122) := currentData(122); xorBitMap(13)(121) := currentData(121); xorBitMap(13)(120) := currentData(120); xorBitMap(13)(118) := currentData(118); xorBitMap(13)(117) := currentData(117); xorBitMap(13)(114) := currentData(114); xorBitMap(13)(112) := currentData(112); xorBitMap(13)(111) := currentData(111); xorBitMap(13)(110) := currentData(110); xorBitMap(13)(109) := currentData(109); xorBitMap(13)(106) := currentData(106); xorBitMap(13)(103) := currentData(103); xorBitMap(13)(102) := currentData(102); xorBitMap(13)(99) := currentData(99); xorBitMap(13)(98) := currentData(98); xorBitMap(13)(97) := currentData(97); xorBitMap(13)(95) := currentData(95); xorBitMap(13)(93) := currentData(93); xorBitMap(13)(92) := currentData(92); xorBitMap(13)(88) := currentData(88); xorBitMap(13)(87) := currentData(87); xorBitMap(13)(86) := currentData(86); xorBitMap(13)(83) := currentData(83); xorBitMap(13)(82) := currentData(82); xorBitMap(13)(78) := currentData(78); xorBitMap(13)(76) := currentData(76); xorBitMap(13)(75) := currentData(75); xorBitMap(13)(74) := currentData(74); xorBitMap(13)(72) := currentData(72); xorBitMap(13)(70) := currentData(70); xorBitMap(13)(69) := currentData(69); xorBitMap(13)(64) := currentData(64); xorBitMap(13)(62) := currentData(62); xorBitMap(13)(60) := currentData(60); xorBitMap(13)(58) := currentData(58); xorBitMap(13)(57) := currentData(57); xorBitMap(13)(55) := currentData(55); xorBitMap(13)(54) := currentData(54); xorBitMap(13)(53) := currentData(53); xorBitMap(13)(52) := currentData(52); xorBitMap(13)(51) := currentData(51); xorBitMap(13)(50) := currentData(50); xorBitMap(13)(48) := currentData(48); xorBitMap(13)(47) := currentData(47); xorBitMap(13)(43) := currentData(43); xorBitMap(13)(42) := currentData(42); xorBitMap(13)(32) := currentData(32); xorBitMap(13)(31) := currentData(31); xorBitMap(13)(28) := currentData(28); xorBitMap(13)(25) := currentData(25); xorBitMap(13)(22) := currentData(22); xorBitMap(13)(19) := currentData(19); xorBitMap(13)(18) := currentData(18); xorBitMap(13)(16) := currentData(16); xorBitMap(13)(14) := currentData(14); xorBitMap(13)(13) := currentData(13); xorBitMap(13)(10) := currentData(10); xorBitMap(13)(7) := currentData(7); xorBitMap(13)(6) := currentData(6); xorBitMap(13)(5) := currentData(5); xorBitMap(13)(3) := currentData(3); xorBitMap(13)(2) := currentData(2); xorBitMap(13)(1) := currentData(1); xorBitMap(13)(161) := previousCrc(1); xorBitMap(13)(162) := previousCrc(2); xorBitMap(13)(163) := previousCrc(3); xorBitMap(13)(166) := previousCrc(6); xorBitMap(13)(167) := previousCrc(7); xorBitMap(13)(170) := previousCrc(10); xorBitMap(13)(173) := previousCrc(13); xorBitMap(13)(174) := previousCrc(14); xorBitMap(13)(175) := previousCrc(15); xorBitMap(13)(176) := previousCrc(16); xorBitMap(13)(178) := previousCrc(18); xorBitMap(13)(181) := previousCrc(21); xorBitMap(13)(182) := previousCrc(22); xorBitMap(13)(184) := previousCrc(24); xorBitMap(13)(185) := previousCrc(25); xorBitMap(13)(186) := previousCrc(26); xorBitMap(13)(187) := previousCrc(27); 
      xorBitMap(14)(124) := currentData(124); xorBitMap(14)(123) := currentData(123); xorBitMap(14)(122) := currentData(122); xorBitMap(14)(121) := currentData(121); xorBitMap(14)(119) := currentData(119); xorBitMap(14)(118) := currentData(118); xorBitMap(14)(115) := currentData(115); xorBitMap(14)(113) := currentData(113); xorBitMap(14)(112) := currentData(112); xorBitMap(14)(111) := currentData(111); xorBitMap(14)(110) := currentData(110); xorBitMap(14)(107) := currentData(107); xorBitMap(14)(104) := currentData(104); xorBitMap(14)(103) := currentData(103); xorBitMap(14)(100) := currentData(100); xorBitMap(14)(99) := currentData(99); xorBitMap(14)(98) := currentData(98); xorBitMap(14)(96) := currentData(96); xorBitMap(14)(94) := currentData(94); xorBitMap(14)(93) := currentData(93); xorBitMap(14)(89) := currentData(89); xorBitMap(14)(88) := currentData(88); xorBitMap(14)(87) := currentData(87); xorBitMap(14)(84) := currentData(84); xorBitMap(14)(83) := currentData(83); xorBitMap(14)(79) := currentData(79); xorBitMap(14)(77) := currentData(77); xorBitMap(14)(76) := currentData(76); xorBitMap(14)(75) := currentData(75); xorBitMap(14)(73) := currentData(73); xorBitMap(14)(71) := currentData(71); xorBitMap(14)(70) := currentData(70); xorBitMap(14)(65) := currentData(65); xorBitMap(14)(63) := currentData(63); xorBitMap(14)(61) := currentData(61); xorBitMap(14)(59) := currentData(59); xorBitMap(14)(58) := currentData(58); xorBitMap(14)(56) := currentData(56); xorBitMap(14)(55) := currentData(55); xorBitMap(14)(54) := currentData(54); xorBitMap(14)(53) := currentData(53); xorBitMap(14)(52) := currentData(52); xorBitMap(14)(51) := currentData(51); xorBitMap(14)(49) := currentData(49); xorBitMap(14)(48) := currentData(48); xorBitMap(14)(44) := currentData(44); xorBitMap(14)(43) := currentData(43); xorBitMap(14)(33) := currentData(33); xorBitMap(14)(32) := currentData(32); xorBitMap(14)(29) := currentData(29); xorBitMap(14)(26) := currentData(26); xorBitMap(14)(23) := currentData(23); xorBitMap(14)(20) := currentData(20); xorBitMap(14)(19) := currentData(19); xorBitMap(14)(17) := currentData(17); xorBitMap(14)(15) := currentData(15); xorBitMap(14)(14) := currentData(14); xorBitMap(14)(11) := currentData(11); xorBitMap(14)(8) := currentData(8); xorBitMap(14)(7) := currentData(7); xorBitMap(14)(6) := currentData(6); xorBitMap(14)(4) := currentData(4); xorBitMap(14)(3) := currentData(3); xorBitMap(14)(2) := currentData(2); xorBitMap(14)(160) := previousCrc(0); xorBitMap(14)(162) := previousCrc(2); xorBitMap(14)(163) := previousCrc(3); xorBitMap(14)(164) := previousCrc(4); xorBitMap(14)(167) := previousCrc(7); xorBitMap(14)(168) := previousCrc(8); xorBitMap(14)(171) := previousCrc(11); xorBitMap(14)(174) := previousCrc(14); xorBitMap(14)(175) := previousCrc(15); xorBitMap(14)(176) := previousCrc(16); xorBitMap(14)(177) := previousCrc(17); xorBitMap(14)(179) := previousCrc(19); xorBitMap(14)(182) := previousCrc(22); xorBitMap(14)(183) := previousCrc(23); xorBitMap(14)(185) := previousCrc(25); xorBitMap(14)(186) := previousCrc(26); xorBitMap(14)(187) := previousCrc(27); xorBitMap(14)(188) := previousCrc(28); 
      xorBitMap(15)(125) := currentData(125); xorBitMap(15)(124) := currentData(124); xorBitMap(15)(123) := currentData(123); xorBitMap(15)(122) := currentData(122); xorBitMap(15)(120) := currentData(120); xorBitMap(15)(119) := currentData(119); xorBitMap(15)(116) := currentData(116); xorBitMap(15)(114) := currentData(114); xorBitMap(15)(113) := currentData(113); xorBitMap(15)(112) := currentData(112); xorBitMap(15)(111) := currentData(111); xorBitMap(15)(108) := currentData(108); xorBitMap(15)(105) := currentData(105); xorBitMap(15)(104) := currentData(104); xorBitMap(15)(101) := currentData(101); xorBitMap(15)(100) := currentData(100); xorBitMap(15)(99) := currentData(99); xorBitMap(15)(97) := currentData(97); xorBitMap(15)(95) := currentData(95); xorBitMap(15)(94) := currentData(94); xorBitMap(15)(90) := currentData(90); xorBitMap(15)(89) := currentData(89); xorBitMap(15)(88) := currentData(88); xorBitMap(15)(85) := currentData(85); xorBitMap(15)(84) := currentData(84); xorBitMap(15)(80) := currentData(80); xorBitMap(15)(78) := currentData(78); xorBitMap(15)(77) := currentData(77); xorBitMap(15)(76) := currentData(76); xorBitMap(15)(74) := currentData(74); xorBitMap(15)(72) := currentData(72); xorBitMap(15)(71) := currentData(71); xorBitMap(15)(66) := currentData(66); xorBitMap(15)(64) := currentData(64); xorBitMap(15)(62) := currentData(62); xorBitMap(15)(60) := currentData(60); xorBitMap(15)(59) := currentData(59); xorBitMap(15)(57) := currentData(57); xorBitMap(15)(56) := currentData(56); xorBitMap(15)(55) := currentData(55); xorBitMap(15)(54) := currentData(54); xorBitMap(15)(53) := currentData(53); xorBitMap(15)(52) := currentData(52); xorBitMap(15)(50) := currentData(50); xorBitMap(15)(49) := currentData(49); xorBitMap(15)(45) := currentData(45); xorBitMap(15)(44) := currentData(44); xorBitMap(15)(34) := currentData(34); xorBitMap(15)(33) := currentData(33); xorBitMap(15)(30) := currentData(30); xorBitMap(15)(27) := currentData(27); xorBitMap(15)(24) := currentData(24); xorBitMap(15)(21) := currentData(21); xorBitMap(15)(20) := currentData(20); xorBitMap(15)(18) := currentData(18); xorBitMap(15)(16) := currentData(16); xorBitMap(15)(15) := currentData(15); xorBitMap(15)(12) := currentData(12); xorBitMap(15)(9) := currentData(9); xorBitMap(15)(8) := currentData(8); xorBitMap(15)(7) := currentData(7); xorBitMap(15)(5) := currentData(5); xorBitMap(15)(4) := currentData(4); xorBitMap(15)(3) := currentData(3); xorBitMap(15)(161) := previousCrc(1); xorBitMap(15)(163) := previousCrc(3); xorBitMap(15)(164) := previousCrc(4); xorBitMap(15)(165) := previousCrc(5); xorBitMap(15)(168) := previousCrc(8); xorBitMap(15)(169) := previousCrc(9); xorBitMap(15)(172) := previousCrc(12); xorBitMap(15)(175) := previousCrc(15); xorBitMap(15)(176) := previousCrc(16); xorBitMap(15)(177) := previousCrc(17); xorBitMap(15)(178) := previousCrc(18); xorBitMap(15)(180) := previousCrc(20); xorBitMap(15)(183) := previousCrc(23); xorBitMap(15)(184) := previousCrc(24); xorBitMap(15)(186) := previousCrc(26); xorBitMap(15)(187) := previousCrc(27); xorBitMap(15)(188) := previousCrc(28); xorBitMap(15)(189) := previousCrc(29); 
      xorBitMap(16)(127) := currentData(127); xorBitMap(16)(124) := currentData(124); xorBitMap(16)(121) := currentData(121); xorBitMap(16)(120) := currentData(120); xorBitMap(16)(119) := currentData(119); xorBitMap(16)(118) := currentData(118); xorBitMap(16)(116) := currentData(116); xorBitMap(16)(115) := currentData(115); xorBitMap(16)(112) := currentData(112); xorBitMap(16)(111) := currentData(111); xorBitMap(16)(110) := currentData(110); xorBitMap(16)(109) := currentData(109); xorBitMap(16)(105) := currentData(105); xorBitMap(16)(104) := currentData(104); xorBitMap(16)(103) := currentData(103); xorBitMap(16)(102) := currentData(102); xorBitMap(16)(100) := currentData(100); xorBitMap(16)(99) := currentData(99); xorBitMap(16)(97) := currentData(97); xorBitMap(16)(94) := currentData(94); xorBitMap(16)(91) := currentData(91); xorBitMap(16)(90) := currentData(90); xorBitMap(16)(89) := currentData(89); xorBitMap(16)(87) := currentData(87); xorBitMap(16)(86) := currentData(86); xorBitMap(16)(84) := currentData(84); xorBitMap(16)(83) := currentData(83); xorBitMap(16)(82) := currentData(82); xorBitMap(16)(78) := currentData(78); xorBitMap(16)(77) := currentData(77); xorBitMap(16)(75) := currentData(75); xorBitMap(16)(68) := currentData(68); xorBitMap(16)(66) := currentData(66); xorBitMap(16)(57) := currentData(57); xorBitMap(16)(56) := currentData(56); xorBitMap(16)(51) := currentData(51); xorBitMap(16)(48) := currentData(48); xorBitMap(16)(47) := currentData(47); xorBitMap(16)(46) := currentData(46); xorBitMap(16)(44) := currentData(44); xorBitMap(16)(37) := currentData(37); xorBitMap(16)(35) := currentData(35); xorBitMap(16)(32) := currentData(32); xorBitMap(16)(30) := currentData(30); xorBitMap(16)(29) := currentData(29); xorBitMap(16)(26) := currentData(26); xorBitMap(16)(24) := currentData(24); xorBitMap(16)(22) := currentData(22); xorBitMap(16)(21) := currentData(21); xorBitMap(16)(19) := currentData(19); xorBitMap(16)(17) := currentData(17); xorBitMap(16)(13) := currentData(13); xorBitMap(16)(12) := currentData(12); xorBitMap(16)(8) := currentData(8); xorBitMap(16)(5) := currentData(5); xorBitMap(16)(4) := currentData(4); xorBitMap(16)(0) := currentData(0); xorBitMap(16)(161) := previousCrc(1); xorBitMap(16)(163) := previousCrc(3); xorBitMap(16)(164) := previousCrc(4); xorBitMap(16)(166) := previousCrc(6); xorBitMap(16)(167) := previousCrc(7); xorBitMap(16)(168) := previousCrc(8); xorBitMap(16)(169) := previousCrc(9); xorBitMap(16)(173) := previousCrc(13); xorBitMap(16)(174) := previousCrc(14); xorBitMap(16)(175) := previousCrc(15); xorBitMap(16)(176) := previousCrc(16); xorBitMap(16)(179) := previousCrc(19); xorBitMap(16)(180) := previousCrc(20); xorBitMap(16)(182) := previousCrc(22); xorBitMap(16)(183) := previousCrc(23); xorBitMap(16)(184) := previousCrc(24); xorBitMap(16)(185) := previousCrc(25); xorBitMap(16)(188) := previousCrc(28); xorBitMap(16)(191) := previousCrc(31); 
      xorBitMap(17)(125) := currentData(125); xorBitMap(17)(122) := currentData(122); xorBitMap(17)(121) := currentData(121); xorBitMap(17)(120) := currentData(120); xorBitMap(17)(119) := currentData(119); xorBitMap(17)(117) := currentData(117); xorBitMap(17)(116) := currentData(116); xorBitMap(17)(113) := currentData(113); xorBitMap(17)(112) := currentData(112); xorBitMap(17)(111) := currentData(111); xorBitMap(17)(110) := currentData(110); xorBitMap(17)(106) := currentData(106); xorBitMap(17)(105) := currentData(105); xorBitMap(17)(104) := currentData(104); xorBitMap(17)(103) := currentData(103); xorBitMap(17)(101) := currentData(101); xorBitMap(17)(100) := currentData(100); xorBitMap(17)(98) := currentData(98); xorBitMap(17)(95) := currentData(95); xorBitMap(17)(92) := currentData(92); xorBitMap(17)(91) := currentData(91); xorBitMap(17)(90) := currentData(90); xorBitMap(17)(88) := currentData(88); xorBitMap(17)(87) := currentData(87); xorBitMap(17)(85) := currentData(85); xorBitMap(17)(84) := currentData(84); xorBitMap(17)(83) := currentData(83); xorBitMap(17)(79) := currentData(79); xorBitMap(17)(78) := currentData(78); xorBitMap(17)(76) := currentData(76); xorBitMap(17)(69) := currentData(69); xorBitMap(17)(67) := currentData(67); xorBitMap(17)(58) := currentData(58); xorBitMap(17)(57) := currentData(57); xorBitMap(17)(52) := currentData(52); xorBitMap(17)(49) := currentData(49); xorBitMap(17)(48) := currentData(48); xorBitMap(17)(47) := currentData(47); xorBitMap(17)(45) := currentData(45); xorBitMap(17)(38) := currentData(38); xorBitMap(17)(36) := currentData(36); xorBitMap(17)(33) := currentData(33); xorBitMap(17)(31) := currentData(31); xorBitMap(17)(30) := currentData(30); xorBitMap(17)(27) := currentData(27); xorBitMap(17)(25) := currentData(25); xorBitMap(17)(23) := currentData(23); xorBitMap(17)(22) := currentData(22); xorBitMap(17)(20) := currentData(20); xorBitMap(17)(18) := currentData(18); xorBitMap(17)(14) := currentData(14); xorBitMap(17)(13) := currentData(13); xorBitMap(17)(9) := currentData(9); xorBitMap(17)(6) := currentData(6); xorBitMap(17)(5) := currentData(5); xorBitMap(17)(1) := currentData(1); xorBitMap(17)(162) := previousCrc(2); xorBitMap(17)(164) := previousCrc(4); xorBitMap(17)(165) := previousCrc(5); xorBitMap(17)(167) := previousCrc(7); xorBitMap(17)(168) := previousCrc(8); xorBitMap(17)(169) := previousCrc(9); xorBitMap(17)(170) := previousCrc(10); xorBitMap(17)(174) := previousCrc(14); xorBitMap(17)(175) := previousCrc(15); xorBitMap(17)(176) := previousCrc(16); xorBitMap(17)(177) := previousCrc(17); xorBitMap(17)(180) := previousCrc(20); xorBitMap(17)(181) := previousCrc(21); xorBitMap(17)(183) := previousCrc(23); xorBitMap(17)(184) := previousCrc(24); xorBitMap(17)(185) := previousCrc(25); xorBitMap(17)(186) := previousCrc(26); xorBitMap(17)(189) := previousCrc(29); 
      xorBitMap(18)(126) := currentData(126); xorBitMap(18)(123) := currentData(123); xorBitMap(18)(122) := currentData(122); xorBitMap(18)(121) := currentData(121); xorBitMap(18)(120) := currentData(120); xorBitMap(18)(118) := currentData(118); xorBitMap(18)(117) := currentData(117); xorBitMap(18)(114) := currentData(114); xorBitMap(18)(113) := currentData(113); xorBitMap(18)(112) := currentData(112); xorBitMap(18)(111) := currentData(111); xorBitMap(18)(107) := currentData(107); xorBitMap(18)(106) := currentData(106); xorBitMap(18)(105) := currentData(105); xorBitMap(18)(104) := currentData(104); xorBitMap(18)(102) := currentData(102); xorBitMap(18)(101) := currentData(101); xorBitMap(18)(99) := currentData(99); xorBitMap(18)(96) := currentData(96); xorBitMap(18)(93) := currentData(93); xorBitMap(18)(92) := currentData(92); xorBitMap(18)(91) := currentData(91); xorBitMap(18)(89) := currentData(89); xorBitMap(18)(88) := currentData(88); xorBitMap(18)(86) := currentData(86); xorBitMap(18)(85) := currentData(85); xorBitMap(18)(84) := currentData(84); xorBitMap(18)(80) := currentData(80); xorBitMap(18)(79) := currentData(79); xorBitMap(18)(77) := currentData(77); xorBitMap(18)(70) := currentData(70); xorBitMap(18)(68) := currentData(68); xorBitMap(18)(59) := currentData(59); xorBitMap(18)(58) := currentData(58); xorBitMap(18)(53) := currentData(53); xorBitMap(18)(50) := currentData(50); xorBitMap(18)(49) := currentData(49); xorBitMap(18)(48) := currentData(48); xorBitMap(18)(46) := currentData(46); xorBitMap(18)(39) := currentData(39); xorBitMap(18)(37) := currentData(37); xorBitMap(18)(34) := currentData(34); xorBitMap(18)(32) := currentData(32); xorBitMap(18)(31) := currentData(31); xorBitMap(18)(28) := currentData(28); xorBitMap(18)(26) := currentData(26); xorBitMap(18)(24) := currentData(24); xorBitMap(18)(23) := currentData(23); xorBitMap(18)(21) := currentData(21); xorBitMap(18)(19) := currentData(19); xorBitMap(18)(15) := currentData(15); xorBitMap(18)(14) := currentData(14); xorBitMap(18)(10) := currentData(10); xorBitMap(18)(7) := currentData(7); xorBitMap(18)(6) := currentData(6); xorBitMap(18)(2) := currentData(2); xorBitMap(18)(160) := previousCrc(0); xorBitMap(18)(163) := previousCrc(3); xorBitMap(18)(165) := previousCrc(5); xorBitMap(18)(166) := previousCrc(6); xorBitMap(18)(168) := previousCrc(8); xorBitMap(18)(169) := previousCrc(9); xorBitMap(18)(170) := previousCrc(10); xorBitMap(18)(171) := previousCrc(11); xorBitMap(18)(175) := previousCrc(15); xorBitMap(18)(176) := previousCrc(16); xorBitMap(18)(177) := previousCrc(17); xorBitMap(18)(178) := previousCrc(18); xorBitMap(18)(181) := previousCrc(21); xorBitMap(18)(182) := previousCrc(22); xorBitMap(18)(184) := previousCrc(24); xorBitMap(18)(185) := previousCrc(25); xorBitMap(18)(186) := previousCrc(26); xorBitMap(18)(187) := previousCrc(27); xorBitMap(18)(190) := previousCrc(30); 
      xorBitMap(19)(127) := currentData(127); xorBitMap(19)(124) := currentData(124); xorBitMap(19)(123) := currentData(123); xorBitMap(19)(122) := currentData(122); xorBitMap(19)(121) := currentData(121); xorBitMap(19)(119) := currentData(119); xorBitMap(19)(118) := currentData(118); xorBitMap(19)(115) := currentData(115); xorBitMap(19)(114) := currentData(114); xorBitMap(19)(113) := currentData(113); xorBitMap(19)(112) := currentData(112); xorBitMap(19)(108) := currentData(108); xorBitMap(19)(107) := currentData(107); xorBitMap(19)(106) := currentData(106); xorBitMap(19)(105) := currentData(105); xorBitMap(19)(103) := currentData(103); xorBitMap(19)(102) := currentData(102); xorBitMap(19)(100) := currentData(100); xorBitMap(19)(97) := currentData(97); xorBitMap(19)(94) := currentData(94); xorBitMap(19)(93) := currentData(93); xorBitMap(19)(92) := currentData(92); xorBitMap(19)(90) := currentData(90); xorBitMap(19)(89) := currentData(89); xorBitMap(19)(87) := currentData(87); xorBitMap(19)(86) := currentData(86); xorBitMap(19)(85) := currentData(85); xorBitMap(19)(81) := currentData(81); xorBitMap(19)(80) := currentData(80); xorBitMap(19)(78) := currentData(78); xorBitMap(19)(71) := currentData(71); xorBitMap(19)(69) := currentData(69); xorBitMap(19)(60) := currentData(60); xorBitMap(19)(59) := currentData(59); xorBitMap(19)(54) := currentData(54); xorBitMap(19)(51) := currentData(51); xorBitMap(19)(50) := currentData(50); xorBitMap(19)(49) := currentData(49); xorBitMap(19)(47) := currentData(47); xorBitMap(19)(40) := currentData(40); xorBitMap(19)(38) := currentData(38); xorBitMap(19)(35) := currentData(35); xorBitMap(19)(33) := currentData(33); xorBitMap(19)(32) := currentData(32); xorBitMap(19)(29) := currentData(29); xorBitMap(19)(27) := currentData(27); xorBitMap(19)(25) := currentData(25); xorBitMap(19)(24) := currentData(24); xorBitMap(19)(22) := currentData(22); xorBitMap(19)(20) := currentData(20); xorBitMap(19)(16) := currentData(16); xorBitMap(19)(15) := currentData(15); xorBitMap(19)(11) := currentData(11); xorBitMap(19)(8) := currentData(8); xorBitMap(19)(7) := currentData(7); xorBitMap(19)(3) := currentData(3); xorBitMap(19)(161) := previousCrc(1); xorBitMap(19)(164) := previousCrc(4); xorBitMap(19)(166) := previousCrc(6); xorBitMap(19)(167) := previousCrc(7); xorBitMap(19)(169) := previousCrc(9); xorBitMap(19)(170) := previousCrc(10); xorBitMap(19)(171) := previousCrc(11); xorBitMap(19)(172) := previousCrc(12); xorBitMap(19)(176) := previousCrc(16); xorBitMap(19)(177) := previousCrc(17); xorBitMap(19)(178) := previousCrc(18); xorBitMap(19)(179) := previousCrc(19); xorBitMap(19)(182) := previousCrc(22); xorBitMap(19)(183) := previousCrc(23); xorBitMap(19)(185) := previousCrc(25); xorBitMap(19)(186) := previousCrc(26); xorBitMap(19)(187) := previousCrc(27); xorBitMap(19)(188) := previousCrc(28); xorBitMap(19)(191) := previousCrc(31); 
      xorBitMap(20)(125) := currentData(125); xorBitMap(20)(124) := currentData(124); xorBitMap(20)(123) := currentData(123); xorBitMap(20)(122) := currentData(122); xorBitMap(20)(120) := currentData(120); xorBitMap(20)(119) := currentData(119); xorBitMap(20)(116) := currentData(116); xorBitMap(20)(115) := currentData(115); xorBitMap(20)(114) := currentData(114); xorBitMap(20)(113) := currentData(113); xorBitMap(20)(109) := currentData(109); xorBitMap(20)(108) := currentData(108); xorBitMap(20)(107) := currentData(107); xorBitMap(20)(106) := currentData(106); xorBitMap(20)(104) := currentData(104); xorBitMap(20)(103) := currentData(103); xorBitMap(20)(101) := currentData(101); xorBitMap(20)(98) := currentData(98); xorBitMap(20)(95) := currentData(95); xorBitMap(20)(94) := currentData(94); xorBitMap(20)(93) := currentData(93); xorBitMap(20)(91) := currentData(91); xorBitMap(20)(90) := currentData(90); xorBitMap(20)(88) := currentData(88); xorBitMap(20)(87) := currentData(87); xorBitMap(20)(86) := currentData(86); xorBitMap(20)(82) := currentData(82); xorBitMap(20)(81) := currentData(81); xorBitMap(20)(79) := currentData(79); xorBitMap(20)(72) := currentData(72); xorBitMap(20)(70) := currentData(70); xorBitMap(20)(61) := currentData(61); xorBitMap(20)(60) := currentData(60); xorBitMap(20)(55) := currentData(55); xorBitMap(20)(52) := currentData(52); xorBitMap(20)(51) := currentData(51); xorBitMap(20)(50) := currentData(50); xorBitMap(20)(48) := currentData(48); xorBitMap(20)(41) := currentData(41); xorBitMap(20)(39) := currentData(39); xorBitMap(20)(36) := currentData(36); xorBitMap(20)(34) := currentData(34); xorBitMap(20)(33) := currentData(33); xorBitMap(20)(30) := currentData(30); xorBitMap(20)(28) := currentData(28); xorBitMap(20)(26) := currentData(26); xorBitMap(20)(25) := currentData(25); xorBitMap(20)(23) := currentData(23); xorBitMap(20)(21) := currentData(21); xorBitMap(20)(17) := currentData(17); xorBitMap(20)(16) := currentData(16); xorBitMap(20)(12) := currentData(12); xorBitMap(20)(9) := currentData(9); xorBitMap(20)(8) := currentData(8); xorBitMap(20)(4) := currentData(4); xorBitMap(20)(162) := previousCrc(2); xorBitMap(20)(165) := previousCrc(5); xorBitMap(20)(167) := previousCrc(7); xorBitMap(20)(168) := previousCrc(8); xorBitMap(20)(170) := previousCrc(10); xorBitMap(20)(171) := previousCrc(11); xorBitMap(20)(172) := previousCrc(12); xorBitMap(20)(173) := previousCrc(13); xorBitMap(20)(177) := previousCrc(17); xorBitMap(20)(178) := previousCrc(18); xorBitMap(20)(179) := previousCrc(19); xorBitMap(20)(180) := previousCrc(20); xorBitMap(20)(183) := previousCrc(23); xorBitMap(20)(184) := previousCrc(24); xorBitMap(20)(186) := previousCrc(26); xorBitMap(20)(187) := previousCrc(27); xorBitMap(20)(188) := previousCrc(28); xorBitMap(20)(189) := previousCrc(29); 
      xorBitMap(21)(126) := currentData(126); xorBitMap(21)(125) := currentData(125); xorBitMap(21)(124) := currentData(124); xorBitMap(21)(123) := currentData(123); xorBitMap(21)(121) := currentData(121); xorBitMap(21)(120) := currentData(120); xorBitMap(21)(117) := currentData(117); xorBitMap(21)(116) := currentData(116); xorBitMap(21)(115) := currentData(115); xorBitMap(21)(114) := currentData(114); xorBitMap(21)(110) := currentData(110); xorBitMap(21)(109) := currentData(109); xorBitMap(21)(108) := currentData(108); xorBitMap(21)(107) := currentData(107); xorBitMap(21)(105) := currentData(105); xorBitMap(21)(104) := currentData(104); xorBitMap(21)(102) := currentData(102); xorBitMap(21)(99) := currentData(99); xorBitMap(21)(96) := currentData(96); xorBitMap(21)(95) := currentData(95); xorBitMap(21)(94) := currentData(94); xorBitMap(21)(92) := currentData(92); xorBitMap(21)(91) := currentData(91); xorBitMap(21)(89) := currentData(89); xorBitMap(21)(88) := currentData(88); xorBitMap(21)(87) := currentData(87); xorBitMap(21)(83) := currentData(83); xorBitMap(21)(82) := currentData(82); xorBitMap(21)(80) := currentData(80); xorBitMap(21)(73) := currentData(73); xorBitMap(21)(71) := currentData(71); xorBitMap(21)(62) := currentData(62); xorBitMap(21)(61) := currentData(61); xorBitMap(21)(56) := currentData(56); xorBitMap(21)(53) := currentData(53); xorBitMap(21)(52) := currentData(52); xorBitMap(21)(51) := currentData(51); xorBitMap(21)(49) := currentData(49); xorBitMap(21)(42) := currentData(42); xorBitMap(21)(40) := currentData(40); xorBitMap(21)(37) := currentData(37); xorBitMap(21)(35) := currentData(35); xorBitMap(21)(34) := currentData(34); xorBitMap(21)(31) := currentData(31); xorBitMap(21)(29) := currentData(29); xorBitMap(21)(27) := currentData(27); xorBitMap(21)(26) := currentData(26); xorBitMap(21)(24) := currentData(24); xorBitMap(21)(22) := currentData(22); xorBitMap(21)(18) := currentData(18); xorBitMap(21)(17) := currentData(17); xorBitMap(21)(13) := currentData(13); xorBitMap(21)(10) := currentData(10); xorBitMap(21)(9) := currentData(9); xorBitMap(21)(5) := currentData(5); xorBitMap(21)(160) := previousCrc(0); xorBitMap(21)(163) := previousCrc(3); xorBitMap(21)(166) := previousCrc(6); xorBitMap(21)(168) := previousCrc(8); xorBitMap(21)(169) := previousCrc(9); xorBitMap(21)(171) := previousCrc(11); xorBitMap(21)(172) := previousCrc(12); xorBitMap(21)(173) := previousCrc(13); xorBitMap(21)(174) := previousCrc(14); xorBitMap(21)(178) := previousCrc(18); xorBitMap(21)(179) := previousCrc(19); xorBitMap(21)(180) := previousCrc(20); xorBitMap(21)(181) := previousCrc(21); xorBitMap(21)(184) := previousCrc(24); xorBitMap(21)(185) := previousCrc(25); xorBitMap(21)(187) := previousCrc(27); xorBitMap(21)(188) := previousCrc(28); xorBitMap(21)(189) := previousCrc(29); xorBitMap(21)(190) := previousCrc(30); 
      xorBitMap(22)(124) := currentData(124); xorBitMap(22)(123) := currentData(123); xorBitMap(22)(122) := currentData(122); xorBitMap(22)(121) := currentData(121); xorBitMap(22)(119) := currentData(119); xorBitMap(22)(115) := currentData(115); xorBitMap(22)(114) := currentData(114); xorBitMap(22)(113) := currentData(113); xorBitMap(22)(109) := currentData(109); xorBitMap(22)(108) := currentData(108); xorBitMap(22)(105) := currentData(105); xorBitMap(22)(104) := currentData(104); xorBitMap(22)(101) := currentData(101); xorBitMap(22)(100) := currentData(100); xorBitMap(22)(99) := currentData(99); xorBitMap(22)(98) := currentData(98); xorBitMap(22)(94) := currentData(94); xorBitMap(22)(93) := currentData(93); xorBitMap(22)(92) := currentData(92); xorBitMap(22)(90) := currentData(90); xorBitMap(22)(89) := currentData(89); xorBitMap(22)(88) := currentData(88); xorBitMap(22)(87) := currentData(87); xorBitMap(22)(85) := currentData(85); xorBitMap(22)(82) := currentData(82); xorBitMap(22)(79) := currentData(79); xorBitMap(22)(74) := currentData(74); xorBitMap(22)(73) := currentData(73); xorBitMap(22)(68) := currentData(68); xorBitMap(22)(67) := currentData(67); xorBitMap(22)(66) := currentData(66); xorBitMap(22)(65) := currentData(65); xorBitMap(22)(62) := currentData(62); xorBitMap(22)(61) := currentData(61); xorBitMap(22)(60) := currentData(60); xorBitMap(22)(58) := currentData(58); xorBitMap(22)(57) := currentData(57); xorBitMap(22)(55) := currentData(55); xorBitMap(22)(52) := currentData(52); xorBitMap(22)(48) := currentData(48); xorBitMap(22)(47) := currentData(47); xorBitMap(22)(45) := currentData(45); xorBitMap(22)(44) := currentData(44); xorBitMap(22)(43) := currentData(43); xorBitMap(22)(41) := currentData(41); xorBitMap(22)(38) := currentData(38); xorBitMap(22)(37) := currentData(37); xorBitMap(22)(36) := currentData(36); xorBitMap(22)(35) := currentData(35); xorBitMap(22)(34) := currentData(34); xorBitMap(22)(31) := currentData(31); xorBitMap(22)(29) := currentData(29); xorBitMap(22)(27) := currentData(27); xorBitMap(22)(26) := currentData(26); xorBitMap(22)(24) := currentData(24); xorBitMap(22)(23) := currentData(23); xorBitMap(22)(19) := currentData(19); xorBitMap(22)(18) := currentData(18); xorBitMap(22)(16) := currentData(16); xorBitMap(22)(14) := currentData(14); xorBitMap(22)(12) := currentData(12); xorBitMap(22)(11) := currentData(11); xorBitMap(22)(9) := currentData(9); xorBitMap(22)(0) := currentData(0); xorBitMap(22)(162) := previousCrc(2); xorBitMap(22)(163) := previousCrc(3); xorBitMap(22)(164) := previousCrc(4); xorBitMap(22)(165) := previousCrc(5); xorBitMap(22)(168) := previousCrc(8); xorBitMap(22)(169) := previousCrc(9); xorBitMap(22)(172) := previousCrc(12); xorBitMap(22)(173) := previousCrc(13); xorBitMap(22)(177) := previousCrc(17); xorBitMap(22)(178) := previousCrc(18); xorBitMap(22)(179) := previousCrc(19); xorBitMap(22)(183) := previousCrc(23); xorBitMap(22)(185) := previousCrc(25); xorBitMap(22)(186) := previousCrc(26); xorBitMap(22)(187) := previousCrc(27); xorBitMap(22)(188) := previousCrc(28); 
      xorBitMap(23)(127) := currentData(127); xorBitMap(23)(126) := currentData(126); xorBitMap(23)(124) := currentData(124); xorBitMap(23)(122) := currentData(122); xorBitMap(23)(120) := currentData(120); xorBitMap(23)(119) := currentData(119); xorBitMap(23)(118) := currentData(118); xorBitMap(23)(117) := currentData(117); xorBitMap(23)(115) := currentData(115); xorBitMap(23)(113) := currentData(113); xorBitMap(23)(111) := currentData(111); xorBitMap(23)(109) := currentData(109); xorBitMap(23)(105) := currentData(105); xorBitMap(23)(104) := currentData(104); xorBitMap(23)(103) := currentData(103); xorBitMap(23)(102) := currentData(102); xorBitMap(23)(100) := currentData(100); xorBitMap(23)(98) := currentData(98); xorBitMap(23)(97) := currentData(97); xorBitMap(23)(96) := currentData(96); xorBitMap(23)(93) := currentData(93); xorBitMap(23)(91) := currentData(91); xorBitMap(23)(90) := currentData(90); xorBitMap(23)(89) := currentData(89); xorBitMap(23)(88) := currentData(88); xorBitMap(23)(87) := currentData(87); xorBitMap(23)(86) := currentData(86); xorBitMap(23)(85) := currentData(85); xorBitMap(23)(84) := currentData(84); xorBitMap(23)(82) := currentData(82); xorBitMap(23)(81) := currentData(81); xorBitMap(23)(80) := currentData(80); xorBitMap(23)(79) := currentData(79); xorBitMap(23)(75) := currentData(75); xorBitMap(23)(74) := currentData(74); xorBitMap(23)(73) := currentData(73); xorBitMap(23)(72) := currentData(72); xorBitMap(23)(69) := currentData(69); xorBitMap(23)(65) := currentData(65); xorBitMap(23)(62) := currentData(62); xorBitMap(23)(60) := currentData(60); xorBitMap(23)(59) := currentData(59); xorBitMap(23)(56) := currentData(56); xorBitMap(23)(55) := currentData(55); xorBitMap(23)(54) := currentData(54); xorBitMap(23)(50) := currentData(50); xorBitMap(23)(49) := currentData(49); xorBitMap(23)(47) := currentData(47); xorBitMap(23)(46) := currentData(46); xorBitMap(23)(42) := currentData(42); xorBitMap(23)(39) := currentData(39); xorBitMap(23)(38) := currentData(38); xorBitMap(23)(36) := currentData(36); xorBitMap(23)(35) := currentData(35); xorBitMap(23)(34) := currentData(34); xorBitMap(23)(31) := currentData(31); xorBitMap(23)(29) := currentData(29); xorBitMap(23)(27) := currentData(27); xorBitMap(23)(26) := currentData(26); xorBitMap(23)(20) := currentData(20); xorBitMap(23)(19) := currentData(19); xorBitMap(23)(17) := currentData(17); xorBitMap(23)(16) := currentData(16); xorBitMap(23)(15) := currentData(15); xorBitMap(23)(13) := currentData(13); xorBitMap(23)(9) := currentData(9); xorBitMap(23)(6) := currentData(6); xorBitMap(23)(1) := currentData(1); xorBitMap(23)(0) := currentData(0); xorBitMap(23)(160) := previousCrc(0); xorBitMap(23)(161) := previousCrc(1); xorBitMap(23)(162) := previousCrc(2); xorBitMap(23)(164) := previousCrc(4); xorBitMap(23)(166) := previousCrc(6); xorBitMap(23)(167) := previousCrc(7); xorBitMap(23)(168) := previousCrc(8); xorBitMap(23)(169) := previousCrc(9); xorBitMap(23)(173) := previousCrc(13); xorBitMap(23)(175) := previousCrc(15); xorBitMap(23)(177) := previousCrc(17); xorBitMap(23)(179) := previousCrc(19); xorBitMap(23)(181) := previousCrc(21); xorBitMap(23)(182) := previousCrc(22); xorBitMap(23)(183) := previousCrc(23); xorBitMap(23)(184) := previousCrc(24); xorBitMap(23)(186) := previousCrc(26); xorBitMap(23)(188) := previousCrc(28); xorBitMap(23)(190) := previousCrc(30); xorBitMap(23)(191) := previousCrc(31); 
      xorBitMap(24)(127) := currentData(127); xorBitMap(24)(125) := currentData(125); xorBitMap(24)(123) := currentData(123); xorBitMap(24)(121) := currentData(121); xorBitMap(24)(120) := currentData(120); xorBitMap(24)(119) := currentData(119); xorBitMap(24)(118) := currentData(118); xorBitMap(24)(116) := currentData(116); xorBitMap(24)(114) := currentData(114); xorBitMap(24)(112) := currentData(112); xorBitMap(24)(110) := currentData(110); xorBitMap(24)(106) := currentData(106); xorBitMap(24)(105) := currentData(105); xorBitMap(24)(104) := currentData(104); xorBitMap(24)(103) := currentData(103); xorBitMap(24)(101) := currentData(101); xorBitMap(24)(99) := currentData(99); xorBitMap(24)(98) := currentData(98); xorBitMap(24)(97) := currentData(97); xorBitMap(24)(94) := currentData(94); xorBitMap(24)(92) := currentData(92); xorBitMap(24)(91) := currentData(91); xorBitMap(24)(90) := currentData(90); xorBitMap(24)(89) := currentData(89); xorBitMap(24)(88) := currentData(88); xorBitMap(24)(87) := currentData(87); xorBitMap(24)(86) := currentData(86); xorBitMap(24)(85) := currentData(85); xorBitMap(24)(83) := currentData(83); xorBitMap(24)(82) := currentData(82); xorBitMap(24)(81) := currentData(81); xorBitMap(24)(80) := currentData(80); xorBitMap(24)(76) := currentData(76); xorBitMap(24)(75) := currentData(75); xorBitMap(24)(74) := currentData(74); xorBitMap(24)(73) := currentData(73); xorBitMap(24)(70) := currentData(70); xorBitMap(24)(66) := currentData(66); xorBitMap(24)(63) := currentData(63); xorBitMap(24)(61) := currentData(61); xorBitMap(24)(60) := currentData(60); xorBitMap(24)(57) := currentData(57); xorBitMap(24)(56) := currentData(56); xorBitMap(24)(55) := currentData(55); xorBitMap(24)(51) := currentData(51); xorBitMap(24)(50) := currentData(50); xorBitMap(24)(48) := currentData(48); xorBitMap(24)(47) := currentData(47); xorBitMap(24)(43) := currentData(43); xorBitMap(24)(40) := currentData(40); xorBitMap(24)(39) := currentData(39); xorBitMap(24)(37) := currentData(37); xorBitMap(24)(36) := currentData(36); xorBitMap(24)(35) := currentData(35); xorBitMap(24)(32) := currentData(32); xorBitMap(24)(30) := currentData(30); xorBitMap(24)(28) := currentData(28); xorBitMap(24)(27) := currentData(27); xorBitMap(24)(21) := currentData(21); xorBitMap(24)(20) := currentData(20); xorBitMap(24)(18) := currentData(18); xorBitMap(24)(17) := currentData(17); xorBitMap(24)(16) := currentData(16); xorBitMap(24)(14) := currentData(14); xorBitMap(24)(10) := currentData(10); xorBitMap(24)(7) := currentData(7); xorBitMap(24)(2) := currentData(2); xorBitMap(24)(1) := currentData(1); xorBitMap(24)(161) := previousCrc(1); xorBitMap(24)(162) := previousCrc(2); xorBitMap(24)(163) := previousCrc(3); xorBitMap(24)(165) := previousCrc(5); xorBitMap(24)(167) := previousCrc(7); xorBitMap(24)(168) := previousCrc(8); xorBitMap(24)(169) := previousCrc(9); xorBitMap(24)(170) := previousCrc(10); xorBitMap(24)(174) := previousCrc(14); xorBitMap(24)(176) := previousCrc(16); xorBitMap(24)(178) := previousCrc(18); xorBitMap(24)(180) := previousCrc(20); xorBitMap(24)(182) := previousCrc(22); xorBitMap(24)(183) := previousCrc(23); xorBitMap(24)(184) := previousCrc(24); xorBitMap(24)(185) := previousCrc(25); xorBitMap(24)(187) := previousCrc(27); xorBitMap(24)(189) := previousCrc(29); xorBitMap(24)(191) := previousCrc(31); 
      xorBitMap(25)(126) := currentData(126); xorBitMap(25)(124) := currentData(124); xorBitMap(25)(122) := currentData(122); xorBitMap(25)(121) := currentData(121); xorBitMap(25)(120) := currentData(120); xorBitMap(25)(119) := currentData(119); xorBitMap(25)(117) := currentData(117); xorBitMap(25)(115) := currentData(115); xorBitMap(25)(113) := currentData(113); xorBitMap(25)(111) := currentData(111); xorBitMap(25)(107) := currentData(107); xorBitMap(25)(106) := currentData(106); xorBitMap(25)(105) := currentData(105); xorBitMap(25)(104) := currentData(104); xorBitMap(25)(102) := currentData(102); xorBitMap(25)(100) := currentData(100); xorBitMap(25)(99) := currentData(99); xorBitMap(25)(98) := currentData(98); xorBitMap(25)(95) := currentData(95); xorBitMap(25)(93) := currentData(93); xorBitMap(25)(92) := currentData(92); xorBitMap(25)(91) := currentData(91); xorBitMap(25)(90) := currentData(90); xorBitMap(25)(89) := currentData(89); xorBitMap(25)(88) := currentData(88); xorBitMap(25)(87) := currentData(87); xorBitMap(25)(86) := currentData(86); xorBitMap(25)(84) := currentData(84); xorBitMap(25)(83) := currentData(83); xorBitMap(25)(82) := currentData(82); xorBitMap(25)(81) := currentData(81); xorBitMap(25)(77) := currentData(77); xorBitMap(25)(76) := currentData(76); xorBitMap(25)(75) := currentData(75); xorBitMap(25)(74) := currentData(74); xorBitMap(25)(71) := currentData(71); xorBitMap(25)(67) := currentData(67); xorBitMap(25)(64) := currentData(64); xorBitMap(25)(62) := currentData(62); xorBitMap(25)(61) := currentData(61); xorBitMap(25)(58) := currentData(58); xorBitMap(25)(57) := currentData(57); xorBitMap(25)(56) := currentData(56); xorBitMap(25)(52) := currentData(52); xorBitMap(25)(51) := currentData(51); xorBitMap(25)(49) := currentData(49); xorBitMap(25)(48) := currentData(48); xorBitMap(25)(44) := currentData(44); xorBitMap(25)(41) := currentData(41); xorBitMap(25)(40) := currentData(40); xorBitMap(25)(38) := currentData(38); xorBitMap(25)(37) := currentData(37); xorBitMap(25)(36) := currentData(36); xorBitMap(25)(33) := currentData(33); xorBitMap(25)(31) := currentData(31); xorBitMap(25)(29) := currentData(29); xorBitMap(25)(28) := currentData(28); xorBitMap(25)(22) := currentData(22); xorBitMap(25)(21) := currentData(21); xorBitMap(25)(19) := currentData(19); xorBitMap(25)(18) := currentData(18); xorBitMap(25)(17) := currentData(17); xorBitMap(25)(15) := currentData(15); xorBitMap(25)(11) := currentData(11); xorBitMap(25)(8) := currentData(8); xorBitMap(25)(3) := currentData(3); xorBitMap(25)(2) := currentData(2); xorBitMap(25)(162) := previousCrc(2); xorBitMap(25)(163) := previousCrc(3); xorBitMap(25)(164) := previousCrc(4); xorBitMap(25)(166) := previousCrc(6); xorBitMap(25)(168) := previousCrc(8); xorBitMap(25)(169) := previousCrc(9); xorBitMap(25)(170) := previousCrc(10); xorBitMap(25)(171) := previousCrc(11); xorBitMap(25)(175) := previousCrc(15); xorBitMap(25)(177) := previousCrc(17); xorBitMap(25)(179) := previousCrc(19); xorBitMap(25)(181) := previousCrc(21); xorBitMap(25)(183) := previousCrc(23); xorBitMap(25)(184) := previousCrc(24); xorBitMap(25)(185) := previousCrc(25); xorBitMap(25)(186) := previousCrc(26); xorBitMap(25)(188) := previousCrc(28); xorBitMap(25)(190) := previousCrc(30); 
      xorBitMap(26)(126) := currentData(126); xorBitMap(26)(122) := currentData(122); xorBitMap(26)(121) := currentData(121); xorBitMap(26)(120) := currentData(120); xorBitMap(26)(119) := currentData(119); xorBitMap(26)(117) := currentData(117); xorBitMap(26)(113) := currentData(113); xorBitMap(26)(112) := currentData(112); xorBitMap(26)(111) := currentData(111); xorBitMap(26)(110) := currentData(110); xorBitMap(26)(108) := currentData(108); xorBitMap(26)(107) := currentData(107); xorBitMap(26)(105) := currentData(105); xorBitMap(26)(104) := currentData(104); xorBitMap(26)(100) := currentData(100); xorBitMap(26)(98) := currentData(98); xorBitMap(26)(97) := currentData(97); xorBitMap(26)(95) := currentData(95); xorBitMap(26)(93) := currentData(93); xorBitMap(26)(92) := currentData(92); xorBitMap(26)(91) := currentData(91); xorBitMap(26)(90) := currentData(90); xorBitMap(26)(89) := currentData(89); xorBitMap(26)(88) := currentData(88); xorBitMap(26)(81) := currentData(81); xorBitMap(26)(79) := currentData(79); xorBitMap(26)(78) := currentData(78); xorBitMap(26)(77) := currentData(77); xorBitMap(26)(76) := currentData(76); xorBitMap(26)(75) := currentData(75); xorBitMap(26)(73) := currentData(73); xorBitMap(26)(67) := currentData(67); xorBitMap(26)(66) := currentData(66); xorBitMap(26)(62) := currentData(62); xorBitMap(26)(61) := currentData(61); xorBitMap(26)(60) := currentData(60); xorBitMap(26)(59) := currentData(59); xorBitMap(26)(57) := currentData(57); xorBitMap(26)(55) := currentData(55); xorBitMap(26)(54) := currentData(54); xorBitMap(26)(52) := currentData(52); xorBitMap(26)(49) := currentData(49); xorBitMap(26)(48) := currentData(48); xorBitMap(26)(47) := currentData(47); xorBitMap(26)(44) := currentData(44); xorBitMap(26)(42) := currentData(42); xorBitMap(26)(41) := currentData(41); xorBitMap(26)(39) := currentData(39); xorBitMap(26)(38) := currentData(38); xorBitMap(26)(31) := currentData(31); xorBitMap(26)(28) := currentData(28); xorBitMap(26)(26) := currentData(26); xorBitMap(26)(25) := currentData(25); xorBitMap(26)(24) := currentData(24); xorBitMap(26)(23) := currentData(23); xorBitMap(26)(22) := currentData(22); xorBitMap(26)(20) := currentData(20); xorBitMap(26)(19) := currentData(19); xorBitMap(26)(18) := currentData(18); xorBitMap(26)(10) := currentData(10); xorBitMap(26)(6) := currentData(6); xorBitMap(26)(4) := currentData(4); xorBitMap(26)(3) := currentData(3); xorBitMap(26)(0) := currentData(0); xorBitMap(26)(161) := previousCrc(1); xorBitMap(26)(162) := previousCrc(2); xorBitMap(26)(164) := previousCrc(4); xorBitMap(26)(168) := previousCrc(8); xorBitMap(26)(169) := previousCrc(9); xorBitMap(26)(171) := previousCrc(11); xorBitMap(26)(172) := previousCrc(12); xorBitMap(26)(174) := previousCrc(14); xorBitMap(26)(175) := previousCrc(15); xorBitMap(26)(176) := previousCrc(16); xorBitMap(26)(177) := previousCrc(17); xorBitMap(26)(181) := previousCrc(21); xorBitMap(26)(183) := previousCrc(23); xorBitMap(26)(184) := previousCrc(24); xorBitMap(26)(185) := previousCrc(25); xorBitMap(26)(186) := previousCrc(26); xorBitMap(26)(190) := previousCrc(30); 
      xorBitMap(27)(127) := currentData(127); xorBitMap(27)(123) := currentData(123); xorBitMap(27)(122) := currentData(122); xorBitMap(27)(121) := currentData(121); xorBitMap(27)(120) := currentData(120); xorBitMap(27)(118) := currentData(118); xorBitMap(27)(114) := currentData(114); xorBitMap(27)(113) := currentData(113); xorBitMap(27)(112) := currentData(112); xorBitMap(27)(111) := currentData(111); xorBitMap(27)(109) := currentData(109); xorBitMap(27)(108) := currentData(108); xorBitMap(27)(106) := currentData(106); xorBitMap(27)(105) := currentData(105); xorBitMap(27)(101) := currentData(101); xorBitMap(27)(99) := currentData(99); xorBitMap(27)(98) := currentData(98); xorBitMap(27)(96) := currentData(96); xorBitMap(27)(94) := currentData(94); xorBitMap(27)(93) := currentData(93); xorBitMap(27)(92) := currentData(92); xorBitMap(27)(91) := currentData(91); xorBitMap(27)(90) := currentData(90); xorBitMap(27)(89) := currentData(89); xorBitMap(27)(82) := currentData(82); xorBitMap(27)(80) := currentData(80); xorBitMap(27)(79) := currentData(79); xorBitMap(27)(78) := currentData(78); xorBitMap(27)(77) := currentData(77); xorBitMap(27)(76) := currentData(76); xorBitMap(27)(74) := currentData(74); xorBitMap(27)(68) := currentData(68); xorBitMap(27)(67) := currentData(67); xorBitMap(27)(63) := currentData(63); xorBitMap(27)(62) := currentData(62); xorBitMap(27)(61) := currentData(61); xorBitMap(27)(60) := currentData(60); xorBitMap(27)(58) := currentData(58); xorBitMap(27)(56) := currentData(56); xorBitMap(27)(55) := currentData(55); xorBitMap(27)(53) := currentData(53); xorBitMap(27)(50) := currentData(50); xorBitMap(27)(49) := currentData(49); xorBitMap(27)(48) := currentData(48); xorBitMap(27)(45) := currentData(45); xorBitMap(27)(43) := currentData(43); xorBitMap(27)(42) := currentData(42); xorBitMap(27)(40) := currentData(40); xorBitMap(27)(39) := currentData(39); xorBitMap(27)(32) := currentData(32); xorBitMap(27)(29) := currentData(29); xorBitMap(27)(27) := currentData(27); xorBitMap(27)(26) := currentData(26); xorBitMap(27)(25) := currentData(25); xorBitMap(27)(24) := currentData(24); xorBitMap(27)(23) := currentData(23); xorBitMap(27)(21) := currentData(21); xorBitMap(27)(20) := currentData(20); xorBitMap(27)(19) := currentData(19); xorBitMap(27)(11) := currentData(11); xorBitMap(27)(7) := currentData(7); xorBitMap(27)(5) := currentData(5); xorBitMap(27)(4) := currentData(4); xorBitMap(27)(1) := currentData(1); xorBitMap(27)(160) := previousCrc(0); xorBitMap(27)(162) := previousCrc(2); xorBitMap(27)(163) := previousCrc(3); xorBitMap(27)(165) := previousCrc(5); xorBitMap(27)(169) := previousCrc(9); xorBitMap(27)(170) := previousCrc(10); xorBitMap(27)(172) := previousCrc(12); xorBitMap(27)(173) := previousCrc(13); xorBitMap(27)(175) := previousCrc(15); xorBitMap(27)(176) := previousCrc(16); xorBitMap(27)(177) := previousCrc(17); xorBitMap(27)(178) := previousCrc(18); xorBitMap(27)(182) := previousCrc(22); xorBitMap(27)(184) := previousCrc(24); xorBitMap(27)(185) := previousCrc(25); xorBitMap(27)(186) := previousCrc(26); xorBitMap(27)(187) := previousCrc(27); xorBitMap(27)(191) := previousCrc(31); 
      xorBitMap(28)(124) := currentData(124); xorBitMap(28)(123) := currentData(123); xorBitMap(28)(122) := currentData(122); xorBitMap(28)(121) := currentData(121); xorBitMap(28)(119) := currentData(119); xorBitMap(28)(115) := currentData(115); xorBitMap(28)(114) := currentData(114); xorBitMap(28)(113) := currentData(113); xorBitMap(28)(112) := currentData(112); xorBitMap(28)(110) := currentData(110); xorBitMap(28)(109) := currentData(109); xorBitMap(28)(107) := currentData(107); xorBitMap(28)(106) := currentData(106); xorBitMap(28)(102) := currentData(102); xorBitMap(28)(100) := currentData(100); xorBitMap(28)(99) := currentData(99); xorBitMap(28)(97) := currentData(97); xorBitMap(28)(95) := currentData(95); xorBitMap(28)(94) := currentData(94); xorBitMap(28)(93) := currentData(93); xorBitMap(28)(92) := currentData(92); xorBitMap(28)(91) := currentData(91); xorBitMap(28)(90) := currentData(90); xorBitMap(28)(83) := currentData(83); xorBitMap(28)(81) := currentData(81); xorBitMap(28)(80) := currentData(80); xorBitMap(28)(79) := currentData(79); xorBitMap(28)(78) := currentData(78); xorBitMap(28)(77) := currentData(77); xorBitMap(28)(75) := currentData(75); xorBitMap(28)(69) := currentData(69); xorBitMap(28)(68) := currentData(68); xorBitMap(28)(64) := currentData(64); xorBitMap(28)(63) := currentData(63); xorBitMap(28)(62) := currentData(62); xorBitMap(28)(61) := currentData(61); xorBitMap(28)(59) := currentData(59); xorBitMap(28)(57) := currentData(57); xorBitMap(28)(56) := currentData(56); xorBitMap(28)(54) := currentData(54); xorBitMap(28)(51) := currentData(51); xorBitMap(28)(50) := currentData(50); xorBitMap(28)(49) := currentData(49); xorBitMap(28)(46) := currentData(46); xorBitMap(28)(44) := currentData(44); xorBitMap(28)(43) := currentData(43); xorBitMap(28)(41) := currentData(41); xorBitMap(28)(40) := currentData(40); xorBitMap(28)(33) := currentData(33); xorBitMap(28)(30) := currentData(30); xorBitMap(28)(28) := currentData(28); xorBitMap(28)(27) := currentData(27); xorBitMap(28)(26) := currentData(26); xorBitMap(28)(25) := currentData(25); xorBitMap(28)(24) := currentData(24); xorBitMap(28)(22) := currentData(22); xorBitMap(28)(21) := currentData(21); xorBitMap(28)(20) := currentData(20); xorBitMap(28)(12) := currentData(12); xorBitMap(28)(8) := currentData(8); xorBitMap(28)(6) := currentData(6); xorBitMap(28)(5) := currentData(5); xorBitMap(28)(2) := currentData(2); xorBitMap(28)(161) := previousCrc(1); xorBitMap(28)(163) := previousCrc(3); xorBitMap(28)(164) := previousCrc(4); xorBitMap(28)(166) := previousCrc(6); xorBitMap(28)(170) := previousCrc(10); xorBitMap(28)(171) := previousCrc(11); xorBitMap(28)(173) := previousCrc(13); xorBitMap(28)(174) := previousCrc(14); xorBitMap(28)(176) := previousCrc(16); xorBitMap(28)(177) := previousCrc(17); xorBitMap(28)(178) := previousCrc(18); xorBitMap(28)(179) := previousCrc(19); xorBitMap(28)(183) := previousCrc(23); xorBitMap(28)(185) := previousCrc(25); xorBitMap(28)(186) := previousCrc(26); xorBitMap(28)(187) := previousCrc(27); xorBitMap(28)(188) := previousCrc(28); 
      xorBitMap(29)(125) := currentData(125); xorBitMap(29)(124) := currentData(124); xorBitMap(29)(123) := currentData(123); xorBitMap(29)(122) := currentData(122); xorBitMap(29)(120) := currentData(120); xorBitMap(29)(116) := currentData(116); xorBitMap(29)(115) := currentData(115); xorBitMap(29)(114) := currentData(114); xorBitMap(29)(113) := currentData(113); xorBitMap(29)(111) := currentData(111); xorBitMap(29)(110) := currentData(110); xorBitMap(29)(108) := currentData(108); xorBitMap(29)(107) := currentData(107); xorBitMap(29)(103) := currentData(103); xorBitMap(29)(101) := currentData(101); xorBitMap(29)(100) := currentData(100); xorBitMap(29)(98) := currentData(98); xorBitMap(29)(96) := currentData(96); xorBitMap(29)(95) := currentData(95); xorBitMap(29)(94) := currentData(94); xorBitMap(29)(93) := currentData(93); xorBitMap(29)(92) := currentData(92); xorBitMap(29)(91) := currentData(91); xorBitMap(29)(84) := currentData(84); xorBitMap(29)(82) := currentData(82); xorBitMap(29)(81) := currentData(81); xorBitMap(29)(80) := currentData(80); xorBitMap(29)(79) := currentData(79); xorBitMap(29)(78) := currentData(78); xorBitMap(29)(76) := currentData(76); xorBitMap(29)(70) := currentData(70); xorBitMap(29)(69) := currentData(69); xorBitMap(29)(65) := currentData(65); xorBitMap(29)(64) := currentData(64); xorBitMap(29)(63) := currentData(63); xorBitMap(29)(62) := currentData(62); xorBitMap(29)(60) := currentData(60); xorBitMap(29)(58) := currentData(58); xorBitMap(29)(57) := currentData(57); xorBitMap(29)(55) := currentData(55); xorBitMap(29)(52) := currentData(52); xorBitMap(29)(51) := currentData(51); xorBitMap(29)(50) := currentData(50); xorBitMap(29)(47) := currentData(47); xorBitMap(29)(45) := currentData(45); xorBitMap(29)(44) := currentData(44); xorBitMap(29)(42) := currentData(42); xorBitMap(29)(41) := currentData(41); xorBitMap(29)(34) := currentData(34); xorBitMap(29)(31) := currentData(31); xorBitMap(29)(29) := currentData(29); xorBitMap(29)(28) := currentData(28); xorBitMap(29)(27) := currentData(27); xorBitMap(29)(26) := currentData(26); xorBitMap(29)(25) := currentData(25); xorBitMap(29)(23) := currentData(23); xorBitMap(29)(22) := currentData(22); xorBitMap(29)(21) := currentData(21); xorBitMap(29)(13) := currentData(13); xorBitMap(29)(9) := currentData(9); xorBitMap(29)(7) := currentData(7); xorBitMap(29)(6) := currentData(6); xorBitMap(29)(3) := currentData(3); xorBitMap(29)(160) := previousCrc(0); xorBitMap(29)(162) := previousCrc(2); xorBitMap(29)(164) := previousCrc(4); xorBitMap(29)(165) := previousCrc(5); xorBitMap(29)(167) := previousCrc(7); xorBitMap(29)(171) := previousCrc(11); xorBitMap(29)(172) := previousCrc(12); xorBitMap(29)(174) := previousCrc(14); xorBitMap(29)(175) := previousCrc(15); xorBitMap(29)(177) := previousCrc(17); xorBitMap(29)(178) := previousCrc(18); xorBitMap(29)(179) := previousCrc(19); xorBitMap(29)(180) := previousCrc(20); xorBitMap(29)(184) := previousCrc(24); xorBitMap(29)(186) := previousCrc(26); xorBitMap(29)(187) := previousCrc(27); xorBitMap(29)(188) := previousCrc(28); xorBitMap(29)(189) := previousCrc(29); 
      xorBitMap(30)(126) := currentData(126); xorBitMap(30)(125) := currentData(125); xorBitMap(30)(124) := currentData(124); xorBitMap(30)(123) := currentData(123); xorBitMap(30)(121) := currentData(121); xorBitMap(30)(117) := currentData(117); xorBitMap(30)(116) := currentData(116); xorBitMap(30)(115) := currentData(115); xorBitMap(30)(114) := currentData(114); xorBitMap(30)(112) := currentData(112); xorBitMap(30)(111) := currentData(111); xorBitMap(30)(109) := currentData(109); xorBitMap(30)(108) := currentData(108); xorBitMap(30)(104) := currentData(104); xorBitMap(30)(102) := currentData(102); xorBitMap(30)(101) := currentData(101); xorBitMap(30)(99) := currentData(99); xorBitMap(30)(97) := currentData(97); xorBitMap(30)(96) := currentData(96); xorBitMap(30)(95) := currentData(95); xorBitMap(30)(94) := currentData(94); xorBitMap(30)(93) := currentData(93); xorBitMap(30)(92) := currentData(92); xorBitMap(30)(85) := currentData(85); xorBitMap(30)(83) := currentData(83); xorBitMap(30)(82) := currentData(82); xorBitMap(30)(81) := currentData(81); xorBitMap(30)(80) := currentData(80); xorBitMap(30)(79) := currentData(79); xorBitMap(30)(77) := currentData(77); xorBitMap(30)(71) := currentData(71); xorBitMap(30)(70) := currentData(70); xorBitMap(30)(66) := currentData(66); xorBitMap(30)(65) := currentData(65); xorBitMap(30)(64) := currentData(64); xorBitMap(30)(63) := currentData(63); xorBitMap(30)(61) := currentData(61); xorBitMap(30)(59) := currentData(59); xorBitMap(30)(58) := currentData(58); xorBitMap(30)(56) := currentData(56); xorBitMap(30)(53) := currentData(53); xorBitMap(30)(52) := currentData(52); xorBitMap(30)(51) := currentData(51); xorBitMap(30)(48) := currentData(48); xorBitMap(30)(46) := currentData(46); xorBitMap(30)(45) := currentData(45); xorBitMap(30)(43) := currentData(43); xorBitMap(30)(42) := currentData(42); xorBitMap(30)(35) := currentData(35); xorBitMap(30)(32) := currentData(32); xorBitMap(30)(30) := currentData(30); xorBitMap(30)(29) := currentData(29); xorBitMap(30)(28) := currentData(28); xorBitMap(30)(27) := currentData(27); xorBitMap(30)(26) := currentData(26); xorBitMap(30)(24) := currentData(24); xorBitMap(30)(23) := currentData(23); xorBitMap(30)(22) := currentData(22); xorBitMap(30)(14) := currentData(14); xorBitMap(30)(10) := currentData(10); xorBitMap(30)(8) := currentData(8); xorBitMap(30)(7) := currentData(7); xorBitMap(30)(4) := currentData(4); xorBitMap(30)(160) := previousCrc(0); xorBitMap(30)(161) := previousCrc(1); xorBitMap(30)(163) := previousCrc(3); xorBitMap(30)(165) := previousCrc(5); xorBitMap(30)(166) := previousCrc(6); xorBitMap(30)(168) := previousCrc(8); xorBitMap(30)(172) := previousCrc(12); xorBitMap(30)(173) := previousCrc(13); xorBitMap(30)(175) := previousCrc(15); xorBitMap(30)(176) := previousCrc(16); xorBitMap(30)(178) := previousCrc(18); xorBitMap(30)(179) := previousCrc(19); xorBitMap(30)(180) := previousCrc(20); xorBitMap(30)(181) := previousCrc(21); xorBitMap(30)(185) := previousCrc(25); xorBitMap(30)(187) := previousCrc(27); xorBitMap(30)(188) := previousCrc(28); xorBitMap(30)(189) := previousCrc(29); xorBitMap(30)(190) := previousCrc(30); 
      xorBitMap(31)(127) := currentData(127); xorBitMap(31)(126) := currentData(126); xorBitMap(31)(125) := currentData(125); xorBitMap(31)(124) := currentData(124); xorBitMap(31)(122) := currentData(122); xorBitMap(31)(118) := currentData(118); xorBitMap(31)(117) := currentData(117); xorBitMap(31)(116) := currentData(116); xorBitMap(31)(115) := currentData(115); xorBitMap(31)(113) := currentData(113); xorBitMap(31)(112) := currentData(112); xorBitMap(31)(110) := currentData(110); xorBitMap(31)(109) := currentData(109); xorBitMap(31)(105) := currentData(105); xorBitMap(31)(103) := currentData(103); xorBitMap(31)(102) := currentData(102); xorBitMap(31)(100) := currentData(100); xorBitMap(31)(98) := currentData(98); xorBitMap(31)(97) := currentData(97); xorBitMap(31)(96) := currentData(96); xorBitMap(31)(95) := currentData(95); xorBitMap(31)(94) := currentData(94); xorBitMap(31)(93) := currentData(93); xorBitMap(31)(86) := currentData(86); xorBitMap(31)(84) := currentData(84); xorBitMap(31)(83) := currentData(83); xorBitMap(31)(82) := currentData(82); xorBitMap(31)(81) := currentData(81); xorBitMap(31)(80) := currentData(80); xorBitMap(31)(78) := currentData(78); xorBitMap(31)(72) := currentData(72); xorBitMap(31)(71) := currentData(71); xorBitMap(31)(67) := currentData(67); xorBitMap(31)(66) := currentData(66); xorBitMap(31)(65) := currentData(65); xorBitMap(31)(64) := currentData(64); xorBitMap(31)(62) := currentData(62); xorBitMap(31)(60) := currentData(60); xorBitMap(31)(59) := currentData(59); xorBitMap(31)(57) := currentData(57); xorBitMap(31)(54) := currentData(54); xorBitMap(31)(53) := currentData(53); xorBitMap(31)(52) := currentData(52); xorBitMap(31)(49) := currentData(49); xorBitMap(31)(47) := currentData(47); xorBitMap(31)(46) := currentData(46); xorBitMap(31)(44) := currentData(44); xorBitMap(31)(43) := currentData(43); xorBitMap(31)(36) := currentData(36); xorBitMap(31)(33) := currentData(33); xorBitMap(31)(31) := currentData(31); xorBitMap(31)(30) := currentData(30); xorBitMap(31)(29) := currentData(29); xorBitMap(31)(28) := currentData(28); xorBitMap(31)(27) := currentData(27); xorBitMap(31)(25) := currentData(25); xorBitMap(31)(24) := currentData(24); xorBitMap(31)(23) := currentData(23); xorBitMap(31)(15) := currentData(15); xorBitMap(31)(11) := currentData(11); xorBitMap(31)(9) := currentData(9); xorBitMap(31)(8) := currentData(8); xorBitMap(31)(5) := currentData(5); xorBitMap(31)(160) := previousCrc(0); xorBitMap(31)(161) := previousCrc(1); xorBitMap(31)(162) := previousCrc(2); xorBitMap(31)(164) := previousCrc(4); xorBitMap(31)(166) := previousCrc(6); xorBitMap(31)(167) := previousCrc(7); xorBitMap(31)(169) := previousCrc(9); xorBitMap(31)(173) := previousCrc(13); xorBitMap(31)(174) := previousCrc(14); xorBitMap(31)(176) := previousCrc(16); xorBitMap(31)(177) := previousCrc(17); xorBitMap(31)(179) := previousCrc(19); xorBitMap(31)(180) := previousCrc(20); xorBitMap(31)(181) := previousCrc(21); xorBitMap(31)(182) := previousCrc(22); xorBitMap(31)(186) := previousCrc(26); xorBitMap(31)(188) := previousCrc(28); xorBitMap(31)(189) := previousCrc(29); xorBitMap(31)(190) := previousCrc(30); xorBitMap(31)(191) := previousCrc(31); 
   end procedure;

end package body EthCrc32Pkg;

