`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
qWIj44uDTKWTZ+1mHcC9GhHtznfXek6+SThg9ej3m7L/Lc/XyHOIQvWEsASy+eJtF24bXBkTA04U
4aubic3PYA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FuHJ2twPEmSQBC5MXoX/q8+spKC4AYXcmGeCfyN3AribUkV3QF0QxpZ/gnmpm8HCvq6wWX4u9Ozf
PC+a8cwNwYkYHBVjw8m2vRVJsxeaTB4Hgwcut4afp959aT0OfuN5FzSNC/xk9bIMDNJrCHMGe1LU
mIh49gA8oUT0QfCnrq8=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
bA3lomTKIBe9pwigCbapcDGETp1XXuOxxiukByJ3JYOGFmb5qJakTizx2sh+MaxJADkn7K1+M9Zo
QSxqSOHgDdn9Yatx9rhFZaVnqSk8zCFurjxL3xa7FkrfQrF9FdC7+1iZq1tajS1eMmlZZId4nxlg
Z28O/YLbPbfWCL32nzE=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ND8eM+xO5f4CH7mpptPfhVOilvME/9UDwNiI+515S2DlbAGsnIgvwtc+ueUEeT1Gip2yjqJAtQy5
hsu76DWErskRP/FiMCOun3uZ4pJWLpuBL3lsk9f7/13Wa2nXMT6qEi5VbRgwgA/7hVTUY80vmhTu
hjcB9hNPJMIoMSImlOczIoIO4FEY3SW+FO9+Rw2dAO+Vtonx73vBhPmugNwHCK5LwOxoJjM0dUCt
MuI/090uYu8cZUhZUBJaE3mSuSE8yMJgsKUPmJLLomUbXWOAghJo/6LZsFqre4gernB/uCl07+W7
n1X8VmJ7kd5bTkCRg6kWVO0ITpq9M29/gDeTHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Q0w9iswld7AxcoW0jbqdJQ0MImkqs8w6MEWcx1Hlwsw2ItrPDzgY69grM5qiTgARbaw5pMBlD5pA
dWLMdg9BWvbTAIIJSK/sg+TR84f9DLhy0Le7ie1+kX9WermOdFZf+mEHKetxG7hftFD4gF1ehux9
ikeGpBLLx4mo8OSmuXT8MV0Ib8A1zcpdUU3lBcU0GHZhtNw32PicrkC0UiHpxn2zj2X8XPYZux8D
9BnhBIjeBcskMbCaPQGeizx9iMEz6Esebm50BImuhN50jetTLRj6bech2vNUYzFuUapR97m6kuLA
BZZaJIJ6j6J27dyWAfIxkpJIGBemZrClfZ/o6w==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
PKkRlaOjodauNK8Etola960WD57dmghcTLLZFk7vLULnB7/rzJbwk1yC5ldSlLVQcGknezziOZ4x
ACO1Af7uQl9DWpR76WlEODfURaDDn/ZzrK/2UNB27nZSfbrkSzF1itCxobccRkILSY5TnEg6K5We
9FAebFO3228lher3DRpq2OhSfNk3yoAXs6ooliqz0v+sSJ+cyGGJG1sWGw14h8Zt6X4Ydsx7PI3z
tWDxi6VcjrmIIXG/HgM3uJtEE6sq2kzwm0EaqPR5F3kA5IPmluVRJUbwvgxQdGN959VHIAV4vpD3
75ny3D6Warg6soJMTEKy6hb/h5opq7Sxq6mrng==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
5QCMP/bv5Wdr4VeA8vX2bYweg7B3xLxU6PN7Jaq8NjJOmXkh+0ZFCVro/WlXot2RdoO1lK6eQzVE
8gMHgDW5p0vAvMKgBIGdBeqBF9d9kCHDAjE1kCxEGu5Z5g/sW2/jCMy7JqV70iUxVb2mh3qjCF2O
tLfIWOd5xbIrajtUQnW2Ko+MvIlztdgT27gBm7R35/IzqrUieQmF7oNBchKvG9Q4bx2Idh9ihL55
K7KY8jAEwGIJNlYVkILrXFehRusezC0kCRVsWztOaJl3LdyfxTiG9LzEPorJWSzb9caeQjsKgL66
y/X4Itfz6Lcgztwlk+asXdw05D4ygUN+Ga+vl/NclVNXf9DBxcQHxTnEoJwYAhOnQnL8hbEusS8v
jKzKoM4QluB/Q/sbFmQxgNK4rUALiJMABz6KUHKF/1oQFyMCuAGFAJv6gexVUtwg8zjkXKf9WzMT
fq4PuAYudNoZ4ghISGQi7UcxLlekW+S/JnUqjl0UL3VFXCETIqR1ivXKyzUMJWmAUKMsQuDaa43S
DVrw+mjmAfOBiJ+R+55qE5N8Ng96Gdh/lQ0JXWgSCEX9oHJuWcttuViSI4cKoTZjnasXJQuZhTP+
ftmqX2zjut1J8Y7go130PraiKyJWBq23fYJFS06Nh1nK3gzEaBmSSnNu2opTfHvm6NgOUs9Jwvu6
QXfuDdU0oFDCFWBtvwezhmX8ke0DJEbS0nAphcXDBHLXzBuj8k6Bp3Pwa5L8Tbb0SI6Dz7ccScv3
bG7BLbsg3ffUvFf3wXEH2xL34sQtOyeYp8XLljGPZNVgFScVfptENh74S2zCCgKK/BOq1HJU6OmG
pJZcOumFLlmkxUSLnkOBFuDYvKzpTaHWtufNaANJ5z/n/yhTFP2EOKFbdoFcBIdlDv+w+iRwFzya
hljA5mKchNyhTwzklvLWveM/mUmv8X3flbIyo8KeS+Q1IwOVesxyJyE0P9+LPPvpjNPH5gJAIGyz
Zo0LoJ2EOdOP5pjJ2LbEFbKmU2oxGGZaCLDhdLfZR5n0KQ2H/z689MXoghfUVtYMFNqrDxLm9s9G
V76JcQ4vkFyiDoGNBcemz0sRkuedQWErKESMt1wBZ8m4RQbqL8f2kimQgrFJ8+03zTymAJPQFKir
y2Fnw5dtxr7SCwzNZpDb+y0ZjreAi0q8jb5f4fAck7cIU/8I2ox1d0SqQfSCBPjIAO5+Y0u3sT2W
Nc6KYvnAyDVvW8aeZMA+5FDgVLHMJU7Y8PHZPxSNm67wuIMiBzPe7yqHQntZ8ONRzxeQOhs72har
bebo2JeDJs7w1duyzW2+1DXLy0SR21FhjXWINgp0EMVk/vcCIJO8sQEy3U1A9JOmfh6E/L2B9Ys0
h+A3mA+c/+xTBhu7wX9bFmCg6yUWyoUaR1RDInD48+atecQ/u/cBjLSbXQKKrpmO3npYfGYDqj5G
gqw0wLw7aXVRWkW4ecI5LHguEZIXfsDpq8qerVk/DIVwh8S//ELVCvxXrnZQK92cejU8VXXZAABf
ZU2dx6B36ubm+4mp4yoQn3d+uhArS6ncUPwZtN1F54QXiiwjqluWKzLAruM7UGhQ1sCTvzR5nNw0
nOGmYlPpMUMvPUDov2+P48s9f29Ompj5uI0L/ZT5KKgidejJoUPbasrSIXSnbRNbZG2jJkUnAwp0
TxSsjlP0B1u/AnSZjHlJPjslif9vNzsMTzaB1o8DSGq9zXIr+ElPvcFG5vp/N1/TlK6sOfl7g19Y
e25FBZXbBY2NjcK5snwtN7K3B6naBYHuYCegPEQZExNCiQ4dfSj+WEX933KcL1km0e3edteznkek
tPeAWb9JTFI/9/nUKG3aytPrdLpsTk9djFqhZdv49iYr7KA+IOS5ZCOOLx5Xszs7jWPmT4dGrPv5
wW1pcJGDYt2puo2pj0JedEy6Orp48xnnHk4wHm65kht7NC5G8JEI1J9CUh5PF4DlzyhR2mB+8obY
QxZwcew3OZN/C9HzlhV0cKTpzhkPInjI8U+tSVknPMkLE5C8gSyhPNreGqd3q2pA/Q6ZpHOijND5
fqBuYMvWiTEviRkkMsh7xjej746Ha06eqpXdDQadY+S3pkzn4PBq8tz735tqcqR0uwxxzpq3sfs4
w8HIwaLXR4Loe5I8I3uAEQ9BP07ae1xwQNOjXPO3IbV59CSSICld1AUTYsl6E6QApmH6GxP9r9V1
dKIwiUutA55wmbRs4/nZC2Rc7UN6+UvowdIH0ao1WEdh9VNg1Ae0Xlkd2rW06+ecYzYXdY+9KNjY
APSb5hdI+u4PJQc3Sh1zvT3CS02AeNbvAyO+jlf2hu6bqH1ld5akFGoTBibU6tyxG6haiEQdY263
rDKh+rikBqLpQFnZf0UO6xVInqmpLLoZ5I2Z2ve6F88vqvzGfVw1fTNpq8GbQOxrEyBeLL/vBra0
5bjvhx8ZRZwY3STyS/uTxGnkaqElXNLwK51SdxlprcDLLiVdztZ0DhLyuQnPReKmnspY2f9C704C
MMsE/p+iAss9IIU7fTR5+EaPmfYmhfeSJxsEWlUUFd7KVMaM8wLbLzsEviKCEJNl85v1mNGUT4Pn
mKeGOSnMBNM47azLWE14VIwvTDKVGo3SHvZCZz8lMY08GGkFl3QTNlbx6zA0fuaeiIcaWScCgKfr
Q4gOJSQiEmkiLGxtI0oUBWMRjv6R6YD39p16j/BB7ouNGfeU6+RmMSG+hwrMcoIU8KJOsoiN3Vpw
qfAuzM4/hyUVGnn0fQMFEyMCTuk0CgDEVelCbnRVxRn3V23ncSvkkauNmLc3S/kFxUcK/R6BWZqK
Uy5afNV8lhOo2lY5moetAhFg6UzQNDId+jsfWdj8O46WrpK0LsEnFxE7N/QJhkV/lRC07J4esE4s
W/fw3r/jO19c9zNWVjENjwWtqEWwc3UqejZS0xfcjEK/U605Hkt6YjvUcwImYS9nK2ik3cRVcZWj
OGd7hBFxhHTyjhgMJHEFmszbxhGAf8G2kQQ3n/jzXnAvnlOdwGBmouPFTkXp7z3NHXqrpn+4xHhN
peDyxPIYbGKvHVHjEqt4TU4vJ9kWkhFryXoDQ3vO77MqhYJ/ky4sSfGgDO7m1Zz8e31hTl/4BFqq
9zbp/kH5sdYoGsDnex52Stx7Rn8jIVreNeuEPhx8Kg1AHa/SQSbkRFR6eRT5aWwNgIy3S6SvL6Js
d+BukM4/Z/UbSw5JYW4uVY6tI38EpqfDBy1Ln2nNXoHnfErlncCGuDXy4HrPZ3DRVMDpNWyrtOdT
z8/BQbaagPngeyE8B2cwe2GXkIh8jORzP7Q3MmnfivqIqAGiMGzb8wNCAyAsomiiLAW69MFfX9x5
u9hxoJ2YFIWPwq9TraKvATlCFkaPTdCZd/jS+hIwdPvZqH8WvaQ4/kSzLPW7SJj1dYpnOTYWOiSx
znM6pig40f8eXtXkomFdq+j1uJW11chG6hXodMcRDqnfcpQkJyLtwuyF/95TEutSR/gvrKIuY/Rp
NziGRkMbyVtjJYyPfyLdHGDANVIrnpqGSdIAb9SyQlP3CvwCyaTViqa4u9X/zkgO6rznSWv1OvAU
3Ogkt89B9FczszpMXgPWAy2u65/KIgcPp3SWi5VUYac4L1aAhU3NVKzvr93g1haIBUitk0+rU2bg
HwSKP8H/MyOhLBbx7OiqRo+gUUNXmpVAvTcRfLzgDFnxWdN8h+197tbXRJgsts6ogiVlB6jPXtPU
MkJI3METxJyz4vfrGOar0teOozgf10CCVubrSrebiyn880446Dnm3TKJ00vfP3gS9A1wSiG0stfl
I8AeVlK5Em5F+svadRTkKJfInPhANpQ2YoRB/Mw9joWw6jHSSenpFM3KQk/4ECWhnFLrhnWIVwHz
jzwfA19NAJKVOxNA3kVVFPvw7VcYq/HFZxXFzgdLBMyMsVstsWENxAQASrX3QUBCDI3UlC1dYBZe
DTQv5W09TmkfNhjXk1oa3AL8mFGr6fqWxXlZND6sAv/X2FoNQs0d3ChFgM20hAMVFqEFpljn8QhE
uI3q15xj0C7dmQ6RzCid2tWa6PnBe9yp8hCogvp4flVZ/D4sbHMSY+re0XVcMw2biKazne5UryQv
Uv+6zdrYifgzyojc6oPrzhOHJl6huZIzfUq3bwPJAmT2hnszP1v0ZnLv/RkFtGyGcO+NSV1eWR0l
TA==
`pragma protect end_protected
