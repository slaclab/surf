-------------------------------------------------------------------------------
-- Title      : 
-------------------------------------------------------------------------------
-- File       : i2cRegMasterSimPkg.vhd
-- Author     : Benjamin Reese  <bareese@slac.stanford.edu>
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2013-01-24
-- Last update: 2013-01-25
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2013 SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.StdRtlPkg.all;
use work.i2cPkg.all;
use work.txt_util_p.all;

package i2cRegMasterPkg is

  procedure writeI2cReg (
    signal clk    : in  sl;
    signal regIn  : out i2cRegMasterInType;
    signal regOut : in  i2cRegMasterOutType;
    i2cAddr       : in  slv;
    regAddr       : in  slv;
    regData       : in  slv;
    endianness    : in  sl;
    debug : in boolean := false);

  procedure readI2cReg (
    signal clk    : in  sl;
    signal regIn  : out i2cRegMasterInType;
    signal regOut : in  i2cRegMasterOutType;
    i2cAddr       : in  slv;
    regAddr       : in  slv;
    regData       : out slv;
    endianness    : in  sl;
    debug : in boolean := false);

end package i2cRegMasterPkg;

package body i2cRegMasterPkg is

  procedure writeI2cReg (
    signal clk    : in  sl;
    signal regIn  : out i2cRegMasterInType;
    signal regOut : in  i2cRegMasterOutType;
    i2cAddr       : in  slv;
    regAddr       : in  slv;
    regData       : in  slv;
    endianness    : in  sl;
    debug : in boolean := false)
  is
    variable i2cAddrSizeVar : integer := i2cAddr'length;
    variable regAddrSizeVar : integer := regAddr'length/8;
    variable regDataSizeVar : integer := regData'length/8;
  begin
    wait until clk = '1';
    
    -- Put write on inputs
    if (i2cAddrSizeVar = 7) then
      regIn.i2cAddr <= "000" & i2cAddr;
      regIn.tenbit  <= '0';
    elsif (i2cAddrSizeVar = 10) then
      regIn.i2cAddr <= i2cAddr;
      regIn.tenbit  <= '1';
    end if;
    regIn.regAddr                <= (others => '0');
    regIn.regAddr(regAddr'range) <= regAddr;
    regIn.regAddrSize            <= slv(to_unsigned(regAddrSizeVar-1, 2));
    regIn.regDataSize            <= slv(to_unsigned(regDataSizeVar-1, 2));
    regIn.endianness             <= endianness;
    regIn.regOp                  <= '1';

    regIn.regWrData                <= (others => '0');
    regIn.regWrData(regData'range) <= regData;

    regIn.regReq <= '1';

    -- Wait for ack
    wait until regOut.regAck = '1';
    wait until clk = '1';
    regIn.regReq <= '0';
    wait until regOut.regAck = '0';
    wait until clk = '1';

    print(debug, "writeI2cReg: i2c: " & str(i2cAddr) & ", addr: " & hstr(regAddr) & ", data: " & hstr(regData));

  end procedure writeI2cReg;

  procedure readI2cReg (
    signal clk    : in  sl;
    signal regIn  : out i2cRegMasterInType;
    signal regOut : in  i2cRegMasterOutType;
    i2cAddr       : in  slv;
    regAddr       : in  slv;
    regData       : out slv;
    endianness    : in  sl;
    debug : in boolean := false)
  is
    variable i2cAddrSizeVar : integer := i2cAddr'length;
    variable regAddrSizeVar : integer := regAddr'length/8;
    variable regDataSizeVar : integer := regData'length/8;
  begin
    wait until clk = '1';
        
    if (i2cAddrSizeVar = 7) then
      regIn.i2cAddr <= "000" & i2cAddr;
      regIn.tenbit  <= '0';
    elsif (i2cAddrSizeVar = 10) then
      regIn.i2cAddr <= i2cAddr;
      regIn.tenbit  <= '1';
    end if;
    regIn.regAddr                <= (others => '0');
    regIn.regAddr(regAddr'range) <= regAddr;
    regIn.regAddrSize            <= slv(to_unsigned(regAddrSizeVar-1, 2));
    regIn.regDataSize            <= slv(to_unsigned(regDataSizeVar-1, 2));
    regIn.endianness             <= endianness;
    regIn.regOp                  <= '0';

    regIn.regReq <= '1';

    wait until regOut.regAck = '1';
    wait until clk = '1';
    regIn.regReq <= '0';
   
    regData := regOut.regRdData(regData'range);
    wait until regOut.regAck = '0';
    wait until clk = '1';

    print(debug, "readI2cReg: i2c: " & str(i2cAddr) & ", addr: " & hstr(regAddr) & " Data: " & hstr(regOut.regRdData(regData'range)));
    
  end procedure readI2cReg;

end package body i2cRegMasterPkg;
