-------------------------------------------------------------------------------
-- Title      : GLink Decoder
-------------------------------------------------------------------------------
-- File       : GlinkDecoder.vhd
-- Author     : Benjamin Reese  <bareese@slac.stanford.edu>
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2012-03-12
-- Last update: 2014-04-17
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: Decoder for the Condition Inversion Master Transition coding
-- used by the GLink Protocol.
-------------------------------------------------------------------------------
-- Copyright (c) 2014 SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.StdRtlPkg.all;
use work.GlinkPkg.all;

entity GLinkDecoder is
   generic (
      TPD_G          : time    := 1 ns;
      RST_ASYNC_G    : boolean := false;
      RST_POLARITY_G : sl      := '1';  -- '1' for active HIGH reset, '0' for active LOW reset      
      FLAGSEL_G      : boolean := false);
   port (
      en            : in  sl := '1';
      clk           : in  sl;
      rst           : in  sl;
      gtRxData      : in  slv(19 downto 0);
      rxReady       : in  sl;
      txReady       : in  sl;           -- TX Clock domain
      gLinkRx       : out GLinkRxType;
      decoderError  : out sl;
      decoderErrorL : out sl);  
end entity GLinkDecoder;

architecture rtl of GLinkDecoder is

   type RegType is record
      toggle  : sl;
      gLinkRx : GLinkRxType;
   end record;
   
   constant REG_INIT_C : RegType := (
      '0',
      GLINK_RX_INIT_C);      

   signal r   : RegType := REG_INIT_C;
   signal rin : RegType;

   signal txRdy : sl;
   
begin

   Synchronizer_Inst : entity work.Synchronizer
      generic map (
         TPD_G          => TPD_G,
         RST_ASYNC_G    => RST_ASYNC_G,
         RST_POLARITY_G => RST_POLARITY_G)
      port map (
         clk     => clk,
         rst     => rst,
         dataIn  => txReady,
         dataOut => txRdy);

   comb : process (gtRxData, r, rst, rxReady, txRdy) is
      variable v            : RegType;
      variable glinkWordVar : GLinkWordType;
   begin
      v := r;

      -- Update the TX and RX MGT ready values
      v.gLinkRx.rxReady := rxReady;
      v.gLinkRx.txReady := txRdy;

      -- Reset strobe signals
      v.gLinkRx.error     := '0';
      v.gLinkRx.isControl := '0';
      v.gLinkRx.isIdle    := '1';
      v.gLinkRx.isData    := '0';
      v.gLinkRx.flag      := '0';

      -- Convert input to GLinkWordType to use GLinkPkg functions for decoding
      glinkWordVar := toGLinkWord(gtRxData);

      if (not isValidWord(glinkWordVar)) then
         -- Invalid input, don't decode
         v.gLinkRx.error := '1';
      else
         -- Valid input, decode the input
         -- Check for control word
         if (isControlWord(glinkWordVar)) then
            -- Check for idle word (subcase of control word)
            if (not isIdleWord(glinkWordVar)) then
               v.gLinkRx.isIdle    := '0';
               v.gLinkRx.isControl := '1';
               v.gLinkRx.data      := getControlPayload(glinkWordVar);
            end if;
         end if;

         -- Check for data word
         if (isDataWord(glinkWordVar)) then
            if FLAGSEL_G then
               v.gLinkRx.isIdle := '0';
               v.gLinkRx.isData := '1';
               v.gLinkRx.data   := getDataPayload(gLinkWordVar);        -- Bit flip done by function
               v.gLinkRx.flag   := getFlag(gLinkWordVar);
            else
               -- Check for first data frame
               if r.gLinkRx.linkUp = '0' then
                  -- First frame Detected
                  v.gLinkRx.linkUp := '1';
                  -- Set the gLinkRx bus
                  v.gLinkRx.isIdle := '0';
                  v.gLinkRx.isData := '1';
                  v.gLinkRx.data   := getDataPayload(gLinkWordVar);     -- Bit flip done by function
                  v.gLinkRx.flag   := getFlag(gLinkWordVar);
                  -- Latch the flag value
                  v.toggle         := getFlag(gLinkWordVar);
               else
                  -- Check for flag error
                  if (r.toggle = getFlag(gLinkWordVar)) then
                     -- Invalid flag detected
                     v.gLinkRx.error := '1';
                  else
                     -- Set the gLinkRx bus
                     v.gLinkRx.isIdle := '0';
                     v.gLinkRx.isData := '1';
                     v.gLinkRx.data   := getDataPayload(gLinkWordVar);  -- Bit flip done by function
                     v.gLinkRx.flag   := getFlag(gLinkWordVar);
                     -- Latch the flag value
                     v.toggle         := getFlag(gLinkWordVar);
                  end if;
               end if;
            end if;
         end if;

         -- Invert if necessary
         if (isInvertedWord(glinkWordVar)) then
            v.gLinkRx.data := not v.gLinkRx.data;
         end if;
      end if;

      -- Synchronous Reset
      if (RST_ASYNC_G = false and rst = RST_POLARITY_G) then
         v := REG_INIT_C;
      end if;

      -- Register the variable for next clock cycle
      rin <= v;

      -- Outputs      
      gLinkRx       <= r.gLinkRx;
      decoderError  <= r.gLinkRx.error;
      decoderErrorL <= not(r.gLinkRx.error);
      
   end process comb;

   seq : process (clk, rst) is
   begin
      if rising_edge(clk) then
         if en = '1' then
            r <= rin after TPD_G;
         end if;
      end if;
      -- Asynchronous Reset
      if (RST_ASYNC_G and rst = RST_POLARITY_G) then
         r <= REG_INIT_C after TPD_G;
      end if;
   end process seq;

end architecture rtl;
