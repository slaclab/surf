-------------------------------------------------------------------------------
-- Title      : PGPv3: https://confluence.slac.stanford.edu/x/OndODQ
-------------------------------------------------------------------------------
-- Company    : SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------
-- Description: PGP3 GTY Ultrascale+ QPLL Wrapper
-------------------------------------------------------------------------------
-- This file is part of 'SLAC Firmware Standard Library'.
-- It is subject to the license terms in the LICENSE.txt file found in the
-- top-level directory of this distribution and at:
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html.
-- No part of 'SLAC Firmware Standard Library', including this file,
-- may be copied, modified, propagated, or distributed except according to
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library surf;
use surf.StdRtlPkg.all;
use surf.AxiLitePkg.all;

library unisim;
use unisim.vcomponents.all;

entity Pgp3GtyUsQpll is
   generic (
      TPD_G             : time            := 1 ns;
      RATE_G            : string          := "10.3125Gbps";
      QPLL_REFCLK_SEL_G : slv(2 downto 0) := "001";
      EN_DRP_G          : boolean         := true);
   port (
      -- Stable Clock and Reset
      stableClk       : in  sl;         -- GT needs a stable clock to "boot up"
      stableRst       : in  sl;
      -- QPLL Clocking
      pgpRefClk       : in  sl;         -- 156.25 MHz
      qpllLock        : out Slv2Array(3 downto 0);
      qpllClk         : out Slv2Array(3 downto 0);
      qpllRefclk      : out Slv2Array(3 downto 0);
      qpllRst         : in  Slv2Array(3 downto 0);
      -- AXI-Lite Interface
      axilClk         : in  sl                     := '0';
      axilRst         : in  sl                     := '0';
      axilReadMaster  : in  AxiLiteReadMasterType  := AXI_LITE_READ_MASTER_INIT_C;
      axilReadSlave   : out AxiLiteReadSlaveType   := AXI_LITE_READ_SLAVE_EMPTY_DECERR_C;
      axilWriteMaster : in  AxiLiteWriteMasterType := AXI_LITE_WRITE_MASTER_INIT_C;
      axilWriteSlave  : out AxiLiteWriteSlaveType  := AXI_LITE_WRITE_SLAVE_EMPTY_DECERR_C);
end Pgp3GtyUsQpll;

architecture mapping of Pgp3GtyUsQpll is

   constant QPLL_PPF0_CFG_C : slv(15 downto 0) := ite((RATE_G = "13.75Gbps"), b"0000100100000000", b"0000011000000000");
   constant QPLL_PPF1_CFG_C : slv(15 downto 0) :=
      ite((RATE_G = "20.625Gbps"), b"0000011000000000",
          ite((RATE_G = "25.0Gbps"), b"0000100000000000",
              b"0000010000000000"));

   constant QPLL_CFG2_C : slv(15 downto 0) :=
      ite((RATE_G = "10.3125Gbps") or (RATE_G = "25.0Gbps"), b"0000111111000000",
          ite((RATE_G = "15.46875Gbps"), b"0000111111000001",
              b"0000111111000011"));

   constant QPLL_CFG4_C : slv(15 downto 0) :=
      ite((RATE_G = "17.1875Gbps") or (RATE_G = "18.75Gbps") or (RATE_G = "20.625Gbps"), b"0000000000000011",
          ite((RATE_G = "25.0Gbps"), b"0000000010000100",
              b"0000000000000010"));

   constant QPLL_CP_G3_C : slv(9 downto 0) := ite((RATE_G = "3.125Gbps") or (RATE_G = "17.1875Gbps") or (RATE_G = "18.75Gbps") or (RATE_G = "20.625Gbps") or (RATE_G = "25.0Gbps"), b"0001111111", b"0000001111");

   constant QPLL_FBDIV_C : positive :=
      ite((RATE_G = "6.25Gbps") or (RATE_G = "12.5Gbps") or (RATE_G = "25.0Gbps"), 80,
          ite((RATE_G = "13.75Gbps"), 88,
              ite((RATE_G = "15.46875Gbps"), 99,
                  ite((RATE_G = "17.1875Gbps"), 55,
                      ite((RATE_G = "18.75Gbps"), 60,
                          66)))));

   constant QPLL_FBDIV_G3_C : positive := ite((RATE_G = "3.125Gbps") or (RATE_G = "17.1875Gbps") or (RATE_G = "18.75Gbps") or (RATE_G = "20.625Gbps") or (RATE_G = "25.0Gbps"), 80, 160);

   constant QPLL_LPF_C : slv(9 downto 0) :=
      ite((RATE_G = "10.3125Gbps"), b"1000111111",
          ite((RATE_G = "15.46875Gbps"), b"1101111111",
              ite((RATE_G = "25.0Gbps"), b"1100111111",
                  b"1000011111")));

   constant QPLL_LPF_G3_C : slv(9 downto 0) := ite((RATE_G = "3.125Gbps") or (RATE_G = "17.1875Gbps") or (RATE_G = "18.75Gbps") or (RATE_G = "20.625Gbps") or (RATE_G = "25.0Gbps"), b"0111010100", b"0111010101");

   signal pllRefClk     : slv(1 downto 0);
   signal pllOutClk     : slv(1 downto 0);
   signal pllOutRefClk  : slv(1 downto 0);
   signal pllFbClkLost  : slv(1 downto 0);  -- unused
   signal pllLock       : slv(1 downto 0);
   signal pllLockDetClk : slv(1 downto 0);
   signal pllRefClkLost : slv(1 downto 0);
   signal pllPowerDown  : slv(1 downto 0);
   signal pllReset      : slv(1 downto 0);
   signal lockedStrobe  : Slv2Array(3 downto 0);
   signal gtQPllReset   : Slv2Array(3 downto 0);

begin

   assert ((RATE_G = "3.125Gbps") or (RATE_G = "6.25Gbps") or (RATE_G = "10.3125Gbps") or (RATE_G = "12.5Gbps") or (RATE_G = "13.75Gbps") or (RATE_G = "15.46875Gbps") or (RATE_G = "17.1875Gbps") or (RATE_G = "18.75Gbps") or (RATE_G = "20.625Gbps") or (RATE_G = "25.0Gbps"))
      report "RATE_G: Must be either [3.125Gbps, 6.25Gbps, 10.3125Gbps, 12.5Gbps, 13.75Gbps, 15.46875Gbps, 17.1875Gbps, 18.75Gbps, 20.625Gbps, 25.0Gbps]"
      severity error;

   GEN_VEC :
   for i in 3 downto 0 generate
      GEN_CH :
      for j in 1 downto 0 generate

         qpllClk(i)(j)    <= pllOutClk(j);
         qpllRefclk(i)(j) <= pllOutRefClk(j);
         qpllLock(i)(j)   <= pllLock(j) and not(lockedStrobe(i)(j));  -- trick the GTH state machine of lock transition

         ----------------------------------------------------------------------------
         -- Prevent the gtQPllRst of this lane disrupting the other lanes in the QUAD
         ----------------------------------------------------------------------------
         U_PwrUpRst : entity surf.PwrUpRst
            generic map (
               TPD_G      => TPD_G,
               DURATION_G => 12500)
            port map (
               arst   => qpllRst(i)(j),
               clk    => stableClk,
               rstOut => lockedStrobe(i)(j));

         gtQPllReset(i)(j) <= qpllRst(i)(j) and not (pllLock(j));

      end generate GEN_CH;
   end generate GEN_VEC;

   pllReset(0) <= gtQPllReset(0)(0) or gtQPllReset(1)(0) or gtQPllReset(2)(0) or gtQPllReset(3)(0) or stableRst;
   pllReset(1) <= gtQPllReset(0)(1) or gtQPllReset(1)(1) or gtQPllReset(2)(1) or gtQPllReset(3)(1) or stableRst;

   pllRefClk     <= pgpRefClk & pgpRefClk;
   pllLockDetClk <= stableClk & stableClk;

   U_QPLL : entity surf.GtyUltraScaleQuadPll
      generic map (
         -- Simulation Parameters
         TPD_G              => TPD_G,
         -- AXI-Lite Parameters
         EN_DRP_G           => EN_DRP_G,
         -- QPLL Configuration Parameters
         QPLL_CFG0_G        => (others => b"0011001100011100"),
         QPLL_CFG1_G        => (others => b"1101000000111000"),
         QPLL_CFG1_G3_G     => (others => b"1101000000111000"),
         QPLL_CFG2_G        => (others => QPLL_CFG2_C),
         QPLL_CFG2_G3_G     => (others => QPLL_CFG2_C),
         QPLL_CFG3_G        => (others => b"0000000100100000"),
         QPLL_CFG4_G        => (others => QPLL_CFG4_C),
         QPLL_CP_G          => (others => b"0011111111"),
         QPLL_CP_G3_G       => (others => QPLL_CP_G3_C),
         QPLL_FBDIV_G       => (others => QPLL_FBDIV_C),
         QPLL_FBDIV_G3_G    => (others => QPLL_FBDIV_G3_C),
         QPLL_INIT_CFG0_G   => (others => b"0000001010110010"),
         QPLL_INIT_CFG1_G   => (others => b"00000000"),
         QPLL_LOCK_CFG_G    => (others => b"0010010111101000"),
         QPLL_LOCK_CFG_G3_G => (others => b"0010010111101000"),
         QPLL_LPF_G         => (others => QPLL_LPF_C),
         QPLL_LPF_G3_G      => (others => QPLL_LPF_G3_C),
         QPLL_REFCLK_DIV_G  => (others => 1),
         PPF_CFG_G          => (0 => QPLL_PPF0_CFG_C, 1 => QPLL_PPF1_CFG_C),
         -- QSFP[1] Only
         QPLL1CLKOUT_RATE_G => "FULL",
         -- Clock Selects
         QPLL_REFCLK_SEL_G  => (others => QPLL_REFCLK_SEL_G))
      port map (
         qPllRefClk       => pllRefClk,
         qPllOutClk       => pllOutClk,
         qPllOutRefClk    => pllOutRefClk,
         qPllFbClkLost    => pllFbClkLost,
         qPllLock         => pllLock,
         qPllLockDetClk   => pllLockDetClk,
         qPllRefClkLost   => pllRefClkLost,
         qPllPowerDown(0) => '0',       -- Never power down QPLL[0]
         qPllPowerDown(1) => '0',  -- Never power down QPLL[1]:  QPLL1 must use GTREFCLK1 when the channel is operating above 16.375 Gb/s (UG578)
         qPllReset        => pllReset,
         -- AXI Lite interface
         axilClk          => axilClk,
         axilRst          => axilRst,
         axilReadMaster   => axilReadMaster,
         axilReadSlave    => axilReadSlave,
         axilWriteMaster  => axilWriteMaster,
         axilWriteSlave   => axilWriteSlave);

end mapping;
