`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YHN5Kx0fkI/NAxG0s0/hJA7uBGtuBo4+NqGn+e+BcuKhfdfE9aSCvWn+9k7UclBN0wmVEoH4asGU
iwAfFQv8EQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DnExLL7Ssie+AKrJyyfZPXF/HX+f0+S+NEA+0CDWS/u3lUJupAXhiuBAiv26vtECKYWGzdrXARNh
obraRQeQPuElImXh7n9sZ02CLIhOH24CJP60FCwwur/pqQqUWFoE8/vveDuDZRmzQ4rqi79hasoQ
0iyyijKe7AtmTdLhzB0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TcaXX36lv3C2Y+E9bnYI9Rn2vCXVD1e/bBLsAwL75mSXhq5m1YflzWg9UKF55ic1b0l0d5THaabX
lcY0tnjYZS9wQ4OqdsYpa5vxAMS7snosy2pWuWtKvhjYKgOSHQwmsoWHE5Ksl7A4DcrAtEYAybEe
xoaV+sH54dTPsbLPPVc6iKp4tHhJtELpz7Fq9vsVQfehEotf86P5CTUR2yI0s/WQhmRs17ffkmpR
EsjaIB0Q6mmxpfhp4CIzgftskbLiWn/ha3CG2yDKmkZDhBad/FwpSAE9R1VeF1zm6D5YYtI6nxlU
yx5uP2KiN7d0dIbft8c6azv67S3zCOSwRLHEeg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
O1k14k+8bnP60ltYZqCFBIdDPtx++Dj5Hw31QRIdOA+IB1AhCTg+vZ2sQI+7d8dav9n+6GwIUYxU
lCgxlxH22NkhEHl9iFFHO1RjW8HgCc9dJ/uaAdrtmiB3g6XJAANVKEOssQ+Nzzm3GiRihz8rQFUV
ms7yb8g0j0oHVhMFFf0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UbRxaw64hdV+a3LzPRtutTdaELs4pP9dMqTiTWnTD8+QNHFSKGmEqDklid0//iftNx+7lnWLPT5t
Wq7/GDRtpmtdOIIhaN1Buju1qOaJYJkyiAsKPL987C2doqunfoE5MeGXcudvNWCmsJqk8AM1S3x1
jDFqgPxJY/7AzsziD3jo3eTxb6s6rQ0A4NdE5OrGui5hRi1Vh0dVjbWd0zk0EuBfh0UaU3/AIq7o
1S+EsOK8SiySV+uUmhXCKnrijC6Kfyh0hWWuykX6q7QxYPVQcNknaRVyTvbYhkAMv4NOCgtuanfB
NHS1uAlK3fuOlqc8ABh9btXkh2nz5sa2n77Z3g==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
us7LX1fVYz7gf4dKyMya/XiHDVSoQxQegl1K7YG5ssfyy+oo8e2zrP31nHQfrXBlBW6z0Aqjoyus
m53NSUCyDrO3gi17guKCemq0KGTz1xh94zOJY9waCkq0T445F6Tal47rHDcvQ5AYNl/tnjS+PhVM
fPgX1FUiejllFfXs8YtSc9UoL2jWvP/3pAdZXAegiuWRbotQ2TWBAP+FJvF6ASHtkpvpoUGhtw6o
URez6+nkGGTBkw2BHc2OaRsTv7pRzDiu0S1nHfgdTyS+B8W2X01t83Dx0ONxz6yxT7d3BG0yn7LO
WKXP413otbRU7iGuu483v4nRS6rAhCKsXITMww==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 598944)
`protect data_block
xM8jDy9BCPdlja1k+l9vJwfddqxV/ouR47dalx5EoIZ+QBoF6oFNXwiSYRywLxbxuQly74Ku1jEm
mgEr9SQqrM86tGgLdceRFmE6nemusOXnTCa6BDs2j04tFLwnI3cv9yCEvZY/3NALbwNme3ngWta3
yTUG2M8A6c4jKFCnMmf9ZSabe91nG1ZuxwuX0LDlbR7CIGO83eqFlf2P8Da5cgdaTdwv1icJn7YB
x318HDEolb1rUMJWdDyyqgqnuXURX06Db6Ywr22ZM5PuVzbi6JtU3EW3GNMue13Cp2VfsIMGP0wC
UNfVG+w4jrxMEUFwVKoj/XaLO3N7huwlzxM/lXIuitzEToH7xcE9XeAfF1ZGmbgzaEFBIJUYJLKE
jl4Tyu1Bp9IFgOpTIRIgrOd1QFgM013imZsOT1dzu7G3Mze9nG+hIjtDNA/U9aHYD693MLOElLLY
lTE12zsqw6ybmj6BDTmqqi17i4DjECvneYsmvoPVtcfAUGWBcaVy53HzIHLsgG+gzYQfuY9LiOqZ
cWalY6pkljv9kA0hhS2gg+u9m6Ht/5xX7jAFJsVGW9vVVKi/xxQHVeTc0MExb7GtiP1WR4yuMkMP
2V3TL8a2dlGE20FkAdZN69zcz/4pgT8qXCNrvbslD2Zu05X0udU31TQP4XQ7eeTK40HvFf7+oJgB
YCHnKP5WJi/6/RNTgno+cgQJtLSOnbCxomHBNXGIrgX11yWeU63PWyG6+WfNziY5wSw8cAvBmgBg
OWvBl24S0YOo9xqwQCvWhCYl7byXZH1wtobL+PVhQSim22ViC8LCZn8+/O3PVXsGuKQmh4GpdSwN
dEk/b05lPShT4GuVdWuZtkXEKk6v1a3IgFlnwi+Z/ZyD83MqpK2u/E3VU3ZXjfsXtb7u7Sk2iFGy
TBOb3Xh0e4KYvILhuE9a52h0+8ecRERBNLmkg7ZL96KYWbzK71821Q8cwYI+G1p9Q2sDD57VxFEx
m5ySdqwm0fHhCpPHocg24MVL1tV5ocMmCQfLAP0Ntu261bR099a18DNhHuN7k3TSnwe2ruB2ikAb
KmSOtn2Cp7Rp1+E/f40y2UO705RCM70SrKEkT1tv2ojs0YKNc2zegoHOQnfqrjScwkSpyKeCS4Ch
A3B/dxTJ5L68m0RDyuphOmd4fWKEIUvndogLZCSQl58b8q+C8/r8pHebpQmugSav4o1PdE5wvFoC
l9aVqpg+hVVLXu4CRsmWUMduTWYBb4yxbumIvdVx6GYJlkR+yJcJb9yNwiNcUa6blBM95HRFlZ03
SENzRuQKewCtgIOrwx7qu93vQe9y6jmTjrHysH58AVEl0juivrcFImfc3HLhia/8Xv4PlvGWaUzU
ki3kXlO14D7fBaKXIyQ5t70b4gysISeK17dJ7qeX+ch8/Zicwg+iOGqm/IWwP21rm2OdMzxUBnbG
sJUgvqFRTMq/oiy7W1077lpU4xH1APguoeV8FfOmkC96edZ8ZSG83uHZDrJkXQFf/FBdPtUZSjWH
tP8+UROkWUu5zwWt6G9EMfvtaxFfXqiK/psvFgsNTM6N4m8JDxfG4eyiIolifVmLQTsuEBlLqdqU
DF+xDDboCGMpCn3ETMnX2LQnnIN1/Wkk4vocg2kZtQ/bwqzecjN8AymfF8RLpB3CmSmdfaEcopQ6
GvYGUlhBeWPNYO0sWQa1+qQRvPu3WXDmryBSRUJUPnV00zT+PH+n3W6GakvoFQHxcKXZ8f768/R1
B3jIlrVrFFK0OHvp4SMPYOlk8xBmdltLhszUdeITuvYy1DnAsUduSn8VyenVBfJtPX6HoOSEtZSG
Am9rCAIpNN1MAZQBbTQ4KZ1HfulhuMIHq6fCSFnth3AcmFHX94DiBrRV06uUFxgHso3FjlZtOK4U
Vkh4Y+r0cblsfIQ4I0EmbsG/jjlSL/oYXznziWXZLuW7JPN/pUO7k9DC7wHSN6Jq2xZS9U7a6nCD
Yro13rZTEZdEsdeIdOGTPh77GbNixVA7US7nM9gS44HDp9GR37h/nfExXV9TEvoy1IjZyk9ELRHH
Y4ltvLTylsFNU366j13u9HBnw5++gGhIZT5tG/qVWgscPHWOhZ4QICjhp4ExIn3HxreHDPfzp7IC
xt/ALePE1kMYHE9IK8PKf0CoQXAzEnTGwNF02pJAIBNt6HhrZkUzmjTPvqebHmxLWeD9svysKFiN
oCwEknlaEaUzMqVKDdSCbC4TNoiUB3HF3zRNIDu31qc8oPWtirJmfbiVrSS4sflEF9cPorksdSbb
fybNqfDdr6YzpetOzHAeWOpboZsPe90EroI4w1CVGtTuJ5RnoPAcFIJuuUzoZhp/KMKI7vvrJdTf
di9L5+YHHoOKQzjEt/gD2wsbVa+weB4iRIV0QnzjomE9OOnQQceRFyuJatb6ZWDtVIPZaKQ6UqN/
+v691pv2pS8lo1KWO5EJ1ZdEou2WjfC17GONBhdQNSj/uJgMEAeJ16xcKVKTuykgKDGteCiOnGAn
Bzek2wtGlu4TCdU7axPZdak8t8P6e0qWrgp7W79awp+lKxNTKqZdG4ewZ+rLUwh1oIF4uueRMErx
r5Lw5cGGT6GeP96IqgJJiE7L5kXiUVNs5vfSX0WfzNpQRPA0pm0pZ7VwlUWE+p64fnl1rYro69P+
J9elGic4eb108WrNHu2qiL0J6Ic8MsUnW62n+wEcbq525Anflabnfvq673/DgnD8eI5+2juJm82p
qz9sjGLhaPSxKwuzYRaC6afvCpWEjs0dTR/KDELD3+kTomERWHLVAQuF7nj5r11UbjcvFUDJrTi1
eGROHwUaUb4WVOKhLz/RJ/KVkLCIa+FJ0o0HpMGvlZaivWse764MU/Fd2ZP1R0CByeu/XnZd4kQt
oy+HQCQdDLF4hdM2tLiUR4JEonwK43dc94p0P51LTD/prnRsHB2GDkWZMUFDYA6N8Hw4M4PDhtZG
RRzjkZlsvduDHJUy4V5naC+pcLb6tyOeoc0Pf9VuDxNOsX7xIk/Fc9NXzv9MIwa//QXLtzkBAyOX
zoh3uPKsWUXkN7v7AQ5tco2rzF2QZTqHXM5FYoeT51PZu2qdiaghj3xdjOMJRF5W389pt1HYxdXr
H/bgjBA6y410Ua9jy0Zm/kEBBev/pnsjOoN3BQ1qoD9D8pEwGf6hGLGIiSnWS5bdhErVYiHhk32n
IkxKzl93HYgFobrbRvcKZUNmFi6UHTBRTQ+jNaw5WZY1NTuwWrlXR1W4RwJ5qr3uZ7fmOoRkjTc5
gAQJJPy9MsdlVhzBHULMaaLWgcu7o4VT89PW7KA41jPPDOsasqj1nUlWv7La5YsXiHHoBwVzFWTy
SYag7eriVzzz7ByTtmm9GCHId855f6FIuU/gDpsDjJQqD94icYuaAqXS86vJX1/vb5gD9/aRvOsn
3iEVTibeNL/SgLJfjXB5PCkqI1MxHx9Z35iulTyJhYJrORW9bTbaCm4VteEcMZRv7wIqw52JL4ul
gNxtZWZs3j+DTM3XHM9Z8kb4/vP1mvtW3gXeoVII+Kf2kJyZ3m9uRhUdyMqBWXwI+OjBsdJ/d5QB
InRRI4xbUWdYMibeqi/yliJgFhDWdJnWVR1TUcJ5p8qyjuikU3Fq5sfDuEJa7U0JG7VnBozylGnD
Hil2JEZ5bNu3gdqU1a1KNzm2aZx92XRRR6Ik0i4dYwmmTeld/aZRdYiPndtIsGEtB9910iV8upBK
WeUd7T6aZTX7c7mMgfXVxSTN4LEpEkIRGbfOM9ARm/Bn++KGsw7pbEuiisJzZ0T4cckulGPOE4CI
u8SzyLPHr1PfcyGoAgPhlWESYvkR0BPZgKJaKI7yIAni/1Pu52DLzGYD0IrPJtgyS5NEvGUtQO2W
2IAQE2mVUAQ43KhGoEgaUqPREcpFS9lmZd38LWHmf/CE6/CD02q7kYjm4nU3OSCY8v1SZ0QOU/65
UaOcc/iNRly+pMx9hIYas60ZysW7c0XjWE91rJJX0Gc9O28mU27uBFGk78+sF74/bdvbfkLH/QgR
BEr3kADU0ntfb/2i7WhDA0VsCD7a9k5Fr2dYukfav4yAqJOqRNsp7HOReugWkhQHSUifBW/31u0v
JkCQb0m+/FD5YD9LS/gn5J/KBJBLGoQgqiJPF0LJVQxwMPZ8E5ZWJh0xm4IKH6kMNsKIDwIrzP0l
3UjUS2hEh4tc/eFgoOFjXt09iWey77XjIyTLm4dTWEhL0Kl4RMEZrBm5cMf1jWfqM2m8N26jI9my
cflZumgaGaJOe7fjq+PFB/XZYdVBPZ0yxW62v7FhjroQRrYekJqijQ1fRb2xMRgaGM1uKgy+4MMe
EUs+vq+LINMCBDVRnVZ/J5b6K3lT6geir1AudiNUIKMWB3ypt1BsolspKpj6AapPaGofEVH7v77v
Ckc65pH3nSmeqxPSr38H6TxbOtBK23KdQKjtNqo/1hWz679wj2hWRJYQRlStlBANsLyX34/qOGE8
EfFT3hoJBn1YDyuzxeeR5/PSVMhTgMqrL2Dt0tEZx/t5LkKfx90vA4v8IhRsXiERHfBYjqifA4Q+
Wb8BGEYlEc04WwLw7gqlEdJMgT6ZdJKh2tHGtkvFKn82Fla17sVuaPPPb/mgj41Qvu8TLegOMWe2
/XcZJ4akmY8s2fMr17q7Mb4nhcoN0nvnz6puSkLItWUr/evFTPBRls/0cPhS+oooum34qZ1FwKZu
9wAjtSMUPh3/DcTbbX9ppvBoG55/KWVAHk9UkX2U2BTzdJ/RmCTLdNBLjSFFHpFdMrXHfDddOa4H
c0zkc9lhWjCEtNVaVFvDdsKeWpZtwVhoXyrohjvvGOKv9mVtjqHspeD0bnO9DPA6UaNxJkU+BPRw
Trw28e+C9OP2CeComKyPmaj6BA9H11SxekDbEoxgiEgTYBDLrTtEv2cgCBs8wFH5HJq2XXOZpc1z
OlVZmo+kkgX1lh3eQHiNajK5HhI1nDu2PjYIgRs3IysZyOiumsskYnnD3J6sJWIVA0YYxqi8ORmp
Ziodf2lxAKdH7fsLOBiQ7rK7gQQ4b4dkmxnFUY/5bx6uNpts2F9twc4e5S/5WKrAXrWAgHsv1Tm1
2DUvlmwi3c7o8oibA1eeZmGQuAXq2ZDc9QUCHvkqta0iZBg6u8Q2dOObXIRdMBXolonCYqRJdRXh
MdW+KFQpJTswvmWhAc7douIu0Po6aqOIOiipQfV6ydUFPzTOtaFax0Pn5MteUdfdN9plR+UF1tcF
GZmG+1TRfTE/8dUSBT4QX36C98NzPXNdQQ/YEihh+o5FdbAoWqO2Paxv845+1v3y3WoOzpAb1Z2Q
E+kzLI7phd4gC4WxD57jw5Wn3N5xqfLyLVibIJgQxzas6VpQhMc2jLNrma3BBoT8dnGPu8ZLEZxB
pgT9t3KCgrsfdrXFWlgL7fBrfgqXnXl9COwSKC91IoRQZx5HSl/cjd8bm2EozC6BHw/97zsC1aE0
Hy0Ioe1HwwoFrLJRvsLPxCL9FAY3Y7TSl0tCOXgNIGu8lJgAMi2CdnIGfanb6euwoKg7yu26fJvf
q4AOOex8NmX8I79+84s84Zn/fnJsf52J52XGFXqjriKr6KTFCrEfi8/c/IfgRmz/pbcjZ4wb5ebe
VCad7WaPorr3qt2zNtes0I/FJo0pK75v99AiSJnKjQl4I9JPTewYAs4WrnwOnD9niBk8SvZlEY5t
t+afCZsg1aBMvxOTIOm59Nx6R4ox7ri6iArOtAUHSzpa/wZ2MH25aJntHvZ6XIMzRgRnuKxlsISi
N6Pt0Xv5BHIcuN6HzSE+cU4xkU6DevqCW1Pu8i6ojWPtq/vmzJeeS/tUiZo/tnosqeXE2dJpKzOQ
WqgvTXCwe8gYqelAFMAkLP8+22DTHk2AewDvTXvQgqlBuZh55K192nCsXBvLpCY/2HW7qxvhi6Vh
YbkTuEvPLV6ENmr4utY4S0sl3vUi7oXSOruedpovKVYxzK1azdaX8mO/kSbaox6+1au7Cm3mYoQB
r84v805EeW6Sz1419lIdB03lxW/h/3MaltsK1F/WukOcaTClNukdWVHPvX1A2ir8P/fpollwZQGX
njeRR8GoXvj/em28gdSKW1Y99u9dsH4RjDhHioLmAeDpkpczhDvwg2enWr17gcfxrIBuWYiIdf66
adtCykF/6+nmJpOSenLbPo2PGtHCFNIZmWiwZdLv4iqAbTwV0kUG5FRNJPokNMd5LI928WU8OntO
JVYYTBu6ChyQU8fvAmLdMFhi+/NktZw7YDPV1zvO8b5VmPzEv9xRq4sAgR9RDHMz4GO/B68jezJF
UtDyaJEtVZkhAq/uKVJCuq0LKUQqUFdS+Exo/auRB9fdSYK4T7XjyQPmqGWUpaDPCnez637TNLa/
//k3+KctIkDDdneW+pd32YY9dQ0KlWY40/NjmkLTEMSNprljPsHzhCCFGZHP4QYmY6soFmA9qJ1M
LM+RCbF7MGRecdruT0POxcH9zB1MKhs0v9pNWZ8NMQY7fx97gUQO3t9mrYJ7YBClYqM8bB6X08Yk
ASSJ+6W2YZEhe6o1Br3gcpGtJVyXQzQviUid4uOuv1lt1dakuCyo7ijuqhwAOyZnvsE84TBxGVWZ
Qhn+tfTenyNjQEQyiMgIr1b7mWHKcsD800BklFr4b2hY7rb/kB1csHMnDS/pUANGBzAJQL9vL7N/
/jzv1e6G4XyFhQdcaJpc5MUlE73W9QWAX6D3PHUb1DPQA97gumG1kAXeyoVm2sdTbd7lzwLfVJ+O
SFLFn/ekSbuDClBpwTBupInIntFpcWNXflHjdpw/JGEjz+Q++U0IXChA248fMz2YAjGHzHGg62Ey
S8LtLC6aEuHlInc2NT133HE41gssh9Djv4JsUN1H8yAci9cSu2TOqu9n4Dgwg3mBqBZrsGB2l5UH
YZ08MUEv4IEjgl6nb0ECvBfIDlEjZKLZF0dcjTAkTIweYd2AS+PNYpsLr9NgaUA0dL6kOKRHtR+J
5dfAN6DJaqrr56nobfNy8wUowZCDte67PNCyIc0yPvU7y71prPgWhRcEFJ8CHENM0sqU46Yblokt
JzmsyYmIVL1c4sXsvxwWlGzyi7sCVGN+GZuB4SVLxGv2KmvnWXHonY/tVVoSaIQmrD0YgKvWt7hP
U/1UDSLq+Qgooom1Brw9GqJbUiX0B6DZ0v19xfEhU8FDOLV2TuZU6ldPFcJjSYaWSsqj5t8AXez7
prHOOTOJa1MZpSwdEJBxfGcH4cPI/uMeMQWH1VUrzVlwdcacggfaCyXr6J37rdO/cHZrjJHbVdeY
MQMPXPtBrKIPQm6yqGj6k3KrD9IK6Qh5JD8sTCzjV/Dnl6WkDSzbKbhe10XHGy0N+Mx1xFKzcLJ3
FrU8tyUjU5Oc1boqf86BQy1EKEt5w1PkV4y3ch1356SJW68yUMb65vqexMBNyPlP3/WTHYbZaQJ0
FgnhK9aPBLxrfwisDT6Qj6spovqMRPKKu8DSILoIzsJK93pAfdRXJcIIeuTHybiybwHrOBRUh87E
ojZvne2ZiSSNPKvb7hJfMLRoJh16kcqhUVDZIUzuHJCTftRNlxiMVsGxcb2X0cjlvG/QHSNYY7iD
jBs0+SMRFPfrjyiOPpMgTJgfifLEaLrjHoCHyv/UKDNI9R9IPydq05zb5ZR0QkefFuMnxC9F0mek
yOPJZtfVYUmIzc7CHsS/Rc6WrefqpXavVMoGErr7sdqmApOyOmIxfMPcLCUwCgqTD4nQJ4wpleo8
lTrQsdsJRYoFpvJvHac+MSIw2zL9Ru9uzYXGroj2lBkloSuMQQlvxeIEIRO3/DLBeXrH3U2z7IjR
h68k/vimP244ohyzeVjNJwaw7b4MWwQyGjBVt2Ws/dwUiLa7oTvfyQq6auqBPEgrMz/QONcZHDIt
vf1Rn8WY94ZK9d1luYLYnXQ1ctsD74IIEbhBtGXZC3EPhgEzwb9hDJftLVDnlg2yXC14JWJPCBN5
p3YimCHRY6ua1M9ddUC7Va9+CzTqQRrIzlxCXmQLbxnkIS9oEx/u+DWnyGEBa3uSieS2JOsHmlV2
hzT8t9tzVzpFP/tVjPNlleEBscHDF4O5Is3Uw7uE8OFa0HmqWf3e8PDI07kSSqBTMttzBfl8r5HZ
M3yH+fUBv4xn6WDG3x4wfZGmhwZuC0IZY6FnEfp2tp510rDwRoYthkptRu/badihpg5vBgwBFtRI
MpTkzmFOdBFPVQgW0HjauMDz51lhHeRAEERaO7HCx6LkQ9ArZTFNMiwgMMV7Mkre/2N6tls9bp+j
0D6MJd4Y7zi87ugTMxcF9r9/EXWn+hFXA9NDcKVj6dxj+Dotxf/L+glCGGI6Xdk4E7m4YZUo7g9T
x1w+S8l/0QrlEBWHC2oq5UoHHcvJRgjMio+fGfWVCm0cNKfyytYGBponUtW0LGzawL4qOLMGwO28
1HOpE2NShqHcJnH2sYp6s5Js/iBa9m9wsyV5Gs5u8cLJMqup6KG5nNPS1d/dXYcwWUoBA7Ldg308
1X7fm0vMEmnb6eAMmGL40XVLtjc/nwUko/9t5mtvMJv16WMvE3TiMKKKhQKFoSX97eVKV096vsUB
Yj0m+qYwqYbJyH5eqtVCIMMZI1xkYZVKQHNFOyYLCBcFy7/W8ZflH9iYwlZeOd73exlp8R3Ri1JX
8Q0tJLRRkR65JQFPiKvcOkkLCO8+919peIfnT7q6b7wW32z1k2soJXMrcLZpzH8zjGT3BH309EiO
gmajI6q3WRaRLNCESPPLGM9dDDl8kzJhjG2F+zIKq6mt9FBrvS49f7c90CpbfT+bU7Y/+6twWfmr
ndGq55ebWfMc7pM2VXWxHlxw8+WWCFwoTESNcVc8jkj09u05zveaKgoS8BTG+EvXHu3RwBEYrCff
aS/NCO0pu7CuYqnDXQaQy1ItcIl37Bc0HTpeIHAPu2QE7MIuoOPubTGWZIy4hcNuuytt1bk3yrKj
X/Tea4YGhRCAzJvxEIFUiIFwKxd/bwgSN5+HYJr/UasprxHkejwgEB78Phez/xMGdMibuslHE4vV
tqBLhRH6NePP2zwLgqQDMVysOe015GW4uYMnmSjABpsO4yzVR767LyusRjD3CBvYowSBBJOxEqKT
PMa+1C7mpMY8E+TyH7Gi9D14sOirVQ0OAAjRcfstXspU1VSGq7lgzCjYTH/uj6Rk1HxrmWzUIncy
D2IdCZDw6W3Tt/IvjFtpXaEE1SDIQmv2QrUbdfc5vXsOFhcdthajkHUTCnli97FrMaKSxtkhQdLa
qubxHq/ucJILua/LLBL+PVYUYFV4jnaO7N5LIzk/gkDjgmEZJi67OZN+sqn1cYeleEet21MZorHU
4rgrmgnR9kP2R9MnXN+byYxF1gV+N6wAMvKztpFLSoB1BmTcOzDLYhcuzJdps7YSA90syJ5riesR
nwwsmoOO5gzBCgs2YViLpcaL51DY/vl1GPnHXCUiFyxgZxYEyv6OafAYTm/8W+403Sos11x02nEh
YgrxAgpQ+zUaAKZlfoTQYhoyrnfgaYDrk0fRLrt/uMt4GDgP3KdzVazcincwlxdcKdTBNH7KDoJe
bBH6sTb5lBD3dE6mipshF4lPQzjvzJGpSAjSKPBHRAjT3M9jnxxJ7xLLrrLXr7uXQ+Eq1s35ZTYv
N1f1gPmdDiIQ2ogPi7k3ECSPkkJOQf8ef3RhDA5d7U5BpNAiZDw9q4ekjDT3hOGWyNqRlKoWdkGv
2ZzCmCi54fcUIN0X/qROt6ldCxms0GMKkkon2tLQ4loJr0Bf288/Vbs8cGg8mnI4fdbgcpjxVtM4
tEnOl8Xar9LVduKjP3+ws0o2hDmmIdafZOOuFSqLhO+8vxYSzWOz84G/CnAfOkbSSwl8hNdZR372
n4BZ8bcxjxJYhgF4FLTYqIx8LWy7lPcd09c0JPrXS+rGrTwdfi7ARI489QNbkvnxCDA7QbBQJqlX
tMVarha4hFFRb8I+2DS/vIgOsMbwRMQeTEowNoAW/Qe2T9JwTYKhURcous++6Be4M4OnYEeRgMAN
xaqXRrhJhV/b/lx/TvJu7ccbiFfx97K2tQPlmivmmjXh9dusELajhk0qweJexnw48zpsmzNmV2RN
k74m/zh+GIeCwsb9cmsY85fnM1z76cN8V03iApmIWY6Y71fvy/+Xkht6T9OjtsKZuF6kyYL/QU3a
bGtQ3aXh8eudMPdGmDHldAs+3EiRlBOd1+3Nvv6vmgnWu6Eu75gadzTuPqzZbp6AHyFzbWqL3L7l
uiLUp17d4dG2KYLXM1Rga4YJkW1wk+mRe5yGxJltRZVNpcZwIrexILd+bD0n1LMjKgol7kBpXbzF
UKEVSctV52atuMNN9AA+2l9oLw8zfEhHwTp0hKgvVYyC34DnUJVWs8K3jiZ69z2uv32RlBAvnHnT
YKchwhADx+egIRiaKyt8jWicMCverIGNDTuQ+dCsX51BWhJNs7+JP95+dEX1ix9g1rtBqKAQwClq
S6uhmvyhqUiMp8UEldp8yY6ZHwiWbGceXAjZPfnsshTmHdVmFceq2n9K9FOUtEeZeJv+dNcCs94b
8ZE+fPbpjjYRnGHfN5tJtBYFSxYhXD6ObO2LYAwbyhSiSKoB0udUXqsmyny2zxcYZk3DNNRDt9v7
DjxDv1A+SJrATCIUyY2qXuRo/pwryKKhscP+jbVCXJZrTO1dOdSoXS3ouM7YKK+uinUnoVjAL5L4
xd/ukDCQYvB+TFezHE6SmZZ8eiHfZUkNIy1l+fsjfOxIAxvtf3priA/XQiQfYaolxSeaIbmFICxm
J3dlpyt/Y+7PstWnATMuH7Gq7Yt5qIZwSeOtNkbIoa9WU4u6JmphwSD3epDaXL8xf4D9ahin1E0B
byMhPE72KzXsybiUaaXu2W0DUYXyu0ObY42dtu20+jFjqPHiP9GWaofNYue/pkLSfWPk+tYH9uqD
f3YBw+f2RN6GijzyXVAGm43+0pdKdo7+y7LaLZApiwCml/jEXuQIwh4omL/u9bIIPofS+p5W4gz5
PDYBe7afi6TiV/G9SxDBCHyTwXc4j1fSwaJUfLYuJBJEjRRyJFtLFE8YQ7nF0fC7hXB1s7UAh/6j
40Sh7x9l/md4xSeXeBwmsXjdaLTpoOd8zPpFAcXSbfOa5NKsxG5/dJUEAos5p+vABGcDvmdsN8pD
I0yBPdVNZCARWXF+Ss43NvUUftsTGF1uijpBuqfYr+ApWKBUWV2oAgOJ/uhTlCe6nx9Hal3zSsLY
DFKPgpZwYHR/xBypWaoX4ui03yMCMNMi0Bvqt2HE6fQR1Cx40vEdR5/utn4zIVC5egYPUBpoTPBC
L4myuZU/IlXtau78kQColi2u3dkErNFC4acWNLLE35sng3XTbsb/8+L0DOdZ/BwtBD7j2vHuj7yT
4Mo7431olMLSTTXCqdXHNrgFuzLH7J13dqwcdUSmKX4qG/VnE9SiPc5kOGWrVNDZxV303j937NwH
Fx4mC0PNGjIcfwwCKeF9qH8MH9fwJ5fRGoncRV+LZq+gwCPu4NWeED2KhnQRagzTbyk60E/4S3sP
cu3QVExFXxU78xLKTi0AYcRMVsRYnmJz87ncpXY1q8qRUBLMK2D/WN/FWXItUAylaWPMC7TA7pVt
tVnnLNYedMVZ+zFJI3A800U2/FCEmktD/eoF8w+x6p48Tau72tqkr8iIFLZrpOycOeTeqlAzEgs8
ozJMX/Q8X3jLR265UJxM62DYO6FqZxu71tl656vjQiQggjnLQ8TIuTVtCRQJDP+tsfHJAFMD0WBz
x6DUDSJIh7569NAJ8adFmr20h1rXoIabecd6ogWbW6DsAhaj+6dH44asDiyetSCV+my6iVoxpOz9
vTx3AP1K8CGHHDKpLb42+3ALd1YkS4OjAPKQ/v6JjOQd2QacPb3nuRpp0g26CxypVHO62l4nCWrf
8nD1j5EIa4nUUni4ait2q9VLQxOFxIRhMlLDFVCDPk7ruu3p+3oMobb/e2UpuatWVlsIf8DNLi/S
UO2ftiQetFliw+uWLniDsk82F0iFxj1nlouB7fyKBjNTe7AerS2hlSKobiVzlxorfFhR8qprTW+v
w04V7hpjj5AKE8kRqBgQrq2WHJmNMkX+Oi/LoI+iJJdo5SuzDUE3cokhLaM+Iyz8PfARTg/Q/uRF
k5uG79/pFBCBoKi6pZOibk7TfmCelQ+M5W8g5OmjIO3FlY79mhdW3aXMwLdW9vCpN2kLCQwWm7PP
wOvKxo0CYvAX74BJ6zPq2bHBiaaBhRx+5HXUjkKvGY8mW1BgrZwca2o8VIE7dLEloiMj/3K9qcSf
pdR11iks00eYeVf5jDRHQwCe0IywdcecpfPTaQmArNQk/u1Bu65QzjoeQo7fiZrDpnECuHF1eEeK
zuNHkVLTjUpUgdRO8aciBNDKsi8LC7T64EF3boEWB4pkJFQL2xom5ZLehnCiC2mW6XSXEyHhzCzr
uZhv/jjv2uOU2DjhZ6OWBC/6WC6x5uuVA6mLyKZUaEEQ1J9XJoRXK7fOMOqKa4rvkbgYJrj61c7N
V8gxpPJTLFwNJFZedtzA23P4NSacLCoZs3kxOJqNjX8LgAjsi+0yDmHEDgIeac6IH2sh+nhfVoN4
RXpq7RIgDmPRXQl4OFsHZradPIF6mkPJ+Cg3v0d6UIgwB1vowHuzrM0KIyFtGhQuSwAj04xYPA1L
cRcfXcVbh6xUTczaBiNTtWmSQ3NTYpz84ZxXzJDNJbcPu9ZtEEBECUEKibHdhIEpOugdgnDHRL57
1gmT+3CQ1MaL1FM7oBxkAyCsYom/kJVl+wne+laZlQU+CNcQx+mW9BMSTY3v26t0uctrSZ68d1SO
emxo731tWGyFOkT/tY0/myQUI67koZIRh5PFSybiQK2VJ6WdbiFscmHw5kcNJkAMy5CJ7C5/2NxD
Ff4hntGS+8yq+LK4IWgw0il/g0fBiOViCqlqU9VpOfyalX1HKhH3mPyiIenr3qmU7c1+YvHYr+BM
nNO4DgfPs2wTOf8WGEVrgSreJWWgJGy2fNhg5uaNUfQ80XswU6zeisIuYYYwLAegCqEpLfbh9hDE
Js+l+MOFddgXcn7v7/b5ksREtzKoOJTfaQq7kG7leMy9jdme/JL2pjIONhhxL5V7W9W2Zjc9v/vs
Gomto7r20FLWi53HJT7nwGxQPUzYDaMTQVAzLnTWhE3NwgrtRSY4JdKRV2gE4mrofDXJl1qKqkk1
6ZAjk/7TKLiuviuKKlg/ZTRLIJ+DJFZHuAzISFpa/R7GHvf/dXN8qCg9TZmuubT+HAy0oMrtiASI
Iar/Jwb/ElEe/el4H5eSwJBa+a8iOOQQOqH2kcUYZXF2hFvrrHmsEWkx+NUmmiK6z8hf0M5p809O
O2u241enM+74AfvkboOW4nvy7qBNti9WrOkQMIyNSTPg3rMGbjY4qQqF8UU2NLejQHpaDB+BImtA
097+rRcLJKjlpUuYDe8/Uoa8e5UBIHJSLDWepxDeyvELyZ63HpjNTAi9qo7gpgtG3OHtMlmOMI8Y
bIgaEa63gV4gurBIzizKb+5uTp/fuXorhmORHqV9UxTLxALjJJyLEEWIUodbCdVequ4ux1LuFKag
e2TB5p/x6q69rOQwczvPFt94ThVrQ/viIdtmrpvLaAsmxW8l4K7sPxDamr4MRJBGegpSRYBeqF0r
m6fxA1KdZYbIAan9eAEkwpRH/+dCbqVixe5o93wqhul7u+xH//jyV7FE8TK3/daA7sq5RIdtmMuw
1Akiop/OHRrcTZszjsmk4JlG7SgOkmdRbAHmelTkcS9Cs1mh0jnDt8VT7WORkL63VkdxW7TrLZTq
dqI+CoTgHOmddpMqffsV3n+N5FZlC3gmWX3V/UNKFsMuPSPGLCk+LLWiZznPknJO+2n83sm+e9eH
DzKxzLRPH+YGuUTLuUOcQL6Tfz3m9cCn6GM0WKiejTyynUt2k0EhjGAYP/5gC6aHSaTK3hpBR8Mb
YxXlKVTwbTZHpQNGwi5c/BFt807G33gJbiKHUzpEXeu1PmP7e4sLNSRkNleN/JlJs2/nKwPb6PMo
/qhLmJGRYGegZDhyTfe0AX2SYiuFZYbgRxF6jnK9TSJJWJFZ1l3Z4QbQPReEqUYnDYwflUT9q08z
IgWZ2XQIfUIir4WqmUtUn0Y5iQgrFEuv/WNsB523j+7MZyNWzV06/TDPxoDzxvG+X7TB8pkmVweh
axuqMySXVL85wvk8gBuNtqvmi+Ayaj9JCIxBIZqAhctA3xYZiXGxK8Y1iQ9gcxWssrVIVI8iA5n2
dyJ5HqqOqbGntqsYmyD1yXzArR6wyya9CJ1foFz73jPRtZEP7hbl36YYNDeRki1m0arTlMlk+Kw6
KFlYnAxvPTYdf2QKyuTPqLZqFEeEL/d/aHYkPSArKh7seN/sNL1HfvnDpAjnaq2Q9PUIcXsPhQWN
ZUJfA/wxyG4yelQfWt33wWUB8kUOBkxSeIRKBH3WmaPyV9i31YBzBWKuGJG9vOQZjPsNSWK3w79M
qCh3nrNR/wGl0IpoIZDqvB1obEmEvFqiorqKZmvGOGaelHg+ctsU/fXUBvLK8LvAhsl4rD0yt8uV
CbMERdg02pWPIds8gf8ghjDm7rURv/YM8QsRerEC74KRxsSY2ikNXxZN+1pQeXUlM7F9g9V7cmmA
cROaIcdccDh422nlqV2WNT2jl5QLksKc87G2iKgvF3GssfeCZKFsohXYmlBybYM6WHXJoGOfOXC7
yWDgVmnVvC0z0ALaG5WLuodSPE70kVaPF+2jdjLYanYRdX73VHEtHfNdf/DdlOQ19MpNO0jigeB9
QNPSh1SOObReOthcXaPZYXvUjv2I5ZvqNnZRVoLi9z9Kb2+uD24u0yeaWF/nO5za70jc11fz13rU
4rwzPXyaVTBpmBRjN3p4KJKbWzKfVb+Y34wQa2Gmuj6uox1vqpRvsRPZv6rNjIih7yhSuB00/Qth
jDXkol3VU8oL8Hqdmyt1lGVrmiwiu4PU2/e5Cf4zIQ51yJXZ1LyPn5J1TKAJcYSH6G6slO+I2Cgi
tjV4RuR4pKjTzHCbnZHFICcpaKm+Egul9LQBJ+H5WJ58lx3ryTZUZLo3jBZqDm7a4FqlUdjNU0xw
PABQC126uPESCMNtKS+a4JUHJ8ACgcgwRCB3aUHPcpdGMl5hWJuLauqhMRz6zCocAasyQ1J1SH8p
snLKGpBONCInHXriVbbTDBmULc2G9ltLx0SAl3Tco98ZZGPMY+9cOLURrXYC/SXSbOpuc4aqHAZe
HmBVDbXq4g070WtYj29VOtvHwmlOFgjGfCw2EG0gz4ZDER1/EmLTUXvZ/RWpvF4XXQgS3nHuhauR
4GtF1MHOMT5LgCFxXynIDKdIz8WA/j2yS7NQ48X9OAv+NTTC7OGDr2tH8WTMghUtqcNeVlHlLfC6
BWFGlT5Im4i7LCTPcIciEqgERqqhGcidOJ0f10LY1IfAOw49oX32lSqAHmkpXpj8OXVIQrTRwPXz
uz3TQgA2vN5R+fiBKA6DeczBdGyc7BchTUILMZgUlVEmkT8WuLhqz3/2OK6k5rWEo6T7e0qDijzJ
fTMULRyNTWNpHY1dp5g2gdD4EVWfQIbpjqiDQB16RCmZPrmBTrKXnDl11nklsFauuaTtwBYIvfQB
5uM28E9kF7TLl+xYtkkOXU+U+HzV3CSKpHI+u4iKk+ath8sH+X0PAFdHrnV0J5A40RggPgoe0R/r
c1BjHEsibtZFzE9YNNn5xRpxUjxr9ZMH5Wfsld9n+q3UU8yr7S/ObapMvmgEvq5Qg3xh6+wSfmRF
KDI1AIfwFeOBLrRvJn8zjN9m6NNtf2GYmOYEWQ1ndOvKQGovtAst1Z9+4g4ePRTlVneRFKSyfRQ0
5dkxnrLDsi1BSAiMqMx5Xa6mtszx/Aaw64Qi/9e9n+aRfhdv/MTguuU3YB7PbVIYStMHtFI8rovi
GDs/VSV9t5uSzQollRwj8UnIGKs9pxXBHexFlIspPDfYYx5j/WNslWfttZrh6053rY00KoSitxDQ
4z9C32bZEpkvyBNYGaxAhwIGy8G4gvUIjMmqjdWsN/sq21I+VUcjFPLTAi50QIPhJUKXYJdfNfix
MVQtu8XtKJlYpOSmhyKp7jDoT8fiON5MmRXQg3lHduHw6lly4q/IV2xTu2nIl6G8JCqxpvWkcnAd
ueoCbV7R5DpPPunCD2pouBdHaqOB/oNnPSb5D5cx38jXhAWxEg35KyIfxkeK9gHXjo4eyZJ1yABr
58x4QtefYXtLOXnVysWTe5KtRfWMdhyl9jx+GwoijnJSV5UWglaAUlcDp6SdL0uJS02R06nkZi2O
Y5YXAGXrppK4uCYEBiYj74rKCTVnXNOdTuPdGHTAxIRpWL2i5vyc7ddzY9XSkj1B4SQM/HOhKiLX
9lXOcFGPfy0+bs9/GnAkps4STxMfpfchzexFs8q7l3/NbSRqvkps2CdNFDaG+DCwgByIg7V+LgdG
rwsRFpLefdbcFQOlPfRc19s3LBHkUVOKQwtnlkKR16llmlhsaB5wO/Thebm6r5HNaNjnPdWUtjCZ
n5VXe9koZOjdKQZLyH5BPiht7uU9B3i+913vgpQEvoZrd10YS9TLwLWwF7Z7S/Ej49MjdaFxItHn
+RGpwSAfsJXX9o0KMja1w/RlC7gio+LMlDoTazUvPdPdy8aibsMJ7w+IAFLmCNOuzTyiqex5jtNs
G+8gYWDZySwrvtzIgrmdb7dt3CyiD7domrB8Zl7XD+hCfhFPP8bbIfg1UjA8df5baTaD9JqqHHAi
yDhPcegjOjfbS2YyxYQQB6I5HQ8Yz/0gUwFknCn4fhU/a7I/Jtt214UlSHlUiXu1HlLHIWu/zLeJ
cnWXLD21BSm+Op9pD9hYOPJ1G5ZyyN5EFHHi4D1eH3RgsMlJGOWnJIY/GjMgupaGyoc2LHTfNIGq
MtxsouSqjd0zhNZeZuXZ/Go17Ko5bZVzxerMUAdouziZ2rkcOmxs+1G7T/FziOj2lKMePD4qeRFb
21H0SuMwGW1IC5jXDrYu+As6Y4SidNyBk/LakGQbmVIx8hI+NSiphkezeJpDnKrzhXs7BckeSYkQ
xuRNEnBQgdDSQzpQIALABPE69dfMyJF4uI0fPnWZsJBXKtzNfEgrOE3vtaTmvD/BQy316tHA285U
ZU6Y6W5O+zZNe2P2GxXcOdn+i4MfF7fxCFs7/eGbJy//rFvN0a1CXkcX/RMgLmpFUX0iZ3sFH9cT
cXCaDcu67SUR92kjXh85bHol9/BtulOGvoxAJ4zE+WeHyaIdDukOAz73bvjbsA0GL1YR+qEL/fCZ
tL2uh7cgiuGDoWMxhW3cLRN2UCy7AvTGojFMX8qFYdOJ41TuuiOzVSAyubEL3+4sRkSFk90G5I6b
ZN2Zarj9iwVr8IdevASJ+Tt9BbbK9VKsiWaheoeW9FqNEH86rJERG24ZNHn/+c+Jj149rJM6LNmY
E117g7dwSHLXFL1Wbw1v81bfB+Gk9jDkYxFjl3ElqdEtuqX1nWz6HUzt2YHBGVg4Ok4sLMecgcJ9
Y4cLWXGaT5ycgXgxoaxHxt38AkbqrjYvsfxWzilzRkprBA9VNGFZyAHDYgLm/HBNBzJYZB09avQ9
sfjaREZDvNQUdy/uKIxL8vX1FhjRbSBV25aje85V0noRvlcJubID6fiJJ3n025xUxVZ4th6wvSaT
QDROamPy6dnJhHrcamlmDO25wjhgFH354Bsu4MoEpivjx1P88avoWvFh1ydyPhhao6v/7Mr+5TIs
ctOrw2ySiRQypJ/jKP2T1WyHhhFcQvp5TLkp5M3dMkXhdw42PKOjOvweqCDm0rfJdaKbvIAHCvX0
xKKVX8D9egZJTZvNs636DD8Rcu1sUk3ImMihOEiW+myNqjIItHhg8tTHyrGCuTG6lLQ7P/zcYltZ
0M3Jg3hd2Ln1cOeNF033Xyyjk66PBXzS2X35yixcz4HH+jehoV2qYlEqARdHHL5qi3OP+pieetQM
sc2BOZ5pqB9npkAG/+KSXjOB7TFo/VNz7/1pRR3ePhFWy78juWc7NLOt4U2sCjxkBqGbSMLrRJ1e
qNV5W/PL/SZSiM+4lBqRcn+OkqdAkV74nDbdMkR2+2xGhok2U1ixoe1Mb/hCqtUcfSBGduLEy66m
1MXfTcpQ5Q5HoFmCn1vzsNnYrTm+Sn5iGtEcLZu3scCGHDqPjB+WxJNqZSqUhr90ozY1wO6WDvTv
lPtzjlNQdvYNTnOaK/XkRpdGXkWVcPGBMlrCOtJLjAF0/+jpx8ym4zlDez4HCs7tvaJal3lUPSz9
gR2QLOwMo3bHdFyE2wYq44JliGW8eTVbkJfJ95Go1Z5dwTT8W1OSJ1wksQN7XFSub0p6dXLYvHVi
zMS0Dhx06DN9GYgw2Mv3berz2gsSfceJ0tg7RufpJVqcxswsqvgt6lmL5cnQz1/kmrlBFsM2eJjI
YyX3PVjYI+cL7IgFAiGZIhs2sb79AEesJZnoAsDJLob1f0cjTl38yHwZdskOfi2/1tm8m7U9x6MS
GjP6cAnDfqQv4zP5I1853+dDHZ/Nqm3gLYitDfiflYAKbZEPz3b/yGM3+YRzy6Ij2XDmJtJMhUF0
HhjZGJ24ypCbX3QNoTp6VxZ5nDaNe4/eqivp8VKfZxBUXjhGto6dxTqodxkyiKZmy7GYavYWuLb0
8A5MPGlPVRVdWeGd8Csjn6+EIx5HXxiL9ZnxjT4x9O41PK/rbEmAPVnOe09USpVxNlBdYfHy5Otr
9MSVl6V6zbDqj1Wl6Bi8woWm09RU2ATCzBHmCCFMi9xbCEZ+YHXDOWo8JCqdn33hnKiSKP+XCrq1
CV7Rtd7nFDL8/v43UGJO9CmcwjXzEszHyUDPFJNFpxnFHJrXoCz424t4UTH6v0JQFwT07Glqfy1S
/x45Y681s91B7natGuIfJkz5PN9Uu5wWEdQSSEbnhb2uNVoaBAKcvpxpHnEDZiXkya4cmrJdwZkj
4ELipQAoWvZqbg+Kj6YA8IXip/c+pIvw/NkqYvLnVzEXGC0H6BCH7QGre7S9Ca4FCUv9q+fv1iAh
krzMbGK04xaq2/O4dFsLxH+JXabmcwVGsRol1D3mwG0/01u0BB3XDd4SrsdpP0gT5af3d+EdD6kF
2XzI+Xlgi5eD4zKH50fHtNtC1mcxzPrrUnu1VylT/WCgjO5d2RMNi0/XAs3Rk0QWYn86UKpwv3uw
QiW5vTM8aA587JxshKQACGetRj0WZ9aPJU3zsp5CFQd/cThT33UKWsxjEyWFnTXWQY+JPKimAu9j
bcLlB4+pFvYP01t8RTlFT3lAlR5UZNxsVOkbGh3TwApiEyVUPbPTVZO14kabZgSO79GyJ5qNyo9p
4CdbGlEKNFcGrUcwbQmptEoCIjmHv0BnB4zBIOcbqdB5PnR6XUPI4A89UKjw4F9hkszW4+u9wtrG
HJ95/Y99TVtPof/QgqeSNz4l1ajlv8qGWOm+qoAFmKqBt1qqfxLCtrXoanZU9bkOGC9kWi1oj4aL
vCJnvk6A+Zro1644GgvsHQZhMzGv6TSa9723TwQTbqis4FzxDJoyMicyYTItbBUXaLbnKbobqAgS
VWEeSlgwGJcttaV1WevyXrb991HbCcfi4rh6nYP5w3ioHnW0EJCZ4V49mqdJFVmRNKoPfI5DvLpz
kPfYeGJOcXdhzI3spd9g1iFJW9cVpQCCZetS1V1VvLGEV7RMwl3B4qrERweSCkZjnlIsmiwYHwEX
PlYfuRR8e8r0cx7JSdps0NQIp65hEr5WpurOgi0h5CdoOcwErUbtW5csGBFZOo9q4tIo3AinTCAw
ZyhVU0b8oqSpKBibHrlO3AZ3LIxWeyKZJhmYGXVEJb8xlXFMzaYzXvg4Z126q7sAD9j7wvcnumFm
WJLCnjXbm5W5MHTh8PfkjqK9lpyxbMElYR5klwh88To50d5Q8ShQJ4A6J/6tHBK57dpjO1i6DWYX
DDxVXkgrgtIy8deAsuO0VU0oYTfcmTMWYOIWaBcA0XAF2sU9kViP5+k3RZEdDd2PN6miiYA6FP9r
v5qzKc5jXa1mXjVLEudND0+9pfwsN0o0vYJuQz7su6nwLdB6SmSp1+8uS4oXitk6ECW1nq+z6/4T
Rv1G+pPydIsLGY2WDVkkbVeFRr+5WeLNcziqVoffL+f3ZQJxeTtTj1yspTgSb/izWzyB7/21Gj2l
IOLKthj+//DYyN8m2eGvbfx1LkjL/zJqHQBMuhcAQrlUZBjiErzcgLDoYua4nGkVJAlgyc92tsXs
lgG+RlggfS2oqmDE4BtbeaMERji9MwseeqAKNduo9zS8XanOasuLX7HWeSetzS0EOB2Gcj9qao6v
0jCM4OuOvMA4gvFCQ5k9ZxxG/RNNSDqPqEAhKUmJEMhUOysQEZjmQVgyuVsHdW7esCYOQ1HMWqsC
iXZOvk4UGC5m8ucbIdmwnMnW+0b52lAc+kF4HFVYWEH7D5J9IipCIle4Sk7rVR8F+Y0/htRrswTZ
BO3RwVlQiwLY30OOf4raNHEEpIR/FFRs0MJ2fiKLyGY1QrEwHLOVKFaS/jADbGULy1AnB9Z7NLmV
TaB68Hzkz9H2p+9xrggX+l+obf9OjmLEKtWrtVcXGhUTKr/TR0AbUJmyzWu+nGR19uZXHvEgniiK
WOxnAKIsSVfRvHXv0ZEStr0x/jSi98g2BikUqEmsj0mz0seBpUA4mxHvjyfJPebEptRqGixa5ZxG
Gskbe+ZSKG+kUzvVz53TSvpavREtdgw1XJBMF7uwjXDMVaX97spX/+SV1kPJBCkjaTGNe5NufNKV
K1KKh7FqVAkDi7PkD73m2JRa5ABnUqBEs6X2/kXm2L1SMBXtVDdTL47fShxIZJ9+M3wdEaYCyHrc
tJW7WP8xFfGPZLNWgSF9uxv7QyDxeZSCKWaLhboPwNajv1zazai4Wih07np8x9+s05yLuk8E1Bsd
3b8UDQM2Q/xsVwe/bs0Dx/BAHBbQ3d7FbhQtrjVrrAVbot+TsfwxrQXE77lKnzC8d1pHAhSLi0WJ
diMLT2gyJlPZzPPt1nZPg+IB4DBcNbTJftyfMJF8+pxstyxfT5kryOODcEFl7XQKxvy1lKQCzJHU
pXsBtETYEISH7uxFMdiTvEkRJZA9bGxVnXbm/DiH4/w/BEvheLC+GT0QsPDbhN+4YLKznNJj34Yz
5m/GRWWn3PJUf3IDFeJ/FpRqq4593fUbkApCl186OQUc+xE1kr9DBY4rGIHrxVdgXACRTd0iVCSR
0mGjCXLcDr2og+k0qDC9Yq9s5tCx9b0nx/jSrLi3v214yDfiiWClZwmZjYxtxPDdHGY+Ujrf8iBP
1aZHLnTwh+zB6XFWfRYynBquaTyYy73UnpWRG7lonAB5EeHOHsy8x697Zdjg4RRAX7voJNdLsVcj
t2pmY/53RpBTgQczi6tuMZIaZI1mhm7gag5D74Yrmkeibm78oPTNkEP6Js7g/WldNqoyGeHvyrZc
YtIWP9ZX2fG1I1fmsWXdn6CmYE3QNzj6gTn4bVtXl8pY1d8M8p2PRAhkk9OVBOFd1ilshOFaHTJA
qCJmfBv+oIFRJ87DE0SSg0Ryst/Ht/H/4abj4cdf4FR6u7wShE2ZSReIRFkE87h6qcufX43SllmD
Re19sAk1eP1TwLqkD29FkPci4BkeyPFxM+YqnHRROpQsUegpzGuO6uYnIof1k7x3p0O/3kUPlr3D
3cqB3ummJMXFtgJA3y2JMUEO/9H9wZ+XWQjIr3jA4izC+4u72r+oQP+KGQzIT2W3uesM0A25/E+I
yKqnlBMMjiuQH8MsVGw40GCEv5m80bkjsZ0j342j9To2WsfKmOGBLSaEDML6INF+W7e+PDgrMYDz
K43da/IWN3M6gt2+ETxFaQbQ6TwjcO6Z5RAKFc9AjFp3Qiq4wpCMCGxMDQ8gX/+J5znZfKKUBn3N
iBGKFIeldkb88i5+hPuNYcQpfDWYb5TOB+HPZsxQAoOjQOSQXmtgsSlngpbqEIinNpRELTjecIJF
ln/AcIsZRAl2po90NrGUrig4cJR80vAWaBs718ao8QNIvXCEH7c0WRfQo4NGrHFXeWXfnNapKAit
qdBWoj9jh0PBcaHVeEqmWOrLtPI8hhOXh+8RYCu1X0Bt0am/SQlxoiAUok6y6d2vz0Kx5HbwdLK5
5bN2PF0x1lx1MY8SiOqbZ2loZ00t4KuI0OxYc7azpDIxY9EIneoB2hnn9Uj7HD0c4xjfKPmsu6KP
IwEIKcIm7a3CvRJCxWPUXKk2DKX5YOyovRIZVz2HBAkEY0VWZbQD9XngK047QYPnUEBjQxE2W3QQ
TBi+BEqryZPhuU2DE8K+uPOijIAj/FadlI0eUGxGFB/Rt6Tm7cT48L8Yvz9njVAYnH792R2mL2RV
MZV1+hUVJ6rz1dDC2seMBURk3WRikE1KKwgei1QGKJtoR6g9lUo2hlcT3qnQ/QG/nmuuKuFjNVex
CJhk382kL4SEr24L/+YG3gKWNGFuQ0qdl9Eb7UzcvKhz53JQ5e0TKD/1yNgedcw1hIb629qSWXLl
sxIStJ0YugVBGZNRSpJmZY4fA/Co21GwauDpO4uWnutsxFXDA8h7eI6YaTL2g0lh/YwGNLx7A5i6
b8/kcVb52dOp0M+qz9QfjS3dmE9bNMFkjHoC41EV/oYM8VVJTgjZH8wU5bxny80eqmdLFewtdFtc
n6oPdK1Xb/jHSP46mHDcAcezKAdWX/dYnUlmhDjfMBEBWErm8T790b0Mrmar99WbDeoNvViDdRWM
TobXNdth82KiPRULc/dZEZV04OjzwXoSu9ovOLQr8WXR6UgUoYBhmNBLsQ2O1wcICc4rflPiLnx8
b9q57DsS6+IxpElBv+l0QORkYUQu57by7c+69lAex3XaLmHbkh2pjEGaHz89fj9dAWvvhyZFtBfj
L7ZY7vLoROixYh7zr8lqruNUlaH6V701FcFDW9mW1clQZYesLftcF+A6jRAZANaW1GtwQVi+B7yT
JprnaKdN3JfWTy9DQU0DYr87ba7FzlBntfjoc0sAmfpYPTvDYEBPsExrwZwgCXWw77yeyPo0V9Ik
9mWzUJQ+NQNcVXz/lg26iMUeSRj99ULTFf087Opb43BbZT4HuK50fq1uvUTmjjGmSgwT3dn5AqmB
P+rPDiVOBPwEPaDBs+a96tGTiaaaqVr6Z+ZPCfMmaep/VPM+p2jvk2q6GHlLghh48y3HmYYxS0MK
jtoLluQH1PVc2xQN+73UShvYGC49Hpf1zjdswD+L0CpwWGprhmDdDORlxHQu6BF4bzRUeWVC4RM2
gHMLHph5qw3ReD9W0bIk4htYZR7i/G7O77FS8Rexl7DyCZ3SvwjBYke2b3Aa/cgu5NnQwPHD78QE
71f27cD3DJMyIfDMWsFo0aCGzbckQiuKyZemVm5nQqIF6l19o6+PCJ/xN9C83rbYkiDocWMfKi52
KNgZD4jQcsUdseIrvwt1tUiSVzC8kNB5o/flLZeHpBxMRelfcjp/PVMxeyP1IkiliOpY94AzHo24
TGprH71ydgshc2NPMsj3RuegwVbVhn6uqRjRurZ8md2XPGyEN7oYY8heRFSSM7FDCSmcIw29ig0y
nOqKuIDbYXYjcvXly55rEyGrp6+4VFmhvwqNEuZkTswjBg1p3Q7X56Ovgznp3it3fFQqX2J57Zu+
r6cQ1q6L8BXiWUyGVa0+StNTFBjQ5VnUr8TGBQEqlhWjoI33MIeH+z+5G44KTHnt4tXrgXS6slhN
7X8pYqk5xQGXbVGgZEWRmcpOSXYcqY6rrFbXwXL07QTwFM5IfTrZbhVMLEGd8SpNxn918wxtxsAh
Dd868oiNrZGYuFA5W9REDomBJRhJ5ztyhj5mEMS5gYE/wy2uCOT/NAQr6sCT5nbYhQlqi/o8Y6Oy
rsUJEwXmX4MDf6wJ59L/81RBd3z7akUtzxsL4a0nEX+9MPCmEGjYzPbTpyc2v2P4Kcew0pDUmw6B
lVJJKOKWgtP901P79wCYbj9LNdSV6PMWswHV1d/CGHDKZVkJGOw0cuKp0f/w5rStQ5POoxkrkqgA
qCaXSFxl9CkofEcM8z8xuE3Yq1N1QvDT8V1Pd8CeyZgL8JtbQdGOmEMVvqIZJ2YcWk7VKzVeH3vz
Z7QKQGEL1ypV9PJ6cxhp4rMeMKAvhMbPZNOj8W2BczO2BgLfWWgxORzwZuoEYd4tQ2hqBpXEgjpH
5KdCkrJRLjGl26k3Ly1ZflyqY1qxz1FISrQSmAaWaCoRNXMRk2gXMw7gcBvYm6TS20UbDYCaD7/w
ZURkeTeKlcyvlmASOrbWHupCpdE0d1FWcpRdNCG362GD9MQUZP5CSBEnz1lYOHsZNpy2v9q9NeqA
XhzfZ5BklLoakyqc/rgyhbuYGAp6rKxXVkXygBCuRC6X9KgFeNEjtc0nDN42ByqF8tWw48IsaQUG
AZCg91R+xsMDittTnYCcfwUUcAh/rR0JDxwBSLdDWbFRI44n0PPqkZ3ISLNDsOzGzHFypU+OKn+X
5Z7fz4KH3RTYSswDP1UawbsIOZP3362TMqDIMrlkqz7LQzjiHVjAwFU74SoE05HJwwsYpPN8/jjq
Hf7G8lGNzyAFV+27zxeEV6/NWBTfg2E7VfQOHj8+EKVeswigf14JyXoyqzoY2fBLkhQ9+iZ02VoB
TdxUFj6ySfwwQbJY1cJebXBjCekbXWRl6O27dvd1Z/IndPCvmic48BmCf1O24TZCmo6JtQ2ttNu0
tn/gGl6LSlMIedPuknf4Xk1HiF0i1dKZnGZdDlJ11LNdFFA/IRqcqEAKxjtd5YP7ThoeFaePbCA+
uMATpCeJQ8axgCsSx6q6cgDWOxNlT5D+K6ZAxVyrqfDb000WFchfGYbFzLNo0UtTljcOlvXVdm7c
B2/YZf09tpxAftgfXgoyOjMMCdqIJ35oAVwgwAgLcHIPLNB4wo39JxHUGz0L3d0tZuTWgolKnyU3
1FoUKl+LxUnGWxlxIyV4GeNwWx7BZpPGqoxoaamJE3KO98h3mniKFodqcCaKWAtSxaPKDdDNPl/9
iQJE2nXCkKPbNzSrBVPxrr1G09QjNwGPiyHgRiuXcX3m5Gyi8MTkEkkaQ6rwFW8JE99vle94YOV5
IM3TZFupDfsuUT5AADcarxOjMrNImpPuJMfjVLn3Cy+WIXJm+A1s6Y8WF0udLHn/gQrfMw/INWPL
HoHLRmbi6kKf36DgYyBkfLyey4vazlnz+NtrivCLBOkPCtTjalno8A5v6aF5j5ezaey9FIfiPjgE
G4AqytoUR0Ej5LKMe8ak6tQ9FM/u0RKJG8Ogk6RrC0HbelksmfMbzZ/nM/5ooSRVlk094J0TDJ8Q
CCljwG2CP/TqINukjVmFS1Tbkzt+YSfmtzWV9rvvg6XTir4TBSfx6iTLhVwI+UF0XgsQdPhMw3+D
cLC/ejv7AxY+5gyr2vbWo58WSzoP/d1MPeEnF9jgpzzYJXh1G9xJsbCpvUCUYT1Go1UkXWFPfXn6
GRKVsfTJADMJPDg90sIXZZFi8ARzdZOb5WEgTzvVp+16HPokKkoE1JBQfQwJ+MKR4hAlEY9PYRSp
i3mxuq0GQJeXsaLh0HbaZEevLwIvfz5qqvfzJJLJ3xypxlprGJMcTBDhV6sllU0viZpArYDrMlZM
TZVCAStFdBTCjV8KulpjcebSiXLFyFU7R3rxOSw+SbtJZ9rboar6ZlQ3XrPmIC2vPVxmtTBbUnnr
FKuzQGtBT9RQmJ6zgbMHMOTvK/pMhtmpG6HEY0UAlECW3Ya6l8KnT9hxozIVGmvfCoNa1rNYajsZ
2iXOgQEugZQJo0rRhnTGG9/UYzhEHShD/t6aWwhPIKVmoAnwQQRDndETSeMWOsCS6mUHu/cRASFq
/S0wnUtolVGE5Pu8YrzfbdemcGdwInxGmz5dc8d2tRRL7EHbHsu1+mwQJo6ZtuoZEDnZzB4W9njY
Qt8nvYA0l6bkdZnEOf495OBvMKi+v8VZoCSPfHQYpfgjCXAqIBSbMZV6hNyZl383rTBVYDXC/XsG
ExIQ4jJF9sMGZnFkKNBcM64zu79CGL2864SIBn8O8cRoysYdGjXNPZHpvE0SgM/gebNal7xzVYaC
lJLrFvL1uLrTBfCA+5CVW8TAKlGje8bazmrMhNrZURM8p2R56IOtgwfmOb3UxGo/MxUQHtRv1HD5
w3rt2j1ysvRaIS5nhSsJIVSkHN8jtf4jJJwF/G9tGhGiAlA2LHVcXQpQ7StAf7eNcYZ4BlrTlmmE
/cmR+MtoQLWiiT3mN9KsTJPv5ioIDnZtY9OCqGRWi82QpyGqWWnfIiIWajcpUNsuTPx9rKIxL7wu
N1UHGRnhrNVTVwMnArOkPLYxo2MxDN+0BiUaUJSsNj7TKN69nm4ZHTFjUn4EDtLd8qGnDPI4asGA
xoXQ5b3TBiE9DZNTlARLQ/qNVtkGN9bKX4Dn2NwvSJn1kcMBJOZbJwQvTf5WwPbOaR/9oFx8azJa
mkJGj+cQZVlSwduy/vzMoAeXnb4QT4tyM4OprSOdHaNEz8YgyxFwC/cBftffKCFumjGO3eZlNjbj
MQ/148MBuWvTQaiRH7CwAbFfP9EiBJpH2RAk2vesdskHi2P3Pethfd/bUNFtq0lkW+AKG0OBLcAp
ekbMCNGGFAFUXiV6Ccl6j5PZmbVy31/p6J7EDTC27t6+T6lPyOZ+vbuN4Ib/gKZ167+FjqRifRVc
OspvjE1SC5MiWsTSV2QMX3+IsWvwQSkPRcbgvsmmipWpQEZEERUTCVXDkMkNiPABHq4fHJ6jmjHI
oL2CGvgWrtBLiGliZE4dY+4hRW2EJHHQQcjQXDti01Q90DEzoTr7DAxmgqSfW0Qq1DIiqxkpvPpm
oti11FBiKnJ7gTYyraFv6L6rbhkyUl4YDQ+s1XFv/BYKZJlOGZMSdLTkWpN9bIiKSM/Erd1E3KwZ
ccC8r6Nh0m3BmPfsUx0Tsm9cFmw4BoPBvMJH89EPMxBug71vIAJ17QVlO7sXDAQSou8NvdTsJK2g
f+JajeYExAMcRNyM+5bwmaCN0498JOwcZsPBm1UzvF6crDRFwb5lCMCuM848HXk+FmzMPbCjK1yK
LXjaqQ3R5vxtBnRbQpaMBJgT6zJk0SOxgpXuGHNTIom0u5OCe6TmpKyAwl0Ktwl1jdZBLLyWop7d
iy3PjMGxOk2lHvob9gTm68Spjsdp6WBwMqxXEgVXqiOSFERsOv6s1dpGip5ZmyhobfQmJcf0LkNK
lWSQOpdtq6Gla+bgM77Cgk/FQFije4Nhsgp0wa0gJZZl73UPEcKjAOKcV9fZb1xgnzU3TYg6JYN9
l0+PV9GUajSh0xPookfcffNMU1C6GssI7Ui2JoyoNoW/8tyzFXwjCBU3NuLbWuhBYNCYEDhXjz54
EFsSsf3sPIQMqXD2iyDObwkxcC7v6rCSc28Di3ztfOW0Dg0qjKGjfH/Jw5Aet6XwBxLH12ofTsAB
f351ghgVq+zM3zZQY4F6LRpWyPyiRr/Omm8IBIM1FdBZAIIeDD7SjMwW/H6tBczaprS6yXqZFSrM
KbGMAGH2dyreqZJ9eDQSJ7zI3hSggGkSE6bsyUVi/165m5gATv44Qvxe/2XM4JMUU4d0vOVHpYYG
pIRKzVXivuNWLAauzfN/WF5YE3GN54c175lSO4CWK63+4t3VXOci2vg+JCTaZ5KPl6Em3gW13yQk
bkxHgDf/pQatQGjLwnZptAUzV7vwcZXU3NPbc7+e9+i6+Ngpue+I1HUEXUOzMs8FqZC6K7A+HoT5
IPFiIB/ArVFaqoSxD3X78H5BkGxKGgASoBI9B9HjDRFjV7RmD14c2Z0l0lfaKj6QaPft8w25zWv2
djBeUd/wNrZUbTenJsCVB1aObJ5k6nXSmjfczHsW0LYCP7300JUQzR6F5nADjO4e3qy1WOy6iX8o
RbTp7GbrE0Yw1cS5pbR15JaDBTSpWauqJSpkFKpvAKOj9aSvR/sQj+PKmDrIwWu8yKGgs+zlHnoP
TM3fYE8T9bcFZyMOAo1JGwmjnVJBcxGnFs2zEk2cbf0tZ+8MujhzzyxiZbXAkWdWOcE7kHEjK4vY
wevBIjZ/qJWVpRaZXGjRcMninFKUttknh4lDQwlVsTx0OHKCpUABk+uqMwzXAKayEvW5prfL9PYF
mrMPJOG7vm/AURjKrTlTHZt9Z4X0IQEQPmJNy26sTf4rExlC02pMqzA48WsW9Mzqc1mwtNUEtXb1
vtVKfEtvbX0EyrOfArfEmXxIdcJvoAs1DkswIFONjX9EpkHkCBK3p0Vf8q1zIAkb6icB97E9dtKO
bJ0Zf2Me1FVIxSL134UYzHdn5kOhsjw5GsIX7wdSlFsKBYXiKbuDB4KBybnrvGO7Hf8zMyNwH8X7
nEo6ap8jpurlKUL8bdS8ZqM9z2fbR4MRYjT5u9o6zasBpRmGX6ObsS9N1tBpVcRQa3fjgf0xMPlg
ZhRgdSiP7pPN9BJHBCfgfaZDlWojaFzj/kvs3B7tSL91DbI6LNaIgPXPsEW9d4ZF93sz79KB8/Zk
0nVYaaLvoi6YXal2Um56LhRZ115RypvBJ/Uwq4NtxylU61HDcV+cbGgGbhN37WVZQhZ2nG2wUwSH
1uxwXNVWUklDW38ArPiYHRs9Yh136WzZygSlAHkNGdinVuyhdnT4+bJOS6BsZyA1WY/NiqrqrEID
zr2bM37WELOOyjSvHj5UomwTNFwoJzbFhLXLdhoJaYwYfIm1kanmnn6d5OMtrVArkqBv+b3BCg4G
PMcnnCSGKQXop6V2ufJblaDN0FykgWzGMpkX2vigYQ0SOXjSRXSQmm4uIcX6VIeuYpiPFUI8kZ4w
SagLMhcuzoVRBHjAvoguzQL6k1+UW7GnAM9GhHsF5yGOmtGnGL296z3h14kl4i+OeOo21MQtED/a
pvfIYLGi3vPhEBgm/glYpm8tVqXmHtyKDWgZqAmWECgviU0jvSUvsFpMDSt8xWxBTH+J9a0bQkDZ
Sy2Bsx4jBGut9ikk16crf4wAxbRv18An9Ao1YtnzioOuiLRwqa2Dpv72DidKJXXCH/2o9ot3bxYW
VpcKsvsJDxUqgAMf0xhF5g+vNIsZXZulhrzvDUSwR9dk6sBivVdoLkXeOATNOY31/EsfM8aZq1IA
EP9aHm9ye/nISemE9BlDGv/hfssPU7KMkenWz1jPwF/dqZIRJOnQsXX7vP295qx0dCpJeD7t0VQM
agDzVew8i1425fR3ujB0ZxUn7v75z5AyUBrFmxKJVgJeRPvAE8GcuaDlujZQPT+6P32dmG7OPjQ3
kjq6c7rkeXgwBc2cepEJ1vmbQoX5XERPhRxMZeZ4PBH38W9YNOJ8uITebYJLRejib5sMVwCiyCuM
Hue+lR5quqkGdKvVpmv2EQdO5EluRYq84rhIX1kRo+QD39XBr0O4uwlriWjRZ3UvlctUBh5HBasf
Oz6OgS8DAq+mcSNTfWpl5mRmvAMbl/baet4eG8gzGSBPLBiCSXKrKks9PUhvxbvK4P9g4FMAdCqD
AWQXMOwnBNsRK+ndgZZHu3/p9gXtARC1zYBDFSAxQ9/oOPFROyJCvT/dS+/kzgStqahMBqvSPFP7
17Rr7fBrIZVmExN6G2abJWvGdhRsMa/nXXTSNvdhPV1+FfwrooTBOJMhjVOjsD0OS2KwRFosLGcH
9twJAcN1bM8/PKz06v49PHFs+gT4orI+xLV8vyrcH7Cjan/OPVwvYX272NjXtHuwttOZesNQsNb+
FrChcV10wuhLYGPSAcN/yFMWy/yjgpjQ4wiluv71yhyqFZvl/3H+wXQq8so4J/BAVg4Ovmiyeu/D
oVe8n3N2oUrTpAeVD+c4FB+qCf7fMG2pil9ryXHbeoD0inpvBfCsmZJ5SYpsHEqQlkkuB7Y3fuMa
PJXSqqtgOxwfwLUtYVDaPD/gD9C4nhgmPf4pI+PVn8uacidGWB8pYUuEqBK11wsYYbqigqLOd+UZ
N0akAlYY8h3fJyMQWyePaLeWvTAdjAENS2Mw3M5LbwsbdbxrtBNt8+IPIYxECsICNZWpnzRJrRYp
SuHxtrRToRIjDTiIiK1+MCscs2AYxQME8Bzbg5oQQ7bbB6cvUMwUi+/J00zdqi9peUeHt4tokkRj
rBq4peOCMscNG3eXsNq/YeVGUd5DFeO5mWWVZYpvawvVrCOXu5xve4YInp2YWgKzL3OZcUQfGc2N
0riygL/T3xpMpePTB76svKWCe2xy6XSn/ruPzLTtL1lLYusjTfCQaNaapDrvNbSfQuLX4d7WZrTA
QBugKZktuKS2bKAAyt3Xo8zvCAMvMv7taUx734fZ2wIRf/bIRQGSApYmyrAB/P9XAuXh/zOvrYEJ
Z1MfmnyiQJ38fWvzGrWGqpoPLlJyGpKQjul0HZLf5PrZQRr9UygWW6r4Paq69eRqxpWvOxMJyx08
hFax0q8/T40Y3XWQyhSOqjhHREttyq7mMscxjvO/1PyXG7bk3aLgCeY4V/NmkXiHjToW4YO4GO7f
7HZ635W3VrBpFTMeyNl8m3E+K07Q7Ag1qyudKreEz+VbnvVRt2fB/wHrD1FXvsSKIVFjys7eIXDP
NLN57/+5WIa6WJwB8vZI9HISHGkeSIMQMQgXp8q9/HUuCG3QD0kJjREdc9y+WdJunphZCOYf2wXw
xi/IYuRI5bYPdV1oCdeZ7DSATG6DVB3DRlUhpL7DWI2u/BukeK3VHzCu8oDJE8gZslKgehEdfM+7
jQay58Um43fiN6SGzWkLX0cBJgc2LTyWJNR3xmF+6hY20+ig85/FRNMUtwd+oZyQ35D9zilsYc8d
063MsAjKyT9f9NzYS/X82zMQSY5JiQigx4UQVmF+Mru25H4DLdHUEBB4LcZMw2MyZt+Gq/2pet9P
E2v/R/bLpAneaEpwnD1LQewvcNc7VPZilN8cyPYClc26gBCOvBlugRJltbf+gLNnbi9O+g6jDCfb
b1ToPOS4KNSLB9fBcgZf0erkWMZpg6GgGHeRa0ZPk1j5j5YzIgtgWJQfHkJauAQ5Zx7dfZo4dGH5
+kxOfw2hiVVrrkf0rBsL3FpL4qTJZVyGoquj3Vzl24NAk17aArqtYIHIZxIr7H5RWEerShPYpmvc
PWDDJlwPmebxZdqgd8swRsrPAZJ0zl7JKjbZPmW0UL6g9rBsT5bpuiHIBVeTJDIvpnGV4fQLgWFB
p94Wi4cqIWny3fc09Vl0HCp0Oqg2KHGrbZcx2Le2t2mJvmuKSpmxK5io8p8tr0sduN1Z00tNIoE1
c9Hj/OnstQaCEp5uTvtCsttpyhZ/oiUDLtSkvlDbSpIKvFcWcFL9k01bKvFRtFgSMDZJFbKYMZqL
q4EgAE1dbTHzmJFBJrs8aNggNbwJp07AkvVSD46iVfsE5lgJgLxEbK8N4qQM+DwFa9Og+phkAjl9
I2cc210dTDOE23LH7DriGPmBFYVkqxP+of/RLFEYwSxjfkSByVDtc9+7WlqSPUxguv03Ly80eUQt
4Vmt6NhERUdPVH4fNcuD+4uOaQIvsORKGx/vu3XorpWGzkJAyKSt0wK8G4ZNCrKGHlzrJAgR0DZt
yX4i8aKal8rwmbV2wahRadfxhge2fpd/Ak89U6JxoqluhPuY/ecAUU1cIQHLLeJ0x2cDzrRvGuY+
l7ij6BmJlwxc54rFm5CO74M6r7yvJ1eWeyixBiK/i9xSoHrH4ARH1QwPCDcbBCUqW/LLYxCQjpau
lp67KrdExVJIGTaOwbIH8oDvYIRJ//ooRlAMRp603ODHqtpueGJBZ9qKsz5adgoJxLbUpJu0tS4+
NkbZirESanagQKy59Z6iMJA1NznXyMhM4+jobBC6MbvFKr414yX+o9Qo/eGHjvk/CPneWlw4mbg2
zmS0d1BRhFQ7OQQ65taOaYt7HyANi9OF8WBfct6jyExyqE1kGkxjDIRnCZYlpOdjzgrtNhb3uuWm
XnYtUv4a/oMvnTzM3b4E3ChQXU7GSYJkr2vK0HQ23tu+Kp6AhCK6sho17mD5JRsCYvvfhLND21xt
97qU1G7htt9t+8MYmiPfiMpWBcKG1sHUAx0SgI5K9a9RHZUWclC7fWMN1SJh7KsVbK3/R1P9wJ2A
Wutn/zqmOupNraUmxmwpfwVeGJuGG6RUE068xH6EY7zLOH2fJOzL/ul1HDQ2P2JOkkFszpT91MIx
uKwdeDoB1KhWJS2DVhpIjzQnUBw3sHWtiYlMuX2QLOp4GbyNHahEQkHda0fqS0u7TXmq0GUqp7xK
g1oYVkHk8+Not6bXEXgsGGm+EBrdXNxuul8E2pb+Yd22q8Iz6E86ERCNbc+J7Fa+mwRABefO5gEn
U/CwzgNkzCv3g48vYzC8cf/jh8K9cIWmRWBvhwsZTevcM4ax9Nj06kMy3jZUHIL1bL0OotKP/4bB
6l7Rgw6isZxAaYD77V5aOudR7wcAxytiElcXE7oWBkaEYvKUO80byJ5tMoZ6bFyUJ0iAQGfxpLx5
DPDybxOWTzNv3bGbmPA153c3HJe2HLGlTeTibZqFQGS1ksDA1HBFX0JZR9X/4eC4AdWYG8frIs14
zvY6ey1SYZ6pguxO2pUFj1ix91MdIqKBU9A/Xn7UCxFLnxJzrB1MjZok2mukTsAlbLNuPsOA/ltd
Xjqi0YanC5mdeafGODuJ3P7pEl34oFsYp1rjBqkKC+2ie/HeAlMhbBLHGgqsnBz8VpiB4/Rqjb/r
TSvwJnY+TcZtc1Dx60rjp63Z3ptIjxAKBJPW+rO+7rIgxoxKqq+NvfW1TgkR3hD3WgKDIRS+aDTQ
ok5XErEf3e77JH+otOnKpN+hhQBXeoSmYsu5aZA7QJTE70t9GvuZWim33d4mkwShEn5hdE4IGOPH
eQ+AUxmcFnfqwlOr23vyFFmq4Aa7nK45fowSTBH7dza1Sz6Vy5ma//2wkljy0Qo9K8/wYFSrA4rJ
RU2o/7U2GjVXviKpmSi8+6t7SpjP2ydJjDaTFvS1sCJ+YjBB6E8kTY0yozlsqyDCRSpGzdPOH94J
hBeUsAywlAawhoYvy2ZKlPx2joPttKqVDIzwIg4Ahy4qQjGz+AIgktGbcEbEBa4zYzbhCp3sptqk
6VNvc+3lx1q0o2Wj5PU2uUNV2RKvsS85HalH+XsjvHXnAQoWZuOcVHeyGMoX0dUZtD+5gcsObb3A
0HFRbTTOjwGbAL6Vhw0h2kjLyXPfP+ja8LdAR4lpX+DXqngD9KfpCM4QP41+3Q/FuxPreezP8tvs
ptwoZEcBiC/dlGt7acuLsvcu0tpTHBPIiGnnf7Qmnu5qfALNpPfFquE3eIpY0EzVGwyeZ208ow7j
uVBC5RKHjrulOZ/wp+VWor6Bud0pCrvtyGylPpDhIE0G/IZX+JBHROzJKnzvniffK+8CugCXIfrW
i1QmNC7jF7L6w2qMFqGVMZTYuPTGrmhWp8Wy6ZJnBL6Kfvcby/KJntpKbRw2udSzTlHpYYXcM/9S
ZsZon+846ZYxkLlDeJlalgH/yv0YjOTIHtinZCu0dBf7repIV6ARTZ4/Y3MxCTQYz5AfMfhEAMOy
Q7rfynu4zdd+YNWvA/AkxlqgoXqq26zxE1bSfDGuTS3jEAMgdFFJbRB131oYdAk3wc2ksH76snyU
Bo3R0X6BrHk9RyKWRTumuiibQqWYyF+4HeBkJHxvPUGDk51HkkkypFRVgLin+dtmWFmXDbZEuz9o
RJPAUptOcjwpVI4EgygMyX4I0R7SQfniNdopl4jsfnacQUFk8GaGJguQRKV93hHiHi/XYrlQmAPW
wifFqI5Il4wgP6FsMXyD6f3Rc3P2JHX1OEcBFOfnwfik58VsMQnIAjs0r2qdUgN6Ed92YhO7JYkI
oREM291HAJrv0djAkez7g7Gy/4pBb018XFgZl+dMCDZCbzHp8mQtTfREUHgHS0FyfyDbS4Tbyjdw
STTPwWveacPYgSAI7+oXPAgGT38qe3kYQm2qa/imPJXKyA8zbpU/YoPNCTrMdirXYYCZxe1mtOwz
ECXzw5S0HWEVRpwUx2Df6rfrxa4ilAnDDI9wNm951z+e/JIogF9ZigAhA1bdyxxjoI7uvwW2l0gf
6m0JxeDGnsaAiPHW1dixkpRahB8b0gRHzqC9HqK9ito/2ceGB5PiKBH0rcZiFl52SS+CGYzbyK+c
l9uub+r4smShXkxjzmZqALNtzNcK/STxRNqVMGU2IAtPYV/yhKqO0Goq7B8ItQNg8RMvr2r0xcJQ
G9dX/1BlG7WDB68gNREuavh9Mxo8uWv4tA57ccV08FJCa+Femp4zLzPaAmEHp0hgRxCSPBBcYzqP
ruQCGnV3iSI7MPAMs2dhAIFtrgd4e8Isd72/lpsv05pN8ROJ3nGUsx7zvMrjJQocFIHxadtkRisr
KwyJbp1dBpMsI3aYq4mXUIUuDk/U4hW6NGSXpN5YuiFzR7T93wsBUsiaCDJL/mrHg5nRcljIgrMe
9M5rCAdUruD6T3YGD1i/4d2e6UYTHjpaom14yZ/T90AwD+OmwBnO8rqhXArB/rJaytp76HtFZNgn
C+S0RGm3K5higqhcA0VS/dXevPmdmfunnweNaGoAaqAk7U8/bo1DC9Wv3tIxS35DxAUr5oiezgce
nk0cX+JPr/lgkAZg0fw5S54IAFGyy3nhsY3isUul9l33EHWd90EE+fcWXfkO0SLTokW7hMYI9Kdc
Ce0VfhmoJsFf70zln6sLdEeWbOtjG49zEgaVMHdEPQKtWqyRGU5ZIpRZ2TuO1SElXCHyZoiF76kM
RGtk+VJXQXPEx0JV+KWzqAD5NtpCm5nlO8UJM7HroLw/121O3+SwwKbiSxacD01xl1m1jfZvrcED
tmv/FlUtiBF5xNFigOzhAo2+mpIsHcOpFUUvz8WW9S3yNDKITyoMe2QI2AFOk3l/MluwIb/p5Nt/
kOgWS0VKOryJRJKb3gFebgwtxAooYkFJASRYyicpwOv9w82/zZeq9HX4AaCAfgx4KzlvXNIFe4pX
NSXm8D52gZBEsgdyLGfBs5Clh6yp4f4lOGsu3HcVpEBLi0R1Kl/gBfpVNfwDQe8Qm+4fbc4LT9t4
+u2vQPWcETPQvcS7yH3SenAyjN8c2PRDG2l9JB63B3fp1XJR/qgMv7bHDj6OE0dLQTVkqvrZPWgo
BdqdHruJsbYkfzQ2cvDJie3k1V6+qVCUKvP9MZqXvzgEUav04I9IPBDBohY8O3JjYp9gjLee6P48
KNw++hxXiT6HdiXvGa3p1u7E30qRE72TfOIaXQYnirqeMe/dG/lmS1ryjk+O4kajU4rmuw6laQGp
czrEBjgRGTmjTW3mcqIYSOPTFzEXMnRs+D0x981I3ztTTjC4h7VNm6nEp9PqebmbgEQDhOtIUUv8
kp1Sk50osXv/rf7/+oAb+30pWskITDPJAfoTTzITuN1eumSrfHOdTCyYaetaG9NkxhgtS1bpCB+L
akU+aaH5mY3bd3b3SoYlbviGgrNyLg+zcoIxJwD3St9AMkWmZWI6DAP9zfCzN9Yo4GPLg2xN8X0y
tTrVFFr3Vcfh0oKI7cDAZCRqLgVkplA/dNC/01EdcIuIh9ztOeOt6t8u0hu1a+tEaw0pkyFxICGS
0dd3yjPrwTG1pT0h5dr1vRD9IH5cdEwjyZE+TDMYFSmIngKQENA3TUQcs13OLUPvRPrtzQaaLyVE
m5vOyRxPeNMoErLeWu4MuQD5rDficC9GA+uBoKjHfEkbmJQTzMd8c3UHA5xTetvC3QN5T3b2bJ/f
1unYonDiW0kRHEHxFjyOTNNsZ3KO1IDRVqNnx75BrC6777f2vz0lzqmbiXKsWyh+r9X3ecq4CWoD
kv8cAtlru/I8ix8TZcwwZZNQ1VOuIKDZ1AFL281oUSpFVvRsSy6iolB3e9RHq+4qsXhXkNcSp6Xh
DT8AY450P8tSlq8PqboTwQZMICyhf86NGSJZhsU9MZynXcZWD/yHzAXPQsse3/yX2BVBd2WAqsbb
Bsfkc/whmkoSWITtuGo6897Oh1gIVJ6e2mcOz/VQMorBy01GzH1HoN3fDIehQb7fTCNU5H3px6rG
ve3RloH5sCNSqBkd3aFgS+zpdCViCVLhSsNAoQYmXMo8Cy47jIkU51Q2r2g3EHDh0HbDJui0ZUal
W/ki9J/C9S5bS/6Nlncr++g+AvvAvAJDCm5NwPRoa0gG4Kl92zxRZ1ZTOK4+Bm1ofGmnEgCz6LAR
AtJq7IRNelZP+QsWq7lJwJANFUJE2qjUVm4dDEoaed3fptRBn3zdv1xn+aWqvIojRDzanzDwxgGG
uWH3LTwp4fSYBe85x8TC6oOFxXk5B+oS0BxOBjIZK7RDEgYDsyV1i80goKQlYedrGHw3d3AQodqo
baPbZ7CnW8d537+ERPDh60bKsestGtaVyr7l3o5bf7VurWtxGBY7ccVnKEqqbtwAFClSm4lCtHiu
Hgy7wpMtqhBArGqk5wi4Sz0jeLS8vW3P9M7HZgjGlGW1jiUilTcR72h0XJQ/qDgYDCy+M16+4cVx
DZxjXvNdyKUQrwQRVovQqpRgpdtlocnty/8O1E95+s1aNfojnVItNLslffU1LZpJMyLB+sch9gOn
T7HfioAHVifZ/t1SEpWv6XfLibOS51eXQytz4Xg0kaqyF85lw6ijqQlDhUJvSYKe5s4TCjcRTmqh
3rc6NHvmqFHetQHJE8CX90goDlaVKhVrJ//p+otwIw7DDNk+lpLDTIa6sJNf9c9PSmiSQTE1LqxP
7Msxl1XAw3lQiHE60WeH+uEEjPazw+cPFn//Og8J5lG+9JIeppZNtE9RlJDyKZTZfbUicrEDR1ZO
pV4K0YILNOnid+rowI7I4yhFlH+PNkq6lnMwdI/gFG6op8ime0mZRz/bJ8vJ3FpBDXAv0ANdrnrX
ZwpQFfNJIZrCeBzjSEFxIiFQtPk/vdaMc/Pb++5VMJZXPjPnVdFEfq1hvl+KyUZzw9VhY5F9XxAm
7ru7vky5f0SToZ7SSWL8d9M2Fm9359C6vM4PRVnVRY8mqyEQPOmnTK7UBlqG9+KmhURqqOR+u0E0
2ToIM+HZNCmsDj7Qbd+gRSj2gWG/iPaRt/S/zg6HavqorPC0dLmqNE72vIRNNrcPp2NHQM9raQcf
uy1MIzCLpLgAf3tjgjAfufP/F4kKAa/vBlxPZ1lWtVD3hkDY1m56yR3xKMd1ZVMJWs8vGTQURAB1
16KRtbrnrrfusp0QYZFqxgpfxwe5zASVjN5QK8DAW7jCbK33xNMzqt5MHyRyEavw47X0At0/uJDV
7oIFtidCiIAd0ByJUuK6+eg5laMnKT6LzxIsL8bd7hMIQRclE1q5g6lsf4AMy6G5qM/BPUGJN9pn
31Uoaf8fZ/006zxvBRP7UuV2RWDlY7EpAEvq2N6PHI+o3XT4lNKdYi9LwNHJlDq0QjKB373Si7GZ
2C/P50mJQDRXZpmdjeVPyaVYrZZOWLPzAWYr5g7feojGbs+G1mADsmkw6YV440E7usV9xW7dJy3T
WSX24EvlF1253nR3yyz0R4K3vLrT1SOf7qaKJ3rf5c2Vk+z/hRUDccLwPyA0jR+9UiV/SHEQK2nZ
DG0NNcIPumMajN6sf95hYQf5yNSznVLZOWC1dhIYbu4/CWCFhqzePAs4gu9MRCoMcqB1orNRwpW9
xzI7wrP3bKJwcfCIy9VpG1n+gWyyaa2yvV75XDfHaQaxrgTc94rT1VpxYe+DDIkeoLnot/wzPxg7
09u2Z5+1T0N6Sd0brNGSIg7KCTvcMoBKl3fdvCvJqW7Q7KBDEoSv8hOuU9ZNWiI+vFr9BxJR0tWL
1ab1qYeTJooOeEiTm76ShfTJGH2nU35bK3TWwRqjUFszEvt9dAMYJNx4ouZOVzDrYNYUig5LFkJk
ccj7kher3S+hfiMAWmg6wHb69Ho009xWXC+7uf3ChMVOl+FPaAgfIVc2G87u/wabFZZzPoYpM8He
EBUfsxkJzxuFetNj7EqWRRiF3rnPpbO89rZh26gyEELW8QVfJjAhta/NKXhXI26OuPsTzlKXL4Gf
PyuMi+7Q/S6ZBHBLJDylWuLgKkkyM96SLxJjp552oH8lIBEDBIYmKxns3QqrAp6KyozgUTyH3Iol
y5+XI4VgpkVTDZd13wWdmDb45c3HvroWajK1lwT1lCvSPCAzZ3wqubEiHJ5NqeajKoCwPBPTGmFT
ZdwrYOV5vpQo4o65DAVN4TmQ+vERJaY0851N6QeteSI+LX7T8gH9Id/hJcatU5pKgfSSV3TrBRjO
gvPQ5/eEMV+5Wn+dsLXa6yPUnx+1dSwXdr6xf/907WnP3ObBaKZUjS8npajyzmo42wQKStSqjxhm
4549+/34GPWkovhNuoyUW3xpuOVqKK5LL9jcRy2Mchmav5+gOm2Vw1qkeNU7mZI05Nl3g0Lat+Sg
E1or1+uZYis5AO/Z6X3ZvyWRTpuKGyPacCQAcWldLCDdCN+SoT446LXGJLjGG1sfPj+WlUNuVOIF
s8i7xtQGKWVKa995UISIaoXnQFVWbejEUvxVz2mS7UDMV6FOBfkGVT0uR5hjKsu0qgxAxnIC/s/7
t/1PpZ/P1xHtvspuFVLUig/bfanKW6i7eDOaldTtJsP7vw8MkOS/WeqguH1R+DSjU5p3wW6YSV2i
jzmTgMW8nOSBo0fXLOhiVW0yq06hGGvSpeuYBi6SwjeASeS/FHGNwRkr81JljCa69nrOIfAcwyIX
qdSBVbsbe9/1993ua5o7FETTdiHL9BzKWO/2RIphcIqIeZmZwNHyRhKqDTNcaw0FJRL4F7UCpMTx
acEYgD7MPP4/93F0Kjah7MudykkrTCIWUX6mKDkE1Mh8U2wCroe/2KHxtUTfWZiA8seKJkDFKtFC
Gxv9QBXBhDBoPrY3BlCf2UkFYEr9R/3mqzlHhQQjerIu3Yo6tyJ6ehvCheqtajXwbrSbrumgLoxz
VBFWU4euyapbgETvPzXq4xN0r6C8seE+Bw+TDK5f6vBHKI4cnS7FSlvIkhL7xgZE+dVIYEx8f1hP
QIHxtnsLzeI+Ql7vW+ABV4o0uKQyHqf8Z5pTBoaolmgbfEV4LHIicibU12XwuwLq1jAE9+kV0Oxd
pvXdwkUAkp6G1dhUvIA1qCfPkVTeWWgXA0bhKm6pMmngszIMw490IKMb+PK1e+GgFnls8qTRrdWX
1x5gEKEF4rEKFY6Z4V46R8FGU7BXnXbpkzev2GPH0FK5wMI6YSggBv2+ioWf2rx4Lx1cHIsS9hb1
PtE+EnikLJQCIQ7HKnkmGOfb/Sqb4eoAReSoTNUBu5u9WLfDm7Nv4Bj8vBKRzURRUo3nB9nKcW2a
JQVk18TimV6Mpbv9NoDq3bOywQNapZmp8/nNGn/C9DWQ2cI4q40oIVbT+sjfCIWTRawbdkdzXf8q
VYHs4TdKwqvDiMz1+aCDqrRjAvNojVP+5HrRQWmpDvAU9LjAWwJcjSq7W6I1ROaTWdpyuLuL84GD
1K4NvGyjdeuLtORsT6WmC34Zx0crvititren20gK3DYQCl/7D/G/8xEIZLXUcXsqb81YWpSVXuBt
GQYuopM/4Unpli285xJGFUfIbXqv+0Q909DYE/P+yMH23iZF4ipWzjVrIsROt2EaNl/41UwxAEzw
5Usu6BJnexbfDYLK7k9ljbJhvkrfBDvdWoB87M9mqJECAPTvmd9znjrBm7QhJAWjwZrbt/pjuC1d
a3nh22NsH1JGBhKubq+sYrhGfudnyxUXheEx3A448llLDHK1Li/pNbMl2lR3Kcfpakt1ZYBgRlMW
fJIrLBgNQOSL+vUNnP6U0E/n7QNOAif8O/PAe9isWar5famJimv+u8QrdcLEj4Ce5L7WZK8Mr0Ff
k34msvTmKJ2cSKd33arf4MENbpLBqWx3g64U4bfBTLbldztkF5zsgjtLz7X6J6qkM9IF9wnbJsjY
2EMLc2cUQAyNb49uMndSxysXNdiJnTmP6L6P7S0nsd3LdcVQtTX39kgk453yZEALaXuHawv8LpBT
V5GImjYGLwkPPUyaDKtblOX6+LZrEjXXO+K6Vz0K5rNPemRebhGvcQs4AYTdq+hidVsKmvje73NX
RpUs4sUnzXKzQJc4K/iKOFIF6QmP7b24hWVlbJW8m6nkyjk0gNn0hnrdDQ5fz8v59z1pMPGhKWxv
UQycOv0KymA6l5oBOFGk+M/IypdYyVW3q6Y5624QT8/c1DBEur/3uWgMijy6b5z/ytJ8jAfD7kiC
QNg9UhbCX3TRMiCM5opWKydRjVtJ6bkRJs83HCC0gYH8t3AursIXSRVSqXNlbx2jc/nQfsAgMzQd
wxU31/P9hNrFYJ30VH0vgDDIyFVUHJFIPvECdKMG293mEvRqsn5ECwWnmnsaOsCrR11mLD7vPBhB
373hDiSjCyH9f4AAopWafzvA1zbKBQ7Edt/13/Vts1c2jXQtS5KVmqRzp3kNlRl4mMX6J98SLiya
VPjsAg+N0KodBmE7OJKv9EhW9UOFw43+5iHgteDmOb8VM/wCzJ2Ww/xZe1ty/3F2r5ZjWQB9ERcv
d1dOADHZi+cpCupT7aPmZT7QH8K1o6JwtPDnmJU8w424NIM+7wRJbRnAXtmJ7k7p0+0SgRPk+2W5
uA+I7qfSByZbSc+16/K+sZzVsi+Hg1cumUWa2HT6X5qEgPTRqbWgmznN9xBa6ZFeWrFh+0I6Z1Vj
zyt1LCjbZZbzhHII4Ekjx+eM+Ye8bDxspzNv1g3iB81AJt8oQ3Scn2TCARpfvXJUns+969pK9Zjl
cc3DG4pTiHCYbfMDIaEoKRxwYj2GTwcDWmOhw1ufthJyGhe3cHb9MI+b62G+tcdjDkati3wR8uZ/
pzQ8ooz3eurUhD/d4eBgqatu6EItL8h669iuM6CpfwNhEttYatHdIHmnZXUb1S+RmdDIWdWl1Jct
FlMnirSjrsxO6m6olKLVqelZHFrF9TgOuRozQ6eL5EZx6dT87GUS7EWbaWjHA3eI8ZEjxKwo1mfq
MRIFrgJmHV0ovkRts90gEDR8ehbMNUVAp3KXg3tiJDhHpmK+Q2OyEx41Wyr9cEnSqZnKS2QUfNSw
ZG4p0QS5FudKAYIdbzzsIzEQXRmdWLt6tkxhZj8dHAjb+XVyzPh1cJtkaT31P9AtVQq+fQHDvRQd
Ldc9sMMCjELz/R1wyZ3SLi9N+tZIG0y4zhvHT9onf+lUO+hb9IMit8N1/ptZfQRr0oPA3J1F9AUG
Y0bFe9UZ2vt1XtKErgV9s2JsWFCJeq0vxoVATg5gs7oEbfhAfr1UHNl46/alr7i4WIKi7IQA4UbE
f2PBkMNYx2I30//4DXNfHbw+dt7EQxB6X+9KflolPgFitcpNZwOiWeNUiRkubhfA4FxMkqN1SIHo
vn3sprE4Pm//IWKkSfiDHWoi5mv2EnGevehlgoklNgtHfHGLaAr6h093Mfb3MDTqsbIucb4M8nBV
uiuKO+KBUsWz+V8awmcQj7/69mb/GSvDt/GQCUgn4kcD6k2mj9Yl9AahO5Hq4V6OWfdMVX18r2Qe
bEvMfz1HnMxiwsZ8snKu8lwMmLcUXVF/M38OSLn3mFDLFgymG4uaBvhp7KP/Vlp6biBjFo8vru9t
OAEDyzlQD8zcjYBCtV4zKFDeLzXZk+hvJbKPH3r3wo7Jji5GCMc5Wh/ez3q2vzZS0IV+ArmWfQgy
pAm1AopW93kUcQ+Quskz0DfxbkCkrKOZ5AdU5dPBuDP22gK7lKXlKcFNmEZUR7xGZM4Lp7aDdoh9
yF6rK5rquIHB/9FIjwfoHxTjcIOK2RCI0GVULAjei4Ls0STEuYkZ5nYZM8U351aFIk763f9Tflhj
xcB80+/3QTTFhC52o7aIWH2LsB86usppGGP8lWEVCfO7JyOxz603lKPIwJ1RWhLyFt5Ffm8tu4oY
EvW3ih3Igqbv9mB95V4gMOwHSYE/hhiCtLNrV9Mp2xxL92dODY3y9Shi8dv5qvhtjjDMRSw6djCg
GpvvN6FtNXDxvxw9f0ybGu9TZ8pf33spwf2ppvRYiftVhAOahpoIMomh3ocC0kgmaFStO7qJLFPA
mLRb5f2JwJDdASIawWgwZBcQGMFiYgUrJV5TGHB56BKCen2SFbRojfh5jIuZYRMFtKWAGiJ0N3IW
Wt4j7+e4je52F/wNcRt3GD5Ksu1nxudQw0+E6zTqmsTJNq/cHEk2FmNsT7UwiAgMAw2SD7Ve2ssp
e9cjwVf6wMv6H9G4XMyhyzSrS1PJ1XviG5gG7mPuucQlgL10O1r3x7pnkQrQnOyENEzBjN8zx0p1
1/GlHuOMdnBeYbCqwdd0ypAlefAAGpjrKPPqbdMWIJPFUx5NhNzkjxIGYsOF5NKIjXvLOdfIoGN+
fRxakeqpWASMpYRzFj3zuqyUvXaMdNiQ+/pHX6wfBo0nz+ZDOmaPO4V/5MVLtdTgaXnPmFm4Ue5s
ZUfPXoW4WVRF0STNcmOe7dlh4fk14CXADJlyKxMVl7H9V9QZB7Egl8mrgzXMwS+6hz/jqdPbElRb
6dvRgJb97rMzBlmcpr7LqBY0urWTSBFO8Hi/shCBvexoUq/hV1sJ6Md3TahGjmSpPzpTgU/yHb85
seyttdrQ3GHsTuNVmOqmBRjaY0QqXn9+BPoAKOH4Ps5Te2R700wQpMX9e9bi56sGNV/qFuqC8IKB
dFZdHL+Ss/8vziyyvcPAYXrASbztLuZLqnquFgeL4I2yRHv+8CUVW8N2mpHqFpaR8c2Oi2EzOVgH
x7KXz+02tF+JqWJnE+uGDWlIOtdDLm5u6zjO/korQoP8MgikauTtnBoy1a8mUSc+nxyMImFpV6ad
V+D8bAcHQ9b5dDxSlGCpbS9uguuJf07Or4jnoHczI+wTRVF15x3fQSJPntkaPmhogJbHp+aUC34u
TekOP5RXKqkp6FTgB2wAPlSyPsGNrezN3Md1Ei35Wyoj2TC3by6QwbGwCNvI0aunxswqJ7KPN1Mh
5pAP9ibzxQsq/++WyqoJXvRT8J4SnmCccgmWMIvTymzK+/ajrUiigYsWxqvLmZj00qKKoWe+VDpA
XE+R6/I5Y/+puk88XqXPA7Z0FJRA/S0JIKmk3tYp6Y3sSSpZ12OffnxQ58NpKA523WYQGgEUkLlz
rZ2KdSddZTJFqooZOIAk1fo8Hi0+khYkDmmrzr/pQQHaD5bQ8wPLi/bofJvU/YLOzrHsoswbt9ZU
USbgz49AcYpb4fDOO/GAs1BTykuhQYgk1cTX4RjK/5owmdbjGz6aK/KRmHHoBOBhQnqIHAJN3RVu
VRnUB84jFLI80/OSGCO3pw3WkoQjhsMQaVCrTL3Dchagd0KEE4BklpHZc/iZKV6vHg6Hp1glaMad
WfQenzP+Z5VyqH9ToLYn1vtuTPp5W2LCbsFuEE79tDAhhZaOqGFDjeZLl07Eh12ufhIVYVvCIrat
lqcau0huwfG8dfPCViMYvbBMzW13pJe3w1mvPDToBvN8enUM5cIqWWM0bSKOCPbFHi/x1Diz6e8h
asYtGVF7+rdFr71uryaeD5NULtOKfu2yROFGYoiaU3HBpt08LzMQxZMKTRmIr6QrGsc4WAkhEtQK
DyODjau0lofhq5Qcnomj46AgAB3UuAPmdn4O0ggSC0an9X3/45/KWaeQnQlMPl7hv1LSkkwCb0ZL
UNCc8CiJgHcocolP5LYVD3lPjJE9eTkz/Uhwh8A56axD74KIcIpASn1Fq1ZQjiaP8LjKSrPP/O3b
LvIk9LcLDj68G57pvL2dXVv1/SbMRKMWjZmJY98fVAGlstjiFkb45203xSQywCgYuj3z919alGgw
MpL8uoHItTC60UiBs8BANMlm9mbH4L5+MuVrMEZoBU7UxuXOnY4Y4difgFCnSWkT8V3nLQoBDrld
AWYiLadslAZ7ZZjUDsZiQShM1BzrDx4rrYjcGOQSrVrFWjZ5hiwNxYK5mR69f44ItWVdB7qir/YF
zJ114Jelqq4VCWWnWLY87aPRS01DtXvu6AxoPpTwn/18oOu3DVBvj+UBFfgUSU0ROAE0K24Yklwq
TAHi7tEFl5R/ObgFs59D60hQ8yoqr7+yeIO0szr41x+zOi8oJlc9NpzaNLupqMoZzU7Di063Cci2
+J+5axft/s5060iRNllolWUhSQsbBy/YS69Qd7604GrfBlgM2AdY+FxhnQ3mYkHfxfx91tzVgb8p
HfQaXCbc9sz7HoNPbD53AMbu0de4VS/kZx+yNpb/sWTRoEVIM+yNomBgtjZpGALRYLwGF2VkF7It
IehUBcJqj1lblNpAJv63SMxOxNcwppiqwZpWcJcVtT/HJ2roziyehkJ/3ybmDNjtBaCNs/de9UsW
LPuIgnQy/ppArL5mmYTvKr9gVLZ3Fn1Qxa7vvr2p3wncz2dGJfl2dm5cQQSuu4l7DE/7+JSWqsD8
ymTrDOBzZNAifEGMUgWn4TwL3crCQX45izHPGY4UAhgCYPxVTBecaaIWUzgYhjKXbrs0uhM4ORGS
4Wnlvzmd2Karz5Jf7M33od8nbXltfMSVoGsGnmuVPGkv9vbCos8FjPO4+oHbGFSpzS6r0PdZna6k
0x8+AidWJ59gRw7uRpYUpSdPqG0pXmmEZhD34iUMdOjlED7Us8+tG4jE3asdFxL3symV/aTZ3lMz
YHPcm/wPJvoPRAFcAbbqE1mfdR1cpyFTDlM/SE68Vb/4tLLjKs38Hx7ijbE6hjUzUFYfJxlUAXfO
crPHs/q5ydCBY69umXSoYjyHXU/GPyOdoU1ruHZu9kQihZsiiRHyCVqhU3x7+Z1RmNEGUde9Lmn9
/C5bbU1LNzVSWEV/e7niw4xLtMXsSbY7oAgwI+KFVke8MoWyURCcjJxxAQIxHihmFIopXEac3jg3
0XH2mp6nQIVtFYNT2vEX4tR5Mc59UsfAQOoZ7wVwEpfD1ZMlxJnDPUfBzBzi2wGxad89saUgTza/
GBrt+v+DebaG+gJE/GvUBElQnh36VuviRylq7ubKkXPZFihyN+I8XW8OHA4fjVyNaKbogOv2k9c0
zOLMR684MeNf+fwL0Jd0Z/Uk5cS5u7CE5X0glzlYnPX2LYTEyYtrJmyY7xj97RE7rIhJ2kRIfZxN
AGP9gFFPeFSJYWtJl2a8LUhRS+mGL3Rmr2RIpOpKr1x2pkrf/TUmO77VPB1jB9vKgui74h/hrmFP
2YOLmV60qeZAgIhI1YPT9ws88JcjVk6NteRPWY6aCnUvg4cXNIpCnwir+fTulRa6disBT/Smo5N6
vNTOqBXuTo2oJhaXoaJkET6CyX9JSsVaHox25yAxpEGSX7KLuRClEaYit1IssTRnxppMg2cDXMk4
Z5ZmQ1a1gqyKUexHxDPRBhQJih8gwKUCgcU2grEoaBAfVmw7rZcMhyYePvuD7KVptnm+uijToGXE
PyzVrxpDTW+b09O13iG9GUWviY0YOXo8XoBSyJbAmL53beANjADXIk4V2BDJEIc/x6k/nvhlyINO
xyimL7RCIvW4Qh/YkeYWWN4uaX+MDGldPCc7/Wau6Px2faH2nT3AjBX357cQcA98gtJlYkPB7M4D
YIbF9x8BrQN3jq4gVNvEUsc/ObtqRLolvVRdq9vFmJp8UjpbxZSVs33OVRF75slCPASND6f+CsDv
mOirj+lIDD2Xl2NiLRirhnoNoD9zNjzwDeR60o8wvdyV8A6thhkG+SVEw4PnBWpPRMKePBiZ+xJ8
MKwZCxF8csP6cYP74ZznfnnT0IHm9NBx1+zCCI0kSZz7otur1HsxklFJ40qSI9C+d9FsX8G3eb7u
7gYhWAGK9xkuRwiSUT6ySm4/4Fx3+Bo5yg7AWcNEqgIWa66reCTTzY0C0qWhpZMNQAPG8TX/YqYf
BBppmMsyfvwML+oDovDQ/9NqX50Rbx2QocBWqF96ByHL7Xi1bRWyCp/LNST4uC/JDF/KstMzZvKf
ZNXXMg0eisRGfC1oZj8bZchH9TRKvH27ycQ3BBup2yZ4fP+drM5z1u4o5Htcu0/MjzpqXgc2yy6l
hgnYjHJwqLp3YCgeU27ScWmagSgXbkzDgsIZyJvPGeEs1SS3LYgmWo0moCSH1xI8SfnCXnU8JD1O
zjNnJQB2E7ZoSjf0Oa8jYs4MuGbFwiUdKVfxWPitjzPMVCaGvTN9hIBcBV0V8U+nKivneE3M1Ao+
63/NKrw5n/lmzi4es/OZD1wPu/u37p4i8M1qUusNQOu6se9qUqGgvptgs/KsRmEOWQ3pVdh23ppo
NP05CVXlehmw6jLrO5JphT8sWhioaB6CHoCwPKSCwoD1mLhEZkFNpMfYyBpQG+sfo3aunfIBsnCN
RXPd8QiN+dsm6/V8gKej40ZqNwpGejbZoHt4R+JLm23pXNBU04SgHmtjuzF/s8A7qgveY9xy8EVz
lQXoGj9A2g6wy/I2ZG16Wn1n5E0sbgDoptn5dvY86KVSyQ2xswEnTcwieb+HDdODG8kwZuSsNOh7
L95c4S+jhleXx2orXF5nEDTV1tjNO2AINo4jcSYhy5+/2DrtkYNxMYXZz+QmpWfjTGBWvkaMdwo+
cOKQKog24KqpN+8kOIDRwHnww3UTRBw6Gasr5c4yvyVzwjAE2TYAD14oOYyEpBF8xQVEb3ivhauh
o5pJXn18+cySXvi+OgEbJ+jhbxS/VOe0nvQuYlY6Xb4TPqRMRUdnlVvw0tzzgaE5OvEmBV+2Q7T8
MfjpEtMbHJFwF69Pe/KjJjBw936e99IIhqewdjbmO2iUKG1UFD1UrCc3ze9S/6tAyMyJvlcTjPI2
/Ozvzf//hcJRToxp47qLaA5ME3hstOc6ZvkXdMXALlJmGenjpldasSiqc5IFd7M2Ud/Y3hCeypru
lPNEzhGJEBm6ec7i4q5xc55Z/3yQa+Q9h3VyRDBrSPdm5Jz+7ZgHrmATM+asuJbbc2RXw09xt/qr
F9lClKlgA13nbnTzxalAe289Laxd9UKUmwOgegJpvGChs/Ueb+1oIv1oMJIPf/vWg3QxpfC1M9u1
AgwnzljYd3Ke7n9yv085JxrYl1v+JLiLMDDVDJI3zt+6PQppz3Zb/2GiWW5o+wqifV/6nYy48X18
9EMQdNyoikPwdBcjmmcMN3rnCTEzHAAramxnoaVgnHGu4fz0hfswkgaZMNKP8HU7UYa6y1LpR5Tm
wcMkCtOtTJjpQG4Iu+/XDIvhnKiYFb9gmymZ2rsMMfgPjtyhoW1cNjpWuYEweLAR8uyp7008t1IL
kwZXDKysABWKTtVlVxg8LLwE2NLINigatZqSHsDsK42DzlBgiWy8WxaExV4OJrl50MsxB/SIFS7h
3ni7KKs6Wqp45ZM8VsNm2NEFNqnrjyX1KyPXI00NLVeniYkscRwlXaCXadGtA7Mav8lvfEvKkY7I
zsrDHtPdQ0ONMQxCL7HgkD1184m1675vwT2aouSjI9BoCFLdjOryYA+jRwFJsiAarvx9/kl3cMOJ
Y/JXiUPxPp5G6JEyKyWTVrEJA7v/47vpeUwrctskFpMAIpyByt/hnr4zUt7lcLKYqEiVODBEaS11
a0wRByAqPiN+sZOmF/JDu5CZkS11QuU8iL0fbkitW9XUBQu4jJCLV/i8eOFySkZqHEYvVnTPrHsz
Xtt2vkkUyWVGk+R4p5KC/huzlIS1aVuBm3E6qFTxEjmVaBx96lOnAdLs7Qll3kfCi+mz6w4ZdSks
O8GIRj7S36Q/pGhUUvjjgfH3VFW1/l5obkWpiAq7r439J9FDacXYbUXO8HDeRDiKLfLYyHS8gGKU
XIEW6qu+qMvnSa1tmHCd4w4aFfdWV191nV8ojMHeHYo4Z0qk4odJSwoGTn/aANQJnosY1QLERaYE
ToCb6D+O141BGiSthxrBy0mtrANbp7t9AOey8ScznHQxbRGAbb2n7IwRWE/CvMVl/+1YZ6dVjJyG
18FHx1e5hW/kZbTKdx9rGg0n+RhBknlekjanavMeDoDqfzKdNBaPJzxC/E8fabdT3sGnKAtJwNN+
OOkvkStkK3r2CUKqFy4a3cR57rB8DIgYivyoxjQUoIK4UD0sjtEZlsFNu7mpLmEmhnrCkk5kvXl1
7202pn0UpgTt1u24sy3H7SADAeXtDMdcnUzgIGHFjcbYHH9S/2GRoHesjt1DlBvVYKcnvujLf4PQ
hyDQ+Fi6j1fQYwCsoX9G7caK+OJcKRjeFwJ+kmMGENQmumXYlsqRGzEzfaZUDMJ+ATbciCpFu2xf
49/LCfZW+jcMhvpHPBcikJkx24xkGLmtqwoA6yIs6VEndsPKQ+8L5zW7NvokW5pIco/j3DRe1GoU
ZIt58QTHtgF3yLWU/f75Vnd/VhlPPT8cQ8f19qNyeKkD4zquSByyw9dVMV/44AKVjYMEHs8DuTrV
kumftR1C1U+8VY5qlb4sR98SIkAFZQuPL7W2EFHoVGTGWDbzOgdIDS0GnW6cpClCA8HryjUAx/vr
dgbRAoxu0Y/gIMH2u5dyNJJVE5DMCWKqtlJj0h/P4DTV4Gve++4m+ZRyB6RhcI1oAQ8KBhAF7Ks5
k8qIA6TQFGjulTzZboUdqiwGMaQggQbSpw9yWK8j0UNrJ++6W0K4DXuonYxA1/8B3H7dhA66w84y
Ou3gGb9mqWme/DIy4zOpl/d5UQHbRaOb/wghJgjIrViH2iS5sQVL9s3EdWGXPrK70wCP7ze9LTaU
Rd2jlMHCUOTvttKuKu2O99cmn05OoWDWlO7FI8kYi3pwbu6ZRuuVzF4ngfT0JopWgilrj0eHuBYD
zuaxn1HcqJyFr7JIV4i6oYTLvB5Ivp6gKMfJM4IMSlWkrcI0RC/PhGPrTa6X8X26NGij1Tc0rM9k
wpiinsfat5a0IsNEeF2LzTpe0VCT8DbQX6xbnC8iH3CJSk8Ssm+IXhdwfhSwRpc2x7jNvR+VZEGk
nzXBTe0/hr9jZUSmqz6CYoo/ue9JB7dFD1FKsHxaw5ch5Ur1BYQjZsWB4lODs2CARg9VShsCpugf
gzcvP8ZV4fo0NmKgHehPaRBD75YG/JUNANBdLuScC7xpiCwDGkcxUM/3WEjAKyc0dB1IxCc0JX4q
CIrT0rr3N0CBuWzCweUA4d4rOC5q4RNQNBDY+yl9xOEDD+LsvrUAxfI41gZxHT/F4gnR2PyFKqLx
KC1Rd3PuBleachb9NbOlB6ML4/YJtlPXD518x9X6SlAfIrN6ogHGaeGZW4dIfLNXLhvad5yOj0aO
izlULi7ZGUuTfW7GD9WW0Q8EjEayXuGrZS+AFf5Q1NSkZ3IXZkzojYvGMMvXFDHFm6EOjWfkTMrm
YrUlyjZFVEdEJlRh8jDdingBlDtahCQHBjv9Oe8uvJ/UUNCqduL5w+T61jv1bSLDP0vZlEtZ/i1q
qBKdz1uZ5N0XaG4cxyNKeFQudKDCQOl1wHbGOz9Y2FSCo5IGeIsShSRVBmq1pQt0tWuAb1YAOIpa
C6Ic/lOikaVXfb6LkayV06d1TdFIUDBjlx89gxhsAecwhkQ/iu1rzoDN6rF+vWsB1fYOYQ12I2t2
wd4I9rNbu6KMre0vFtXhJckh8OsOHy68iVqslrDAO16SroiXnDmCwCe/n5/Nt66EcCGEz5IcQTrm
ibou3Y7Hi90WA7enmk8iS0i1imrjBYYGZA5QlbDZaJiWks+ub6yTksqRF2Dcq1v+ZcmX9WiI7FOI
HvpxuHCNNtJ5oDhjrfwhBe7X2q8naZPclFr+i4zicwzc12A0jEy2r2hn8UM65Iu+jCgx9ot2faKs
/aDR/0ekE/qxmKbQ9idLAeeWzjKWofKsAUwNosaI5kJD2o99JS0wJTmGx9oobZ8rbFzCWkQzxOmM
DcIMtvjqGiUEn+JL7zJfcKNpts/4zF+eO2XxsTxF6mAviFSqNljU2BSSav7Q5r7pFfgXP2NauZj9
9w7N/niogMFo3foPXCH8gvCtBIeAVwwgImUTvcZyyARJioEZz05PQt9Us0YMtHlf8ND/yj5FpEvN
r4B680GiW53r2YaKZbR42ZYMZIw2kSJ3PVrzaW23JlIGQhirR3LwKbhQeTESEWdob7KfaGeBRosc
YCMSCJdJQ1+l1dmichaFh4quQViEgQf0p5Tt0QWH+j5o5NQ+7eiCUuiUejfMo8dQHxPgSJzJK91J
vziNy+S9H069LNSkEdnlGqLTd9m6S8KDkuvaru+dkhSomHRS0Ntxj9GnM1HLM4cOBWDQp8i5+pYm
q5/DCaS5Nsitsy2aR/Xw/cQz/snD+WSpfcjikIcvovo3FaBZ0UVVvDeZ6msiedO03hMClwnSFk+4
lKuwX9PH9L+g9bDleaLeVZq0qGDaKt7ar7cPM9BNF4dfc46BccaMuv0GsHYlET2Rgya4RX7cgqIk
ZMLGQcfL/XnyolmkNUphT+FPf1YNefgQ+BTJp0Q0s8t6m0DnbdKr10bFOy02209SoE4vz6o+HsP+
TkS9TI2rIh8rohjbJoM3Wrfx+8d6sKRkJGlEBm9VtEbrFqeW4QMcTMnDfi0yFXztfQHth3pi/OhC
Rj/OfRZFeAF7xtIsXTDPe/6Es4Wml609orHy51ZxRtoDM3rfrfhhFBSa2rgBvkvAlx9LceUS3bBK
r1p9asg/YrBsXBM/VzZkSLfW/BIwiGt8mQ/GRipK6XsEh/BaVw5NdZO3ERYJC++Xejcxkhv5eYKs
SYpIqqjemDe6XXH/XC8Lj2d1NG5eXkWufkOrPq+hL0sAeqYRHeDtM0FVGxk7CEtv4l8Vpnbm00bG
8SIF86TJBPBSQifFGHe/s3HdsCXvt4h9cVAIRwFPFntZtOOfpPeYVP8yC0ydVwoqAMKCbOHPl95d
iFM4jgWXBGH2us5Iw8UVzj3XIioUZEEfLdhCT2doexNwAZ+mkBUg1LbpVRZ2gKateHr7TjNGOJBn
3QLHgCZkgjbuFXWWx5DzudtfAuk8kI7CtUn5/LSR38W4bmQb+3pXuXD5sWPE4Mk3N1i383GEdjU7
d+B3UH1BYqLHFnsuOGuAWFkaqLe+iIsGrDQj185jXEYXp8Mdcn2wuIYlJ/5+kwVf6Keo65dvXXE1
D84Nt5NLOxJ7l2D62/tL2BSo+F3zBjAiYU/pSGEpLrw6npgJUuC3cBtCo3RedRJU91QhYLW+2Ts0
AHQo9zzhfNDN716BOd8XLHjtjjCArnlgdsprS9I7DuuuBAFOAESTKqnyarKPLbZKiZV6kLAMiPDa
c8xhLwg3y/xBrEdDgcXhwLTvHozqr93W/ytlVoQQ9W8dO5upuKPqbXSfCSSkzpEz6YvTEP6xvvEy
ujoQzPCqm6/of2ssR8pNs2rmDRo6oY8EkPmLjfyK0dbetsjp8d/Xaubj8p6xRN1a5spNi2VobEoS
d+ifxBmfmkKAsy8ckbJY5pCSSas/77NczczsLaNKwytfKL9RTZbvGJD41GUP+ermrcE/dy2yWEng
faBmXuAQBKt3H1H+U7ZM72QEWxyeUR43UF2YLKI6eyYvGx23v2anEh6XSE0Zw2xGIrZTZ6zEhTOK
NL0vn2q92C3hPXVsBEtt5QMy2tV7hc8YC3bDk/QNsxYETuLmClEQ2mTUksS8iqs9uEgDoyUlgSyd
CTkpzN9YVd3To16I5WSuXvl8RF1bIF2qocB0gUQPm5K+zabVe+PnEQU8zaQ6vqYXTpdoajkPTwYh
jSvstcp9X9/SwIfK+ZB3SIXO7cpE7Ooxkw7XuOjkecJmHTV7QwYeFfzMwFZPa7DyPyldkZ3z22L1
DhRWvbwLeMPCnKDND1P0DP3hwOrvmcyIi4eLkrENFDdcDqSNhDd6CmQiHcTgrktDdh1z/OJF/7X+
d1y6zbc6WqOVqvUWyzpQjDjPGpnb7A2MT2wW4J5S92bHNC3RK3EI8biBBLXNQgGJUR8nTIQsHADm
Q3Uk4aa/NlzHmZNRbzryoCslTjyOSSRb0rU6M5wR/FeXojujgxZ0bFMzu88pcpnQWCGedqLT+lHj
+7MXA6l8aLK+9cBzZ3gYoBvq7wjIlg9o5PJ5374BieN2NVTJkh/N0uFELmElcD9fyg0z6kwU8VGH
GY/WCf873GmGSrIZAPPlJ3gg+hbb0rqdK9aUolht3PHQFDhw2ebzh+w5jPsGdexjlut4edyGIrsF
yvHFVb2ZVV1xtRXzpWcdTXCdKXq0GXRwKSkRKMxjdw7Hw41Qnc8nRpyLbO2y9jt0mvIEDqH7wyKN
jnWcTcoAYsBQDtK1IMGfZGEnnsIVzvjjWHx8i4j3tOLq3VoqpqBtFSMUtgqn43qhXKetwNTnOGiI
Wd0BIopLFZCV8sCASz+D2wB1qbSc5WzSnJXnF+2ynfAc+vAxaSozR3pHNA5PoEFcvcRSwXoqX0ab
01NBBznyTngLcDhIINrSCm8Y4pnlB30hifhBCug1dVAU9CYvluXevpq37Cba0OfQklCKLyDPDWHQ
618bf+4SthqRG3oe0uQ6XguMZIPy1+Oi3/LW5+UYfE4PN9AsqPZY/m6QoyKpuTAhRc9m/BuK76yN
anBpCIb2SqgnKRoIVzZcntyp4MIYudDJ7IAJC48gIpG6jZ7//6AR1eFYDFCvyBxfgoG6gWFptbss
9Ly2q27woNKv7CwiQulzJ1Cid8gsfSxyFFb/ZGinsqtRzCZXlT0eoJfVNdNP6ST+KVelfAgIWxBQ
Y7zdPpmpNQaiXEbPjakDEL66LZQRWMHLMPTE2WZ6NdiTyND/KRchtkQ5OGq9aw1npIL3kMy/Pwa4
tCw7aq2xK5hN1cFMF3FJ0JzYkbn1HmQc0z7DIkv87K0FtpNs//RxODSx9C+YTOGrs+Z28RGa6XV0
a/RCOSR4ck034ONUPDnT+8LdQinFy2VOSFqfkNpTxUCUJEBj8YAohjhmH091ywOnPmL664vb9YSG
/tVjC/X2bntkOvDxftP9NMTE4YybaW3cjDeH01hSZu4fVoOlKYt9qRKNi3BxMnriZyu06yJUZ7NS
Vnf6KCii9DaLofB5ziF9ZTE2H/WxQk7ijC6CHe9F0/x+6lOXeRAkcqUlpVLitnsC+M5TikDXEYLF
I7HNtngxdrAEcskkRm2gbce9r0lL9qtRScwqAUIxv7I2ULm256n1sIB+dJXgyqd+9hMi5hHHM0ZH
2vafIYf3f9J6zg+OcYLXEydDyzDEkGgQHRo1C5UAdhmoknSMr2boXj53DUWL+Lbwqie8PVvnEful
o/Ref/sUS+rwIiD+4eUtLZTTw9FR9/dp4VmZoDdtHQQViOjTpb49YvOGbSaLf2YNwHwd421AshEb
efZu6gIXrE6XICtRiVdQS/6Gmr/15hUdBPRX5PIIKI8DIrhcMqoxFdtvzmzSk+2DYPDxcZk3IZb4
YoOs/+V1op6B01pHsZUhHgwf0IV8GCPRzB4ezKfRNdVGF6nOVBQT2JdJq8B575dfPjNq0E+ghW5L
5gNk0XiRZflKqrQ93L5EyRpEr2HP1ktigfDIHIQOU2/un88hjlKri+wSoTsXccFYfm44L32FY5qx
mAwaKqor2inytkPdopT70kzs1qTeefvaZmASAKnuaTF+GY++lTeh8+gNDy2XnyRlqkoltq+idvuY
uyVGqjSCPV/OoyR7a1t/nbTvuXDN1eNImfKfV22awjvzfFuvOEOLk9u3kTTYsINIorFhzGCnRfP8
oUgnHmXk2YiN2rkISfVAN0JX4hrNaArOkfJmXzudIhS/JPqone70RlEdwcGOZjMkMUNoSk4gEDZc
EoCGjJUIWO9tW8e72C86dAv+CHc5jiC4s3UIBnc9QQZCuYyi1GBEh+UBZpg9TCbwjVtXDHsficVh
vpPYP5sSIMTj1aI0JiV897YZDjPMt1gA2zCIrYwQxo9c2mqFZc0DnV4RZBYQ8UqsCmYuADcI8ePe
5zCIGIk+/K7FsANkUiaqx8BjRg+gs+Uto0xCiPsU3voEwLRgjfhQZMa127UT7Kf+znisSHGhkdJI
I9Y6Pqow8ctC+tzUe61jMaNpzf9rClbIY4I/2aQPxOrYv4ae1HaA2laiLG+0Mvd3yIDnJU9VZyHC
aed//XcfX9NLm3d+xHQh7imue+L3ZUASYna4j1sedjFUrNcRxXuzfhIByHqC08QLb1/o8GsWOPqe
30Ctdi+Gglneklie7iirB4oKv4R8jlDIWjKGJW5s230/n5ke49cmqCQmfHxsnqRh5oToG7C8fO1P
PdoBO8uudG81MwwIN3oipGdQ02QjlZDNanjyrF7sUIxPL8abIDNEHRsViIuKJVnYCpnltit3K09w
XAQi2liC/6NxYaKWgkErODiRLdn/O5KV8Eks1JZRqxZqH5e+JtU0NGNz/ztPf1Gi9BbT+2+aI9g/
Jg5G+5p7HlICSHbP5XMS9BGj5gQXjjm8gecM4KZXqyVcHJOtISgblY95yG3O8Q7hh3v4ZUa+2FCt
V1v3arKGPvlLCO1g/rh+GcdaZLQbbbxmLa/2CCQY/fuRildM6rDsmD+DQFcdL7gxYAyxDf8hlvF2
XPPVdHBYqbcMuzmePw1+yXHmrb4oJbYnHDcTB8gokegZsA7hCKkXaKmCjZDDvBHH8xveCfIxGwRN
AdwGbfSXvenyb/uoTuRQ0HXsODQJSD+r8KBxh+rN3Y5G8PlnrVyTSzbEGWJiyod5H29LfFHNBX29
0CT2D+ZenRzEV/+54bWAWol8W+3Q2Cx4b9INEcR285OpKQKQx+FoPhkG0q3uG0fXzAJSSAKlGa/8
/drk9qdxZYEgq0acA9vCTmsQSG4IZq7Jvd5OEObg7rxtjpu1n88OSdQX0gSf9pW9Xm3E4jiyd9hz
NkLDKpAGQ/rp7At9ziHw3lDzOV5NxLlnrAiE5qAzvP1nKhhINb6NL3XZNXwI52LEUpDV4SHA9u5w
xksNrdYsOJGUj002hLGUWUnRzsynsv8VPkWE8hRJTTDUzsBTIhUz6qUkK4lgxDDcJf2Ym58FsSlt
YjdWD4uUwhIr7Vtg4gL3OdwbWssezczlB4qeP2W00nsukS6RTcwsPt/NZiEmy+Zg6TYSzOJN7+96
z8GwLMgVxrm0dVbaVjNlgwjVIOTvuP7Ehq4d8VUhZ18ue4KwgImrybd2hxfjfUVdniQ6Uyk1eR0p
lZ5BbU80fkbLmc1AfDrgcA60rKvwxXL9tfJkZlL1vThviaac1oJT3gWZopodq/pA13yY7Utj7cRR
8pJtQ7gRDVJ1qbYrzTfy9UgSNVMKenpABhQLoo1m7HUeLWRrFyVKvD4ROYNRtWDQaYDJwI3t4ecs
9PArp+7AlNwW6TXOEiCJKr4C2oQ0ZLVdtjrpyL4s3l2S1OV6ewoetwp61MlcJHAKJ3SsupSgzWUv
FuKwy32Fdh8soRKYvNT4MxJbDk2G3OpF5Ff9Dy9tkArxmT88McfLkeSwtumbp8XEftYM9rHRwnc0
afWetRyRdDeUxH40X3LVzk16nYdnu+82z/p5lI8rX1W0MpYgeY3tBlt7p8eYEcOuyjcc8EdcqDed
q3z/zRYwS4fJ7HWI8bPW8xXxfribAPaqROLs2HwHrzyXFQRfDrWnSR99fwvBuPCtaGZ1Ru8kZjkp
cmiaM+OB023L6nE3CwDSis5dvy40pzhmSv1rMPfExYuHtX4f/CukgWzkO5RA0UdkaKxW2rm3SaWC
oN1ga3Osj/nNfEaEv6R/wteq00Dxw4c/IMj9erKMV9k0S/B1yYHUP7RBd8+GLHiG4TTeDjuWMtPT
zV/LpoYJiwl2CQZzl5gqA1DbElA68WENFEhmvKCUiQ7SPyUvU0uQBitw9JAe9mH6+yGIyxkWXvm3
75PdsgUb3v2CWUaKF6ldPGCBGoHH4h75t868KylFM4JiH1d0MpkwfjpJYIf8uQH8WGV7dxWFX270
8i1HxhtAQqiQGrQ1sc/ESqr8V2cJjhsOmp1dQ5oHCunhK4magIptnn4nJI4nPUgHxjtmO2Z44Uy7
yGYA2NeRW+nI9Mes36nEFr8+11gYpMUgn1TobJSREMr/r+uo5m9DNdnH3wlPMfoLwUMAKVi2zOko
jnDtxblIqh/4fcPlGMYKhpzNk30LPYPGEM2t8G+oMTLragxgn4T3+z+uSV9RbJTisPwpCMGpHgTq
1I2aaIpD35X6QOXOQeBTKQNBld/mGeqEQ10+J8qoWFUZFlZo3+zEa8LOw0f+3rNhmndjZLT+TeTD
8x4hrh+oEeS8O+jk+9iCb/qe3KwvaGeTzpwULapRIIKq/doD016jfwTTzYDcq5vPTbDah3XcsIjv
IuvlyJOsf+YeFhvAFhFzgVkIBaF6btMdfrYhjiEHt6DFlTCXRZJALF55jRin7GcdGE/LxEl97Oaf
XQtsZz1X6uHZ7wa7FeYfhTIIS8cNFqS7rBnsGftkoDVYtwITKo7KkAfSXKXIK8h6xWKg5mKZpc2m
HyMW/MAzKgAxKdpBujoe7aLSPzCax01pHLGeuU2kgYkzUy4FZxF0t2PmPFKxBhfkJ2brOKWJJyAy
OlvEMGATNI9i3B2fWshkBM3cA72LHwlQmEyTpuLt4+3nxNXG80g0dmaY+lLTXjQAo0AcjhvmFigk
IrJuumFl5xk+6OUNJgCBS67jg+WUq3fNgzI9T8DudZspwA6vPET6sgCGMYoEczG8Ci12Kmk34PSm
o7zia4eaNw9FeiyoPmjW9RjLif4PXnjRX1Gpi9DL4sZ9h/pvgiTrqzXRofns0w/aSLOoE/5UvBsP
ogbwGTm2jrOPee80YUX7nF4ShbTe2XJVwOGcZVWVHGNMmvJA9jiDnWV51cyXI4whxydb0U9g8rp4
nPliS4j6UibKerwWjkl7u11iRKuMdQ/YBk9jDN6/DZ7VLN+aUMKNelwhUPFJ9FHMNB8KwAZCSKDi
Ht3WQECH8zOdY6dLrKXlFPkuan3JIbjYluR96cd5BYLbPlXMfkYfCDG0+SdtRvWDjTHnMFbcsP3c
7fQs/6AngsdNQyYCJlQgc0I35KLCd/CQuCkJKMIB5rPOPadRKPOotv0O5GhAWprkkVbVTK4PBxCr
Scni1OTGozLpx3fDJsmTM0bGQ9XJan7A2ytJugr5R+sXYE0iC2lSOos6zBRGYZabb7SAsrd+xNmr
lhxcUhinF0gwhNx3rAhO1hJpu3MSzvwHMYTlldYuciuJpB9G69igboTiAQOcB//2GDOUoICdoJEg
IqTxc7uzuLoHs5qMHoLjgTPRYNdFF+5Ft1J7s53345seYwnZnWo5iMbdemLL+NhHWjTMussyQh6x
HFGYt8f+KbNfW6q1JcXGGVIRpIeIXHX+bTYspx0hvJoHpAX9Lci780T1BWqQGnCkv015d3zz707T
/0ZVmJCu3NEsQzny5QW3xq/EwDEAQqSQASENw4E35jOmmWrwFUAGHMNejsQo5Ny2ZwMhtaO4mpAc
/xKW4/kh3Ezohesi0jaAstLwafia+T3ZzYCtcinqnG7P+MVpZ8JEGKhu79JsLsxFtVPdmNzGuFvb
scxbCPvJJqdOomMs4NcmriVZAqUaCGA3VIQxJcLNsUCpaBZIabmdIS7PB51XGMetgL8NstlaDlSX
4t3D9Z2A8yMcyjBkVESibReytmudxKqNMvvODRP94WP1hAK4rAzl5oI4Vt1RRRvSnb++J02ayPi1
ibxC1g2NgI9XhhYJLnYfI9lVekEFvvhqW6NhL6j/gTp1rLbiRDcDHJgDX/0pAaEAyeYK4voQUGWr
uD08ynsPWDuZraMMU8yraGZnIEq0xzLKWmm4PsF4eVodzdO+mrRzn0TY22bBh1Y4jiEQGatIOpep
dkhvCXk3zmw0UESPwt/p2mchkCc1VsgE9BFR16Iiitx6pHUHxD5Yj/f/1GKrrXE151uWQ+7FK86k
NF/iSbkG0wOYzAn5nG540JF2a/K6j7r4ihmIlBx+wutLunh7MQtA9Usn/03Y4coYaN5HQavhJ50n
B7ItMQoxBWoro/AW+ODjrAEimvZQqWhCn/tOe6pcfGZNSu8fnq2ccv6mKGD5V3OUwkycjnvylhY/
TlpTk4M4rvalfSG3dkPVay7uVJb6Cku5b5aImaCn1eIF5x7w5B/hRdrl2kz27PbluBU9C71/+U8M
lyQFSAErWSSVqqiaVR7NBQcGBDa8pWH8EUDroejT09ZYIoOjVR/ZBYqgdBNooi5ii2IdxcU32qrS
HjU+c0gjSvU3iOtTOFqjmrNA07zpr3cMdgFypGIXgqUi47yfkodpxHwbwao2wtUjHfvbArlUgO4V
+g3ABaQahKq4RCTejA2A1DMnqnex/9Uu72AnZeh2efkvt4dmuD+FHw/IaoeS37xpvl/F8bthlBWp
ljJy8TkuA43si4/jhZIwibmOfE2ar1hkHT8R/iMGT59mK2qXd+EVJ5Jrqm1J/tGJqT5LZaPKEedJ
e8yrXafvtxm1aIeD1rt42y7qmnbLgg+2TucqQCiD1rObEflsjLdjtDuq0ZmjawNqizMj3jbjyVKO
//2X/pwum0ESG9OTqgdP6zurI5Gj2z07/y3+Y+tu68lQGfpWIp/RB/Q7ZnmLURz7tq/kCY2BtZlo
EJDcOd89yL9FgRl+GHENXCtCQBgPTVyaeKRCfvmqfpHAme8Q88RDZZmaU6cdlZYaj0NickZTPAgy
IRR0mzAnNccCXeWn8bVl/eZSUSesDerCSied1GGcGPBH2dySIM/+f2hiSdiyc4VOTeG35yydQ5kY
IPvS7dAjxpDzVeirECvVyl7hvEVBcWZUCv7yRn2MDYLy0rM8yoxO0bGgbrMLSA0ueuwuIujtpMMK
LQ249Ki+PtWPCHW2WfJUYqhGwoaemhGTQF1y82shj7OVgNq4Z2NmBXh9y08YicXPGmykS8IjoXvl
VU4AyJ8nsyuLB554YxfjvGyG2vTh+oe/IV0En9iGsYQp/1ClPoEQsy/e31CIZt6OMnixkQrycePp
TsgRX9Jz4m7T4MzPg8wWDZKN3YsLeRlyINB2KrgNvb0EsIR4juW2wUhPnG0cdq7Gdi1XUoFM1kOM
X36OBHJDQ0IYXoInR24Yql83hxPEKMov5+LbTYvTzcBvogoVu6z3DDapRA+8qY13Ni63Ln8Izzha
+EMOy6hP222NU9W+GvTGoyE0LBTELArPyV5rS6ISr+f7gB++A+1tbXsXkzbzSV6YQmlV2i7jbjHB
Fdmb4D2PFCgU2uqRWLh/OExgM1ZxGvBv8KBxJ0RgJKxRIfr/rPdHbyoY/QWn5sWnDObLWJHL1Hn+
5QYXf1DG17K55N5ysmvyrIBSVBDN9bsEtA7wqSAwkiAGEKIxxP31Vq2iOnIadiWbxaVZ+j/NO312
XOXCJLE4Vs/sckQ56KSXgz5ZMNSuQDN74YY/KY5lBQL1GOI6yqRIxEhMLkeQScmpovYurloRfsEA
AtjFiHL/up/Pu6odcP49o8XQKtIgBymEuOTQv3uRL42jWoRvfJm4RMpus6KoyYDyL0mrxwa6rmta
m0Wy07uNSJrISlZbDr/fQkqnEomuAaOk/o32eXACER5YJN7GRYk0oGn9AoZLSMN7TfveIRcJAN2J
eczx9ViNd/SZ3YlxYaC4Y1Oe1WYk/bgzrg564KkmnH7XNoOgMEcVGtILnyMS8bRVMw50wESkedYq
x2SegIZV3JidQoVz/ojM1hL/CZxxWkAv/DUJFGm5SGaFXAzHEOOZ5oYsguhihJLxWjICneIHvNrk
Kkbe6dzlIe9aB6L++loDLYz6HdcxcaDXR3RVS9XLEQbZmay4CoIyL003AFoUpKz7OP+HrgoHc2oL
Q64ev1Tz7o5OImyx6PBBDdmzV80hz55y5Blbn0+ZoC2us+yqvhX9G6kvsX4/j/KDEYncbPoEjmT9
wydUe1fBXiJ+zYFk7fHAVxmFANYBUhtFwfEvU1iJzLiT65sTZxo26pIN2wrNLV2iDOehmUPBixiO
H9QQqSXPzBG/tGIYspbHTG8IzybaeUir+8ZPIN/0WN/86e65CS3Kam0xQ3ogDzSKxFUDnH5hcCha
mM25qfKZBJI45+PSF/QZGWtuoNU6VD0fMEfal2tX/xfUFBtYH9Bjno4bnhYuEDRwFNciLDD1mjUg
uo9UmsVQAORCfhblVS3fJfHfpxdh/8QmMFFN01hYghc7F9KKOk+oTrC7+pZV2WMZdHUjpFa8bhbU
v+ViLvfj4yDQOv0WTZO5ZH3N9q5PgC8S/ee8nb64OpZ4A2opxZwtuWKPmt4ej75DkenK7V5WhL66
B80RK1By+SqQ8gCLdvvYiIZaIc1FtMqIAnAm1hW0fei2I+j7Ig/f7Ja9Rtuc/BxNmGYesFK1ji8Q
3eLdOHPKaE//pPe7yKuOe7UteU29d3yCfm0QE7WxWEJSVTxPECPymuhuERwJI12VeW04Rp/ccjKX
m8vrcNzpdJjLACSsJKJe5WY+WBu9HDJBbdUYc0OPdm9Jy9bKbG9eCqo2RV6/HIHxmDwU53imWnHR
NFbz3sWlYMKym0/Ui1V23L5025umNPCiCxqDOumrSEH1oKCNJe+Zz/cV4gPdWACuOb/jJivkc1a+
JktzLkGLm9LAHz6ETVgeZEIpLPD2yXTHXOsKIREd+2oMsh4iKwz+hBSuJNZltDHLONwyTnZo0RqE
XHYpw4qgf5nciNq4GmOQPfl2w9Red9ODPkiCdgGV8m83kX2S2awXwlBnuscXGp5nFtuP+tjEZeXI
+OvsbeYbopKM4MoG3i9hfCTxqEsKdfVTae1+FWQiGct4kwjICvSaerKoa+ovvdZYjKgPj+Vae2Se
p5/y/Sg/oZks3/1DpWAxx2E54L7uKjgIfL8b4GGevKBgexGbNR93VYrGqmAIcbbk96TJR1sD2Y4+
WR0iTXzeWKvJrhxDJY4xunvoy2xwVoPjI8GP+ttd7UP8VMD3GLzN1lRMOQEowYBuVSNsm6Dbt+2g
Pilg9U2HUsbGI0GRXx6NsWz/TU26sLklSjOXi8RaAAvPIC90/tvRJwYJLfh4yMdUnwydnvlXwmZX
az9HsvYV4T1SjfdHWLNwIevJsAku0matHPkNczQNotyi83EkEWssOoAZVjohTNez2s2v2Oti6VSi
gnBLHqd1l231B1GtUFj8BFIPDziyCHxlW6pP56oLZM5w46uwVFhPFrkqH8m8djlp1kEhYPJujb/8
tWVUrrxempb+S5qRfzM+IkOXAsjkWznyaeiHHlU0RMrGsspLB2fVrq/QVRPGzSYZYF9at1ozgG1a
rhxoDhYe7uw/uVJ03aCPw3HlhWCoo9/ckHBqm5k1Z1+C35cMRIvL8tuJd2JrExbIJrLmb5Hcm4J8
G8OQqgToHteZ4QDywSzKo//vSc8NsQyELCWO3CXxRvLc/pbD3nfd2lvhbcAq9J7JgQcOe+UDlN1J
DfEGvtDQ7d1aD6BjeoD0Uw9YQQVBxrHY4jypbgFGKGJ/IGoEU/dDN7hRMk2LY7pabZhA1t14eMxi
9b1lYShs/EkKW75iah7HGMQOsMK2Vgm4oFR42o1ZGaWZtcxHeHaoem5qgRZI8Oba5DA1fX7m3Zp0
4TQ9A25CypHRQ0x15W9Rznwu57m4b/FVxq1OQbjIjg3aElmyewiTFr9p70Rv4EaO6YW2N8v8rLtd
MRQ+nXrfw+BhKreL+8sy/ZMGXs3rGxpm2tpqslfnhlPys6Cch8hFN4aDfKyDpdQTP1KpDeOIqhdd
n/D6ZieDN5inkvXCWcyONnUb+dZhb+aDrUxpN3OJHeQZz+uGW/VC+0Pgd/zSpaExNMOUkuE5zoVj
umHQKITvhp8Aveq2V5r93uyF8N+dRzXYUkbbB8vCSowXcRD+nW08P9D/a1gPIPM2CcBByJfntIZ6
Ud2y3ZTjuDvoTVkzHNS3+hNIVbJWk7ZPoWhNozNw2ediyFA5oBCdT18tH0JgwylABkdkN9fy7zMk
QZZClgptSttgPTpTpzVAsfafvJIyqKZOkGx97UIr0v6yoY7GDrK35woSAXA6IE/xqg6TvJYoqHlw
g41OyCKsyMLmKkaPShUr3P0D2ILUJs4YdN7tMqCMzz2vPpupsSJ6AuGclF4jzBW1qmPl3UtwEiLK
t4dbJz4JdshRIJrnULieMDd4l+TID1TYENVpFH1bK3cUGKthyNg3bFnOW06QAkFyOrI1IMUO75b0
w3Ez3kaDrWWONaVSSwrlyd7rUaluG2lPFvqNLFxKAIMXD9h5KA84Eck62+6ZHJSTvmTtqQ9216kJ
ls9SbJ+V1xcV1pjgWDh6umq5PdgKNpbIpx2Que4naAzIY1G+Rr23aTj7RsN2Knij7PW9fxjUJQRt
6WfV6yeuA0YwsFAgoBjqszQThbjxiDz02jC2XoE7qzBk4cb5lnFLtzRkrojgFtnC9v3uifUVQzcV
NDUUl5Jph1na/FmWspes+4mi+L8x00qZugin82V6iRHT4PAbdzjcc5Kl2/jUk0/3TQVXh7oQHex0
vPk14e96GhNsVzuarRRHEqdc1c0KdeLDpLb239ieqBz8Nj7GqnYVMDblYCd8VBONTpgdZjLsXrqA
uz+RKjKbBfVHWzBO6l5KwPmlTs6cSWUNr0lrXOovc2eFpugSGrZuQr1+sSNV75bkuS0OVMXaP4T8
ECzJyHq75vIY+0zziWlp8uFac9jBpM34JVPD89/tYhkph+gWfGUimQtIZxF+sPLMfiNlBaxCNJSP
/pKIGmFNPhs2lhl73819QCejv4LlD4rcVRX7UtNN1Mj0VXJYKkBYC62SDW1JsUmdy8NiWKqJt3Yo
wuJasNB91fDlg+qo+2B0E+yhiyZAyUePmKC1gDfThZlMhPNNq1/IUmBIe1OZyy4z6Uh5nzJUBdoh
7jOHN+QN5AIlQ79d2QDIQVfcfXyJ620LNzDLo315fN0rBFzZ9CayDapy3VCfNHINEju4vzoh2zY9
51iS5PlnogNz3EezmJQkBuc4/oZlhT9A2JWzQiGuXQPXkpwc3KlrwaXnO7MO2D5XqY9qlQWpT8Xm
clNanQnYgXV/T5wI7R+xtn0NUAnvCOxcDUNy542IGTxIj7iqqBcfQm0LKO6cy83JcdxFah75qzBb
i7oxRKrfWlJf0GMeJEtJUUysPtB1cU1iy6686sz5+igQ1l55IQqRoiy0mMMbo1jNDXhUHEWKKQKx
aryOAqW6Qn6G6PI1sEKGi+4xJsdHvRNtCDyDOELIKVN7rBTP/Zl6MQLuuI/DWIAMQS6SDFVX9sDL
F1cAD2GQjavfA/Af3d6QE5mwZt18Rzlr9UQkP4UW9b5LTPtai17Mof4memT7Z9wwEO12S2IMQUVf
YQLTIzIPmU6mibXrRoD7SQbigppafPqLXWYxwFdm6KZWCQgJ1swIAcAlkNTMCRnVryg/YKGK6yFP
zGc1xICK1x4+heh4NEmtQotSLw/s26o5T5a29s4Ou5ybs9NhW61tbdlYs+i7IG4gdwN2M5AVLJsQ
Jb2fCuVyO/0EWk+h2weg/7JScMVKFF4iSRo4ueyWlYCDdQZsBdUnbbKj31IdVNLH2zAph/2d/pca
Y143EYDbgkVVahpnDQb2W8HTw9b6WYMUUI4UsMi2jiKka+zWxzM8zEF6ORVzkI0VDSO1D2JXrO3L
W6tsjviMmdUPRm6fmwHS7m/2lZ/U+aj0RwXMorI83DVIyr2PYi+LWwI2vPCu/IWoB1z7tS8uw6L7
J4zX6RKav/gSowpwfyKTWqukZKgk0gMNg0vJqPXXWLBeVyi2ZPbEO44EGGiSk5yhjlTCmJCvdKiG
9j05QRcLyb6+2UHHygRBs3iy8MwG1Jqbu4J8kBWuGz3qhxU4dghgi9G9hJQB3Dmtza2J6RZ/DKlu
qD8L+Ib4oL3uP0I9Jgv83fjUE2pIBCZSqQKVPyP0I1O5nGlvnBp/sLtaHVJSUQJwM+6841M4RNry
PWVczM4nARLxQkFPHGzUcsXrJa5OOXoCS8l084u81QRN4tFf8m0+O7vksS2dF+8Qc5AV1NL1s0CQ
LsYayxMQr5vu6yz9pdaqMtc5a5YfDjN3F/LGd3AzCaEH66R0xRMefX/c2215DQ/DTKJedQPlLVzh
7zwZ9PWMsIJ5IOn96d1fej5zfOkgjsfJ+ZdHuj3DjdObAp2J0tS7pbbXse65rJYTC+seJycz1KZi
47fj4zb3hUipD8lWSkrGJGCgE3I2440q7hajNwBgtFjb/Fb5dEyP3N4g36kcVHJAlfjmJLAJMU4H
+Db4Ch7AswN/1Hcg1XkfEdygBZdyiszzUqEVsRRmZMczwmMok8rm1W3gymVCGG1jlin4FRKYISqm
pZ5cEoy3K//44ASGERDoo9fH60NJQa46INs640tmhVQYPHyfg1EbTHct5sG9cQcHOrs3xHhCCpmV
jlp1Bp8zPK6KrKcrwKHk7I+rEgHsFvmgqc83kPQfqHRGjCI83DvFWqTFPFHUWN62x4a8IAsw4i/W
IbHTEG/YWY+qOeS0C7ZmOKtQ8Rp4vDdPa9DQlwP9Ufl0uJt/D7R12JnHjRksvkyfMu+jMHV5455f
RYgHGLrEFFCdcNo9YyUzbAoQxoh3b4ZYLESlVrwM7YhUV0jQgF1r1pYZ6JqR55SsqEaf5YLyjz1G
Up1a1uCxg6371ZMgQW+DQbbZ1LwOzao+w2dN4ny18qqyUFoA+9rBhiXMLVX57qHsWFI5W7jlPIHI
QeSx5iuA8qAmfqEIXYV8L0goJb1tmEQIKJ0ivDPnh4ikwtsbtxA33trUv4QkXUpSvnQKCYinRP6X
X3Q7cchSQzApyra4rtJvTfkk439y/NoaUgLgKMX3ar+QbFjnfWo53EokNOqSnL44kItwMqfM4tOr
SBd5Nfsd/GZ2Xgao7KOTCu9vkYT3N9176reB3UGdRDgih5Ae4U+sZzfzCEqI0epv15ZUYSUzx/ZN
D9ipOpYyL4KyWvPZEmbMKmbq4o2nrE9s7Y6z5dd/HR283L1SXSCcnUzIT8h7OAFZE9qRgU1w7J1I
qdkSzpSn/YTOKPhoxC1xZddnO4U1nurbikT0CGoCShE/6xCfqPOOSQ9VYecJPfRC+ZZW6hCFRbbv
VzwKhYGyNgx9EFOUZi07wK8xS0lzSyc6p65+nGDV0j1zWL4xdXvtVr5NVD4QO7PnQ5fr9hN/PBqU
wRgBZmZX4JsT1inZbnnpjai4joe4s9tGH67Mz7tzxjvzmbJrJbZFLKO0uUXZd0yksV+kmkhoEwq5
ISZG7+9PG5WpQdERnIYjb+tfm2sF3yQH0t4DbTWIRyyVCWL8uoQLGYwlwczi1PJ1/bLJBE8uRaR7
b/5ReLcXDbShN7kkAd5EmbWF9dEwknSj67tUt0F6/+tor0gaIJnPq9KefZ10awTsHOZLXmIEULy1
xY2VOHauE0K7aw7sLdn0ZslF7lUw4a1R6WrnAt3lZNuf0s4oxQe0tGPfN8PREJCIqfYyMQs6UMoB
iaL42ZbAU8Q67bPSRrJS08XFYIFpM2r4vBuAFpFFbB7hTn8jJa9BnWSvGxF8aasTGVM6Nm3JrxKl
tT9djCoIYm2uG1k0oLEPlr3k4+l5h87Cf/NGMQ+jU7ezVhgUkVqCYw8h4iKK4KRxFFk75pgGdxgC
CaiX7kLr4yG9t0z3EyXjHcR5MfocU0mkEV5Vxis2ktIxs3I9ZBQdk0bm5SgMrlyxswCxNNpnSe/Q
rdy/4trtkoCJ+hZsESsjBKvrFBAQtTAaD9XTlUA3lWwTZjj7J/LkCrPTsBUH2I2W6WPhse1npXNJ
lQbttBEq7xj7wtFCWqvDq1z8SeTYoiexvOWeAPyywYNOsUAUDdb3kVsV4tqUVyyDgpx/idUerLCo
ESDFWpmwNJeiolFUS4kb5i92hnufCk+ge3fHKWqVqIsJE5xt+rnQgFcXrPUczedHUR3haU1B0hbo
PyOLZxToqkg4PfwhWOHUTswCkMJYNu5noDH4atfGAaz0mYRvXguryxAagrYmu/dLijc/JPufGs0P
JIyKmJibLw2c32c2CvBL+aPdeCXZagcgDXRxDOpBLJCqBzVFTMFUjOcPuVfYeRhoI8+TwfSjv8Dv
SNYay0nQCFemq1tc4jF07d2Y4gUQiBolc6UdhGNaO8zg/fdtnSLuukIZNlbhbYcdNfoCDa6FTZaa
CJknFciriLgVaSsvkGJZy8hD64tCgrWrJoOzovRZ4af/5X05bj5aVtSWbdJxGljURDRLPPXDo/4+
4fPzZvRbQUqhykCSpb7Y5R9a6/pCBXpehjPkteF+IlSKw8AG8deA8mx1Es4ncEnbjGAM21tlawsc
jA+5z7kUMp0zAGZBKCbo77OX5pqtZ26Mbc49RYmsLZy8ZZqBLT0dfd3iGDLQa+sOBnYjwJHnzPQO
UvLT5CKNoemTKAUf9ZGXWARXJrOwn9n0hVJZHUF4CTwG5S3NRwhgH1PgrhrTlK6MvdSP1H3huF2N
3iIaQXAMYSTjIJaGJPHbm1TboFom+lbbaC1KzB84tvSCGo0TgFoqmJbsYlQ1o3yn1Nxkh4G1jc+Z
M3dMdmiJPXDWqVRP5v8Fs/Pvh9y2Jj67g/kozW6GxrIiuF3Gnc52P3WToOb87Yfab+j2GbfyYEy4
cjtzQU7pKFEPjaPMIFHl/ChRVgrdaoMr9cvnteqCiuAc3iPUPmhkoaAkIy+NnA8yu4GiO+W3q7Qh
OpPRiLd2FiLJew5qqvbeJ/A9lL9Croja+Kf/iuas1VbrXf3lZmcZEO5wesU8Z5ikcfgwi+LxT8dh
GDYGaZdFMLJ7+01qZU6z3JzbJBFhzfJ38RjML/FwmrzZFQViTkEPJrg558IkdpxzEpdv9zQF28X+
lCIHknPx88+iwCq+P1/k/HsWtw1nlicPYqGxjyLee8aVk/y6/Wi/jaO43upezJt2ecY6MirxXo2q
vuVwZ5HPNtugjxR3L4rb1RGbRRWa/tM7snDnaI62RlPjonZdFeZqnkEYMPQXMHAlv/B5sniBUV96
Vgfnr2HSU0Klnk9ZWZx5pHsAOuV0ND4qwFlRDQkR/p1CqXdEIVNwDRepfR8ji7a4sygTCkSng5VJ
+eFt0zyHdYCQdxeMqdf34ZhTF8//Ss7dS980Ticj+jeEGDSygD9yXCV8Ju+lnFcCt9E1aPs1Nt3N
6Ocuz42ycrWLtGf5q3S/1WEUusDg1wGSpfqiXc7l8+ER4GoZLJbeH2fHu7g49R08KSEbZzTgEwTq
oxTRyIYZttHnWyzFJFMll5gjSR4xWMDzeBTEj1jQQkUzkGryaKjsdpHjShe8K/BThi3GB3NXMa++
TpvViCOlbjOqoYH5BENFNxmEbt6XGfzZZB+TrH/u58m/L2v6ElXR4U6UT0xwDtYjCaxJV2RzWlhO
4dMh9NjekldVg9bZqY41sA/LH5d5Y7v81CJDz9m3LuRuJqIGDVVJSE7Kx9uLrAS9b0HrdRmhlcci
5H8ZgA/SkLlg1D9HLUGu4RNifBi+i+kd0zo5ZkZ/54u3RxU3UVP2C+D6WBUBYrQZh7euRQ8uV6YU
AM+bg+THm56kkCWFd4Jt5g245tOTt3Cx5yLSi+dIUG5JkRDtnFR6LonKU7n+0xJ83M47Ja74h7LV
eLIzUoByN2q7KShJEoPH3Ct7z6b7mlvscR9elX3b6Aq+x+fwgEfI7h1j+BFCX+uRyZ2gzexPsEzs
uZMk/6/vwJhaZqOvsC7x5GkMuPGgy9SH/+G7NrXcs80OLf6G78p0QQEcwAcKGr2sxDpZcJDPxRG6
wZ01pJxvuL2t0xWCZO+wUuvPLVMbA69IyWKiDe1Kc6XAmxUSbGI7qbzhT892icg1cIa7WBlodgN4
Wo8Cd1Gc7Bq6tWr6tcPyQabduYizzuskpmJfqgI7XEVs8td4w3p2IYgxDGQC+vQ5KIsa9bRV6YVh
ojZzExdrPKwRYj4bXo1RNeAB0IDckclHbIZTgMMh5hBJqh0yEWvqJs8aZ1IqwWnadF/ZpUqR6Sna
gvKtpuXCbeq8OrGQQAXwXw7UVLHcbygCKMqLNcaRxnKW8b3i5F2hk9y1GFGBxIavujzg2eesxD0Y
WMNHx/FNht3x5mmWLdWpCtXkR93Z+JN+AhvU4fXa77k2rlAXSyKWdRAEYvZW6lwxcrlFTM44N7PR
DahwejxM7LmtnBzFc4Tg8TyrE5fzhR+wVyGjWsPBeOBRnmT523EBtGUvJ+o6trvX4rxjtOp8ug2Y
97G60gqarMNQKYPOPVuFei38ORlxIz6PeUUY0/7l6KkgjBjkXx7F3z65/dTkIhJb1eizsYdAcGj+
Aa8wYCDb0puol/OazJEWyu1ZQH5FVm8/O4RYwXlPhbKFhB49kr6/ljO8A6EP7oXzMsIcUuXaQlZF
I52OVBfrcc31uxOqWjP5N2yP7n8QVmJtFFEWf4RI/O9tKszRjL/g2Jjs26uA2EXHbAaRbjAWda5X
k1uUo1Y38VB3ZzkGE4mLckyhGbLAa0i3GcoBVxOAwAHtQf8dqiVvqJKxizoO1iOe3fqsuerz2yGd
A4DI7DhyXBAl1/AAud0oD/9QIdeUeSf/R2D822XX7u3ebzCTVI/DqsAYYyEDt4MDPdzQ8stwJwJ/
EuEw49cztH3eQiTl6TK15YAaEXpQA3w00sniJOQwz8lYv1tLfFwF9W8wbM0AWjTLVAkBIM1oh+yf
Bovp/55U6TYJozhasOMs5lDm4rJgluG8yGW+uZ40k/2PVGniclaPU6cH78IKG3P8x/1WJsizQlgC
3AIAeDhxH/qvNxEATMJtD/lubaUYQNhzEffjXSt1Yu2VgC3XVH9jGbGk60/VuyGPHy4rDLLmB6S7
d5hOZp/aC7ze7UnI5XLTs3gjNA9ogqYmyRzHgG4TPHyHsamBbP3hiNqGR7q8vUIYtadspIyQoCh9
hmD5hVopCMlGCZxo+8Bj7foMYXUs9H7HjC81g2IVK4PGJXmWXHkmgIyheHH90eEwg62sCHVPWrxZ
VzjPQg9k7jFvgdZDo3dd3i4xjD67HHBku91z4lHoaLitNK3JW4OdAU81LtzXN9sKlYfczQjMMTRm
5a4zHJpwqxQQeipNUEod7gDKmCMEpTcu3f+D6nbp9/aGKYyWZ1+2UMCudnik6wtJM23zkMwbW7r/
MpRQNlfIRW4fkz9/1SqtqPxiP0K7GAH2Fvw2UWnWwkvUIzCu9hbOc9jOiKXXFB6weH2e4ZeV1f/I
LYEE1bWtju+HJfNzJFXe2ZXACT14V7Q61iyU0E4lk7ke4QtDVRCqg31vP2lFG+oy6iZkoNsMwJ4E
V/cIxMGP0MJMRdrUCYNY7FqMR9/fW+MUTUn486smPiGy3nGTjOler67Gf5xygNcojlYehMR6Ofom
p9rroEgQY1UyCo6T2MSCCfOFXn6O948jBJ25YNyI7sM4ueCf5BXLNAIteYsfmEbEnQyuIc6R6Ks4
7LZ5lnQEv5rE10u/XN1tI5kaY5y1DV9YYb4tvtmMHqNclSm0hYhjMkRtn/KFYc91wNhSXEa1Ftpy
XZQiIjABWzVwKBQ3hoT6fHyzEZnZphVS//k3ZpzsPTOrbGr4hETpZk6cgrZE7l+wypLxyg0j5p5n
tdyNWAE1EgieS5abTu2jYQmP9rjC11sA4La42sHyWzmvDhI1EGMW9W6gblT7Cm6J++hFcc3ugpeD
2Jmr8FaxWfWy9f+Wgd4RQkEED0Ld2LJ6YB0abJdag/XTSnrYrV7rUS8Ex1CNFfVFo4bYtHMHN5mM
OcYA+HJBuMVBdO1DzktScPXSJlGT4g2z0KDP5ZjmIcYSH6BFt3CuuFQPaScKA6qZiZUMU8oB32fF
3sg9SSLkuN+FC3ksrxoUUM5Dk8FNlJtutmOJ2BQYQ5vFhI350iv11+3Mce4Vdm7D58TJyaBc9y98
vMgptvGmAnyo+uRWIGlaXDVshOme96Fnkxh8/EDLtXA9hacD7RzevdASDlEVYAFAX3pT+S/B54yM
NS+ep++S2l7C41hig8a0+FMf+fm9IDYGMnUE4eRvCTR5i74Ya2L5m2tDuA64pJqRiaafAwDxMXfM
fSgsCh7/+0AvD5DertJe4fSV4QjVnAa5NMsCNsXtBAzaqT+wQvNn8cLkf+BKId8vt2mDSikDklN2
WcJpI4Y4+bzmIrWhysFbZN5wtE3wtFvdCgYYwPMmU0Bdszr/mNWBLor8j4iAunfdpqlV7lEHKARR
bsIrPgFz/hxrQeAmDL5MyzGuCwArXSFpLyxvzLeXF7XnmA75ZPFcFsQRvNEcRxd5PWFRDigkHUj5
dzy1PtNK72LEqh6BseeDoreLRgd+/kQQrFOz4eXkK4StfIjnIjsRSbGeaLMZwkUBCdXWG8R4XqIY
GaHs9aB/aqmCXEWhF7GOfBi1MmicEtd3umEVFVnIvc6ZiBHZQ2p1i1pqwGK04sf6FGQL0onnLZVu
OeVhSgalzKoDWh1VYKV4yTcRF/6QGL+4nKSOckGr9qnKCukP1/ahsijnbU7pQ9jYh2vL7AWYJ9Lo
OeytWVkdkZonqXAUjYrZdpDD06m7Z+RDGsoGulmOtXNFJt4THaDen1asbjuqt+vAuJssa9pYihZB
WAb2uKrdJT0LSpw3/FrzVl4ecOfT7YLIOrItrhP5m6SSftaRgo8eska9DYDxLlY+aLvXmZncFCLS
ttVLhA/0i8cDYOrFHTuQ7nvFJmklmf8HlgSvEw1xASdpam/3dq/5r+NAQ+5lDm3dQd2dOtLJ0Slb
CeH/CbJH0xT66KDCftogSK46TS///j2TxuTEANS2uo5okCWzNrraCOFc1WP+RrA6p4Jl8nMz4z+4
fREgJkBXMQeZqwrCkqmN/qUssNSXES+59lXX3vjqkpUQbPW6WUOP4hcSV8cd0gXTgn6Fl/DSoDyP
TPmWdVm3MC/OZHl6he5DyFVctIkuIFsST6EmMJ8mjDONb0YJsVGDmxai1MAl+mvn9JmRZ7c43796
S2psbEX2zLrlfvn8ujdMnwJ4CTWv7P5UF61qBWlPdTdxdx8eJIrgygJnpj1/NZqD+aQVbApZQzC6
wLXj6gaB26hH76icJ2T1afAfYun/wdbI8t+1Ygnli6V/2iwpwYFgYS7g81VyDuv2IQAzpZNykyUv
hIVIxAiH/fNvS/m7topjqdXKzyQ7Y3vjYAu9hfHrcWDiagKbKdk/cV4ue5SnoYYwpJo8Sjcawxmj
AihLoEc75bqazc00oCRb0m8fVi/RndWV5An6dyj3txRu7mlVWwab2SpLMr/ZqTLjoQfb9SJtFmog
I7Ogw0mbz3a1wqOOpkA37MH458Mts3o1GFEE7mdMurycBnN2aCq2fAIrQxnYxc+RqV6F1+7ZdXV2
8MM8hQbz8e95OGdoemKjvB6NS2AimuYnGYR8SKAs1PFiSBYMbtJw2jMg4eH4sLa19ID3HiYd7cRu
+xrEG3o/Sdik9EmHUH7a5y1Fk8yAJkoJdNgSqcaoAcgw1Swrlgepnyn/UbVBzlGAfpu2X3X1kwnV
Ub2jyd+aIF0/Y1Pnb6AOXFa51D0ooPZAnl5r8pNKWNiOMJa2Dg+ri3EaYTvF0MKz289/86raQeGz
5rJq0hjEPif3aW0nZSdC8L225wQgFtoxDLIwJHyEUmMe5V92RlSQQVhs6D8fb4Q6tOhTZj4kI0EB
buiuHukG4FWR1VBZ91KGHmgX+hNh02SJWlP4QixnfvJv+tyiNi2qNsSh9RCF2jupNa3gnA0XdQwR
UtKARLkV2Erw3Sx15z5QhS2qwTxyQar/EhXrw2ECQNKFkBx3WgBSpWNTdp9/SMrl7hXyJQnYptfP
+t6b3nfS0bR0pxSjL8BSHaWZqfkKz8aSaE16qPTbpQgjGhGak7/846ufU9QTx3lITWcRTNAVhOxX
HSFzYDdUQ3ZIC+36aFr+fpHZN/Xu50dBH9aZd/hwNyQGjLyYiAqB9H5Uz8OAyDrC1DSo80hIX1Ni
gGekoras52Nti37TvxLpHWAQwKz+xL6BZxS9T3LhP43WyaweT3DKk+UJzOak/JBv2J3U9C7E/jlz
HP5NsGRlA2G/ne85skBBXq8A9fLkzkljOLR3C2x5iw00f9NgR+fK38//MMTjXySrYRLsngOFIuB7
9ccHnxQ49v7Dq4QDsLYLkOX7aF2SmSZIjNWeZ0HS4gvTQpRsOXkUndVs9nSQIHy+jPrRW3szW8+f
BA8zLLLUhrIIGfoydnNcJnH0LoaX2RzxeOIS0cMHmmzm8r2XvF0N68tqBJIQ4DhR9hSuXtfCdYTC
Egae3s43YctZlYj+Ur072fxrFmvKwTWctMiy54LU+VVSIT1ix4kzj96Uxsw8jnGSpchL+WaYAcTz
qVlrIeve4gOoBnhl4emp1cJ2j9sZP7+QiPrVqmxLAIQDNfhDCwNrJe8UBd5yv5pSq0mA6jPnclIV
Rx3aVQ64X7T/KchCgEbhQLOAh1YQeZfpJKwYayS7kOrwX12QkKYa7yXjSH0P9hO4QEz1eJ+y3k1j
Phcl49Lp3jXTxTsHhrJxuL/HTGcyNAYrOSZFnqIGEwz9CvAmI6m1Ae8g+qOA09zye56MKsRXiFZx
hngTdH4bOamc2MREcwG6UaHigFjB5i4OBPsVjYJVNfM+mS86MzyymYyU1aeV6OZD4MicjYPce3aK
neFzvWDsZGdCerq8EFv6Rsq0kNuk5Z4k7nc7I4JEIa+0zNrpDsGwlZyDhzy0IwyZ6GutidFTns9f
C3fH02Lh66b9OM+kUT/wmAfeiaqPfM0AsHATtxNSBWtpR37Qi7DFgg+5jPP3mmhN7+kXAEkcz0LL
cWgo9Akqh/agSEUC0D5d0ch85LqMqVyWLvtNi0wyVvts7ojVpmw7K/3ntpoc995tjhp+AN9gCj6E
o85u7SVDb93niuxwb5NbneO+d95NPUUE3gXxhkfO0N88MBupUAoUtIdfpqrAWEgiikzGG3Z2ji43
Wn8hc8QpWmWJ605Q9GIBsxRp/TAswbX2488gqciyWi76gjsdmg1ZFmXW93XkDYp5vL9FGfB7Em+s
W7DtIqs35swBH5ltFKJWuq6T3UPsCPAAApC1kqHiPfqxksnn4Avhu2CR1V8htH0g9ojrPNeNvWCW
cDCGkhNh/2ZQe5OqnMrtwt4kc+WBvAK6TOyhSNk0qTXjnNlbqQa/ZZ1tbzsGtDgujG03vSaA8IV1
H6Z1DTehpvaqgRP//9GG3btdlk9/YwBrUw2/ENXc/jnKKZd8KIXPqydJDagBBar/7DcjKes5nKEN
mjQTjAv17Rc5A9J9GmiS8ZJrUvLjnku404XXjbanHOwnhewtRDSn50eEyUwCzVCe70yQwKza0szf
2Yw1BTdzlENbJ6TjalffV2sZshY0GcL0NIcaiF2dSF6Ro6qup59c5M/COWcY/FMjI3s+7xFbcrsW
Zdw8IQzADUAzbztad4v3yOsIrXS4TRwIqLlGg8k8t/bctJRwIUxEpN0UsPswuEjQR8wNipzeTBHN
+atIMcTFnTo7kwVreTlNavu3eaTnM6Yf2vTD7/WYqKalEfdC8aYX3MIUDvlZPEZSUNljb+c1emD9
fbi64yQ/3pKlP/yoIlNJvRQQo+cRIVR3M5JJYWY6TdeUXr554QyWWs1XJ09W3RxvXYHnuHnax/xS
WduT+3EFY1y3NfoWWCQBsGCB/4gUU/XwfMkNsEleaVkiIR1KUP9yoteyPTqAV5aGH+NSfTk25iX5
lMoBsCT84ijC0tZ327D3CXSYRx2dFzCrJz12ooBosld2tIYL2WDttoaikTKPBB1+kh85JRV8oBBi
NJ08npx8wpVtPic0UmaqtmD2Z/FNWENHNMulhBVWcU5LwmsjMkLEytW86Cu6tQuC/eqtMKgoiTtD
EptLc2PhZhy0wt5SiXqZ94irkZvdkTorFQyjVb8dWXgL5i/3BTXZdh2Dqw0MCvJUa8Ssf7CcNfcW
j3jMIhnZ+5fuW1Y2fUtYOhPtxD259N6x+VfFRrPlrF64c4LeC3fAh/Q1HX9jkwfRPBnHppbfzpat
KOl/8matIDqLLa17392y5h8izDYho0fGaDqpb8PlfkRvSIYQYIgpBhpg/QWfa0N5AnBQmh+JuFN0
DS010lb+/snZrgY3aNX6sCE8ilBIyDqmSJkofSxEMPaYKp3No01J60ZIky+l3aN16fVccWyGGXzm
gh5bpLDTr7isUZcz6+3BvMsszrWQXqMcVGPlC12XPgWHOPu1GT8m5soYtWyMpy407kEPc6Qcr30m
nDmwSL3ITk7tcWwSxXDdmjw9qnn7WDf/dmK9PDdvx3taf5cBrF1BmQ6zynx72FamJlsZlfcPB8lw
0qfIX1UTKwdVirfuRUP5/6qIUl0VTJetXZtot/SK2bNQbV+f6nPbcg1WClBnfiZlkLdymwqM7l7a
dIyxYGLou9ADFa5aiq28ldKJ8R5XMowLDYs5pCOT4PInUltCJ7p6h0eJk1UY5DdFrIHJOE7gT6C0
7kOxBqIM/SPxSdwoT4sj5nkaiuCYFJNxYWZ8PiWjzToVIPU97vnxhgqidk33HlRsF9W1BTfGy3q6
ZdlPO1XV53ExW9c5FQRaUsIOh9LhJIHJtOAlRDfOw3VbCVIXh9G4X4EHCRmtYSmoELjWVgJXAJBb
zTPGvCpuOyuMjQdV+idP3Ai5XD60ytruN0aIvI2e3BO/PO/JklrCnUgj/ScVbN8n799EJTpwfIIx
lFAbbb9OewFhvPvEw7sGFRkJEdPJwr8U7qRElZT8pUQDXzw2I+WyicxCmZUqVbLonZQzpkFFbvjO
n4moQKC0GnLKRKFBxNARSGpqRtYOo3clRgsdNhw1AG+jD3SfsQAwrM/NdLUy17wPyyJKTwMBDp9q
UQEOFB86ZDnS+ju3fBSGI/JuKDRn/yEKtThNYBJVAtLu5kCzl3iYVVmIr3DhgaDcwU4vKycVDfhD
2VovGst/uWH7GOb4kusNUd+DRmHw67nelHgIiA/CO2VG5LHFSEXkgGaaBxq7/3HJlhXnNYUZicsp
6IN0lY65KG+4ssD9q90a2POI1Pv3t6Y6Az+3wrQKPBv07AZU9Ghq9w9FUzc1KWxtqIZgJ9zJ68xA
dqCACc4x3LWnSb/2Dzv8FKJbdaQzvMGqy+MVjVqPFdNKoSvH1ekvyKJdkUGMnb2brK8gvhCA6cRO
S2ducY8071vQvkZXB9oNX+4vHf2JTmubn9/YdsYSDlMo2+56hMzAM+I/ITauvSIT2LhaYDNvAli/
uMyODTejwsTg0+rSLfcViPm19yEIF+zU+hzBQGb2UH61Z7bGnDYFi2CuvFIU+KPWXNGXatFb8Wcp
/qL6L6z0arzBggcgd+RIJ5O5GsT48YWPqZsrR7yIEQ+LkbaX15EH3NYLVbknLEblByayqFyPUMq1
RGefdWIgzKW2ODnp5W3yAe21XSQs8KXfg08YkLJRZxSWryk6MHxjAE437Lvt8HP1zDoUWs49fOJg
B2euO5/zOf6OJuy6mHCAo4g60y3zCZheabovGDy1cjq0Qk4kXP4rzWzPmHDpaQh40N1mg655q3bO
fNH/WXzw49uSxwF0VVfpEjzIabG25QKImpJ1CJIgT299znD3dTfZA4astRovwZ1Go20HnuJsfcJM
RH4jDMIev2aNN8SH+i5D7HkrKt5c3rA2E+g/G0JUPuy6e7KcXM4RGUil8oGYrniPvltZ9oE6Sxxn
He8mlqtCMgVxUMj6FvqKAmKJr2fqKTG/shzm4KhkoiOChdLi3kIBZNtWAHO86YmMQM2yiznDDeQv
LHnZh4rX7YSi8pDh+tedersX1H/gjH2BRe6QJT5s2HEktS52/ArDl+HDzF4y2a6Fnslulmu5cd3K
dBfvQd6n49t5+g0TfhpPCHLbtQZQuc5iTI5KMHl4RrvnLPp2jxjgXcVmsLvRWQgpvF2LVSqI9O6V
BwFY09KqWVddgRCBWQfuulAE7aul6oonlSO+xDbCuotvHsAZVDco+8JetTfJ54oFg+9OqDf19KpC
JbDjIgW55G8esPpxN9OjsFUsZHHTEhweYnd/vSZQ38N4ucARKRfhI8+fJcEQDE8b1VVsBzvmHsyw
DkjEIp21e8Tcs+eS+mLgBTXuibGZUigGqNTek5f0/lvk8yDGZp9/nw6ngd4L8JRwqB6B6VMFR6sH
2Pldskx4AfbZ9z+yrLfcJWaMnGfwUOG9ECG/qIaqbIVzX+pBqKwZoib2Z6a3aamg0mhMqIQCsx9U
WT4sJ6Xsc4HFkRMkzMMnEl0IAlwEwxURo3OyrRYSZBU49wgwCxcI9j2x+hP/PgHLhSEMis0rC2k1
jyGTPesLlwakah72T0EzZbC4+xgjThRWkRnaXy2B2s9FLSZi9AsFwqjWTb+Tbx3Tn1uffSLkT73s
TGOABQRIS50yJyv3P7E+0kMcqXlf4Fl1bsBGJy1wyfacRwdjrptKFmiiLym9uXUI+hHKrrwRaD20
MV3imuj/HQAhwa/hGi7ljdwDmqPbnNcllzcX8gvCvtIMdSH1Q4zA/e/UaRGcM8zHlExD8kkCmFHI
VQ5ygMbYYJbt0kugOdK+htzShrQfM+LcM5Dr1F9nG9V+LTvsyPTHXkBhlYRLUL/zCv7rGERsPznb
e2lKtSgsuEaA08ZycIrBoFCFrbPjFX6mlRltzs0rWgv/nxo4x3iX7HafNJNgoRCWHogcoDDfQz/9
o06pJRjV8Cu+MSyT3V4U0/Y3rvX30GFiaprXs1o8gqozidyK1yFYjHsVKYgicjoUgzr9bEhItg5y
EkLyUz0Vf4/KfzaoHZZqVW1PkdXAua28gtt2SvKfZKlR3GeofqSTDpx5jEqUmtdrxZ/4ga0kQ68w
VEaDr6qWrS3N5P5uhVCB3vcDXAGBx8QnYfaN3lI+lZSMh7Xb+GgRUjaP0f85Xk6Dr8/jEEp3qyCF
xZMXGdlZjjWvKhPpE3VZkOA9sZ0BKqlqFqq7USzxbCzezvIsoTMzXHAxlmbvWkANEsccglchV/UT
2nKgtjyJnjfxzDvb7q8/l8epRmNFTmij4vTbXQECwdOlfWDtW9E81nxqq3V8AnOfjtigLcH7WlJ4
RfmTHx51Lt/uaRxqUau0NFlLA46YK1XtZnzOcOQOfzxd4HOuCvEa2s84f2b7glkPn1VD7acPmIXA
DoORhXbfEnkAbOZftcTIw3bsl1XyHtZCluD8NAWRrHOAvI0R6Q48R/UfEST/aXG2z1CVnAAO6eDO
iFCWQXgKjCj93dOLaVrtBAYF/70K4S2nfHDmirm0Vgtc5/SSbyEbqcNAhyJB4qTX+FzeMXZMYvUk
aar6mFCoWg1Y3j5RCkxGwxYaOkl4krQ7zcGmSgQ5xHDkNnvkHfDCFyOWN8yb6Lx/6z7GsN82ZHWz
bjIGEKaWVXxRSX5A4zwWsgAwu9VZpEHjySdfBaGPyJwPRU8Ze17muXr/c5Hr6ICmmLEjA29937HX
d41AQrVPMoZPf3EfMhg0lpuZJJvriLiFeOqkxc/02zx1UDFXM7LNpyLEeX4TZQofyEZ1+B/Oa0Lz
Ti1NYcn7NpQBW4k+PnIlFsiGBiv+DuHIiUO01bVmv06ciQA1zIF7jNIFzyZm6KcLy41ZGTXV7sIc
ljTzuJ6+eJykGJsFzW7y1m+R0MTdigjtlqUZH4wTRoZFLQsQAbKFBfYv5ZQt3xDE3Nx+0HmsFTjt
pn338WrlIrqPuU3tAljMjomUwRO3BqAEb82nR4Zg85NULXsQdNQrlVnPvX1SHDrr+rRQ3ZCDOG+G
uJxtHB8Qc3vLvJIS9WdXQRpbLumzrdgFj2GgTIkCGNOieekT5Kb49ftWz//d+Oco+x+chWIrjKNl
OJfM7ykTC3Cs1TqI8eZsPXU1RnARFflwcFtbsGuKefQQNL9VkWn0/AdHuhh+G4+vutu7dxgkSoay
B5t/Avc6c6aYfkcNrHr1F/Y3fMbqqrmh35fRBF8NwS7gyguT4KViodHWrkUn1TBLYo8ciPvegs7U
vTMd3rHYP8xdeiL2Gr49jBbx/4D+fyeJEvK6fAiQfxZdI02YxpceVZnGitvGkREyCPtBlZb0xEe/
wuuKgLt8RwGHEYqE1QmFZeKNCwEWPbeNddXi3LGvWjLVO+OOLEQj163dJcpGvEy78VurRtRbPCfI
Jd6yk9+3qLPEAsa37VorFsKlrlSOYCocbr9nsXDQpZ1byFKcL0MoEuZqhYnDng0T8VJaENdtDm8q
uMLVlb4Gp2shwySqhDOSXSB3/4c4Ua2Ex3UyqY4i3jwe26+0r/EpqGR/jrZy0FAoEKx0mn4wMqoV
5AgfhrPFl2kOpKUv4KT/prbHJRXfYzjoP9fpLM8CRIwo+K1ZiiEZd9vxOPU9mdhEzeKV/xQ3rY2e
ZAPNCUdXsDPiZZFMFDnuq1xJqJPhJSuha0rdqCGZ2bMJmo+9q7/F4cYGqphQtVNniKzem1WjQBhy
XRWZJ4vI0vPWaN6IdSMbbAvLzb4x0LCMwF2niFXn0FQzh+Bb93Ia6pBaNstRjK29gGTKd9XWY4h8
sW/3wNuAE3v/XN/68PlXP70BYMpHY69Ikbspe1T6N+7UkycZmLAvCpzmWXcrlk2yvzK1s92aClaW
Ktc0U3lTAvl0rEWqfN/VKUaTbJb2Z2PgrKNFTjZolK98IRm7xjs1yEx1x9JlM3FiFfAHtWIrVeYH
Ob0UfNeCsW+tXJpx++PCgLSUMjw0EUoW4KeX/FW+lsyyZpFSN0sAoJ/iElBHqRs2EEkRMME1xVL3
Zk/tDW5IBeexPSGJVDWr7q4QjjiHI+JHcjCRTbT73e9JEHXO9uEiln9TfmoGCx3tDGK2a/pWGvO6
UAH+tKffJlVW12KmgkzlLxSquVBjENSlxR/iHuyvN+YePtY9cR6KHVT/sHREoZ9WIOEbNYJ7/3SE
IeflMaJHxc2CqVAiWbrjaOpuEbsN0QQVnlZB5KaDvgZj2LTZU/4MyXVXq4muqbyqanXKFLtUwFRM
cHtEQA3GkEmFRx09cEEPDle6e+WJnzxPAmQzPlN5vx8fxuz/EEP7zT+MyURu3VejnD/3FQ59PTeU
3JYZ2xK4MLzE1iSdzWNazKCkHZOq0R5++fGCNQbZWMhc6HWtA6pzSAy82ktiocWRLd/vn1wBUa25
2kPBpjtM8g+ytMPoYVLIzqNEEGvNgjhH5b6AYcmNkI1yq0zNtUuga4Ux2lwCXfYOT59W64c6jIFe
ZPY/1D/dUdOz6Qj0jr1CKl6BmEugtFwlZoScZbTaDurpg7MVohAi+CkNKua/YY3ulQcH3PgzgOqM
KLsUgHdBffyvRHmeUepcpswQZheVOAJoyL64xeimV7/ujn+7OJFSCY5YnIbOg09D2hmx6nHhJQ1n
xBNb97hEAt2JiWUkhJeVA+Y/o5M++w9j2vLgLKc3DEQRRphaTBUwX6pTHruTj4uEJ4dVblWEotCh
KZnZBesuHhyrNdCBIL7IGEO22MWD64TG7kWYpheFg0evO6jT3V9LIhAClZgRv22TaxpouTxnfgvE
yJjPnUDu+vr39kfeyna9hoq86LaSBOuS7xhR+Jhlvq1tjRCjlgGlWjtO5yWt5c6RXl0RH33DuAWl
aPRZIHMFbOtq+pKKoN1PdE5PMx7Zvflo9lyk3MQDBi7jEmM1ELNRTR/07fWaA/HD9l9wcqR+ObhE
LM7qNDY7KGZQjwxfh7LEvEJaVif4QxGqT0yl1CjPNYGJSJkx8B6QrjVCOgJHxSCDyIntFAkCtMoN
f3gUpohJ4cZDIv+SV4cqXMKqwJ6U25NMpGvk0pjk8H8b23edjRWLZ57rskuETdTKDhEsJaxpGy5m
yx7veMB0x1fVHTuOaalWUYbYNlQSW4owM2zBHn2BuSuw2q3tvj13FPbM8eEam6X6oWsMPhmKyzV/
eTfyq4OO8D3tXOGvJZzEV5mcz/y/rrLFf5YmFe0VCO54h1mCjA/n+vxLItO1p0+Wb3suX0FRj84A
2dApsQlxaxab+K/8UY3H7JpBXsxChMARe8F0A/H6Iy5Yxv1bzRBT6vqDDxBqAwowC9YVoZXBRpS/
1h0YToK+NbdqZipMgouuxz5R7YatcN2pXijO4TAFYoAeyRF4/d3EZpK1gFzrdUN4k/PT0YBWHGCq
+u79/CqI7QMklhlZlooBY3kpF+TSKL0K6SHuTxxNnFmJYUiep3M607g+qlpDVUzhf08QWhwEYQsj
nEBrJb1jWne7tlW8AvVYAzeTNkbKEyuSppo73dRxl4E0O2V2MvqsQ8FadgoA0+ttSIIq1a7/TKL8
aN3eooNlVY9w1MPJv6tHyUciQjiWSjWqh/EE9wrJ0asFmqs4AhvrUoSF8nw0bvyXWNp3m3tqyHvI
wHH2A+hK2MjtPKSclCNx4wR4XlGgaFz2H3GiC9vPN21in3ROkMo03o4VGpM8F5XW7NynEzBSORhW
jJKs82rLAJDTw53Af7FwXIzhdZfXW+thGvFNaqmXX47hptbZWWm2jRdTS1/oi8Unp8DYPH4z4zwJ
RxutHHdizyn6b0A76K/UB8bhDnU/+kzLvuaQ15c9uGda5HFQ97pPDbJWjoRFQ5+FmkvY60Utt5GX
/FgUEZHx2urRkKbTgKSPU7BI+1Nkpui38WmNBrWQ8B9hoYURui4EyVgzZdWl2FxW93Gz5EkbcGgj
5v6scJBes8cr08f7ybIiHfCW0e8WtrMHz9ylH6b4v5QZu7GkO9riqNt/Xvtl9LUiFtWlKfDnKmMQ
JZym/n++xENVpclbEsGAEl14HBWPNxKmV71r9nsj5ilNGCuLe8iAvxa88RMFRLruTJ7IZtgYHr80
/IPzNA1RcOHITgp/DJCrBNUejwUviz7TLoNvpQ2blNFJ96gDSlkwQypvRKICoyOQ/UFcSXEdEpxf
54nK4Hy3nEz8vVcZayLDclPPRIV5fHucuGn+c8VCbHNCjM5rY/c0Wp3oeZRe2c/A/nr3P+/hqM06
SSI5A9vyvC85s3fVtcap3CNhfGJGRfNE8uebuHvVAyyIuUWM4NHFA+/kT+3cbI6RT0KNGtd6kzvY
PVGCp6s5bf0fGB35FX6wwaN0ei4J4z0v3axcUuavoMx458ixIDmaR7wve1z5NAWhlr6yYOJfZKQo
H3zuwgJ33o02z6+J0SV+QuVtEU9+Qw2vscydJRqGhJkUkVfA5yM9TFtd4IjShPLZa4HSnioNgIUM
aXICENcOYsdx77/TRPpsdu+No/2VeYONWAZXEQf4HoZ9em15iuhyD4ZeE56Gp1aBk6kFr9X3a+eg
1qDUtlouc2sNwH2NF0EO5E8544d8q+8K8niW+GtQqRAsAo6MmuuEsrGhi05LtKnnJIZz4ii948Wx
fvVvYjFEbPTAf+QmqgQ8s4TlryFsAx04tSj2PtF7v02vUB/Lnz7MfBm8sg+sGlF2wEIPBwljszHo
3UMtBg2t2pISMOTiOgwA+phwiKRsuT7rRsAWtn/Eg9ENK5/VInnIGWF9rCOChN0iJIQ8/wKYtGaj
z+Er4yvY2fa+VQnC0GinAKDEQSdLzft0C14/Z3oGLhGtwvnPNbdXSwVhE2JdV2fVRY7uvpn6LsjD
AlJpVoesn5zgFWFtxNbcRXIO3JiBS1Rz2UjIixu3TtEDvXj/8QekpJjkL4CcUc9AXHcn9YGrIN4O
G6bzVMUjfSQ1W4YWVEuzpR2uEauJNppffE6FxEMzHFi3CakoGtJYFcBf94xSys7loX5iW1Ql+RUf
1ChX3uuDcSBTjxEDLanbzeNsd1FPOfCG02eVU/hEvvOYCG1+LeGTKsA997CTqZb6mvGllRJMkPBK
4mdXezmh2UGh5fmwkT2bcl5UR2XCVdTI+aTPxDDHxvVZqyGiiYqcB4DIF9SWnvaMnhsb8ZLH3oMs
cfPWOY23hYbW+JCXy4mUJhNGnYAHDa+X1rVAMUbKJy0D6bxTVCAiHPuqeAN+BSrWv4oPvzvvmQyt
N7iauuutq/fuGYtAdCIaUxgiI68i/RoqTtWTVmbSTygvXenucT0eFasTlUkYtYgII4rLgPDDbqwJ
Q0vtoWTt8fFh5PO8rzoIcwxfJ6EJpE0U8zL34SFvcXyocR2/Nb32y4hL0kbMBd+DxLd23Y0ApiY3
cPKTQ2cvVVH2nzg/FuXPtnU1DuBO1EXF/shHy53Mic15CJ9t6tn+qVUP4jUIdDbtpUpEvIAD7cNt
jVC5zNFMDyaGc2Oa4rTJ9VkUfj4o8eaMcgRRod2RYWF+aHigiaIDR71J+RwO7gGO5Z3QOKyonSBe
XPzTnSKuLgM5Eq9kMw9Cv3a06O5iKBxMeRrZCdgzHXNdfWZh/VpHnuaTBxF507n9HyAQmtuQ/As3
tFJ84MEkd+h+kpEw3Nl8NLVJXCivHQt8/yClzs7fDPLe5kLskgb1TcCq95f+NxsGfn59CgM8Evjk
hfOqhHfTAybmYb2m8PbFuSnTI7GKnSeTyS4PfpsQNNM/NLui+YSZILXeEi0vFqDQ9DG/eV2yQZ9V
7M7xPfspMDXecaubn8QkV40QTzZAaHec9cCT4Qw4J0kh+RNIw9P8gGlGWcjwQHVzJasPtJ2E1kK9
DI+zkbGboStnZfWXHknIucToPtMIMNdXBmwReeL/eBGyZ8/qvLGXXcoUX8ILBuav+TZD+FxuFOeV
h/vVVTwz8Du8Lua5FzjSMZDXjYqsy+5eaCyo5JKx+/dUoC9H7BUWJuUXSJGNFXVbHn9HWvIj24pB
kx84q6XeoTJNgdWCgMUrIOHdYxPFsp2jMGVoNqXdEMHc32fJ18Bof3ji8w3nbLwAEhFoRngID1Sz
q1saq5ka1pxBSqSnUOGK62h7h0HnXccXrbPcVTpqAqevFIthwpV/AE20/u/kBUuzieb1vxObOmnE
wLkSso5hXGrD5mlzjYigUSzexLEZRvkaYHWCDs03LAx7EOWYWgMOZ97gy7JCgAwRaiQeTNYjUKpU
HHHCqBQqX65wfOdZi3LB8tENepN6iAt8qLAwmACz+c/mfv6OKsnsLb2MShiRp+LZ+ioAVfZqcaYJ
hXxbjSyGApx52LA74PYm+ybC3NDqQMMzwgHjyZhmJAaN4DubD/Lthl4yOGmSWEQmPxoi4xnfdO2u
FR8IaGrVTU+FxqxMwwMsf4PMLLSb5+ub1k7Lwgw6EmSbaTDq94NKNmq2XWr6D9DMNNFI0LvT/z7N
BvmQ2Yl1MuKRt7o5adubrj3NqFfXX2wN83ZMLfuoXtIot8ZQ5Wx3E35897k+mDrDk7HWQyoN/Fwx
NTPuol4eRVa0VspKtyNPoLcJpmKG1tUxD2vNNz6UPeXvHJiVnKuUC8TMEr2dqfuSUvKKlcvcNpoT
Q9q061Dt8Dwhoc+qCr2STyBdVT04pmGmW277bxsa448APZLDJZgUF8+QtDOYtwh5d3janZm0u2X9
S4HiJwpEZdPpqC1HradFVSllvzXmayMQTvsh18Og9e+kBzKCez5W5XcF4Y3Il75/YhCMW26rB5vu
tuV/yfFOwprHi8w7qdkDGYrCJYWtE3rRvXugwmeN3G4O1kDFpNQ3KUwcFU2jy3/61e/IyAFxje7Y
DCKWKIc+a2uYVh8Z3wy9Fq9tWwdkdyN721a+XmbYVtx5tUiOh+B5FrkQkU0bIaCYYtaI1dw5k1UP
OOy40WXaYSOrC5ZWdsmSRwhQUzm5kVoKBFdOJTTnPScwrBnVil5Yq+vItSZNLMLUZx/Wa31W9Gho
DcorXXxB3IO2wx8AASmm286BnyjU1bC5MXasN39c4rgODTLdzZNh2nUKMR9hCwloPAEjSrLCJEkb
YatymIaYVUzeg0tHhzwBm2YxPhWxqUEg3oxL3MzKrELf2yedN4lnXSP+Fp8hWHVsdI4Fe9K2Ll07
9wm2pFc7xbK0/s/Vwp/QuSPYqmSb0uQsSpWVJfHmBloQ0eGMzjpkJ5PRK+OnozCXP3kvKi4FO7M8
8tATrN1KTaQQB1gYz88uEO2drdRSDNe7lUk2Jed5adO9VKURR5AGQcyGwhAIqnlGSN1CdZBOERxx
VcIprb8mfgCnvRMVEChcE/SsvTfzC8zKUMy6jzvGPQN1yoIS/RhlhlLxhDI5sq5SqXYnDhHRaggo
WJV35VeHdzKEAKlC0bfI0IF1J56udBfc4et4N0JAuEXE2YAnFVC3fmNxCgAUF6g3yOIuw9TyZ8Xy
WO5CKD//33VYE7kO9iR+wBF+gBsnxv70UmuMcul9gMuDkhQk9+2xP5YpNisoTibcFVyscxEYmUWB
5WZCtgrTyHgmW887ZW5M6TEXojS9rUav1Q3lpmOne+1SEl3rwSjN43ba2SoWswB1kqgd4UoZ06HL
5ANScdrvomT8YwbY/5ZnZJsZLIAlkJzygBEUwyZaes8eHS0QjPj3+yGHeIbXQJo5DcssPl7sslay
2zgdhzig1dVBV7rFQWlg11dchh2GLgEaRmlpNLAqsSDAZ4lliM/puXzG0U8dJElhbzSKSS4LGLgt
AtoCdvzEl3XegLBlBi+TNxBzvgfWaQkkJAGMEan60oPgLQrd4eiirtHxHDjUAvk2SpWVlAtCGkx6
K9f1IkBYXlN22kInTzWObECaBBaKavyUQASucMDyeluJU1ulLHR3S+nMkQ04Fxpvlmx4FFZ0YEW0
PyYgXqTDNRzdWmwPUl7eGdhwOqZi9KKYHtIUXafA8ivtnY1wMAIU2r9OL2MPjQqlTFEenq6Aekfx
uIj4WT5f9br16y3TaIGc2FNL09jHrso30r2DQB1/8upfTJ6S0zJHLXwPlqdD7osI9MfFeDvTvwUe
4FuvsUGZq32a4bmOcPwQanhOAk7Yyy8Nr+s3w3XWC97X90gAMXGHFYcBGacOmRWxkvd0xcMk/1LY
BTyinDMGQBFT6bdwzNP0b9Gf3rAViIF0Ndxg2RNKmWkQ7IhZ5RJNeS4lXs8GtmCRVYmaOfduQZom
nelKHERsSaYP8H5qwWqGJhJJNny9dAMKOd4hdigbrNVok261jFkx52yxDdCNpNGbf2rxVUDNzENy
FDezWFMeGo8WFyNkJT/kIW7h8wsEF/c6QZ0TxncthaJGVuwj8e+HR8cXTocikNwR9/VcCxR/Sl5f
HwleTeMd4Z56XLlwcqLK1JjPETpGDo/ELmc59t3xbE5hdLz4Xu/0zaEnt/4RsmopC9u4uOZh+yhW
XepaS2+OCM0mD+HpQ8LEsHAiYDIbtAlWwoV8g12lIZXduavTSda9YFc9cIGsujukx3w/vSv9QBQu
NNBR1FPFRyVaSWC8Nypl5AnecFF4Xc8RUgJs9MF6g9B7R2RGIROF6h88alv7k3X/CImqRUry5vou
FWdYtLkbdwiArHw5QLKl1zjVtb3aUVp7rxhnqWpWNJ2fuf+MJVIIUGx7huyuCYYP4WN5q+J+pmqd
ai3u22v2kIZIgHgO9x52FoPt8RqlA3Be1G/taeFchiaeGgFQXY30JgX2dVcz4nfLJ60ePxFSxbVe
7UPMvviTzzMj+5WAN1WcMWkPw0+/P0gEC2FAdLF5i25m35VSnbGSjIk2d2mmEe1LNyNWV8U3H4jz
slRV6gq5zAvzYJAFc0pqLno0H5q/V+zWA31m7BWObyaXHunI8EKgtwV56agbbwhf+jKqXKWZahw3
WZpsu/cZkeqv0K+ytv5U3yY3t4Ay1yJTKVtIxmAWFB1Dk+sL9b55CIr5TQ0CPgLqM2c9OJEhUai5
tLygW2J63AftDrx+49vIEesqwT9f4w4rYWzrMSZ9Sik1TXSCv2l2wBMkL5/7ADmbaD9LG6YDy313
B7h1hXLjo04MAqWwui4LzVVJLMCZJFtury5QQU3XumNciYXXIMDLQS/fxBm504olKNW3i4zpcpjE
796dZs8i59Ji8sILcN+0YiAd9rCs13g2Eq5hzbr5qAFeWasVZ1HEmWZtYMoZqbE0clDYSPop/uvN
4QljsBWSavSV/3e/hSCQZguQAjaxIzSY6uc3PSzd1QFYPMWg3QtCWxRS6zCAykssJrS1Jo6bByFc
VTrcQRlXJXw/GEwi44hqH74I5UD5QicnspqBf0lkTGebDdnHftS76IJLejCuj7ryZTqB8SBWrXEj
26dgVtDI/z6qTfqJ61rTeP4P18fTL6xOvjEUiJCBXLArm6NhpyFzZJeA+DQkvr+yj+ntgf7caPPh
U0JjSpRU7p751OocT5YlrziTJkV3iieoshJv4J//F1vgTTf1gYlixdQD7+KxIUTVjU7mwM1U10po
VYVUZiKx1ec7mfiMozlWyHpsATU6b78nWf+jVj82Ppyo3V8NV6vJTa7WeUSErhqfzLorZCs7UCvy
fl8vxyHoLN3/iOMp3zfB8SVavoix0NLS6qTFPIQbjgAIyfMQiZ8XZJFPlXQmJQ4lmwf5gARt/y2d
LeJV8i4KGxMW75uOdGDtZD12ZdHdR3cHkKmkomDdda4tmQmoI4Hyq0Qji5uHKmkIKm/26FxFrZRx
/BBnniIYLy8cYqQqsQS3QBIFLdEomOA9tb9tkulUqMbjqF9O2IxuHJrW0kiro1c2p2paieJ01/Ml
G4pV3rlHxQie27f7d6ONwhL03Xo9HMHLsQVI9/QhXDo69Ah0gjhYKDIv7Z2dpX0DJ4aThSzWDw24
kjUFFoXUQPh8ytiOeBcywuwnSm3igq1Qf6h5WfAyfTLhm5qxq7ce7s3TdM3beQBQUqEH7Oko7z4t
HupVrsG9JOzZGctwx70xFXrBpJXUT6hy3BxG32GU3SE6+wK1Elv/6k98LPUqduE5Xg/7dB/5zCC6
f/NIXtHw1wCQ3sGQOIXnrhMjSO3UvNuNfzxs0G2lCK9Mmm4gpj/xuXoIGjKE+Rbf8BaifhyIRz17
6cyMFgkueJNjFqj5yb8MEsTCC9WPQV+TeM9dx8i9R3wO4Lb8niGMK9xgv9oKlBX7vkroIjWKaxmb
XGqpM9ynE4eGxh1CZ77RbqwiLNuZNUcgy1mqRe4jwuFZ+lux5TT2+pLiF0TX9pyDxSJIkt1MtDb3
TfvMYK7a57qm6L2oQ5T2bKnRg+MLzuo/NqYVmp/b/7/jJND7R7PgOjwiqAsMpYIUrDAE+9+pNNz9
WAKzWUk52RpkzbsTo+umoAGOTsBwjp6MstRRr+GnUMSWZEzpHzu0O6hEeY7GbW3eIZgqhjYVL9eT
uAJ6vVODxIb0Iim1CfVflsGK68zeGsScO+0nxw5ju+ancfLqB9PstZNYIHYyGqvr+BxKwCD2fu0y
pTuyE4dO6IY83wLfbl56XrJY7lvUpPl3xNMYCMNwn6U0DEkaz5yQWm2E68CNZ56Q1vvLmKTZEn2a
h/nxNtC8KXLr0x0UZ/QBIj0Mv+BkmM0oH5cnJ4qXeJA/XqCpd8RHgoZ+chfufm5UdJKXUWP++9wT
jK0i5YRNwScD2EojUEvbiQLace5hQ1g+SdcZCmA8W7UcY67+Z8qavRzTYQpo9MjnByMIbFQwcmpv
ATBmfOSQ0ZMMz9lzbHgsqTfDIHwPsYWe1bqrxfkFWH0ro7olnUMJE0i+LYrjPklWfUFdnJHeti2Z
8BPr/pyeHGsCuZDtSpHHMhFoc7sdbEGvJOLU39pcz9Jv/SnaWs+ls6vEdx7KHAdF9tKDnd3yevZa
21IjBcAPeURyKdiaccj//Vmxvo5jZ9LqCaeE4nOdfekfqyV1ciqthA5h+43LK8A3VwHruxLg828A
tKl3Dcwb6oK9X9g5mQsY7Ng6xFb3aiQVjeAIYVvSisGVBEwRpE51erEuKJ/x/A/pax49vzl8cOjK
DDYgcqftQ4e7hjiEmJXK45Mw6h3o74S3ThAeUhAnwTcHSw/C57W+KdKRlnIT98Rja/yeXuTW1eAz
b6OWBT7JcPGPa6VmvA63V2ol3ceuPaTHO4relQbtw0poTCSbsv6hl8QbqGuDGdi0f7kgg/Rjjk/9
csgnLTiwPW592Kun4hzysF0/zACehVg5PgAQ9kka1cS6HK14oWTzUyjrGL5ZtnmoZpZwZk2sLjt/
Dcm9odFp95kQEzy/eTKkoFpf5BghGJbFEwyZYYtChQYWp020FCkjwHPseC7FQFQlY5s31AdfExF/
7jNboSE6MzOjxTH01gY7yHyp/p2hIqQZ6I3TF4+HmWwOLGrBJMYTjRVDDVpALfLgbMDGZX23dbqs
SyV56Q4h6KQCCPfggmliCeZNAF7+Ba28tfUrHthgVQCkSU4+8Ar60dZbwGBBTn1zLOgek+Oezep2
PblIGJpqKjQGlFjsP/xfy6w7HjaFR1TjRYRpBRAdHoS9XgmuHLD39KRJZcBXmMrFB4tNREjmUl+x
MU65Oe3iso4NEGzvSQwmK/8J2QFiSXxRBps+kxlEz8EgeaniBCFSHIIJTdNlx8zpHzgfS4yJUIxs
lSWReblGldRVhQPtiaR5QjUgDSqowqsAQmzNrfR9yTZkGfXlYnbbsq5YI209EKrYazayCwtHHGl5
D6WnJfN/h/MpDd9pr7fPyFPJtLBOFbpDF/EAfOz7HtgBLyZS3tTwzOrFpxt87XQVqaFIHL0sRCC4
Lu7dvwRjNzlk2nJ3dWesf9P+/CASa6QjPYGrcLR8vJcjPg/jAwlQuAEnwT5i6ZJOtr+7LO2rnhKX
hiUc4IWYqhfWyqGHXv58vJyDUSl1qieWC4cp4ShtjMxLo+q6o2f4lyePk4r1XBb21R+jVpEBWYH2
SqscvOaHif6m3muaLnF7EYmqjAtKmI16c1H6KmPsN9WZlBNV2ppF9Thz4hDy+ANkTNYoXQIQiiny
ldIbM3Y6090c0okvt8dAXwdkGCeTibMxsfQ2A0TlLoGsowvsABqt6nwK1AYD4Zvpn+6gtJxkFO1y
zPNvglJ/NjtUj1OX2uPtWxlBhmWx90/NSUGm2QIgnireNl/LmghcKhKvctMnB9KQ2r5RmvH4yU6K
NsvLepZstLHkuzh0mu+w1Afsj/PikVBGe4etusW6YKzmS8TuY/qfjS+5PRQczSrAlB2Gyx++mmTM
sgPcIGQgzIQUsgqtluV8my2+kVLZMsrUou2ECY9c/rCKD29sGoGuhZbbp5DiD+LXom+z+z5FYyby
4ct2Hbv1U/lEoT6eKjTEyOkp13t2Acaji7yyrTTgBIPw08S8dXvUnAg/cgYc64iMXRBrNM14+akU
JrUkQRQWbLsSR90VjmtqmC3DD7rLbEUZH/cL9ffUjdY8YTEf7vBRYIXbjcEQ7c1cuU6sOiUGZmHU
aX5XY/mlJ98Bixrqqqaj2jSsJ4qClLx7Jr4F4QTmMH/ML3Ms7HTU0MWn2PV9BzXvR+i53uW1o1P7
y8RsV5lrpkyHtPwnRofFLDezWjyyWt+UZ4VzZt6kkRk21P48lBeqeXuAHrPVTWf/j0pB/d1BcK/9
21yTUzLe6arV4WXjyUrptVbWEeIKXGQejXvFAvNaJVqkXs7QWJPkgKCFHk/G/yDnCMpfExMoHvY1
ybPZz774JgnTkTGLEns8CKPDVmduapfhGFbgCKQhplkWje8ldaKsmd9rhkhGaWoPU6GPwX5w+STw
pBjMhKFUBaFBVVxPPV8XMQrfKPZ+X7qZarPxcd6O6//ItpstBmOlerp+9sRUWCmV255tOiIUx41P
uQNykh149s4PwocPaOAu+ly4tUZM86h1EKar9MhRhRDTUhEqMbYQwOadEpt+1B8LBC5ob/CyxxRD
5GQfwsojoXU0YugJPYyV/40NiVByI8yqx9pCqlXLe5FkS6FN26YGZjo8io/ezpDY+GIulQklMKDM
w4lVT/SecXxvi4l2ToLeJ/XWKKJp9TZYo6KDRIMmYDTz23pjfOHGT4Gy8LlvUcyxLFHdCz/Ps6yq
bGb+Vt00ZaDVVusnAgrAoPSik2JIIQpQfvRGr9nINDj4j26ZbT3GW0orpYSluh73gifUSubPuCsa
yKOy6DdFjQkHU20ymT6A02rBVd4Vn7nniWMxC3WjV6sQ4uB7G3r/bVh2MXb/G3eO9JQYKKhkj4YP
NsKsTminW/VUZEFyHgrmqBVnRtkRItzhWocKubr7ZY6QwrHgtiTx8TH1ed0v1zcZHysxI5bMNL9n
P84merFYZYD/FN153AABWnwy1oBPxI3L9f1ViJtPFWwxxfVsZSlNo/ClDvISDldGluTWT55ElZWk
rWzFz1Dg+Hyvv2S+9B4YBZzPJMe/kVH32th26t233ThbA5KpIcqWBlmBzxtKSMtXzjVYxxLe8OBG
mL04coDTuSXndq06XGYjp5Om+/RqRcExL+r4Cysg6mVXq9ItPkT1WSkbTuypNzI3sXEe6/pauqgT
nO+SKMMmrAY9XJgmdeuqgT5rUjqovmpLerd8MMWEoUkCt1HhzeQ4x9P9GjliCZz5Kc5o1S2myTAB
/McXhdchLJsQMl0/MtX4vMl4sIDhy3/GAlzxQVT4goC7qENlVHaugWkB5ZMVqm7NsGhl/r70MsE7
A//lfCCg1Z3d6xz9hWlnyI4uA/PkZ+1D2UYBOkZsv3UJ5f8LXL2f8diFU9EUwEcr9FKhpiFw5c8n
gQkng6SlYbELZ3XE23fl0w+ju9g7i6r96idTSG3X/5o2wXmTzfq95ZUKuZGLvYif05Lc1C4tyDnR
994KTk6NEE+9/aP1yVhxxi+wF2jmHjLc6HWxEG1IwP3uaplU0K7u4QUxdyNHG9cl0nSStxq52cDJ
CIMl/OVlSD2zgi1HRMBZuiDNm4bqPncNJdUSfOAbbrnf9T8GfNLcRyEVTQEIyns2x5qM2YD6l3PK
3X4wvDrVoo+gCM8JBVvRR4ztu+So38ILCPg4ddory2kDGpSRWU5tKQls5NSSrMnuLFF74ijDdMaH
MyCS14msGJhk5kFdxNe9Tg64hIICIZRghuzXfz6pCoLD05udmg4hUAjh5KEQ9WtHsuHgPkSKyUW9
Pu60uMYwHC0tN/7/9jEklOAXHZQ6wmZWWYA1W5U/ejnKOw7LCEKltHQ4CC/7VlPjoV7bRNLzYVRA
Hj4vKPy1ubiUuINtcrTxCHuoaMLEBIZsphYvqkZ0np1YeeANa8QKQnhZa3L9JJ3QmIwuZLsylzfQ
OmoPQjV9lpuiQYRDqjiIhAOdWPAz5oB+AjzJHddK/vmL/sljkl2Tg2FF2GW1hApNoenFguD7Ovzt
XCgDn/rQYSRqrXHSLiRdbIr4WKu4S12ZLbIusxiLqqwJ0T6tsylVY3BxPyT54/zm8Fbkc/2hKUAD
L3eaGhQyfOELVyI4i1k03qio4x/cGbf3wMUwrI1CFoeaBJZuYvRou2sYeatO9CTtGZFiKsDuhn7I
uHmFVEyCtDHrVI1/3+fcdP8Rb0Rj3KxldNtey6lCHqoRVDDI7YThO5OGhJXitQxynBHvya/P8Pqv
wbVYTAPZghy+7cFsEppx/SJwX0reMnEA7P8EtZ5dXfDyIdkQ7Rp/rP6RP4FYCXZ6hCX112KjHAVV
cWILpyyzQE69I5m/VrdTpUemiBN4t/MXdDVs3SE3wlt/8AaGI1vZoie5Yh4CFWd5KfkevpDFUZh0
iyEhsXXIF03EEEFv7cZc2MVldPl2dJOkE796UNBWMaHng+iXSAmAuaqVL+Lufwipm47gj68xBDZs
KWAMPlre1ENOz86WJD8njT0LXRl+e4n3+R+Ao7L34qTJBJRc/Awh14H+PdP7H7jjwIssTT38kZ2f
AKeDDQkN+P8UiVirpmjVyjHIpGw6j2qpAtLWHmthfYOOo7CfJPSruvzKv8UiVATyg+udQHv7KcJF
UNEfho3xXHvL/iwcsx9N47LSDYmOw0zrpmNY1j/OKtL8zp1IVVITACSHo8BYeVFUOHN4JwncdHSp
D2sQTJ5oB+fEo6WsY6NHVR8tfFFGP/jpUChKjQUD2LQn0KxHatbQZQ6TLms6HpeUVtXhrzW6ZNrX
UQ1kgx4oUIGHUL9eV06dvLbjO5JkxOmjsEm/n8e5zaiZqh23wbHKPoaGZB2i+Fc1PgYQD6BCiYLP
4sAdeUn8/rpCaY2atijSZqi3loC2A8Joz0kl7wH/klmEEgcbznX3PIKKeZaRD4ICTr+N7J9lwqtY
SJgyYYCkR4M9vvkEwLXeDEPDj/oDX8bDlgPUZG3m2jDnLDatnothRQyrooXFwS9fxnP1o2zm2z9r
hnpFw4xmjygw0dXaMjxphh8Iy6+uRsaA9KMziRzCnVKFHgu75/WWv57KWnTkIcstvFatZmbinbWv
kOq/b0UIoQ4lzUZTHhXpfH79+zisltMPADtnWDlBIyWfXdChwXwNk2T3yr2jpZ2cK9Xffq3YUAS9
2fxAFYqYUgyammj5dHu7D4heVRj+Djes1YxtRb703hqIwRxugxMQLo2G+LDZuy4wbl75uBX6O7EC
51lTkTKZq/A193o9cqLEpqUsaHEAWlxQZsmOLAmZ0uqVwykxM/56LdE6JtA2CTRsoxKhSCxmF+jX
h433F730K0m3CtyGjmoorM5IXXNL6G0cAgvVg0MgE7aTHiWC8Rfo18W4af+fpffuoFckPlNdymca
nccuA2ja2ZP1cYXcjyh2QM/SlASsSp3BtlInk7xwHVNYRwQLC6ytEdvcAf1HrrtDbJ28ta/L67aH
w4A43EZMfRh6DjtmBaJYP2uqVjZN7IlLPoUtM8BnAXoqBPy35aqkHdi+p1GPqmwbWAdB4AAzvkgj
YTSLSGFdPIanGz86ylV2HqaBVxfROAxvdtzV3JBfEOiThrmapQLcjOux9KCZQQjqE2W/uRO4Gcc/
KolIemFhe5x9vqa6Ru+Tgi8S+fFJPlGCabHx82rGA9eR9gpa7eyzYE4txrOM8WQZr+ICZi37VuOa
K1VymVzFnKggYMu00GE0+6MTZ7wM0nckxkm0sakLSzvEw0k2KR2x7x4Dfd7r20WOhnynSfhCmT6j
zlNy8HOf3DppurM/wSKYjeCsFjdfxqAOScGJ3QTcAeqOKsy8OPEvfXYco+jti2w/fKKqysN4Nin7
OBvA7r+LePRhtGFBMJPc7O9ap5E9/m84NU+gKq6ZB0lRWyO2qm2vY8J4TRt2imehMiOXVW1o52w/
gusXbW+LxySQOyt9tbltTi2HBkbWfBhNUvomXzvB4cYUjl4VRhiuhRjGe74wTJwTGN2e49F/CkST
gL25gz908jzne0VQABH7Mj696c61Qr6HmA92ALZKjwiF38aOYcuJ/135RhS4hNDzgnS+GTr7/XDS
sw0v7UPQ1Zg3phUuPwr7UbXqxb9KKxSz/4Vo26JmjN1YW3BAsMI3MmNBycjRT1wO6SmqJCmpWunX
8oTtVd1VIv8bNiviX/8yepBOHmRke7hkHBjFKy6VrCVpGoIDiiMtfKIfpb/aLB+5r+NWXz6DTIbK
hcriJeO+7JTTQ3XvY2vuFGB+FAvpet7vT7pZ3OwWDjhckc3B43eTB8jLgCIHHxqmbcrzao6pO5HN
Vffworjj+L71maHmjKV5pEGGe5EJRimtOsdFqYYa4P6/wu2wPqQPPoH1C6N5j2sMw7/yck3sErc7
9nii+8oWSLuIs4W5dCd8+TXVIVvzYiibn0dJ7gewqghTy53FMUCRHnNpYg3uuE+NqB9llVGXvLZl
m0y8bSdyIMJHAyuyBzaohWO5g38R9WoMiR8e6GN1aK+LdckM1UMKYhgGVHQVB1CNBIc5p0M2BUsF
unqX9qaxh/Z2atPwHSMqh04dAJp30DQhCdWJNIJrY9TpxRgIChkQ4LfU+ZvQx9lLjyOxMzkYRM1T
K/dCnEbkoEnMtzh15+D/xS6naXhSydZi3HPeAeC5O3ktvV44C/9YjzC1zwbW1iiw7YIhREpkEm9B
7EPXx/qm3tmDxHSzMeQStH3KwYLGbiptvaqjgoPvABGDeLktga7V49RSXDoS+JFWuk3gkyWSSuDK
p/kkmFy/xAkMgrmM85++OiBKzW//+ad7zJAPaNQy1P8JpCM6JWL2Q74Skf5nlbnxiTQAdKI2s2wz
jRHcaXbCJ/2KIkSCSuMULdBggg9dT2aSP9brGuktePpcDAEOH3N4E2tcjdq1jt2uZFUR0c05uc8p
G/ySJxqgtF911S3oiqW0U4Wr3aA/TCXzlzilE2bB25GEl8GWzA4TKpY5pB9jjP8DtZnE+kByyc66
t0ag1T24XJGNaY06iQIjYjAtQdiafZ3EMQoQiEuKWIB3YqwiNSsdausypO4LaQl7Pfp6P/UJZNt/
H2Kj7soxODzI2MbRLA4NIkDWoUm1El7UBXxKkCYXPDlnafCI8DHUzQk4+oj/fULOPIGYKSV8uTel
LpxrP+M6uPWAER+aj3AcpJT7jrz671Re0i5IpaDejV3RCed2mC2BC1X8AsoV+ZInCizjOsfoBK31
/vO1y5+1BzlfG4X6TP5rbKtd3hDP+V+/E6esNilKwkuv/WlnlypGDY7M6jD24r0DrvyLK3cNPGtF
1NvfBoSOnTTerhHIhibOVKYLbBhIzsVjk2GoaYIRccn/dCHfdila1ZcK3fQaUg54E4mChZktZEfO
oZ/x3PmHlecwHpbbEK6iKRtfevCsjWotQkryxhgbuzDkRG6SWzTAH7O2U7DyNoF+VDZn6nMYSf6G
GiEqxbtwhfh8IK36xqyCDfjMIr5ezyrN2HZS6BRyJqSKIjZvdrwnK2wm2YMlqU9P1c6tQeqv8mr9
DrsWXdvh3TwfKwoGRFnqbxfyr8zpFhNonyEPMVzSituFVldk6YIrw3xvwK+BF58c8pm1l/pmhTR4
osf57wZ0z6ZngMQlvS2c0P8Lde+5xwqZ3S9dluOoMhuj0wns6INJ0ZDmniCUfBsX0ZjyK7qugKdG
/Q3gBwd+dEYJEGl3NkAHDzGUpIYi2S1KGINB3TOrOLsufDfRJOHCSoxThNX6/E1IWfyOOHmNSuE7
QgesFcDoox7rvAyrrK3glVIl8YE04R3BSkfyHaKDecU8XH7EDjHGvAR+hY2/n/sxn4kvnikYU6Q2
eZC2u8FwYR8A2G8wMrF8SYtv01S44Md+NrmQLNu+t48n+3DtzPe4vklJenfA7jh1Ovx5eHroW++0
5wRvYrXgeR2H/6mpa+g0caw1j6UPidK3SoerFVFYbN1fEz4nNJkAOw0qWZhU5i5gmZQB6YQWGSkN
BWNt0kXzid+BZr7Lz5qLp5DFDuy+dLOQmRLWZwqInO2TGsxkBYeRZHDr+09l3Bh0C+NXSCiJ5hbD
EILU9J0DOFeOgKSUuU6p6FEjZ3N4NcdBdOnefB9Gn5rkGsDU7aeIF13nmg0lQy+Wt3Vx0c4/pF4a
Q1KsiFxbbgTaQMuOwYEnuI0EIkwWS2APttIT/uEnvfoxE4LlzkbzY7zWJgeRMpfW4VwEfvTtsqed
sx5WCEaCZnLUth1dgcbkWGzFI6tAaVrxNOQ24iru0ZJ9AU4p45FxOS36DRlVpaswj/783LgiPgdD
nBsU7iQu7PM36jp7x7H6CS7Qr+t3ZDsd31Qc6+QH/lZ0cblQyejOK2m1lt/zjfw7Zn3tRwP3dwtV
qtW7lvShdXuhDKTaG8WTgn1WspfcTWDeBAzgM9eKC/G8z2q1npFzezHicxSpDHjEgw7hkr4PY3ue
oOQdGfEWRi7RmRTiErAtEr4TVcuBGcoExwEyAnmaAGN5u9HcQFq1e71tVq8p5T5btVnfs6aNUQ0E
wKaCGlwvEFIUm5ZjCDluYXoGfITyRUbBBkmWk9ulQunt1y8NDeAmQkX81aGg5+Cq0wuaLXMihxXB
W3hy6FjlTCpUpp0GdjEyvYTAAwpu4b3zSvk9p3PTYqfB4js6KZiqPmiqo+9cw1bvIVVxOUFhAqbI
yjAQtoqNXJ6Sp4fG0FPwdHCXWDM+mUp7QArwqgvEhlX0Qx3RLOYt0x938oFdpDpZuKjlQBmxQczD
VxmMjEtg3Zx1Ky9qtaJbvvBkTBewAKjgKAG3DDxCYgOZ1Z5v7ZmTsEwk2FhVRYpDD7olOigy9DOR
MOx+oOl/ehxueOUxXlz3CmJ7dNtjqqfXXiCJnwYwXmpqQz4lsoS9lFKMn2e4sCnTMi5ytHv2Njv2
ntZcKtcNL8qpZKiF5+KanbZwJKhQDKO1vxqTvqB1TosJKJqtuUzIhsnwqBStmP4JmjtzVhQTzEhl
u9DxKoK5lJm3o5NDMs6doZ/vIBCy9bxvMFwVWjKzJrZpl1NZuZlwKtwR67A9N06Z0KOB7QlyzsPn
QPwICg5kI3KPdYwMUipQCLYgP7E7DT60Xa5GLghTWyNkaUUAZLwRKQRP9Vfyw5CpgwrTdV+8Tkkt
jaJo0vZleiH5iAcnwQFOQlxgQTjD7MkW26C9X4kCGrkYXeEhxlWecV9Q0LtF0oClTFqluzOorfrF
Q19vLoX+A/iweIcQdCRDbCiYNtOtAQqgktnvzdkEk3b8OqBh8SHiAfXh3laYZKws12skp9ihfHeD
LmzYzb3rydy/vAyZtb2JJlPIv/Ns/PrtpNGgvOxdtw5ug9p6LCBWVz/3+3jM9oyfs4ema4lrk+A4
Q0FFBW+FZNYk6A267TwwfPMajVwuW1lVgCCrwItjvX4YAp/5sJCP/W8Fg68zWfORQFdFTMIrC8RX
fgvXemB8jf26+dxIKlWSb+EcKvyZx5FL8noaoK9LsgWL/wyb2nEY3jdrki0udfJBIpSuwip1Tlyq
faNWg23zoHfHk/T3MX6e3P0ySSW+Cat01OPIRhBzyUMf0HmudcdXpgL0+MRZ5v8spBNxIDhgBzLF
qpwOXjsdAdsblkqFMoYfX7N9P3eVbt1cVnnK6IILnqK+2+SnkqMPQEckh977XU4ffHT4iRvTvw3X
xrxR/1eQBQfvy2IDs6RXrHyN3E0LLg88mIWKbsaaz94va3Ta9uCL2Br7xG/ReckFGKcgyjuO2q8w
lhJCektngKTyWA7NFw4rtV+eQcZA88EHotIjIYACUAQVJ4Mn+vGMCJC2yP/XaM1ndDNb67ood+Pc
+OQ0EyxHbZaIrxom7Iax4qKvYeFJHTNmjL6ZFYbJ1XYK+c2lbiTQ8DFUTqyUPCGf9oGLfKWAgQaB
iscz3s3tFQd4NUg0Wco8k5SY+JbexbS1x91xEYMOuzbUMSIL41P6XyQuMMEmUH8gv/R7EM/WT76V
zMZEKpjsUntuMdZc87C/WJdvxx4sCYBpo5mw1rIoxubrLMSaj7i/dmKn0nIsJ4Xx8oKT6jH0Jn71
EOxOvEZtxmezwMRPI0TR81+y4/VhCS2goiU6+FRBjbq3xMSZVWrKOeaEKMlbGTyQMdtycIHN7tUr
fR9KptpustWgn8R97iUOhJlXwDNyD2wJ3N3+Pu9ju7g6CT1KJvImxas2PDQwQVvYnmsRZ7dr8hTM
a8dCrO594PsOWrCf+VtmsFh8thK3mtM8/vknwSqjJpbYeQ56FL59lZyuL2VBzAqmRdUdMS0o5z29
q2lDw8KwFcjHqYuZ03DAeGw1li0f3IX25mmTsEkMO0Fmiw+j+O271mLKyAHZGOU4Cutdi+NMnNaa
Yc9lbxeooRqWF/mv0MAAm3GcGh7+Z5IUyU0Yw/ZE9ArB/Aq9lBBBNcVQyU5hW6Z7eH2+rAc6F74j
81N9cCP3CAmCzPHsYSeDD2jXxJ35Nowea/ClYslx7VyD1oqRLvvejTrZG5t0AVG3A8RdjBQv072u
OFciD6VV/wypEkBg/jk3EkKNyiWDXbW98XuPVUMvjI7sbhLZB56fFlU7ScjzwTSDo6mcR+VPjVSz
Kkj7lV8v/g9pVeYj8rb/CDVQ9t8fY8r64+y31zD5EYkgM75EjWMkYUrF85mPnnaFfrWguSWVPh3E
NNXHLTNLOyU7k7kCY3riF80lVcYkaRJXCvfWOFTDm7d1AJp7A0BIYd82f87n3RLjVY4i1MPqWvl7
eVRKdCo8ep5TLFtMOLQCBoIq4x4YwZN0GbPE48rGOz9fZthSMZg4pXgEgzMBDUc754Mw3dzIPsGH
7d6hKau0t8XvZo5b/u+7hMNpHgClKP8TfKGNLANZ9D/f71csFE5oGwBGCnYe42Sao6DrX/SMmBy3
zLEbGzaJNSY9xGhuEuQPDggHX2jkBlFvFADLFDU61FZVNT6XpBmqO5VaQ5p7hwWA5KLTeADPCoZv
njJwm0oOtCdW52FruqmsxGCZosrayyzQQcK3sPM7jXm5HJe8WCJVVNstEH6SG0ht7MtufENyN0ly
boPSTtRpk/ihOxw341B+QgvrgnHFa2L+XfHKk9oe9u+aCLa6+eJUT+bxEZ/QLUWDqe4LEbj0Gsaq
f49Lc8wJJWtOiBCgThmivMJWeTmWL9xrgpRyuEtQSvLa8iAYxSWZJrMw64EbDsmPxz4er4LMHVdI
QO0wa2HIOqgIfASF0p4MOHS02EQ9kCadn3whXb+M60BAI72mI2HTADlml72+RPqULOTtUtAahTsU
v+I6Ye0oje2bIyCVAe3HSVStrQLwTUpjOO7dogeNP6V1xCIN/g7QlWpOb1IqBaCLjNxxUjV/S6I+
UpH81XmtBE6RPh5M4KymmfpPlFy5u0CFBFGEQxK8boSN7TjqM8GEjRoP0LWl9Y8DHGiv+nS7LztZ
P9ali3+1yn+80aYRe2DoH5l7rvuOPMGZYTmTV3/E2lsNi9NvWValTObA18tQPgjiQ8Njoa0Ge01B
ASTBN9/42EtThmP+yd8l33qPaIR+fXddamJxA12rRNHPUcFybdtWrKrjw4V9WxeWfqNFcVatgq6n
g39p2ZSTEVNYDK+w86Md5ZfXzs7jWOHB+8zKXp4YgrqLwlVH2QGtJkRdgeU5whbUCrnjPEUTlsnj
1zwIrmtp4MUO7pdyZxyt4QK4nPRU5Rgvb7Cw0n5Ak3Fi7dVwS7+uHOFkcV5MeJnGgfTMij6BujvW
Ak9wJNxmLg06GevnVCivjGyI0/PQBoETmQssapndC7QSVvQfRkhUXfb/AMOUwyZH85OYApwDA5aF
IXvnF2cq+czFpUYo9gPY8OxM38WeKFylMF9i2AR40NPP/d3LmvGcqRQUbUIlTk/CAjxoxzu+QfBO
facHa/kvJjVKjFj9QImV85tLgPNYbFAu0qCqo/S1GZU0B7KAjGFSgi78FysbwTWPMOKemfwLbLBX
mmEeyI74etd9XPx3CcmnjqFVvmypa0RDJe2Vrmn9M160o+y4xLTdpaW5zMXffRYRU25xme+3WiEx
g/edcww2Myo6eEqCeY6NaJNuz9QxySdheawvgSaGllLOYuRccOkO5od5teZte68Kzlga+ceuY8x2
R1J9MDXu8xx1vN/ZW52IqSq8m93rmLqFAgcfitcFH6ulwJNz2JXQax900YML5+trN5PBmboaKKH/
6UBKOFvZjG3n+zbsFBxCVWlkHbkV2LHF3Dqrf2UrawkAaeNct+gnEmBbLPRsyW91FPkLqq7fq110
i6OU1MzzKs3w8QjykS/2nb1vst3Hbl43cn6KTraScqVigh4tomdhsfDmfWBm41pFAqvx7buHSMTx
mL9KjutcCgO6VMQiEXUeKonI8YSattKu+h6y2p/zNd1sGi95q9nq1qQJn+/FOo7sBd8cvIchTkr6
6BzxFVqKdfjW8dTB9UowbsBqA9ytvK5uo1iVYJyVEhjhR85LUMKo9IysWjoNhQIq/j12rwn1hnY1
LM6vcx6NFRhdH5ECn6sDn7wRYqkVF3oVoKlPh3jebbnueUpatiPACONQDH3zHBnqWAjsWiGULO46
t7YGhahEWtLdOBvPf6TkzF9y0DrNIerQvZBMiECzUUDCGO6qZKJc6zrlG/jsm1BtWzS9R0TK+JS9
2RjXUb95xWyggsm9Sg6blYHszqnxPDbIy7gTBUFyjOj0D/klp9H/3QOzb/52oxSxGSpYPkX/I9yV
ldKfqSQeeeKB20mmalOJpVJbspGdF4wY+HVvTWKsglytlFfmGE6Bj0zDe4kZp5xYU0lbFsM2fUvQ
/DmcjwW9YdtifJJ7aEWPSY3MXm4kf8rNJXzQjN7L/jmPE8GJeWuOHz75amuI7SQ2qtZIcAf7LJ2U
S73XFRmbNyOMhb8psfYsJr95+UJ26gmHtdUOsq5W1CU3nYFUTwErfIDh3MFfSWAbJ9QzG1AElnpv
FeEAOkHDUC6t38hjh/Xspxo8tRzGA5JDVdU1zj+Nrz2Qk7Rz5hI6PtfC+FL/3G2iSbFZmKeKK0lm
jeykFg7my/56zP4YBwq/jnltDmUJBWdmPAp2k3t+gAnTLLhbJzmSV+jJqapUDi3TN+jCNKiIUeOM
DXfkLPDb2h7HxOP04Ye6geVef+AWkQG/X4LAtqiMLp8qa6efch3Qp1eLsk0c2UpV1Qh0xVzyhmax
LD/3+ApY/ylK+7O0J2gN9rLDkaBv6eCKHoyStM9by7mEoOfN/ZImVpfM555oQMMw5YRDaxYJOTxI
ezQZk5K2NjJtY43dyaroP825uevMMlL8IstkfUNlVs/BjQ9xlUTYJwAOZPO5dJSARap2pVp5/sQ7
vNKeWP+DZ0wyZ1ryYz34mv5y/eV6sCaU7Ffv/MtszWdrXd6uIppdmblX5IR/s1PKAjB6gfiahRoY
KpWEhfGdF5YSVgi7Wx13qDbcK/dq89wrLZrUAu3KMigrdoXwNakx1LkmZVp+LtklSkykhjW41VFw
8xT5lAdl3RAt1d5VtBFN4fw0FMBFNY++AwfIEbB2s1dWA/5JwLzlMCQ4v2V+JStHhCjuDuRAUW2L
3veei6bHwf7aY8mIlvi65raRPIoYVgdMl55iUZcnPqUg913IG769elbFMJtKFpRVc3+FkG/bnP2b
a5v5CA6BhhPL7zvE2q/3tiyHfh3IcyuRlrfb4nj0uFcHmBPUdkPhgSBwJ5NA9IOFsGkbONVKtH0r
1Mr7VhJvSVSd5X02f+ynHCpBWykRXYVqqwFY3g5y6pazhY8kS0YN3l9+80MHtoWzKSyf746YVlez
0K0YflbivaxSWJ3zkYQjSHlBrbHKwUxZ6Nh2atvB4Ubdp5s8gidYfThKYMutqmWxAsaXryStzd5N
f2zg2tWmI3RsadlglMs+8nQVrF8KfttTgxSJg1nZm36di7Nm5eDV8iYPjQA+VFqStjkoQyE3cvG7
dnWVr+HsuiXjKsqICevdk0TZPwH7IFacSf8VJ4s/DgwguOzaRR+8Pqqx3Q50yP3aqO4I1mRZzFww
+fgSAxdYITcm6nma7pAhwW+DUifX+ceo5oTXmlf+5QjX10cMt5DqurcxLMlcjysMqKskY7T0XHMB
7tc1NxfHb2qumUCm8oTW0TBTcaPiokcdMbypU0igU+hIPk+zBIG4W8dTv1POWv0a7Hsufe7Qt9aD
r+K0C6sz8YRsgg/PcdDpw9+CsSksU665I4WTCLa6vc6GArnhoGJVlnwMQ5ZxsCsu24lqe3/XVxT1
9oSopE9do9G/j3H/C9UVt4SYN09ab/gIgfBRtDv7wouAdBt4kd6aYJbAVm9XPOG/1pkh3kz0BbmW
NmEUZAh25HEh04zZiTKftp4yq6cxcfHKXNCNFXaG7obTb+hb1EWEYU184DokHaoYwPiKAmv2BqBh
jzACBIbItnutb/T79TzvHr2PNe8uGn7hMKVynyf7/xKz/grKApgPfYJfqEvq2NWVMF9+VV3hgIuG
iCh7z8cV/0b59llQDxjg7NE8wXiHd+sKgTK9EprllreoDPnvgYZx6E21nQzovWIF+BneygENaUZH
UZ7/nmGWdSxtBqdpQhLTEYz6XCHqVDAJzVENAUNFMVEbqfcC/HBv01UjpUAzDQQ2IBW5lTqEeGhQ
OwukN204YyO6DQ+lQ7YcZIskNOnfF7HatDRsiRoxLCCvXoBmwL/7A6hnqRTWygwOUVgNMgv2fdbX
uEA9nmkBcwD+Wj4gmZBxFNhfJIQEgVpab9HXFg7Nkoe0VUGjLx28ETEHLs8El5vUluqkDPe76Ku8
43CCYsW+rFckxC6igXk5VhGIXiBQ6KO1qYGQ49FAo5f3sm2En9t0T+33Nku6zfyvllPIiyv61K+R
UAyj64A0RYLNBwOxqjP52341r2Ybb+iCm5IHwP84skHEftT3a9TQiBc7hQVDTKyX2RIan1XctHf7
qaSE+WzLvUcIBs4N3egMD06KwlxqXXxOXTbtmnELcvhbV3veZ1K+NrcV9K3iV6aivDQxOK4HmM1F
h9PZQXMkCphKvAyT4u1m+sJ6tASGMwwiAGJPdQtrsFJwDmZuc6AVrPR86y36Mh2tGrLN2CYliR4m
ODdqq+xa4wFLPkqMcOD67lXpc8UeMN2eBcD6yf6mmLs1AfiOqNxw4SgrniDRGtWpDSQYzJbMZxP9
G+/mIlKcbMjwmInH1anPXixctBOxhqxXhz9EZD4WYQskmKc7njFxr+zsHsK4xOoM7r17umVAgWzq
Q1A4KoqWiKtudseNfgnftxXCvHu1POWNP6FoSbcj4YbdBtAUw1Byh0ZlRgfw9A3uBOvLxfpg824t
+/ffHV2Su23mnnlg/zf8MhZvKLU97TwvNPTFdpEs6w2pv7KY3pPW//1lM+GokLfrAOi5Kt1WTaCq
y0h7bJ8TebgC5yKpf/Ha6z0fYZEJthccQDyNPwr4PaL5zeXHq8sJLrb/SKyQ80xLeRCnoyfkvTFE
/sV3Zg3uI+DnLcoCv5I8hNkVmJMs5S9IHKkTKjhvWaMQ2VH5j+SMgBI0lt0TpTFJPZg2I12L+WmY
aPqT44BFA8pGdl5rnwUWf2Jk5Vsa1cBiX8yBZTddOJGK21tdMM/dkhG+OxtbGvuXqV8bNOQJ2pOi
HE790gPrs8Q8ZQOKopimNXc7DpGf9YjB6dWFFx8gybytaXpnR5fHpOOyNjwjJfJiKmVdZuLNAfmR
jtpjKWANIws0jivCDau4qKkZHW2iz/HpeFnbl2nLBimJbC5w1vnfD/MoUtoGo2VOhdkZnbg+NM8Y
JWRdUaGiX4bi61Df+2CQ/DDfpsRh/041gy9gWH/HDSboySlgATIWqIMh3mnUOH18Eut+u+jj1iVb
xkS357l4eRTWs10fzB6PqQv82omQRTb03/H48OiTvMOtsesTgW8fmZh5zj4aQMCcR3YhhJIx0egp
XA5TK7xwN187u9MYEEQon/UHjI7HFUYm1UMZIxIX3iaQ9BWvfbVPrCRVz85M26Gi50PzLPQGWmE3
dTKFPXhwabjMWzw6tLH0q8o5BiPXTCth4VRconwh4rM/K9DHigg0PYMVIJb+sa4xr0CmvTlWUtq1
avqm1YkZlarLXjuxNDwzW6no8y9K2s9DHSy/zGZHFj1H87bl2URvAZDJQWYsaSdi/3z/rMoNSkZ8
oM5fMy7U5fikG8mlJfUpP0zlRJWS+Z3YcGgcNhMMNW97a/R6b6aOFlEr3jVOlMhiquE4sY1URDgp
K4pZ2B0n8C6/CmCK/dy4ihcmV+B6ihlVTMbfER8hKNsPhPYCocEDNCe85xSNBSBbqRbvMS6EUwY/
zl7Ug/XtdOk+Mo4L+8ZEA+LHUemLOQAVKvGrP7w2Bw2O0QkSOgiMdr8xEtuBCPiJnngaBCFOBOaR
kD4etGyLxC/t+YBdE0thRq8BUq3904AgeLiLTaH92E/4p5gXQJJbqcmycTMDm3BeIo1JcjHJtrS+
0or9e8mnAznP6Sk50jYO/0PvK1SadAfqJ1FvMi/o1zUymsPJIUORRWmddo/Mx0kviSNOpg3UQMlK
iBG4w7SMpcudQpsY2cjvBg9Zg5Y8lbKh4wqVVVqOt8Eto5AeytUNsPLTFbx8B5RA9YircwETQbMj
6CeInMXYiu9pelpKCTkMpsWIwszxTIeFD2xL21Sg+LE4ALQ1Ar6J7OEzKlkHm7acD95BeEgf5AEH
F2TSE/kYp1h7euakucksRvAFjvTDQM8jl5ytPUHKEcaRsUUyarqPdJSfTCU5sFJAooJ+ew5XyOlo
Waubs3PWUivkd+ZYS0JIwOCQ3rn2veqY0Wy2+y40SkWiB8yyuTHe84izgNYNorUtVCCpxntxJHtD
p/2p60J8JDm4LBKNemy2tbBec0yhcoVwmJSsp+uH6xI2d0YwuWF6hOSkEQDABUMeOV//OoQaj3jE
ee33YMfWj0xc/R9UeMA/IzjQpGhnmEQhRxkKZFQ6AhD+of5RS0PrzdPysppgVPohIIQAyVV4Kyey
XPzObU0w2gTmuGQAo0AHwxD8pbHK+3MPJPQJ54tKaYHLUTWoF1DB1/Rlcga2QZNSQb3Tk3QONnEw
Yg3afloxmKrYmfox6LQ6c2Lqi17kNWmXJRoDBYJvfSWrirZmzsMThcv1oOlAXQANNSNpnxne166f
bWxZfOlKOAQcxfja8BlixImfX12Lk3gfbZ6Nk2n3tSR/uRo8FFkXHtoyVvYGdDb8YicoM0ILxHbd
bBN002CndsJX4Wd/yuezTkh0CR56JhmyBG2Y7+QFJdOKoRfWXmFkR2dAppSla0RFclVb4BmrLUjU
WcaMBQ1SbCDCILAnVKDQJWDR3atq3mJhrEVGyLZdktx3n4ppm7n2UcWLfRQjI4cIYJE68SFy4wuO
eWg1QxZbc4CvK1RQ3d0/+9jlk5UPOm0Vk199E7r8LzUvHLl+WQmc/Vy0bfebkqsyQ+XfuRSycbg5
f1PUQKDrEIBtZnRx5GvwiCLBEH3u9r5x5dOPSwNb3OFMhZnaQwMtwaB4bSQ3gcTWuAuv5yQo0BEF
0KzhjB6FeO/2c7DMZ0neSC7IHjgq1v7C/1xQwq02S0ZcoBZwMjmlnASbo2VW8p6G3duq0ke6/9gk
b52Vl0/k6/FLDuV4pJVyvglOjqNkwinKIq6eVkr6SsPXVN4nkW+S40Nj7aya/kUqJ4QeV9Ssxfah
mdoOs5bDSM0JGv9Waa/+bc4w16xGZwgOYqoXB5mbPRWEVtrXQ2aRkLHUTi/OWw6dV9NcbO4jsiuH
U+Fg6/hiQtSySJ0mrgHKrURuCoeZdOFxnuC8tX1wwzYZQw2GPLsM99ENDqNXX0mFet34ZTlbIDTb
VWn0Y9mM7qUXVbtZOFKAqcJuMdf+blRN2EfQJbugscj9ROaHZLXnQyBaMcbSnC2gRAqIHO62cMJA
iUiWeM1nfN/RP7KS5YPALtsIH3tbUyoGguLKA2O0E778amZ6Wwn+pZ3OM+gjSVQQB6NaTZR7hLhX
mDQdDvvQ5cW46vX4fYXzq/ZhOUtaSJ5LNYNIxCVBSTSMP2CEnXpbpnmzwj7KkGq2dqsUWu3xlz+C
8U+urA0s0TadfRN+nfN1dUVrMtgf8GEmEJTUJoTCZm/zxjZ6mvCS+RY+5i4zH9Odz5I+1syzhaWq
ihKH7H56BwBczowIxIPsGv8UiIOUAONV667U4lStim8agICNhLxsTucP5JibKA1znaXiWI/QoIwp
DDR5GGjTQ3T3c/5FwUwfFmUUgMhqfFRRqR4Qd0YsGOK/ZpsEFKik5v6BUz2Vahsb9yUY1y8Sgctk
apUbCsP1fSwK+2f8csqZhOWvDpOxO1MpDCAYaLVPHNvZXl+xJOpYVRGueCb+7AG9PGG3PVEDnDUJ
AORSlcWJOA83pH8g0hOSFRX+rDtf5d+FpDsiEjW24A/ZqBh9gBw1yohcSgwAMch7km8ONM6+Wsuk
sUC3kIX660psYNQuPMsJN2txbq84m2DkWXjWBHUhug+mxzN1E7OiBycg5rvGaptzgzzlQNF7oFlT
J56hx+kDkHPBZ38d+3t/lFCvPpi/SN1cMVkoEnYhsseaPKg0jLh2XSs5Oke8dAFBovjEJ+tBV7zB
FgVal8hgrZ9H76B0p18hf7pYGpYnW/L8HBUIa5fb11Dd2SXJexI+m0/iDffZeslC9KWnBTiofmNi
n5BTfhNU+QUlGuWOGq7x5WL4p5e5IpqnxRuKDslp4zJbThvQ+MSfcgE5GZAjO36ZneVcqbwZReDe
0cQNki/Ld8DVbepkSWdiUCy3nm77Vl4MzAJWn6uyRk8hWdQox4Yt0NemZp0QNXca2Bov2WGGKU6S
YLCM/gyZ1VsCGhKKKNwUV7zWEVv694HPvbb+t+TgEsecDCx3/SwhkKX2ZCsEtzi4l32/YUIF8r3U
/aTz0n6cO4mGrGPhtzjKomEaDcS2v6T18DYetrjYLwHqbpS50GcAblTCjhbUftPvUWiOpG6ZNM5N
vqvlxvcg8L9TKLdKK5VQgAWpXEDiXIQM3g8bPK2RfCHfRxBLIBO2pCKSGNguRKpaeVUbhlHWDjV3
9ZvusmWqIFfk3CWjdtmadEMOlqkIWvKxBPFwNsro/Dd0cSzqX/zfZeQtjRpqxoOYMyqbe4Ie9RMI
HMoErVjXjfeC4pbuxCJahqaW8bw41p7QDtpey4WmiGh39Op5e5lDTMK2tWEH7sS41khPFrWfvd6i
6TIvAFVtDVS8tpNa8AIZq3SLh+y1b7c99nYOQ1w143LKfO4oedcSnEXoVQuUw8cBs3RjBZt27NNU
BW8QiEur8B9+xPvAAXs6ChxO1HhRF+EBVqaZJTbGm/MIWNBFZDM7/qazBE0/ue+KjBykNIfcS47U
144CHOa2jOxNs9m+7oyCVCrjowz3865UDfwvRYBJ6/OvKgVRdvTg30tollp5IwDm6pCeCK40DCT/
lc8C5OZU0MhN4rxFtPqSP0GzLMkORXUg4MdSogsaLWiqUHDIztB+va4WMW6Rm/R0f3v/0JM3X6uf
503S7qYG8BYkJhEL8dRXSfu0wK8gcp5g7amuW7bjljcVYpJEhIjCu5GkksjZXpvXbJTVy2zycl8Q
4uIXnTOHU1Txp9Hk6JOMDDUYCOXyL6i6QY3xkyMW4ds5gzTwShH27ukCCFWoFMPiiLRIGnqbj8/D
elnNzqSjodHrmVLdS9/8aYahIintJM3ZPzEzZAxOjjeUQk8Jex/nWgmOYA6L7TSv2PePXhobcG1A
AbQsY+wx+IrTzA92Qhj1erVcYoUmv+XWMyMCWINZnM56Lv1eHTh29Ct8NE5QCpjkJuJRmTKkfeex
vYS5rN5H4/9y34V2VUW5BJu9TvSzq8u9l8fdnBZXFyN6kEJYim9GquRGopOoywGRUG2RCgF6uclX
jc8WEO18nfNb6eftP4wuiEfF/2FEeAqZo6oZAZdvQQfjCWz8ObOdZKeclZbRJzeY5rB7k4XIvmv6
iirwm52+Uyg9BZfX4vUD9qkGL0fBIqoRw2/YQIoqbsMw/zRIvUG+7SYEKNdhUSDtDz0fQFAnqZFh
19R+Hl7e37CbrchEglyiLK0kqBRZIX3xC9+PtN7LA8mbCGaRlfEj8TWE6PWcW8eaL304rVv0zHsR
XkM6dlSNGXKxfT5sSEvsoUVdQXcKk1mYsVLVqHu2tkV6HvLu6Y2doHyxMXyugG45SoWRFjWk773E
J+Bpl8lVvR9tSaS5KGaacOoEjMQSl93QxraErJbT6DYGUQgJxrSJ+9bClWJkRiRijYVwuRlW5jnF
n7/+X8B4g+cGt4Nybp7RqCsfb1jpBay9fWRD3pqdC0DImvK+BpmqenotZsMqrGLibZ4f9tgtpxcB
URZ54RvDAp/EVaK146wmVSbhK0oTlZmujuYZwreIUN6Snx/IzdYfea25cSuqh8zhteHvtpwn+YvN
NTQfq9EzxoZnqwAk0oE2VkknVJje/O4s8M/EuuBTh1dytuc/Aok2j1yYJ9C53Eueax+VJ9Yp97zw
O/wQlB8hMOeOD1hz0ZrM+fm6eugEq0lyLhQp6dn9aExGCtfUvZ/Mdz0718vHsNpeq1rIXOgK5syd
TK1L76M0Hju/orb4HcjLwNWk295Sv9gE7HtbnoKUiupcpvovKRDW7IXj756hpOAuMkUnKIyD4pT7
kykFA0+5DiSuEL7M5+medYHKfO+J5jLfGUzEugKdp7vVRMGVt0VZYWjV6tdJUKMabQE/hmXJEuhD
XKK9w1T4Q1e62uO8v3O1a4f4Ux4Dw5FZs73WGSk3Tqr0yflSfeJ7AC7it2E0CgulvefqsF7AP0O+
3J9ahk9awmtBFLWD7DMd3wEHTy8nH5aCxTircYR1NB7kv8dUpBLrdQUheXHs5BgKx2mT9tMNjExW
pwF11HQbh5fT+pWFssh/6DH5kE1zTrjBhIgbuxGINpuA4EIz1RS5CjkDFg7s7/6B2A2d4IXR81Fj
xUA/0Jq2SOJOZ3cgoJFj99kOcI+yIEDUqq9TnaZLsYyO5islTFeC5ROgNr+uboWDe2/aVhYSajrV
JaQkJYKyEFOYnuqmFHwgLEQYwz4L/1r9H/ZAA1bhppAmzszFswPi3MiyYl6oK3Bu+7zHN2d68vns
GZPIzzRwVDfHwpFetosqNKFSMcz/EMRDf9R9yvZ0Lfzhs7WN8Mrsuu9EgJpfGB8ohppQ8OcAPRye
ESfKun3D8GJ7zZwkvVHm5L9hnStjSQecG468AeZNCh/zV/kp6m1ABxXIVX4Cai0twknNmjxY3/+M
feDqQcCT7X0FoYeuoNRhUJxIISIQWC1u327eJTudWbs7zG4PCPhtmYr+atjF3JE69VMyp0ODz6dp
cqb/WXKgIOzN5mUFMN97oHXIDTxAYoj0/z5WOYGtsEPdW027RKbD+JsZB0nGapPFjSZCrkznhnYf
AXKzut3Gbo4WhFPMixl3mhn1ie9UmA+UU47JOgBKs9ONG46DlLJQo9ECi5sLbEZrbHB4w/GObyJT
GZTRV7/y7oUfX/uVmEuA4IPHCYDaO2BgRVIzNgOZSUK71521TCM+B9vzJS6X79/D/QCCAsPOxtd9
nq/XIcpmp7Ya15qZOsGz83Wn1JU7fpZeMyehZL4beeqRQ8V2ajaLJxFz6Cy1HYBaVi6AB1lhcExv
AAWzZubVkklOQCqxEbM7QT+uiL9mnxP5Cmb+BScd/U8H5qppDZr14HskHqvL3uno7t/QuR60KB1T
/ZYXE9DfvRn2BsOXJM581CggsUS0I0VL+/mvTfp4CMzPDDqQIbPHgp3HhDkaJNym9oZjo063TK7E
6PvTxb30H/Aur/C3oXknOwtNjzBcWIoF+83jj7H4848jpHFteLYOl46MebYkeHdiORcYlsbutL8n
RsQRymVsvDLqKHo5oQcZwRitq6eigXRRzMvg1ZNppFEbPXyaE/Z5DCjkdZraknes3C6zlpp4VkYs
0w3ak8G5v+iDjpPaEYN7Kw8fG1luEvtWifKgRGOlsSPPUxTs7tSyoQ6RpTE/1SSXXfhoUQ59BcHU
3WYcOFzh2fbo3i5qwcBNJ9suHkgEn0lAhfBITPnZUN8jD+t7041jWE8F206dUq9iVauJE80tCltg
7EmM6RVHewz7ESbLwA0LrSIq7ZkLKrNnvg99cDwHgLDYqvOUVQjjKf0zwJJmy8B+zH5d+mimuzXU
Wo+SB4KL5opewmf1NxxexXtI3gMLYNnI+3aRcZEQdmfHgWiqfLygpJuQ119bWJr5Vxrj4bL22ZHv
Bds1Sh45DTfBPtdODRlPBQy951lTXqfbWtuHUPfgmdnVDnLYyFILrM8K0OROkucfeceT7eZhVQOy
f5vCGlYi7TVg9BEztMuD7sgd1kZWtUxjZluAqahpWaQPAo8O4uSDMpRN61AMUsnPpp7a7nznb4rf
Dn3PpJNWFdX7Atv37NFOfeeSCUzfOtjbKDIdNt6Di5sf/YLgr6njehoL9XGaAv9h/X8m6a1qhXAN
ihZJn5FBwLrPotOP3jFgo+NafKk9hGFghWWJr4JjHkTjAmE72vQb14Yzmk1dPeIqxy9cGjiQLzjg
8qeo4PwVXJ5ErXwNBHAePcL9dhJcGx8jg4JzPXFdmxu0BuDop2Fu7k3sGaeWYh4Gy8PpwQoqoaMm
bVSNIsV0FQT6trK2sDrr51rHiRGddIAbfrnVQY+PiBQifSLumUtKxVJXZDE19So7hbwBCyHB7FV/
aSY4sTv6ptdnN8AHRZNPOFNg6ZuAUYCm8qpAUTAFz6BYB5Dofq5Cok2hbIoHoHJ68V5cM/MwX5AP
F1jdbE+If/QAnSBYnEjwKDrc14t9f6YrjW0/8ikGLe1R3GdkATO3CWhEEAEeDbVFsSzwvv16uEoY
XrExXiOupaubxKh1bh16btQh9PPbMFbsNCujVplIPZca0F/xhEhVTo8lI4ljQCh0W6hMDV5Tl2j7
4RJHkhgcBanH5Xe76klCmlU1inltFwfYTrXvf737BmAqfCs95asaljb/1s5bWuJKI4dyAbmPb/hh
+mTW3Q0DtqqMBXSv8FJqUxqu5GtaWsKd82rPlBpFMw45uQnwYGotSOX5FFMg8lbEFb4NpqKO3xcM
tRxl6grrA1BTNI4B8lXAMSoO83eG6UUjrDn6ukPeFEUhK6LJ5p+c00ri4zexHDebcJPuD/yLu01a
GRTy5DPt7taWn0L8Ox0hFYDiVLYeSWd2Dis29uPs3wkuJAwQMGXccL4A7VvJKwv8QSEc1xLzH5gQ
3fQW1bDP4CxCl8RMnbFj+0pDK1iz3eVCW9MxwKsnFf7ncbHHQaAdjPGWuH/2pwiBmlz6YSmLaW9v
0p4hKkSQnm7Bt805WDlCEUqzIjQBRDxsdvlGxL6jdBBfj5/OTgyz5NMxj4rhzataYP33O3KDtlEl
YVmt7iyvYexNzYuXtni3zm93S/YgFqhFi21xfxyG7hUisiYb4cbYTUOZschrh+YsG6hUk/yUf9T9
nKmM5OMCtdlqMnjEXY1eKd7LHJP29afUMbRRXFWM9kxQ4a4N9HldiY4tz3JWp1rQxL5+4Mr7tbAg
/3qO3cFsU+8tZL101nJLSCwyhprfmF6FhozSr2FQbs9LAveiwBmGWFghgpKf/eMYH3Yj2foHOel3
4EMPxhoScX3WfF+0Sa0VDaIlPQJW697KUJljw52syc2e/buIFULpxdLljQjjzeg9zAQkaMrJ47Lw
MbIWKx2J5jt60Ft1Qzt30OP3Y+YZ2rggd53gYHBZIvil0/E+VB/vh6herCEFBPIxNxeVfdKwsgKT
lB5V4zy/AdhdFsbR+vEyHxpP5pkZLcMWmfgxP3as83EgOcwbR/I9A4RggPUp/JUMTJPdsrkm0rqd
t+o2jpS1yx2YsmUW3y3UHnNvL+/Werv+1PlOP3sbhn/08bpl07pjBSp4g54JPykdmiNW1QqVAZt3
u7iHhdYlIhUooxEKbQxz5nwBVINmEU1NFUxi7uImvGv2yRHmx6kPOdhM9Igb82Kn8wB/c3rIvsiK
vPHENhJYxOlJibCBdgtoyL/4M3b6ZwlSAtNJ1Pln/YcSrhPRxqasYakKb8VkHu3rahKm4kkrLwgH
fnzWQ3nCVbfH9xTlq+DzySvJz/14mGhvd3uO6+DG17walZIV1+RbiPeJGlod8mOzWWSy4ij4Xh0i
aAWPk5eed087Ed+TbnBuQOAV3IEpbLWdY/1LOUyLVMKInfE/407ugikKq2UdiMFC7tSKkzxjeWR+
x+/fwnELVwKDnlmfiMqeqH19rlYPS5TAWSDeQkMAleFGMMavJGFkGQHnVZqEf9QRG8NcSJlh/23S
qlxFKmtBRVIpFh19lkel2ZHt/0Fvz8NCL6NSvH+utKBmfaxqEUS0O5EszMmzBh/zwGULdVhPdDv8
1AeBjK8626Hkx6bW2/l68LAtZXmOSl/2PIvEb9snoEecC5XyMxyqN/Vf9EmVTALbEPWbYLB01yN9
lTWoeUlLT2k88mXNyO16cD4L5SnIyeZM0VLK01Rf1RBB89Q5BHwFKDMJ2R01+FEMK7Q8WwagcbkB
vEzPkTjrjPYXXrYys/mKWTReysjceie+N24s+Vr8sH2IzZyjWD3KNus/O9FYYYqS/duJfiTGPBEl
pGUVUiVCW4wuH+HlMOFpAKpBWkbRs+SjQGY60AdZ19XM93QfZxVfA9OYiClbSbG+25FJJR40KYZO
uMa1qPi3dT6kdeipOGXRn/LgtrBt1pGNHU/GobSlJ9paPRqQ09FcKrpjfJYY3sGVtz3MX/bkJFEV
wJBYe6SrSfh6Gvrq3py9RF/qT2bPUvs9N1jl9J04FJn4WhhFZKQc3Jj65xCbCHdV1vaOu+RB0TVs
QqiKdkQAzIC2nROmjdRGsMnzZG1Qw65YKv++NXcL75RsicA34MWQC7sG6FNTKbcn8hn1UcwGq32k
OKgbqiT2dilGAj0eFiqx3t6kM186DJ2TsWCkjj7jn9DT6x6z8Wo5HnASNmOJLfX8VUK1lrzIJb32
LFJTDGyxwnE9EPYUAKCHpsakZb9TBT+yiPpmHU6DHCHh3amUDxY+TnoIqWQo1DHP4a0gs1UrzpGh
FFAcKHm3uq6rbGoXFEsqSNtG/XIAScB91E05zk71v7/LcrsXuzoLMxuEVKtU1u0ju5GlwsmOYo0e
CjDIkhcJQuV5DUWK6G26978/CsbnQvyoMtOxHw6xLm1+r+NIqsexIUbjQP7HiK1dD3wKO0m3ATlc
/If3qy2VUW+l3YsUxzf+muyY3X9DPq16Ybx2trpiuecVxDRa7v8wFgQXq7aYotDi/6GlwNh0LKTN
kqMV5vrPn5bEra7M+7fZ0lK7pUr658CV1XoQ4jArR5BuunMMlbWnhFM90YN00bEPPM7jsUqsoXts
35MUqJtbzYAadihqJDbNpuELS1sQXAl9NPo4dwAF5TR97WMUOZeYIIL6+5jByd0zHQPkLLpYsLoC
enCnxuLuP/hftDjFiy3lfi8ORxbH0/++35/MTlvJSDFy7WRglVlWcAvLzn24WBHEIoRDvVnP2Exs
8KvqGeOAetqK7EuYuzEcPxcG+P3nPBkkkQFp7BW0gEObaToGxogaK5yV1kEOQaUoQZacEdiQO6yl
XOtmO8UuA4gwL8hWZDFCFQEbx36JBahskhwo5m984m8wPsnljXImehwLvwl3qnhxoi1QnYfNur59
N6RmvHqB81p57aLqbg/V6Pmana0GFoLqJgzw7PNsZ7DV3rCuMSNnK8q3b1T/Z07OA8X5sVFlydnw
bPmMy70fRpcV7vPmheR1vJhFjiwmKEPF05TOYFlZDdJ4HYdyyFl1MmSTUaPKCLDtokMrxD0J5oE0
Rm2HddgEURjIWC9hV0huPXVfRETDppcFw8vag/Bmo++KCwY2qIgUJazhSLO3+00Vsm4a2um5JjSK
SUPLm6P4xw9rICFY02jyEpWb+nFACGM76EM0s0xmuCwNIttFh8ubQWbuF/8rc4a2Csaaumt0T+rd
ki1Esw4iiGNC7ys94UsxZhqxKc2NlQ1UKWT/guvQHGiCiwBJnjZg0PzRPiicySRI3rYjXmWf7hTd
PFrT9MSn2jGvJEFK38yaA6cBu1qHLblsZuo0gVWXqeQY/MPRmGdov4Pjv9MiNZLU7xp6t/snGnGm
2PhM1TgGRKfDw7W0PgQGVmhpEgIAmTiWC1FwtwqTkOff1SVjmd16rwhdH3N+VTsXyZmJbwYtTiss
PzBU+O3m9vp6BfNlJqTV3TiLGRHfLyRO5txUNe6hYwE4ylCkbxR33EaCO9k/L5xzW+g3765xRHVR
4TDs2wR4pCYjsUOMhatIpKhnJr91IoJfhpHHKe4jConbOaohQ3npV7KWvNUjlaLfQj8Q7ICoFFdV
L6Fg1qdiLdkEfsgx2P7XczBIjcYMacx5ru3JuO1tqgBQTsrgVh602BvDScvcYdVx3G+hDKNj9rKh
adw3QoUJ54euSVkczi7rTBotqyA2EkYu5V6ekajDDPAacFT33e5gGh/ZPJ0WAaWtc6/2MY2NHsM9
bM8J1kXV4qedbXAaYPygpM2L3b2lvoGi+Vku5BIXUWfiFkFCvY7gmG/t44xGhIVHoJ4aWBou6SjS
XoXxU1XuPBCYMlQrPDjclyjvOAQAIPdbxmLvJcWsjA1NWW4/+O6U920iL8XfnH3Mcr11KkkqPXHX
4YhHy5h5geQGk5ichgRAvPKwKCA2PRXNOdUYyarlHVjR9gOOKyk4XyYg8Hk4NLOMzm4rTw+M+WBj
2eJRZIiPSAlt+nScrhWWA5uyDarxezlL4K89i8HgFrgy35rMJF+KzfDBN1YTWpMcR8mVuE0Gu3Am
xk8MIEKxyYFtKhelJp2wIORMpYQPRZkFWjQmJJDqOpm8mqjrspF/PG/7yT26y/QBE5DHhk9bPKWE
EA6FGaTxHNRFe/+5QF5q+k1YOVLgu+xM1+zD0mlob6GDBfRDZbNZZxS0atjBTb7ELhnLwHIBT69b
Jkj2lS7OAC2P7mbgxv4dCs4a+AAGmKPbaX4J6HN9R7s+9jxqex9DCLkFgSmRyhwDqC6mCu0JDBZZ
wyxmXmiwz04VTlC53eYRVaSXoB0oax82v+VQTYhuCscyUI7YRfRz1Q43YCKKh8/tIiq1TnUaJUxU
GV7ll5kllBrpNTzdvi/lI7/WpzcWyd7w7dVQHmPiPqrJI+/BCS/Llq8dIKLb8Pge5es7l+XELFM8
oT3nBWAiRyRVN95B2tcH6SJCeweIQVa39ikq5bfKDjfLEb9zH73RzZMZFz3pjrHJ4ENh+D+Jlo5w
/fvGHY/8gMinCtK8sE+kDQ9o0zYmyL3jLsCfZn30i4tdBrSXMQrWQ/05m6hDN+vd4prgJWhjDmi8
w1+SCdvmw06twiRkKq0LZDDFpOVIgVBlycSb9D9AqXaulY5rEVYL9VbkPG+KVnit8dnlK+QiGdFi
7YOpRyUOQWkHkbZrmTLTe3ddImM9AxRim5rEthriTp0MQbb1M75oVxzpZuAwjMFEGWgx0TMQWjhF
OHCG/XL0X7vjy+bqxouVjBd/Xa8vbBopjRLuIq475KwRB3XVdhgb5KqAnQenDMi5zGAIcXzpEbmk
MA0jqqBO9oYZjN527O8ALSuI9wCqKsIvUnYoJqxRJ6SILClb8IhP2Gcy4dN4+vedXwwDoBR6DwbO
epZ5M+GfLuGUmCUWvJMuEXr11M5pN1psMQghmdv1eARWoue+b8z/649689qbIDBs/RLwofJDkwgg
T+LDCNvyoJfJ5y67BsW4u+WqBoOhTCRFeZk8rOfmgdQSQiEXx+C4fTm0B6O60IzEsRUxqGjFF+RG
HZIs1nEs4vSTbicO1G30SJzWQGGYOeu+C1Skj9/x0RILJ4QfHihHu6XZgfa8oJ68pMpz0Zq/Ezr6
0w5Oc3pEGJD9Rl6VO/Zt3STJkN9fB9ZnmSmQ8Qj2ZLcqyckZ9kM2t+rFujKuAHec0DYaBsZQYrtE
WS0ZaGyhMP3ebGq1y3aIvMS4JklDQyERT/2e/H8UdrGN4xnFgNAI1JtybQeQDaniOxnPLpD+6lpE
1Jg6rNu55uKO5zbuhc25Krun0MvK9MP70dCoaN5exT8hpPyuwDz0x8s/3XwqT3eg6qbTOGXuRtU+
AauoouFcnaAbMhUaFDR2dt/x8P869AxO+BxYDvdINZN+QZ0aAU7B7ofPfoFaJuRFG6NCYN3XNf6i
Tm870ry+S7UNaW1/z/6y9vDm3/KJPla4Lzz/Bt275ut4wm9SXc0VM/6F+QqLxgaQY3nO3q4ZcdNG
CIED7qLDBTSWuV3A9zPykbOuDsaqOD7+9ZAIFFrLgC4sBMD15J6UJhpf7g38gnewBnJUpN599W8R
f8IjiVxYoKXpKaeVLgJZq4UNqvQ3ixW7LzrR2tq2Sbx8W4KUUOORoilSIBTyf9x3R14/QuQ4bjIn
nuHW+ZDlAlqMSRiBoEgVeV7Hp/NkNppKJ152cVdM+znWSwOFQGrfbI3FgccLA6zAAoXwmVak+tp0
FWGTTYqsFj0L8+9DL5q8+PXhOgmY5kiA7Yslt9SWOwKJmIll9hhI8JGL57yhmby4I8u1uF9dF/6d
QbEc2pQv2AzXeGO53mCLG2BsjptEZUrat/VYWl2R1HhKKa4HP76IIRRkuKoblcKmrJA/Fm3zNya7
edOldIU3xpDy6pvkWB/oaamDcGdIczdFWKE5C78J05SIb24sGYYDLPq87ewyDmBj/85dM53Uxsxu
YZaSMBRywe64oRFSrkjMw5rFd/yyzAi8Z6GERxEJZ7cDL71gcfo90w1g/AVUaU6Y/t13dW63CIpq
RMPSFMtUlz+daLMlcxn82Qo9Zku7bCa+rmdHP9mKPGKUbi2e6Wz72z9Y0ZnTa+Ndd72ATtHSZcTU
yuVB4zHRtEdY1Wb0mSN3MeGlL0GOq+M7QwBnG704gBZHSDjcao3t23QudOxOKUYbzz+Gcy4aaMDP
4pSre5qfex/qrK9/lCWvMBg8R3uB2FdTO3H4L4SGBNTGThGvNI4UDa7cb2pcaIDN3Zq0mp2+OpOS
vNVayqoN8HCayoX3Pjigf21f4Z+Rocb916lfAVc05nQ4r+eJsS0UdfHay/50leFEjMfV/MQ/hwJt
nYKOy/pxSY67feSDQWJgrFIvXDssNyBxF0aZRql4kl3it4HSYhRfnqd1EAXcmhQTwui/HZ7QgLBj
K3Tei64M/K3Xyqo1SBa/HzGAk7sA5Ql6A832Lg3j/M8J73ZxhquJJXVO756qQq51623m0p98U3Iy
jO7z7SYwbtUhHa3LjmJg1huWKq1dfRuG8Nb2J3F13zbxPQTDTfnDrzNPKrURVh8Kf9aiPR8iIl9C
cF1AOFGqSTH+eZhuRqfHIPIw3NgkYTjDwzpE1K7v2nV2evLMYgdRU/XZJpE9LT1FcMRo0RQbTOeX
r5gglfqvvdMtPEza9DeiXn2Jf2sVoCRhfJZpwdZdVgzCowfEkH5TveJ+6o8FE5lE5hwT2ova0nzw
r+zqjQtjDV/9YxHd5Kd89GcwI5wyo8HQR0jAldfy4ldNMeD2T6vbnIDoNwFFPyruy3h6MGxaGGpn
09Whn5ZN5qWGWg4Viyz/5uGuOdy2muu/6Ezc+yZAJMO601f6thMR6rEYRR3N3i2aMzpSDy8njQkU
3hZQH7t4egd7XtZ2RXXJBQJBosnQqcdz85VIFh60mCYXb6loB7B3iYa03Hbh8lPC1Ppubvuz4+rp
tzF5cC8088n2rYFWxgQ1/YCeLAvB07WxbZB7ImC8p0IF2gZvYUAQcAW7jmHSftRpHJpXDQ1J4Jbs
6WTtqW6dq6Y2PfjYD5ZhaYfi/FoGmYLH3dR3IT6EBVXVeQft1vj9mxWxjprKz0RNSSNKOA3sTq7I
Q2+or8VtDjQpVPFeBoKCp3aEj3guZHodSDS9VUuiWGe8ziWhoxkNX/ANNAAqygiSKAwYZXuE6eSk
fIASxmHcTU/ByDZ4IIysKwDt4bHTUZtdtUG5uX5OM2ttjZm5Zcdg8ftm0p7zL+3sFL+psF+X9/bI
2VdZs0tet5ZSBurGOv8W/AaLIObPRsNhFKCmCfgmpWCDMyyO8r+Qf1G3z8JmfBk7Xtvgug7AJ0g1
DI8UgCql7F/l5t9/GOduuAFBdwjvp8krF4u6hPCSwfI4MgHa1CHc3/eGOJ7KN5z/dTdOkonlRkmn
iziSKtUyoage3ihaCc0mBQW7Fgkm3aySecq3xAfa1cLWwnfRDirU8ZdTN5/I2VEgI9d/osaSeLby
fpAy36AI1LCsb089JG+uD7a+s5843+xeYVKAkZSWN9luWcVQgfijSZSnq4UT+T+semOD2ZvCaJQm
xmgAUhTzZGkM7zsaUouPaE7VgSe2OtMfrAzK9r97PQfVnwN0SY2TWjJTetGTDzePJkyqB20kVoF4
jSuzNgHDc3cP1bplk4tG/7X+hRZisc7riF3AIon9IZjjPhL2kDCT/rtPcWTRYeOxtLVog1R9clpb
G3cQEFauDaWpRCIdLPhAdigoP/qwraJvTeCvJuin8Gbb4SUvQ14ubMkKRq9eRuHARDyz3Nzeb+jh
NdeBWsxgHLgKp25QV/E6o3Mv7hCyw/7dDbuCYIEnDbs3IF58L5hDBHTf2M1f5nJoP77HJljcxVqc
ZXG/ks913E89cofqkwT5LTEEY9Pe+rILN3PbyEjRraFzGVVoPNAUv0JZ+B/NpVavX3oeGzlBQIaZ
AgUGuPOEbO/6vUtnpGKV+GTznvvOpBcpLdeWiGigsVIxCkG6CvpIcz94QFPRD9fDZWTON5i0a1Yq
VwUGQ+8U7qiQfiyPQyTG9iub3LFJFJanQJj+PXTlklMRzKaK8Y8nqzrGZ1PPtV688e5M4vSXNoU4
xfuUCEFJKsBluewjgRytaDAeUqa2bMBTEaGHsgu7ZeCslkjZCclGg1GHZTwlwSp99neVK9ssJWLp
E8WYDZp5QOYXpmmcNESgDf+YJhWT4tlw/5iSAvy3r7sTCB3ItvjAAsOch/O7AoJn2iZ74c/bRyOR
UHOKDyJDai/gw76VHwi58vv2l+twil1omn91L87tmAzXV8lmQB5/TicTOyqxh/FRuNVYH8s16dvd
xWjHV6xkqIuLOFM/iRAVVGMMHQhBjnzUS829x8mkTrYADJEl+gwd5Nukev4SyUjuGLaSemaW97M8
iO2EadXfNbrGI/vhI33RSeMlLp0+18WkkklONxk35kvknQ4P0ouI8OGjCiimqOknK0aFh4squkq4
sFW8nf9ZuHB58ADLgcFQPeIDufUlQMGNhs4TX4IWHZt3+sAb2mIwQCsDcQqtaiHpRsqUjnVZAfCi
roKS7DQ60UcnNweteUZKce9lH5pcrR8F8D6PE4zmBG5D/v+EqAFOERn/bJ8GsnyYvC8UcmJlsxLY
CmMxyiV93508lQYBNfnLMUSv1h5KHGDkG2E9v1Y6ISxJnbicLesofVLl+Vhdw26SGew2rP5E6Yrz
riqifN3j0JY2dIohaoZ+YwxqKHMDlkH6KIIutZDfaN7cTL5IF6rBhns5xnAzeTbEpRd04ED/gQLX
R9warhXC8hVuyaOOOmgKMn7gLgua/2mwoo+rDnALAHCzIzfx5gV3bHuQBidAmbEObk8q8IhtpvaM
ZvVKzEwVskHehf/GBYycQ4Hink5WRpYXMqjAqrfZlVvp/MI4FAPlPCKPnHl+5j49HppoCFztZncb
2NM9USdvJSzDTh9UrZ6kia5x3H0pTCW1Xri+F7YgTP4C4F6/PkjH4Dd8vcyDuB34ppJuOPaSqlJw
L1UYyO1oO3IOyKK/KgbjN+pUxsImWsix+Z0Y2akBRDC/t81Dxb6x8skKaUSARLCC6YpplV8axWsb
nqtCctPrituB9AUW9hgDJ/2EjywSZEzX6+DhKvVD1qCx38AFawtNxGkYWER4iirKRzcoQ2jYQfFX
ywc0sFpoqoiLIx3MX6ECiucKaw8KURROoT7gtiN8UIpA7ZZJaEVDkj5bLcVl8KXyu0NRECo2L4kz
2nZoNQXY918JblAAAOXyI964ojUfiFwo+nKA9K6BpL9MsGs1UKtp5JyxB+VxrtzoVS7VSrXhka7g
z+WucM9OCbK94EG9BIZUMApTPr3q9yTLTN58UoI/4B4SQ1MfEMzG0r2NnN5W/vnBB4QpDfCkki/6
xh+hCV5Axc846YNVUZj+fC+BQwv44XJoTV6dKmCRUDbNwaELiCdRCIw8VCmUxIuSYOBMVIHdQY+m
FdVUdxOtjmpGEQsJ7uXtjH4RCR6oPpQDzrJl4YRAnEe/2FNu2FJnAcl/rQPqZpOvZ6OJrAnpscD1
QP3H5Ws0myXC+ITIEthJ/Brm7ZkcIfdjMHw1ltfVaq5QrANgJkWJ20iId5vAWyuLoDA1JTENl7oe
QGzTQG+q0zSyBVIIio2uQ8m1DTqeAXbav7YxlrARivSgOGUb2FFA+ykbvWAwTqzJyx28rY0ek8B9
j/p4D1mMu8yJHHU8kL6G9mTSZvJlOhtKbC+mM3w4guRsrlDE4AkYx2K/5uPk8AmfvVxEwp8UzIo5
0Uyn8p7FmCXRlHSFFDEa5Pp0q5axqLe6bc5NK2M5lmoUl3MnqSF2tDxaRY+5bUzjeLX3d+IscaUh
HD1vWY3N4fxH9+6g+p06xzF7BOFLr0pnG6M2778Qygw2/LOKih0WXaVc52sYpYgH/9xcRioyc7hs
QS9SfbpbtBQoqYJmXNQ5kcYXnb2GGXLOUO9gV3XDi87n/jUa0XXhchgoB6aQZWlChh3OztAgJSJ9
41q/br3rkyQZEh1AyMjn0uQb21y1N3rLuHwPFWxeNG4IY+HjF/+rEF2rl2X6ycRtTDGbJN0prACy
Ysk8OYayD3PYF0M6tApTdsraXGZQNfjji3FtDkXB+BxWyvmAWJ2P8SiqhvTHbCfFdtqPYb7rKrQJ
6bbydZiHlwDbKuoyKqmZSujnl9FasfHAmB9XcoftxSY5sLahMa19A7kel3X+emVArBZI7ibv3gWx
+xbboV/0CuUjFq9h44wpSmtm9vbwaN8HSB0lLl+cSPNHTPpUxZSEoW8t4pWFoIOYgWD1tzew/Cm4
xTGykp0DjTXpIgt9+MRouOEMdsyJSxLDjXtg7oXY9kb2arFsUIXtTwW8/835ZphHe91K7i3lvkAw
LVdQFk9WEKegBM1TOxuoy/XhPSgjM0tqBpeukEao/rbRy18wFSIujbSJFbZaPnzCbAEHyxBe4tHJ
cpiNlwcHHFqRY+uGAUwEovSFSzZr/SgsefH2Li7aDqkYgjHWGDOpLjjv616Ul+W0JmSeBEuahJfC
NjioWEwQ1cGSyVKEuItw1Jw7ozhLD7QrvlBoVHMofsYAFII/0i49Pg3sVxRu+e0hsCzurShmAowS
5Rala0t7yf4FOp00oU66IBqmUl0pYErGRm1HdQVLkxdD0saMMG/EsEfqLrPa9nPaLkaYGlY8UR2r
tsDT0a7POrS3g0o3VWiZjhTFEVYqpRuuXWDYd5akVz2Nqf/TASeWZiMbsw9ur1I4vrKPWS2qXpHG
0l6WZSeTnGzs3/Q5aEXtlcrZWqBSzYrHvZXmY34QDXr4aYQRjNOfJeI90w+hp3J7JJhlnz98DRw0
/Z2Np3h86aqQUcMsU3+yUOTo9IsY08aySJPyLnrUNholtkk6EiZpjzRgIiTxbbjdGi0HyKW6BUay
onVTQcUvTj+DH7oyJKVIB9IjO7AsdKknpjVSyCM+DSpUn0yGLU8fOmOIkQqMQYIUJaiO/xE1KHvn
ZsaQr0s3QeXcJyTX677EewBtQGPopHmMcIGYQU+zyxzRD/FLVUFvBzXgtZkeGy6qLLujywXE2QH7
+GI/WdO+R9rpdWMDd7/WrrlpPneDilTyIf2b6FnFm3XQPrDDgGpbBBZM0BDn9tmYaKyHMhmyncFG
TGoBEjp6ejs0gidfbOecIV7qByIvNUEOyPL24c46SYh/i8mRcJ10VEjzEEDRf/aIa4hOTdSymRR2
yjXfKV8KyjowFCbv64HpmyP8Leo/MheHVi3XswN3V2qp8+LXVrooyFrcWQtnvZ+ofNHp+dJ0CSmm
rFXvwSbLsvZ+08BRBR8JWsB6fahPxGHYkmia4kPeGA9RQNiv0cgNw1imNAniuclXjBGhPFkLyYXD
Uev73MpjX9p3ReKPiGGtC8LkfmAW6Re4xPHJvQ2foSNnsGReSRk1pIoUleBxd04pdyneU1MdlEZa
T6P7x/J+2GmSQ5Z6nS8CpWej1Q85C1Up1vZCh8JVoC6GwDCMwzlcZq/silXFd4D7K00SgmCHSeGW
d83lEEeyxsch5gH/UQHc9wwOlSh91FYYCSrTut9so2PFPmgquBKBriniMQd4rAGGAcNrq03aTD2c
dpUcQ7k8xSJN3aI5TdKJ8tIB3NNliE4eVIg/5dxf5QecGJU4j1P6/FSPWUurlLl863qSP5roZl+I
xa/Yecrl8PUg5TFwjYkSJbI0asR+C/qiyqIrP9PsBWKKteWD/LbX9TxszST8y04RM9DHDeQ9jHZl
is/mk5ApHIXUw8G9aYqlFyoelhsqO/WWUskj4Drae8wCcjgG1E4tgY1kqIox0mIIfAKEeHC5+qd2
ohV+gkP3T7ifRD++DfZ2tS5Zi1PD0cot5z8kC2LFEMzJ61DMj8o9VfUm+PDaMBUJPsLkUae7EIb9
m+y3rMbxbISazcW2Fmuzk+LhWOiCixWjvcTE+IyZdtSd4snBxe1XBOhHTmznZIz+vZg2bv1CB7OE
F4DMIjxTtBAu6F5XcKH4sYWl1fS9ZR8Ki95n18TwApc30abqNp4tks3ib/rR1tGN21OKdoTdNZmF
QnPqTkSNTUaNYcPd0cl3SaxT6qPmZbBijDCcH4KMQt8CPfxKsJ68mD1opFE66/aEjQ0ajih0B2CO
C6Me8IsKBP1oNV6vueb7rjaLHGQoAWVNghvKuVfIT+EKtbZqC0yfTm8jTsxzwVNWGuItCpecQVIq
1attUYj4cqJa5bn9aDM4bNr8tUwn201l9DALWJOHg9ocxL8GNr5WWYdG21DoajsbEnbDukDSGsN4
aUE/XHZ3Ufom7gZqnKVSAXM/4RdP29Z7zRFZDJCuJtNaYGJciy7p3pT42okCsPLGvRrIniRlALls
DIR4+7kNnxl9hwQH4zi3uq0WsjwVL20qbv1JX/VcjafFwf2XYI+sEzIEVDpDDp27mpUIPj+Rpxcn
XUhtz6nJen5yDu8R4TTZud8mHuthm+UGHMP0Xm03Vv+DjSBVo3I0mrmlR6t7Uj5NWQI/j/GI3SqH
q/+lekiuMGaRvFDdXWtrLSs/GKxCKYZQzIdA5z1P+m+tSsqW8Lw4AFyOpYFRSA/X9qxXCxneBm9l
VSPLtyz/SkiLTpNcBouwsjuZAO58bcL4A4vpcXHQSPC4IZZ6OXFBrSdXkb73q55HVHPvEiCbjTka
ue98GvLYbyb/AjCpGyfklWOiFwkFgzhnc2oFQ2RLNwDzIspVvzhAWUhvApU7R9cEvvqEV6Zr+0kP
gN1TOG5af3HdPdArNv/CnYqu710dMJQb3ze3pP2m6ZF9hxEgATAPxfyARxFmiMngcQg91AUzRm36
fYzptg2GNTUFMujYygyUmByrXcB6OVrpBHZkMJ0IS1uLcLLm22vFkHbeXhnZ9S+Zlanoa6uEBrUY
9+PTEDsxcjI3F9w0r3+VDSyzhRr3q0mvXHUUcgzdETJWd1f+cbi7L0gNcQtSaOqZ7GO5z2NUYva/
nbft4Ee6n6t2gfCUDTFZVyRdFNVaHRnKO/rt3DmwWSLSB0YriYEGcNlD7TssmizGwpvwbJjd9iTD
SdB4XH6AZ8hEXuKKWPXBtTQXISPxFmXiMJs6nhwu5SpbQWRJbu/8HwnbCnwlUYbHSaTTb3O46inK
DOO+DnwuV16XlUVUGwcHsphgblxzWklapUzGkKR8z40sHZaPUvMgc/CHJftIszNOIU3VRvGSvG8Q
R3F2pL4dpzXUH5yIApAb5jU2jZH/3xEX8NC/6h7iOH7R8YWSlFP/4LHY3ru7AgL9PS6SGMfD2wq5
SmVenDPmp+gCufzhwVRS3bJOMzmpjgYIJ1jUbKoJF1ABkf4T957su0b6ODyJs44pF5s9iS9u6+vY
30tzil/RegqXgC/0QOfqw5lJK1ClmZUMI5N9GlnJttrXrw41gD1sC6HHH4o9PVQVDUxc8mC/Kxr6
n1h3HvxniHJ1e+XdOnAwknvUOlGhmATUtHh/VnUBiioCY8/KGpz6qVXnnEWnZB3wAlTCmTvD0PYg
N1IkvpzjbJ7XV7l8FRUZuMSSpL29dZo3+tcSMoc7g2dIFahw9mx8WTkYnnZtYnNaTs9TjrLtp5oi
qVnyj7O3Stt2AtiVYT67RfU8Hol7VI1rGmuTGNVTTExuQo/WYQSeODmh1tSUkEKTWUf8hMnVUcaa
TadfspeQHOoWxEJcojdnu1uAr40fa6vJUGIPl43Z4/CCCMyspZGgn2wQdwM1JOM2okx3cvnT9K2S
vbEhnZQj6xNxYa5Rkohhet4NC2nHmm7ngzH0JZqruEICBW/Pm1GcyhTo8FkRMibOy4KHYKbN2eED
eW7l0Q1Stabl4cVpHqGDlE09sw9xfCHB9xMZRjTmlSY+OB0Tm698mxHL8oKO2pYEqOON35SECQeZ
8Xl9GL8nNLO2+KmS+ophmJI6td0Q6N3HYdkL1lfBtQJKKyWrSq0EHRx8S9a06er9ojTCj1yVvQzt
63IRmGCfnCVKciwTlsI3WRM3zxvUiNukwf+g/vV/pjL5YclWuVRCJg7dW+/JdLetS1OyrTl6yxk/
5qMsTEgl0NStpgh5BsOgJaQcePaMM7SkBEeqW9P6rjiKzQcMpXFZEhaFkR1lLcxFnyHzXuZMd6QO
kPPbYtb8UzrHm+lBwOsQ8BcaN9DtbjPYnHj0gpT4sMUs0xxFFk+Zppmsk1Hv4uaQWtdJrQsCtV3Y
MNL/8MNHpj84DNs0TchscKmkQi2zSPnZaAKCyE71taEjfkPV2dPl6X/jg5ha62d48oxUhJvKuRE+
AJL8eb4r61fQAXUsjtdHF8HItRi0EB4sDV3DquTKwgEg16VrZ4fCUfFBp0VS2ZXix3F/5/uH2ymp
BUXK6JTW1JLZUodU9a6MOu+c8GSpBAwV2ZBruR8rhtsJMTxtIC8AAWfJM+6kyv8tTxRdHQCpSi5t
WUiRzWDA1F7YWQb8nKoIkFHlVkPF6/8CFZzKwUQtTpgJNT4Uj8Qd5kx0ce3ymWKqVwKzWSeVaGto
7dLSOJTNSFo3stzDF/NEkTyIJMuWOwOnIMEXZFZCOnSpqQYnr3+3n8MWw3Ml9Ju7huYVZomtLaDK
1O9H3eFJxpjdFdxmULAmNtdLeWHB4qYLCjwGHwe4X+YldF3pfC6v58NboDgnlNi7SOsFZr1Lp26U
hFDRqu5/NKujY/WxB7Fn9SdHFA9zjJfLn6pwoR+N2a/q9WIwBnW1wrKbJBhBgXz2ZHnimQgLPkKZ
UlwU5MB+eiZSZnNhkeFZ2QGR6HzgohmWzHKx2e6tYmlSLtA2leXHg2fJQG04IF5z7Xit+f0Ox6AI
uhLxf6vBkPO1EzrMKsnEyLPZpmktm5DUyJnxDEePewJDNnaMWB/thL6vSx5+33Osx8nRLsrvqqJU
HDQPgNIaBjqhH8y1yhAqH3GsK3DQGp3WgYwoelZDffmHqtrQVOaqBcVA+qPc8U4Ll08AKBQEuKAv
Tgli1/oEbBNb6sKxLuDHApO1edb8CwWehPrmo2MtQ8aLoTkf6kLzXwQxePZLdi4HI1Hwy5FMOug9
OyntyAQJeePrM/iUtRDK9bsQWiwCiX5flHkJFhfoDunsVHZlE4nFlKRgt8D5txa4yU4wYy2+2Vfo
WRpKH1WNTEmPvRrxfacxKGjy4JzJV6n71rzhbaSCZvrz4SMZU0lUcugfliHB7YBxeSXLmkRAhlD2
U+YaxCEJjHN6F15splDG1EbxUXHyWmpkxvXEhGbYzI46Oc9IJZFesi9T96V0dFpyk6T/cZg0qf3G
BD1X5tM+Mu13hUtmlwyDcHoAw/DqYtNF7fg7h4IzNWrW4aYj9JGCl5gjxioA7rR1IsecrdzIJ9NN
i29mZhg8DbVSXENN9ysrlJmr3iCNBw5GmXayBVsCHcQWTLYmxpemA0K09pFZblOZ8iYIvFBzGC/p
THWbeqIGVIk2a7qOSIwelf7/nGGp6/iFF3YDNyvVrUaRm0h3El1feAonIqWr0DUVRLIK9lRLZQj7
juo/0ioOeVy7ePDHXpNquj3hS9fTNZhXtspSa0GlRjSroexCZkZDdApyr2LONqyU2kxJSr4ZpRTn
/j5CrX2uAIaleRMEdwU2rgWtkU5Zew64NKsnvXUZXnUedMK50pAy3PSoJrhP3iBD4Rdnatp0Dx8D
0jJbOeNF+tfDHYJ/phVZ7duMHMb5Mc2RDnCdnYLoqY573ugw8wIkMn9YWi9xnLkAOutD26MzTy5F
F8CkiMfxVYAM5c1EZ4GJ72UOMOkRh389a4NkLAqDeKn5irtz5xHlaB6PWJGmVfzwLlrbwHkAxoWP
LrSiSV5S0FujyyRluxs0XdWjMcTeZ1sWJNCs52Mm8SWUVCSy/CoyGBKYHl17uNjcoIc3Sk1WEKE8
76LRPHGr+aGvcyVAVucRJCy5qsIg9howRYXjZeWAPEpjYQKkmhndpydpmJml14qYaUti/ypfjQi6
OIR3EoWgpzUSLW1yCCNXVzZr20iT8jET+dcy0EK6xcVCGobaR2KSSwOZbuwULykDaWPB2ovmVzR7
5KROXWGr/u0B1gVy9kHdXhodX8wauL8kGWfyml0mq4dHOs6rA8sYXoI41QhpcnCDbyvi4ERUeMXz
kLeKQ3SXt47/UcHmYZUGsuCzfcbE2nDROpKkvlW4mGh96jBoF//h25iMR3ng3pxhBjQqTeKikf3q
tIQth8FIX9r9iiZ+1F3R2wIPg8Lviifb0TYwGmu/TV1Jg71ca/wF+3H8M0rEnDoYBx394aqZtcXq
SUJLpzJTrZhU3DP13a97iUVTzlq9hcy3Sbcn05Oabn4edfjUaLRLJ6IYuITGwUu4K85nyfny+nXz
nq+avTbwjjSac5Z23qXMjAuRs5M8FSWBPwThSU3Te0r3Of4X6i+llmGSKUQLpGikQ22kcCdQyIMT
HcM8k/X+XjJVTkSjFaVp6wBSdiWnIQrnBIo6qY5Y6phpAdBS7l8L+zMDjrV9+CfdazEg/eLw48st
88yY8+XXfANOV29Xt/zO/EdQCyf+k/FPNdtGugkNVcce164Yzgw2MvinPj0p1nTalZEaWmcRsLaT
BR+tYOcUNfiJsFhnndR5SN9IzPBTzI+wxdn4q8b/BUPFOoYF2pQhhY3o43zEJ+YlX4fkpZv4eMS8
/QFwJVmC6S9SBIqOVPRQPVLEpupO91TQdfeLDe+VM/jsI0Bw49JH5IwGFmn66WTXiyRMoMz0kPD9
Z/do149pqQdStOSmERS+1X0gp6+t6gqXIwjl/H8y24ofYKcfXIdBu06A7SxyTnx0xWkbjm6Z2161
8OQG2ynfNh78VXvj9ChDdcrypnelIbnU3OyGO4QKoM+7BV+xdKtbyIRb31rAH/C8asHJs3lv8CGW
fsXVrKP3u/Jyqy6x9OOgL8Z91wvxn2/GgenCDg6X99OacB2WIbEb/reyLBgWAX25Buom0KnKUTBE
5/FKxbukmC2ImCgUraTvVoQkqGzsb0KD+2BCeK8rm/Lr2JPIxHfKhkiD9SfBDXmS4VrV46DRKU3A
MX5jkM3foBUSsq+fC9Ygw2GjQEnCmlNh6Oi78OAgNdrINx0QQN0FXhDhqJ1kv0icynfwC2T61Xkg
2j7JeURIIoqgOlvDRjExmtuh/THUtoSzq+vo8/aolEKb1h33YbixHug7esrLKsSuxx1qKhs7ypZP
GZvG0p46aau4F2V18E01PdP1CZyYd/cu5O4HM2SgWG5MsVFw2FiWSwtLiolYdYZHao+8hV6Opl2V
lIritMurB85/GeglGYDE+/Bpcmi04KEm4BgXDuzqS2SCYTPwBISd6JBdozdpVLdBXK9UDftUWiFc
YXJodrJyPpay9Pf6Uin7RLvgI3yk7OhWv5dInIYi2iiZW2HONysZmRKYimzrPLbPg5uMSCu9Dwb5
bfJry8rkECGfPmBDroHRS/iozaVxc93SQHmGm8nDK/MOLRs9Nh33EjVICPL+PAcG64TLPy/A8tSP
d8rdUvPcwPy2CUweoBuaR5twskuZn7f9yo6R4NDoD8L6yaWO66NlTFpLOAiAaS85flkdGjURzrho
6njq+F6ICdWJwnBxRSvDJggN/7CYWR2hRWWJ1Nhswx6cH++vqMIH3MqVROGeH2Su01iklIUO1TgR
1hXJXVDn7xZuF7updV2UXlZE/eodeV6ELArglIdD/0Np0ea+Z5q6XQ2Y1OLPWPBsw2Tux/koHuTn
InuaR0s5xjSPVCkd1s/Tx+f/ZD4jH6FCJFcRtMRALT3nEnJ9ZDCfFYOSBTy3jFEz9QF7i0HA2a9x
DYpQBQtpXkIauQT6vm7d10mnXM/jaTZW1xKHaQEP1REiGbFnqYDp+18VSRQkGqLquuSRydhDN/UI
dFaNlgq6OhowwKWFU5MkjocAxLz1pP6vPhNfWyGNKk7TFxqFz/q8/Sfg8I20Qkn0FFuE6GiQRPc3
YnlV4fD8BF+bQf8DdNCc+GIymuZ/xCt3DWSCBGJu4AbDPV3HNJZj+RZLEIU9ISG/q6tWHfTJG8Hg
w8Z8TnIYNxmD72uYEuQWAtrGCnsqaxFVWDx6UxXFyv2mZmcur1Gp2k2cuVt8YSlBOQE8TaCu16wV
EoxN1EF+8L4Ji9vj+N99CvWEgj6yYyiAhELz1lCJHSJCotmPgJJl7hlXw+cUph6Din5YWIjOqD6V
/uKYk6WRh4QmdCIkvAltmeToaFTCwuu7eG682ahSnIFOnt7vRQhMoxL6psmgA3HQNa0uYtpjS4sM
yQ75ON/p0RGolA1FgiOOZ7eEEvZ9LALczBf9iDnNYEqefeQfawhnV+BPFsu5P1pdi6DQF2uxY4iD
7tnZFdkhO7i4J3Yqk4efeN7OG1O0gECmJI60ZVmufXinXlCKxyoSLxUJCpj9G4U52VrXrG4nMu6Q
+TjQ1btoOEBg4CKrlFJO6v4ajroNVc4u2jXgmz9p08ZnEEd0y///o+zDpT3MqTbYJW2nPfmJBPCq
n4OGZoPfCnij3LQnYHfETgfhkCVWgDjxLzOiDO5Vqucz1bJv14wA1UF485cPIkhQGxjfOZNvFZaO
OuQgPHdC6mgYG2wWlm/Ny4flPjR6+rapwZv8VS+pRPH7Yf10EBiOdnX5XNdvIJoBQUKxrxaNDxLk
WWJiE0l7uT+NWyN9UVZz64xJrJeDxWMDLZknbxrhACzTyhgGDG6w6i12dWXNg+L25ayG2kBV5VoX
RoennHMu0JyheAsU6yQNfLvrpJyBs+v4tz0gsLRo830JaHAV8VbRiXbx1iUfQgO6n6nYsohTI+/G
Dsfks3Nr32Mqk+45GlOlunhl6lcU7+clRiVogLBifWmhaiNamvkxwgYn70YP07JNxfkCBJgxQc/d
kFeWPlQsWBvUvN4RxQRABpLYJ1mFWd0dqeKL0ffKEaxuJO+J6RMXpXRJEG7U5gA/JnpZlgcD0zc2
4wvd1L7S2nmnlln2ewq6WsQpXUhVUrNJNdO4v2BTjEoMys37s05aX6zfk+ofHRYp6zhsMiquWl7R
fNxhQRSjbSce8xnF87QD7FIdIAUEd3/OIoIfKIDHBrtIPJCu4oxQ3rQqCctiiWjl19AP9G2PNbEj
EYZaT/izbuV4R+joV9vEwWpuaWjoW8LzjW1uvEDL7RSEvAd2cNNjanDY4OfndDy3eFIno2TT1nSl
52Nj2Iz1Wf1PyGU2RCf10TmuWczLYhfo1YjLORiU9tDz6Nka9TE0tAZHr5huVfw3tYMY1hB3IfjF
WgiOsR5ouiISHEU8/DleuAyHRS6YgUqHQc2DRK2++Z5KeamMsG6emLF7c3A47Lx6MLZEGbhmVRQS
c0qKiy3FWrpnpL9nr7VLl9JEcF0LMEM+YoyJtzQ5GwjHqH4SrqfAAm755CmDQmjYOnjgFDZkMjm2
kTKcrj3w8FsLi/whtRxATLh0QuRyok4jssO/w16CrGkHXaTejXretU7/cxQatK4h91fGab+j1zrj
TCl0DnDgMlMwj5xcYy6CEtXFcOpsXkHDM1ZCGKpXT31lI25muRTrl6Q4IaIqwAV2gvl6fXoq1+By
Oi7/yl+OCmXyMEQUu9tCN3dlZzeQCI45/913++dFyH8LCyLzLqwu3H0xWD9pD/kyVCtGJrJCEi0r
sm7Fk8MB7W1DoBikJ7bXxEO86h6pL7q7f6WefEqF65EICS8j92TtA+k4zSIVhAmxsiZ5l9DGrxsk
NCoyTRRwvzL3ImzHOY1q8twMq+QxSpaLXTV1BL0Ul5htGp6NgPoBSx0VoC5/kIp6ZHZQklSYoLPJ
kvV29tlckqn785RV/ndWqz5hR++5W2/1McXpBVccm63lQe+yvzMMZAOMXgVe/yyJ5vcfEmT/ak4n
Y9PAjuAbAFoWffeiFvqEFcCa+l6eJbjvonRXBUFfJbw0ndt/0r94Th+A8pO8MervaqoeEYZ1Aeuq
tmg8idpoewLciVVFuWD6UItGOhyA+QPAIeC7uSRXSyh8+iiIKvAITO0NcFtF97zHRY1HxenRKGbX
UoyCYOso4oAASyM33S2zrm+dP7eDabYYsJC6DmigkmDHLip9hWrn1bGpwItENzANcFM2cR5/0fxw
tQputWgrffilDWQ/smARtpOC5taOkfIBAe4VWL3kDyxWySMdiECfOh0qxCAIm3ilCFJn52+HG5iu
BzV3bN3TAgefr+D+BceVZLFPlYYZ1x4sC0boyocFhNVqXaR7OqG46ZaKbaG93Sn2S9pFdq/GRr9v
7sqEnRsHMWHtsE+YR9t5PYSN2/+UiPKV/2SZfKcRqs1+ar7EmBId4Wu8O4BoFkOBmetZe9OgFLpb
+8OKYBPZnz+reQF36BVmVECFyDecIBVJvDlHzCbiyXD+Wp8Y0/fAwi+F6SGDiXPyOHlPEbKmWN5O
1VXg58E6cabK2EnvcAUSjW/C44ldQaLnLhdlhKes65j3ATazozbqELMwcDcMFRF2ho8b6F8XLA3P
zk484B/fhVO8/xLPbT0uwEt38Rom4t27bjpAFHMqQlyMfciRU8Imd95t7TySw9AvYK8pOw/JohN2
anvddavDn2ut/DzDlyFdtn4lrEMaMqwxghi7EUKSSy2e1flKHe+taXte+NFHqLpl/cEBKq8eNIIE
gGITSupYwqlyWlyq23hyYYNd7rLtMYx2cg7Kkt4tzQZaQPVUCQw4FzycUnGm0RXltW/6Q+T7BaUE
QjmgTVQrrhXxznw+fi+rTroG8YQugY7gpxO4TPC2U8khiF+Kf4dOA4fRBlpW2ba37CTMfCwVL6Ag
MA+jQaNZTYlaTbyvwcwjh4ykZ6ivn5P0IfTleP6rfd9farE/XpcZMcWNro2/RCRP1ficEN9RdDsm
CunCs9hvuj/AJASiUMuvWv7yzHsx9Y9LgaI3l0JIAh8hFJyGWGPIwST2h5Ifzj6jPD0DpWcU8tba
3xEw3kmHuuJBU8Rz+NhWr0AIiRPqOWQj0BO3WuaSfualee8kReHQ+iK8y/fZzN9eLr55JX8aykuu
Q3lFEGW/PuXnLs4U0zi/Xhk1ut8lX8vMLb2ZYG/WurpE1tt5eJNuFgTokkRZq2uB68+1GHBap4K9
U6AyNCRbQVgWax3CY1Y7EkJd4EZTgCsk+gRi+eWbVgRvxL1n/ZdpZ1uDHMt7QiySqYS/iM3oFjnr
WXixsMrKg4YehSUf2q+0z2e721Mo+wg7NF7x3yefQdo778dEaApAtnVty3Y1qEDh4hsik/vS4ZZJ
qjw8fwtTMaf4OnMYbKyiMtc5sfqwLuARIdNqe0ytvk6nwoSD+QIm9WhhRi606hZyPS/y0bQnLPf8
wFFE0Hkf0DGuICCC3lL2UKckhtv3WUc+Wrsj8+RHG/Uv3r70/v8bwjgdBLFmuXRmH8Yv7R/CoSD/
fNlbhNvdgEbDb52gBlfb4dbeEnw/XYh+AvefHe78hVnIXYOlr5Hp5vnXru+JJ9BPCWUG96B5celP
bRQKjPnr25k9D1K4xGPl5pT5SDiM8m0Nq4CRN2eYZJ5JrIMrdWeYNr3rv6E++NSp7U5/cHkxEQDa
J//8+eHRCE9SVlmYqA8gn0btCLOFwnWGwJh7aRWR/B466qqnL7ltjIKqQmqwUI0fl/0cotPic1Uc
NB6nl6o2lNBC4wnUnICxXUOxnkBM4qsgN6Gg8AjxctWCOpqA6rCKZCbgDbSArIDu3L2AKKsLNgGy
qZQaV7BAuocHP/IYQYQawfXJO5Y8xUOqLTGAdkqbG5lSofu8KU31hjI00M/BVfB6G5w00rdHOQuh
Gpl6f0lWKfqWgybKhOWGOWsK1bB7huzsLTxLDa6giFCfuLmLqbyROgUQ4Fdl3MY2KrnEO6xi4ewZ
RxeHE8VqPPHHcPc8n7WY4beU+DTEJkFmQ/6RGYkrmdvdXW7LUI8KQ7hJKpJfLgURe5WaImuySbEi
W5qUySK8jcD+WlCFQDXXYL594G0sB8f+90rCqk9BxhqCRoNpDvPUdz697GiVzN9TPSe6/R+FQDxf
0wGnoGDecl6hiChqdDtjZr3IsxIgwgj/pIZtVR78rLxzQHiWBxSAZZvTQ05cbNYWYfjldDfy7Zj/
gfDDl51eQk+9mUt9XamkHJN5QJu5yib9d71vjdOnZrszvS4nuOW/hygc7f81EAW8nkBABQsJidZ8
jzdgOTfChWCDFMLGHqFKQ1yhdfEEZfrFrNaJ27K8BX35OlpqBkTxBzALQP9iWX0f5En97j7eTOhG
zUqChZegobdyeEew29WBUs+pV9t4UHnmbCFtbGaxqTO4E3vOS2gzVIYbmaMMiXxOIz++1kDk3OxE
U+DNmt0MCK66sWNXEjj8yBV6YDX2t8oUPO781Kxf8KyM3BCaSi6qTC07Fc6B5M22Fr5BmBilFIts
Vn/wU2VCWQ+36RK/BEzfuVV5G48NAZ3dYbpn7qwDw8kcmH4OFWO1nm1TL46mF8Klu4xJEfWKl2+p
Axu0j3qWClHPxvUIFYvIzEUfUdIRtQfP2D1h1uSjMAlDLJAHkExRtqhz2U39TyegucQIe4GlcN7c
CnT6KYD6m/LVuDM6LcP3ZPRlqeguXM/dB2DzfuUhNeMlHv0fmTSW9r41WyRt6O2P6eVZoKgO+KEZ
q8tVT3LD5RwlQ85B+bZLPpjDsGkrzTfVDu9E9G2i8SgUedY7KmEbMYzF46px4GYlfVApSto3kJut
3nx9icU49B7bbDFga+f6l/XC4Hu0I6WrMQlwmy2JCPsIAEVPrpoIQBKAAw4c1pLMro7sBXwRYBSX
CGo5ARkntFeJxOwnXvhJetgjcJycN5L8UlZq5OroPkchho7VndGSQgFBsGmYlvfC3VGdLoNTHz9/
ymghLQ9s/KdPV0GFxY0dkP7siYXtxWgm/oXniqWYRgIHUNT7pfvXD6U41j6vABR0ITvFJ5JRqyWv
uMsGyoSGvYg/XvWZKPONiB73tonsffBheP4iDRhzQmIe5JVt8uECNnuUvn0tGNe+AX/XVDOv1TsK
/5yRjcQIUU2ueSGJ6yzgmy1l6Qf+eCRdB0M5C6MkCOae1cIwYonwOWGwngOe/vuJHaIsuoB2g0sS
GpOEdVSeEO4g7NaCd9kp4tmTS2NDHQtZhHRCXPxRDQrv8sX3/8uD86I/zbJlnkNaIjK0ltb9wmUD
9UE1XuZRoJxBWvqJw3wO+PufWESQp9jgeW2qkyNii1i2kSaY2f6wkU0Bi9k65gVe9jPj+r9ldQlu
43vJ4AYpRq+gxIMARzy1U8imwuJJWiNwSA1DPgGmtb1SHQEUUpmBr6w+qSdwEQG14TPsZm+CduW8
g3X0i+NW90tSmTqON/go3TuFT9kvzcxMXqmXMcJ2zbJoOhWBJXvfRg048/sec1x0QGUlW3lnpCG4
QiiDLzL1HQV9gGBnjM0Vj1C8KhapVoczEPdEsHOyhyBj3TQjtxj5znK+PJZJeUX4N3dnZGFuTcU/
bbRyKnGs1YtaOf+DF6P+1MD2g/IqSBOmnZAecWYa60rAtwjHOZkD+vUO8Yy5oQqyOGrboW18gG1q
EbrG/3hZ1LNfqLTsJHPu6deIedI2DIBDc8BZcM3rpR/pkPEOvK7N/D4gziP5z391xlFISEx7akoW
/Tm4PsW3U/v2qeqEwa2z4Thb/CXAllLUu2jvsRnR4TwbTLlrirWoS5UOLZH/IsjHMWyNMJLpr6/0
UOqw9p/GTzbQiSWF9hinE/tAvHy8w10EGncUEISGH4J0fYXXePOrnA1sl10lxdr8R9U6Tf0lZC1X
/sLfaZjl0SfzCvMOSSUCCuCjARg/BzVqPe9wjusGP2i6Ud6/5ljAcLdL2z8zpH5IJ7XDb8h1L04z
EdjnsQ5mytOPZ3O5kcSX7OzLJ/qrkiuqQec1LpFBFHuu4LZC+s8wd4IDcYDfsjoF8qPiPca4YW9o
nyBhfqIb8E8ETgNTAUc1crfHPazMVP8zC4dMcrJwxaVbgXRmBuYFAWr1skil5Qb+DU6iD7lcVRpr
8FIhYPL3z3BUnsg/2C4X/YE+XQjK57X4x6qGVaW+FeVzXEZDJyHp5PGG5rdgvhoJOea+ct6pxkLk
VXGYp5idK0ysJcmPtjSkshDaxZrwiAz2Y0zmfLQlcNaVe9d4afqEGvTb/vtkWaQl4onHERpZuzvL
fHDMMRSg5ceisSkgrYFaYS75nEk+uDVsVWXf/SE8c86DpYRx85GmruvT+0NK+gUraRsSwxe3kVEh
xzi+5E9Kur834LAVp/ZyurtMicEDY35zZn6YVSKKnpYQv+tTrMGlaf0GqGlcv+qCWOUWQgQU5v0b
eUglqxR1vmjX6grKFNWQAkxrmAUF3kAmu1In3opN0U3QWR5+ZfBQPpO9Ww1CjiB0n5q2P7/kwh9b
RAlJD6l4fnit1T8uQSGYfqoLFmFInhjQ8NQ65RQ5KwBlwZmQANgAsRtJe50hrE4rwtDA3XZVB1vT
RsKUfAaVKW1DgEQWyiENEKAvJCUcy9YRc54fyvdtfrUHwoTj4rydIEfvbqta4yB18CMg7YhGmbHO
TsZlDvAuY+KarSuWiWxYJVxHW0/OPDYcCNsBUD2twbQZkv8Vq8vWFQJl9jd3RxXCsXj7TX4rUA72
Zy2jFXtO/gayikGUnGvxO+lbzUxuK2/sAn7hd9Qs1Af6OdrfIIoyJs5KSU1pixSzn1+fKhmo36J4
31NVa7gwVwIee4cU8ulZ9Lr5DEpLPRsvhYf/0zK3cwTeYv80fdVKewRJoe6BG4k1KkVRqygKr7lc
yD+HA1fntxgsUZTMJVglAF4GfbgwgDTDRBz7G82xKV+6w8bsKjmHX1qNZcVSJyJPgg/2NtU/KINB
86IWcBqaKQCnzRh58prDi6jfpxJ1WYlxLSU+HN/4pBOOiP3dq5bptvZ9j/aa22xku1+Ad9n697tz
Qfj7MW8psO4lzfl/gcBi8J5RuK1NTMelt2p1kkSGQzFnGXDmGKIBr+II/jgKDnSnY72ckDg3Bfur
R4t56AwcuYz1dOq3Xw5Za6JytXzrCkdShxsiUJUlw8hcRP/HopoSGpzkVLBS17NjlE2/3/S6KMk8
JunMgUREn7VS+6uNUlYFMvjgjWM7ZuvDJVKrY4FR8/QKkyms+fmyN0T6ujbbDX4sIr/5IIqmo3GO
wXg5TRxKDQh2zeJdrRFQJdX0t6kGlgV+TT16DC7nib3ZSnmxZ/z9ab56ohV0Jtm/NK03+4K04mNb
AYWYtH2hfjoiGLKRfQhcLZdMDbiIrK4PJmAHr7fAaoPjD5YDl3Nm6iIkZbO+1o+hGbkyW6PilAlM
T+WxITe5x+zvt3T7GGPI82LKJjUpKCmlq3dSFD8ZBoOvilvtaGRO2gKWdwe64RRjzyeR6TW89ZWS
kSEt+7VQTSH9ywVtXGIfJ7rLYNq4nsJATRR+6xpT69USeQsLKvTDktCmv2wZZ05LnlSpUKk+E4g+
6pZ/UH/2Eulhhl8goZ0YiRJmzFTxNihIUBtvkNWUJitKxgY7gKRpezHymLp3DSlkVZ3BvVsK5k6v
jnd2bvwhjdYCBd0EiFg494uPsrj14iCE0nAJxG6pB9Wr9XFwqgNNTzihpRvzjEnJ8KxgMR8fGEUw
1iW9JKXGEx5UlEvdcX+gtOgbMpdKko2GseDBEdoS/eUMOY9ZWkNc2zVwGBvfUxC6dLSl9TSbLtxK
4rFP0a+biTl7t4zLwmgb/l4OmQZAPRRv9Jvj6wvlMgDsAwPDL2UZoXYo3KzaGLAPA1QXz/jY3pnk
q76XPUyxiBljEEvLKAZAK4ZZnHa1s5400zAeahoX1OOVQBxX6A6iVbN7exvInWVv/GVf72cLN00g
Ao2ab3wWEgWk5u1+U06UyUY1sshWYdTPpJiZGrx8qIUD3YLrqiAu1gX1EbkFpySjAeWwejiej93k
NN12hJk2d/uo3ljQGYzgLZVr4YCgG2a30eh/9QRAHiQeiBJzjCQYTZrz3xo3M/GOJC+LL/ubFUDI
zV9kW+a1CRRTY2yoN1P5PcE0CO5+wtk6cytxosaKyXPiwVYoRrwidVPI+9K50Djh+D4vUSySpQhg
/BecOh/nUM0bGyqjtK9ZxUd03Cuc62o/DsdrpA27xD7PGW5VSHalXb2a84d4CfEs8rRFdEuKU3Rh
jMLrsmZ5XgETHxSnPeHvvQbLEhx4+IeKZrAT+D3IRjGxqcszHuLysQqCD89Qh6zkSNXo0BmG5duR
kytuDCHprhuZ7zU0Wr4o9Qdlfx7BE2LRl+kzYB5tHGcqZETJdQ5oIXqUeHRxjfCr3O//WrPpGVDP
u0yarpgnjFQtH6hFGwTXS0LWiY2hPYXFI4xcv8aBf7SBkK5K32BR/6/3qIKC2dxnDs3yRYBYiD5S
qNs54DHbsZdVq21UzJM3FyViahGHYR4n34PQF+sjJhZeJiyam49nV/CZWeWUz2LZMWr34hZmz/lS
ZudW/uhDKWoXlNtzxDzqA5xVqB7mKFBQC0px2UG2dowAwGOu6LrCKZm3bARJLzNNEbPNN8cE3gfj
x3zkbKR1MWQ5IAIUcQj4QqJjbA9cAgi6LpmPWQCSpxA2I/L0Cnd4lKD2i347Dq531KtlstIx1Cyj
jaGBdY8X2svCyS+HYP07wQEolBoWgkqlhw0FGx0tkGJ8bCvydjG3kIhTPCn5NWjq0liEI0QqK5oc
b45hMHwBCYC0aNNA2jN1+oS9Q+7w3tjUYZ2KNbN45EQdxKxBEwP5v8x4rqmHoHDM5psOeHo5TbZk
x5vnGr5liygQhrsDU6WyUeSkEle3l91w6ni8XXYOG56h/7yQsH4WX1xJ9OdSDGbk3XLE+j+chWMj
mxk+0pak1xNqPI9leTsxadVFW9wbv6rPFZJzdNOJy31CHe5Htqdo4YJrmk+sc+Jr+IO/4CwfdaMt
xbPvFUV8Ip39MhPNCksKcME13vvu88vAgrsf/p+IphfWpA+Om0TN94QgDQc0iGsqQZVNJG+jJgKU
L9/ZPa9a41hR/tt9zgclYd1/aOqw4PSHrfDOU/g3tl4BQOo/exv4bYzvywGM4MH/yedkKSVecnMs
ituO4gm0CIo41s1ExMrEYyKkaOxo0Zctrclsrdv799QMqA0vabBnu09WG+194Xu37SdBiGxcBPRT
+3LMlX4VFPu9c1ajOUngNls5pzQC2HpArHGY4uKoxFzxUF6bcGQZ0TCky5Jh4f22Rct+PR5cs2hl
s3zknP9ReGyErY2sXxBxGVFa68B78DST2/s3F6YXVEaFj+5K0zN49oqHsr8WxDreWR960rpuSlMP
/xyO0MQDG2mnwMBEU3xFoy1VwV4NB/RtVPPb1axfEHALWZbCXOzLVLV82DqAusc04qofMvAtNBoM
j0xEzHYtLozQOJskwfKQZTxVxXxlhRWVLDxXSzQqMhuLc3v0KH8IOptKT8292UWaCZdFk1d7MZiC
2hpbmfO5EcZn8rReCGKEPLEuKvtfWQvmiA+FdvGZ5nNhCcHrF50sGS3MXlHoinWJX1St3gAbSwcy
adLfA+DrXITaflhKM/SPUE7PK85x2ODToMPB1rMk6PqW+Y/GOcUSePxzQdGAyjMyXWimMfJt1Kzp
jRzLxx18KeI+4Ommo4V/V047vbWBECLTPYIy1UbfiLWszmpfH6fH7Dt+xu+ChDkKz8Kyhp9+qG6n
/3MIvR6VyAuuu1fuC7zER0rQd+RsWmk0xypcE8rH9dHoNVxwR5QUyb7G49LyuMyeFeiAKs16cDMN
TDRzPtHYwWyLAbxFiR3b4IyrLUVv7dn/7h8+gqzjO/B40Ravk5aZjLvGSuUwgUgBP6NWUL8HC48k
HTfmey6YSjdPPmxFbPnAGL+IYroLbpYczoFjQjsfDg3M+YpWPHc6CjQIoxGRfebHJ6gxKqsXGpn3
1SGMX9sPDxoQfcgMu64GE0XOwgBdulp27x2CyYRYuIDp2T1Im8ETOPyWZJ+aaESg7ET/T5Rrb8pN
vdClyBVB9VM5fKjQKn69KVNX15aw1sYGIvnl5dQxeR8JBfzHs6vmHbM0n/9FOmYPSvnJC9h+qBU+
Kcw/2RTkbIrisDlojI+3Xh23ORuCaFSJDxeqZ0VWyq11Q0TIi24ZMphgXjP7vnm/UiT7TSvSleWY
wesW+uWQ3vEm8ZFXVbjzL8ugGl3nqHyBL+clGuGwpOwYgEgA7+HbWcme79XCmZWXVdIjr886hSfP
KbDt3OY52Vm5BLe5jzp2dRMDS8tENiXs8P+9DUhQEKdG+c5z8wfTL6sLEalO4fzyH06f7mFuIc74
a07Zos95e2h96zm7mejkyW4zBGyyFB3QxljU+5BAW+rh59+MNpsEWqLB3GRroVhrjVxt9IGbgt2q
qv6Ulc0nIGfZGaVfXMwLPQ5hkRUxUeDbQEG/ZwU6V4bVvvFWR2dfTCb21phoPvacRBhQVXQOC+8i
Gt/Wtf9IvxTX5VOakUQaiCPCvu2e+Ve1OyrMCZao1qHOdZsIg4/MfHHU6qS+yn5zvuFJ0S7nU+1X
le3BgJNqzA+KU35XH7LoDuviaMaY81xrvLTwlewpBO7Rji1ZblDVztS6XYkZFbZqc+1Rk/qBuAMq
nOjvoStZlXku3tNeX27xbxPw/Xo18j2PZrNrEKj33JMez8i+BpKbnYpC3wym5IiUMxKqr8MNovNe
yb75FEQ4BfarQq2hklDiGC+aYa3YIsVOylkkr63IX7NG75J60yyt1LXxG3FiSRb45TsfVW3ioPJK
R7Ye69jUgCSjr/6kSvv64US8Vwr1kfH9yYe3QUTiOSzM30amPavzXrVCSjAY/5zl9RtGnS1c9Kc4
LMH5/Tv0BSLkYY1COPdCf0ssVWqi8iqLC6NfVcUK/k4KU+0X1kYOPqT1KIQgankWP7LFmHEfM1aQ
ZeLHkXvTu9u5swiFgfXsUyhOTYfOM7C79zzrm73y4nIz2M0zdmhnh3cnXgpQEQ3CYNI3ykz4H49z
O4btIJfzF2YSSngP2Y5Tn+qeZa6UybJkEmvCzD16Qkk/P8hqlQU5V/IJr7A/VhTrFEXkY1YBbTTX
/0uryrslZDFC8FLKaE2L5KhGaOhRmefpMM91o5i+tcvTKNS0erYlkSdhD1JNV+GMR5wyua1U1ruO
k/REGdd0iUIfLTtMlGCbQjhHHr6eQPnvktHuV53Wsg6W0g1F6VlfO5qDRowmq4bQHU4xDzWlniTm
8SBpiZ4Cc1Uy28RERTliPOSWF3YeWsN7ZOkpTgo7F5VKGnIknJT+Msb9l/vWiczx4SMz+3T1cVW5
aP9xVHYW2KdZ9i3HPEul48jGZxJWdE3Ayf5hLOUB5gBZ8nPeS/URZPZ1G6wUybjtcfm0N7ct7FwB
EqJwjQHryVJK7dNLdHMmE28KquEPLnzm+8unI+3AMwLQASBOA5ZFStUCigwsk+9nT4G42zbeKBME
pMbpnJnBOlA3WV/0/tT9ks5ylpFlfXKLIv8tRLEqvjWxbiHAoLhGWt9vBrhyGbOEETlyMngabCcx
DxX9IHjEZDVG2lno5kC0g/Z9lGl0ipJ/xbRc5Va4UkqHdVd5baI9wkwHbG1qig8mJs8bDp4KA9kd
IrYjj+DaQJGpBLP4LQnWbQn5aszfK+roMRl/UE1Yy0SEHv1aNC5k5chOiKhPbq4fdiv9xtt4QlhS
G4w79uQd8SbcUcwarBk7/aI20N5nFbacIZRwF+oJwSWYm6euBzTf12ZOKIS8UENQ28K8c68INEHW
U0ZdRuBdVy/Wx0KxKvx3AX2K5eus8vyjRv5BwRNGgHAGJ6u1P0jWn0sN34SJOZNHsE88lthrcGkt
xayvw26qDQNJvu6IgupXwkxB0re9WyREmZYt12KD1f7UdWCq+b6+s/tuvak9hmF4HMwPmXLy9G79
g1SSgnCaU//5eReSgz08MK0LXwNJa8InN3swjGM9f0DTNYs7D04p3LghebmIkDbYRx+Ca0w7fr+m
6TwfdLsXiJJSSa67tCxvkte5y37oiu84Cwb+NsDdazLP26GOm8WxFIeR4HMCNrWdNVAOnyNFSOBj
GNwYtPbjZwTGrosINKqP0FiIlQz3ncjg7m0b2F5yPrrQ4grzf3lyYcOaiFgPIsppqVQtFiZpSnjB
7iPDvcJtvlD4sedg3TC0UTd38ujDdwup2f2pBSjvwLf7a5xvcql4OuicubqO23o6eYJY+dJwVbha
xKTfdXIa/iWd+zKlrL2MT3EYA+2ztdLHW6iF9sjpbn2T5OWROlGj13MMdO5cK3zWuYqL9U6peky0
3ivarXT1qNxX5yheTS1Asn9Ee4mUvAzfv9ZBCutz0tnTBU9KZ5tpw5OH6gBeqd+B+Cwsy7ScatCJ
/1CP44py8aKHM1etViTMIAsO48zQfnwcY6FzEmpPeIaCA32FGsE/zJo23L6+TgVUJYu0Cz9HDKgd
mwDqrOeICE2RMofmUTJap+B/vzwFPj1qe0GH/jye82vPruEhdsnFDIaakNBg6+BGnLxIGLE2Kzig
gOnGH1DPJsHRhOGQV3R5kqUdCQvCPL9WS8VBV/mWtenRWoFzj9indgut5wot0NYnGqYJJu7/eaik
xZ0PG515u1ROAShUPiOww5bof1QaYTAkNju91R9AY0gvGXD0c4RHLJGZ5gbQENhA5cPwxfeXnlLM
c0Ey7kn/7n6IfRVJLPirou4N9S9hh70JtEM2uiQeT9jHy5Y+KgGj8QGMiimyOwJhclU4bHKPtu5C
xG1KCNJFGF3JzNYhrEXEiN3OAzQcjfIl1AYeKsAXKAUgkn0gY8GpmCbBuNWfvbkYjdspnUEMLH8e
MH2wCzG8yPVdz47IrJwDL+2EuwXql3twipXXHJfiynwY7y0pYj5CmlgnzdV7gHArz+Ga+0ek6gBt
g/K3ncglwwVk2PWxBaOpWqy56qHH2A0xSW4vlfkYKJW1ERd9GTpfYBteYJbyGAEgMBpwUDrxGLuB
HXkmcYM3cvt0haFsQfBxto43BlLyGGdxpT/M4lEp84Flps7crRozUc/EdCexTP9/WKXoLmpehgP2
q6FfDDHtvnysZq29Cx+l369NFsji0b0zA0i7Wjfl26LQBtihZ9mWl0MhzUfsNMEPkmnCWKb+s/ru
2+w3RUo6GgfriL/xHRep/p2EZf/VsBjf5oSbLgjLP5Ffz0L8wteqyiE/PahgrlSDV9JVcl4qRh3J
fnJ7n6ktWPWq41x3G1b9xGEDFmbTMogRbFvcA43Iw2ofoNZdx0As650FOqdQk/8oXA1I0/vzssgj
aaGqTP1h3GeIu44W6loMGWdmM7TkhQ7b2+zv+87F7gUD9p8mi4ROdYMTJ+FddJKL5Svf/Wqdpw5i
WYMPZsPx1dorpbKvqOzH7kDPBK0CrXyLejJBSvi+3KNchdSyMGWHoX9T8HxPwp+OT9MPhwHVpBrn
S0wJ2wGETW03/8pIxwEHlo5bBDsi+8b6sIVDaGkoa/7T1PG2yrXCGuKn7v2uQ7BJHoI89KsulH/J
8j3gVNBrTkNqWoi4YPg8/uVVmyO7U29OpkTw2pPKr+0PNFtSGcHzdo4J34lpA606ytEkUHwwauMh
oTNosBWujcZjN9gES1OhR4MGCSL+Qr7BVgOuQcHDOxFt1Lz9PW7r6I0MJvjMWK2EJ/wb1MWDp0pt
GUAkDsuuUufCxkuoPcHi7PKYvQlmt0pUG6pbk1nhWyma7hHkCET1Uz40pO13dDX5F+jDjUtF/Auj
sankQRPPP5n/DdjxmLKAS6kcHPNXN9wDI8k5Xbe+aHTf774pPJRMqMBeeQXxame7hnHGJmTFROkP
7mGa1WEtAhnfcC0KCbvoU491u/VCe650J5m0DSgEAooc/JjdEdLa2qYSyjiN2tN8cNPLIMFdy40h
lU5qhYKRQUFDr/ikRL3bFCfeHu+8QxteUQ8PYD+OT3uaB5WDVWbTIhjyD4UJC7GeDat8Mh5jAHga
GRyGz91u0v7a+9mLCCBenYNaxHFB4xaanTZ+IYm/LDl4LErnmLp2lq1jAfJgsHYcETrA6WvcFyw4
GopfgubDGzpjMHDjc15Oq0VmcVX5Oz9U/QQk2tlEyLitFZOhEcn3RrPmk4fX4rgEQQZYpQx3Os1h
ICRXoLUL+FogsMOinohFRN7IUKrRRMDJ0UwakF5rxopE2ZIwpKTUeOuaKNUvSZ4b0sTfniYDzyg3
lC4NEVwPDNLhcwFsn4kNqKVPbu0SV4sBTHv4IrSmd6uzJZfvLdyHEpK3CvYTiL2vHGcWFKeFLlER
elMHPL5lPJvBTcTMqpYtKNnI3SB2Fh1wCJ/wYCCbNP0myz+gFlNea40DromFDkyQG0xZ1zPYCYbJ
ZsGRnEr2wKV4OFYgd1o1Hjf/npCQOPeEKaMBx0j1oGxTFwURJ+17dp45CWyVzcopZlxKxJPJ96sC
SQ+HccUOSl9DAGS8X5h+lHEjbe8OvVCln3tc6YbGpDGdYZ2LpzHn+QF5dJVtWHaOHRq9AQTitrIt
o72mqbRDVaydJdNe1poKdBvM9XprUzhsFXANz7toDeeCzJnlKmnmdYZb236CIFKN7c9SxAqU0rqD
MhifXiOzJx+42eqiVE9ALYQDn3GQjtO2POYxoaofuGgTQaN2v1Q12kICcgNnHF/G6CMAifqmG7vw
vUR8HG0QW+ECbk3kfyj9UYVRnBcRGAko9G9w9+Yqk+A/sPwz+F0bFTOi/n0s31WPm/hzYRPvQDly
r06x9it18kGZrIy18KJTR5UKuBubRnvKOO1d10xn2J/CzBcAWhDoY+anvhTLcpyETIwyMIk4WDjh
opAP/NQ5cCpnNFKpSTQOxu1krGuNVpVGaVdzfe8lNrIfx1KGN38bLX4b3lHB9goVtoQCW6VMQk7t
h8CynkryRo9Dxza2EJ9zaFt3dDGKd5LOKyOu+DTnaPLZfgOrgy2gsRV7+vHwewku3oNbNaIhbVmO
wTs1jjY4iSnGU8jlXgRywjks0EMvVPRYptFatXy/FKGEgPvZ+TWqmyOGypFaAvzEuwf+qKz1/f9L
+pSXcSo+sgmHBlPzGKpwRXgRGvVco5iWZzs/k8gzXmWRVtpyqTMPurjPp+/+nGkYRvQbq4Gq9Ef6
b35a3V4KfZByTL7WsQnB+QpMAoI1HYP9XFnmAx5qGA/gB9Y/GLIhbqjN3aWbGE8WgTPbxHSHj5Rl
GWHhx4D0Q4VzknmfQX9+7mRwrBb9SqjZ2SvQ5+7SHQVdS5se6fU1RjifC63m3wWQPpZ4DyI7ZAMx
iNms8cvv7CD2tCsjGrLaCZf5fJA28fnSPQOnUGtdL/yDWqxhYRPyWBe9+P9uVSt9IYwn1YGgwQA9
RdWrUUWvUWFjgD87kNTfwIyP28W3PKh+RsEHq30qlNCdJgTIbAOCajsdH1KOyHG41kL3R3OxUGbE
ArcNxMYzwIh9Ge1hiCtFQmBWc17Ko6VbitVmuVAiexU00hT8E2ImT/P9XaCzNHabsZ1q21Ldt8U8
R84pDdmWOInX9EtaSesa2gBRpkPI29EDVA4EQyvQPpgTGGx6BSrbl862zGjz9O1lVMXwossJp2TO
Czl4D49qdCW1Xtv91I3UczgkzKAkIkITUSQvx/gtJ/mRDHlidu0sEQYviK+CGFAPVLquJbEt9Uc4
JkndbRB8tXMu6IVG73PvR4B5R5YHwm5Gkfz/2/R9YC5RnfliAkFNOjv02TaQOUv+m1vdsv3IL7Du
4rHMWNAEZA1WqEhLv1NIOzMu6D0XXJRZ6b9DuRlglHKntL0DYm6GFialcfW3kqC8N9u7XsGecbRj
MfUz44NUeFHcDApY6aGT74oEBD5Vlj+l47wPnpLvwp2edSpg7d5PflmU3c/WkOk8Wb9pWCypt0ZW
X0rsXZL4nmVb6iXOwZnI7TIzi6OC+Xco8w7Sjrha0piYGmxlWTrsmz2bD5UFG6Fu78to9TWzYiaS
yPQKDQa3FPnowPQLl9bNBDiLHN3JZKSXXacbe/IAtfzDGFxtw5uf+qN58IiehEn19Pw/vnq01mEM
q5SwDpa0QsqvO5+HVFFLJUAGo2kkLyaBsrSJcukwDsr4fmP1BGztYyBZkJaLZ1RAqYzYDTgIEvNM
SuCj1MkKoMGuGAmT+7AcvFtv38gUhc+EnAix6a3Uh//cH2ytQxh5+Gfj8WzCfXXbZxSQC319g5b6
UBTFg0Bl/RmGcUlr/N4aEFWYU9UBpuqpSolU4qtzBYSdgsBr5d8RZJeQ08yR24EMYXr3SG7M064d
2z3Ivr8GZZM6k0wpXIQZIPbOedueUXGhNNMYT6HTtEfX8cucseONfUIZY4aXI0khdoVLNiO6UObU
FM5xYKTcrmlhkK8S0rhch5c64c32ULc95qeDdSaOP3F1lKv41gEQpJzM+xN6McTEv3pJuQIGM7N+
wgw9y8b5shSpBBiHG+bqpa+th3BLBGmd1in2VkIZrAk2r2Bw7r9L4YUxzSAXyn8LZZgtYAo/Xl4B
KtyE6pFhhJvwowrfavjXUvp7mbRuktjkwStSYQ/1KzEj63wLecI1BFmNbFUpNYzl74euVzZWNw+F
JteQO+LDvPnK1bH0mf/Wv+ClH5+vcEblhQix0n2Qkrwz4ZhZVX+N3MbHKhRXU1I7qw5Pp4KNbpMe
2I7ECyxb8HXFKKYYVJT1Ev1srezUmIJKotu5JOmU+wBcAgkWhdqHjfYHbLN0CjVIU0hC/uBoM85I
C/afonsXhKz5eu8dy5fQwrZgI/m+x1rU90+in3r54H+oPtLqzbwnhyhESYKhcSpQkfQvelueMZ3P
AJ1JTBAN9wwvL249dNxCuU3TKzXxvulhFTyQNJzR5ZLgyiBHvZbSRdvedVQ2+K1MohOQ3922IfAA
MozWbqssRF3kFOgOHmKaR+zvc7OI+xLTy4SfWEk/dW47SYHLw8UQzkHmh0buEaixkmffVhxV46jw
Ap/t1sBws/Z0lXgHr0QBjAESQbVOLOPQGwrGrgJuE08SbiOOZLBDMo90EejZMqIbt4/svi1gqQLf
JzvQMUko8DmKue5TwCB3Q7zFThGaiUcgpzC7s0ia8OPekq9IH18Hj0usxgrXzqmlOways6ihTjyz
NPrriTEPPUglTuRbUe7Dx/4PeQ3G9fyvjRbrke66yfCUxn/sfthtPm7REd8Q17vYrhswmpADAkRu
cAgDwln/kpeBvT2L4okcLkrEFyHsVmMLvXdW0zL8VzoHuoHM4h9ZblYh85wGr8kMjyMabu7R1WLw
DxVnVLfl6KEx8rCO4pV050OLWPnSrsPrNTMuPeBULrpC8NURpTxRWIxQ3fbc4inorLbminiznLSB
RtsVpp8tgaRbdwx17kQV60ITs6cMxfGz/O1k3aHvCb8ur0Zq2XEV4WZM9tsoTnTU+TYWvJbAlp2l
GxtxdxYAcKI6md4M7PoufpWjwGRgUmw9ErCOC11YRBp8HbJDdNFly1F8kRcUpIlSnOUDqsg2xCZz
nZ+XRT5mcyIZB1LYdOIKYdVVnPFBR2AGQISTNqV7ZQZ8Ip6Da2m/Jl7QFOcdXNIk0a5fS6/yQ72h
d09iVAUVHoZ5XlHrh64RnZIP68MmNuGHpThwNgsugCXdBQSfto4lDjSpMZx/EUgNKK/JIEiPIlmX
jB3+xv7eg8OdFA4ukQT9zTWedDpFpH4jFiHVM/Nele/vP72V26tTN+dgtzK4Ju3f0pASVd/kezmv
eIAiheljEYA2Is1p0979DOQ7oujkfHAPzR2Ht2ZFiwJVmrMjziX++UquxbDH7xvBOevu7hE1MceR
BVwJiabjBDcqfpbE75rWdLG8oodYW8SQs3JLkEALusgS4NqufV+2GYBksyiycnzPSI8wawLaIcId
4f7JX9NmUjuS3ewFMkLWhPW/Cn65JawoeI925fS+Jk89T7JegXzRtCV+KVYOFe2o1UNzFLiihZxY
nklaW8jL6jRzzKygA6c6VL60qwJqDSrc7mCWhiohPbdpVkQu60aMXppzFYoSxXkXvz79sTVJ8r6H
mTPzeyUqkLznhG3N9Jf3RmEkk3NwrHtGOJqDTfiw1pIpXIsks9YeqOBNggR35l12jG36uMAoVOao
hQNKZhHuep+7OhVdTMZY0leW5ZPHwSO3arGXKJ2f3HGXN6BJxjnxqM+H3KWy95u4QJnTuSzeH/0L
bUo0nFuTO+p4R7t81C7IAYHx6d9zdKCytvBYip6w4y7LdWKTClt7IrudvsaNS8Sz7Krd6HNJoQKz
VfHNAnoFo66+OucSxsHdB3GFuarhMmdCyukVP+iF4aD6LOV9rwXTXtxwZyow7fw54zDxcGSvR1sY
qjZ+Ccvk/YuAKSFjotH46DeqjdwG4P8jiK/f2dWkyABQyFSq5/ZaYXUmX7jJQ6ysqEna3bbjpH20
lyP+G8kyATsG7+CvkX5g0nkdx6vSEG3dl/gu8dEP2ySEbHJeDKTis4DYlmXGb0ShCO9F6QN1wkWW
jaPhKmxCbnEIac4sCVFtG0etimCAWptUvKMF6TQD+AW0t2+MRsaboG7VJVZYTxcNlHac38zP84IK
GlcQjCg7uG0krRfRK6+R/aNljwfqc4Ufdl/mTtFYtUv0y+8RO1XmHSUiXAsOZwR+DEkvycVkkR5q
QlsGm3tNWUB9vEi5W3OXGK0Ux8c8tQmjIq+TinaWVM5K74WAEFeH8ez+YrHBFmcEzTWjuLUUf4e5
Ew3vA8cLyvDO09KWQQtWuTTtGjGHOP/HmkzHbwV//aqfGkAhZVv2s7z3yH6xl0m4hBn+F85qFtWM
sgZj/ic9/U0yqo6yl1oaizeRPdoda8Dw5Eh/51/xipaKpLII65Va2XS4ovYZK1S5+0tFK/ZuMdcm
KwhOUhNg1V684C6YYnMOW8AZalRI7lwLINMkPC2TUk7ontwT75PUBa1EYn2blg+9d44TExtbKVbL
7GlmVrveQgOx30Ah9HOiLJfRyYO+HDOoNXLZbiJOqZjYxBdhD/tQBkW/SOVI5X16cbx9mJbg7OpY
Bt8lvyiFOu9ihn/JzmV7KamIaHvW2XRXXfdQ/bi/en4c7emQLLAMnlOa/qcj9pHDY2+sOBqxX4AZ
f39z61GJIdheRQvSN5H6cztXOuvey3E/vHhTctZmItriNsXXYc/jJ2GHDQxPaWCzN1sQWtTS4rkQ
gksVfA324/3NM85g74JaB5K+7TO3dEu032l4CSi2FoJtluCRfOnW7gZH8yoRQ/NYgeYlGlh6xKfE
JYsZUQA5j12u5Q4nZD49ELBWFBJM98E95K65+RNBLlTaKzy1Dpl8xLTN66BK4OsN+7NKzn5loUPy
kzOpPxwHf94utaF2fdf6NLh1QIPXP6/EbbUVWuBG79HlO2PynuDoCaZZwgh7Ylq6XFQtb9cZQaK4
1LliabOknamXVr3AsmUJGyLcklBAq+wYAPKWn4xsEuxMuJOG/u30w1tv9sKE/sDD9onJ7tnLXwpk
8SPzhbpNXj468EAQKjBar9iqUh/RX08QYkO+twtjOHhRlR1XCKHcq7cUyngve7R48Mhl+o0hgn9p
KJWE4UpYMO+85caLwoynJCJPIKTjAYbyRCPnghTPTE1AQpT51b+YKv04M7eqtV8Wkonq+68IV67M
3j9dsIB/ecXA+pSpCP2EjdfGvKGI9gAcRg4cAxx9Pcmrpi+eQZHaHF5fGHxxCM42UA60l7VeZNS3
rI+kJ3k/OPAKZvgGnFbyeUiPgRsTYyjl0jLsUfgUPLt4CedumhA2p4MQyWQvOr609Ay1KcVxGj7P
gbRywh5KA03z3X7+Oz8BCjTHVlsw/EiHDizZDHpNLr5peuQNE8rhne9X9tMOunJXFoRn/UFQhbDT
UT/Qj5hbsjPbCzXJAnWu3mOK80Fsbk9wWiGQQyJHll5mBW8WBiaPZI54WGiXxtA9xCYQTd3oKHqi
EJVCR37F/BWdXEfgqKUHavG2SPNXO9q/xu7pflqEhh0BvKWKA6cHPFyKI0nM8SfQILp8+LPPLptY
Y2g2lhgy+wR0sxGSf/eTDkpv3Oi4zpkJT8F6atlbwauEebRTMYomt1OTdPqSQCoOc9GZqNqZPKA9
idNidrMi90QpXNLUnJMQXbj2LFYbEukgCSgaVzUlI4ZTQafAq/6gdQp0v2vGjc4d8t1xoxGtkuS0
wCAyOCEwCzgBN9hRzEd+fKggxnVLiU3U5Qatp1zNpl9FK+Ui1wFRN3vQ7kShaeZoDvfOdcu4cnS4
uqv8mpmtlIo81WQcZ1CF758dg287k5TfC4qA0DJcLJ7inTsXLXwkQj3fOJGpssbapmJEKp0QLGH2
at3T+TFHERQxY82h4vVqWFdJh+B1Gg7L8eI15IhdbSbGEGRpA/fVA4hzF+GN2yasxPJYjrz0jrsk
6WyG8UPBPlBuhpHFs/dpKOEqSMJYOdpb1/0L7cIIoeD0hYw9lAWp4idM0zZJcr1d8FEkAiEhOJxr
ptfCmYE4o7f+cSit34o/uBC+xO3L670or2U5eauawcE/6g3HP6grjIn9TfllNRoNG+B8ATgpYEiR
S0Bvmh2lZW0IoV+dG5adZtJqdDgU35bhHBrAA+9eZb9gVMVdoyw8YgqUPq3KATA052LAxWKo1C/X
G3mX59EpS+1faGfT0XTYstMUs4CdXu+5+CRs9rlo5a4iLTU7aYX9eD1D81t277MGLSmMuwIcjU3+
DQxGTOTVAL0GqXPAHGPK9zY7OzE6hDkSiXhQs5DdHTgKfqceHdDR9+eIJoDkRF6eyBLSaWa9J4OG
BI9dZo90O/7yljOpL03qEEORq2sGGW+DDuLVQdB3WtMcM66/po54k+NygNjN7X8w5tXXNh10Ea1F
WuyeEo07XT7XWo/Q9GAi1dZx2z1ZaIIDfSuaRZFZVlVl3preSe1gtFGwhQ/g7qLFyE/B7ON7M8g1
Gf1eS0K5wgP8KR8mVj7tUghUa9N1p0zeTXtRIborvEcwSLInaP0oMS1ycGrlDJoUHrYhJ8SAwW88
CVMkBtugwd6HyzfztsdJ92TxdWiU4YrwLquT+VZ5aD1odpDr8DguFB4pDaBeBKVbsNjZFVqXzP4P
CPnCMYCeupOY9NIJEQ8oHq7RNFmoMy+jNXTQsKd0vfwhGLkwjpMYDiB1oHf2lc4WCHUCtyv7i1CW
sNE4RKD5W3YSbT7MCdV5ioN3YO/86XcNgsSBAc8rFhfg/aahVp7D2i51P2qFZ8gmxog5oc4ihWKU
e7OlPF7CjB7RVxASxLIEfteSHmuWr7oMYFxVEXEmzRQ7ETNjrIj8I8d3ROky86kkWwkzK1QKDHrc
oGbsgIfogRzyH8kZ7lT89bv2K+4X6DdXDOQ3sEhACKQ7Y7EVao9LC2aLn6/85O1sCI4EGy835+mx
N6lZAcI/uhbvTHwxM+076nY8B0vRD1gYlL5t58662fl8R+MQDVUCQ4jlkQEcVJJTwGVN5zC36eeK
2UToTDXy8B43hsN1uk1MFXxM/oNpEcQz4mkt7D1R5B9v91B3jnRttI3hf61CPCNwIz/pikruHh97
/vyj/apXa9u+HxtHkwoQm+/SXItUgPIGjptAM3e8KOCn066Z8Vno81c0R9ErF7YhRQGVH65ndDHv
8inmW4HXE4KBy18Y//hmiewYJjEo347XQwClSCUUpswEoUHw6Oi+80l+oc2xED0/7osMon/qKa8K
ZMpkbLyPOMq76Rrned9zs7KVgNZ2VSxdEbijegb8uPCtHufWgKfoYQHfaxM8HvaTW0FcwDXjiF1J
TYNT24rV8f6qPEOIpb2FcuSZWZiGIS0/Y9a1EndBFZJsgEgbLa02h9Znlpyh2eyRsuwJq/+aDTv1
BzG8CR9U3l83OHjMkBw6Hdnsf02Y7qCJ7h5/WF0e5Zz6Kp0Kq/w3/bv5aSekCPLnpvDfH+vp0EOI
hJOSDoCeHWaZBJbneqptx3OgAaOH3XuFxWbBKqntkMH6Ep590WdGvHb8xU/cARzZfcKe/cz5AUcy
m9/DjdLieJGvPHupg679639rg81UaNq9YARNOLfnT9lH2hmQHwRmBoBPsfPY2n9B7/tNQmvKR5Vj
CITy1+1ucrQK4mSy/HLcTihqEetY2u6bMwVcrtuzJqJG9S2n4NukurdFFpQdJTVdA4ZeCA9jCNWK
aUNg7W2YohYgv4oLbXaYy/QAyvqFi71f7vyNE/0NrSwG9VxhDpVGqmQQSRezfyDh+ENvS33b3z0W
gfdtyPA5qVujZlJZwpgKD6sQXWAPP7YxDtRbXzgO7qQthaHeN4K8t2N/xsB2SPMyGZvE+PRwr8ff
Oog1o+MKkmIJxxBiOsydctmPQoeNC1Li6A3dhJT+K/7jenqVGFeZV8veF7BgLH91rBoeU8bnWBu+
GbphLVurVAsnNrWnWLTOiKYI057emc5qs8pm73GCSvo691UMXcffvSLiFJDpS/sTdVljgSOQlMlG
tWFTyI5Y534MiCa+Ae+Jpu/X+Yir0DRw7EGMa5lwC2vqhef50YLvR8v5WLfnKLFr6PhNRPySm9V9
8A5zzUCorxqMA7o5cS9GR2favwnnupY7XE4eq2S2ZSYI4IuZ7j4eV0ohxfjuSy7cad94amNmBZHN
wWodpfrodIrjrbpzTObRJnJrKQvmZUy98KCvvtqGeCXLIq/ylziZiXqppVJjgg2Vh52UADT2qD1p
TmvD1yPwUVbPMezhQmUi8xb+RAxhXba4jWh8jWxFk0sjEFhonE5jK9RM5FkO9jV9S6/8+0/NvFxh
Cv0VN1egE/uLTcmwc78LXOzR3v4gX+HGWyJQmuAkbq62fAOQkDS4aujpCKkjt3+hRpqUFrIO1PAV
hOUgYGGvBECMlzRIH5Ih7J4M2KvqxQS/DdYemtIg3TqknMBXOH9do+V8YlHOzTvFKMjqD3rzsGMj
rGI8ZM5Us0EXKkT8BSE1sIB8Vn9emXoUY4b0G5fNYLQUFQof+j5TWdzY2cVwN/7ljwj/Q9T4jOsn
79QIHFz1JbQniZSk+d+JXLQm8aGCwETtQhW27W6/bxEAhsBSmmumOK/oQ05BxRCrIK0qfeaA3Xt1
kCbHMpK7pjBYVukeyXkrfocPTeLZUE/JuAb4A5TYCxlk3eI3eZKbqtRdK2dRx5vxV7198EkS9TEh
VjLnF8tbNCSt40i6d78WqFQKwp2nURPUDmFe7JCMJGzVIa1Zr5Bog+Z0urvoG2IAluP1cnRVbCbw
mwmLX8a05XI+U4D2fSJdk/fgQGt37rk9gImowtjJsACJfQB6NM5Ftiq7Aaw6p739H5DN5UzPa6i/
DEW1ytn26T+J/Vpcp4SahX5ylK9T1uOiUrVZF+APtKyGWNed09QtLMNewfrZdWQCUguREjYH8JH7
T0TKOu069hko+7woYoesJXvemX5DWYr0ZmHXJzeuQob+gqlbXktJjGAR74muD+qE2SQmXo0gfik/
4nKrx14Opbb7WMfVqqctRxRKpIK0X/LdWrAnC4WM94g4NfEJ30v8hgNRDLBwrqPd/nDqRPqB0R2r
ISdIZqUVakciUfUDftjWUzQ9Pc9ST7DOt2FudmGuRvjljJ0XcSYLjbmr8bSMiIP1lD6HWjl683uf
MkDFpD/8l80zGQXD+yHNQ5CYCOQFozE5xXXkFZvUegEkyPQe5tPSi0ztmutVajjiGZNqZu/mRBBD
xqaVgNrm9YYPUGjBrT7emobu3E3KAjIFUWl4BeyWE3Tj1CIeiMMgtmOmhnejxFGGuq7KTUIdxCco
B/0cnlhMaawsY62Bva2RyTY71WN+FHqRVvULT0oI5zyAikkdFhha7gxvAnt3hVHOZopz2wsKkEz0
RIfkJEmETLRNGwDl8uTHdBKrPFNIoFKp2DR3vg/sP1CDXKEMwsj9PmfFFp2e0/l1DxIPe0JnETJO
mZ0xh8zrynw578TxfUN1UPICrcxhGUyDx7BvbYC0QS/fNmYg7b7DmGhhjtclSKFzi5YKGnXMs6mZ
5W5nAIFHCeVpV4MSAtu9LG7hIsSoSt7eL7Cx6ft22Ymn7GDWxnSbFukf2U72DXKUrsYNEk4A0bks
Q83MoLhMLWIjCoEn1pIvkm5dDoHlUWzEGdkf1ymCl5GseIDwXS9Rsfswh44Adkq32hYTp906Hf58
zuNzTMziK1D/Bbi6aR2WZEQi323vWTN27QD8zOI+Ki3ilciavZ/6FbjP+MKYq+0rR+cy4xq9W+u0
SaNax4KaRYua7PCvl7lbsNcG4rLmWeAPHSa5T5vBlgEb00fjjhoUWcj0+8GngiNDzOYjEyJdoTSo
9f3S5SvOsJAfWr/9V0j5LvR8wtuM4b5/lHQ1gXSFt2pBxVuGrpAA7yfZWVpQwPkNGnkv+MtEH1Tr
RVGVTnE60hWT8z9SZbiIGmkhdlo4d62YU57MSiTYuF7dvB8FkmiNX5qs4W2blSeNxcHeTF3BDli3
Vk9qYkhZTfdajvJBhOrxT5WLVIK9CoS+avfgLYehQwqOnQYx/hoRONxnolAsNYLBnU3jUNRklqr1
J9/v9kGkcvtUPATxdxMuK6lRUlXHEy7wc3QqhSppR56IWY/OvuUl2P3ERwmEtLjVoasaF8JsVcbR
45gviCIZ2ruceZMJjlccful+n7kyFzUoZA5xX7PZHr0r6w1tLbqgPTdafKo1jEhLgUR/3kZuwKRL
7Q1zh2Y1LY5/g1ZWsqmMeqKX47ZkOmowiIct3urFJRKlKPGP9OF4ZbP0QuLow6ReKEUoKgwH2hHW
+FYkQAI1igFPRbrySj0DxgeYpz3zT+M3vduVDzkEtU7YHlLkR5VaVdWfFjO1D2plPzFN1vs6bT5V
nEs7WTqfxkKdJefjtJsykfghKZ9ScK9fnkgMrK4VFYeUOggZx112wJ9Myn+S3lwlESaufptPQ4Go
F2zr+pthWj9yoWrL/v1vjavxRLeFHNvOxLDfmtoLwTFrnJ/ch56DE8z6c6RKPoZWab3gFDDR8IDG
FoQo0ipWJZwkqbdA0dd2wrVSv6HitZR7QMVfIx0blkM6N2XRdSbz9YV44tH8Qh22rPfv4FvpLNkU
uDBrVrkCJgXqolljrjC2LItQVEtG5qrhqiJu8o7phRrQSHxFKkqMTgPgOliNxf1Cx7a1rESblv3E
jTEKhg5/9UWOja3Qo5v6sT3NI2ftuMvPJHAUW7Y+0gpfSf0oW0H2e1EqkVCDPOSU8LWVsIVqKUF0
MqDsDEPc0C8fzA+URSA2F5es3SYwxqsPJWrLcZVcI0eQKCc60PgBetfAhrCz0o4APsTYKgHTfbSo
mO2YcoOwJrF1n5HOocKgrLcJLLZeBEOyUmI/RIOTt7tBfGaTPSk06K8OyjN04hHNqaGlRIPDXKJj
jbWgo9kso1ALPAZFgkipNfCyudfQ1lQbUVDbVL09UlEEu8ZBQgRGUfZG8V3bt1o59nvGPNc7nNG7
7Clek2DdpoCLVJZZNCbm/YxWcyACBk4JDv4+uffENQxc8wHE90XFMGofpWRup4K8bx0rz3pGYoX7
vv46kxunnk+3cCJ39h/XX/f34kFbibHjOJLLKVIzF3/b2WgnElpo1PagCWLJ1dWneKfClSnmB0aA
GUFjLwq9szJz9nLJ1fdrpiSwL6rGRDGOD7IfdZwZf8rwhWX0xOMaQRjruAiN7W6u14ddnnRPYFnR
hTeSvqjXsBYmN1hv/7j+yHhbKu5aeeixanjbL0HyLzh7jJkr3lQWzf0SOt6rzM22Vi+w3WDDAOSI
azjLegXP0zrZ7bo/NfbaW9sSVrs2Sd9Gw/7Oq3oVkiRho26jnAzfzKyASBf6pYFY7ss9qxJqDil9
CYYctYzHj7dXHnh6Ym5i3Gth2Q+5UcyWMn5g2hOzYCRH6mp3hbTPIded0tii+nX8w+KnDZR5xuJ7
uRg1MXXmh6WPexOHLRgCrr0Nb9I+rbinuKvU/paRSX8EpIuuCxmPfflwFvWloF4vexw2Hkc2cJUa
pnA7EJrR5pZlXNomHoUjsV+2kqzETUkbSOvAc748pP2XYNXBvMTkTSV1pPfmqV7fUoMdpetYyArw
2GFejCptuLhhypMn3J+ZwyfmgIy/fafTnjL6/IjAq6X1R2x3uZAHdgZrd+gd2ifj1smkMcNz4xhy
Uxos5tg/7aJBT8QTzfD9qIFWSsmnSlYxhBuBap10qNJZ+dqyYp+Wm/lsGl+H2L63c0uZ6AsJU0nF
w03aHqn/0yMrAHAuK2V5eLCtxoCdUPuUeVKDEPqGZ1tYF/NSbPlQjkgjluXl3fgBNFyOn08S9Vrv
rcMWByNrnanJhgaEu9mRJqFJUdwQ5ApyveHgkpvT1DblTb/z7pSwFOahrjNyy0oYrx9h/tYuciyh
uDuiunP/ziFgZ/K2T/zCrmyJrshc5CrML0fU2FwguHIXOjlVyoRnKa/kYVZscecOzrWrhaxBvKuu
9A9KMZE4Q+T6vKw+EB/X0uyJvIWnb9WIRZHqOGWCXDF9zo8QbEvJSQPfTvbKPQA8ohqVnl5xNshI
IHNqFFF09nQfhT8g3AMhSFcv09YO7yHSm38kK/nV//CL+A4/bEgFHf1Yq2GGesjqfFE7ApLbgC8B
uDGHXrG09+hUceXi64yGJNosJgbQ2Ia++J39KKU9CIoc4GZcz3CT04hkoD2p4YKrhyidt6NXSRWx
FvKNiGzQHjpGZ1X4tz//LrfgunS6O4uC4b3D9BCPjIMoq3lUKqnGBcoXt/sma+h+g917fxzwh2Q3
e5UtoxM+RgHMMQ1uqLeD3IV5VWLWBLFcBnCjFg5AGGX5BbRPBxQXI43qoKCGi6CiTvhI5RtTJzMR
rND0/czrtKqKp027JXodER6D4HgEQZK6jlCkfEBMw4fTpUYG15blpRvPCXyzDJ1aoYZP2MzjC2lA
FLJ+u+28BCoVhBQbkzKHB3AH4u94889/wvbem0gJJK0XRvVQdb5nT2WXkAAmnEEA/po1AAKY9msZ
3WZ5EO3l7fjJhp96snJC2e8KN0w9QNycF67YGoa3IU/nqHiCLxqMZ7FVj+kdGCMPmZD43wsTkZS7
CnesdMtfphWwWhzyTYnwVNtjLscnwxOBoU/AiBx0W5WACG8elvnudMmk8yKW/Emp5UMLRE4+bdxP
qkLRYnYVST8pwEvKMwMk7NX/ACmVH/P7stFwKGB1Ia2PzNwgG6yEpmUhIMwrgjzaWkEH6aUCtaUO
W5Me78oWJEWUz6qugro/Q84lPEN6+LF5BRBpXUixyiVgW5agkbOKxWnpfb+LvUsdQJkqbd1TvIaq
3L/fXnkpWbXyGHMPoOsVaDqzD11/TeL1DDN0TPN/PFkMFoaDD1LMdzQ0/2PymYV/oYPtVyYEghuB
ETJvKXMlBaiBTDg0DOYG88fKKapPL42VIGYbTrd1tNnArkFFmQavmXIYRQBTXUXSaGESqUEqSSWS
g+n4O2qho8ocKbbvdfpBKQLKER1Thv0k0wriVnvsuFSSdIH/bO64JDoupzCER9fIFbtQLUMUtRgE
9I2lIEuVygD2qfCk77Z0FWiq9wKqbXgnF2FYIEHawDY6KRtUjrMpIn/w/7GqSa+l6oZMuvOUlmcT
CwlvJIheMrFLveLc212UcO5jP2rzBP8bKvgLF8LPIDQYlBiJ6F1No4D2nNydEeRID3Wu44wFrWGS
6VkNA7GCVgVSuC2H0uYmqevWdVt47F2sWoKJeda2+JaiCyuLefGCH+IIj5+YEhD0MxqGsg+NuQ6L
SUQaS19vPZcvvOQB0fxymHjU8NUmCHdAHABALcV391yLZvjDB9KoJbuq4CRQC+7PMDjwYcBUbqfa
rHRkQ/+IWeoqgySsFfB7SYwO4whRhAYyIcrv0rUdyWKvan2Qc1uFAgM7SHuhE4YMCUOj2UbDRju0
etrpSpbiXCt2Nx42h70yHIJ1cn3bHXCBPCYMXDWHaHdZdy6F9LuH8d+dlTKChUHtPzFH5MQ9Obbt
bcT9NltVE8/Xzpjt8VMWEPTftIHLNepCuWpXmkw2jM01dwDsz/cwHe9Z1vxYEybCzf8zUp/IDvqF
ARiwuioiXTmCAlkW9vX39uV+yCwLviPevK8Gp0yayZcNHpiaSXStre3mOztUqRZlj0rIV1xpLOsP
XI3i8L44vNILzg+K2JCxKDvxgLpV2mEjk8/FKnOP/nB2rKEjnTHwXvPN/k6X+0CwudqLDNEzYJSp
FQjwMgrKE3APsjkdYa7Rq6RkgS7LkFsJvMKaC/HY/OCLD6mENmKBSFaWlI+ZHTcHt6/zHBzNxiQS
bGM9Ii7h8ky0Tu9Rl7AmdHMJKWtZef5rGk2w2hyfRTbbml5VY7gY6PFY5XKgB8oIhISjneF2gtuJ
4PiXM1Q2BokwR13sYFdCU7Npj5gzeaFTKbyLdAlw2EM1ccKnjIL5B5v3YA/uYqRIgO83BAhwHuux
/VzgJgNx1WFqbJKxvoIv6pW5Yr9j4TfjyTmMgu5R7+ar4VXZjHthTZ4RI0BQ8vWyt8w2WE5knYRf
Q3ERBKT5KzJeKPWMdfJFn+lXVB7dg01YmecW30mfIk+ha5Lor2vd4MzzDyqX0gkgFJwPbE9Tb7XW
Dl2qHiyP9jfM3wUHdGnxOosjsfOvTrJOCUlfudD0y5bk9uxI3RqZ4/RgRuPuIZV1pGmMbs5G/VU6
Yx/Qi9lm5by6UclOr8p2u7AeKjIU4W2cICVCj6hFM/RzvxHQ4NpcRlFbLxa04wbgWBS/f+fNy2Vk
gYjRONjPQyI7DasLfLXzjAchLzg/2VGdCzgmICNkf+cCcofsGcTrvm4vLfjoFx8A1fm57YGeEnqE
2IzATAEkG5ejS30tUCmJfeLp5gg0kcUqVrXXTt4CKYyZ02SxmwPRK1OVTmYt5UpWuraSNeKPztwW
zRWjVO3DwBSGQxi3ZNZTVSPnjeP2Rq9iKVlvFlCEvoGAGNv/fKZnWM+p6Lrus8RByDlo7tZ12SB9
c1T4WVHtv29kKzrZHGZhG7TT11x5aFU54p0rHX6uP0S1ee2n6CPA5zBz3K9gNc/s1IKrB5s/DVJo
m7rSGiF110CzinOG0WOteFLnn0y7WTHG/QoVJ4AwzASplJmeL53vctGI22JsDjOPGgQ1+ccTWgPx
ZJTNmf+xn/uXEhUE1ztH+ZOEHLZEgI/nfP8+jZlqhoNy4ti2Ygmm7dSlPrkkyeR5pmM0+K1/xBru
3OaX2ZAjSu8S3jhi07LB2s6YADPoBHEmAG+fZwHiD3lWOjsiYs0e23bXNXqZwK/vEejpJmkRpgtC
LDanh3vpFSqXZvdDKQqcxnqAQgFzW253gvIM2NTiJ/PNw1l5aFDxGgH1w0zHR4dPZq1O/edtrfOO
eHe52p7e/SouMrkwa7nwhgSAD0J/sxTw5/TvebRFCDsXswK74EvDmbJD2fp6p3SMr/tqOQYHd+nE
TsLKxEE/sjgO6uPJhYQ3slN2j9uF06k+bKOd6C0wl8S+CWmgKQx/lXTADmdjXd1MpefbSU2Q5Q8w
IqCISzOkhEGKmK/X15YvAPEbn1d2y1CZL0ePRSChhAMeugara785fWzo/RAAJ7Hgmt/5zyEdQg5J
N4rdwvzWH9kN9chikKsNmApE9+SSTEi3V8E2D+UIJfzLpqWt9L/lyg5GH1oLliVmJ/+pPTDOAtSZ
yRj9/bQIKGo/2MAb8CB6jgIo8MqgTBklF6a9kuoOvchiMRFtjXd7wNRiI19Y1NioE5XmNot6w2HP
1JpvZfdq0jp4ZKLrYZ7m4zypxT0MSOJm2QR05zPfA14Cu94G0YF+jWqn/m+8IvtwPgD5MfA30x6G
odM2K9XqqhY0aegrijBi2mbPqN6j/ht67vemFL9iqT0y/Ns58dU3uK4omTNqlhvIXHc37S/JnAOc
WzI2e4N4q3ZAGEbEJ9N1xBi1J6kG+RL2sTfHBAoWHq/UFvih2K6wXrV/2KFWuU9AF3qyYyBlK121
rpnVP3gBt5dfhuxiPal//QI9D3Ybqn1l4PAyor0G9U2wwt787dk6muYAJ0LNnEoGkYn5kSWxkosj
OLeYgX4DPAYjwP/+ZtrogYRx0KwexqFMsjRexSnVoWb5MEyCvTE5mdhx/2uIgI3ZDljU8DuwdmbX
F0dpaNys3fz31pUAtR2jxy0H+y8Z8gxsh8G0ex5Oz5RGU2kMNSbe6qjmAerXsVVVW2w56XblXcBQ
4u8qcD9cCuFg04uZ421+Je88G9m6iH3TA9o1aRx1zXkU+UQzUmPdl6Wb9BCfEDsDDp8p5/WhzbOH
qrmhVRvIKGc1vbTx8EpPGnbb1yzHibg4+5tJ9Q4YbjcYvWGQZZnXmvUWu0x2XNVrsUfi+tE0ZRJ1
AngvrhY4wQ2UFh+uglnk20QsKjUnkV+y26iK9rqRLTTMI7bwimP6PrBh2VGYT5zpAE9dvss5tw/g
hH4WlK7PRXGP57IeFDzGkqh9qXDahJcKOqCiFmTF5zgfYTcb2L0JhKDuwvol4MQVfee5ehUF9tSQ
CliJF3718C3AxJly8MCbBuM0u8ZCtzmypSyDX2gwLUhjoLTtQdCJeKnyvFHU7ofB9nSXZsT67bi2
5c4clJGXmvWm1NrHpBPTroDqBWs3dl8SswxW9+wlQkryNFIusoQCuoC8XIZUXdNWst4wxLeg+Byw
4MsuOXKT8kbp4i56zZ5cxPl15ivjDhkwOvhO1dC44JseNVaMmDY4ei2PvqVIEb1w27NUlD1+HoiY
wOuCU9PPOh89x2bYsSuM01F2dqSoKkAUO6TQgQYhrTEn0/UzlP6exa+8ljigCKF2QU+pQqr/ir6b
JGSxqVtzrYc/oRYErfQNTt92xp0Z34xCJ1WYu2qAIgpzQ+iLW8n7bbDOKmFzzFzHxzWp2b8SaKCv
JU3/3z+ngEVPNBTih6fEh44jVATy/h6eyYlS33JhzzplkGVbwm+4LiixTMUeTNPo06Tcy7s/VjBC
lF073THnjZ9b0HyNPJIATGxITpbzmPPD3KpL9SOPMiiimUeKULvGYzqAwf4JmXf5/kZqm4vYgNLW
vQ+k9o3FkIx4Oh456IREU1LE8ENiinSlgUUwcBlz5ZLKP4QHQVEaqsnKLBJhZ10rlDxGHeqWLKCH
RTDxasa5DpTGEQPwFo1zzB8mwRQGXBFAs2X9xwBjA9+pEPDVRLAPS0x8U/XTgD1Bs5RNBXEjajcV
1KmQNmzDIqg5NGz/pSjlQ3ulC/f5KRTfXCyEm41zou2zFLvW8zk+UcnhFsWmYjuuF+pUInlnC22q
fIYXx66FHnpK3XtrQ41FpC7nuidpqcaI83YgwwhYsSjhkyHy+yqIZHIC7NeXhgCIOD5Uhio5dw5/
tbQU4mRaPxSoaXuiHCnWHlVcl+gqp1zqDeKZ5Qi1L+WCllGyHNAvOpOZe6mvJIDyU0uj2IQ3IWcF
bf0ttVG0BlWBVCcBbee08qqh8EKT70NVa2xStbzB2JhHuOw92tF1t0bWJM+dy3dgQ5CI2bmaV8l3
0HGnSvsoLNWXzRwbwx/QkaprD1OqS/aJWtAiqp7fM6ZjyVnZkDUAUiMnGGd0ViL2MmIm1dsiMxsN
mmR2RwPWHu+wdDRqlponoXp52isQVRR01QNu2zXyZFROGUSZY7dS4etcQ73axnzUOMoRzeDZN5pp
3gX8gO5LyLPKtVYgH6BlQd3XgvlyKtbeHo6iaow5esUl/23WgYLE5TcHvI8NyqvM5l5h1Q1rXxn4
OdutAy+x4oIhw6aaV256nYYj/jEdin00tfCuoA+fSul309+bMox5OsueZM8ENzqsd/xB1lWyKJeI
YJwyQJtiylEVm3qOWbJdhESm2PfWgDbGaMRSr213dalxO5bOYwlrQcOmxGh8LXGSZkrjQJ/nl9Hp
Lhf7vlGztrEuUNLvteeILqtOcKBRSbOuWLtJ3BbvGf/SFZq12MbLzJUIKGhVMrTvviJsPPhlINQ3
cuNmpPr1fnsrB3uYRR2VR8y94cWRNqmk2+2eWYCv1NsKKNs6KMoCCpbSk6dqaLcG0t/QMFnhJn9I
n1pue2wnssq7jcO9jxzxqBRFfr651z/3oD7O6WSsbo37/g3LgE8JCFeEmWVO+6120tT2cfXMZwHl
pAvpAgarprzOhDeVnLo5eQS6PNuiT/Sxxf3OAcDlDa6oTeTA437lSbmxDd4VFviBrY5WXOLvequY
pGyBh6AdXZ7Tfh4yBhag++BJmZS/D33ZMCq0LhTdPr2Pp9qXxSglBG09IsJ77VTJhCXg9QCiX0Tx
PKcqUptZJHw+c102TTRbqrTUhjvTzQD6AGRkk+2e8gaMzL1DNdRX/HEThAYGRGZQTpUr/Psc9vNl
toKtMAf9W87hCT0SC0AG6QSINvo/RFpHu3L19NDqOLQbUeczfIajAXswcBYpwYYC2N3lnrW6AebD
smEFF8VM9aSNKOO8yzd/oqC1MD8jaYMiN0WSFSUhlgBi0KoqO25q30Nhbj9JM+SFSuv547XVHSwO
w8W24WoA3lu9zIXVB5bdKLwWpwFROXSYoP80eps4wymKKevgCxZqltDIgf/tYgCe/WHMf2NPoeeK
Z/JP4Uhf0qYd8CagOMtTnGp6f7IUVl2VNVfF7rLEBEKpa6Zbv1oy9j04z9m+yXznO1EllcDszdM8
MRqk1j6kfZ48NLWQ33T7R3UiMrtdmVHt4ewNSxNUpUrsSpNExGWOMgzXAa71/sV0s0VGLA+nci0Q
7WvoiQGY4sos2y7ZGSZcvVF5SZouhfeNLcCAO4BBFlFRugq/Z+erVBTjCDNZE+eceRwn8JaOElD6
q6LTmnWJBlT9TGTwPpAO/A/8fVjX+a2m/QNsGKMp4jaDVgFd04KWzTfqGg8Nxss5jLagyLyiQyBc
qaXohZaSOOVtNV3IVejUuZMuJ8JeJE8w4RJuepmCo7pLYdvXuCcOVSyE6X0cJEcwKoY62mEVO/JL
KqmH9jEKRZ28bF193cYiEJopExZQ8rJIIQ9CwnJdEP6b/AOqTioT/Vo+jhofHJEnf0+3yaDG5kwN
xab3SG3N/kkY4vR+eBC2fEHjgQIfYHz1qEYtpP3t0BrIXSFQqBgvxZW7S+11YJGt1CenvLl7edp5
Nbf0AJ3CDyPp1puh50Jz4HskiO6vOPFo88bFds9tyIFlgat/xlcQIknb8g4IyFcIonkgYTAfStlI
RouOn0XlSqmewZoih3KY1DXiNe+COGUycPncnxBUTRs6e8SE7LcqB+e0JXvogHXEhn0ekxYRo9pH
FZ7vqxP65/1fWODGjfgXQ2oJYEBtuzT5eCEvJgVtD2di3frZT5sf9HdCIPgK3Y0RoBXsSU79Xmnp
Thw2AHCONXPSokRH/XYvsE14AK1/Bc3Snzhf9RGLR3jspjOJn+otb+SFxA+eXnf9KlNSe5Z+xpVU
lGo6RJqINYA21XkuaJMGDIPFmpgUzOEqfk+CvYwNR7lnkJEYgIvTp7JehdA3yE/JrH+4/9FZ+q+8
ADKTo6ZPJ1fn+LwcYgFOAtdclj7T6aO/u7yRJAcdKojBf3iMOBOjiPF75LrnLRJdDVZkXKeSK+Kb
uHmxLM3BSYmUISJ8FD8GITq2MJPZJIMadB+spFfSshGOlGmQ/ROoPhgrV/7YS7vtKsMcpb93ZYRL
YHuE5AkOw3p3vUgGzkMRK19gx1ahUZITpeL38hB6T8nY16G7eYz4gcvUxJ/oMEAGGIhnyrfw8b8V
a40fU/Yr7WK5YzaKr7UovRnB1GBRHMwdmeHWp7gc3B44tok9X8TEZXhYLzCVbt4df9l0GSAEd+wB
TO5LawHr/Fnb+ttC1u6Njpo9ypJ1NnTvFa5r0IY4JNl1TTTE2+8/17Amm7QTIqMJklgsPzJ4MZdo
62pXpvcxUtNp32x6Fy5o3mR8G/pVgb2AgnXcbK82rgB3lacM6OHIBZsB+71QIXedqtdL+My9e5tf
mzChXXCsTe710HIlCqrAxuGLuhQ+/FG+mXBRKo215jNc23mG9x1u2B7Xnb9AZyzHQPA9GFkTfmVw
CyhqUbXxW+LbwuGvNJLY0UonQwft+ZAZ+KHtSWIs66mteCv/+s+j7PIx4Qm/+F6KzmKI2qBpbAWx
f/fNZLWu+CSkQTFc49ZqDwdsPc8SxPbaKHt7UHzyXSsK3yWArRtKHHTdXe4fULfULeHZoQKl3UUq
pM5ol8WY1GsHb91nTHNy208ubJhz/36MyeZVyorixmNu1FxvX7xyZznOE8M2nBhNH7qDmnWpD2l9
TSL8Rm22KOct1nAUvdkRTMV+le4Xrb54v2j6RUF0FNofibtJbnD1eWwidRh//RC0g2QqiVBkLFcE
rdw1770g06yt3FtT7WdNEhrLU95BoEH1jRJzPkvT/GSSsWNgFBYxAmA4ALrUVihUMs9QE6uZdH9u
wU6yBR1doboPbxH9X1NlRAWEfYuSttgujkt7/b7O/6WvhYK/WdqhfblHvCxTbO9jfDVatICZsVA+
4Po6RqfDFFKyUbV5pAFDrLn0oi9itrxEbPMqChl5PBjXu/4I/j+rqBQOoc8gxhHSUOulUD8Pg6F4
qCeXpIu9qmbQ+Rlw5x3eZp0LS2CiB8nRQ60aNnz9sZnhlKh9MgoWXykFT2AuFNx0K5oF9czv4f0F
AZJgqLfRz7WtjMPza022jV+YHkrBkb4q0HS1PIAwUyputFyCzNIQ0Em3E/AGycfEJSsM2FaRQIn3
XIcNXGm7+ciDoIIgcGh+R+eSNtikoRtzSxrTOOWo0bTfESPBijG96fViklh2TbKHrzRD2AyU17DC
GWq4Sdfo2G439xGQ3a9Y+Y9KxlvySEZhufJFPLa1PI6gsocVunNEbRIvITaPXOpWDiLw70pth/B9
z2goZGQ7cHJgyKn9jza1bYo5G8ztvb6zQSLuwqUsBVdRUvTSiG4KAEPk9Zpvpc1tjUFkPBW34O0q
LkRIzfyBRBlTi0d41rZXg9yAZ4Y8vMTmGvXiqbelTYfdlP2VZ8aDdfhmAgxaybeeY9JMA4BIauD0
zLxYP/dAl1g6Ljc6kdxXajmatCihdRGRlYg2U0PEE1PyChDa9IQP8t9VwQnxS497ndvLQ4BHztcI
0jlOEUlE95cwmpxLkNUQl/7Y+Z/s4dRYgCedHJyVtEIP7BNm+z07u2PmkS6TI528ySWnnRrktUzl
SWEyksrbySV720zoBTUUT4TTtNrQLhLIxeIdbZS9AIeRNvRIWON8DKRmWZddSkUjsxQn86BOPG+a
xez0kncc+poarfhObkENWfZ2AmwFod/avl9Y6dMnkUrhQ9abGA+o893wC7nHce2hodxrTtPHRhoU
Ftxp7nEKkxcl6iO2mLLfjXb0ltNa0c7LaFN2Rb8Sn+e7zvObh9CM/XzhEbnSFjuC26GlyvwPIW8i
+p7SmAjKjGQDnG1Q1YI8uE09dbCLogzycnNjsCe5sy5NOsspNvrfsYnNlp6KHvwyXyAXt3mLzzun
4Bv8NZoD886H+Xm5gDxcmSiqzgMqqNVzhzFARowGYM0eS9+B8McW6cqyEDqiv5/A+o3i/Wp7eEgi
uu19oxHrJdk2UfnjZBNW8HsOIKlnUt0nJ0lLs71B9lQI0EUqJT6JBzYgLNNB72CqIW7jsSD91zyY
v2mwa3B/wMGtMVRg4xSabXMZPrp8PiZ/1s3oYtU1bDCK3cGQs95GaAt8mNnDO6wRhYe9StZGG2T9
8koZ25Us2e2/4/vxpYfQ1HczfrrsZjnRZwp/wTtOhtyqE9G9yF+be/K7zeOl2cfqxNpu8hVAZM8Y
+LzNvIQ7liVqQGwp9l5xeE3qNkgmluosv0hF6WBzzVtyYkWodUYfq5V3x2M6SegC0CI6KjuPCexi
TZFVXDBa6111PuIavbC0/JMrkNeXUhsLnW28pjS5BrfI7pTEjPrlEFwhUzFmRDb/FdZgFEQ2K7S1
WPKBi23QEkRIYHIS1zmrMwUjMEOLoeqm8EONgh4roAcHm9bK3tuR8iY9OQaX9DB4mIj3FuvJapSB
+sTH+GRA46ANZODyttYqZR8qRzn82YT/AlKqpdo3tTCy6TLkMC1uwmZs284o3WQN/486ahXsbE12
8V+izfoLx9pEmbQIG4pHTDqNNR8LwOM9qVZIiDWQB8vM2agFwsf2Wq1+sgiTEm+neQZ04jN4BJ9Z
i6TdfEgKbRnXgkkc6B/q547JEmrd3zoFQMhLy8FTDYjzBHjlKfIcs7tqPeNHRulGWhB1PWgW0zrF
iMhRZuOK9q8FG/QQStbti+H88u8w4fb2sYF7FE+z4iSaILOfWGOllIoQVZWvVL9g2nAF5CwvmSpH
31aut5wcJMlEv9/Xlnf+0udHqnKLSFi00hzjLXL50rm0haDGyOwd5fKL4geG2yfbiH2Ra2aHuBu2
7Or7ofXtZxSwFIQZA6NwCwikrKJI3lOMRBg6bVmmIsrpTcR8ojPfn4netG9kpKFERFavq/z1gG8d
sNefbKFNX+kx7/bXDnvBpeFJwnLx6ja3yWLpR0Q2p6/3N85t/x6BRRuNZselGcAgzxdbNGyC/iWv
uhd8GMJGO1Hbn5+WexjnahfpeR4nqmEmjZTUcBl31WoPdd7fb+CevxL+V0ARX1ZyQ9JvtCLOzssQ
NubuTrY6YZRdCU3gdyZK0xMW9ikXxfVDnOQwcgYKqecqLmYxSYzjyZldpYxA/1c40LM6UvavkGPv
Nzp060ciTZalGcuYxSc/imLwla5fR0klMUDeOSGNGhT+YwygME9iCZbI1g1hEaQcmbDw72SlytYe
YLDwcSYrYT3jjNVc8AY71lfAEGtAmDdEFqTN7eWneRL7EUgepMr/RGlVVQVY/D1HfctU7ncC39K6
oJKszsPBqC9B86YThwi+sj0dAeiHj54I4TQra/cMmV0aUo3EmoFLZ1pC5Aa72pqfxs0yMh/cGb+e
wVbrpE2tQBzVTUSH/19hvNdp9YdUhx/VyoCEujC55EreuUaqWEe+BPe1qj/5IvVWaBVP2eTLvrdu
sF4+hRSxRA9zmIhPqE4jhsKz2bi0gDK8aHAeEGN1mp6J3d+/IMBUtsc5VBIEs+yOtA9pa2ByvAII
hSQRhmrXB3F/1Mteu1N+RcQb77f+/WDv/dSRkPrke4aM4rBS+4hg5zx0CKqyyTaUKl1UEecqrFSN
QkbMjiCXo30S6uSf2H+diwtEN9bdecPr38XMhD5gqDg6OCzVZXxMn7nL/0Wvk/qOgjq5D9hVHBMI
reZqkqLJhfpHOSNMTDXOMj9CFhMt28PwyZz8oKHwg8A6N943NjT7BayLhZGghX8+A0WyEvX3wcOz
TMd8dh6wTMWU221Q0gR9TJ9WACdvBDJSi3zcPIhgB3E/xKTy+ZlodPyqWXEtHwWloyiQS+jGT0/c
tH++A/bhrdblLxi41FZ7rqrIxg794rsxTDjF0XIL7hL6TcGI9pqyvVTI2nfDRpsNANeJJ2cA7MjF
f4MdAJ+CUFxirnykWHp67+c6y7HaWijmYQR5tgsfhGAzVLAx0wPsWpLEcSZwJKz4NtMo1yX20IxP
x6udui18/vGpeYIXRYrgHsE9kj5acO2qnFnCZOTzV7nsiMEuMXaSJ7p3aTyiKnNrRJokrOQ80C3N
CI4caFfJ3is5GqT/M+C8PEROFrpEd8Gryrj1clgFrMV+2NAARHxNNCdg3018OBnu3POOHVmHUb9H
04ReLBvqzlSVS+Z0kLYKOHMi5cadEWXTUq0Uvy2YUufhR734hEeT6O3H2j5wc6ucwvbHYWmZ7lNo
Lu+3S06A7zDXgVPU2S7sjDLhh0GH5Fj2ysoOn3xcyU8SU1EWINeP6nMJDyM4/oOPBmFKeegmNXZG
urormf/61oa5lppyCjMjQ6U0hkgO8p1yMuA3NJG4EwaXKoGXoQ6ROHnM29V4wDFn+jwB9PmJuDeW
SSyGuToHkavqGN1ctjT+PEbcKTFnfWUlP0HIyADcg/rrqGLT0tfs7gFqKGPcWL90Vmj6Y3xZ++LL
7SNcLzLPj6a83J3kzqaeT9cTGcdRkXlAUQAvo3JxAkV8LHmMS1T91JBCgDmhun2ugbv6e5SA/JMB
ln6lkONmi5R8ZfW5rzDAVIpmj8X7f0c3KOkLtzrMrZmw3NTvVT9pALbXoStG7LvLoGqYpWGJH6D6
SkVjyj+1fVSjH8PFPkwmj1x8ghkMqtmGA+lTg6beFHPfeY8kdflxAgGtnh979p1yl4QQDTI9qvMh
sio9UP2J/HUI59DvSQRxkxU4sNEeepXJrnf8+GriENoEDTYs1wb24Q2WsT4GKjj/ZE4HhA8k2J5A
yItVv+6zKRkcTKYyzGgrmFWS/liycdJy6Sw4Ug3CFYest0EANjP76amp+A3JhuV2+lKkoEp8tNy5
YPrcD08e+eLXm/n4uZbHwyauoqtI/qaAk0nX+asyf9llKDVniF2wloamynZV6kG9U76GC/l1tQzG
F3A5NUTXUR4y5s/WaqYkjGdN+S9oCx6craGaQcm9qFkYUBb6BtPeKquFN1wM4RUhUf6zBL2/VX2G
gAuBl0nwJr+tX+x3lvnwjp01vOENQNT2YLfnj3YcATFFqoP+ilDOZs+bILuNUT2akUZy+evLGkSf
+BwYy0rct/pRvaEe10p47GwrN2xqdVP+VB91Gj/P94Xpi6nmoQPbbIRyz94AtNNPXOsSUZJouPRE
ugDkcVukLvDWU9h9hN6nbei2GwaXqrTvUSn1XzESxpOBMXhqefvKwx19VlGEB9VajorQY0MkhJUS
eHGOw45sBysMR2Uj9zV+2FgwhM29g3mAJdSXGIpcj9bKC7CipTiu2LD1Fp7YACy34AvoM3lid3eu
7RYXXU2+3q2GnRETYJXfA8AOZQ9DUreL3aUZvZw8gh0VXeWlJPSnJpVoGpMo55Zsff5jxiVO0oCk
waRhmpjv2J0eLJx7b/H7SGJ6OI54SShHwBME5HH1+cNmCeL8XOnjY2jtHZPStEFN2LM8Ase8T8i7
yPQwEP05IhahYqyyGQ6Pdwm/We+XSTQcOXFxmLyAUYO0KS6A19t4rP7PHf1zG8GXjE6eX9X2JatE
vRqh+coDt87Sn2rShNe207fEXrUvbQ/RJGh1B8qYvcAdzp+so0nyTTh9zyZhnPFT7N/bDsIOQYlT
5mO3X4zKxxDCizgn9I7/qYL0xIdN/eIJAHxUBamGXuxuy62xuxmucY1ld3CNR5+1CcTstlYT6wve
vAIMCeFWNT3BpNfecpD+5U17DHA/NkHdU3mv7JFdagXU344wZ/bhqbtUyALYbbaK6CMG6FK2E3b7
fnFFtP9NOTnQs9eMusu23Jzv0v/s7adsSThI0cnxRrkJXba8iZVShdeeyRZE6NcGPnWpkqwTOTYf
cj+HihDF8CkFy2K0JsQTbAzgtVFMJvRWJunrpRe0NpHEC2RYXVUNNWTV67pHT/umgsTg7ImkM6pD
WP4pvmWVrrZAk5aQsKBWqDYkqGSQ1eGvPhIInSOe9HYSD/wVQrsMYnV3MTk39aNnccN2ZOpv/DmJ
HnowqUbXTgEeriwV0VlCfDn8/wEeRrz8q/hSMqT5vtQcy8UenDaLCUmKrHJqbt36Gce8Uql2n6hT
r/owEiPFj8m9oaMtjY4TuHF/dMl0H7RP3sToffcdDJLqoc8JbCiL1gStoeKKWcuI47Nn4gSBZpgK
Q6d1REuPDHLQp6/jOC12xGwUwwWdW8OgXYxxlyNHwi1BQbLN8+sf82ti6g52eos2QBY8fSa6QPhD
Bb2TqDsoJB2JBJl3vjNaCMO5hEKt0lLL4qVAuLfZhh2fhNZBV0I9HX1J6g/U6tmTqtmBgjJoe//u
07Lh8VTaoiMp3+/snBjLU1rCBZzWucx/Dj16JCjkMi5gEHwGRtFF3NhkNkGPz9rAx9F0jnbO+QEi
1grTOpmZhZ4Ea2lgL0GIuN0SgpMMrOTNNCHzUXWWxmJUJACc+e6hFSlw1bwHM9abmMYT9xvTyR1j
XYyQbFvpayrSH2Qt4OLVYfuogOf2DhXZBBZ50qSYCalGapAZLZqH0VTYcDpzvZNKXjpszwQaHA8t
1Vj4dGeZuT6i7G954oUXgtbyxJ+Sui0jyqPHhZ/hcVUrCL99oJPiIxI3qjfPKCBEWfpxsth8n0P8
ZzZQshfoYP3nYZjibY8GsLM64DpWcFKYVB812dWfH32OIixdOORfI2ebXIZC+Rp39ZQHjVZHZQ0j
K4IWXJUkf6K/2p9Jn5Y4duMJmmZJMnxlgHyD3YlIJ30c6iHxywh81KOGln41TB8kS5xT6f1zMplp
cM4H/GeFzt6PBVk9aWNndnMpLyOLsoXTXn/6GW7T36eMERBfHJb9Js0+yH9krUps9vcITjSgAafj
V3pfutDRPEak0unsAOuPwHvMjpsPa1jXBxdAt2csnRPrDSuEpcA2lHAG+GzV+oQbTiXc2eRfRxd1
mX2OHsw1o33HmciuRjT2mlyCf3GUMOlQ7z5jkom4nJgh/83YNTULi9T4WigjwKrWEqOldHCB3Tek
0FetvG3VIv8XLZzIexX/bASVuJQQCH2slRVHLlMhRmMmswZ6ZF7sgw3LBCPkibA3F5zQgUQoGkZa
pxWuIGAySh/MmzAz0lrYHUrUXlPKCuRIQO2w8O/UigJjlDZw6mCS8uHUijEIjCJ+2Vh4up6G3To4
Mp8UrvkPAi+IVWPjA3+LcF0JrotApVoqPEJe0rjpqB77HlG9fMAYFV9ifYeeW3/m2Dk0+uisqFym
siPyxNzIvzkLROz/FtaSGZs1qOuebwhnxFZJt3Mr5jqJ64QUJnCFfaroJztYf3roJcM39Q+vc0Ug
klWAD5tQhYoNKA5cdaWvd4q4Zt6mAUjt6b4EZ1R6pxtiVUIA23ioiAoBFFQtpFgMhXYYjh4pYXta
kmo5ocp+HfiODhHEF3gSOVx/1YMYqZD4mbtFSHoSngCNXhvXKAP696GjABKw9yzFFzCUjeU5DeyL
B7fc1wy4+o2QfmryWCtseEIs9vNcWWseKXD7xHo+OVRrfKvOdWwOzrEBKHegU1Xfwg29zImgH1vM
IlowGb0ijrPxsMgxf/zncrJvHZcbZN0cbwjCA/tmQ+m5R7PALo+KUPCMbjQvBvnTZyvhJ14pN3C4
kK5kTJafy5oMH8GmQSUA5QKaHouDdwpY/HQnrGBx8m3B09ku6+8Z9Ew1u1Dn2Yvbt6XRF15G6WCL
N9eS+RFjDvrCDZajGdqPOHapIXBYsx37RERQbeRasOa0ymZ/wswEM/XOlgp3Qvp2e4b6t3Gkf6xg
eLsKpj7j+LhfNuQL/iLgmK2TVLZQOgkJTYSoDZbDTgfess79aAMF4D9+gOe9E8pASx5uA4CB04M8
i+LkoWya2MlEQ75kSrCb7iOF56eQ4JXGaSN9MyM72oNPT56BTLy6q3L7ZqMuZRcy+QdEe/k1d4Ig
3mz78jpjx+MxnoeicnMNJTMivjN6/DU16gTyllKuuUp7cxspOess+HzGZ85OizKMSuIlTmnoVEAG
GJJakcLcPm1IgyzMiqI7+IUSsbCHW/RdJlKPkh23kxrijwYTPfuwqHSF9tejI3l24zMywK5iYdpB
ebbWVFmkt1hkg45h+Q2zgUqCZUff2Qm5PTesRsYyqYEqut5R18f0bKPortPRB1mVv0oYPA9cf5Cn
YDxqH8rL/laPsSU/PYGWUtfwTwXNIrM7qJwirOcxjdqKTmoLHYnwdovf07gWvPvb2AF2SXKXXDiL
4l6NLdvsNmAtxtkEySD0ymwXWYeLaeIJ0JPVXK64QCDSMO4+RRrPt9GYZu2L+1G7pfHgo5dNLY1d
SXixGn7V/OfB9Uyc5q5r2RHOeuyUnQN13tTWFEjc7Q6sjfboiTHt0LYEp7y8ya7+DZhenOukO3wa
Dv+evbUwtrY31Q2M7WrD8HpzPVk3Fib4Xd09laC4DXhemTZZUX5JSIgD9JwkF2GLIqJjWLWFK5+E
O0wE6JxWYXiYW+H48H0J4L2HHZpLXqmzsDFdKbOF9PIgD3fdhvFPPrWGmKg2KrFPVrRmVmWDbE0w
RqdK2VjahWhAYpDDvSQ+Ey048fK4cYiyLZ+3T+9MzRo3zJQXxuipVBK0021X77GplJObh/r5eh4a
fRJpTthHwXpK7EnFJWvnwWAlPYe9yMl5lz8f4lOYK705fFGD7JvSOZQYWRGPBzka9yxAV9bW18u+
WefN02Z8CRwxK2XAQ06xa3QF2gOIq0vDiPRDRzFQFcX2f86AiRSLoWAgwKy12Gs2K6nXkOPgjvyy
VK3c6I8a8KUqIir+6G9/o9VmM+yGtwFeqRVTRh6g4zNftDHQsITihguEA9w67wggJa2cnTDEe4Mr
CrdNi88uY9TJT1PRX2O9+YqOcDPundnWwl4ndObcCN0fwE4YvEeRZ6KZL3OgBQTtYo99mAV5Ck5f
YzIyEks7PgAW/JeqK58pyWCtNgDaHqSAZnBKaaEUA60YLeNIhyqtfRm65qxgu/xog4DIZKHHRPyo
KImRYDDy1C+UBKc3PAJV7OjywEg9aLbIyKAkZIkYjzxQ4bK9EmEEgzMbc1U76TbSP/adJ9ksjk6U
08ZIjw3jufbURjOhXdjx/1iodWNFRAkcvcy5/Jz2lkQI+1Ycs7XWM5OKfUVvA3EQK91bChaobMmP
e9nB+bU+d5sBZe3FmWi8Z1HYmz5IZaKuSHaPbWU0/H0pxfO8GrH9FkLoBBYk4UaR83iMqnl+nKRR
/M5x7OV2ix3EdJZDMoh88UNoAnmJzsVMNGD+wM96nZO7k4SxRT4VkEZYTue1OfqwgqnFVM7Ch6mg
kbRdVRShqmyJX2ar/On6uK/RXQTDuRhoIYLLxPsCJ8SnwCp5buE33KNImGsOh8w8g4dAL4Io+VJR
X+i2AU5jAkiM3aKV3gF0GYqbOo+o2NCU32xOSnUq9WcK9wbrhCU9VeHnpIZY2JcPZa/1mNwsO7PR
ctzM2Z1SOKPEX1nyvK6fp0sVjWiH7XsVzV2D/z5wsieWXMwuI42bSj/jK+EXoaVEuCXWoC+0tmjZ
hBstq9pOP1b5tIJ7BhAQm9PWuSUp+BkHaTd/fhiIXIC2CfbwSn8XrlMce22fkha27npOtloeShhA
BGzB5SfnjSRLxnRRKkizdXqX2Bi7bhheFKmO3G/xYkySu1yQaYX/E+eAsMiUs1btZCerlvlIMjNv
Y/fvEm6M1Q6fa4mm61Ol88X2TB60YAbGUy4wCB2utUKGGVvc+VXPj4S4XH7FxgxZ3IA9+MS83aqh
LL1M3rEn/aNUuQMBseElpf0Y0nVvS8GSQraIQqaPH99rl76ptScAo2KTStCkw/kNQByEhO4qQjMW
t/yW2s+Tf13RC7qvvkwnQM4a/4FTgBJ8fFGBC8KwGNjFI1krrngdYx2oxqkiyz0tOcxcbxta4hpl
qNsprlnreZs7QRKyfXdI6WfL2SJ3C/t3+vYgtXtTi5K6LsKCo2Eh+olxNfUqhpZPKpFwTDgEiL7e
S2aEIcz4tZM4H1Tlo/96TGPQvRWxOkuqdla4o6dIbIpjMnRoaDyClg7otM3fj9rWDvpnQWZgSNtH
HGsooHG5PkWSMFJQivJ1fPUkHnFoAr7axPLH6PtuGkf71BR+9vLGUUhK0446+JuYFgkK/blfWtgN
oZFj3QN83reKUsF9dKvx84zTKtZksZoOk0UG8is6gck9S2HwDK7wRY1I7/mDo5VYJE0Z8tjRtlIb
19QuAkmIGJ3GZHEUwfbgk1sUddrNfni7tIr2c+Z9Yf9SkKN2LDa3iq7caUrd+Kh0GnkYfQBtMacm
bYlk9vd2vdNYMMumls6GlG7vc0NcC9bpmOwtJKajlFtBrliy0CfNxX+3xDFJLu7Sxw4du0WlMa47
aNDdVJ+P49xAvX/K5t5FNrVN4iGDtjFeTRgqZ7K8GlywQBDWX8WlUXi0MALb25RtF/65reuOQpl7
SWdSHeq7qOowcg6cnPoMNcy6DiHkk028/QY0ACnJcMEAAiLdmVopXwsdV5D016124HY9MJuOmC2J
ZvzsMABgPbdPRpTAJaD9UD6p1JFK0TIBXYWV6rkYWn/2iOzae00bGLWy+x3J8rCKR8itCbHmGuzg
isOA3xRl0tIzCo5IyxThHn29tK4omjIGhlsbBjbA8wy0sSSacN4f8WYtFeLXdqpdxxQ9o6X/2b4P
UOua16yNq9miMuB5qviSWSgMLYP9iM0i1WsIZfTEgCwfV/K8bqVEpe6t9heUkJI/RaMx2kV4Tx5n
TBx/bunK6mDkT9EGF2N/okC7Mi186zExusCzFmcIAB0N+D4Ynvo9jBwLQGBC2rcUvxUGLELqRkW6
DCVDNe1hpkRcn1yp76PlqPtCpoWW38YTvWPeFWGUF8QRuOQejXUR1OEagOGwzNapSqMi/udayztm
ZY5DhLQnuoqnQAQCvVzD7wDVlJo1lh/aXAgryi4pEcnHy9vCygof7XY82scOFxNvwM9Kjnemu6nK
e7m9mFsoixg3vWqVpCL9XUmS7dC7yYe9ktHuDAqnG9TKI7Eyh1RWkp5G2GdiAXOfSTCXoPY/b9US
Oos4yIaAV+h1AYMotbJpuVNQb8K6/C4+cZCc4P0xFMcphIvKiNYyPv5GS3LG4YmRzSOrlTgBdbSP
kh8suBuAtW3dl49jLzPvfZMSPuVSNIn1IbO0IgSOzeYzjXrtztu4rCqbEVzguFigL4+Jan0T8Yk0
NTW6y+frxO/QUAtfay5LV3VFuC/sZcHghKmWP/pdTWcW+f9OzhBufaAKyhqlCEhaMTlFdaf7VGtW
GK6RCdJv5egvueci1Uv7bwPBsd4K6D4gENoabn7Emhu/YPVHzL9x+pb3DlYDp99rZSZHK240vHvW
X8Osc6+/chGwx4lh1qi/IvGyuGwVd7E4xsBps1FuIMdq1eQctOzxZFfcHxDNVdGF7DPPq8VvGmRV
KtpMveAJr7SELR4Jr37x9iv4Wpm1yz3pNyFieCUKv6AkF6q3akAv3LOZu1RhxE6csK2pfN0HPN7p
HzbLOf9k0Gi1CDAHNzpSizpy50NS9AmuXvsxYQcQwkhL8gjvSCxmPk7m6Ce1lyx01EPJaZZGZbz/
lXXcKqQSCCJ6KMsgs4scNiraNoV8Rfjd6jyMirC7/JuLhuwOAZVy55XLHPXdRVrtV9RcvFYFyak0
4nu0bm0EiTihdSjaGpOPIb9q8XJrWKDPXSMc9zowCSTecuIs29fxeqqxir9eMUrzKSNNXSHLtgiJ
LQETNwDF4F3RaX8eRfLJgUdLuXdoxKMLIU5tl8DblRfBkOMSNNgkgR46nYEkXRCPLZft/+s8wkkC
Wtl55SAj6yPzlDsh/nQM5X3Vkh3INtet/1dmDJUHnpvVmhJ1fLavqtX7Vi02/dEX/tZBAVllMYob
OkPLR22gnCQFqPXoqz9oJ/9UKZ8TTTybuhIQRAIf66l3yfh6coPUoYHK/YVjsTpECSmfotLIFmNA
9CjezoZrJzpQpTTvbLKvVmXGCwWo/FoxHaHUWo5RRYPbKD/4wJjC9LSZaVQ+S/miSuTN9MX1vkyj
GctfmNtsP251+BxT+Z96cGRt9LVtD4dzgeYvZkH9mPv2VaZzyu0zQyyU01aKHA13tfaIuGWw5bPA
MjXYL8R7OgEJVZZHtbn/6VmazD0CGOLJOrtvchrwtP7jHy2DYPBDkFFLL07DsV5jQMgjr2XtlsT+
qQJ9HjDpUi8duBVmOiFr99TPJnQ2ZpLYB3/rvKJuG27cC88tpOs5GpbTxqIhdUmV3qrXwoEMiGBK
gqY5l9XHg6ikNRXyB+y9xeLpiomWopnPpoEFjt1jjrAATLW6J5ydBsQ0dIK7UiUyHOjfYWbQ57YJ
mN1bJkMF8tyqR1inVtdIOIzA33qC79EUrLYz4mq7MtusjijlFhEgAqNdLYUk05WUC7oLJDdX8RBL
fZILIcpd8HNczAB4hTOR/E/bfbd7X1c5Oje/ow+TheZJlNPW66vv5BAnSa5bDrPbsAI/bxGWIic0
R6rAb7UfZ4GTstXCWHaV+vXSnWZkTijVQdE1jXiG9RJtBpKtYZTSwhSXhhiSzsfYkTOhbtQWXemC
NlPbCJGeRfMWixXEqbLSiwqgGjMkr+PE/lpdJ3yW+DIISmtErdUN3pLPneGmEp1Nx7GWHzzij/fy
KX90yzSALmRBdJGvOGuVFbrfMtRCuSKf7rIisz6fwh9bSt0mTUfsGqdQDkysjdPIM+KkceC+ZC0G
vySsXX3Ke90/wvQPvuMphuiZYz/2VhkCMnvOWa4toxaKLy3c+VPODZ06punJlmeKYJEuhGU2X2Y2
j4amk8bZatBF7w34EyIT2KgmiGlasJThcYeaS3CKnsBspxMGV7zGpNiP7u2IiM1llUAGRfsW9ku3
ZBJmA4wTuscyECrG62aseJI8WMAVpaeMZOr55Zb+9HStKndmxnNOxG74az2pCM96zogPUSADeCfg
ykIpRcR21cH3pVA4NibwSbr3S7c2oK7RWTCaESi4UC7tKTEvPWMklYmkwF85TdpJQJkgym7wlVPq
0hzsCIasL3RDG+xf4KasuI1GFDvxeoz6qXfmeg4xpAiiit6acFuth216iVL7zfEwOZq3qeOwdIFi
m5NMw1iHaiG3irO8ULaYY+XaYMGu3nxPiik0+BInoYpxhe6j0DzbYOJXjU73CnrOYjCJbu+Dk02s
NqJBTKGykr0Pk0YrD/HjS3gbMs5YzQ2b6PfUUSG90uWyJJI8TFWXK1RXiaEtd/VUR1oOTJGpP3WR
5vaQTJIfXN3Pd6S43WnBDlzeCODsHaGTBkR8t/a0krd05XQXW+UA7bahzs09tc2iqdbhaQqeIe5c
5zpU9xvdXcjv4fSa0qrd8vbo459Zh9XobVtpVnxSUBW2M4xUtIPhhhrj323NMH6+dP3LySeTdukR
MUEk5AcBa8f09NcbqYBe2dM+opvKbWs17TneunlW2J+6b4I0o4i88sKT+SRnvOQ5+fNYgHjLtRLq
HseYX6a5T2t4ADWXpPKGKzoIUVGtS26Wzf8CK2GNlHwSNBzm/Gaj2ppwnDiEir4yV7kLkQBo1eoF
mGnKZITQ5PTcfJ+Iv713nR0htWYilgomWxX9G3T9d51JlPTGFmXpDa+3v1kch6kd7m3wC9/O3XP4
D6yJdELX7e+VuBiEmE3gmd+kpsDS+05cOoiLZiWN83E3uNo48S/frDSgMLQvONLlfH6joZHZfpXl
yAlkb9IE9jXeWVpoUN5igDzyFBc+YvjYMv/xlfnuE4FDMkLvpSU+jXDFcpZ/8EgG87hzC0uYUCi3
IJM8l7DErT076R7aSs2ybAE8rUTD7lM12VG7BhcgLETeTPWtSP9tGW+db4FMi5OLcMsQ31e3+aRF
yb+SKz4cVXfCrTprJAtirAbkE5hw2Rs+H7dnkTLaCWbFJ+UQjs5DtsvIxUWa8jpTn4Sz4hG0pMYM
10GEEJBRFsvbrrmmIDOtrOAWa9be6+impun2WXwNH+YawUDHCm99qEz83bKKsi+9FZg8a7Mk0ojJ
WLy9zjHjPKRfr9Org4wapIYa8pb5aUOA06paiiTA4k/RdJ2dCOpVUtc3CEIrla9C7yGiA4DJuJzB
HZqWmfpKYtHKzvCz9SqnBdrB3Jb+KGhgLMpx9mFAWYj/p6O2ssqt1Qt7XQJZ9c4NznfCS1PwpTYL
yYoG7Y3GoNmLo+Zg05iflv6Man9MjP/ay9rjgJB5Hxaw/EUuSChryIn56hLmmq5dybNaZCaJyFHW
iMNdgS0G/ZU2fOaG6L6kje6KZoY7oPNJXwD+t5kkLf+UlS4UL11W0fT3AGEWt+COyzS50hcM2gdG
MDSc9434RHUtVtdruxU8YPLCzLReZwhZ23FTZdqNllP34F0se7HouWNQewakZFUWwXNS+MIMC7eb
RNIhRd2yaANgftkU0j+dV4AAGQWqcNRnEfAzHQeYfTmXclcGOyWTRVt5sz+9Dyf0bf/La5EjsLDd
gQG89iJVEQYVvuWyjQSLyvKbynA0p3LQDTHWYAKCz39ruKW3KzgdvRJaLmn2CC+IyfYPelDGs+b8
hy39/JisHvNwl5tBcbT+7oeAULj6KWJ/Ew9/meYdl7eBy7tVFjdTHyTvmG7MEL/4+10AP1x/6zkG
UWMQJzupQsy0fJgWpxen/Doij9svjRMKuUHugqzGrkU4uY8Yizoapf1ofkhHgZ+IkhijjgidjrTt
elO5VDef+0SPY8zPWUgpDhTZRCUyKejHn51iwNzinSHeeQntE+Q7RO7PV6EiWvm8TscJpuKGXkGq
lnKr4260tYz286obsq/f3f/m+tlSlygP+rlSntJGLbBK6jOxlBHoCIQT8YWMQHE/OjRthbUpepD8
P4jsCyMa6BWb3DDX1hbWVdwSpyxoFDruG2RaNch4gyANKXWdz1jNaooWCZDcPcUOENGRGqj3K+yD
DP4xDoQ6TXJoHgPb7F/Gl3LZHtdm8x2rlSsa2+0pV/7SsmB+0WI/2h1yTcdpNWLiE2VV3nFafvtu
rkgRHU0FXbsETvqYODSJ8s+NAyvnGvc7pEHhkrs8fvHNSkVXhrQ2bFVva7bsDB2/lvNJ6+qQ9Bb/
hXxXk027h/1fZQfdf7zDUPSmfqLvd0TjX/P+DfnzpVdRc58VrY9o1NIX5hofr4F6oIUau8a5UyxR
eph9/dtoUw/sNVGf9nBdyhCK6YdsthuBNLkS+9Iu3r2JOnn+KWl0esd6VyYwRLVaZqYqbThbasPs
C7Oshp2U1Jc5rsCgAeUoqtvq8DY6P131xIaPEbz5GO20chQWFVN/FSLYrY/lcCKLbfnsTGKZV/e4
KoyoYYT4VS9BCdmd8C92xjOW7MXYGeI5BbuB8QfFZptVGDqIlC+4XmYA92rE55Jsdo2z01cVXUtF
OAKuLQI/2htDTUpDHufTDx8JFbWfa4I1tXlNrrChyYdO9n/JDQ/uDHExscpzITOqwQsGkIwOehnM
TTbdUgNd934Ss3Xr18nKulUBGbfzhxm0hFfbBr6MpJpRdBckJ8Rgup8uwqZP9R7vFZbtV5qT1TCt
9HEmZ4cpWeXzUv7h5ALdN+3qKpWG0MqD3pt6cYNe3zXCGGyrBdB2Vp0Ksu1dQ/w1bpL8vqMsVP9J
g+FRkF1MDAYpGsp9nnlIUS4Dqvpa2Ssf+j/DVpuLMZAYsDWT53bjyyCpqW62zyt2Bl+ZLSJgDFXT
VUcAJteRFtNzpr8FP/ZbUfqB67DDqqMq82W7JpD+eHlRh9X2/7q19xa1TRVVjB/6a8ocn6V7jng0
rJ/DZ8LCX0mbVZBQO6W5hJpw8JeBuus3Ow3d0s7O1g8UOe/NcaCbwK2BuwE/asec6zan+fkDE2Tt
gsOqmR+ruI0q9y/X05SaLRCN4vLbdNJf3hQwn/wDp8NsTn5x7nWS2nKaLy61lWkCjegTQkMb6WBu
RqfVXxMMfB2Y5H2HeehMkmy8XoO7rj6A+nefaKfxbCzZ721B9bvnSPUSf5DBKb0H/j628V2Qe8uV
LGPu8UOpdk7oqbJbG1xnxHNNkJnxhAaahCEz9j2i5KzUVF/zDE3mR45xflK6aIFXD5lFTS4tHhdB
ujfGyOJZH4mN15OSN2vAghpd3YSPFqco7dJVozsDosZ/u4w3iejtyztigJgnsxFHwyMO3Sen26kU
r/820fxWLk8Qc4nEaT8Ogq9pY2HwI4nhGFCrLsOjFulz28usTZyRyA+Cw+6WBaKt+CqFS60VFZU2
D0PagHTXxpuQWi/gG806hrpYklEZS+b2+RHhoavX27xg4SybHVV3M5/PgmrJeRlhXAudTN8C51tw
mRlCUviDUBt/y5IdFUK/9wykpwiyrXJKzkB5cdn63z0wMXpJOd0RI7WLLsDQz06cB8ZjPzhijb2F
sEFesFUR1ZIjUoFgF6Bd42dhJ9pARXGFwADFfoifyJJHftP4/EpOLJq23LWc2ATjKGPik2NPM3yJ
BU4RtS7jJP2zhfG1xR3pixmg6ODAhyn+jx5tL4fqxd2ALIOy8vpO6CRmBZnktvEXxec4BBNq5fwp
DlRAUDTLTIMm0QrTBLS+3gjHJKFCDQkclYMEm5BcaJxX7kpyqKagkL15dd6E1Q2iYh47dXDKjswu
iNHAa4NPXM6HaX8JNgSDHl368A+mXErg0mQauSCGDxU8WGebRVNlfpej8PyjHVsnXahplNf0ZFEe
t967b71Lp5/SjMvV9GKfeKGPca2kre5rOgRWJSPQGh1+53KY3roBDnAwSzChT64JlUv/jI8jNPcD
V+qw9ufvBhVvd6E52RmqLC2JevRl6/85GkS3Vb/Fl/lg/Ok+ziHgG3aY4g/YHoF6rqpB2K0RJ9/g
AlZLo6F18ozgyKJKh9nbGSNCfhJFhapJNLiAry7z+kd3Id3Xz1PQbhNJQQl+rFNfLxJnKQZwlL/O
JqZ2EVHYBG2ojW68rtqMUpWYxUfJY6aMvnOjp1WoRt4vRueh1y5e/B3/PoJjSXSmzsBVw7hiZxsY
G4ItgwKENbCXnR7QWDv96UlZF8TLnzUqRu1yIDIoJT5jep0jGjVHxTaVNDeaAxsIyli51JCJGogc
xpI+CIr2384/ukkjVzvkPiNzzcDpWXkmhMs6b4p9s+/VeGZSaWfyqDloi1igUlsXHQeLsipLFspK
aLYHrh7RkCGJz9sZ7liUivIyBCtnNZcBqEzvUjIZOfuNMqmWj0S6euib7trELfh+6JqhTI9gM1ii
D1B1QwpuExR7/D8WNs5MLVphdH7EE2bb1tTLw8z2XWeCX7RhOcv2/CaFNIDZP7fD0Kq8hZGxdoNy
QnNO8ovwXgkxPv+xxrUCNrxPcdw0ZuyBCvCOs783q4wNkzqsQ0l6SEFo56Y+QacKpWlb1PrTH6pz
VcUqXuxsLarfCjzzfedQPXjuwdy+L8LCFaVnHlgRezy/084mZPTFwD0/BTUBqYAO2f84bsdsvf+q
HUU3+5nk4zly8Snjlts6X5ZAbtTui3EArX6H7MlfNhLgX5BVBcMHRnNC2YgV5+3i9iJ4UKdyof25
9nHxH0qAVdDLM7Y2LGGx8tBH2nyHq7xsud1TCOdXhfHC/YXUF5wd99NXmRBEHweniI99LtJtX7c4
bdwVWkv2BFKaGtZhkRQvFjyUnTaYtRz6wy6qeKG/3pEzpHkvP4WvdDVRppfFbysDgBVKNMKyW3hd
bKnXaXXL4IRX+w+hqfDteFtKBxKP5tW4YnYITwsQ7Tz0IwZke8cz0sJwM7hYLdx2d/H+W1g1Ixnl
UY93wf6ZGIGN8/UlY8kNC+sDiFKOi+aUf43uvDbRtjmfkqE3bo3be0C6T10nl++qjHwvMAJfGPBS
D/u3SEgAAzwJNbAe9fOsI/qLZuqObB0v3xZ4/WpjaxgbiQneYTXXKsILvfuuVt3S6m2JGBKdqVaP
dPp+lxFFxdI9jqlwYbu9FV1vYawXdR/gUqzbvR87phyqQAOffxR0qFxaBpbTyNjcrbLTjc9Vvl57
gdvm+i2MJ8GjWWirGjWetIVSVlsmjT4K9SEdRrj317DB9qcP9V4+X7O5B458Spy9ysXkIJB9v9oP
STfZ225YQYYX7pZ84XhQChgg24LfIbR6ZHL1Rhd3hORBRx9K7o/MgehaB7GMxt7I1H3L5ucQ6fZK
2kv1Obbj3uHRtNj+ODPzG1+Q9Qz9C9rMNWnMmDxrx/Fh7EmbolZ3ym1GVyDK6FCoepId7Vcsfjta
+Odyc1o+wkxt0PTFAPZ1/Uzhdv7BZcRggSRy3euobdiiNequsmXtP/nMfKLzqqQgIHUOzVB7a7H3
+fKFhUxp539QMfmVE2JF+DjxZk6GSbpU32kEgKFwrfnz+gmwhM+fdyaGwdDkN7Y3r71m77VL9vE9
7Hit3cUAETSXFBRMZrDVZ3/3mhyfXCcL+HiJE/QbjG8M4Que+S2FamqEaxxDbnPbA8ntd1vsfAVf
WJK+OhOaVVEBQBZErL6EDiqAjBjB9tvEWRoYIYAgSa9JwQ0JOO9AZ76XwHWXTda9f1Cksa7jjWTm
gHAp6lYD2ns8Js5Niz7teXwRs+jsbiwxzJoA0dKDX3ftPjha9SvhtIyAyz05fqznajpLok1MZ1WO
S9WjYLVKye5qc91GiYSl8FHBHID5rHAiXZXqBYJ0W7S27sUmKNpWkTNNUmu/OL6xQvaRCGCahH5t
4UZJFg5sbFHJ2Ug5xnr9dclp9e+aiQXgijU8JFg/dt/8bi9waQoT8GDo6CTNu5+MIVpVGE2rwPS9
Aj4iIGM+i8WX6SBZXsolcdO3zaLDcuk5AT8oHS/WcYaayNMcSWNgxRwA0G80p0RvxXekjCAfu/lX
+24M1F30WX0xeTfTuUwcs7XA4ViCiUDmhVrEp5Qv41H0elA2LeO1zhoeci0jxy+8UpWzrnPwnrjn
WLq9h7gWZ8sBL54ehrinA6lfGY2Elmtu54eP9qU6Tdjgx3BRFzb/JlSxvF5wVakrL3xQVhe2fK5i
biDUxFzA8aHtX4roiLwaDyqQcH02J5Dh1CRah6xaHSDNSMnnbh/eAJ4DBETwP7LUmzbVdKs/4nAv
ijXAVu2kYjKzFuymSG0W5yvLkc542mYTwvEN7C4kiagRRs31tZrJOTXHilts6A0kx2xNusaGbBZb
8/0ZrMcj8LY+TypVv/dpLicLODkCHGB0tJdQRLINqUEmwQxWW8azQYTpy59o/JYpFWvDheesUQHK
HBWxbhtjBBoMQHA4SKkMF1qvlZSFdY1vcz/yqTyVarpBK79gdYt3rWdGvNpKS3tprSAP5HUAyXoc
hypwzL+EralFG2xDNY8IEHHf73RXElSA3b2QENjOQcrxUohgytGLCB7bhAxyeA0LaGgFQmnNpEf5
SLoGtdGHjzPx4G82idzl6EGJxQd0+uy+Bc3kyum1bSThBZK9GrjpBn0VbyRtExb4HNaZQi0B4RZw
s6fpTqEBOqvLC68rgg+3SGEjswHOnrJF4mT6LgR821KWtcGFsczuA0kz+CJtxWC5bU69vQVDFqzp
74dgzXZ+YnlA+dcclP1I+PSL45CRjYYVA5IPRr7sh8JnIeUj7AFZ7maYSiDflF9i7BZanwMFEylH
htvrFrNCVjeVMirqXp2Fl/BmyE34wkHjOrnNaqbj1PpHL/FrJfa/InuSd+IjHIdUO1yBJYHENg7i
8aknQ+Y1HESqDqklraHTWFD7UJYzKW+W3DrxT38kBrqwEv2D6QTA9bqdm2io5RNFm99Xj+eIcpJi
Y3gX6a92G6O8ZZdLprkfRLHtSonakvoIzEWXPYsObmvTNoo+gi8P8oFxCSeJAyFpaKRCIxhPUpUv
3IU2puhlA1FYb/nN+JhW2WDONjs1ofqsXhvyoRb41qN3jJ5yqvA9WD5kX4737All+JyoWXC8SIej
/g/eTcDQbme0xP8mfxFIkSdQqcyiCs/ipYYaLQ1Ck4fY9zyL+g7nWkJTLn+ae6CD4kFPs7n67K27
EjR6ChuFmHPsLnDv3nQIccQc/eXA3DfJM9rugCwJ7P3wC6Bs11gPabiKJai1PHd3JRpQbgq8Ultl
qOmdx3ODRQAq3oE/6n1yncAgoqu13pIpcsaa4g46HCPRubClVnrwAHGH+Urd2IW8QoJCjkWzeO7b
pv9BB5khVXhw+mQrjGB6XIUGLEs2olep63uq5Ycu9PjqgZMXTc3VdkOYhnAfMvK6WQ6IzH8fWbJS
PL6zg0C0il+yM5r6M0yx7WYvWRzHNsF6JsDKlaqDcTESeql5g6Xwfz/ODCwcqZdAZPnenmv8okFa
6Lh0jfZSo6fuhfvM0aF5+mOvqsDs1j0nUgPfcZHWWRqP6B7C0+8+E0MiiQmLiIpNoOIJC8j+vNRj
MsIYQIn8vyaXPlRa6jTGUq+R2PP7B1L8WC+S/MWLL77AtAMIkKVQSdzim7NlPrzFb+veu8KEV4jN
ytog9xvKRiRstBdBQTGugmbIq+oLgXvpHdcGiY+fnACHjDGrIv26VO++xFS/4PACU2VV6ZUu9dX6
WQZkCD1mnApdkdQFuZ2F4b2QC7wDul3OXzaxUMNA9XSX7v9dJCpCKu+hRdqiQf82JghR8JvIpg0a
DlSUlwE0B4IrojZ8DQ1uUqFIWyfwfHxoMpvs2ZI/2Jx7yRbDb1sF8NwTBMNqmcyYZqFOiv3EG9fA
UrzpMqpKa2BplAF8Mz3PycJg3gQlCKJhbCUo7EeVpuo7P1Jz0EuT1gais/j5DzG+MZYVfEOL4JDQ
rGp3GgaEWqmzO/RWNtkrN3aaSlE6v20CD7AZuzfWWHiwqGj6gc3HfdYPwQag4zxvEZJ9+noV9NAb
E/FuTNxjBlkJFwvw9+snX0zinExT38CLJ9U7t+3V4G3UuV3sQ8OCMzi7WyXP0LPxqjWCTI3AsVCy
oVJHIThkEY0gPmAQ5HUeFwvkVM8VH8zcGNofrQXnqLupI3MqU9WWycses6OaZBc0mYefTOdxyOFO
Ux2wF6KBHhcTq2NPtrVy0Bs8l2aHdmvp0M7r015DFTDD5hKMoZiYHfy6K6dD63LE2396TjVn2wLm
piA9TdGMo6/7aEQsJpYC+L3fzsq4d2UI6YcKYTi1x7qwcM6kJ1VEVe0x7ZZnAihpvRNb2/kQFHaJ
t/zG+B7lG2RwopoLZ5rqg5zqW8k/pKFtsM3Ff+hOWcF8zd1181g4Tg1t1KuHzcYpjYNhRhlIWzOv
QO2siWifqoJJDLdfyFXSRjRq+tOZfEaNgzXdWSZ/k5hD5uG7ANsk6me1eUz1VeiFTCWq7nl0UUIk
u8cF7g9yJ3LuhiQsDNDQ+2zePBfjyR/evIV8sy8nISWdgYkCs4NeUcY1tMF2d9A4UsT0gwQGBIgH
8bGlICVwvPv/M3h9L2OVzsIKJxW0KOxc/u07qaoN3vN7brOJz50BqGKfWbuS4fKsg1J0bJ48Qzlo
VrwLnQDac169+8s6ije/rt64QjtcHtQW8XH0AYidd3zNTg74CZ18kjhHwAXsu+gjL+djHP5mKoID
Wsq2t1x6zaKRCGNuxfHdtiakqpnxeXXYKAUoytkzgw+0/TWCHvm7vB/oNn1rIvgrfcxg05Ay1tgM
ulxBQGfv/21faoa6q5U+71v4T8eaz+EnJl5D8qpU028JubjB/3Nfo7dle7b0uvnWInpM2tllYBGM
AgWEDMQat0SsJyB43z791BjqFceHvAF+1f1+NwO4jV03BnLNVPReRFDWf6ZtWA6e5y2wC6uVTqd2
sJW5hQaEXtq3jMFDpTHZJyO1pBZUVLIorvyGjzJViF5AyVdSz+5YoAV/luKt9EO7U99g6upEOZQ9
UezUSqurdSljoxY0Z6xNbH6qpKjeg3Y8x3bPQPaxg62j6LVcKt3lubYE57kiGqHmdm++PDKAUEF7
d2aqTXIuvrQ16dcvk4gDksH6mQhQJQKB94rCQqJem89skmN2Y0ewops6j+TZPErErNXSof1ozqng
xzkkTf35jxy0Ag0yhRW3N1wMbDuxbd0lQkQp/iEAmcCWw85oeBLdZ1iAeW4QeeTrmv/x7qP9STaR
WI4HQ65Vdabv6ikBu7/MpRTN6aV+cmInChMe59VH4VjdzOis8m7s3HSGAJpUTW6/55hGu8SaqaCY
WpvrIeqoMLZFAsMk6GwbIF0MV+ihzsqAS3LYnGct7brvZG0KddeegBPbk6+GZyX4U5iUScZLqQ8o
18lP5i8B8CiMxPtZspNHL+FJUZifbFqWXW/HiU7yuLeMBbmUvVA4IF4PIxuwFP81nMKflkakifIR
eWSJKVOf4S3PDhMep2mbgsSk1T3mEs5pTeAb0APX859OABuzwnJc8oNojMoUfowdUvQL07MXufFe
j/b75P2WmWoq8PbuUxX6TXEXqyNGn59UjmT3fLo4qtViDciG4mx4HzlqPwpwDfcffUCyHCak7ig/
8qU25GoSQN4NJA8hM8t/bhFf7CKtYgJE9WJqKjQmE9VKgBTEa7DZwsynYlAsGZsQsFK08W7R9K8p
fhX+x9RF2qdV7/zVNeLj2JuDh7U5IyYlh2D/hU+q1PEYqwWH7sNEibcPflxRqhO9RgwVSK2FDyRH
D9dnEnCAiGLlwqhsVC99T/NUYVf2y5pDYCJjlmqv92GnJ1t+/T2NqimJ87PIx5lSGwYUMZ8OmUmQ
ZwScOpNK5DeAweiKjfhxIvWvDP5wYZUWje/q2KBI/hjX8gMt8LzG60kPidfDRJlejS15Ac/PCAUZ
wKFEjLlzL6cqOKllDiGUhVYymWT8dY/FPYYdJcjV2iWXapMxZQaEGb+oE7+e6q0K398YvjbR1DBb
VItQAu4+oqhO+0SRHx+LJ3yg0IXqJZ/TeP1qNg1IlXb/++bZPPRK8mWRPaNyV+a7jZh7K0G7pJEQ
nBeDAHGukvu4sUOTIC/Da7sRw4aRqrwMAFzw9UO7wzlGfW7BQAj/aNT49kMBXa1+EtKhekS2gruZ
o5M53KGzdtf8zyoSk9ez5hMjEIoonHKC2ZoEDEnUiE5V9xGV609KZTYs4HdT3KhxCafoj4GBDupI
mLFv+fXt0K8oRgQzv9L5Ac81Ky2GVtWGYVbtBEywHCQ2Usq4+kiRIqYm4ctwl0gCSn1S6QI70Qzw
+piid2bNp2x0SeSRs5ahxOrYDPomX9FFIY6oL94FHR8nVYVbaHXyu6sj3cicQdkw9hQJsEfAEorO
eOQTAHYTipbO1y/mio0z8tevP+ZWP2uRvfyMcykmUDJRNyyTq+ll+lqW5HO9x+664/ScHTuRwxkd
kftOi3anbkpM0b2eeTpti5LOlR5BdK/oQ1O9f0cIBMkLXVxivqDW/dTSsTTKHfvIwfYQybluUhte
zWEo9bTOwgAxlYWaA/AIYLnAsABHuBzP5gEJNuppcHArlAIAxOvoSvacB3c9AjBSU1TZvBxto6Fr
KCYPzGrrIGdBQ1wr3K5FDsPJK8aSGFho2WYbMqEh/hr80NNbPeWqCVpaZN2Ae58I3ujN4xAYFXHz
oEKOUvmQq6iwdZrQDaIhoNf8vY7pZRS8+Jejf868DfQKv8BRZNgOHARRrvi2mGpkUyb2b+qkr7vI
ZlSClSryCOd2suU8hKaRHo1B1UD58MhuY8Hhd/vx0ynj9h6eADpLH/9U0jAhqJOfRXknmlT3rElN
kTolHounA/8FuBqxXdnP5xkRKnO6xGBkJxa79vkaYCACWfSIL0lXTCAlSasE7vvIxo7CRJBaEqec
8aGyJ1qWoCGGX2QhZnSbzdNNaymluhKny6rdpjqJ/xLptXNBAHC9gi7zGUkRB7w7cYc45dsQP48w
mMfFmXFJrDZxZYX6tIaNB/Lw7Ar3aO8R3dvQkj0Z1rQP2V20mukX9ViQUw6BBf3H1N3mRrxFGgq6
HXDIDMf2Wph8QtkpPh2D4eHn8WXUvYaIHIU2tWHM67quaLM7XP6zMhnHAvp/yUVcQxprkjervXxI
ikji3Qd5QfSfxydhX96SRiPGR19DFbUJNdk8WXchATGJMxvdaBgw7gDtJvMgJIiPfhh0Zj5AVBsg
vMO7GvLkDDqWgLNhZSuF1znv9kSuNawEljIbdYZdpGOmSbO7WDoDEOM0cAnTlerbTCfPHMDmgx55
kfroAIwrlISk2Cma5GfOlXcvGffcr1gq5gYxczegEKkpv/UVQG6gllaDWXaSAA4ybSWW9b4cDCWv
pS/Hx4CKiu/j7t26adbJ5Q3GVq0O3yZW+fH7MhVuYwDZsdS0UO3403+2nz6EKzA20XY8/CKWbqHP
BEDj8s/DhvLl7oD3k68hJDRSfhNxq0bO7vrKNDOUlPGnBKOCjEMvlsT/Tcowlgm0QYxNGtv/QJ+W
Xbqa5076E995pU008trTKAd36VNmBK/KWAGyUpcHcjTOxCZRDem59Ld4ZrVEbV0FCvDDpA/v/BaK
zN3CbmozHERTdaKZwz5cWOt+oBW29WkmpPQ9980gtsFBSJHkmdKL/QqgH79L0JQ3moa6WFMouLyB
/C1W3jSjwY3kDB9NHW4Ina60IeESIAVB9ge3twNGEBORwZigbR6vFaiPbVDa1cxZXQa0gcGNzOVW
yxRrf+Q1vzFts3gb8KoYbeHYadzOMw3zZ36m0XLVJ1TSD0rlJO+AT3gvpElwTBFLywHoWSmAEckz
TEOD9972F9tDqp1inRNY1RiqshbtU9Xy8IVzM6ZyNYg+pK6YljKYw/oNwanN6OT7Wl+OudaUUcJw
ClBwlS55/h09BnGG/rgBQ3lA/w+MF0ZYO3BTbFhwmXLSWeS713U8JB4XqEvHPTxtD1XjVo3xxi1w
L5B/x0YUEd/IxDoWt2Fd/DPablWsADVNRHZHg9wO4r6QUd6GaPO2dd0fdraEcyk46AFhm2y8XCUd
ZbWE0Kq5ykWvsybUdmL2Z5sLZWxmq0z0+xVvniDIZz8Pzs2QO5a1tA9MjAqI85v6klvcbCWsDs3f
e34FN8djrbkFAJBBOi75qs68TSOzO/wA3z4U7LFQE4K2mxbQh+0nH8Vg7U1pGCVRcW2TkVG2JdHm
f+YNVFMqlBudQvXiOcI6253AMKBXytkfEGT05ukdw7uYqudDKIky+9boR/FY+cL4RZZIIZR95cJu
bHjETxLiFL91Qm/5lNeVQ/tszWUs7u5YTTQUsDtlt84BX3+RyQFI5mzCKUusMrBAjq6LFN1ADpam
M8i7xHy/uta9b543ucuOfx0jKfhpE/8YKl/nkoFhMaWKXtJCUn++F6OiWhxUshDDIGCQGVDcQgTI
g8vomvNEkCugbL9QqciwRTC1uw6QsZY9IY8j4nqG0quhvAT2vIJx5FhmDUPkmoThkAotZZ5XwuOb
8OgGHX2jrzGcdGyfw8h3uh3bp307EamTxWUSy0mvZyxQinAbmfESo5Oi4CMHyj0X4TMoHSPWvXZA
FCaufZmEbLulAAysaCCoMqWiFgEGIi9Bp+KgPuKdndNv39S7K8cVmK6v4SaY+X/EOWYIFxtX00Fz
hog1cW8CZbn6BMYmfkAM3wZEqBDqNHlmxnCFFQwxC4SBsdpLLyKgPGA9kXiSvzzsUnxbf6C7aZHU
z+I2+Y9uSLp8u8cJMFk+JA42N3W7godfyP8K9uKyjXPqpwWLome/23F2A12+CsMaCK541ARJwtni
QZejwDQ0Tmd1I3Q+16X/T2yA9nAUi7DQXEipCMHse6rEzVGzddAXd6xm+hRoxCiaMT7Ab3yyAr76
w5TTsckT+dEfsP9+E0/9i/rwL7BNx6I0Y+dynqYhnu8+4sy9akkAH+g0++UQXx2UjLKW4yFjRis8
l196311I0KGhR87zSExKyi7XWtLSt+BbRleuNhZQH4Nqtq/CPgBlFJnXUDs746CILUXL8XZwzvhY
etea80KtHJ3C2CbPP7UTtpJgOCYyDd7yV5hs4N06G0wZOOaS4G0G1oBCRwtwZ/Myjt8tyDrNru5c
fJIFWYfz3X46YC9EHD60y66hFvsr9qhvhWoBlH2prF4dDu3YGX4OKwDLX7dinvIFtqG7pWoTJHQ1
23qIW51y066yf0NvSnCUBxyJNXLEDFe7wijAty8QHm/CdQUu2iPn6XY6vhNWUdmnIokvJbizlV7u
7mYR1QZXNX3RIzyZNG3p9PJKRsofIMTAdwqcIypjMO8f2Cphh647c7h0qgB8IEojnZelK/2QPka9
rCAkbBnYRlDL9Bvi0VPPGcE/M3vO9UthASfoKa64xlTfa43ohSduMmZw75vDpkJIKNUwpYIZr16r
/1YOqeDbRdQPvypYxwZr6l7jzXSzX26Uk5SLxAMUMyDMaL4Go4QHxo8wQLZFVUNp5ApExNXBWSOr
sYpyGXv9x5fyn4kmS8EtPR2JRbKMrfDsJ1o+8SromDrTiJY8gyJZxvGAs97NSaabGd0F8zMQce1G
+1deBkkQzGeBa/17glFRLqbMA0Mafvf2bSFyI1IlnyR/TV1KRn8VeQdaF0e3HiHBzPV4avfAzDBg
KSUv4vqm0Nlv3DF/qiXFM7AgXdpfOnHy+alHwPdio+s1l0DXwH8cesYWk08bWbp1S7VP1ZKBq6SF
wpuKcKuw+KO1R5eiRzelIBNsQyiOv2SR/Bo3iyoVJJcPHDHV42mKanqyTtZFnRYwZ4JPKDYQCWuD
FwNPCtDnINFvZNeshitoachrBLpMfTCspvrLCxp5tGnpwUMm+mmclCkFCu6MfKDwwLy6hNpYSev4
8RnGIew/mQzvQIbf4YWRbxkdgWhmJwYnaULF9T44GEqtxcu194SkcVEbiS9JHSgfK2WwIvH8ga7k
ptugRPtxcD4KYSdP6Wi445AYTWI2vWpIwY95phBWUTnX5ScBzcSlBDn262zigFKcxtBdP6BTgg4p
5NH0LOFG12BMLHjF4GgKJbLo6XzGC7io6JFEMpv11HrqbaBSwlpuZjNXmE75fw10WQoFX4A4mYfA
8xNA7cf59Psod/LkJ4UrQpnqwmQvtD8BHVYc/PsudLIDnlJmJP1IHhrk67ryMDI/79u+GGX1rrAI
tPLYrmUNVX+jS5TMdaR0JbcpNv4Q9vKWw0h5p3t/V4lQNJeb1tdbBlRDlHszmLjBOqLzK3KbfF0k
PeqYZPPC2VkXOaxzOFLqU6sBTfgmujkzfE+C0qil+EnnTRiz0x6Aokbz5cwa2qtAaQesQu/cxri5
vsQ7wmuLPceoxhmK/iH8uByORYprmuYUsgW906gL/+73ffr6trJv8gk3/zUEm9FWdnye7fm640cj
7Ys+HyBrM3DVBkAuqXxgTSkZ7LH8KtGHz7nHEbG86gSAW34+gsUxRS/qTrAO01DGOanKp6NYgysZ
uFFlsuVbnuJ/ifEMkPyPCmi41XpKX5e9stRN2CLqmkeiUKzjElNw1FaL9KPS982G9eNJdKJdYT9o
C0Y4B3VOArmtK9XoE3R5Uo71WQG4ghM8XI6EXh1x+wCbv5fb1gTTPoANz/3wX6+CAv7yKCuwTjdJ
rGAT6Tgxj9zidVgFY5PfwDNMJtuqqnNIOb7A+g73PUifFikguxO54iZgF13VfObzsLLLpkuneyfb
265QB//25t5M0ch9wDtSD4M0cTreWrFrHqLRoeDd+hLgSL9/kcgq0J7daW+uBYpU3KNYR8xFxT/5
xERGHBlr0nDoX0Zp6qWQ2hgmksTWw2V96QUimiRP9VAxtapmZak1/RxtFgyW4FMpKprU42+JTU9q
tgYI8tJBev7RiwA50dJeQHl0J9leGER1qK/tIHMwwa/bAcPgiRhLyHjUGfuDEck2UxsB0DCsmsdw
mlnSbMeDlxsioZ8l74g6H+pypQD7xIEJrgTW7K5fvSNDl2CKtJNbvLxApQhDVzNpGfapX1gIxbWs
Lruw6JcgZ7Ij3U6k4202oT191S2KI1j6yWGaTmbkNflet/Y7tnZreGOmO+yG2UbrJcGVFBtRKmQW
6SM/6jWj2ElY+cZAKkAiXeRPeGUCzcs+5ahCI5vbFXAMT6Im+C7mnlICh2h2jflKiFEkhYmrkCoW
nVImON+uKY2PiZdMtYq4A4pN4WZMI8vJf4W8fdPTV8YLDrYoFpSf26Sg0tIMSY+Ro+DMNU+GLj07
fthw4JDSYCi/seqKSINJmx5Cel2pb+NkN1yWnmugqkWJiv9T5MZolUshHIRjr1PU+IG5QU8O1Hl7
9Hz5GbCRh1lr0WU3aOeiPy9NUvRQKfmHbDZhihf4WCa9Hkr0TdpNx1ItuAm55CnvEubeamOJP2LT
waB99nMS+3i5uNyMA+KOB/XQvgLGqVeESZu+K/MWDP81bbBeRklzUqioaK0MDpMDn7+b7SHNocJM
BK+gtaUizK2R2dKYgu/OlmyVmV0bZkShY1Pb8lCuzhrM0YfC9rwKv54NgyE5g1WO05Jrnj94yFJY
1Rr+ohai3IfEjQ6Hxa4UWvVIsvbVo67bb3mcMCvjeiwhtuVsyGLkdQ2d3gMG9utDs7uImHae8Cj6
f+gweYCXXVyt6ICojzDG4cVfnjACpU5GIAjUeGBFCww1DwYq93oA2W0HMaejAPEZb6XYZLb91Jln
dnP5O3Y9z2iEv+bnEFO+0sY03n+iBpo2+D7PRAG18NAMlEbpb4hMmGGtPMMs0huEtCUySyKu6eCM
iwRx1SzFjECkCRE71D+z6e7UBriya+bTAswT5CswpawWhDE8AuxYjtfr1Gvu9Wpkkq2EeAr1X+uy
weM2UiNWoV/FDr0/CdCP8byvY6XevoG83atOBC2xDYsWw01coIdTgUynGKQpDf/YXUpYTuy0cQOO
J6+kDLxGptpVa26Q/BpLekJZP3ZiSit6+1365US9+FjQ5D8FC+meMXnor5zsHRcNgGZse3j9Ow7/
RBScRgvkEU+KyS+rTLDA/CUC3VXXdOACozwQ6sXjtevA7sywJ+Hd1uwyaXjWIsv5QsmchkwrjnrX
nAvSjSP53GYdp0FGhrFZ0CrtKVcKxUGkRiuCIqaUh+Izr2UCDiyeM6qpK/vI6ZnyCrU/hxWIsiRe
G+RRr3nNAecCdVjTLy23btE17YzBuj6XPp4zKH5QpgzKeT6QbrccrVvuOsBwUnAl1PcKp5X2IeMv
TTiIwqyaSn4x4x7gH8fg0ehgBa/WgfxALuv8R2xnst3MNxdDoZwxG+18HI3UyCPADXehlFvkeeqt
yH/92+5Bwg4POx7frexDz17jLi6CEyC4kGbKjFu9u9HQTrEU9N0GQkX25vv+7aeaeJY3o+aCXOpU
5TUGmqEJ7ei8FtIOPF2g0aNEyPTNH5RjymBHcc0oJXsAqAJSOWroHEhKBc5NYI3gKvFeacUxOVsc
GnC+/1+R4FjvWD8EXYbBjGlWVlm9Xn+egr3WI6V4WWqFAuEKQVCLWAsnjZC5SjB9onJNHeH0iZJV
FWY0wVKjBE9zH+Iu/C3fppdswAzvQaODTxFGbeVg4sn/8/eJe1Ihiy7JcbHqMKx2oTFd05aKV06C
T3NWg6UwOfGshLDU636HY8CtfagczPLbwNJzdOSJJKkZTDcUfV1uzBH+EWhyTrZcN/QUsUlpVahS
AzNx7PG7hhBz2xABtY7n8jVdluh43jRY/EDa2CFF/MYANyBgbBbnxkfk7utz1l2RBC2+YDMR6Jna
GI6Ejv/XlVfNDDnOJmvNMI+rfgWK2EYG2nR5XkFK/xhaEDG//3UWX/H9m2UXac/cMWkgU6owevqW
tA6v5/SDg5CN6bgCsYsS4IbMxNXTw89Ue1et+dbcNFdgsDRF8nSNhjWZZSU9MqZ6Dn++JeGa3cLM
ITp84N/JIsK+JhAOsXQ9G3LwRktWcgiYWuDGouOZnVifOGuqevSMe0/a8e6D/vzV9f88N4pfCZQi
LiCC/pNpuy24+yiw8sfkrrdlvOXTkwJEdpfjtdeUZMcjr4RmwBdI++CWxkvP6fSyfeIyztlYppIO
nGlZaqsjgE+cbafyEv+DB/ba45e5Rkyi6Hj4xfcT4YFwz3OtTNZEc2qMduL7Z9LmhuMxzWFmv81Q
8qHWUaZnpDY9i9006kI4cws5J8hEp9z4n2zQgABqAvrbtxggzki8zFg8ZlWi+THwXRfRRi0gpG6a
TAYbYUV3wxlSuQ0PUdnyqCz+CGoLdHEx7xbvwus6NoOTwmfE/vLmbuXZKZbRPa1kHKNET8hqOt3s
w0ftgAErGJPgOKvChvgpR1WBvjftDpszy1ixRDw3NszZCJjqy01pB1e1v83D7GE7VTbXmfNEbjaU
kR/b2IdqOhohSHwFAuQzClVUYRvMlPHQpZ0rZvtLSoyrJHY5vKx6QJItRF8ZdLIHO1O3Kyc24py+
nLWVgHi5Q1F0CQmw8B98B9hdLAZBvgABSBntgovvORnhF7txGGbqPeXA/KT4MR0kV8mBxmFHuEIy
ktH4HSb/y6KqxFK61eTJ4gA8MEWII1SjtB99lbPlGIOSssXgUh58T/EsJ2bFQFJiciy1N/cyKh/k
OXwmEIAxAygHLtfRwxmafXCkP6kLMEyuXGGC79stOf/xZMA8sYnYPUsjR9GhM1uZmeCEq09CwCoy
8fc/Zko8L1KaN/7lPXoy5TFNqYenkvWtCKcCmfwtbz+9RAvgTPOn1SNP7puHA9Hass6zvMpkhg9D
gyixdL8+l/g+CCy8G22vco3cFFcVmKWW3P9cV1iE44SgdfBK7Uro7WfQSG/hvswwmsnB1Zsk8xF1
z0POoyntpv5kow2tyGZy6UiQw8CT4pMLcQKqLdYXs+IuZGyZBdOOsS1qQffOJD7IbLGHBgjdtl+1
HnbXxHC2JQ0ncaC5MOW/nM7KETG9hIQyyEu6iGZnnmjvg2D4tgOpvD7yKGH7kQHz67HyaPssljcZ
IEtWGrH8RYD+3oxI9Q++tWjcymXPbSlDTcyRtJfqHSVmCIONFLPk7H7H3Krz1AID9/32nUx+jagX
kmyCSipI4lWDO23/Nqn/26TWY/SoeMBfzMGR7II8HkJJ2L+b5k7VizOsbshDFoNd5y8TZ6wm3o8g
nurZ7JLQmxCvNrn3F8vqbtzlFrBj8MctNBS+PNlcuwYwvBl1PwyZO89Tt6pNqoTnR9k2MyBgENCT
TVRScFRAqf77F+3OyINQsVgXudhYC2KNLl4V8Gh3h59grl2s2O/ChgWFA1QoprZM0SwPS13jY+6P
A2/qgUr7KkYW2sIO+D2fAnOOE5/uVOD2L2N9lIiyNQLdM/v/rbWtbwoLImjmZ6JdE05OaVMSesQc
zXe8ZZteJk1/Y7omXuzOoxHYL9wd6pOHGlCQxqwwsmBtajeazSLvuUQSAVRxG+i60l/OSh4/Ptfx
/riuEuE0VQFqKLyk6dQ4QiF759t2piO9lkwKoc6qJF2YC5qU4bp25R54+3jJAPFaDSr3M9adMVvR
TubD2kYDnX4ZSFXG+SvMCC+GPDQpvjgI2bB50iuoXm3zWysXo2dXgZI6HN4ZlH0sBMYJIo7eFeyH
368/xqDBCkXTsweVyVsaPsJvYFppAOKxMPQ708hQUqVx3Dl4EttunOsvN9uYnOQ5RbSRUGI7whNf
tdXakqL0cs+tO/9EGGM0967XQFdeZsUDwMPQIVUSzodVC4USnCo0aQ/Fek4TfYaIcggUo+nPUUHY
YIdlEO2mDF7fDeC6ak+cig0M3x1BQjr+l2VHNa3DpXuEQ62AcXjfZj4LMtYH0AMT1z9QASnZr+24
hXPgd2aqGccGr0MTHB2GoGGoPFD7L5IklayEud55PWR5u23NQejidGkSqh5XTUlqqO9X6v2FO7D8
628PP7wxFXeVAUxKMOCO+VmJQnNlTgq04Iu0915g6vYOKapicU769GjS7k1zvynUshCo5MpGI6pt
sPqpEmKodKWr4lkLgBMQYKEpr1lECCWc/r+D5eduqF3S7275gm3QCNQrjrohv8XK3Bl/dDXn7/Jh
JHiD/x1u7heYDvffXMOKtlFqzAmRmZaWDGfO4vs9Tv4SSDn31QppjnDwP6W6gug/PR283cwtqAnN
N13Hqc2suJ0AXRZqt3qPQxWuZoO7yGA+/Q8vDnt3wH3T378BfvRlmGmos8x+ihb8eR9DItENn5Pj
7BkcevTGZEAd67lvN/PKWsW1NnzlzTdWGLKzJ30Bs/yimqq4r/2lwQT6XxVpYvavIBQWQLWvbD+b
XCLDKGlF6b9GuZcOHjnu4Qz/UoHrOcyVpgqt4gcg8Zoqpdj38LlPVxvmurXlGIPufW+t9ykMGCUd
rKNfjDQSCa+TgyLGB3nZX0kiuMi7SmAHG+9gABhI+TJqKQP4NG2nMaonPiEFF+z7YeDOuH5FEUo+
Tmvbg03DxJnqzt0ptdJ971BxfNLRZ+dLlhUKO0E2G3qxu/cpwLv25/K0hJIlRi0gFiuWP0BZo0EQ
TGNJdfuzA4ZYpYXHSJHgFDEH40i5W/pwWMwt5x6eyAZuV2WaoyWj7ouhGZWgkh5NJEN5YY47k2m5
DNZPocLuQ0w3z4Y72255fdylv1atGRIRa7UF4w/Z3t6W3j2jMHtZXtBMwzlT65GQNRgA+DBtJ++p
BERHDgZvmHymZg+APjvSlfotilkyoRDQOUAxGOo4yDwl4+92qN4OYHa3jlmXQ0RrBJcyLfBIlUNq
eg/8wyJ4yJW50G9yp0KB9xTaeWJy4yEqCFG0O6aCka9sYFuolExCbJ7X0JJNSokCDpo1lWC7vPaI
8VTBHWoMK7OoMGeAK7BLFS5aQL4RoZJB0l9IwnIuKNC1qIsTVNhwBEHzJyrShMjNUty7lx0IBv3e
YJKuqijisKZvNL8ge6N7qONo7dIpvwyGkmQE+s5Mato/ORtX4kSndMGhhhAeJbZT+G5G53SyKtSR
vLqx2PDTWI3qzNl6IGup/3Q/QMCJINAkp/dZYRwtZjfuRSxl2mZQXFx1el98xkzput0wv0MTJiPz
c8PC41LH4202tYYIwi+vepkRdOnJFrBW16oYMRSbwdyPuopMCCDPKRa6Ba2jj+ickusKks1Nwv47
QiRCIMQ7rBJwH6eUNUJyyZb59H1j+eN/OpBdSZUPLvXzDQSiKIKBd4fI7olnGHWG3VzpokxJ/TMo
e2YKep38apt+i0Oi+bseuZoxNlKOhhoY8WJKdKGMSy4o8ZATVuosnYMjtfpo4myf9ok4HmTrEyb5
4RXPjU05mFlPZzDdqI2CYCm70YDoyJ3ixVCFXTQ0wRWCAsRPlnZ6SzQwXNf9QRv8zN+xeN9ZbSqP
+OczrdSu5z2tgtnGKDeqr+vXSrxIeVBTXCB1s1iSNDaWL7ahrUKC+jD7NRrRWERpN0fdjJKUEDHy
t4BuAor1BoFsLoU2iCiSF92/hiLR1oLquC5Q8yb8H35zqK57jkhMNdoedDS5ENVYqXzlCohq5uv1
O3Xy0ZHYFkYvLmQYEhD3N9x3+HxYHX2Ckur72cLDNq5FavGOAxtutUOs4uA0hzuf+XH6FhVg5kxl
k+Su81KcXeAMvkAa3pSJC1cHyc+eIVdTnK+X4gqHm4VsXWCpAhv+/yJU7ym3jkY284OQLIjTQ+fe
zZV7TYp0kyCEfTA3Oug7te+TBk+dFNQ+ZdMlRC2xlGUkBiKe6ht0y3unzeyHvh9YrMklQvCoQvRn
F5q/QDSwhKcVpdTCD5qaxajo6Vf8VmIrKr2fmSR3Jx3AHvKZBMqamcSJCUxXpMhWAhF/tNJz4z4v
G04X/xHfIhTdJfss7oC9j5b/joVMVXjGQA+PB5+xXg5tcfFc7BLmCtzEooQGyTvcB3T4+HjZeRGQ
hSGiPknF3xns17ec6LV7BLvTYnFn3DNut8RacKKOmnHJu4suUWgXTGitH2pEwToi+WUs3zQHj5I1
uhaRTUQ2bV4LiInhwJD6c+yuumfhr3FC6LPaLpoHYpDt8bvGpTbo1Poo/gS9lGLtZzOOWFTfm7Dz
mZwlsjTdTPMnf+chdC2KMjyQ2h/3b/ZV2UFvn3+5xapPuUxPPY3DlR864KKdEpWISMeDzc40MljI
ytpl1ho0RUoal5Vh9VK7I9IXOcjWmILHHP8whAOjja3iU3T1MgOpEU3D+waFLxdZlf0VvfK5Lkc6
YKTkQ1CPimL8gAITZqCmE0kLoQ0RIJqxdFVgtmGm1tzyzcgHagPDeaN+TRjvZSe45NQRTQ5FTy1b
WiQu8gMN5r8HwwWH/xn2JZtYdxIlVN4CvqHogl56w/VBK337twOeyblgQ4hCI3IWX5bTAho/MMek
p3TFiUfR352CJmu1/Evga8KFj+TB2BxR9kjwu5XjidL+smOjWDGbcrxY6wt4cphUfPJZpandSnkK
zcEWamDTWIh29a5vMh//+9CFj3ngt49OPOri7AlVFuPnwNwYwZrdTXM6fcVVSry3Q5b17UJRMPgL
AHF58sNPwBYT/AGeDSwsYyXPmxAa6TxJecBLK4h5j07I+rN1QXCQoZagUWA/YnBn87geoLCtge9l
FsrbYceBRZXRMmiUBajI4prqbyDLKiunSnErdc4bJKIrsScWVaFAsgh+yHCcvMs2FHmNvY9Pkt7o
rags1HbpuSYDHYXUWJXYuCWr+lykmMEQfambr0tQfq1neFarPghMHMg772wpkUA6GK/GAvjEqlrs
TLTJ0ptzSEtnJ0pto51Gn9fr5VFRWQ4yoXcp80WRx3RCHT+wVwKCr8WzKDw7eKd1N8o+EFmDtHfb
MB+pE2nJGYBywyXFW/gwPu9DjQF2Sut3tODz+kQ5sHlzn7vy67Ib6WhnDyIwuacMH5qvKSGlNug0
HzgpG+tBnXw0k5/Aw8SH0AfZ2MY12MtjcNfTkz4VH1hw0LicE8+RyK9/3wjYNUnRsUvexHhPaQG5
640+f+UNezA7WWpDnZ5ss3M4HZ6Hwl0ihb/RAPa7NUL/vT/Ik20D/uLLwSzehX0SCisryx8EVjsc
3OSw5XWtnOrWu9uwRIfVO0trlwzkwcdfVrHoUkkTiGvbuhKXmYF8aJeUMo4tbPl3++Wjfu2ZyfH7
NHlhA5HsCIPOvSgCp4Ki5aXDv+2M5gUYeYE7kfH1C7Yg9wBJXQOKe6udpoMt1L28cIl4Vi1wX+Vs
sJSzYKMonUVw8O8iIz9gi5rsoBZzvLfYWlpTSux0u72l8DuaQEDFTOa4jVCOqSIYk+71ry+BoHKF
rjfzbPMU6Pm2ypt2/rkvv7jxBl+2HuU2MT07RvbLAPJPF58+GV5IbDrt7tl+qhRKvYkRE53RF14g
GbDSTlVXZYvafI5oTD6Ior30Rn15KK9zJ0gymM+gwmAeW1BTCn1b8iPiaY2duIuqDnya35m00EcI
847p5wRNQW52C/QMHykJ8eineZ2anM1na+I213BpyrJMmgbEKtlvy8Rx5tpWIOYaO97qddF/YaVY
Ib2Ag1b0ThAtvyAYwdTVNbz6Pt5LMVacQ7rQXMFHujccUhwfUq7xZZs0j/t3dC7YOT8mr84dh1ei
H8yQ8NGIJLjUxzLsDlpwdY7Vqwv3F2dLVucUCfOWyRa8dTFkd+qSxkLQNaiAMollfAr6f8cu6w/y
B76SHrbVp7pnkG5VtUitBKvHR5kLwXuNCuqGXRAFnLguga+R8OypjVaVxAhAIFSVY33aqkfJvJk/
22toUGjd3To9xz2zY/R9ReJDiKGiTqTPe07ReUrJY2NSzctQ1bEnKSPcv9BN6EBqjswRrBZq7Mpp
mLdsMUmX4CkINnCH97dWrmrtRVkeESw7w3wTWdggVbUuV4SaZbVKMTDwWyBhOsUPpO9V945PiStG
VltKpyY3XGMz9J21D3c8kW/PpqpKyUCAfsmErIOqK4WgxMHGmU1pttDg5roLFxk5CpvJWGGniNrM
x5vSOIW+qmFjg6jLs3ALTxYPbQ4qbB+3rglHPBLaLI0dwcgr56/pxS4KTaaqiTQHrFZ9/hH1Bc7c
v5TNWrrB8UT6hRnTZpD3sU4HwN6jRJf0+AMQs/7neUWjTZcHJI2OqgsmTGmfOI2j+5WHGX9SGIoR
D3YckYMgfuGU7h3vVxtcPHcs71v39PaP26hbustmhxMY0rqeskWfdmarVF8x04DpyjUMSxq33gju
vD0EJDUYLM+LW2Q8D518ZF1wivj/R/yi6Vc/8NEHw0Vha2A06oTj1MxgZTtOWZ0B0EfjydMhHDVj
7YhNHgDYbIqKeDDUwSG9011rAosWb9pUPoaqNXjpw60jNc6lVkWEIwViEOZk6qFtcsgO1kV/X9ma
4CNjxJVlvt3pGWHZGePNtb6kWVigt+XKDLO5/VPxwOvmQiSd1yEYxb9i4bcV5otEl2c3MeEZH74A
0EHSmvjM7BOPaqPEXpx2ydvMy9USeQi9CixRpZNqGCH5dbqeQmmFIVEYPP0zJD0UitpKsD+uQm2f
1lpg5gkLBxpidaLyMCD7EJDSw0jmmkrg1GCmeUi7Ggqzd++J/OgL+oDq2eZJ80K47eWD8CH49k7+
j6ZvZ3R2BQX5Yv7nVTK7lxSDurNJmhQv1tRv87Iz9QrA1FXytS7/ODEP/aTPVp9YJCchVB0FW1+1
K8SUEUA6I5Osa05cm5ZWvinF5rJuR85yf8n/pr9AsfoADPTKZq83AOOHmU3r+sC8gDvk7JiEimPP
XMgd37s1Ofi26tA7dOQYC45it2JNUzFWjSnk8MKLL2O4w2OI51oBhFhQQ09YUMnfaLDg1hedlkg+
DUtXh8YXk8T6ZO9b92xRthzuhB5LlgZSE+2YDwSH72MObVSmLxvjIW5DIUqXhBQfmXZrZ6+YppU0
hGLQzxRtXWxQjlXzMFGVorxaooueGHyODfQq9yJx9PerTVTTvQDWhpOJsNq3Mt04tyyLDCKxsHTM
uOCWNVUX4nByk+RahR15ao/aaS5ZVEWiSgvS5sL4ZJLEIXJMOt1fAdIB3z5wdALTK0i4ul3dLTuD
YpHWqAL+sQhbCHinnSJUv7Mzpk/7cV/HqTkLTafg4XFL6XgJzJxbN3QRQGBwmqouVTAxEWYHjDFo
mYIIGs8x2dpr0udSCaJ/B8PzHDLtmHB6t7X9DlgnLfRmIpMVReSKy1i6dSB0go5VQa50q4pRRIJl
xMJjz2YoMsiCxNLvykVOjdny2nbIUn4Q+UztWwrlcu0XTolZfY7WXUVTKxmv5Gz6p/wucTQ3g2Db
j8IFxQsOi1qwPQQZWQmDBc7k6eG4v8I1Ix17DiWIjWEDByk98ScK5lemf3+kT7hCQTRnbIF3nvAY
znesA5wU908cb6zw63U5GSgeXZH/Ae66YyMeEE+iossQLn/s2ajPaaXzqVCvomN8e2PU9y6YpguY
CUC83kYTBKnGpgwWtBLF9QqBHcTLdhoN8q5BqLy19NfwYZZYkZ608r3uaA8mr6xKj3lHtiURWZGL
5Cmutwk3zIxr4Hd4LaSmsGt1eXOTu2gTgCj7kuu6TfL/c/wDRwk0SCpFHzseNCT26v4v9V3nWsXd
ZtcC4oRXtzhhVDKQf1R1YQEVKk5aeIfWmjEk6XXG3I6I1yt20+yH0psISYiQ8l5pDQ9nOfVfIs81
odJD/4A73ZvW3q8NSmuTxyWlzD7ePcYyTn/RUZew2UnS/6nzDkiDhYhpAwvLF8XfIsURun52deff
fsFZXTLj9dsHhhfeB+JtXepcXg/evv5/3m2vIqvAAJOaZ55U8TDJKHYYKQW7JVkcz6oRuIP4HFRj
iUQK6WtfjLTx0gZqG1z9fBfkjzzQGE04zf0UcCy1p+X6rIP9K5hn4XQt0AOh3JEZ/BkeCtme96l7
HQ+1fUa63CFLqCEoye0365vHR1zqqbRt/dJAQ7MzHNZZmc8QO80YfR2SHiOkoBr76jAU3m/DtQMU
EKqiZbxhOSpwDOcRns112yOnLj4XWA0qgAjt6ZZ26AicGQwk2eWNwbXo6SXMhcCh5Ky3a/7A7wWy
uJBemvFsVHPI8FVwADeUlhf5VcaFd26yopQRqWVghQBBv6DY53CVPwfox3wOW4pG+i9CfQrWc2Xp
KtER4Bqees/FS6u0uCdUnuvHWmG4iJtS/APY0FK/hsjhlCLgBpQYx5K3YfeX3oIKSAMt9qu1vxBr
+Sk5D7wZ0D+CNZvssvKK4N3zHeew7V6WKI1/8VTBSo8We8/q83uT4Vd1pXky+1Jgs/R4mfnANzVY
2zcRZMXfnebr0g7M+1I5ktBzOrJTgB8hWcfV6kACOatzlevh3+zVRI7TzORv1T48WPPuvXmRCFbM
w61SeAtsmGWeAHcUOTyINLCtqGhRxhrLlA9KuRWdswLVOc7F2HNEMR8opj10bwB+5Ik0Vu+7btPU
rgSmP7ZIkokX3RWwXdsLU/9UBLhMN8P/EJFbevS/JE7/PgYg88nuGCV5FCGGK67l7GgPXK5iCkLg
16Ot89M0xf4oEx79dn8sQCaVg7Qk2Dt6smYHK2hyhMof3UnX4jxZTAXhvwu4GPXkPdjp8C3mcYyc
vEgmnaSkDn7Pp9vRTPTsVRRymkh4xnbDrFfkiR4wb1/fqUUarSW3rvjVzbFGIBg6eJUT1ejwJSZN
DHSxNIrplzM9GKqA1KU02/qvjDdGRIcB2CCWvo1TdXLFcNAhAOyD1rlbteMenISrUn5g2kBtOxbq
9fYKZ4HoobDAXB+TjVVACFWWmjFF3XPu0bGiziBaLyw4a/GqE5d3qW7HNO8i/24ngOVS5Zu5SJeh
wCLi2bE6ktq1Mu5lsSTbBNTKj/5FwO8aq+Ew6BDWqoPmryFOSxdCCRmQMKTn9xXOMGZG+2Pnm9e9
aBsfObRN0QOqsYfg7J/dLambCr6AwclBg2LiRgNnQRKbkUX6CmODsg07qI/u19zShcAYQgDNwfja
eomIDd+qc4acLthSI9CQwiA8qxL35m8c4ArANF+iB+MjP8oeTtAPjLb1dhzaMjTs2Br01jEsh0YM
pZv6Eb2PVx78r5evqK+u/LzAD9bvf4bYZ+MOzjFk7+0B33nckou6rGCkNATNEhFeNzaUo5MIsTIu
nGhBCmwKsPUTJZshtdBTbiJPlnlkPqmEzjsT5ZFSpYdd4or3Nj4aXC+wRQsqUzUK/Bi8ANOzgQcj
N0sgNpAs+CwCU+E4IHxYkx6o3qTCz2wWhpYuptSiUQDdd9KNeZPHIuqS5ll7t44+Pc0JhlG6OpTy
fAAUSE6GI10aKq/NBuFo812HTp/baRtQTBR1I2QKnC9mvSnlNcbgT481rwSr2XCZfLcOJEpmGLCv
AJN9wbvwVKfHpqhOlIZHP+Tl9srv9+r2vWeWq5f8Q0eF7fEhloSuWGXCWua4HjYMvEkNRG0TT9H8
FTpaUzypsksyRS+ET2yaQbXugECip41MfS5Su1Csmrjc/imEKQQP/0Vpib8fgM7OCZRf6ioPZEVZ
H24BwjaDX5Wqm9hT5dj2fYwuzXk5sgtdGoH9+T++zkoSsxcfjLIPC+hmwgBezbQNuXSGM+oSZHOG
fJlm85P1gMnHJMhjEKh9bB7qNahi4QDH2BzP7zy+2NF3ICOF4R++tFarIxN3pbuDtHHry+Ac5Hxc
McGBjnORliT4sUYTaJzRoz4mzbf+8CrC60WHoemnedccZnj6eYw3Ih+/K92jmHrxrA0Hxk7JJYAj
nULrK3DdhxQYtlSizNGpwShtRn3N/oIUpbe4Gghd0k5EVi9fWfOxeFWdqsudtXczPiUWphK3JUVr
e4IMHlA4PD9RZaa6eviH2KZspjCVjffoH1GMQkkwaCuoetmZElD6LlXachhDXyopEXF+MpHGnUhk
EM/T4hEhdQRlOh7RC+F+HiCqr0hm4+QdNPelQz2ra5z+KUv/IXXH9/TIRCaGQ72pyNlU48tl5h8T
cznZZ1nNe64oM26lwBNN4msYn1fQiDlC1FYwNyYcq7liu1p2ZdY3VJWdU49YRDrmwIZcjP+cU3EA
WtcRmxUHoofOh/4H4AvNmVwzhmGgkhSue52Djc/Um95Ceqkfq2ca/shYn8k6DN0iZP3sp7BhaOs5
KdJWipvkCOp/9xr1Zy3GkQ8vUIn2q/wD0/vLenq/QAUDGsboId1z/PE62q6VUKA88JIcSK2K3rzm
z+7HyIs5mM84R6SdDQ6+Kka1vdJHZtK5RH/jbiw7qTQLY/prmy/55VaWQ1taJ4NqR6vLUBtglpKF
AgYlBRTHAlnLyxCt7UAr1WT3psoF40cKRvBMZJokrpmkEkjrwus2NuHC5fEuGlIhsQBIk2l4izAM
pA8/69DhNBVeS/8NJ5qqQIIv+bRmSoXDxvASoUmSMDeutfc3CKzY+kdH7o622Ma4ZgoUS/cLWz/w
LIuuJ2UsJscGeaip3Ph4XHSRjh6gcjtVLLh3wbLlSSrNtLc1ND1IlLZKH2jyTNjeI3ZjlZK+7Xct
Ie8rPjl8Erdzjhwjzfc7eRmuzvtSeiknwX9YCywII6tl5ybLzD4Nm26tyx9zSWKtyTP/IZoQVBe9
xEQvY84gLK/XJHVxjek/eMMDFLc6i/yoWJtCtQiUNtRZGx5T2aCXZsNStQIfdIhY/boY2r7ME2z6
i1j9FV5e7/XdscTaXRVfudjOHWapLyNqP6lC6y0q95RpT7enOrTh1u++4Tnt1gmtxqE1qDSK23Ep
FMzORojb8tHBijcVUmQUeJAGUfY6AWS1TNhrxzFrSzPUNWzsTOHOY14eQepN6zTA0hATVKU2HvAR
IUWei5WkzLenDgW8iVLm1U6N/2ptX13xEHzHcyQnJmEyO9YDWvyn9qvxBorWtJzeIz7UVS8rKAsi
pfc07RyRu6l4HZsYI2MsjqOS9MjrKWrmO+F17imvcaDXC/1Y4CvbBix4C949IyWjl93K/f672cDI
kPGoJln7OHUBtUkswwZK0af9gCxJneKEXWwaf8sKQ/NK1wkGsxp9IYcCLW2ruv47s//TZDEGu9zK
xRKo+lo4RQLR7fe1dF/fDESgwNXGqUVQ4g9hPou//NYWFjrTGc7BhEpFO30WvprVAhAhRzHwu3aj
kgGfnfE2t7Ke375Wpfp+ggp7cq2UI73+0nDxM/mqcPb8QoeG35TvVZglv83cIVKqVpgM2Q2h/Rk8
C6rvG0I7QKdJpsd4QtjwSpAnjEE6yo3yKK8nEchUcu2htSF/hFs5yeOWulhVYuPAspWGGRKiC5kt
S7Iciu4q6SnMN7+oT0Z9V7xuoetfTACxTmbd6Enax6CCAIMyFDblRVWuXt5+vZdv68ESFV79junF
HfnR0RKElexGf0LudFlOB9FvXu+sGJbk8JXk3nmLLZNn3zbD4BvGJ7BqA4U/R51q0byIMhlL+tLF
YNSfPfemiSz8gJt64X2AMMtw9qbSKIn2eciwWfHJgdGw1fX7eSy9/bLL+a2eR1HK3lEutdL8gu/i
7mMMFgiTnqR/nmcJADXhua99ldBSqRm8cUOsf8VAtwHqd+a63nNcXcUAwhnsEMaUAsWoavuvGTgh
g+NtQLAePiESZTqa1yscftTe1qzjY4Ek18bwcjtI05IrtdXAziy8Y8arRZMNe3/ULD9GW5Z1XElN
zCKHNh0RRKS6xogvuG+uKHAjUNRA6ttbAPBX+cYOsuNweIBiQzHX6cZSqbwH0H/V4imoelxY1UlW
p+8Q9IO7Zfbg1f7BVOPByJ6L7mbQJaZ05Oai//gmUTommAkrEU7IJ7DfMBsU39f5NzsF0tpAjWEp
ETpYqmvMeOqg1pSFftHdRhjKcyEdC1Bk+nOSPv5MhCa2KMfXlPrZ+5djbsB+fWqIf3OR0QKCzMpe
7orK6ZKRlm9fHJmVJ5q0zHlrFVLDiTdggq1EfZIsxmsOFgpO8nh6PEuaB55RNLJwOLySM1R9R+GG
Kj22T4IkZGBQoQ8xjYvklRq/EEoe1RhDEwLKShelcFSs0kS8+zw1ir0mC1eSglT0aZAM/ywoRShN
LwkO3nwz/r1qqm+w6mxkrQs1pQYRpsEXYVQBYM3FYAtwJydrIV3+o+Q5M6a2AI/EPwaHVIYq4H7O
USkcp1HBxADjBBnOstOl6NhwAFRipn/UoWTMrdF42uiPkIwBWafjkTgHzwgdWlKJIDIs6G2Q6wVs
3UPAbSYW32gsIC5x5ZhFQTvIq05gB9F0UT/h+nnilGXCbYs6q4k3Z1gyTyvJD82GQn9MzP/5SKtb
GLFNeE/snkO2STsnEjz6d7/dC5pkPMC7Cu/jeMfyoSKPY6RpaYDOlp8m5tMarqqbcZKEWXmD0Zqo
jUVhQg93qridhWot3o6m12TzYZL4mQdupl8YB5U8cGCtVpvPJzR/GCMVe6vMHgfeEb4BONJRXy7D
grbkB1QTlnkvU26TpBuDghoPotmxKAxsApK2XluqAOKcqeztURNYQJ8FGhlhCgrmt9Fs0AHhGQXO
qDycL4v78ejO93hGNxF2NLeVH6XXYBP9Q/yAgq6fH2VdpvCtUr3HmJJEsKXWe1jz60jwlvjLK53f
fQ+PlILlL+hcRIPgpfZ1UI6cUyPqw4UMk69Z/ggZbmwtOxpMfBI6WdUHbEpx+3I453N82wzKJCbo
wVsoxLywDaH4ml96N+0EORUWmKJyCz0Z4eXOcr2Er40t3vlLPQvq2lu27ZQQtHu1lKpGzojd/Bi4
8NdRCBfNf7esu4hDt2K3Uk4BR/HDvpdW3qDsGA1gr59ugToUArgAlb3mbIRsrFgWUdB36rEepOlX
SdW1pcDGaXnAEYSOrnrpWtSbV9iykKKdhRVlAAarGjOUTH6ErOLBG3CWRO5C50vomhPDoNjZV5LJ
Cwsk7cGDehQCZrKM45Yqdjl7sYWYYiv0CsQxaMqvXWYLvRQS2mjtxIfyozJdQ2V0qGA/myw4tpBj
CLkwmLn3phH/Sj0jQTWUKt3zOyr8XEOeZjvoe41QxeKQE08zsk9WfoRrUVxegI36JtRGigrY1Y+V
ucqODqHrDIfJ9Fheio4Ejm6nPpd6xLn80lNeXKVXrCnTIMM27Mhz+jzoYktm6o7gYCINdskLNvn1
+qMn+fzGnX9IFd3GJRshl1YEmEWE73/gaUm1cWPtK5kh4JU8f9KeWNAKkF9WSyD10MZoVEVv0H4z
o3FB6pEPCs0vp+G5YywJ4N8z99A3VCaKBw2Un1zc2U9hz1wnLIDGTPJLb8FJc6UXqzBOtb7EgGnq
1M+dTLcomCTR9RIL9cQSNNLW3f6g6mxsYw7r598uccYKU78Gba9bx8P95EoAkCPsN+MbXInoced3
gTdR/sJzLcyL8rawos8xS07DhCT+xfUl41XhQI+TmQUbyY8SY0DMBYJiKbpVk2lrvxqOcKWc/ytw
EXAqlTMprHAdqarZXqGb/h7kUkdyfuFW+3Ymv+3F/2D5sSuhOsTSvfOcdSQKIS1JUtBsH6v5OHQr
PdpWEYJtqrZnV/YeKIK4Ztnuhe/ORgFIHKMwgj63joaf+R5GGz2MWi78Ou8prx0IniDMalZO+hTq
xb/dvqV184wOdpODBKQZHcY4ULdNgLyAp/emYL0V6Qmpa/NON+dKN5F5Rz62yBX2rzl8W2KRgVZW
k+wgOT5BrVjmzJhp425F36+z0Ne1F5UNI+YZP9dbMrIn14DkVEOPqDoweWLIq79UoUEHlK7/CJzG
/u9cZiCqGcA6IQsv8goT3K1RwG4PLK0SKfFxEFY3GwBKNgYbAB4ZO4iNF9Bq+6ij6HzfXirwHTpW
Jv2IiwKygf23nVF0rTm01LOrHCG3ro0AeF4z/LOXU0sawAnCA9vnKGMN2fJ4huC/EOfic5fF34Kg
o8zmjdR/9IWt0qNfsMiv/M/ENb4RFtbnje2jm2C957ZLAvruDXDV8m76KpDWmmQM+Y1xNRUbYnrz
U0WB5Lz92dDcZ2uyZ87Ju759qCrG0xhSMt/dpLFTbyQeZy1fobFezHWKqMTgoT2c5EPJnIfU+fDx
NZtBd5Uq6+oYpwgFwe+mYQiSRYzsR9uopfGb0i5zUXMIIuMztuFN4Yv9ftv5AYOBD4OmbwRVz+8g
a3KHR8kaTofaOfXZI/tKsrB786GuGf1RPPCPbo36QpS3ZMDI7yNcPhVYENhpFumBcbe8sACrYyTY
AwQKkIDCtiiwUdUt3PIaDNw3cu1K5tIKq6B1UeUQh+8ac6aZzruQaljd0jy9vQAbPDbKQxFb/vtT
79UHfCQQFEw9+z+yxCLW+ZEsZt7Oveu5p1nmL1cbyCiMVCBAPCN7v2h4ROx4CrEiUt7XodqyRg/Y
w0M0jRqh+e6cOkPgYxyReerJ5Kibel39NxpjWKKy7NbeRMhpvrE1zQfkwrqRkMDt2zrfj1yBZgel
vfKSGxxhBjVYU2j4GAUYZhIhcjyLhmnooEEg8BcjCq+u227rRiESXI/Assv9x5obUf8Ohmtf+dQu
LVEXnIHU8kCUu3CLzrV6kKLWJ0fI3KgAeSxoVECIfirDbD9yOjmhAilG8bNEfAydAjNTpr28HYX1
AQ3yj8IjrOnV/tNEb3NH5P8MDJxoykCYB0exvclBXZbcT+pm7/kjofjDejR/Fkr5Ig9g9nvtGi0C
8LKQXGknbUfjoz85gA8H1oetxGKINF8N7K+JriLRHbAu9TQjBhJrpDgPuL65NIjSJB/ly9ELebvy
KZ+TDQ56mxqxCNOg8o1q8+16KXmBrSWvuoYW2zr7SpZRnwwzJnNVV7oyfS9wBm3afQZp7dETJfJj
hCTm3PK4r1DNL5Kuk4SyKA1G5jGGwfRHx7fqhzxgbThDCKZAZXG3wU+iaFKa9gzohUq8bw2K8CL8
DmenQRzGy8BAY6D5OmmayduZNhSfw66+J7IRs68WPmE39TPJUqFE4/O6QdHvK9/hCzTwVf6ZOIPz
1ENbOLoa4zMpBwEfXo4hzixdSiJJq459CzqKuUdaj3MK1OwTc/pw2DyE8PCHHalNlrzqmdJd/9Xt
QLMA55vIeTJbBFyimpZYvXJCkBQBYm8EWqzZOf/p1Sy5GmAhS9rQ6VAM87Dsjog2cYC3sdlE0WpF
4prGCXtcCd7vMTcYE/M7+uBjNnRnNyDXmXyRkEwGSnl0TGZTbG/ujJ3p9mCnvGNZ4GwWosq3Afge
dUXSi0x7TEu96UO0ITIckZHjWmz4j9UcI9lz5shHVpfcRxVTpOmvuyJXczw4RA3KUqkxn4HScJNT
bWl9WKjSgYPAuzYLT8tSJSEwLUTs5Y+EZwWWH6BZuZbpMVOZKWAOI+QsF+Yauk2+JG//+rsgXIg5
FshHpEdJPK8ILfftrrD/GSumA4QfmI9rgOHyFDXJT8Bx7whK+CtGSrMgk5t6EZLbuqHGk6bFZqAs
AvJU7pHDyw6CMAng3fR+n/JtOzvIW6zrRJbBJ/H5XWtNvENPdPgVj5nv7LRbRgbxm7gzBQAnvrpC
NzmFVYK8HbwKd1RSji+yNgz6i2au20Ore9MY+lvKB9Fky+zKoaBv461irdTqw8jIf687wWOKRpjQ
g31yaKMXCi9rZVX/0zohM0zjkLzyyLYs4Td0svFANWeDfzpIDHYDbZKzDBxAma6AH/0JDb9/sU/V
JSYsD/U+MnQeM/CCw1tmcZhEyTn4zbKTIilBvnz+TdDhh68nzCdkWZyaJX63467ONOIL7Wsd687+
rwGbWS9E5DyZV0jTxCHlwXQ/RkqmiGe4JMPBCndyUfLue7Dn4o3fhFVAzzMlGlLgpeS0KnoKkZBO
iKpzeVSR+HxUHaNK85+fQJqEILEbKwa84rCRQa8kOHKhjWJCHxOfZYPe8V9B5hvn1G6ScDNk7O1A
PEHRE9T8Ob7j4EqYChwywTrrtQWgIAjN/ykPr6m9LGtdh/zB1Gc2PA4x8rh/7m2Xa/YLOXzOmBF8
XyUmuEpGRpzA/IVdxDbRU+gdmNgJKzseb/9BX1aj4wzg0Se4MTsBGaskaJ3VpWF2K2fcHn8vsoNK
O0GFs3y1IhoOhjf4vU4O3bp5dGV3VVljD8Htk7PlDW6YeA7hsFShCtdrOm0xA8C6550BHSJrfgdS
SVqYCm1m/nVWUX9EZUyh+5pc1Za9eNgY8y+W2Uhj6cuQkVN4oPGCObwcTsz8Zs9rRf3yC1pDv2L0
tgomVpCnunxzoZSz83x5jFdpv307vdHv5RQsPgw7yDJJPrl+KkpSd4C+51OgwnqvXvxb+dfwdPQ+
+vvMdQilZHUAWZsCg7V4DdTRSQ1y1sJoE6EPoIFrFsxlKPHONPFSNa+S/ejV/vUp1mae7bW9vw4I
7ly1wF5TG9UuiL3dzfxNTSCwpXdZuhwVQEuRYOpKAT7HCup1tESQL0oci2QbrebtnPIbDoWRBoNu
2XNmeKMloRruEUGefyVkh+y4pwlrmsFxqxa6toZCfEiDmTQ8CJIhaze2oQkYDnI10634R7WYFXjn
QdGcaErawuG67AqUp2ZvYPJ0Ie+KQX9B7VePbwY+A6h7dKDqtvex+JMyEop6gbv1Z5T7bBvgsaqs
ADCAiI+XiZbp3vWeMMJV2OAVuiKu1aN1ST3QUzhjEbJyp/OROZfZiQGB4T+07dgaiIbBo2S7XGaG
msQjsQCoQTOLcJY8VtFAd7GCnscu4dcr0OJ8FZrTYNcqCSTWZ/TmiJRHqQ3x41HOAVSE8Zc3+iU7
ksfjUzvg11ilfrUXYzxUtePNubX4oW0acRHFBIbnFYR1WuPfWCLBePmX3kkqAcYATUVWTqkmtoG3
IGEmAfCCb/1MeActJNnKRERXl+SKlZWb5sFOPj8oQbF72fO/V87eMmDAEULAg3tmeFq98+tvANMB
gKwAYOE6BwFcTRbhx95Yws5GmKMCm4MOgY5ItnS9F5eBExqoLEuSYh0Uhng7QhAvw6jAbhag9bFX
r8UyRLFIrPMJqi8C0aw1RiJarcY8OTGC7DzxiqvpmvrCl8yMBk3doN5g5Sgrzhvj0V2ymIkhN5uj
oc2uxzAE84d988OA4rfQfkAiWACytaKyiaJwVTbmLvPceV1aEKlI0Qa45/1ezEwAMy1Fhe3Fr/lX
S4EiH1ThvV/H8kz5rRZrQ19y/kXG0R9qVIyPEl8lwwPbMF8LEqdSMK7PYhO5D5D+RVSPDhEROgMY
5y+O5F1PlVz7Um+Gb2ou8RYo4hqx504upOg1rPf/Gol+rWeos7JUMKvg6CpyBUM4Olla65oUH4Pl
LQpaIoVuWeR8/tT3XSD9SlKk1cSr5S2BU6h7/5MgCG++Gi8o+QFvLzBZwH48ncDvUEJvyvcPUJUp
YtmF3nncf+iOZteJna6U2lAMfoE1Va3QVTTRxGELqEjGq5ANs7oMwKhKqZzQnorbE+XeJvCbpdEH
8TyZRZ8xBpssEX/TLkbunngpoqb700dFxKm6TDNlZOSQP63o8lGVoFFRMGQlom5olNc2r4zahsKi
GhP5VbPSyEFT6qeN8GaamreiMdDBD6siND2xGvKCOoLH/27bZFTkpFueu2LYD4b3mdpmdA0P7vAz
vt4aooGli3FyF3yF4K2AVucYmW8WoYoLTrNV7vhNhwB5VaEErPHxBa83vmaD6ivtA46wUVuhnvXO
fgAtHrLo2UEj90QlO5m7gI/B0MVgGeysaGPYEuaFlCtiFU9rm1HNOKc1tQWVjg+GZHvQmmwSC60j
NIIn8uh9et54syVtIC1cC4LBf1I/WnJVX0XUJ3tJ6FNYs1h8umtGYymp3WIRckZEEjmMX7NEkNDr
q5aF64PnPaIqNiiVB1JTlTNRAYcDE8qs9mNMGJJxtC/MqmwJBGYbGmevgBTErk6cDFZPN2gaN0eD
ikT3JYjoxFmorA0vKw2njUrHX+YsUn6jjLU2A913cOdPO8+N5qT+7QBvcjmIyY/HmH9qgFY6DzPQ
XQ8lzxEzCSBHC6p2Rn9iHYfxS52M+LSoW+z21RPwoYbJkJOwKtaARsHJLD+vs6L4O87K6+Hsisgr
A56O3QLHxWpjOKqdLz2RlB5qoh5A5ncxGHMw4RIqD/Nkf1CIiSFATYQfPVYp+wvrtWKZpaTQX45l
Jck4r6Cq3ukM9C9nQrmK7OVkw7lThaf/Rka/EpXl4FQV8MvtEqh4Yw91HdmIrjbIiRy0WZDkz593
IMxqiZlXETZ1j9SocC/q4Ldi6Wp1teU8n1dzV0AxGgQEfLHXEQPyvL9VubJaX3FkpOzo1KZEnGuP
JxqR6nR9LueerK0ZsRSrEqjZMQ61W//MnfOVGenrzLXwR0kIVzpf5qJ/Spkr93GnY789YjGfluXa
IeprM0WQQZl9PYb+XPOjO1kv1wAFmNR2pJ/K6pFvgsk8yGDlOaySI83NeFqmd+Gtx13LZs1SyvRE
3V+UQjHom9iWc39aKicqOnzyyoJ5rKSHPGF+9stf+kCWgUaFl6sytbqIId/P3Bn3rGtXxoAktcTy
mPmGhxYQZdq+YrDjJj5PQdNDqjqhV7t17H/ovuGYPcj4KDcqEXiQHC2bAMTGgXk02gWS8ixjlwJa
E0N4RJR5Ibw8pYRBjXSIrYNXNfDuovCtIDILvl7IQ2xofHi/byKVD/VI+YeJtSuoY+cKRIcFqf/Q
fWpyBePaL51j3C4OE8glvS0MhzvXnSSSEsAoHXJBVCNx2YLCQZ0dQy6NWhTOFwwEy1oNrvuvJnRH
Y8GQXSgeMuwoR86k6CYEU8QE4ukCu1+BtFVReNMnCt4/4cXLZ8hhTEIFNyZmkwSAur3C7234unKN
eEZRT0HDaKEq1x8sn3W0uYVNLR4WHIA1UNduEbqVcx9qDEgA4N82c9rncC356R2NgVlFAjj4jCG/
gkUlNAXVrhIhVo8Xdn12lUseOPCzY1SI6a0nqe8xHEZZSw8cxvW0pDXIJT6e920SjUz/ojhcMiTb
LrWWZ6xacS6f8QHs8vUU6unIPHKq45EazwplosRmcVktSCB4zU2WWfuTZey3mXvD4DRPT6g24NeH
QXqXO8r9MGmDZ3d/4VsEpaiguRNgt7pkaQajYbIWZvzytrLG7qhkvKtxGZnYcdw6fVq3gO1CveHm
ua1NMS8300Kd4AONtIZOW5QQMQ9izGCq3j3q96o/eL1L9RgUPtm/+XChL339FgJKqp/tyi9TGhPS
0TXm40ECtlULRlzvWtqrsgm7N5zvSS1drCr4HMbs09OmuWdxue4goB2mcxbTQ2H/fbzJt5Prx+yc
liNpacONHRJJWI3CVwshyi65+QMpUvzRGW/WndUW+uymcSJDdFM4b1oLWeKR3Rff9z5Y3m2GQvwr
dIBDuJS/eWax1yeNTMGsKzCRPaD6E0yVXyChvBWNzrG6YjPCh+h/0Q13GM/wuVAzkypnefhLSPel
u8+EyHWaqX3JWvs0V58N2qL4lbx61ueip0HZOwFN1ymsc+LUiFY96ckdJ1CJHcDrAXV890CdK2NR
OvGxErirzd+MsRbBF6OoM1hF0Q7d9MPkl9QsdOKTsVBjKvwQW6mnP4IqvhW1RLL+2tJ4Tt88ScE8
RdZ8x7ZsCjxFUGDRKmPavaX9LNfQKfJSjNHzapZYLQYYwDkO6jI4+YFCooogwnmjs8vIjyQ9nSEG
SIfjGRzD801oziTiNi/bvuFJ0FfA7lRU8ofhA+7WPfRi1WcNEY/wV8w6VhX+ffiPGLNT2tjN4G3o
3JRnE4ABJT4IOMl3ksOYRUTuCOrzbm5Fx2qsEMaXWUis0ErvHuDaia+V/tk8/+ISiOkccCEWfF2G
rs0sOBuByW0FARBtYg7CWka4xNuqXf5d7oNM5NAtlSGHsW+qpIbSSv7KRwkQCw4EBSvKSUtK4NKq
ijBUTqv0+K9Oev3AyS2e9tlA7rdTvKLuC9PlUbdKKjJXgLp7yonJjqLcUYv/VuoAOxb/+D2q1Ibr
VCbQPyBQWKWFQZ6vuoKZUutd3s9G4RTCTxkqIRsae0rKU3unuv6ceS67N4L659MCyQcW2DpHYkbn
gu4Q6BTEuK9mzQVZ3uTSIAzJVdvfrBD0ryjbuMfe7lvxAlsYOvRhmFVVyFl5VNOrhc0hmODEC0EO
ryP5zviPUhBFfHQc7dbNLncPX1XKa2wpKS5tQ3My+u0dYCg5mzTIEvf1v965sXOEuvKoYCG9Apxx
42ADPPpp9fRX2UcUVL89xCHpKjolMQ1czXtskue0ToTCd4OEkwkYdjVihwIHkYwxbEyi22o6dVab
qquYV8gXSpPQ7X4TCtlu2igrRmylVSobfnxJMTwiLcSzhNnyGlQI2cube/qO6cPakIvKenMJ3Mn7
T5KC+4zYTvx2AW8954oxOoLG8lq/O7RZxLbHtq30zsCCPpgS6Keex9umV7EdZ+4/mLW7sZVAzgbQ
qYKlVOgglc249ClXY+tbdwBazEfBslHysAlVh2BP7PIRS6TT+hvX6whoibILnbtRdXbeWQqT9LKf
S2qUDw0U20ybx1bxb+qQuF/5bNGTiye08pM8dAkUDm/ojzu2PGxiCCD7/mJEyeiJfLaQ+5rLtik2
NJEMSvTpSWaysVUmJvhW427XLZidUwfQa+sEz9a1ZZ8eVtn/k+miDGrINOh2D5WnMUTvH82177ny
pGxJGHFnQMMUJJvHCy0K7h1OQDeRs9vYvVFvfuboDGvKhVdc+dHuSllJIqxsblvFevSeq+R6fE5U
CvclKiQUmZxhDwn6hnLOtav8iG+eoh0YuCoEHfgww5BO1Eqr31AmJ9wza3vILsfQSctrpnSqcOYb
ZJHHoZGbdNMdeWA3C79KI0bichQPMgOan1UlxPpPVXwOEj5YkFe+0aArUgiE9eV4WuhtzWBcAQGI
2R53xVa7PK3PEaODKBOVjJC7gmbhs0pt3c3NsZmD3Xq8Lg1oy0VEYFPdHh2Nq6lkuq4ruDoLzzFh
n6RFg2XS3yb2nguU6xL5gImtOuuSQv5CYQp2G2lPFxhSWzZxaRgrRJfsgabAplAHb0Dq91xoIm36
49PzbuXT5Kg9/vCcMcUcDVpvhEuTQQ8gJlqi8Jg4JjhihKko83Hv1XLhC3IGaSdxv/gWZTqtnhti
iL4xMNv9kEAlyiiUIHzOx3BGjEniOKj+jsu8NwWnxVLp9r2ggGFTWP8bPYz9SsHx5D4M/VXP5pfs
re3eyjnpfwiN9z6IsVttoZKrOjm41VR6vmQVVFN6LzkLo5sjB3C4jlmUbivBCEICGsVg28Aqsai7
EmjKP/cSVmNFusKrDz1rUMOpBVgvnPuPhg/8ByXRzZc9zLfNNGrc3rVMvjO82rqk4PZvWD6b0rlB
e2YwhfyS8gnIWR+zzcuH77lfwnPzVvUsIiHCIofKQlXENqo5Ur/+vIIxb6eS2yFDOSHCu3x0RehX
msmtZ7iDTcqNKii/WqhXM4zIDMw8pHVQnAe+jOUpKGGk9shz48agmffGa0FlRz6bLvIs0em7q+ee
SCN11BMjCNvVe9UJreqgSzA4dYuFdjhzZZwsmofaTunDxtVrJLHDCBy8v8mRBHhfkpia61Z4K4hN
gm6awEDDM2dtDnuJMmnz4rGtMejAPcFlSww95tWB9ri4V7nh/B8RdDtxKrIJN0amtqF7jkFBio2u
c9NrjEWHkotOy/QnNJ69TxwMnuR8F012NwT+9e2Rh/bsPew2CfdlthkGWY0mRc1T17FGhRS0Qezk
k+rjagt9iPofXingwSs7ur0h2z1eRRRBQTH7bprYCU7BkF+5sP1mHHhIHLTUiiWJ+r1tgPfMruxz
7LWqWiikTHOVm9NeI7z7133BvMWGfqQ6l/zOTmtSzCH7uC0ukASdprfoD0/D372d7jGiXxOQEQVI
rud1FZbvyNcFlnJb1pA2y9vnO8v8YgFLKC3ECjPttIuLrqw5Y14UHnBleD/f27APkUc1T1GBClRR
8jZ5suI9tj9eTJsdD1VHc2UDRHOnDZsRUEG1Li4uHGGhSDmH31sDr5bGW7ql37K2A4hr1VgrTNzL
mYIeIFM7egQXuTbTUFmv4+LiJYJI2FKI0PxL8/AOJgFztJCvi3SOay6S2CMHILApUUeQ+bNH/If6
WWPEfeahqtqcu1raoIymJ8Q2A8yMFRe4GaU1KNf2HoQDnJJ2pmi15pyO+bnqSOZbMcIN2Y2p2AQO
LT2tuVdxTzOX6z6BIp0mremizq/2aDou8IcNF49OL59hVE2rXZUQo4lV1ZNA2F0r0yzMSMfKEoxL
DPajqx6AqUxmXhMpia6Pj7kOV0DRbX0HejbFsI7OUHjM9EHZLyb9fEhGD5s4fcmzMqYvYtxSpMog
BJiwD27QKzhbvo0w9jeii/QsvxqFQnJ1Gp7E/xtedf1GLtHb35F4kMa/OSs9K5AXRSrVarQbPGM8
BMoMTDbC+5eJcNHWWBYRrr98MnKliyJUAQprNMe9I6dVpvNXQEwTmpkW1JYWLUzhJOBG6vrGCy65
e9A2fj+/QhHOkc2TfzEcymKC99+HigyJHROEqfHoT05SDtDJPThOGH1lqKgPmUP+S8SoxhQSW2ml
ttGlLhTCgX6Fc7gVtesdWKoYaXFlpFA+YwC2tnr2B+4mpVQnKj/ytVHmgUvWhSx6RUzz24jpHnya
9ePHAdl9JizSpTnpFxP/F5Dc9z4kk68Dkh592n0kQJIB9MCPkI7NvO1tz6ktms8K99tuzT1Iggvl
U4lf57INrBJV+/p+4EVu/Xx06Q37avigL+0RTY/g+WP4KHNqSaGt8UUiO8K+qH1BYmLt9SMMs0Pt
qoN0knjLVDAQcfRRD4XC5agWbYaqqAcVWUqsmTR/fVKuibUjdot4uYtefUDeg5TuSmyvGd6t/Qhx
La3uSVv9/gzk6d/jcgoD3g9FKiOU5Iyb+BQOroR0lKsQhdY4vnSFV0oGCGO2qLYuTa3GfAi23hjx
d+HGZOdPQHhthEIuznr/Ped87tiHsL7l1+dBfajhqqNcNbjHy8Q4eaMUxFcMMsSGdX2JI1AJls0z
zv2UFASl711BAHDBBAVVFpZdA0OrupOnEXtUuH1UZ5TH8hjQ4e173o70EMaZ0mRbVVyT89xHrND9
jbpWRoBMgJ7qODg/J0FImJcIHc91HQVPTfdeTkqtiEydd04i8Uc1P6ZUXggv7AzcFjMQYoZafBrK
O1oiol4wNtuOyh4RfELEFUgun9NxmEyFxnzKuNAXR3DXVhkO3BfhqFjpQTYkDMVYZLl012Bzs/on
3Mo85Rblr2NVc6+7pwtrUEeVku1h3+7r3nhPcTQrmHuemhH6g5AZda/59jiMWasc6W/QmwPUqGSs
ZR9K1vcEZfCn/5EOCG/9tz9fQSPE+0ezczf5Dn8TC9f+pkaThcd3KmSiCY1X9E1py90BS+enszG9
esT7JkfHPu+f+fbMNF1VGymcbvjh3H/W0C+iXHg0GFhSqGVkTW22VXmZ9dx0n9xn1jzQzkmDPWza
J31MvADcIgaj6AhFPcvAebd7qozWdMxwIFEUNMK5Bm1qGczzyg4WBtyiGfm2eWcH4N6JMd+v10/w
/oKDGE2xF4cjgLaJd0IosulWz70zS+0upQPi3llX5AQi3WVrxUc6+s/D+GO5CEByh2OzFG1LM5FD
w3fv5ffSM0wqvqOq1Y+hNod8dZEohHBczOpn7HOCQ0pfMwd/rksriZImB92gjBF6TCP8HzTJKMK9
2eeHJZmj7V4VgCQFsxVJoDhbLT/GKc/CiFf7h8S/nRgbTbACcCscFqTAZKILbhMHlWQ+DYn4j7d/
t7U/6H33atqUASjQYagg4bNQs9VRevqii/YwOljTgCWr1zGVz5+S4LD4IxzmqZx2hXl8OCrL4nCh
AKnP/IhCdoy9rFk8fIAP5L4ZsBDQgOkAq6KkS6AsXJ4PXQp4jQeqPj2dMzHNK0+EtE9H34RfRMXp
VFml+ogBkKZtLwgqIGhXa2Fq7QqSZN9v8uOu+tNt5vIrgxJhRUT0ZXWYFcBRA7gFmWFUxtL9FYuF
qJNbBYK9AL1juvqmOylW8MHmHqmo4Od6E29gaujy5O1DZJm0XJHGbgmP1sydX6PWidOQMQ9m5F+a
HWkpKsOQq0kBVcRB4YRwnLMrpDDT2eiavdZLi1zIFSklWg6aOaF77+CINigeB6FA1hoQcoqvhN2V
3QWncf24b9xepCiO2vg/RQ7xYYqtTOfsqPZd86X+EVxG5unjdm0usZbmGviQeQ+lEZPYGE6fqPRl
/YECYAq+JafK7r5kTJMoaEbmgvV5cc10NncvgPMtYz5++aqH4nmHtTqIZQDKjLIOdEo5dOa2J5kg
Lcc60BCljXDtUJBrxK4FE76gQWGC21z73JTDqQPZv8y8RRk1OPu87MCNLAYLW5obXMopCNYpOojr
P9yg/DXAyyadOy3CAt+bmOdVWDCtemZcPTOsHmdQaedlA0FxV8WhiVXBroLQ7sCTLU4/rPp5Zj7U
NVwDMjJ/Mic5Wm0yVzxv3hjwTu5enhPTp76z0PoicG2gAjnPl01S4YkmT9OUssfnC3Xxk0jGKwSp
a9Tn55nOPSpjIrs/RCoTUaXD26azyu4hTq+oUTjKP0WdqPz6JY0nsa7j62JOcHDRrxVyKoY6eVK8
taEnvSFeKAbQuYdAgeka+5SmdXsuFmpIq3vZFHZV169jASsx67uif2kVp7FOcFNSkSMs7eZKTRzl
YM8O0VRMWbSm6DlHZWUA4gce0GSFFXNodMv+QZ+z7AXgUrNzSJg7c0IJE/G3ln/7IYJyb9yxW3+f
Fdbar6y3x8kDqG7cF2PubKZWEb0rl0VNCiFuprYT11Q1fthkrK+M0fZpALIrF1GYWnv+EAxWRDV5
uyvUcv/Sd4pu0dYxVEJp7B7xUeHCi/57ARXLxUQD3ZIniKfXOXgu+Og1gNoMCf4UcR38XIX8BgFG
VpgEKfpulmQCdaU67u3ucyzKafJ0kFmhdR5e9CdKwsvbdf+cYmQrAkWPLJJ7ICLf+0CANdsJLiMo
qmysQiDrZ9AHONaFI7SGWZXbiZdPc8OTQkAlF8R7chhQ+1UyzRjzTM/VaQeLvbqx3zE2YOesRxpr
a5m33ZaNTytlB7bFjgTuEHImIMSohcHcMDra783gcSML0NLKHL1aBZae6FWFZ4LmIRD/FFktLgql
v7JKV9L1vn2sMvsifzaiNeIHgFTVFz6bUOcKv1iMqa+vyw61qx7vSsJ0///TbYw8m6Gn+jH78M4Y
PGPy+jSsW9OwQbPI9X0LDaSPTr2jiPXz69k8y8LnZE6oGc0qE0xf3ykyjmWQIZwLYBSU+wC/Y40+
5gQE1qSg6BJYWbU2s+kaEd34CvafRDyijpEi/ze2lbuFquysfwHx6EeKENkV/MSikNRB8NtuWkxA
JZugAVkMJYrAaochq/kFSHmG6yFI9UYOvSWu/vsureVbjKtpkpTaq9/Xa0+zS1pVB/YRKCObsSbg
z3bgzNUJmmbOcCuKylHeeEd4CHei7+BSqQ0n4L6UejFEGj9uifm/ir5b6AlrV7mj0vgrAMbvuuji
mUJPJv+Rc1Djm3cOG48lw2GAfg/dW0WNRIixa8Eu65qfITnMFIjRVm65hz9h4HrUo+NSnAuDJNmU
QOJunY5ycuvMN1j4HyU43qOmfrPlIuQL5jm0VNDrYNr7Z3QEoc83JhOzjouhfBjb3MFA8GGlxst3
uBXXUXCS7ccvDVsQDcVvmPqaeaz53Nv3L10N/rSLHcpj6U6lqR2pcjmylcfev0MoUDpYAiluQ7fc
+oQheStvK3NLObUmi8tNuW8NvW8srRaPL2GBx6FnvJblPzqtm8Ed+USVfGcS3aYvJpSps7rmhMhh
bXwwf/PeLBGDRxxdpe+RDUQYKy9WY3RvHTD7jAKDqkUB2TNJeoCYFGAp9eao3nOFp65rOneUH4U4
cHPxUrxTaPsvEIQAgpaM5ZFmPLVNkObIkGyQZDBzI8zX9mWznOTl4kMowsdWbXxPxKsdXAxGoQwj
TSwfAkMBfLsW5ZgoP4jwm1Kp86sC8Tj+ooFwMbS07eEYI/52ZKbRHnVvD8AUKtSW25gOS1L4rItp
7pUCITkeNTmrwrZ+DUGrIjgiywyyagn+HgdNIPkfl92FbcmDE3NsmfxLK1gmYt/GN10bZurrshYp
T3eX60Pwn0LIdeCoqffp1LucTP08yxEU/3abQh2o+qP3s3efQY52+ttX6ibjN23T/DykTCpkiQ2R
oVV04eyhwvvuFSf3q7xtEYJPl+A4YGiz7cviJzGkEVYivKSebKue8i7b7Y89NnajX873jhrW/toD
yyNT2gfAe8jlnMVMw5zeB/kpjySl6jc8Y9qVLjNBSc0rDs1nrN3xlyingMOb08QdUgeDwRSgjO+8
ae8VpeK6Zd9s/BuKiUyuF+FuiDSiocpeJYn8OCGSJWnXULkxAqoO6uTURfleblEKDdjMRUKp1Z8H
aBEb2vc4qZ5doTuOho34keZc4KiCmAY6AV+JO3N4AzgyziLUjQuV1cmUK2BATJ2F3/9KUgHybB0U
CJ9RKW8/3i+5JJ8+HXiQBoUhW2Hsph6AsAz/Anc157ESA4Ftwy8UcC9gTEHCtBxbp6C1J2yT6W7o
ImP8T5w4iF/p91sGZ2y+xTuVduieT8LwdgfO41Zw81VwbKACnTx+ixASd06UP6AZW1E7ToDRM5yl
9t4wOdFZHKWYOW4RfJgqvgEo9MVga+iCrL5tbcNPUN1fDwRRbYj3H433xuym8AK/LEtOEqQbuekX
y7+5HjLaAG/4k1MMJOSmRDwWmZacwMdPFOUovwE4Tycv2C06iw2o4lJ4E5ECZh0+v+BjT2yAB6wO
aMA8Bi8P4oHkeN6F3bMSH/85im8gU10LRgIJh6RSh+n5wZMkw95OwZDaRgrVgtG8eHNclycZ3JUi
oqGzTNfHHKai7IvmavzUwkod9k7r9hs2r9th44+nVRU8wqyCKajuw6chGmb+ab5XUzw5BHQtITDj
hpkPvq0MGQMYUmJ9fVZIWNVXzNgRgv48hSOd9jxXVH9JZk+QWXWCXz4Od8G3yGxfxyKusXdaRY7c
WT6/dgNQ7IuHAD9EM9n66CEBPp/cHrHjHnO/HnFMTdh5U2734VSBgbNgxSXkNE4I1eVYbIGta3SD
bB58Os2eUiYLhf3c3M5kUfHyM5458P63OAvNqledmvHBDPxuQ0CE0/QPqNrWffJbbNdQewfyZWJr
7HATdQohiqtx+ei0tGC3z7qhmwCd+/Yva3yW7xGEeKag+y6GQ8voIj85s9r1nXZHE1LZZzVk+APP
rK68R50zcxTR9r8yoqVvzVFUQzq8qiCmmfKq5xxEe5SbLPKCmip8zThnkJDXOzL0dO5zz22vVnPM
Xs3k4ZH4PZpMvBNeH2f3KNPbeJQGRJCeVIFy8klfr/PnRN4Uzx67cBji50QWww+5YjwwZIaTbjI/
AmL2wa/YFbxZtFsrVykkcctMI+EMpB3m+aZA0ta9cIwprogQc7PonXh3/D+jjh/tAbFCDU908zm9
tcig00xn/p8yiKdH2ncCKR4oVLTiuOxO0TByRw3NcW9iXvKZu6JeoSE7L2T+TtJDZEQ2VqqzwEtn
XLnJsyNJO3TcnHMYemIKQDq8BOl/a1rhVrVsHH7NIHXRX8zznEc7Z6RxdVFFPVAFOo12cAIqQXgU
6uuuozlikXJ+wdvBZ2mTNCYUN+/Mycu/tvk1ZoLUsXhlRHaBfSpqRJC+5yu0jc4062Lb5h7UefL8
rf7o3TbeunEigVUEZ+meDdqJ0qZvaT/jXYKAYmPVYv3J5kb8QcnY+5FpQ34qovW6VJdq5UTwOUpC
lqsqThxShjx2uZnX/HkLHJrh6mth/Bpplm+/P5BufEHH2w55QmLfOQ4wV1FcXmKbyufO3b+xFySP
4EdeT2O5nyTAg8R7XYEnMEayoZEI7oQpc8HfRipSboVho18C7+By2KgS/YCA026IRIf1xqSKqEjt
N6/jD6dNNOxEC7td8nX5s1EP+Nxy3R9CmOMthCSHTU6u2/YHFS9HTN/cyPehyXytHBBp1dwylAoK
lQV74hmNDn1aObAY7S7iejIzBTAHMMAFQ+FlEimxQI2Y2nKgkOP1WZLxqAHEikl1Jk7hlayaOjqh
EltZVRwsNn98NH70oRWw+LjY5zdnM9IR+nLGQfowKGoYPv3/L4qve06PEmVpaEN3lSponSbjm9cT
D/p+oWZvg0aUP/UtNq7bn/hXsE6xIGUCiBTs5nwlJgx1WH2+hJuJCpnHjCDjXLUxbzFRV/eE3Wrd
zH2uqIhR4ci0e56zi2GgwLIWZlprVCQbKg6XehW7Luc9EyiBIDrV7J2aye7Uaee5rKqVqOxAEDPU
a8z+9HBdSBW09LpU8HWFW6Ft6NVA+jtUZVFgvirXfssMu5oPqH355GvGjajRhpNMlv8Hhp7xt/DP
an0sIediZC4lxxxOAG4uR9Fwvff+uEzAd2S6zwmWa3vnPXtaA3GqlIJfQ3kjYKlW2lA/W10btZcd
mN8elsy0Dl+utlMgshoDusFkZpkZRm/vetvv4Q4uoXzhJh1hUEz6rndIFYqI92The0UkRQpRjfrm
kBxADsa1P1Tj6gMfmpqncKSeVT+OG89ywUqQm7ncJAAp0vAhyeTumrX/UdD89/ic/HQk0cYxr0Vr
3dzmCVrR5llHAumfrPFmwTzCixCB5oLVOH786Aa72Qm2l39C/GMjTTd63X4dD2vjoaUXqh9/qfHr
8Gwa/G0GWs6T3NgRBmLEH4Xf0DnH2kr1nSFeyOwlxans1/nPcRHzqanz4acrgyeys/Vqk2BsCm24
aslLwMr1BjcE8xmgZsRG9gXrY0lfkcidFxqMASOIkBSQmS+hiCKLlYvb37J10PU5oZMfmrnAtuS7
BK5dCf5fGLOK6FZwWcCHcE0G9p7Q+nyW9PlZJh43jrKEvQxL0GflYgAwfvFJ1MeBV/8AHWWdQZwc
nI7NxxAF5Bl3tR4JFCMDi+cMgrCmndXY8rzuAkRmtCb1ThsMbxL2xEMzNuiU34mNv0CjGlqUU7V0
sXUcYTaOU6DZF0qtRjwpdfGuTtKqSyKzaGbUnDELAHtpPbtwT23TtLpsFUtvFl/LWJbgoiMQk8v8
2ZqFwzMKvpWX3drnQuy+bk1IUdP6dV2cMv/7tXM177/NE+QLBPzxLTlv4sMG7/drIvc2pq/Lfawm
0UuSAYi0gcnCY8iUfWKHH9w0MVl6Xz2HGN20go6DMXvPBJ3jHTmmkCz9+tMIVHY9MsGdCAO7pSe2
YAEOaz52+Ku9NEcZAFyscYSkup8DyLnVEbAcyJqg92PNRTRyBVBgXSdHP0klgaRQB0iltfw/NliR
wWH2MykRdytzv5U+eVAr0Z25JyR4CdCziaiOrU372WIFpYGGiAaIDbIBpSlOJKVXUQ6J8zeJTj+e
cSAFciODAoTw8G2uENaPhfketGZLDAhh9yU5NyMBLp9tOCfCOiQQpsIQrit/oaCo6RMQaoPkmv/f
IRA3p8vgezVAZDDPlmBkwxhMdspJMxtVZYLbVUORHY7HTaBAV/EpYy5dh3Ip1LPoTOxiaHmRuPWc
2FSzo66Qj+cOHUAy7g60Wf9jmcrTW/WH1Y4QcAKwk8rHL/JUxZf7gnml5AplTgOypDAxgCB+nOT6
tDIMKxu+M6m5ZKvKoMCElzTXnOj3myHOT9QkiXFVUODTdILEGSvXYwQvFaj2Hg+hVMEy5OGZ47Zi
PpzAOAAuOqkz60cNXA+KpUM+6gGCKr6Ax2J9ml2R9Ostmvm9NFfygsvVGOCa+K/NO/UHiZiEx9UM
PFqKwHIbJOUxQf8DeEQSztQaFLh0LMSyIZC2R08TLFOvXROpcJsIXC/Ua924gNfu9LpEJzz3oFtN
GMykRycnqtEbX/rxbi93M96hVukSIprDvOzB7WryhjwQy+638uuZB7Uo2FOmZTkqop5Nt83Ltif1
3oYZcUa6wSYrpigLaJmtIB2eKYTqaNiLhvbrGgdFlgvBmCugkx+2KuEPH0sgTheYdOFF1rkhIx6w
Qhgmzj9gcPluMHJT3KihLDC7dmXSxV0t5A0Z/7qqeeFarJN7g1mHyRKhi2YPZ/bRrLNLvBN43U16
ex+PBR9qyIZECZ4XhVUZHqGZuLZ26ghaEvZwliHc7+2N0rgtZKxHJqKOXy9iEYFoI+/wVhK6utlj
7+YAeF9eHz+0gso+mIsuL08X3fk64wj5Bfywu7J7viulFcmhAT8xfg6ko/PMalP7bcWJ5uFBANVc
is+OGHIcyNKsBJjtubct2R6Zr5VcOBMzt53jsdOTLjHAZoriLGxhbxskh4RcD9j5xZtlio/XbU9l
J7rd04D1Iv0pZm6OmP19rMB8RtaAUAcWaz5SrA9d5659/JbhZ0PXy32eTYJ5ASjwhxBIpJ6WVUe/
jP7cXXMx8O1QaTxBdkcFBNV/GrUs5EMtl71elQsIazY29ZnIAFPpD2sZAwAdy7zKgrI8aXegiupR
epHsntYtq2rp1avICtxSc9J/x0Pq7HjS5T1gAJZ4a5H1HoeXsrmSv/kzbmzMIthhle5sNhpQbt0v
ar6KminF1fpbGCMrdwVMjXaQx/pWC3DFcnz6W125t7pVpkl/f8aCTYs8pQ4jyRba2Hr1goRvq3S0
mXTJvNnbj2NvVszlG+JXwP6YLHQI7ck4eK3bz365gRztOMa42MUy/mUXGXtD2tjPDKIrtOqxya0T
XY6zGrWh/F7uVDmcpe8WcE3UViko2/CWlow+VAD6fDFVBWHys/zSmbTGfu0ylkCJPV+Sy4pUENVD
yvr/QIt+77nLCX9SQRFPH59I4j2KUmPu721Bg00+uhw3dhg+ixXd8QC8JOqfVYnDOlMlyhwdZMpO
lXPCetuYUCcNlztk+QSxKAHck6OZUmcyTWznwcnka6Bv0vDBta8mwpjp0q0pY9pS4sXoIKOHj4j8
jURPdHpHqxX4hxMmkfySDAFrDtb/rJqdljZzCktLawG9SwWRnJxyaVbDh28A97WvEIDf2L6ZHQ2C
BfRLPsW/VW3dyPYaLjuYpzVnk8RtVc+OVhSqLNBaynCrH2I9VX+OKnhhYG8+/cKtsDmEiko4nGBg
zgat59X5ayskpxXXrf98ImTfv9Y/rz+bk4NyCAxGPtjdjJMtYUyU0NuopIB8vVWYY4I7am+yRhkH
Sw+L4jDy2y85FdbImERiQFZHyaUXFiqdnc28jbsAGE3lBezn6BiJvMTJWKAq8cjbulPOG/70LQZr
LqAt8DEqF/rZYsQ8SPKAaY/KBEm58oMTOcjEu6UBB94bbkvkd/BcXy7C3k7wV2CmF8A/7lmyZl+4
LWPMTN9e7hV0SodSUiU5AvVXIq5e3Mb/QYO4Jj8odELrLVbkW1Q9NhBqRJLf2yiQ4/7gsUFyGeqv
PLcdU7h6KbF8oQxv1cheSJKSn5zRxY8lxHp/FcKhfUHXS4OWfiCKH+Q6bPxMPIJxoQ0hv/q45cxx
pCWxRcdl2A7tNH5XYRiAov2VjYDDj2/GK4K8GEeWif+cFJDaaRidF5O6rifhfoPHCHacrohNp5uV
bUXUXIuStMPT7VQ7Xmd3s0lbggOFtjgAbqybEga8SYANjpy/22KmOLPyai9NXZlpl9Lq38Y/Wn83
vlqLzcIAS1UfNw1pgBvApVPdtb0Zqi7GdibjowjMZQSa0BP1tIlGPP/GmPEhIVJTZdMX9BQgxluh
W0se/S39i4//2hvrBehFALEDzqP61n/q2xGEjMKfsMb3VF97kGep+bNBmTXF4AZ5WxQO4NKC1Nyo
vJ55IgFfHq7UhFIj63YOQWScVXeyWPM0iBPkh2PP+a8TIEqnGSsUTa17pC2Y+OBqAcaFzSPUyBbL
4b6yp1tBufwu/j0w8GT9zGbbnC2WI7WvtAIjHNZSA1Ezqcjx4bPar4+dx7bwavdeA1nzZA9N2sIO
k72vpa2N/EypxdU7eA9hdWEsYisugnQ7YrUxKYeL7w7eCrgzTryLtXQB2o6bA0fjbAXsJxzkiXse
VrW0Ec05RbfOaqOnpHG7wbnGRrWcPcJLwPmtws+I6krYcbWL++Ym9wmd+g2VKER2okaLLJBcq45b
6q2TzajD6G8Pd4YpPX/0vyAmsdTQhj2DjOlAUDtKDk0F7NsAuqAJtVX4YazB/3J0zD7FDGynJsQn
5co1HCAKq5ciXbuNwaavxFaRp2XVm1H0J8l9oTbKBjPIMqD9dJFfYXHnqt7xusE62w35IJ8iaC1H
chf/ORInPQ0N9AQEV/ywtzjNyLHQ/b9f8EEkr4UrV+fndE6S0TNXRtJC0Wpk8P1TPDUgfUf/OBY7
0pfQQsqBKYSp9LoJPJBEwxR+wcHVOcon33amZlC2GaEfTfWvFUO70vxCp8V5Z8B2oGXh/eorD8U+
gkT7IATIZQwwmkKX6m0yTc5ItBNUb8ZYWdkGM8xTUXBefdAC1EqGYkNY/DAZrqJv5vYewq1wOIWe
4gqs76iCxBbU4QFG49t/av6km/e36lo0wkIl1c/Z7Xuu3ERJ9Mi3MvUhD1sHnOIBCXZWYwDrq3SU
Y08UPaXNS8kZxUGizOfLdRLql8evMtOqzTnSkUkddULr788HdLgOmuGTQ+pwDtS3LTw+1hZC2yGV
wRAtN+pN29NpBYiqE6Qbyn2W9U76JSu8q1sgig1qMiR0xgIorXKk/DbcmcnuIwn+6/TOhzknN6if
rtVbUpYYpvpYpji5l8KL0MFRKsUywKhp4KRLHmFzEVip2Ub6GYp7plImx6JYyR5+kHLfxz/kGIDz
C8ijp/Dg4k1cKmQjWrpHYfGiKqE58t5eezDucuWCeybrynK8uyD8iTEGVT3Gday7FDdBbhPjXvFZ
eix49XnuxtGWM4+VWJl/5l+zi3120lpRoQ2VcLMmcegpAknCIukT5mfkzpy3f3JV+RC/qXR7N/VP
v+HRGdsN/pC8sWXqfWWaxtk4Z87UuwnYvDb3doIubRfDYdkixObZiYExb8qJtfqiEJyo1BBbW4XF
DF54A4EwO2ahjf+E/awTdzySKhAuCSwUa0Td1uPwUI1I4gTkHdeNaxZ2mttQeMenwADM9GKRqJxH
ysEEFXhANxfi+4igIU65wZQvnzqLLGfWyFCLSR6d9LXRz+BeztsIXAf+X8bi+wHYvoxF4ZEyCqzK
qdyfXLHiecwGKtSaET8+4VH4YYJ4RcjWSS4CzSi90B5vksvyg1uAIx6x9SxlSTRAu46OV0ZKFWnO
BQENvWM/GCzn/BiE92no3DfD8A6bORkAW7L7Ie2YsD7w37qUtxX5CY4pedmBt/3ntiR0lL4ZwkO2
iMez7mojpZoA0K3m1p4kx3guxyU2PAl25Y2BbJZ03X1sipGmhrTdhqb8zUq66IorTp6RTNakMVs4
kleRnOpxk5AF20Dxa461ej5HRjetfku1h5dBUw8nZf7KeB6tsCfnvPDfGsk7odenX7a5bz/HBaAC
f4k9XN+rWoPSFyNCMV0L5qgxJ2vZ1HRMHvOd/Frm76fmNXVwPARMKzLK1pwlkXe/raIuV4OV+FPq
fBtoM1VI3Cuh3Ly3bmDTWrrEHU7vAbJ0DQ4JTJsz4as4aqSTZV9fmJakmlRQjhU1DcwFnLzpTYC3
DzMpB8YtIj8cIo+os7kYx0QD8SLbwkcUU0kekVqoD+JpKELj53VytO3StYIOt0af6PIx+8MnA83v
E/vEca2Jt5EBKjo0PIEIFOF0h0AWIXE07PIb6plkYnnmxwpgc4c9D8AjUaFVtW/3sYbauUM6EpuI
7BfQVTb7hSjb5InTmyUV6DbRNPShrzYVFzTR4ukfCxQMNMxqJsvwezQ7i2pqkbLc6GH8X9pRrKsW
jMwPl82BkbU5EE/t7YQ90/2vgYpddgN/oiiEsWxynAVx6d3LkdV7MZ9dyGwbAHTjgYsv8mZ7DsbT
bP5U1se+m6+vVgAgzCUrxlaWzBhVUG3fV10MqmA8rIKJrnKEBdIgiUdwQOCCgbFAptButPYOcve4
cu6pDBjpvKAq7C4ng08zFDGET/h8128alFVQa9lM7HMPtYZFAQwK5JIA26rIMXDzOWPVx3uuYlda
MEtIs2N/EaiCjWv+494WzPMltuEAzfoBhkj3pkqnyM/6UYk2mhk22CvEEhx3fnpxszvQufVfZvjp
2ONOsl0SEw0P91DfLuklbIxWACcaMiiEnyHWKAYQbTE1luRPoZvSKvOmsQxfz1szb4fD9HgCmKpg
JB7uU4luHR7HydBBCABQi3iGj9IoB2BpQGEKLUgMxmxJ+67JlF+kAdkdTg+Y7zTFc4I6ZtU34God
5/HvOFsfmuze/GUndso5tboI1+0uNrv1jSGlp/lcOomma4rGN3tpmspyabz8llWHFELrNHLKOtWF
tfYoWUjTF83D+y9eD3l99ZzNO5+5wRn1vtn7+wRi4QsnXLvN981BiA3hPKY7Gzr1FdDNBL1YPm0X
5VJmZ75HGdaVVXLN2gfT0Pr8YEPp96HypDUSASpujpVaOZVr+nBNGYr51kgUmbsBJaSzPofec8yO
FGb6d0y7pUaNw/IFDnxplTsRrYAIfyg2dJM9b/hS7Zx//Ko/fzciu1HBK1PTaf4ZFn2GL2C98kHW
WOH3gxraw+0+PSmfP/1KXCfXlvrIkQpV0jOG64Tj2fyizHV03vSiSpcUyhbYfu0EAXz3iP/Besnc
oK8BEkUK+nMm1Wy1q8vTUyX+nifcwFrLjXrZRQs9lHfgE5GtJsgtGJqtyleJ21EEAedLs8iAhNeG
PHfJItFeD4JnHRUlFBti/BlsR3WuxmShHRKFt02SzQhLltF4RvjDkuCOQ0tGwpVficTqS2Jz/gkA
WswJ22H+87++USKeeBSCiO/OGK9iY5fltFcH0HOAM1CKj0uDu5maRhFD+akur95eWWItXZ1162VX
Jx7ANIxJYoLUgOw65hfXZj4WFJorlTHMiZfvmxHZIX+3QgzdH+xwgUfwY30Ahj0VdD8gkv/7UZf6
oAmb3f0pCnmA70WTWagqCSdl2JgsY60Z16Tkf1y5oryiU2dnycnW0QsnlH6wSR1EYY9T/cpHXw2W
4g9aMT7xq/sFaJCpqXT5iexEcjJonywiwKGUZ9sZ5zptyX7p8Mgj/t+kqiCn5dTe+CTTriu4IdFu
KQs8+X+mt29LkBaFy0d0ikqbhBEqXU04p6UNi41QoLFJu+rqeSngLHuVwPtpQajoE2YXl1LHkXY/
qYJvWoKhUTv7TlKjeA6QBOo4POw+A5xSkaWlxyPlIZjSxKToHB9sVpkdaWs06Cino2oNWVIPNiPt
FeoP9lXl8oiLVf+f6GORj7bUFzTmXTMoYOkRhxpIZ5AdbwDhjo5ZRXiPgMyexwrnjfwEZj841BfA
pG1i79Ki2LN7tCCLRGqS87rZfgWmg0df+38aU4Was+v4TSsPVd+4XkHcL+EAgFLvHpfjId33RRU3
Cao5P3pXa9okolJIXHZ2/alr9AXQb5fz6fr2jFdGe5Aa7YznRT+PYK2UggUvDzhFUJ5atGejL8+k
QA5SQbWpjodfZ4vDQ7+bFOuXHZ6U+1WPUsjQLNOHLhLY+nXyDkvfl6AJrtuY5AWiLxdpsQTbekVw
OWyGneXi6x8KpbE/vKAtZSb5KwBCGEYzR29JPCF12Lt31HCLh4oFVyET+RAZ3XvLrdYfZdu179Q/
N29yvVZ5ZZI0mpelrsuOg8pjyQ0Ijozox/8rmWd93BrVwnwEerIwXA4RVp71h9px58X4VSXrz5TO
CcZpgrYd6kB57vzEypG7uBSeTu6b+x8yg/Q+QEOKks++htbooC5tk7FM/JX13h9rNQMPUr2Ckn18
/fFwarCN+ArHbCCaV8yEUyq+eOjLd89oeiWHm0CTnOt5x2X+BD6F0DmPS/RUYLok4XdDrC22kK85
b1WW0KTeT/JQvVMK8tE/Q4GBZWgTFy6yS3QnkC6EpM1JJjyDRcVQ6yHNaT1+cGMQGrcqvdUd1xnj
zH/3CtPwkWwsfpB8ebR/gv0h//cHRc2jy/pe+j3dlhnuPJ/cZutR6ZkvgjRyd666WPq99VESVptA
EzbrZIwzovMVdZdWEibFaXAX7fAkUmx1+M5agVmE9dXk1NTgYHB7blITGLsKa1cHJ0zOmQuKSobn
cSQRe4upbghkD72sqTRkGgZqosL0d366xRu3swYhnSpzmymR/R4WmH2jvpNEpJDoUOrnSwFFk0Ur
ZFPczCkQYfD6XIa/caNnr1sdR53XKKXIRPysbZuW4ac13baDQFlNIcXtsBAnYc/MRSxj0NwU9BVN
+WH4DoZuTsD12GhAybaIX9WmxPIR6Qjg+F1FztH1wEJNHhNAoEljFdE4N6AaEBQqKwtwxvtKQlfb
ZnSqNBz6L610gz+b1w4TGAzzcrv+Hgn1MY6ntr4QfBRN5ncn9O8t9IJwzL9VzJ71bh0RxwXSz+6Z
8Z4hILWjC3d40zxkjt5X8/p171fiaTBromyJie4LAmeHjKOCkeuU3b97bqK9VD8V75IcoPzkPmSA
1zsyOXcyEae+s/F44OxoDXrO5lz7CHdcEFVuVhapSPLLSF/MTQCGFUMvJB9v85mMDIg4KXwvmsjT
7RQxCWgQ3+pH3/yDb/XW/xPJwbTbdwweqCWFFvpWrBdJgA2qky1sXBi+1OkAMm2ldUWlVBK3PzTd
9k2tyTN93a5Uy7I/6Bg5dO9dT5bCuTVlzM81J9b9w1luKpkp6XCJvXplkFsA3kDrJ2dk1VH0Kd8T
0ib3QO6NFr4rkKD4jnOc5FHUAcuL3jE8nW1u4xRpfPRHueW3EUosaeZ72GZITszwToKAoOd4upAD
1lWXieZfCZQ/EGULVVGNNli1gspoXMblXw35h7lW/mijlUSFjtXRTCcRZujMS+CIxM9Q6p2NKFUt
iLFKDK8r4YtWVjp+kltTFi8uZ4qXqwMrnlK23TNBec/RBobuKBYLYlKbUHxPQxz5HizgmhLQJSVn
9i1vFz94XC+nXOC1ewo4oGkMDZgHS4BSp+ZRye4qIEJelgCnLWxsJIPOe7kIXGOX7/LqBBBqOZHi
puJVSIaI/AK2HuB1GvCZvBYcmJRahWugtSK6J/BYw5VJZ3wsdhWDp+V99y0ya+tn6YEtTyw8ikVy
NknC0R6vNbePKXCX/XptBwMcqPAU8HWT9wTplGJzGBp7Hyd9haqRG149gZyOzZBzPoIZZIEiA3mw
QLh+YyQzrG9iIkitLgpiWTgz97jSafhcOYaNNSZyoVaJeilsk7/HB3uq82ksaAyTS8I0Yb77sx/e
9x1u9vzKeOuMsfFXj5E3E8+zcy+GdNcSdFnWWOUyYHgxXfDhKm4/XhPETn/RzzY48Vx8AJkfSFnU
kIXH6DgpIbCyABXRiGv+RquxtTHzWMLp+KdeSUu6RkJ9SmudElh/oeyyMo3+hyG1RpDWBzr43Jo2
3K81LNbcNysPLLCXIl940EEWbz3iD4yRXyiqlOegwSghLoiHUIhVQ4HIQAosb1hhCreYMMoW6zK3
zlhToeKJAh5uBbDS9bDzKEFUnuQCBIsA7/UNuDRb8hDoxDWAkAEKzfIiuJtKxUL2YrU8uJZUKs0B
YHw+7M3UNUnN8inCN5sRd8Mie7lJXxrCibKNe4/l7z8TOaEQdWs/KDqnC5lteTYQz9UncPh+ZQxj
DoihiXbUT+lxtDn/jE/TIEgOnLKEJEQ+G1LHZNR3QC0Jq2XIaqc1PIDAJvLESi+xo0L0v7XHUHP1
havq7jwIyI0pygnDMjfoq8kx8ILEzvH9k3JVsy9r0zZb32+O4YUwIxyOnjdaOTTC8u+nb2p/9xTM
q6IQrvO5UYCirDgVAy3KpSKX3RhAckHD4Nle6e4kQvdV74mdDNta4Y1OAAtLBKqzi30HWmYkpzNR
v3BYj3dG4vCfxnK2B72n7xdomiR/rC9Zz5t5ZLf9U8ieb3BPAVTAXSHhw/b0X/GjQeTp3d6H2zqv
QDnzJEAazx9NbLPXkCy/Znct5FQG+GtT2Gs2bhSbDqZR2+kOEAm+zHcZx8P8WGVKKX+uKNlXGQBH
hJeHqsYpvqhC5Ghovv5XXqpwE3o77anY5WNgE3dO+iFXZYadv7NBWLnEU3nPsE30/LeaSIw3nkQk
Zq7jWNWjeljiz/AR+/I3AKxFvZoVmK1Vremj7YJoHQdBlg1QdQQAfTbZ8VA7Fh+/HmzPpbrIVZDz
yI0FWYi/9TiLTrltkAVEO/QouTXAbEfSAMy93tJym2hWtfmoq52bmVEv6KA5RxwHe5Blevprmifk
O5dnfJDZVBELmV0RWZ+vHiIhSefwGqq5l1pXv9ZNbCKaXvJOf/8Kpz+SNyAGiqCSFhVOYjnlMju8
FqJNSSvZY+hIqqiexst76TC2Fy5tts72+8nzrMFO1rbDk103YauTbxo0NUuj/btJ6sAhNl54Fvv9
xpfYGUrV63ULjJfIULNAatuvn70nOb4gx7tiDyKRqnhhqOnMVYwO2jtyc4UO4ragz3ceWslryLxc
sZsMtwEZS41kMKpqARGyYINGh5YE4mph13GLhZh32AKmYZe9UQTs0vs8zr14NTgvUL9Ch5WTmWhl
1OhoCG7pVyJQuu9trC242WxW3uxz0OF/tgkRk3nokjw/BykCOqSWy7ByIUOba+8zJyjinvvwt3rD
z7RghPWyq3Rw3Bgs74Rr0t0+M/HFv2Codck3M0C5s90kRRhnPyzYso2DmQIYE7N20Ss95t9N5meT
OvFVuVMoi5bVUA6cyKXU8uodDzbOQYoQYrT7IzAkJevRtwGxBVPUyntX7A29nw5epyoMspi5v3Qo
tGg5La6Tg/J15FxfxfYMM9+FWyelj13xbWIGybejBHuFMUDGnAULp+Anp/YuZgTtFy6woMUc+sib
geR+zNXSQVefAfptGnMCZSj3YcHv9lvCuDnhIDMuZu5BrVpf3zS/dDC53ZpawhlsLax95PT3+fX2
WU+kUkGyo/T7RWflYQyfnsaesWME8Zacdr7URPZ1naoW2RTJuXpriJ4HsN4xXVNI3n/M1bL/Ds2g
UMOUVUNEKvbOZwUWitvnKzsjkLiLD6pcLvXk0M2pZoL4q4FafgrlNYu7aYIs68L3cCK2dwM/cFlF
bk5rZsORFtZBtWz/ooGtiHjrwLEQx4HisPHReVbfnlrjD59x7ADTAAUGCHuPIpgE7qZc9iORB3ww
MswMhVu+hH+qyzECIyRtIALVs2xZZD51IvgY7ZjIwj2QXHhrXyeGmINc2XDk+QkyEfkIxClGBP53
SS2K46eR5XGVZu/UM2UOG0Vzbr7b+AaWjaa0xoFdUGlgCobkCA1VbPqTIknmqtuyEdhvlXq40xy6
RJBYx+lPYPfjJe/UG1Bm5qe1WyHNtbYCQcMFXhbuAH6qKHUEefuwP8Lscz0Ubl5hAO2eC0nuYUTY
uZuCTl3acj42C1K77MGiN8F1mjEyrJQl2b84uL9MTmdt0oAz50AIPHnmzWRxaC56DL/GK+lxajsz
QrD77hWupXX343JjRH1IdANOzoW/1njXhNKk2TYB6JeLDUyCYzOuFAaV+m6dkcbm31NPIjwZOScN
IRT1A7YR9e7IxJxdOxFDukXrihT/tLqawHPzkVhas4V19AX3pFeVz4WXomp6c38DHqB7iJTQy0fd
OMLzlWljxSA/UBbBO8jY6N/H/gyU6OlbyjU42o4bkIa4zot0iSXdBtD2vFm98IJ0HFS4ozYfPk4Z
WCyv2EF9T4v41yXa3oZbwdSZWzFnOZ+BGVWGtPUZCwsM5vCkIi2O0x5AePGiXpeKdfZjGR0oB4du
2+r1ucD4fqRMQn3PTE4ejZZiH9d03MwGv2/mEeg4kmY8V+zmjFLYC3g6wQriFLjRAriDm2/bgkbs
muxaOwzP3Ccia0wd26AMTOqwQJz7Bhq4dlZ/ZF7t9TxHKFREqOdIy28ULPWK9D+Cook5iWYVu9RA
ajgo7nPW6P5oPSf6tO1uK+c3GqpJ+R7jI5FvE4rSMNuejrZx7IuZZpa99A0H6PWgiBrdE89Qpjx6
dHBewA2NhcYSI2PBp/i+quTRfdhZASOkH7MCq3/HELVCfemLSgtzSF3mvkAmPvv9SSJ2vhMv3GQi
Vkc3MrNBKZx39P56LA5Gxx6nRP4yHP2HNueStxjFQ7UM8a3B1wDyj1RqcxsSjq7HsK2Qwyum41/G
g+BTUj/KGkLPn0huDwxu5TBVAGUbWxGhT7AvbmL82mpccqPZMxvRIv8ClRMCZN5hDFGQq1HyfPd3
yD8yDqf67pLuqEkGb7NPXjehIjVU953oSBzY11du7UOrsP1QulYnWkCdHN6FzxgLpRb3cWEhjJBV
QxRBRdrAVhNJVL4u5VO4N991i2S/OQTn7ZAMv4EN6IjXDu80YcOgai/gKll0y+olDa+Sx+X/QAva
wXuV3YFzrcFlvFdNii0xGWu5YVql686WvrvuMhCWX/BrzWvHrJAJ4VluB9FkUOGtonhdIqkMdjYl
Ap9QD/v6UEhrfQXRueJkYqvXe7k81amoMGARgDic0gEjR/xx6sgKdrQ1cWKGp0EpXoKc8BsqB4pG
/wSzeWDuzdxirFJuJ5w/OX0eypcEMFSEGmsULQt1OoRA+0MuzjM58kq64Q5OG/Q6yY/Fci5rxhBH
7t49qe1NvlC2niUmckKgp1ahqH5vfTNPAbMuvLZXK4FfYze3wsCq0oilp8WtITuK+3fFPVTF/2ul
Hg4QVNM9zBMLllzGheSoBCreHVpdR+VzRJQG3VVp7NJl6i+YGCVS+ctoPAOOeFVx71HDofbsK1xP
q2MQPNgNBBVXjFtRP9KzJmUplz/xlDDiCPCWMu+/3FNFVG22tlZrFMRfOFSzDKzdlef6C05xs7TY
XeFa9+kdcKjNRaIfWfpBITfyzIWx40x2CqxTENy3fnujYtYG2I/giSu/yV+5Zczg7rL3Crwrl0+9
F1Q4jKJE8tPeDgR49IlO4qe7wSvn+aZF3ni+TNLG2j60/M4LnGhUsf7uWdEalOnYU/TxHjKJVhBY
qU+qXvTagSECOp0fAUL6/AnLxCKyOFKirt5As/J3zdlzuLMIwhVi+PWndwFSB5McCNcfU86igqUq
uUZIyOHBVPVfdQn0b9Kn83gGqxBN1Hfojvmfoqidm9dD/QwotJo4+v9okWBxJdJYRzZKc1Gs6lQ8
U8AbVs55i58mwC2l2MzbmFTjIqJ53xybEot/qJuVoJKvXyIbbSsbtB9tR46NGHm84vhKIurmJEZ9
kuEKzmILobK/S/oG9LaFdSknsxinT7hEpZ3gVPzxd2OkBNL9x/ygtMB2mGXREiBYhLXHqltqXDTT
vt4wxNrurynuy32JGS5uqOVqP6lOo7MpurZDwrxTWsaoK0rZzd2UvlBGIsz1uFKc2eIKGzeH8fPC
2htY9LK6emsqgYd5XmJAeijlBcidLK1GZYDh1a5T36nDK1TH3+cWEyddV5FeEGK/qhytSsBaHqrj
jws+UaXSnlc/z4i2Q5GtCXjm/yWf7ij9nnMEofvgUXJgGa0ZO7W/CLS7VT3D6ib+yEwoIHcDgT+R
pCL58mRAsUr5hA6bGm/qmMdvJi/5u6eiQJID9hVsr7DvXtUUWHRgH/A9OpEG/QJ6dVeBWa0/MhhZ
TA0exk7vSh9Yk87w78mz6esIzXnAsV+Z20sG1s+3vl+qMIEz+0+eYf2SQJvo7O97rEuUiTCKb4Ct
7LWXT24V0Uq8nzKZVWP1r+rxGgOpZpO8k8rWUr1ZSshUQ8U2odne6sNydh2f6xQm8U3gJ+CXnic/
6hLDhe9sViElmBV3wYocJrRRWkZ4+muRxIWyVSuEdLKpUcpFsVQqfa+m3ZAqqYv1+It/qizVxeok
RW+d2g9rctq0EuS94OVgEbHsl8HNE2Pr9OqVa/FzWkMkiBWt7pSwA5j9/3uIKNyF0CCXfVArTm/R
uNDpq5AzqX99Ep7Zli7Bqu5nGlXUBvvbTpjGv2h4/Zi3QPTbb0oVJKvgwMyoKpjQ04MzqaKDG2MS
ZekrI+4LEpJx2EOrNKZcvgYao4TcZvFq4zEJygdzaJELsWx/AhR3xigGj4WQc55FUdabOzP3e7i4
Sb4R5sK/0jB4q10mULgpI4Xg9k9gJaSZzWQ3ZXIwPdyP3iS97x4UrTESkWqRbm9VLXRc4REc824G
jehhRMcmYQtAVXGJMBhmiTfC+c4s0FxQVxapyQq+xzvUvqI3QjCm3xVrZyeUZBChL/wc5BbVBkTG
Hj1vnuKg5i+oYStIhYYIKczo6YlSDzwsm/24R42GehLMXTJPLIUoN1xSHyvRak4o2mhvhA/2ttxu
S+RsP+8Zd6hE5Cq4tCiw96PfpxQxoMEY+SX71d1njHUUO5AeuJAYmZIG+G/8uySvML6H5AlaeuAE
xT4V+C3Jpuct8QT/If9ctzqPjPi+FMCdhaMtLve+wAMbbqu12Nwp+v1tiMyVMiTHM877MWFk3sKG
+vNUnSmMfg3ziijluv9rlDXR1mGbwJDLUa2/VmJqeDVPw+Tubu6EQqNG7aGpryvgueRWnH7irZp+
ZDq+LAVOdJEKNBhaK2U7lX2pQB4S6YX6KfQjvMeonQX85uJPGncwE/r3OsaEa+y5AL6ZQRw5BkTQ
FvfjKZsI6UoPgccaGSSSOuFgctIx1sdgZ4eODHlF+2dM226mgvQJf16JulBL9obEyqlnnurpMeJw
kiELKqgavY/GIll8VYLctuI6zYjYBEo2P2Gtp/+ShanksShWUwFWbBoYPTi4wx5gG6fuagcZvlyR
XBDhF28aFuH4eHOMgBRQvdbZBX0vpRp5STITuu+GgTPLlul5oxV40PE8f6w4Su3IElTxGwrZroFJ
syVUWZrvOX2TtpiSQOJNInfNGvMDSAuZtxAE1MEczyzaaHY12/IW69ushnfNTXojidOthYZlMvYV
18H6/tkObtMBRWM3mNvxKua5iv5PXViOzfpaAlK9zI2JY+iFkaR8hzksAHFnQaBXNalhLQk5oKil
YBuk1jw33tt1gWa0sKd1KK4ZMGE5ODeNVB0h82LDtkzMUGBEk2XaMPpKfqjplrUVNoYkcaOYM7yV
nccEI2f01hoSy4E9RUHK7w/IOpEEMWyNmBgoXRRuDyvOsAWUCsmPDuGr8VNjy+h+X+0U29Yq3p4v
7t0dgrI1iMov++5X9ZXFVdrg53YbSwLbj0+dDIMDPquGoSn2vAPS1yYV87+8GNa77MTJsImSQqOY
p0ESi1TtNJ5ypsb18sqRGoWFFsC4+wOdeY1YvUHkutzyeV+2zW+nbwU53gaqQOZJCvNT6YKHocKs
Eufv/hFX2slYBiWmFcn0LtzsVvZJc8ybOY4igeqHAcFds97mWL9ReaLbCTSq83MURQl9jMHIgr7F
agxkwGMKaWIZ/A1nVthkYynVHRkACVxLviGLTpmOKOGOyO85CZ9r2DPUHkr0Zb4H9g79PzeE5Tr1
DaNM40jPSHdqHGxgX0Twx0JoP/EP+kGKITrr9xAwI64sJhD98IN97PkoNbtYInY9CNpTy2jg69fH
p2VN87GVROLhaL6Mvs+Xx4AgTQQwqaiPm+3n2Bpa/BIrVu/9PGPXMHpXGYgJVTi9Y1Rdp44q+o40
iUxp0thFM24TwL3J6hbGPtpMTfxdCzk40WF7vUWIy56M+NK/jnhTMW+3EJ9zacZ6uDr+ZDrsAKUN
rJFgk383InhlhP33VIWz+9FCkFuydy3hDxIPu0ykU2mZJP2hWK8T0cLNOeZC4jvQzkrPEnw734Yb
CfZ5p/Wd/oIVY/TSYz2IGJ5xgykzzbTQEhjkxn3Mjn2D8jnEwJQG0EWoRxv58hgME4ar9fJynaTm
0kJjTaAKWiWjqXFi0sedAn8FquiNH4z7Natsh2/ex0QvRVKy8+cLwLrN3Iem8AltmlCyc2G2BbKR
hf8Dno05zxaqMWdsXAw4LMbjRzjL+NjiDl+dqqgl8/cSl2SqBS05BEWMC1AMRi9giE29punYJkDc
xyMY+C/qRv2eG1w1FDjG4Im0prAaKTQ3Z9uoJHoXvFWDEqRq7DkYVGgPBMSfOTG2o9RD2mrsF5Ty
YQCk4dabCEM7PiisD0++s1QRIPMhppnKbDmfAdNOywcnHw4AADQMBWQVZUVuVorrlQ3eUC3CejHv
monOTO0++Q4ozE3KCg3Wd05p7DVIdKad9CkZXlpWAuJrQXJr3vbZ2IXeMOMjoUJZU6Pn2yJj++Qy
WgTfxlKU4IEDxnFREWmY8WkG/3iYDDh6fvxIXZ1UtBFdaVLOMthfahrn4NBt/BMGBaxvDyda4PpE
Nin8Fuk/hcqnMuoMWucvmqjIe2/Ulq5+K5Otqvs8Ms2AmUbvoCu13jov3qwiEHpkmbjy6SvvAXvS
wOCOWXoYjqnc9fenMETREpBNuQ73XOc1xDtzLvW97dIIaH+2yus6Tl+BkF8+uWCiPdMQD7cGaNtL
4BjFG+/kK/T/fbADuFWLO4OgroPHj+fkyC7eTob2NtGBkIHSZ46XK1k+zXNZY1aDWSBC/jj32nRk
q6JVMULhEky3dYPBzDP2w+kMY62LFoPp3Rgvh+gKYdK4gZ7fHzqaJO23L7K7+q5OU/aEQ7wmrlM8
it3BmDycXPUNxDt4r6Tc2bV6zAMtEfvQ0yJ0/b25O87/Gx04s9Wkp07ib9RBU57yKrdFSOnWbpCB
sbGT8jcjCmEEYNrp69AxRz2AWuOC3sCdk8rELSNW0C6CFHedXpvL3xMWH45QoSeodbn9rn/YAqRo
+1I55knwzO9IqXAZcCBs+AaJzb3lTyZ2VB0+loNDQhyC8iQDQg9FMo4jViKfwc++RFYKb51sD0It
2lxiT6phoUM4JyzrIc1Vt/kRdtO6JZ2NixDv3KkEbO/T38mD9qdMB4r6JtcQQyWmvtEyKIvGxHI8
DR531BVvKsnVdhztXYyKWN/UpRtypytifn6lpiFz+Uarqpw0uHh+JVHa2FiRnsY2WjUNImKhl5iC
G7do8z0kp3ERVM1/qoWZBWXgNFdUld6UJfuGuwyRuhv9L/IRuiU2lBEKQ7P1B5S/M7XBIOu0mlXV
a4ZbwQgLM5tVkeuMJC2gzqFxjhYYhc+zqup9Nd19DfNMizOLQoBM1KJq0PvB2KVGSGsvQe77ibw7
7xGqVJFwdx3rqCfDNpcYMt/9mMrq8M2lJR0DYJuYdiEeNrU5EXE/oP7AmHN22Fz/prXrlVkJ+Dtk
KE5qsyVvBarKmb/Hk8OT6w/QmS8cIUOsaPp1zi+9dziq3OJ6Tdlk1uNBBArbl/BhjNvWOSsnnHvL
KHeUtoA1YN1pGOqoZnekchxW0KHlh24I1kl1t24CHIFf7tGl3kDegwYhTR9bj4drk4731G9N8R8C
kqX0QC4AmujcjWS0UpPFRefWhS6efZsBOlkF7AYBMFrsnNR9O2AckmSmn4RJJaSecnC1x7TkwARI
eSrT0L0kfbgCW8vQTpucoMyZn1oWGECIO1Py4LwAHqZ0i4CqvG9lp1Wegd9fwW0wMkL8XcrZ/fKk
Q+HzaD0j6pB2/ltGrNiLBVMg1FsqLqUTdQYioNJ5+1USQ6Yibd1ZWvmbsyg6P5nWy7ROPGRD4as0
kFuXqTFPdeQxVdmiqkvmsY7dDDbFMHjGK+gH704M2DVVLz6T+QCQh6Sui78yMEGUC4Javlh+xhh6
0RnzjkhtBg0cpBolBx8EalAXJSxSLmXysoCydRyf1hBIzVlN9lYTC2t/KE2JKp4j7Xk3Cy7R/KBq
tbfIO7cMBH+5lGxYiO186CcoJKOiDGYMHoCmWoymDATnPFf001/IgzqYRcOuNXpGM+a4KS40wa15
LKL8CGaWuoL+B1QoQrZQRKZh4MUE8RPy8xU6pfZKinJBCkshihhdQUZK+F+GkBUG07cgc2cNxAwq
/Rib40Zocx3pKDXhWDKPEG8nykA79OLWPVvaZax3Kk+wIf/0zMCTbS9MvykLMkt5XfRELyqZ6DYV
6KtPgleUBdCwo/zp3NToUNPOSZBWzL+4Fd02IR1LNczYez4IL9zUgFy2btdhBYl1Vn718hUu4QI4
GnorckKV1wskBR6R9tE5O/4zj2wZp8c51OUV8LxSxFN0ZcUuVSunfREGqQ4ZZ+a0yYEhpnoGtRij
QOOPTGS5m0NFJrrKcVL/v1so5Hj4ol2wI/x7GBIcKjuBb1UDktKFEBNxy16qMjFEAe+akHzLmCBR
qoA8mYZixsMSjQljKGwC4ssfdJKQ+/7FCSlXqXoIKgRzRFx145rY1ydLI1Q5Hv/rSBxCXg0c1Jma
ZMEt5EWuyn/z2PXfP/O1K4PbNAieZBYC+h2kY4pBl8Cmu3yDMBQTeG/GGOp4CI8VvYXji6SoW0QV
AZtWCC5ogSOBoqNsy3Kg2XlqXmTINcd8/ZpDFVFKmDWq7172sGwklBqVoOblPR1OV7v4MStyCIoW
GKl5z4adnDIW4QdunL8HIcaYUOmZ3iz+ZCg/mVSJk7HH7rDSm4Mb9WIL8FgCHtCW5XGtQbtbWoAI
wSLHIoUtYdgey3LIuLyJgdqSoYVBoRO2buhOF6UTzeK3TXbWdk/TlqDpFx1V1MeWD1/zmAmhDILH
pDQufrSXy+6shoB9w67SOd1FzqjpdRbZjhGdySpXbEvzvVxE3YlS3sbQqxDlGdNkzk6SdN29lrVa
LBxDvz4F/IZoJQ7y5ccuLhK2Ri4p3jtaFJVsLESY0cLsG924e8eeSXolNn+b8rjeQaWblNwXTGJc
oZIKlX7cRnTxz2uOjtKATxZ0LBMK8Xi6dl+IavxBb9/Em10rO5k4I4mVNHTEWlPgT2xEbfXLda8c
x/6XxdjRAmM2D3dY/4ua6v/dTw32kujBAx9rN5Cn2yVbvy1l5j8/O/nIuNGXcx427rUb/ukbLm6D
sINSfPwQXW7inikcDn4w42yg6kOKHFKN7o2quRqcZQzBBhi5fYdjjPw43EhQyYOZnV5p5hlNJImX
FOhibk0cdizEqToaemH7LV+QRrozA7x0DWRBesiJWlbMhTrxdlVnrQUhIv65gFo9jSGn9ifl4GTZ
Z2gbGXWkC1XzhJw6bZzf/Cyu4npfKzQgGggWCOnhGvSxKqa82KMD4SszRe8ZmwK61vPtrM7rXEcU
uYsYfmG7w/jkVBrJPqpfiBtLRvqvktCspNmVuL4x0A+4TZHH5Ffq97KTw1QfLDTGjABuz9ADAWhc
WOeoSpPBxf/LkitswWDLOhc6VY0svKe12mjl0BzxpHShDoNQV3eNm22/KMwZldi/+XYXOib7yEek
vqOjpujfPjlBWKLCchbGyGNyKbwjWYziwJMoY17PwAEaOwPyWQ3j1CqZMP9AQl3WK5kkFKxqIINX
FF66ZD5lN/U1qxYm9+FUPcZ/aAZGwNQ9oFkEQkI03YMBMTq1pT/fV8+5d3v0EM8m3j4BlABsbvkB
MFe1/XnaEXqPA7XRa6090Qm6pFhJd3cw9op2tc8xiF34dwaXSCPF+HVfs7l9tg2gTipCcdjX/q71
S9QoiYV+Vvc4cv6+ZkG2leWjiDw5XFZkpljMYI4fAhdDEcRFVC8fzqCM3F2PG79yXWOTRrcDl9eO
h/WKgouQdt/zS7dVUlpQ5QZTan7fg2hhINuoOyxjAAdaDMA8d7YnYzNEJXd0K9JQ+nfmEg/pI3cZ
YomDQPoVKrYeSm6bRPDJaqQEumUG67k8Yl+BXMXXuPo8ee6GCaiYLxrrl984bgL8vu8cGFaBGEAA
54EJNnw4AIMj7LHoAxDcTuDYYEOyh+E03Ye8TerguVynjtkpiJAlNS6+Um9Z61X8fezYcjA8FWol
RkF7NojjNw5WLXt6AHmNdBci9cd0qhpZsDO3jvJuA8naNq7LFNxPftBg1Ukid+linaeLkRzZ52bj
dqplf68VuJVc4OEdTJ2uk+D5GEEg9eYvUB0cWpMkqHxl28oRXZ9Q86uLYQsMziSn/b6KzO5OvmVh
GnDOU7HqOJITFAvq53swoXKAgsassd5zeNDX6u6CIqQiC9Vckeyu7/42t4V7otmoJcX0V/Ay3RsV
O8bq2+QT4mvBqlUwwMg8bIsLuWf2reyZ6Rwtj6H1J08osviG45W4TBcisScr0HOVyskh58il9oKK
NQH44/EeYaKb+0D/dTwGmPerE4AGJ5T0Rg37WGde9ae351iGhVZ+5MsKbopOeu160zI9435wd6ff
Dz3Zg+FrVntdxVxjAKvalCqjMXj2fl0rQ6rEeZcS/BQxY41G17Nlbw7+IOOpaQf406vFp+K+ejWE
KNmuAWzJWugpzGBGUCLCibcLicQ9dkemiiUbBbAXjhVpv5zIPc9eWbC+8aiDZtzzedYKYVVv0+Is
bWr/D02LzKW3LJSTkTfRqgxU5Zjo7UYHQNwQCQWgiUc3R4aqb5AOlHL+KIuUD1DgHrV1IhwDZSgA
Jvq1VhZ56+WSFVQ8rB9WoTcP+jpNitgxaj9+MFEalFY1cxLeHQLvWpYDpEKENOz1u2v1hMVC7d+2
XVU8eoZwlit5RT3qnd2yHIHzzrrz3a/0SdY+QZCV1MbnJdVuc+11w46blq1yBI12OKqh6bdDBkt0
yqlxwfgkIjAp6mDKnl0sB1uNzML9QrA6GyewXqyfXJPQSLBQpCyLV9cy3zu9qq5rROtRyZAQ/AKW
RVEo87lYkGqr+0p8tSowFyG71S3SNCHxke62R09Lz3Nc4II7GeWGmh8FmntkAwV7aJsL+SLva4ar
7y9JFb0QYo/YldjzPqos/1Ds1EeEQdzccDLwKwGIGIPFPiObWpy03zReMV5JirZNB7c9lonN66D7
OAmYyM8aJxZrr/EeLOYlZY96oaTHfoq8MqCFY+tajbbGCC05uUaBOh20DvyndS/3/pIpapInOizK
qHhaHgf1r5YStpvnEl3lTKuOLFWwNUdtyxPNxnTpAUbdlC/eMcjP3hdgV6tla9BUWH/6qQ2LX1xi
7COnI10hlaFO0w33mJnPiDms2BvuYyqTOjX9F9EdT/WD4girwHwLRRxS9pGeMf7YE82o0n5V92Dg
ZaF1SmropZwrb/3FBZOC8nszQIUmG2HIH5z+8N6Yoz7JdrQl5Nv1LsjyOjiOwNgUaT2+aQkvYhsg
lBnZxEfM7hKNMiyHM3Qu5A0/OlKnshWsNIzmU4eo2NA5RLzQkMFNBqKLC3WYhPk4AT7YziS2vfIX
hI/CgSb9QP3OELNICRNk00w6XadLCHBJ0WFgcw9jbXM8bdKDCFeCl7HnTwnqqW4IDCOhTQY3WCRH
6aeFOZumt9JYNKnEdnvXmb2YESgqFSKo7960vqrmjv5t5kenNHnQKUAqiKUI4b8LCPdv1RIvURpJ
eapMN3Y8G3efni66i31MDMkZM8zrSGMmXmldHQeDl1pUGmGQXCCM9luPheZoCI7qJOIPhhL9OFoW
pm4y2JK9o/UjueStoBILySITTpx5tKKBAybdcUmgf2v699yQaV9SQt/2ewbNLkDpmxIqbW/HY4Gk
zR8HFl4p6Id0YqsINUDKCDWdHQ8xZ4/gKZ1ZFr36/avjtzt8GvIGXrl7uSb4A5SwOH1KHnat6qKf
T6PvmRxeqaBQBCT6Txlsy/8k+HW33OXPF7pPkW8F/HrLAW4YUAvNf3pRwccSgovBQ0p/kdJFGlui
4APQ7/mV1m/C9WbWKGxAbkLBiUEtdk5qwliqDblET4GfQ5zCM/hhPTdnpuK2QDk3sDueTrVEAhAI
TSxPjz5aadsAxAOIZ0S9rXX4Z2ydx5CbTcosmxF8VOvRiv0QBGdp827iNm75hGo3TbWWeNaBzav/
UmFzuszBqk2n0nYt8Ye9/Z1Nahth9+OyjpgYin9sDRH1dVFa/fne8Zttg1ol5dLcxip/1caUv3dx
JYl/Fn2CNXcpeeyOdP82HHLiSG4inTzhAsOHsKFqMY4OATHzSIQI50Uy9NZhDyA7wudfGpoSLI4G
DdFraZeSht9Xt/xpfMb4TutJl47V0dFV1F7z7Hd/iRRAdrWiCg1i3gO7QtXoQ3PwQi5Om3fT23Gx
OzfjUVMsTthOG6hZaro9wQQV9kmYFdVBE7TdYRWvLBJS7eKssZNlXZxEZkg6NcT5ka8oWZH6zNLF
29aORvQWVXBafWcCRbKmCXtU+wFWSbmKzYuHZijdx96MHQYBhs58uQ8Pj1/gDjgKwnTt2AXSFjNL
0p0esUE1iBCBuknlEhUOTYlcsG6a0j0O0uCp/J8YfS/68bBCsrPEnVxopSLmgQrEzO6lN/O0wlnK
tPNLQ6fzhrgo/wBXNrVV8pC3iQt3mCxSWfO01Jh3fO4k3DMvrUOc+1jHCa0S4+TZwaQ5+3pk3SQJ
oV96mLTMYl90oV5/W9E9MKQGAz0YkXw653DLdMsPR4Dk95TsIQ1NyyzFGXyU6H80l1PjYE578+IH
tblyWfQq2WykPdd4s7SPAN6zKhj6u1EwDN6ydN7MuMwTIa8ULTJpecqBi7sMhPPgZf5zsjt1k/Z3
7d0eAkTR8A9ZeYP8Sxm9GfyJPOXV8n4/42y0F7mcltOy7+D0WvWoPY2TTl98epWOb9WNhBSIqxvf
341GJm2YZJ6pUm3DzanFDiujVBEKpbaaXf7czXwPnwOF4uzgBEwGH30qv6DxKRiFRFNVaS/tx8Uk
PT4GLTeor7MVlUWJAntgRlN86aVbI6G7JsqLxcCnGH2vjn6hWbcZiLpPuw2VFbmIZpg3fvkRmeQc
1KTJ/bTW6oF9CzXR3c0vdx4O95Uqi5SNff+lACEVqL9j9NV/s6KCwfu5SaddymVZNqkS4wF5WmAl
UByyl4BkIY38EW9nJmqdnPg2UtEaVAu/J6gUapg2Q8MFPHiMTv2mgi8XJ+lLAMlu07jfRUz2+04g
iyS1MjBIPlzTLEIHslVEvRnU/kMgt1+8bftq82nWIjHGehSKs8MuqzW7b+yE2CPuzIzxhcC3oYQQ
/9igDMjYqtmEiSFHXOfqgiAw/gg5/Mzqu84gKN9XotE3oxtEJff0R36/6ENGEXDZgR05shCqIblG
6xhSvl8YqdO6JHIH+ACS7IruAe4JOjbS53ZHo7PffUl6RSkbtWYB/RAvCgRZx3UJwZWpSXL+eMbQ
Jwtamig24nyZgs4cuzlKx3Xktx6gqpVMfLDRv/mvuBjk35q+OWSABr2zof2wCikcPP1W5vAqE4ii
UzKM7/H1I/r8lTJ5LhyxEkiVW7bd7UVD72o50mDbr572VYnlRLyNrn2gyGHfvlxEu/kJME6f3jzq
2QYfoKYCyptPewjZbn8xCnG5dVwrgAOMIRtdF9j896lBgsBvm69byLgep5APxa1tsh2QSLPvuSVz
gvPWjNo7qIp2NoXKTPTDeJoap/ArPo2c6Des7nxMlnfqMpXa2hpop7BvUu+3/PpFpvY/5Tc65c0Q
NeLyOQW8MSLjZvo9aX7UYVRqCeRLThnaCHtkccSonID6/w1zm5OI3WSBauSdnT/RTOtAH8C6UyWY
cQ7gJwmaME85y3I/caPpFyFTx2ECfQuo5vhJfHYJxKRKOQqRf3/3oJs1AAiHfGsSzaXiV0bDGWFQ
fKGvTkrZVXrBY4PvQBjH8I1GMOYuRF+LzwI2lbRWsrIl1vZ1QDrhi/vH+mvtke16M1hXweJduIzS
QoOLbt7G4U7Aua3X/ZTfOa8Hn3aS53isiUJmutGfN6d8DFOmJDVA5xVXj9w0V3WWyO5KGT75PhcZ
2HhwgUkEkddVN1PGYZxuJY7upBxrb50XdizFAkSvSl0vnhBGFE9cPq2WTAx0Zthja0bSfv13FOXk
DDcZvoiy/WvVLSW7O1ivhXdAhw41TxhxAF7LHmcj74Ae3LrxftRhGytuAofP9Xj7KPxOCYTRqxjK
uG9EPkdG96CdJ2pmLQLqwuA/kTuABl81OOEw9k5g4TKClADJ1si+XehyjPUZ6L5UYMn3L9/kIKuj
aLrx4oEe+HhurLXwd9Bk9/F1rjAd/bBRRS2j7jTidu2PgTCBuHXXBcXvnuWJvRVypI8b2bpk8evY
HJ/QxiBDGBr4bdIp9tlaA5y+bOx23Psa2Kfb7rvrggcSfqZ0BriOoW3SItKk6EGbgzaREmTpQvQE
hv6bI2Qxwor8vZUbIMZypnYsaGUgBaeLXEi7qP+8Q3sSYckRFC9u/N6qA5mywf8aJbJzpcSYgk9l
6uMuPzJzK0PTI6bD0E7F0KmGGms6x4Qcrrknlk6s25UItARqf8RSNtnZLH28cgJHUFp6Don5h7HH
25+W6OV74uu5nVTMmIjII2CU22Nu1ZgBy188OVu+VLxO/Gs/Icuq9YMCZd5oiMFe2r+xwzQuzqLw
e81VG3nscG1CgVOhtQIXk41qGFu9j8DyQngIXHbdQnRLCWfbzTlV2Ujve9Sk1o5azdNZH/iPqtPm
Uw785ERHdMGgvQYMW48G4oAGxVF7da7LxLH3WHm69jGqm7HeCYvGUycRgdfPsaF7nS1PQhsGA2uZ
DYOzllhk8vAJrucZegM+3ylqU/wov8MBTCD8HdauOShKHDniuA5iUOphFXGgQNVYcbClQwKCyUy/
3UiOcEEULOLxah49VBoTbLl7EsgRe5zwoynreaBMpsm4l5gNUREsUPyttjKXoUB+YcNxJIbxMQAe
BmFN2Am0Z1S6LcR9Zw3M0ylXr/SmcrMJnQbRREKp5g4kn4plImu9WoKWCvxAY9lQAdOR+uR2nQ/8
fijjNVjzwifawl8rEplbav+1xl7HOiz26MqpsaYWo5nPSH6uQ+IG/ISM4OqAnJ/oDlpEzAnCzgL2
tDKYhzzlHS/FeOJKcG8iJQ0mJDXywcKTyLCjj7PfE09hFKmVTo3FmwGsKbEQV9NknLkSyglUomfE
Zng2UW//9WaGIzgrfLrV2zFNzqagycD1W8PLjZ95tI3CYejzbVH6fW5UWE/w2MbqjkLvLuSfhqW6
HIp+Hi15ikdTU3hwH7c0XnqwvhrSCC83ClZdeRxuvw89gmD/6ixk557mFpEngpD6PrRpCPnnY8qy
b4tMkMgYEZMjtBIyckCLBjOBs0Ui16rU5jP2QtDgTgGTNYfRhSS2w5BhmGzRKnm52vSKLm2g/cpL
KbMm/A8lFEOHIHSxDhL8/ltBrJxv7oS0R6+qYtkxwUA8d5JwzSSiNRgWYdgBlkPNTf9Wj2Yv/9QW
ZXNJoe2Zf1FseYZBJ243YS/6aCILqNuNjE0ss+iyDC17jj6pfkJMxe4uOh4rIU8K+jOA9+zgsVVD
qtU/UW/whOb8EVNLP028avh/Jew3Gm7PqguablHLBkPaEGSVlXqepiO+pfiirkrXV66AQWELGxeE
9R/JU7WmSHrKV5+KNAbWmCB6cvIj2ycv42EcQf6ivwMRWRVdXvB6Iufb/r7xM6VhBX6mLZXmLMqW
pI9JjqoHbJefVssiz0SCCK9j/Wl/LQvS7XuPZtCh9bLNKA4to34k1JrxQxyymNov4Qv3mjWvm9F4
5xOYD90lF3MA/rm3zYB55Zixuf2fkTpqkenvjRd/aS+D9WSzLSmVmOzqhvLGTTbwXxocBPQ+3qIY
QGb90d/V51/aNXQnz/l/Js6qa3nwVbL0d7hFKQ/naLIn9FNeNVSAXHW6OlITJfXAcZYd0BGoPDCE
7WXpYqPWsuJY1UZtAUvb7CGu12eOgMU/smIbAcB5XN8gngubRkl08b+W1Fw8QimPQCh5sEtcZYHh
U258+/WQKN8gmB376MG52k5QPe4GNrPMTeyD7sMTE1kMkxtmgc0metETshpsfLhjDOB9xrRAvstE
tdFsaDcpTENcQ/nGLULn+aUISHGw489z3GkU38r40UkyJjNdjjDfN5M+tQrkUPGykzXq9iNY1+pP
/CkFOrq68RKSrn3WEyJdrfbVZS4fh6nwNWz+Sqmhl0k9leHFYb9p+3zF7YLQ7rRunXbooonToOpd
HqUNrhdVgDooh/BNtA76SowacL9or5UfNRviTHZ2kc42/ZuoiKTgHVqIwjY1FQo6GfF8MIiyETSY
0e7xB521UhN5FZPr2nlX6qFXFJU0Gu7FDGmQCdxlSHWCSLyWx2Y3jWtPu/sX0h53Aixgr0QgKRTD
JkyLsYaskcC/jWhgfJ1oeW0uaKRp3jTN+Gv22HNLg+hLCpR67SDVpSR+RwiqSI7S+qPjw7HfNTax
EN2j0kyk3c8k7dla0N08TgjP4v+u5zc6pkLlFmNROuidD4C8yxORPe/5ovp+rqk7O3VwsOZraIVd
3mld9BLbuZyFBv0l0g+K6tytB+PKP5Qc0Tsmg5ZFqWRy4ZSdmZjMwomO754KyFAHLZ7yIkygQapG
CWV5LPlRHUQvGbXnZTnGKRiCrCjNvQOyYndCRp+GZcaouTLaQtABVF3UjLSOGwxWnccWCd/1+tTB
OZwhFduaGAksBU1omt6xqVBSONisL+PU4e95S71ziZOERIvlAxWNxyTuOKveew1mMuYkK91gHpZ5
J+o/ZVLQa9YDaeGd49e7uU1FDwkAB8AYGrfk6LwIkvhgQzi317RjTpqpB8ZKuUyUiCo2GDpvRbML
erRzq7JeFOGaZ4hKcvQSlOYJybcYWvkOkGY0/WY/2htKzl6v1RbhmcWufQT5/EC8SCbPbVZoMLel
z7KV2r/Fwt/KkAS0cYsDZuAAzZZkYjev8+y6xA0VZjlxNUFjFE/8YItHINL/tR8JJJyFFTW0EH3R
cSSNevrPROg/BlycXZmY6qpdaHkZviOOWMo3RA/6DdxoIMiv6WOxxnt6iPmDO8HXIi/b97gOiA93
7YpdYQ5s7X/zjiTSMhrVArTwbH/qcgQOWBfl4r6bn7uCXMlk2iZLrp+9pjzypNIZsc+r20oTQQsN
uPshB0/1BGI1XMIP//EtZAefcvXH0vgC46UrDMRXVAwApSR7cJTy+BWwWjFNkb4/hw5Pq20kBsYN
rQaY+LWL/B62iCRk5zIRMCMHcwbjTHRy5fFprAlzMXHNlt8K/RAjsQ59zbvOtoSteKgD8JPzrs3Z
lzpG2LNzIe/jhhUVesjfH+BO4A330G/ITeNbBvTwuBcgO59Z3h+dqBdb2xmq9dt3fXg9bnZXU0Rg
4g/aWpVls48FGHRFLA7xGmpxDDuEBuhKiUQW4MdBqE/sHQsaulUeC+q+5KNphl6Kl0RoEnHLYAj1
VpLTviwWF1SU6ThQw+/IRK+GYuVcpbWJ1syVgRp0XoJjYs8PCa/YBZwPoAA+U+phfyGHgK1y5CT6
aoicDHLb8hPbqvavVTXmkB4C+Ur9NHM2H5nnWxD1yrm1SKr7Fl2Bj1vdeKHVurpkX58sj+yWV/9F
rzyraHq3rie9cjZbxNntJtMXlf974HjznuOhndxF2xxtuyU9eo6+e9uy9RSAk6YYUnTg9Ys6rG+V
tRudYONiVOdtcETlSZ6wflSyv3ZsgvnQUH5DTWBw7HexwPT8wRQprVP14ZeSnyA+N5AYS3Z6me29
eDS1U0xix9DgRZR0HRftODWXzFAT/PiH3JrtH8G2Pm4MAc4AgUFn4WgZoCyRfq1ZaHSu9porT6uX
is06N+KRgEY1Z8C8VaPYPlgt8q8erV4Yzjv9OWPkc/xii02AK7J9DikSE+NHumeAB7miVDBL+PsD
GuB5Wm/P9FSnJ8nfg1YZbtzOR8eRHdZJlvb0FReTC6fNeXHJVFlztBZgvpZRhgrR2L3P6TlicX5o
NcIXRw1pucYHdVB3WDreZWo02N/qGXyDz/keQb/Sh0buXS0orKvSyf1hWAeJbHH0x7UsgKevr78j
O9dxaf5XQparF8YjkZUZN+aWWAYEk3UlGec4SZGtuH7aoLg35bs4w/p1M51T5iexzfJZpesV45cW
1/9tNU6A2Ggx1HWttN9ySCsGJK9/96WJTWBcCLZoVj4JBwDKSM0KZyxsbWBMgZVfDfBFgV0wMPOu
BaZynT2fvvrYgBWNLeiLb6zx3Gr3bV3dL/l+z3AMyn4Sd4FFp69EZZkQP7PaypJXJyw1IuW9OgvV
R5anXFT0ImYCEMTPscGFRzfA0ly+NG/38r49I3QAaM2CklUIyLkh2EEyAglhY1MB1BLzHhuOPTcf
vYqsQRyivYaQ5qmUQ/Djm6xreIHUzUvy9Zj9FO7+OxIvS0rJp0bKulvG4QDhmirhkWyMbWFp8n/1
iR+5Hk/ZxlU3k/v8BcaL7t/MxEUqzAILjxAxLZppiCFq6LZZNA4+iAMTq6DdWQSpv0QP3RbuWRuE
kTAFN620vNRDrMmuNonH+5kdzhe0NGInN994q0iQ1QQwpUA5SHQVC7Qyxw7Z+MDlJqL0E4ReLHME
l1qsNO9pvcCODttiwsvaIfb17C5ie7w12u1dEqNL7Iv90TQGffIzlmC/mkbZWXUTbhuYJDP9komK
uQYn68usfxKZ1Rjq8ePLotGOAgEXw/alnRUT/DK7jHmBZMtDjqJYVe4c5mwjmk/EQkcsg4pcfCEV
y3cE/3sosYjoupTfW6GUFa4XhbG+puBYj/mwZKU4H+JxpSnM3JY6KrHZ5hBtbMBfYRIMY0p7IhrO
jWxGl2NU5frnXPkt1D53GaDYJ2URSr7nwCZKgmqqKRO2wVAp7pvmDUSNSVkbdX9aT4Ya4N8ZDqUe
owd1BAm2fs+OSI+C4Ai+yWBWtkKdGQ3SUHZv96J28jgO4UdM1pa84yDpXODE0hQMSnaEetjIUZu/
+XPLI6Sq5zKm52HkKHXtdeS8ed40TAEt9uzZB9X8Zv+Kdv/9GY0FdLNA0W05+wgnO72BmGAqox9X
oyTMzjjuWkvD+CwofNO1nhlbMDF0hSXpTdh9DfEHk+x/eqlNR8y8AFUtjV5Rqzyk0rK2A/T6a0zA
MoW8cjsBbPe7tpzHxRsSR1K6Y1I+vrJUgM4v1UB1we0YK9AvdnPHzfX+SHnIi9lgvWtMbsuq+SEC
1Ezlw98xatBl5B7sk2G97OhxodPkiz4BNzAOEMDyseQYt6wih4eyc8f9THgrJsI28sT9gBsus3K6
HvX2AuskY4SSpUgs3M28eUYFtnOhyX83hBAFaZTISJsJoeDw85A3OyRTh3f7sIHqwnv9nyGgOZdP
QvSWW7YTc7uP4ziDzmSpYNAhkm5JM9n8nGYeyDULebj/CgbKIpUEc6YKAyi2FlUAId7OD1lU6cb1
cIM3hnMsfQRFI6SWX+Gwv+OjfghgioBmX9X/A9WcAArqRqqlZv5VdIk5aDnElQGTvZwGgRX1hX44
XLkbHQF5EiUjCxLiTZ3M9STuvaIEwfv+qaSW9F6V7TNePFWb7YIHdNfFEEMvDGX2GItMis1XJsSv
RMEpNIIyTTYfWsH8hP6PjTr2JMtQ2o0wkJzpGql1SkEfPZ75xYV4M+1Xki4QQbRGYPo1UC8FHJQ7
tOJ2R7MowiHfua10fIi2SU2y7cwYPcV/aCdufJPUgrELZ+MoWIehLH/hbAKM477WK95ZrsxaXvK6
FnomlEWcanE65KpJ38mMlyiy12xbYvcT2NmzLEzqeHPowbjicjuVs9JGJ5y4NKyW2qmWCWy7RIpi
vKRe5HUseHMYtd/3zZpX28qYUFlX1sKa22tCejHvN6L60UtYJ5hhbVn0Gs/piOJkgVZ1dkrAQz2x
2vQmzdSMY42AnqoIOG9Zui+3Bvsxk4wF7tm5/6i4Y3pFDh+wObil27iJ9o+ua5wvw1HOuU+1NMWp
lOWUw+tE7oW/mioNoj6fYw0GFhDfNhfv8pfZgZDXE4TGj3tSI7P/1oz8hyMJ/EeAo1PBAEXgn4nG
M4XH/H2ZaCibgAGbcpLBey6O5tm7Wy5alhBtVhldpn6+xP5MVYZheiJAEZsehZQpHwS/L1grvjAy
dn1SSehpwa1MQ1UpCsl4ndQG8EkEiDb8iPcTlL7I1JA6uyrRFxcef7MrgTE9hjtyfNzgpOuixcb0
L+ZjV8tym+Rqv7q8jUMzn6vsCvuJmqdctKmm6BUi0j1HdzmFqKgP9h3bmSh5G7PZeoIuZ7uVBTp/
+M4LlWk37B6NbrRIjhUJz4M7PxaFklP++gFByAHfhAH8v6FZWz9bTyZRwcnCP5nwKt7q4vM5vJdi
Maym1jI+/POQUuurgjSwEucPI5AH8LtTcdHosbyZqjUtTgNEf5VHY+zYOFRmvjG+Z4G4VZ9HWbzd
Q1KUQm1P/DtKCZStuhxrarMhUKPCjQMI/Kz6rsSnUdLQ+zIPZk2xgyRwrDGUV3GY881DK/5yLSqu
FgtT4MCVRRfgTnFKTX8f/72WvZ4p0rSSLY2S9mSIr1yaIanYbk+GFWP6iZyfkrTYJY7EC9IvkQC4
G0BoCuCeUvQrynqbYYs3TrscQ4Gy1RD5ElCOItIC/VYXm35WC93x85iUHATHKg2y4aRfV6UfaM3T
thb/GhQty8s74Xa/TBVAtjJpqMUCuvDId6mbVL4zAeCt0xhRvQ5tzhf8jsXonV2YBCtlL/96cfwF
2BACaLsVxouTrAeajS5Qmmhvpx6YxVgVxSkGAau83zL8gQqQlasQG0wRzkhGapiYl9h7n0lqivLZ
p+of1gQyTH55gSuGqzHM2/XNq9WEN0fZPZWVqWALaZK9k5dWMuCdD3ZpTYtdtu/svmpsbCcT8aYm
OjV+udvq9C5x0Imj+0UkBzdAxaohdcxgt3N1Vs4SDUYMgqP46R80bMApRZnjBUseirkalxDbWejV
4j9dG3W2ovI7+pBhaUbQR7bpFut476Q/6tkrRGAINeW2g6mV1cRDRZ2ZzdxD6y300usEGxLjkScn
VJ50Lqs6U7Rp/SW8sg/9OlqJGlUBp5zcoxZitOK36ImXMxMH5CFTekNiH8niAfn7QaBht5/uM8CK
7ZOKgOYjMvR+sWBtsWJMXUFHh4SdUzYhOAnEa+U5EJ2r9CnbP0kykVeNGiaMY0nHowQgLcgNLXaY
hUvwDZosneU9Tr+DOGYEg/YJRLe+tlA6x2XWtLMoXPc3X+z3Ull3cJvb5pCXWaU4Wvs7zs2Ci+Ch
tVso+ym3xBt+d5uZNNpJu5cGSBqZg1TWwvKRu/7M+4FZs8ACe1Nen+4ykwfdBKdcCyydD3kcvNs8
ykQoSNoklw2eAqaJqBreSLtn23bqhN7gS7fccpJaY5EAaTL3k3j8J/ddPvyqDn4mp2yU1Q/ke7xK
eFyOi8Ijm36H+EiivzpFxDnPUgxMy/Xc1Ubf3+o5j+W01170UBSaX17WTlbjr/1QLeF3i56FRYP1
onJSLD8zy0dKwlFSvJWXbcXH3wSNy9ru8Dq1FiptBPMYtlB+jrAb02KYLOUUUorLU5W/4AgPTh8L
NJnSTNI1q5QYEqqAEItfsPHCcJXiERZRdDCDeEaoyT53kVYriLsndd9RnsKj92ue582nj5pGDq/e
1vls/xBldKVscvgSorQ0lQjdcFqtLF3g88DUuo6X9R0Lr+wZiXg9DH67cd2bkRyjJWES9EOJMDcO
Nl2+diuhbp2Pjzcs2snnZsF+jqzqq4vm74ev2LOlhLLXtT6KSxh2g0hTcytDq0VchXKbDnWQcMNd
EWLiwzIcR+gl6tRNfq7ezQhl6H8cg+Y3fG1IHUe0tNmkcVIRaytUAwb1B3YHI5RCAV+47PKJSUBU
A7eWSV7UTYIbL/nKHXy6EqWht93CdXJ6ahfgoaSw3vYcvQQ6Dx5vStRv/g/Q5AkiWOnElLKDMIn2
BbaecxJR+0XMX63SISQCCkCxFA4ww5s1FLRVfVLXahqZBGjbyPUCrYPtW6vHZGwff9Z8ozi4xMeo
W5iikKVZ6y9mq/nhSrI+zvVqYeXpUF+cYwKpFTpnBqUCJcFyOEwPFw1lm+UHvYcLhetLE0z47jTj
cVGmWrMefvCB1R7jZVS3IhlpeLuLHAD8lDnXIO7uxr5qBLNSY99C3QjwN5ZDKQQF21nYVNLE70Po
6cQ5sJCcEu/dP0uDes/ota2WCq6NAR6mEydjuwR5WQ75Sf6J9XP25XXGMPqVnS5slioqNhwkCQHV
RL4lZVRnkL8S1pu4i/xKHZQ24/dkgt8GQVl1HAZDsURdS3faRMhjLZjIKEs7G6mlevMIhIyVwlk4
LwOS3Z8T/pRCviZQ7+qDbR8J7qw8Zp+PAf9+eJgP+rhXZOR60MX3uWUC7cTWXexUMPKf3572cae5
RhwukRGjetQ9cQPU6fij2jLrJy95CJhat3+URwW9U/ZCJ4grpbadhnbomDlwtFJ0KU9gj+raKpiI
f77gnEdQnMuvNe0xF8aL3ZpHaynS7+pvpAn0zF2tqVfISlu8u6RTezfjr4CnHiKyJMwxo7iK9Naq
Dudkbcj2PMFtwTeZRlQ25ai/55k5uzKs7avLc6911g2Vlb5x5zMZNv0+p0cJ6mhMuwDO6eflbGHb
/2DwatTVWNCJQzywDJpdPyzFXo0T9UFMMQw+8oNvwx9OyrDtw0kLb/0RNpmyzaVkGIyr5SA2xyRP
Db4wk3jXsQ+rM3yh4Walw3LNxvPk/sLEu2FmocUqRm75ihBsAZzL1dQeQ0khXqYwGiEduj2J0zoG
fNlNWQYqFyrrqkXVlTMDDkMpKW3oIj6B/afGB+cn7hwvKtwW2OwxKakj4UWW7i5DRmsrc6ulxy4m
21RpZYPjjt7g6kH6mhze3cadlPLdE6TsK8Ckw7lUR0Z1j9rbdapcC8UPbiyA4wvCG0zDGFPZkLVa
E5EmuPLCjiN9Yo29oIL8+3oYnZEXxFiIZTzm/UNLoVZFvMTWuHXjUfERUf/B42nplPQxL4Kuuvnn
hHXYiEPhYxY1ftJs/pY7eaIOyqkXo5NPwbv2V6AkP6fXOE1e6IiiYJWnG0aHlrccBgj597JuiIwg
2aEe+Ay2V1NZt+qJ3f9/8cWgRe1u00aW05bQ5rgh1HHuBNvXOkcwvdPtRLMGdV+aG3VdxLG06wME
NFmpkLSGx4J1iCY3dL/uCz/s1QXefR9ZjY0YbVMt30txvFr869he8X/nxUXrcYhWlL7fZ5uDR1Oc
bQPdUOco4/Kw0J/DQvRGz0PqmCcxRZ0anFSwptIwDRB73xsh4sUH5CawgoQYksaXoJ3CRpsNc29S
a7QaIdQ39qQaxPxkEwZE8A0VBVCoUx+T2NM6hNecxctsOY7wxd2reGSBUQ5Eg1hYmAsarKoLIRIy
cWA75g6nEuSftvhYI9A7oa96sA4y2d2marwtueZ7q5b6cWa3z1Lkj1hVWZXLNetmG8By5N6T+WoS
cQFH0TyZuCfOFCk+ovrWqxyknfBOqaDJBFo1SZLBZDaDheCPLFSsIDL2XLCD1ZT0PTzWhBz2uoGB
z9Vg/9FLAcOvggv3CPtXirB0bXFUhxwtEJ/v4+jYarLcnJ3MSRXvdELPrDKUu/kqNYaYT2ItJJaH
VI0g50qpaqnPEWTPiHjF8BE2bFzz5fA+TklPeF2ihTVaJDk5c2h4d75JRK9PKbo4JPXbuWIzoPxv
3fN22PaU6S6KXiMspQUYmQI+yB76B3ovNi1n8xeo9WtBIaZaNIug/Tl6qsonB9Ttu3O1omL614Hc
1feVUlzXinULJ9fqvP10P5LobfCF1g8bWiqz/H6Pcut+URfX2SMB1xgfy6FBV5aXnC9US9NofYOQ
DhhnLAjIVkq2NieNvVQKKiha2D3yUDOd8CbpoJUAzobI84kKzKQhcX/y52736W7CkZ2tCxsW8mR2
EoYFsu2hJVpfwKUupoeCTOE+hTPxtvhjDJZqJyWDqe2i66tDqEG6YZ/0YG5XOfkKeT5yfFInPWGW
mjtYDC2F1bC2qYG/v/gFBGYvXnZ6LA6XReqQ3g/YRog/rs2pqJk7K32VuBPmcYGsHLgRaIs0auYR
cFn8l8lZKNpeGCOoStx0j/KNXE/Ajuf4AkwZ+KB2BGh1E96zlH2OCbecQ9lCOXNHfzkzSjgqfxDT
o7BWk7EvHkBa0nlmlgPiYwZH6gbkmic6u/8bl2WYGnIMm25S7aakOvk0vgcjqws8RYr943MEtVgI
ZW3dGwazYWaEQcKnlm37RPOiCrcavFCV7g+sDn9caiBN6bfFAtF+8GrkQxyaX1oSJ+r2iqoyK9Yl
nYQ+j9eZIh5kFGQn8iWADtk4fwQRJc5uSFRQCta7pxTzMIAMXiTeTQ+8tXUYnwcJDP+J8RRim3Ho
DnE1l349lkJ9Zv8scKhECItowJB9iCGVGBmOA7ZQo/TDXgD6ZfnJRS7Svj1cCm6+swxZYpinrq15
THvan8tIt10A7qNgfvTFUtiXpDvtSkZ2NG546hyMy1N2Ej9/A5iv66777t1+m5utm+q+ANXZ9rnK
B8GrApZko08TVDpXMwa5IwCfi6YqQNE9ORulWdAgnpQvmjHdk6A/yXIx/B8GX5gYuvmmLvCf/bXH
TVOaGcB84YZncKLCWwS/5R0GqcnfrbHMtBompn70to96l/xTxOOhWasOz/A10uYzkld5ujyeToh+
RaXkBoud8b7IjyxSEwwSjVxVEDVKqUEOo6VcWg9H1iccfjGc9fedn5PC1AFf4bpL94Z+IpqijSDw
55IX3pTvbrVsns5Xcts0GF2v/5hVmU97o3o8eHhIkgQUJJWKctwa9Wf8gRgBwNx5JbQM+4As+jVM
q+ATclJa6f7S8GmEQi3WgdJUCh4Ne0lut97yqNf8IYDQ03rR+qT21a4zDCrCyQBKSd8CpFDVfSkD
Yw3F2mpevYn0uMQxFlExHYCj6xpzKBDC8MMOopzaUTBrPAB4YtvPHPlXDaaqoMOcZxGJh4exmIwJ
kfuU4voWaEl6I0RoUh2MkI8xjfbOSW742a0X9JQltnTZgyY5LVYSPhn8DKh1BeMcYK2ju2M7qfpx
Ay0zL+l1V8WiXdSLwjCNl5St1YILcbYHEuQMHDSgp+sbaZb3+hRir862J4sWTAS0ODBLRfd06O+O
wfHK7BekOLApT3Rn8kxjJxWuTeTz0E4YLbu6IIlcVnC55r52qyyO1zwYdlpIgz/d3zJiqLwd/5/0
008ndZaI5BJlDT5XyvKr1uNg1njQ58flklCxyCATkF6AHcfgHoyZ/cAgyIJWA7VFBDIWMCT7K0Bh
WHlYcsJA7HZxvZEhFWrqNXIFyNwmarJU+bV4+MD7JHUN1VdVBOxrTlaJgOrsUgjd2AURQUp44wZc
lWCn0KSQNESBbzA/Vqo5E5tXjGJ6CQei0cTWc8pCJ7II8d/YGJD+XTVFqL00hPwhB7Wt67BH5heZ
i4OaweyTPzfiLGdp9zPbA3FuUDIe7nxCCo3TD0HrhpRvEIvAi3yBrjcFvZ+GJsou+FH32AZE7+hd
KT+nqf9GaxCFI5Vc0iu/7lOsTtgKWTTsiRv2+xY20gUADoNTkBwL4e33wKSqmiIYi5lMn66oHJrB
vsjI2PEmPyuqn4N2vRxHcNOx74Epm7n2sxbpCxXFR6+dnGbvJMimUZsNIESLoLzCYvPs6WQHMPSR
Zz5yDD70IG309O621A+18vSMZcV5L3Zmj7aiJy0BCDsfq2EY4IiNIbb1yya7c7I6b9hJQIra3h0F
6ngtIuDSPEwYaDbEjTDelMUF5oMYRPj9dgDkAoihBUSo/XBbNYXE1X1ND6Jy+2ceiWf2gk/XPCwh
MHkZOSP3/PA2LY1nwKFZwf/WErZk7n7+RkaA30I/TgPXk1XWlMjS3LHciCCCQYODSh6whVkHxOES
mRHZpZCoUVVgmlWwaZJ6IhMKh3jth46wejFX+BhJo4kij5zXhleW82YE9Ge2UUXa3F85xiChO74w
s3Tyf5Byllp+qqFMelHGcViwGhOGvr+6vxtnXdE1j5q6BXH+10S0PY7ZgbvOK3Rd9NFqEsDHyMg4
AN4yVFkmZwKPucEYxLT0c0WY1I8kBqbvXcjmIuqvgQucpg6qgXmeGq94kqDmERmMIdQNpBJb37Ma
TEem9u9yFbdtiWPlXFhzWf3Tjvfp+4hQUNODPjd4ab0lL3VdxOG9YQP3vyVVSoZi6QuXCRYXHpcp
c4yZAf9cJbYiImZp2xI03YoXXXpuj41K+FtM4A3GsOzOnnXkHeG9gT79uc2uHr0klS+bgSElN2I3
cwOa+yFAH7QmdqBAikLrld6sP2KNQqJn+a0oF9/MJMIKptrTr/ru6fCZjnLFxaUTTnWNa2c0lu4V
dfhgHg0IWldXtFrJny2xK066vXjx/0V7aMKtb93Xp/am8yHBupQ/jXOwQTMVZz5wfro+VyneF2bE
pqhiWsF3VxOBwMqwV4SFdaSAiR3BmKG+Is24wlq+WKRzrrFlMaybtgzRLl8uUXZRUjHd2oQ62/lm
wp9j123TvvgSNhdWl50s9VbEBZgtKYZYLdbW3OnUzPJ4gbR8/Y8cRg94nCimNwQ9sFWU7LXHjvPq
DSvX+cKxsh4o7+0woN7wXvdaGsGrIMT5qx7fDHBdiHV3M/KP1TXq54q35ezD/25sgL3lR3C1gtXK
tug0tdOB+LbtzsbY0le7BqP9mT1x3JUGyQqyzBoSiEh/hZOEwMzozms4R0YeHrm1BjhETc+eESjT
tA+8xJewGb7i7Gi5KKApb6A0gn8iTCoNPiE1bFJ1NiN6je8p+n6Q6ast5Eo1hlG0g596Wn5EgKWM
gWj3Jboi6u904t9rLn/ilnIbdWw9HQoIQ4pFZ8TPiRt7MB+m2PJy6oJeDwVNBp2mrQsmvSpiveyu
1nG5BG3rgQiYynvfu/7gNsvckffc8d3s+KfuHqYJXtCQjcy1xiOzs80yrrYcEIkKYvx6uIPGKD6w
xTkfVmfJ4Sa+VL+N9ShEjCQenDW7H8n++8lPYjFx1+LgwGQqEDl2PzzHIddraFbp2MzdQ58yL6Po
yHTC7LSZRcg+lrND31OvtGfPablCLVCWa38H90vx+cx/kfAiK5HUlcz8TfKFh7RoIecsxRfJe0Ua
q2YtIKAhW8FCU9JG84PMYkNyTArZcTWO13u29CajhlY0DgRGn28BbsltPKHzcQmfLg/ZX/lijRq7
QARqn/d429XC4yRkCtiiaQ48OQAr7jdyGCaIiludh6wfVFL5fTS0RUMNMDv26LWd7Q0ykU605+3T
m8YjCh1jNfvGIzro5yEkh05ewFpZ056g0L7UsG0uc2EVd1Dm0iQIb315zn/g5r4K/xBETBTTqeN0
vMCQVTYe045HaggN1MsBCmCcZEs31ypjHsibbdg93EMdmTIBFks6CtgIXv1TvGmTk7WxlmsAdIWA
O35piqGO9B4ehm8Ps6QXW77r2Leuyuk2EUouUHSz38HHNzqm4n609xBlUGrGjVWOXaT47T+72ilJ
m/EqnC7EoOMVACiXOmApB0D67aNzjXw04/yMZOKQz5YgnYMzlaqXFoVA9jmfIBHgz9jEg0WekLdB
FeJd+7X8nvIMjQr1lgWDDWvRwEQfA9njC2edgUzBt6ZB8KEK5zbqHrSySJJQMbl64VLzVmMuDTCZ
sJ2bz1UO8DHpSHt3X/e6p8429r29vCx7vSin/0h8HQ0YUOtvFT9/6qFOgPNQyOq/9FVtp6+cf29s
NkpupsZc6sEWKvjfR8REgxgIAbT4WK6/xCf5njETSdId/0JTYmnEWBMD2WsFrLX8F4qxOx9gSafM
xXbB/ogDXSjeJBimYLcZj3e8dR4POIcgMJ3n0HygIy/zU+2LlETrmjQTNhoCZKL3QPiLsQ1h3jhx
HTx32DgM6G5Ghi8/Ku4W+G2/PAga41mc5XBrHOGYxRmWZLiRuBkqn22qVBoxLGHJyv1wRP1mOjGN
JLX8FylmUDfvm/M2gRj19ZjcUTwdPXH8r3DZyVFZMJ7+Dd8kayjKcFgw5T1tZbAsKuc22+Ux/Uas
yjtSJRz0Tw6hZshLOXTQvMGpnwvb3vabMr0JjdBLyAVfb908NXW4HGhuEGJoubcRoo84iqbHDeH3
OHkXLmpHQO6EBpMb1nKooNNh6QJ5MMe8oKAgFb1INCFEosI8AmLB+h95mwX7+1Autr5wJVkUZL5V
HcX0lRkfLpAsoZNINy4al2Gh+n/c9nkHtZBGLYWHfs7NbXm/So2FZcyY9WB3Ch5O0ZvaOypbKn4/
mJ8KXmuU4rmg0wgdB52Jg+C0uIrNIipClgx7yNmXZItQsJDs3foAiSkiAam1hMNGhgVcbLhaErrC
jHukd/vZpPlML83RghEa0zXfHcri4H3+GVTw6OFwr89MbKNkiFcmxUll2tDgsaG7uJZO98hZa9lB
lAuNJfSWshyhnuAhrwDiNJEaQwkQybLSuLrFxZFA7MufTmBm7px4rSFamPWIpytxpJzpTMT8eXqK
W+8H+fMQJ23VeR02QrWX57Jpq1EAYSJLqpL2YhlOWvFboqYm6ozb5Ko7bq/pVYYaSW8uia2zMT4C
RP4odJriYoxhLyn2P6DAHutBFZgYrm8g1Hs4k+y05QeHQyAJI7mwf4C25SwmMD0fBxYO9bRqTToZ
01Sh9DMHQbD0wMOgpinKdlwaknG47UggGMkv8W7VtLEcmw9lKpv9oSFYoO6ErdVaYFTQa7bSrJBQ
nIR5RKqNh1yrexRLGPrvyfAA1ZDfvZ6n5XVLVr8xVwz/8SKbhWWhBbjyWBjGfLvsbN5TS+DEsCO1
AY9fstG8J9qJu3zzzYXzNRFGSH5UfsG4tyJIW43LNwTi62yH9hyHMxMYylWmcK/jDfqq8+rmrnBk
qOli+XTgITYHxJw0lMman71GY9jJ0+K/BtQCZvSQdoH5hCbT+WuHPRmRwybfzndXqpARkdPl4ath
cMX+ANSpUC4LHiIfZFs22q1CBcR9+eBBxZZqdTQYjm4kBb5N27YaKOHzizcY7BY1+fuE9UcdLrzW
+VqPEQAaAikSdac3KRFku32HHF0K+pYNBqb1Gyab6dwetHw8qYphvWp65S4BUerjC32QapS8RCbq
m2m/ekDCcGUMmzPbscfm94VkAuUgHO5sMGvLKWtFL51lh3OvCk9LNYHCW/mfKqO6vNRPPDgrlgu1
42or4rgxCTOLryQIlLAiAAHgqarZzzPRyJKi2efEa5apY6V852xltON1ZwjbEjDzvJnjCw/PoAn7
VAnPVl5nxGgesvMqu+LNylE8momUs0INRWd2nUTinmtwUcnWVsETRnIrfYbpgwdW49ldHWbQD4ji
qU8VpVr+JKXvvtgJrL7n2ellYoSuQxJAnhEwzC0G1f31xbeBJEajP3vR+hAiJCtHabjKQv63hlzP
srwcSu9IrM4/iozXyS3ryDmls7my2JAHYlaNhayBlvxMKlWTu8+EEdExOW08EeTR+w+EuC9NB1HH
6dFxcGOHWGO89RwyE4e1QDLOD3e9zvTS6MuIxROOwb8EpdbAkDj0gxVWkgyBQR9NAw7XHf1MSXHy
Is90OH6iTzeVDm2uwdrWJLAEJIhGoZl/VlwjD3Nciesh3Vhy51kXObifgNAu3taE2Wtlwqxu4Tbp
20eyfr8WB3d5wC/JWGPQFDGYLjguoko0D2iya4aUUkBIu1wNtCmXiBg/Z4d5301raSGjvP0AnUnQ
vVxo+u74cDpI/C9p8N4QYkvZL+NqBdpYZ8DFqgbXMWOV6zxEpJ6yQS/AQDUl/1bsu4YR0Wkt0qpJ
woUebYW442eWvW9msKMLgmM/NpAvohMdCPDORjPuOSvHsnANrnHx90/faSukeSx8lgV8CpkEmYhO
i0GndG9mCvD9N81VMZkOBNiNuzz3AnV8A7EdApHfGqhOLRS0SWCC6oujXQCHsCaXPctxaB7hkd59
85Z6e8fO1/R5P0R1TEhVeqYbxYMNRszy/YW+IAcoNXKh+Jc+kNZZ+rhrKKTuycczLyjCXtx9Zmtz
KWyPSkaIOzSVMcU8SWXv4xSjYARlJoWinVMzU7xHDxy7zZpeo4XRrSsXwSz2Xti2HIUXticD07Kx
/pAKUar/IiccqfEdJN9o6l+kAgJebzqsK9ATZHRxMZBhNPxW9ilf2z1B0Fngd6fEh89n+3VK9aho
1yqzRXEvNYymTWux3rkc90Ud5utq95oNovzx6LxPVBW+3CRxfHfhycRBCZyRkPju1GEcnovf3ks0
KX34kiWLo3rISV0kXuqk7qD2bZLjpLMuUXzE30KFqyXR1buI38oCH1NRwgb8Ixz+DiicKb+dYUaI
oMkOi41gtSfIxmxxlp+2XoRdLmAEWjtIsXYeALohcPYqXd3oJdU2w/dZDt22EBXrbstuSwLIybXP
Kd/LHOXDyL1Z6LuswLCf8d1aF2Vqlj3sUGDuweqLiKu+A+REj1f7xew1ApkrTeosVrOv0kcc+l0H
tvdamWed8pJStbnnSIZ1UtNOhj0XkJXTG+Uq8dKUJJ/CfPOeC5UmGc0IbFnhNAc+tdq7z/IYVGpR
LAJf4KpR4Cdz/Bywp2VEqDYycyjaOfoZ8yjj0mUrewZ+fg6v2bN47dpNxPUX5YQSJh+Au2COBth3
0fnftpoJZlf8l8Z0JsrG6eF0j9PgexN17Upt44PN5J5llxNtR9MrnYH7dyS3UDcm9XJSnxpXsVPK
Qwc2ocR360wKrkyHxRwPB9Ua5ySv4fx2tWAsqRiSg9mhDcVv4Tlr5ptDTg4yS5AvN7KX+8foo4Jm
qEHBOE+Ykj03S6HFNfNSGcaL/tuxeWQ/F1FdY+GzUny4ibFimDxU78cCf1xPu9cfZjvCUcnPLbsi
471tIwUj1jwwt1dRYXJ0LZx6m9gAtXIxI9j1Vy0IgYjZk/2dWwZYmiUtUslj7QE/yvDrhIfJXZun
LUvp4aQkx5FJ1yZa+UmJZqIKrfWZPDeBhvLyojh5FeEzKH4aFkjmiwKEyvRbvKP0W5J92uPkPB2m
5YTcXjXQMKC78O77xgH14BNwaN2lLADOXCSpqzeA/AgsqbG+2AL5g0F7kZUuzRYpoLu1YMwjA1hc
7mH1VOfk+IJZKSTLaxRWr9mU88hTSlfJLWrcTpM415gvWRsAAgKNpanr5QVxzVm8dKbIPRHb70l0
JbgZfe/+Fn3+I2fhHCdFWeDtNvDeFTlxE8Vz2cHNe3pQ6cJqk3nTezxPDCrbu9Wn8WNwcqEuSpjF
O0ibZD2A6USmyBm+XOYXKCFiLVnefpODkKmJf/rdYpStBRe06xBh1rtQg/Ix8QQcBMxiXEXLLuqU
P2NVTsQQTLQA1bdAzNg7An9W+QeH34I3qgWkRDwNPeYqtA86OhfhDvhSK7U1+d8Df6KWsiHzQ727
83p3FtF1hSbGHpqc3EUsIY4AvDOIeayy5zAcoDD0w2uD3ip7aru/2E6wdz+X5o31kZXBj14tvp1W
Yy1ge/vYhiaVlmy4KM3A5FN0+40qqRhlQtEog1VCQbNZLIYBidc5TZKtyOticubN0kfgwkbFZChY
0RVgPnWmNa7TlQLaoRYcMmd9+xwXDamH5DDgYW2w5wHpoQeQB34CaRi6WB6f8yrqzEWhoBeabJqv
deANqPuC4rVcwfE3bITu5TI+toBVEwhFKY40Z+e+Poyy6pCKdv8no96M6QMX5Qnax1fQPOBb4rl0
i8nOeDmvA7VMOGEyph7c7sYvWOUK5VcnFZjX93I+PWtsFo7YKahBog/Hw6Vh7VboAq5tcpK8y8/3
svEkRtKaMWviub207QL5Wy9taBT+ggiDYD3CkRuc3c/4y6eYSl0Ch1Gm/YRzC44ScJM1grhPNyz0
85dfjcf9Atk44NpagM75PeqFWOYjwkNDsz9AL1j+jr0lcEhBz3nlwYYC8ACpRb6lTKZJVfz5Twy3
2qMlW+UazmlsQrp/d5ehY6cCaCesPPJg8cGMQbhgO97TsaT23q/I9VITzieMi2VMWRzb5PjgYUh/
MgfBgzxRRnol/WamuCuz6WsA+lisq7bYL3jvcf36o2/SQyc5xfL0susMH8WpT5c0hLygwlsrXNXS
N2mwQ0rGmLTB65whHS2I1B2xD6XEAer1Jv5ffAC6XpJejJO3+uQe3cAGLYMnpMZJ+Z8RKT+6JGNV
u7/pc9NavCboMqrhJiCbBBs+25Z/Sb2ARI8p7nSGLD6aRSTXSzNH146Iibuq2Qvm4DCMzcd2cAVI
Xi1rXxARVyncUWlRBTyVMtwe9N4RDYh2vpANizapYny0u06+02lunE4XD6JPBmNTJMTaLp+bpnDV
PYpDH5mY2xBJv4jL9o7RT3qGqq7yu7fJ71ti6ImBXsYWATxID2QZvkEk5eqj9ARVaYVKViykmPoS
weeihg6eMW57NZ13GVRfHW/vAFjPJesFcA6b+2YUJkygRq3Qo+INnh/yuTy5Rgz8Uwl0M6+qW35n
lytNXT8KcoNSe0U5I+2TtqtRZ6cctCalkMgi7m/0ytiPApuOW+XtBqbjEGTVnRmTtmXPAD46q0pH
dQPgn4fvTnlG0kuQB0DPQDiBJyPWWOqx1KoW5ymnXAEDUJnBBsrELoWDUhzzmD84o9ooLxIppFq3
yJ/ARvqB5juF21ecTuhazlGGfx6qwk6Shh+H5ISKqAjHNya0RVtbExvsO8BqlogWaVBb8OJDBVLo
zEwS2UwvZ/rR51Tk3vu0Q3+8wVwy6C4TllK5TkT9mKlooL8RoCeEYGasYZ7yTjFR7BrONC/yfFGC
wsZFhJ0Ku2YddCPjEDIMIrhXz42MczF3RYd51ZqWAbT4mZhTkG9r4A6/HQTfWxlfX2cjk1IfhHTX
MN9cr2bBsZL1mheQYreYiAVd1xCxmK8oF8E4UD1cQgX3TbuAYiUqgOQ/MLg99WswY335X/WyhrXU
0gJTSt/1B5Gvf6CPRXjaxdKEzrZbcJ4OIoEEvZbqJTIGstUXrQRwAL6nKn1LV9iaBLbqBfWCslzq
+Y+Szm67FuhCAfZg3zd+SxZ/1/NDWwYuEfA0h2a6KUcJcYKnWnF7pvkBeQb4IOy9a3lNqucEhfnU
vpWF1hoPi8zY2EbaDCbRJFvo26AzUVQB6Ezd0f5KVJhJdKB/4NGWyzX31RuneIg2Us76hMLAVX1V
1Fl8gYMtb+3yfLGkSJRt7me8/M9ayD9M7/KFktkuocOTAru4QCAp3MfS3H4tlt5ss3H8vv9Nb8oU
6KfnbP0nmm10o3bxz8QBirACKAhsAnL6jEagn5rCJHNvjiQi//sZUp/mN2lSQxJhUQOn/VYL2wjC
eD/ogAPAIRlsqNp6ISFHuGBdhfz0bPFgW/ueCv3H1s4wPe9bzm77dbb0Z+lB3idSPI7hhNrAfCAK
xYLNjvwdzG5u/DzF/XPLVCPgqmIfMncFR2SHosp+sldek1W4rzhzeonfQIDpOVi1lXKcjPMTK8Q4
TkpWFqEPFwTbMRZHoeUjfMheyPKzSPcS5gQkdjwahElSLi3sx5CSdMhr/wm2ojW7OfYgLa3Z5LDD
IJrWzkeIgq1RrKSeYc2uvpGaIxPKbkp5RYx632p0OTBDzW8UoHgdqBYXaeiJqaSL+tCz/b2vTBYd
CSnhfybq4UjbEn6w0yXo1CnTxSpUH4d3iC9OsE+RtnmeGevFVWcMsnE6DLo7FInOsgJlgsZhEtcQ
IRumtWoMxbg9LNrujQ5BaC5HOLsVlN/9ISOa9ZwvkTCS7MHdmhmnlO/Thup+qn92GbAF9V6Bl7/X
7tYJI4lxDrzurFURmXKTtUW8NgTD2JyfVOChUnvouUwTtKC0imGWW4oUf7LOdUQkdoIZT2StX25V
TrtgjYandOAxmwnpcQFzUwq0wcn3xACNxnWt2qasR3NHuvVTyiIHJgU4qNN73SLjCrecCJCbn9ki
kYpNfp1RMg0hO2ick4rNXnymSC4AsnBgLbiXSSK4mvfc6GOX5gTJWVm1F9J2g5vuVJAHLsWxtzm3
3Hkoou4H/3JIiXC1RBlygVJgMyo+//L5VH2N8MlVd+omSEssdh+HKjk/YLYqaNw7g8ujyjUpkHUz
Uxs4sxNvi5nsFd87ouCEY/b+LRqKNzwqAhMH4AwQjjVQEZHVsk9rpeJrASqmBt/R9Wj8JBC4rzxb
XVXC2XAexNlv55aZ/7VzcsYLNNIS5M438FZFoRPLUZjzDJzk5BD0UnMxQt0elTXWcimqPBJkW9Yl
Hrfrfg6dRCkVhct9LMIWaxXAUSxsRJYU6fOlW0OK03ZeLiQZkBYR4C4Ne08SwwyDBs50d/U7buCi
pk3UZvsPsZxXFHW/j0zF1HWvqKZhSVqT0Negy/EViSyBee1fm9gWyn5heblt3V570NqeuQ1Lo0P9
DptMzHmWpZdFeKny6zJRbxuAzYjV22zATxWGLORJo4isN92u7Arkw+5Kjul/TPsAhg2Kwlj1Z0U/
u8tJYZ1Sv/23Nl7CV4zaigHQnMCQLNXcNE1pqff9Vc4UbwsZX7R6DnyNOcvETiwdzSTC3Xw9lS5v
6aFhabPMmouTXeXPD/v/CsvFMriVI6qvY2Ri+ZGulgQj3CGsRdkyDa7Zk5pXiT1Davj++KeFLr83
f4t7d/PGTCGT5PfTt04CFLRkXS5reK3jC84VkeO/xSfcLCEylm2mJJlSG4EyOVtFbTTrlbeGwToA
DOwNxrLkGg3Jy6oyCb2dYfV58Ss7TE2uTh9pNfIOzrbVFG7PUY1VnDVvfQEehFyA5YmzEbRiy5i4
yOHPlaMvgR6sBVcNm86kL5bPmmbcJakEnLBWuzGpcqwial1Uh6WAOqAWXgNZvWkB7/KbxC3myGWz
zf9CUD35UuXqMTQNUxHayS6bnNEO0cfqaOj5drGS7huxGoOmyJIYbaPa7upwQ4ZpbisV4iuHNt7Z
ZDrcTbczvtwiihwFME/IJWvTURZ8VipWMp3TKbNCWaqunjejNSWZm0yX1Hbisxxpl7ewRlx90akv
RuRXyb4sCbPYgTP9ylIzeavzrBtQxjhouzPkB9jsI4VDbzAVzgH5pOHRWhxeQdn/bMCy2KL/ac8O
w/XteklWJVHkXsOuaylhpZ36aQX2SO7hsGiUZn7aB5yvD96nl8gAJrdO2ix1hhcjwsVVxE00Dnvw
vhhdKPkhJY7dMOmdPOGQl96Ci82ZuOw155GJW71mTT0l6sRTwyCu1Q8fXg5cnwWkYuJg1zLt9ZOJ
k7x3Y/Rb5Bt+AE128Ze5+ddqRtXXgvKzS9dwu30+Dg/uC9j69BOXUiOPbt3uxY86ik+tcMTR8ToI
TIkeD0GbJ3wUJizfP3pzUvHQEAM7YfTFk7kgMI4UU1PIXmk68pkmPN7bnNx/QNUZTSsfIgSP96iz
YYFTneR8bt+5YaTa2DMvknyyACvv4AGg2aaWdTVSZCHV0Dpg7HfkycnNsoGlKAi1oHQt7cFXASUq
biS/pEACTqbO4o0s5ARSMApr6+nJ0kbJ8SbjosbXE6lVsdT7jgtqdjN9Q4qaqFlV/2ttjO9ePP2R
4PXOdM4MIAskZInR6zOn+NEE+pD/8d0ubU61QPi5YSyRrA1IQKr5CvXYSyAyp60ha/idJJOpBtEp
JWEdJuxgXCnl6HXWz1Tdhhht875OX6B88DdUJH2nqoPX2k1fgR3Bnq5h2NLUo7G0vVGrTS97bm0U
+YL62t5+LRIiEhiHkTjLf+UWSFmhwH2b8tnV4UcR44gq01SrOWLNhLOUabXV1KoPVSxws7ZZkobx
3py4OxPTq9xPak6XAI73EOfUkaF//Z0lglX87MGY7k3HJ4yHpoB0adyEUcghrp61dt1l+x3ZI6+R
AmdadtrG+bn35OAJZu3amgjgx6CAuQz6KzDoTns1o/mjNHU0aVeVavJtmgFDkTEHRVgG/rINRU14
9ZtN8duOB90iYU/AlXQ2IkMZ5KHVnOuP3usSnckrVYyrYb4uU4cBHKy41PtzokkpkVj0//4m11rq
SB2PVI6wu0msjORS0aCdd/xX2UP9WRYZCl32Ck/XBXEg0UVWNTRnZVXqU7XS0Mk0MCpANfqSOmrW
tkCheW1rppQ+Ffh8LuA6J10RrkKdksgGJBmfoWsE59POQ62e86VDom/4QiphmyxwfkBSW9rfZo2q
FIB/kgxgqhWPOW4YS1gd0zTjhOrOhTGeanKFDYWYDiO2iX01vtNVybiyCAXuuxpUVD3+YznmbQF0
zVP2JDdyT+iLcKKRrG//WbFi+XsNlZmB4+RQuPcFjJtd/B6zRQdz/1JZmKCClYydXCTMiKo/tttE
Kpc4z6UY//1MnuDjLgJ10OXiw0AG3ZYmVLMmhdMq3u3l8cDyUZ6F8mmbzgmISQP8oJaj54VUMMYI
ex5lre4+yTS+tECCWjRCM+yp8qG3fn69o0bdplyH2jD15l+vxdXifkrFTSwfx/MpZZWkGiGhY9IZ
m0L+ughvCf3sHeZ/2vVth1nH9kg6TkhpjtAIh+NcGGQfc2abmHFYfOBC1yyVaG5Ni9OUqDU9jKr9
tQKFLlt/bwUT2qRjiuTPVkZD5QtmUMhEdIo9LgTWDzmOzJ/jLuvuqNUSE1UEsTu2zKuIJwuhay6w
nKAhGq5KmdtyQxRqte2I2feUGuWdL5snJJmlVG8uJ4IjH1aPHAjXdcliHCx88D+R2PUFB5pEbnkY
Jq7ENBf+DPKrfZdYGFhyXYsTpuAE52iwuPd3r/3cWmGdMQu4c3CqMDp0miVx8+77jHZ36JhXUi1x
ImlrP8EZwSbaH+jTEDdngVfVYtWizPWRe3ofiFTb6DqoGhZ6l6y2x6dJmWDYJdCP0VP1tUeMDCZi
ifaqVRAumXpBlRyP/1FkItyQq1QdqzpenyPfmfGp41Z6Skm5EZPw4hXtvv/V+RlhPbPldMGFA76h
4b7lCiViCEJbtlyVTNaudk+B6cLlvMI1XpvboaegGt2hXRqvX+RIXEvhMdef79GHT3Q8BzLsSzEC
T833rF7mbs88GRdG1qsjI9yElUhJReQEJxGWKX4+sFHxWo2Lf+G+3gMPiXvOIsImynbD7vd6f5bm
q0AqOL0LLAjUe/5qtsMeLmaCiLi+yP8h99gpzl8IsE08Df5b5awahSfZipo0gmVhGKeY0jBzRmxF
OB3i51h6q4asJ1bsqANYIPGzNEjG4ltTu/77QBlHozJu2VtAw6lS84kq5R9mUP047JL4fS/92pXF
Y9R8xFwtHe5gyn6xTH16RuW+GfKzDOBWnXBwou5tI3flE4rcBQKm1NMEzvRX2QvQcB9EmN95tHpG
x900skfOslff/6X06NIdzBN5ahek1Rh9hZVgmAB/mDddM8mLhhRhb2qTVyc4vJGTg6WJ2PDs1s2+
FfHeXd2xm598UNpEJ8IOnVdoQTPjiiU9JbNA2jQCdSOfW9tCn3dqgYMouvozozjxu99wrU9WD9qI
FRyCYie+6/QybTSafqEnYq5ltjH+9IvdUc729LYqqqBVInCeY6KFW6XRyWn3ngfDbHC018uj46cg
jUUSi41Z2+HsqzKmJSGbRdkXDt949UpwqPrMKGUfnRggIXCA7ibu2DZp5tY7sqgVZGBKTottOoSN
EdydiaXPj+MTap8kPmFODooqzgVP/kISy894yX8RpR9OwdrIGPg3CBuIbtQ1m+gOIIi+1BkQHa4X
MZ4PClsNb/xLE0D9Ap6fXVL0GGs5SQg+AQ1BiarhxZ61V4Z20tonvetGPCsH63qhn+Rt1VmXjPm3
NXzzK9YURLPEYFVUCbCoEXFT1R0GcD7iGn96Dr+U9x0tdXZQHZgtO6UZtIyJYWyHP8TwLAhEqdIq
XaXJxbDzvHYYC5Zdbsgk7iultDd3lWWZlkPHrj+epjL0UIytKUmJuQieCf2MBl9+2PkQ0/m0NV97
eR2oOUt+nkYwpNcj4P0eLPhJxK+DXOQi+L0vyYj4csDKJBBHQeCuk5507PJtirWu5BYTUsuUQ1KT
6ua8p2tXRbpHLyeImkKQcn3l8/ixn8euvjSTiuJILBzXnzhkvMETSUbiHT1ItrcrQpBmEEGUb8Wh
9boMXNHzJUZ6GnoFmuHi+jCKH3uDuIrLFoQXI9pIf7yFQ5AflCJ5brEgGQYuk5l3nx2SBXNuH9Ak
FQ9EvQ/KKTdKdI88wZUiDH7QROFLdrQnK22v8imKL9fhOTGOo0X0Hlj3PLMnW0ApZHL2zZOZ9C8x
OluKDtyokE2HuEbreUwQE3aNzSA5Owjp3I/Ik1cG4ucgc+CGx1Gt4hGHQNYII3YnkJLsG/Y3Vhrz
b01xjljLNAradOu5LlSjUz7/pClybK/h86AJUt11fmP71P5Vr4Rsn042/2af3wPkiL/9rbLlLC0P
6YshzOG17p3h//CC6Y4ocbiN8sY4N94fZYxxzR6l3/FthOjacq5CTDy92WAwuI2hmo4Q85pOs2bd
p1xOqnbPHzaGEqrDiz4Un0Mw+g2vxKnPkIBY0uZYD1UEoyeSq1/gLFgHKpuK/blxg1VWlihVdb00
tziIPeBdpnv5Y8eROBE/grpGyH2aR/qokQeakn0lswcN4Q6anE5QZ5rGebXaXLby3Rrn6oGjHq2h
YRVLkLU5C6QfQffZi7nRL04cfmrmeWSH2jBhArjY7QkNFPcij+xo2jdDcxE/wxMXzPJ/iuEMD4f9
i0FY4eSv1BMti7R62R8dObENv3CIlAfsSboKK2IwOOy69xATQ0kG1gvJpxQMUiSO6k+2JgnEn1t4
wCf2HbWNp7/mze3DuYMWX+7kNdNySBVvX5PykzE0QQtDD30RPzANad7hn5iXzB3AZZu1MUmaDjzy
Br71cSb+3Nr4Ft7u/e0tX5r3m7ay8k+lJlQHLYAnkWvXw61a1h3aDOYHJ/eNh9gZiGs7BCvfJ0UJ
v7flGLz0+bVub8ykoqEC8MXuvAHOho3f3c1Gj9wwgHPQT8jKTvuEGDgDw3zKgR2VLV45ReT4pM3R
yonWftS4QBH/snKuc5NdPniIFmHWjyltm/g6NDc/73jyCg3pYWTMJS0QlvvMlNLokaw+0XtI5L7T
iv2v5bPiG4/3T+LZxAh+/TaxbigiSnONn04jfhpqFz8z7WlIJFwyNdEjGx0Hxb38MZ9fqxqs+El+
CXJfLwiFBNAUjITxZU/YE4fmT1vMznP4AxHI6p3A6AFLpRy3p1O5OPAzd4fkH6zf+rmGTRTcV40f
H4UwAULW7tz1KGcyCjMIhiOSaKHhIdZeMhA8TATlq6iajur6JRRS1PaGxazFu6Fs5fQsedannYvb
Lvz6akmJ+IjBSh0bwIkD1OTVkAtt+wxzLM1FgnPOabLZ9A0fVkOYf8n5hr8Xqh8NLtGdT55XCd04
02gyi9OCAAce7dEoXxaYYK3+ZImqPnntU4wUiLqzpCuJcoIGlfgjLC2BdOdcPkm4hqLwTnfkSASR
EsznyDLC2Y30RVrhiqp9axWE1fm5EPnAt3jMBMNZUBzudOo7rlMDvTD1Vt03kNVoAkPeLqGIAwJ/
nDQKT+iAwpml7KG5okoRuBYhXeXfQJnB8rMBkX6aUOB8sN8IZ9vUDMmbdpnFnvb0DWPE2Aog0H1X
BbhDZR+wna5MhUWZS66E02C6kTImFG6pmQM5WVJQ/A3PFKyXjGEe9R5+5tFRQ2kXDsw160WVHjsu
9IjbtiHZd88mrrkepTQ9xVXrTYhMgLk2jLHfP1JhSpLxsPyVJYQM87tupKyuDditkRjVd80YVfkZ
1D6wND9NvcPGFuxvIpVmCq8NICSBbE4Mas1lkIeUenjFONPPmt1SPYZJsyevw14eXux2E0J530Pt
LbmDRI5xBWnp+vu1p4buUN0JqMY9G1IrOhNRwDrcsChIA82c1QxfPq1WGGcoTrHardtVHhwYdpoj
Y1YqYv3Ekut+vX8dBh6fTzW1GW9Be7WzECQkUN1TMTL32Rb8DrK49liDYdA6Bjqa5fN5qCOGVRK4
2MNw6SeRIXMpQCIC58qi84E6uwEh0ATOpatEa3auhwetPsgILlOS9M4m3N6dDX7LqLwLgAkyXpkq
aAiu2vf9kyfxkB/S0bdApm0rmEyJX2FSZ1ZoDK6t6Zt35vVznn+GCoLL3J/s3mXce4iSEkQx9189
6Y/M67Z4hJ9/NJ/1Pbni5cBqVnVPadQXEYP+I8UAWrOWJyMvhmsfMY2A0iOmKyk28yIbT1SjJyg+
hUdnhoMuG3t8n+H9fn/qEqSHCv+mBHP0H5qoxNGgG8Dhex0jYGn+j7+5gRCHLI2W5gm05T5jhkvZ
G2soJxs8sJgp1dPWzLdCNbP6tlWt6x7xtwDMOuvx0jJvKajBWTtNNeMZi8udBUndXwXeQOf9Njx6
mYmOBDiSQofqVDYYYfe4tetEzIVcde3D7odEKBr5wOFKIbWeiI3kg84P5j2o0Ic0Gab5whW0pcLw
LuaN441vXRAsc+aJ0qhE5r8cKwXf2QlQX6vSRzPbVDftwzS4xYan0X0a/eNvROrQ75BArIJMrxwK
Pbd8gPSv0UaVIRepa7TvXjwkDS2J7zESyp4UV+8Cq/0y1MUWLWxpVLFaeajRQDGx/T0MT1bppXle
0tCKbSzq0z52BOpw6bSgeIhEeEl2oSB7rRnX2ZSxHrHVfoLvI/YbMQZWK8mt4FP41/h7VigrPLzr
NpYCS3wGYWpoIMfatyJ37Ali4ozEMDsEjyCH/zvp6j6EHUolFgzvCxUFcXXSCb1nA58NWaTOX+76
6NgOvxtaL+LSYVPJslaPNprdmoSBNDra8dtT4kzRHdwotcQx/Z2kTVC2HtiLrVSSoJJSao7kQe01
EQ0pubS8pB+G1AJH8j/yn4GI1hecLyx/m6OsJ6I0C0mB2HIhRqkTMcqb71SQozq4pDRq1XaxGXDL
KaYSErQpCTBP6iJYJ/eCDEFLNf0CrfPL1sYiunWgBQBNfXNn8qWvdbAGhjFz2dPa5D09HOB6Vyj7
CkideIdvS58jixjy9fck6MvoENMG8++Q97xuG+R3p8PYW2sgqPNd91zs5y8+nYXOjjat23UMbwfi
NNrl3BmaMplky17obMJL9ykP91rImptYSB7MgpwvNc/JwDfpLJyuNgay15p/a/mqAdX8JPG3Ff10
umZb5ayeFuNlKF12RYmMie40woqngjjiN3C+3mplu7RzwVKoWcY85PAjs52ggdmPuhjeg0ECYzsG
sqHoNtyru52RK6DrY4n8qKPKRDdk741G9Mow3dEYWEEGncvyJjDeiafla4QWYu8O3J+hh3NJKyAF
YbVI7ymZ1D2Jtie9PAX8xB4L+MmD7gRiteXnkYmUhHroaDlRYzioYr/19QAY2NfLD8bDyIfgsYxY
kFIwxDIjaujX+oeyrUJam1BOWcEzRt6qtX9FXINyKNlKddGdCqRF/A6TfVJ01wCvcTHylYR48yO6
j6frP6TPeOjDqgHSDySQu6FiZW4bphkA6Zx7qmg54CALoYqQT2YpJTWqF0XxsOu0fCCVv3rAP+aw
qVZNj5xzO5NzTxfUwDId8c8vzVr/oWycPxjgg9PlTONBV+d+BZrnMj8c6RU0zqTSjmiMKfGsUHI4
LM2MIfREJU83cy3S5+K7YJ/PQLsX41S82+gl6ViJp99EtB0qMhPpqxT5bc8aaPtmM8BbwRjxxY4T
o683DKBCvVwPVfPiABperQ/SpUalc56EIAw/N+huaL7c0BUbDRSDX748o/x3M/dnHigG+64uavvW
Tg7+USxIuYFZRw/yol1aGvjNch1c3ye4Id6lZ3T21xuPYVVmLaW2KhzWHgLLrUCiZxFy5W/HpR44
WqXny4tPSsuqMW6iGIqcdqHqkZx9A6uB5KH+5sX+4/6minjWl89nqMDJeim3ANGDa3EHU7jAv4Hp
Ks29JXVHFu0YpB8OwR58MuhYpBl3ZD54oD0R4ftSASig04Arq2keC2F0G28rYH1SFb5t2grO+cO2
5rlHABgwSaoBjeHmViUL5EeLX1x5kgA8SutWuCH0WeAMhuKCCUouo3bs+l8010R2EyIzDz80kuL5
E4bVOt1hOcc5+inf0WwymXYI3lzxpTvEmjKCM93nQqqbYHIcrK0rO6fK0p7TqWz3zgjyaW8zP8Q4
s6n5t8235WItrfxQa8L+G/hcouBm3NEuNG2AMGYeV2oHpUV8FK4e804F2tiJ5Kx21VrJCqP0PTNa
scsuoGdAP6ZzQz90g8B0A5rK2GpFw99IbccIoeJa8swl/JbdVBz/mxUVBFE7fTAdHsUUveH/+3iZ
5hz48KcX0mspl+3C3S378DIR/apZ6VRJtsNb7/tFMlfnhw8DSrxr43GFDllwzn1+0kSook5b9QwM
LdklhGsU4FmKLvfO0lSKnC1HpxgvRZqSaHrJ2eNPZEzWBn4378He8dcgreLNNcQo1wp23hrqkAGY
6vZjyXal1g69JI5DSs9v9lmFtQEf1vbYiG14+ofLrgythBHsUKmAXRRQpAbRQ1XU0JDY49ALxXfA
T2kk7yXZ+CfBkNDbzXrWo5jvLTutefTyESTT+7Ni0kxPLK0pol+6BUGxp5Sqql067hlgR+Lv4O7T
9jtUuBGkknkvjY+903ruqsJD5f+VfDrDCta79GsWV2onqL7UyoR3868GKiZMZoiPXOJzvzxCS3jN
GBkcco95OkV9QAsUIbuX1y3SjX+g2KmczZARKeK2dAYZff196vy4Iezsu0fAoCOCE/vqllcV2IwH
uZ0xS0ePmD22Rj7zuri/uEANb5key/CdFAYm+ijkefbvXeH50GdfNyIU8zbY3lpegZdeI0K4ZM5m
LwRLF8ict5T7cGtQAaFidPknNsb1mlvzJD+tBQDyCehT28HQsFc5th9Nv9XPZ8Gpvz6KaWv577zX
L8kKgefra6vq84xbndiOonzS/x9l9hvCq3j8hQdMxqOOXhox9egbpkLScww8zxebo24LZFd5JElk
zF1MRolFZydrBgi9s/EfwXjzV3l3voXG+bp5s3HGBF6IUH5NeQO15t9RYmhE6d0D4TdZFwH9yxpF
XvwXQyvUMSeUPCHNl29qewKuEln1GpZ5Oj5hlBf7lbyubHS0iOyUDwosgqMP5Di97d+PEXhVuyv8
EBkbd+BwMcv/MlpXC3/VeRg6ePQBROd++2myqG3AzrKd1l4Evlp/Cat8KFRhoytTbZRD8LS01P+A
U3EDZo/7fxhRG/X7Jj4zhAmwVdMKyPll7HnAjf/DNh1vU6lD1O6T1R3AQRHam2HtLCENkq92/pC3
CUsC6qKHokJhmSBzLAK6V4+bxXTobLuoeZk++wimb6VeCQwFk/2J7IwDFf83p42S+eGiJH5NYhSc
1tNL0NxcC2heUGjIVx3SrEO7ptKSzCWbVrEcyfn7m2ul0HST/nBpPZK6VxQQ9x6rH0pQAr6Ggc+W
tBAYOeN0fljXfCf3Z6dkIyg6tVwurX16O+r7fXfPUMGWDumkwlugCY4cgoK6ZiTHsEH3BubjzhsK
X3WEfKV21s1+OZA7upFYQT9rcV+o/Xv+Iy22SZMgUSaHOMfKnvXpj0cAFFzspP/AtcLnYt9LPNl8
E4x0OOrdOOie+PYB3LwLPZtisOQqkDfJdDxEDYSyGSLSpxH+g5q4tNwr1oSpx/Mh0/xWlNiyQudg
cO3zFJbYugcaubbbZj2kUphgfD0GYb4Zh2z0y6kTa1QjXHEwQxEiClRiuiWnr57zx8PQoI65547r
1UKCYpFgl2W+zy+PfYO/G6Gyfuzc5l6UxCQgtAvla9qRImontwthODI6NzFMiTvbW2pobx16h5G+
8pS1tT7RMVmupp9iX3W+KodDD0W3gae5/6m3csMD2MA0IhLjydyPqBi33zAvyQpo20v9HSHrvuUq
dCdx9d6mhXAmnzv+2hefKa3HyNgyd00U5bIOnEr8ueLTvEYIglr6SXwuaBlUNujGEKbvLewk333i
P8xhLHX4k0SmW+cyGfhrFDCAJG4x0Cs2eMd8gnT4/K62idH/3av6TZsQBjV/S7X6Nauogc9FYJeV
K8E0jMLJkX9froSLeUoVpS/Ea4BHGOQItuatzqIGsl6s2PAr8HXI7kNKVSBEYKKJlfaIDSY6YAhB
9FsM66XOx8oD5rQoNJKKTuvc4cGyqWADfsRmC+lNLmjLdypZzZ8jgowxPG24zl7c7bb1+XiiJ3QU
Vu7rk+aXCZ/D+PTpKBVsg/tPpHuEnvAEbMn+dkt67V944GFjUS2mCI3UXNjEQ+M0t/iDcRkwO3la
gWd3pf6YrhQcnm7F3sWzk7SWAhhONAax0n09frk4KKGfVxNgH8/HPbPyopyDsSKYaqf1cvVRng75
21uq0qjm7bm5tlegc3qLPwro4wr6xxmrezrmwy+0UcprAmSbYzxBonwXhKPO/Vq8Otx8bi/hhVlR
M0Ymz1NsZBn84vyMGne3rTTgkYPzkEWoCUmqX8OiXVAazfmBPqOqMK9vM1YUhV/5F2UFydr4pE6j
abXFhcaUTJ0mcm9tdvxiohnVXe5MjgtY0bvxYq435Moz11AJPk6Uej/qveU7vCDWn0R1YlgbTWq3
beuwTS53A1t/xc3iAb4zyHaUvZfFpuPZg6kiCoaKrsxb/AxhzmzrIhnATWJwG9QmA37Cxfz78mLz
uKeOilAhZUtLxIEUc5JknkcvvbiSaCPpD9FoysCexgzIbQXHWu4II8HlhJJMQkBSvbGAOrAsQdEc
agNI5o56J2zVHyw54vjaTd3NRXXwF2BNAQuvVDVIDQnsBzc/cqYFub91eYfox3CmU+3wp+68SXyU
q/qY3dTigsOQCumGfqLJJbiGATWcmTTRuRHTmBuTbm7oQlHBLAaVmbeS6+4drkQFB2O43NAeoozp
/oYxFnW1F17Ie5QBryf6imQHqFZ9WTYVs4Df7dXO5dRSFiyBKoWrXkthSzF4rA7yo+Z2UZ3r7h94
j/FyNE00hNHEbIU9WaD6yqC4RaWc0QduPD9QdDUD7UnWw/nsEgojMVpgeVZa82viAA1VVqjq5hPs
k4coc+kxt/8C26g5KR76vq7UPO7AtHbHqPDuaykzv/lLVIYQYCUlcHosqtR22M6g8Bg0kln89PDX
C5s5rYsWS9E5RqzNgK0iIS4pdk3XxaF5/tb3psiCyAc1xq4o4agtsKW8XpB1Sxaw2zaGwH0udltm
k5Bxxinvx73oHGWdmXPwbDJtHxbG2JU/T4ltmwhLr5ivam7xmmTzq+9Fl90PZuwX88qDkZL/oIZR
mI0b8ZChT8iOlJREr6UUbZJ3HMlK4y5O5PsMprAL8RHm+18dL4elrpXoM3dLlbBi65qOkqZUvsWO
nm2UvphZQwmuc5AlO3hTRylzeWR4aKDqtAVb1hivqAHMimD4VuWXVz5iunFgXZsnXN7B3SyBSO36
vbxmCrLUeqRzV+7KwMpOH3BW6iVnpxFukI0q/BLKUNu/L/TjAm8SM5GQNobQIcoQydLGuRjOOx0T
v/dDsdtMRmXSEdoND/R1+97lQBfDMZ3drWPGdqaJhlZnC1jxQxooHw3MN0DGV8T3DmKO7d7dNMEG
fCTux0YejTptTlonccsmTDOcGJb6hSDfotJWiEGYf/oQB2ZaFQJtfuresK6dQjtbteHGQ9L2d9ju
Et2Q628wDI78gOW/Fr4VTYOUdjTkiJIsa/2URbBR8DJEcm/ZOYmOMTuymI+drY2t1S9+4umCAvBP
YusatovuV6Md9mOzAht5NR8nSfJsH0JxjgakZagWcngIU0yjjJFLnd7paTDgNipSTf/3/cm50IPy
05zuOctG+GNfG4GBFabBYltVtP1laERTaXIklx4oOL/S/ao4e44HHFeoX+a/95TOx/hpqRB1PB5s
7Xm3DSRkyJWrY68XCf3NxI4w1DlOjWbAoHoS2lZiFohttUNUMl6NXUO8blLypjGM4QbMPLsip3VA
97XM5vc6XqPqCY5i8chLkh4d7IjQhh9wPRUTP4eGYtcMECOMetaLooho/QYCwFYD0eMeksn9kFCO
XHaDMy60VLAiqflVgOEod5es0mhLGLJtLco3s2bCaUPGaWeJD5FJbd/I9dUVosZon6pZ7T9guPhw
wuQfbO5/fKB+ForSERsDBiXJRwmTAUfNd+nhoK61rEtKnTkjnBmuYD7smEBjMJg1OYxMdNP3O9aI
QNeL6Q1LGnIOjZK5TLDqm0sHvHeSxSHCZ85ToCzT4nyjttvuOaixxS6PaRqSpJy5aKZKhjb5AZpm
bfKfRW1FzYMxHasBAFgOKS48WmDA/8rXawaitRjPEi41Styhf5c9TTYxMCkFSkrR4A3Pxe9621HG
qtA6Wa2Ub5DtreiMBRWxITFYuR2cQGk4dHs/5g3rcTcrpBYlZJMQkQvuoMIRH9+QRlfzC3NgF+So
57UURjh5Vdy8nIIdeRBvY6viVPQmsjzYho/iinBSsQSpyXHh7/DxVHqHJ1MiwtBLiUETRCltMHZW
hunKZ0HgYISszIV20x9woYHGHBo/40ScJnVhDqbZj6/BoFhomNa2vjmK2NINqa47jwjIc+t3aQaQ
DDHU3bNP2mLe5dykZ7QDBNq30nK/6H6QF9p3XqZS+NvrLEUUCr59QyEcL1nhr1+X5/TWktyPQzzx
p6HPdYjA4tXd9I6NnHjv0yF+H/c1wtTpJ74thAYaMM4z/EiHxOnRjO8f41iXN8P3ToG+NYy7VXA4
g77Ab/84+Bid66SRjT/CXY1XB8mW7foHLxkogafyGFxoWQT1kN+ysuf8zU6NbGZmrKcveefxfKJ2
HEXwkSQSlY7iBqgAme2zNkhOcgYJV/5J6cf9K+/29fU4hBGqhAo9YxXbeC9zuqRix7Bl61+PExUt
vFfvd82uSbD4ZdhAYhD4h0A5RRJfDYi0JgBtNFYsfe5XwrZN2ZQDpspogGvHDR51IWVNXHI47xX8
8pcJr86ruX5RCOhqSYZTZipxnwSqu+jNidKSOoHB4hxqvm6GrpZtN928Ooy6pdqsRiKaX/0gsYw5
IQb7b9V/MALvnS5EM+lC+CFtJ2E5LS8qQ/uBM/TlctSonxsfKf/B8XG/X+3kAHW79TXSSWdUUeA5
2ObRJ6N7NHj8wd3acsef6gaJO5cVfLeCTZPHFLYDfE0eCu2Tk188iq3wKNUtEzjaVOC2kGbXqPIj
hSmGCoXAmdsJ4mHjeahJ/pJ1/3RDHfEtz3OWfyzW8I7by8aSt7kpC/jSHdd9du1F10SCzCPgyM7o
3j5fXEhfWhLXEL9EGoaFLcFR+/ntl9y3IGyykxOIHnf6oFK9uP/a62Vc8yjzLrCDToHCguH2auV+
A3twtK+cj8IxEy/xDL619BtD/mUVLXBF9cEG/jdIOcU35Wy0mVXBROknbZ+KcN51pG7rIlEu8Yu8
+Bq+iS75ENZJglcJduzYzCUHzjzWCTq4GTedv2WREin8nY9HbpidfCMYo+8pwduMi5k04h2VgDt/
HtsuyrQbGMVd2UxZ2heAYBflfmaxJg6QetbWGYNvT85OL7FTiFBr8CNJ5VCxp79+oiAKnFIwRNYn
c7EIr7MjKjOSiOri0Am+Tu9JC5HBH0LyT4MJQxJWTUXR0Mjb+KgM9q7uDteF8pGeU39alyC2ONyp
LtkoqfWaJIM2zd0Ti48Ubj06I+QM565AAERGdfrEtvm3vgQlb7DBPhn2hRZnxlv4CPZi6YFf1F/L
rc/pR1ABBpHKBos4gIV4YV9Z41PX6kX/x/FmJLZxsGZR/mgQiCJaSeyUnwK2YtADaU+aaQ9qMZhm
f87VWulqhiMFz/stgQKhIa9YEQ2ijsWIGg98Yyeg9gpxy887jnf/fbaxcqyDupRHzuixHSQ7b21B
BXIR6Yv3w02tutfdjeWQSxjE+TSqyqd2QEUkyl6C9sOWGjcRtYP3ZZ0nKYpPb2Gy7sIfmTd+CnJt
l90jdX3ZGuo33pqSXCSUoY4nBWp6TvlZwMj+Br50bv6bxaW4jo+z6cr5tcZ/HXWTgc8MXZyhJabk
5ZrNGaGLTTrmom5HF0u8uq+q9we+Q7Q7oG/nXMpJzIYDVX82+JmDL1mdvoXXOP05sstB0E9k2NjA
W7hS5LMoUZxItiiQQCubM3vv66GoQl0T3HTnZDuCEZiibM+ccFiiBsbtyv7WC+bQ38CxovEUvu5D
+S48ImUmyt37fSr1oSOdXg1x5OO/3HxTivgPQdNnXeiFWZFuE62NnZh4fBs3CeBfq3qjVd45hArk
7BPNyzfoEGXf/s184A6wTE7nrnS1uuIAwi5c1UJMSB6BnwsHfF1E5c4iZIrkmu8AdgxMPI6eqh9r
25ubkPEZHu4/WT9XmMZtuBDTwNVcSZnhC0Y/QWPDZCV9Sxb9Z3yxvLv1z1Y8aJxB5YpMVT2w6r0x
YzIK0EKi+PzaVDlzlnu8a5QbBFuI+sqvTpaX4Ij2QZDXD35LXP67IHLygBAvvUOZBxCLiHB+oBM3
RH4J1DfO5zaDs9jLUMkrTRL8pr5ba43YFwfjySx5neLwjO7InOKhwEGvpmt0m1UtjUv06cNBsDnr
53FJZq3npmeZRSEhJ0t7npgPcaM34T3AAbb6yODkR/KqYCZNYqKSgdkKkY+WGqlE1nDuBy5zDZRR
LxHYlruxdfgyGGlKhwi5hVXfeZffaqwTG0pix17BBonM1g4tVGnlU9NCph8rfTRTExq8/9bf0wcB
GJD4W8S4XVY/698yKj+PaLZ0CTDzDWMVqRkQYYass9TCByXN/4aHWbz5UUsU9oVKR/AZlsgz1LB6
QIKd4LVpidQvvSbOBkLkW3Yvc/BIv6KRN0On2XduLw2rbLYvPki6DHR8vA9oBQqPauXZcxJU9zpV
nMFFOgBG+F4ca8q3H5wQbNgdm7xgU9CBSfWkW3Gf8aVGAkd3PGHVxkxMDhj2SdzWlksg+bcF9Bvp
U/uHm97cvMLK/efG47TEwK6/HypJFOraBGM+ypUw6uKTL1+zCOdu6yTYsksDaUvLB2c1GaILYz9a
Uqr3/BFnJxY5sRvj6b4I+E0MCC9VRG3TVBpYp0RlVF8GhUJw25wv2/p61NzlMK3lEv9UI9L5uYNA
vaLrSu0KIMK1DYnCyiFk3wPUAU65uDit0JKEh4ZzVEiL8dWRv6LCer5dvHJ/duA4ub9jnC9azHYv
CcGp2pRvufJWzoyx7NZNKiAsDTui5NxPt7JJ83uyOfG7VpzR5ZwGKW8eOG/HchVF9TjeiznheGRN
ThVvQao810fi2Pn1MW14vMFaR6JxQlg0+CyaV/kJV5506lBhX+65lfM1fCcdorEPe8JDFPJv8x3I
P6Knou03I/6Q+CtBP9VbIppfFMdZSdiJjPXnWnSoptNUI1CLsaHncRNUvRwGHwZfHYND7QNDAmMp
jpj6Z9l3LZVlthzT+a+PK9HuGbCDKbOHjz9wWyui5XE90JyQ7Ay1x/4EaSHRjZ2ofvKBQrQ84xOz
zDvhP4Y4Uf+ilk7jDgxJg4CRDsWdTD4XOWnpzzHfmhUQk3QphCU38HaOD6W5ePc6AwSs0MtfCetX
sfZS6Z7Sg57ecIGCIQOXp3u2a9DgYtXlOWpLNdS8WY65R4PaXDFfXusJYRYSJLMMaLEHIRtmR2iw
jthyhpL+BNXzf2CdeCw4lqxgPsvHE3HyXSCGdheYx1NfkXxIAUDjbPWqHYwj36Pt70zgVsNZhm56
2B0fhBQaBeWnmHvqeR5KTR6V4snw76wAiHWBasC9VfWSvvSEQzTXpn9qJc7HYck2zc5LcyDwhnIe
YEX9L2y2EZcpkr4p+TxP7QZYju3Cnj3qfMbveHoEpWr5cDwlNJ+PPcMH45WS7dkqghzOngkZodrs
Z0bQFXMZTEJgDnfW+Zaoyou4TpemihTAAHntPH1UiUtyU1p3HK23scLDvbfWbfCWmSOdzVOa6xWM
BjDVkKHw8MLz6zxTJBfozjcxxsO3JyKQ7KltDxM4Tdv2szq9MX22KMjOOqcEO97R3wEs3Tma39Bx
5wzORzaMhkWUuczWegcgnRwnxJ04ANwcxVKjS74Ys0IAG40VieGRIxSslo3/BCHvn1PAjW6apsc3
74hb1v/zXDdS3KSSg7sxHN7yZcWRxC9kenZBSVSEZuvFiBDaDU+KQVr75w5/jeup42Cf3RNkxMM2
A20YPq3dV5WtHblIUe4D4MdkBHbVl4H3tpszeUtC3zJZSAMBUFb4RAqxnN87rKZK3hvsX6QY0WG4
nSEdeUlUeUamBML612CErq3+iiwaYETCgtt7wOKzwpzYIbyq6EPMT+aY3XwBahrU1MW/SHX3IJFd
Km9nuto1t3EQ6VUMS2hEQnbewdORqID88YEtadz7B8RrMBnoqrQHlo+zlDQNK6IabQDqSboGsMrh
LYIgy1PMw6mxe7vj979DrHTa1RD2DxULmwR4QGZYWemWPgEUf8x5/ZiD/ZSQehXElicjHX0ogN/v
zJsDd2TdTbGa+fY4wuqFnBikwjmoVLZQTQtrt0mIesp/2CamqdJVW+dN5vLKowujRRZkCbb5Jfpz
BnnOauHW2LHToFzpcpmviTx3kD/kXLn+8ntc9Pz9866FnJEdkW7MWAa29vyOZxERE4jbscAfox3C
p6nBPH6UIj3hXbZWdHzZeczSrQgw2QTe3fuF+r3JUn8OV6jSxW1Lm2gnyESzil0Hq0+pnPEZyQZQ
kMjvkDOQQRK6w/Mx41Ct3MCN7XUpkGomFA5ARI7PamZPBdCBaSrzF9bywObz195N6C2OgYVC4P++
TGy6f1RlPyBSAgRndL8QxCIK2eOGiA2gjeO/GkAu0Isl9v1XF8zKIQXrbbdisXRPBLmK1Z5zp9K9
NTDof/rt4Or8WEl1Tk+acX43x+kA8LvxaKYb+nD3e2nepemYZHeO3nrg01dN8xanyRYcyjZQo6XX
aMClEpbOdpH0nJ9kVwTemgzQDHfp+dqFBXJ3yTgAkx6m37cyFTygT7ZjCrp66IgGQkYK0ywX6oie
fxYg/9T7yjF61SueHR/I2zcYAQagwUypLyBSMecdFD+uKU006YUOA2DVDNL8oaY5gG/Urvalf3As
YxtwcNp1aYYUT57OM9805sShplLBtJ9Ap8ykEYBFIHSStlsfl5goyNbRnr2yW4x8owJkpm+28AEJ
QSEF1ZUB5XIq7IP703ofXecpzy1ZrPvgcqkWP48rLVTqvXB8usM9An2wbFwamGdlwu9IRjv452bS
LZV8CZP2OX70v7H/RuQ815Pq9FlPTRu/AfhwslzZSFJWghXhMbqzta5hDOBVmw4cjNisCB/CeAIO
VNMjzgHS5PrCvrn9Bg7OhS2EaeeXYzXjfP6putITY/m3phjUzHv3DSuApL2Cap3m5yBCOK2fiD0S
XSqP20rt260hKnafS8VaZp+YLMXDZVtzCwDPcKYA4P0rXLqo39aaTqBhuqHlBeSQMW0ceTs3RtUK
jNo6i7VLG5OwZDDiMBBOKTqlreHscrzTySFzuY3pQ2sMpfUjg3CrYUwrc9cbF9GtMmgkpsw8etNF
KjF13600P2iiGWy9g4CEiBh1bgYLv2l63zOA2QDIb0zKuFSey2gqxJBw7w6YzqmdpZj1yMvpEtT+
2qh44ky+6IcEFv0DaM0MrgYAP43veIFsqdFHkEqozU0gsDcC7v9yT/MVimiyYoZ+RjPhc0LKhAM7
KlylwevVq1yzhhv9wz9ta8T7HOLUZph3PRuww79Q11PQhP3FCnx9Ecss99aoDpZLCWmF9lqzx1Wd
xOBeINNdXyb1zZnnvFiirzpEkVoyKjJKHfcuYIpU9ord8dm4N+2/uBwo4prjo/vRTZtZC9Ew08DP
U2U5kqK53BPEQwFBBK7GSA85HPCWpa4/AgN0G2XDRtjOSXllqqIc62RP6b8hB6N1Xn7OILvddT0R
q/8uiMgyxj6iT+ETrKDv0ctRa6MYlgNp+0H1sz9WjL58uUOTO/dzrqlD/5gkctpbg6AuJ7NfJ0hU
2OxeISPQcxDqex+wKMJDP87ySNnO7FLNr0mL25keHxEa6HCg2N3r9gceolzi+97VtyLSxjIc4h5j
xJkqS9CqY4fjIsRR3f+8cQUq8+ZlOTUQxavxNde9oaSgRwOwoQlhlo8CHp4JvloUUC5HzP0/FvFz
ZeImnSvis0eR3E0rSJwH5D/0s1LDBaiEZiGeogph8AXhNpJC/ygu/W8W18CRM5qLJ5JZDbNtRBk0
wAdeYmg6slr+9JTZa95kftqUVUNd/+DXHuErhRviqKi2Obr9PI2wxH5uN1uzbyQyPPKZHMH5Ehvc
kxrS4Jsiik+Y/INIuM+dR3ees6GqeDsSDnYMQfGGDjXibC0d1U6WHv6Un8MiFcS/xO36Ftc1UPPQ
/AfLwfGcjjmQiHVctht7Zt6gGqQQa5zwODsFVwH6XIVthA/RFytRnXwRUSGMWHsK02HGCwvGbo23
+jzfg7xEuVIqsI8FAhJugGK/bJdcA/+G0OoLoviy6zOWJdmNZMK9os0qES20YdBZ4pShEoq1zIxz
dWauMbRMpZeK30sibSHICQX0k/5/lnChNKJBPLyNJRgq/8bGZRo+RDXhcDB6SS82thy7bCVhuxrY
2zl60izPkML7+lcXMiMMGV3j9ODhFmVlSxSBjjSZZYuYohWB/h2E2JJqVNiHErtWxVilIw9u0epw
S9NXZqALLK1cPAepzILvfS5Z2zuFblUPzsMLQGEVlMMg7GQ2W53AE1zGn375+A+IaXkA1b2IaXQ1
DCM5H+PBpySMVMNaOqvvl3Hfq5ZE0GultmSE+avjy9Wu6QPLWjIpgKKUWdaJgUSB5bQeLOp3eYoP
+GcrRCDA+z4rVcMk3Rqs4e3VPj1Ac0HI0vVRNniBKTGjDpJe52AMtSegcx7QO5xW4j2yAzIgj0xj
neiwTh0Q/m9TcD95JkgLo2mm3SzDMPsSkV7wgfZomCBKLKCFLhPKoWL2DLsfZ90No/PyYhFMszV+
MG/kA3PVpHjNW8pTpUxfok75BP3b4qocWp9uhLsDNWbS/RD8pb5ktJiTZaAAJPC6FpK/PMfT+vTq
nhWmY7SqluUTBZwXfNwVlwOEdDlfIdYD+v2+ptXFyY/ADl8USbZoAnAVHzAqD8bA/lbYznsCMsE1
+iHW7SgO2dSn7INVzl3jb/OMs2Zz00OyfLBv6fG9yKamypdKyxvKEWf4034QAYouSwoT5elBZcSn
Q2mENRtx9IrjvSAT2Mf27gkRdiwVPW6FX6Uy5V8D3CgtbM7vrPVkuqbWR/mZ9NWHtxZCqu/dHBQE
m6uFyiN/wiybFALjjnU+xKFcWTW6/Yqj/be8yvnDLJCqBZ9xYrtVWLVDHzJt3XHX3eDcBVp+ZZz9
XdKaa6Ve2gumsrGQFIAdZRP+PNlH5GmlogYDphlsE2D1B53ZNYfCZple3LJhXQvfmuPNG0Zn37kY
5aMrIqqf3JwmIJjtOb3HUtLSlZDiPGGTIFaVMJb35pNpmOv23eVbDHStG705JLkIl8jjnQLGnoLZ
kXCMj1nTHXerlNazAhKXssu+ZL5QsGNWvgd6Ft+ymxNlRtHfTW139Qak+jZstFk+MDRFNs+ehWel
1737UJvQnlR2pnJwW5wVfD/AvSH7SME6LKfMDwqfbjM2NokWB1aXItl1znVphGem44jjlxZX8fLM
K7h80aD6iPEMl447WkYs4DUPzlebyqZUp3UvC6rLR4KMrtjbGnVLBc2t7Dy486NmJuQ8xkteoLne
SsFaL1CYq+hjkdtxEIcat+X06eppz+8GuN3024EyMy6gdS0/0MnXeIBuuwEQ5eJTEmTlzVxnX+Dv
KmnSdvrJn+JH6fuCPlQ+17b2MaT6ecB6txNXWrBYOfzp0LOu0dSGc57/JgAERs/V3IOiGzX2RNXP
XHaO4X+/P36S7il03ZFD8eUj3DO3i3L+b6aNLCzxZSjNQdILjA6KUSxNelfHbQscWm1/xtx3lgwb
ALS+hNectPpAt4tWeT0x72urJt+gOq1KxnI1lhRfR9YpjlvSODWG23cVgaMQugMHOatUFvY3XeBZ
JNeO9smEkiXzhW8Gna6ueaRp2xnnt4ajc5fluV51YdikG/LupfjpD0sp4hvNlhA+RW98jFae/vVZ
Ct8RrCjxOtnkQCH0gWdHj1MVh3xhjfEV86cz2FqeD9ivNQYjnUtWPDqlf6zu4TbpOAKwuSzuqjnu
TWlEJpUWrs8CLrUlwd9ORtNH+aUMSSGific8SA2qBuDl/k4otCf2tckbdDqkg3jUKPCDf/Aq/gF0
m7fOvOIWQptyrQs2+xJ0a5le6TC3nKBjZqhpj8tj+geO1YSvZ13fO44aeJjEIEebrjGiLl7RpBDV
7HtN09NDnW4TP3ixMU+ClgawoJF4XZpx163JVQLmbJK2q3o1nyWCl9Lt3bJAMaDScODMSF59pr5z
fag8ZOcpO8KedXRbXZC9M4GMFOwmH8z4DH2vJBeldmYn3tryxRiY697lc3obZztfl7yKy7Z0YC1x
xRTBATB8QSQ29YtDiJqRuMhMTKIZugC+nS7s7AAufMAlTVV2xQTUoPy5qGfdiW9fwplkp35c0mB0
l4FfY62uSFgEkXqiIBgF34iHisa8N79ZsYl9NUoR6FkY+SfW3A32x0sQySBl+bVv0YYa9QQ3zGfP
+5VcM4pc7fiFk+fTm9B/ZOuZTVH3y1jJ4wuPWln0mruqzzIb03s7WxrC0q+ydFHirwLP0bxI348I
z9eLno8/anIjrO+QFVpf7r5vTavLHZGI0/RUfqSc9/GeGz9cJZPpOGwE10fAaDvuPxvmU4UoFfv7
2qXXjxZFtquRHZMaeatSSIyF9579x1elcYNumkyixqvnJQGir6z5NqrKBtvsKLHn8aQtY8zpFECi
7OSRtQ+vepGk1ujr3ILwpoGr8D2eV73KB5H1N5HeXqZRmxl397EV45DQAn6y8AyMF0ZV7d5tHmli
MOXYp+h5mqpvJOXvgPXrOE3DQLbe9WvJfoGnP4jWN4rChP+dyl3PdLsilnb/JIcYffzjeQX7fau1
OzL09jqvtIklFCAm//QloT5z+K2YOh8f+XJrUF2I1FlWk4fXHYcdPSpN+LG6TRSKOJycwiENodZg
TTd9WU/nDFkmnTrlvE9+U0GfXVWgVTjczHndKTPPGrnsOPOkk6w48bVVVKgWy6iI8ub8Vh8nh9GV
hsxrubonixi30bNRErZRhDamBDxEVadlshMa2OZnYMD87nggHSDcNsHK2hxnaJ0sx/3i5fMwSEkU
1lp7zQ9r/HIi4QWocAmZsTCjIeAeyZTWnNnQM0KgHh87E/axNsU/IDSt+umbOTCsdHKH+1QJ37Qo
Jcc8D3+f+0ZOBOBDwcV1qog/thN9IDBiXEqC0K+8y/w/sDD76VYxl7X2P3JFt4lCS1pBiUwp/Gsm
QqrSjtosSIpoKR74EJStImGu6rPz5DB+S4zbjc1Py4X13zOjiudONJPbeTRIsNbfSK4qv8jy5JQ+
r4dxuNTkWXlQegucK7aDuM7A0HMkPF7Mw2OXe8BJ5B7lBs3V+oC6WMErnOcSCvYtuOBmGo45FPiD
p4w/l9CKsY41wyIE3yKWht7oDjCdwTbzq6lk6mdUXavvcqnoYaIw7Dz+BZiE+UipezRUC/UTScwk
onQpdPe3ZDTVo8TXr2/oIkSuH4Nst2h7/TzqQrvG6q5t8FY1PzmuqURxdtBb3Y2Hc6IwSQqpqtFl
GM9o3NOYUI/AFPNQALQ1cKPjeoS1C+indyhHSd/W0HlEgwH9nwvWjzjw1cg/vzrnb2MNwJuQY4R4
6WrUf+aqgEQluZx2GbK1Lt1SbRPPK8uUz/nFVXiZzTJvforESOAtJSFNgXyNDDLYVhcg1hQkP8E7
BuJT8dbcrApWu51DOXNZ4bdIxR4J4QxhAQrD7RRCbXvio/cVDhrTz6Pw6Ejk6iPQBVH0zlTyzqvH
TBtBT10RKY4DsylhvLtwP6QYatHtFxTdFhhhP/XAbalx0OcCftJ4EwTpX3JKwR3e/YF+bmVocAKk
2COOPH3U9AIslw5dgzYqK/usu1D//MbCFQZLd2oQV8pyEPC+dU9kOdkSo51igf0hHli8IiyIc+2U
mzzokQMJffpOqwFt+DnESbdhwSIrju+utAGyenw5L3H5BNmQnwAQR3C9z+Q9SASrnsQbZlYDdLOb
cnZekRE+/N9bvXGWNX3BH6009KH1uLDRaDEmLYbJ0dmgfTYpZ+AwHRzCQjeiHMASm8Lt2F3F5aRA
urFKv6MCUP3PM8pK57enNA6V+ztvZe1D6aXHrKRKwC+mo9vfbBYxv1sojYva4JD8JJfxc0/toyEK
JzanNQaqML6SeIt49xrL64W7LBa2EK5cPK0OuVWWZ+GBJEj35RnlEuacpkOp5QRQ1lkNyD39pr88
vDCsvcBMT77/rkcB3yBHsgSceONbjRMIHigGf/JfOsg2LA5DZEMWzOEJ8FicxGKbbTBbQUAvLqQQ
EPjz9KlXuCPPqLu9ZT74+5RT4WE/REAMR5f/4L+aWiOe3l2k4iXQDLTjrdBB+4dM32vLK3H+T12v
eRIVVjW4flMa3PTEIRhHMFuLWTT4/BwLBG2an2OGmUNOe4yTrDp2rR3FeowK2M8/g5zOcVlVg8d/
R6xs1XOsGAdbHDxyvaVCHNGl+UOFGMZ2/AqyX6ULAEJawop6/jv92oUnRXzeul4mXnIN9UgEbE5+
hTOwXzm8NEUqMceLdautrpRDRWP8q5X81gbZ98xs5Ll3xkVg7X+6GikhwaqwpJ+t2P7XuixKsbzf
YkCA2NQGCiOlVrwEycplhko9tmLkASLeW8nYDaXEPIPkBmSRnXQ6q3LtkMaU27u/Y/v7/03zvETK
E1ePCXVhJy0/mJTXVGzzm3TaGFmrHPjX1b8IDJfHkkzoKw2MBfvTgvvs+KP/HyRmGPflg2SuP+Pu
7j/IECM3lFAEx+xr1CMUIFgBC4dXV40teO46oOEZexao6id1bVpxoI/sydXki7cW5nwJ31r78Mps
W8TcVccYeeHZmnZu2Jh/EQV0fqIvkWAWUJXJx03nphqBoUV3GZv+1eVldsT+TxSFauqGQBHyiQ2x
1E7tjQ8RXhQgcqex8tK5KdS/3ngHxl7boaUlcZZCV6Fna64B0NASbosl9bpH0vHdmJXGAHVVhoB+
94l96PVf5zgJGGEgO3TQXK+Xvqej21r5IWrSgh6c09+ZSwVC1zZlZp761NM12ZA4nr88IwDHWOm1
bQ4eRC0jGFWyP8ef7C/jEcF2zG06SfYAAiLPjyZGLrZKuukPSLi/zOm9EoZf6qCEigjHHfC5R9Dm
HQxBeZ0PBRCUzgtQS51xyaM7TLD/4yrwmurMqfEnvqUVyfpSOTXy/zlKcxvJZmttL/oEuGTxzdNp
m5TOHMuDzHwMWrQGEjuBrju0I+6fAlH7A1EPI8KP80EknqmUHvZ7+X9HvpYvJeNrcs180UT+/0im
uzyPhGUIggjAjzj92nU6dzEs7i1QvbQ0Yb0CQFDmNJiMf7wXEE6SsUArUR7VoBjZrtESD3Up1/Qb
YMfnJVepTPQAUz5c/qgWbxzq4j9VIomcpkjADBtm9WijiCNsxb5HkJHEAf+X/XGUHMz2LJ9mIVsG
oNqqeT32Dgl6ZDwUzFyKiAcaDuHm20+j/D4YBH6BuNUSKs/Y1rqyGlEpAh8cz2mF7OBSXOp4x3y/
45/PDsSxYSij4b1ayP6k5EkIo7UVgkYzI7hYTq8xK9NP03zFJpfmIs1c3HljMgTvg+Shv5xIyhGa
4nu0rG24L67u26UUAkmgecef0gyRZurcLq9aER0hUkj9q/qsSn5Nm04oluCnrd7BsCUaUaNX7huo
vQm5KUdmWFjcwmk28dxTXQGbt6TmgkO0rS9O5Q2Gp4qwdQEyB+MOKU6lPmvZreLHIRnZaTLwUQPI
6OLuJQw4b5RkUsMcWn9SjTgeN8NBGC4UV4oDrkc3AarLS5v9EnYJAEwb63xL+W+zllZBXY6suQTT
65NIjgyBD/4ScLTHzx35UEyCiBPz9DayoWNrdpprjH4XiSCjzA2BPsEIFsQqhvCp1N0anmX1T2NB
LJkwMoRvUjZmd0g5bN2Hc1TZuVLfsax/PS0M3qsVoFI2pyAoC6aEZfeo0jzM6Ezzas5soIcda3PS
4uQtqi46LDqWOTHg4hqwHDE0i0vL93SOPY9NKMB1J6r1/fQy1a0f87SbfrVNfSBcseHbJ/zuBauu
6mQyhKiHkhjEnY9So/CwJdJuF9bjfFv/LdJHWir3g32F8AKURu9vODGlNM3h7tuNkknIIMm6Uzkw
vX/mHlMkY6Lqgxvw8OykOjaQLfS2kGSbu1f8BGBo50Jg8fC8yHqBkbI95hn2UDCrkletI3jEB16u
dmeU2bD5TEs2+B5ljDAS0dYYVZoICZbDAY2LHBk92Rh71eqTgPXkDMqrH6fqeEbDJLK3U4J2CjkM
NIIn2KBHYI8opUGAL8/lUZFCK+JhVVZKuFYSr9leAecN8tt5q1xf2QVBIMrQ8GIA/ke1/zu+geWi
3A6rDQ60r8iB/j4bcQKELrgx/IcS36EnrdNrxKLKNRyaOODfoulwMZsVOcaJ9q5QEDMOsow9kKme
F2FwLHicWikZgD15cbw5xs3ceUniC8RAaP9UJJqwLSj9rOx3jiaZ6W0Dx2xsNLcLyU1hnCnqVUbA
xoh3+/NvfL+cjFv37/3VIy2a2pE4gkuyuWmPOU7iw59mdgbrzrb0RRUMS+56z/gDRfp8lrPwj/2Y
xkX0NDUdlNOh9VuKHzZfbwzzptp+oM5yKG8lEzCvv0YnTTyuhU4R+1eoPKxBc5U3eUSJUN5Xkww5
0B9uFTOOVoQvdxxphbZ53CN4uwqaHpqIit4cd7kA+Gw3ZHudtr4L1H684LNujsmR2/cOpYpGr1vs
wITLBGcco9EF2yF6pG/jLCMx7ndJHY4iOC3ge4DJ7NBs6yh0jqPa2ZtjasGoJrC8J/5oJwpmnmgZ
Bv9lmT35lzSXPsnP+dECeF4Skr+k6FxF8isQrF6isC+VXQnSQ8vA/h6C/jtE8B62lvj5pmpR1lhZ
/Bmghx8eVUuWkHjZDyKiFOFhtMaVWs0qmKmyMtmL7/NY2JQ2KtaKdrRE1V1s/5wUaJr5v0a0J/+4
x0DdTYSadY2OdEKcyyU8oioGVVhw1erWcDBuP+dfMQJhFFUTRMpTJXw5iVvNvrNr/7kyfjynp1jb
ChhJmeZLpzj7M6qrWuJqf8zAEUHuszD7nICyVD1tppkLoptp2cd1EF+KQnPJStrq7ZWVB/LcldYG
uD7NuDxaNPWI1fPNv2CEMwfD0NYiJ+lk4dJe1Aij1Syd8+Dez61LqQigkO+nM2gb01kW7TZrSOFu
4HEYiGDNcJ+DhLmCHI+IBVPtTPZWeCIA/E3ooh8h3E1NK/Y1i2/uL3ijW8iBexEpt21+04EsFvjt
ibyKCgSlmn8ER66YBGC1ff9bwhFVuj8aWKUDFHF8S/m6XxrS+Sw10Ij3oG8hKbGHT2MQTaNumomm
HYXQyxcD5oH4FtbhnJoG4ho3LtbPaO579asebZobeE0PCQotzZ4KLm1tP5951tTkM2NZ2TYgdXvb
qZki2eUJkx9v/FS3woRw6Quk5MVFw5G46zVtFc5CqVCK0GQu5sVDu+tYrW+gWCxKt0sCEE67sYw/
isZi6dTDQAH8Qeb2aDwXKZ3MC4X7wl0kbMLSi2ZixGCtYqVHZwP3GZxCsQGRdNCYwrU4JqjE5qkb
H8fu2ch1KWiFuU7P0l37Zyrbh4E/tr/8j121rqCNFAQIoM8BVLHdb2CZ4oUudH+ckuTpBZAQmhPi
fwoUAtsYMue1WFHug9Zop6XFzDl/C0ov0tllguaasVJbSt8WgZ+K4wGH1Kwxqxh0z4Tq7+z6tPTI
OMSwh2ZJF3FixxAdwFQ52CxOVPfz7pfIJIHo++epZOa+RLCqhhK43y84U3oiOPFZJ/nPoYIuWjEl
mL81+yyGCUHi1ZwT7kqLg/FL7r6zRfkUWDOP5dHBaSPH80FeXQFJ3wiqBKn2MOVW5fAjOrNQweXS
V7fhSBJOJPcO6xHIca1O7KCUQC1/Vy/m7MlfhgrxQvYPTQ3ymLOFNDzvupMUtVHYwNr3tD0iVPJz
IcY+WUyfrM0B1Ug6+yDC1HWLCYudfbH/30jcg/tbx31QgFM39+S/KJODy+iHHPgnCRYckyOXoiNq
b0Pddr8lTi+vhvLw8E0U3Y0VtevKuzeiH/8mE55yXP9bPpnri2ys0VkV3DKPseRb2QZfjJVIKsEJ
eq1Bq93AXX0X2An663RGCHdRotaB8acpxDqAIiL/i4M+dfVW7tqSOCw8Zw0VGQlAalJv0nVtRz7S
O8wv2VVKX7YuvI3c+lMqfp6IUahRWthIe3wuipFb8pmSP+to6lF93E5FKT/vrpdvUZ0vTyIHUX3T
4DFDyqoj7CDViuICH7xRtg//cSBmlUkI5cNhXN0UfnWVjn6uV4nXrXF8K7cXbuO9YDJqHkpChFqJ
YhO6K1L3EYKXuDdwmVlZ7sspV1dBTGf0DJxnRWYYM5GKVBydYjwVSc7Ci2todVSZxQ+aNGPNGUrJ
fZx8f6qYpaS3Y9Xy4/xg07xD4UXbjCRkbBO1m/h4GWmSuF5fNx7LsU/c3+R2TXQBumJp3P0w5R2T
raDopNmzmxLsIHygjfhwjkgL2XPEn76mjhh9q5VRg+dEkP+mA7gupXGTRER9p5vC+DXIzSqXG4IW
6dTBVu7MzI23MTaPSUx4D+JNDutjDTB6HsmFZLoF9l59W+tVTWglz/fs+x+jBAnnfhYfLotmRvCA
wSRJhkW3Ap47O6RAADVdfv8y5Cu13a/rWa4BPWsGbZAoLH9/WgbtwJtf71Q2TfWXYEE5k2XQezm+
XzQJp+OgItR4lyCS+GfUhEHsKi78j4sppMjV1xCcSURj+pAjq2vcCa6qtOyUgzwGCFTn7KRBFq96
Na7MuhSlxtKETouCNrgMDYhZx51Rf+fz6azfJnbwG0E/QYng5ipGPuUrvxnpd7hbiBs5gq5qZsOl
WcRY4VHdR3/SDAA6JjBSPc0C0MZWChNXe2iWBKy/QJ4Ncn3fBUSwON1baJKNfopmU4Wjsnt7FJoO
AWTqGKVaswOXzFKpTmMlNTMaS3FwONJFWUyHPVxUjMhjomnzQfxMCUDFf0KQtKfVgU4yEzzcqQkL
YMOeqMrSPMwGLsggUllifZkv1qUpK3BJ/6sr6+HK2bw/qq2JOmwfNQmOGUUloXdnCS0dSaE4nZ/b
QhxICirmtLTbJ305AtF61EQ6UFr5wvB5cM8ghY3K6jl9t4dB2kDfM/OplGhU0SYRnwW+/XoYANIb
o99D+dBQXKSpU0OP0072Kyz80NEdfa6LTANWiHk6Ud/EYdJCyCKQ03B1vrv563riILr+gR6iScN4
q+VhlZ0mzlR8v81OqSuMswiWlu7AhASAmOHUlssf9eZ0xXynmIV3eFMHPL7y6BuYoK4XAo0tlTD6
tLLF5JdPpp4YBS4Wx7S4Q2BsxznN9ZaNKbqpdG78TNavZixpP/nbkmNJdNJUxci+8ZwSl1gf5t6S
lT3Fjdtnu/PsyOAZbP8+V6hwepqD7l9fHe+DISLLF4Yu91bEhk9Rq5CGrc4CELyYGOEVw8w73IyL
wnvigElU7uX5YxtuG2nYodwuYRBhnqlrq/NpM7SXilPSjaeaLSrq+mtAaHMJVbLppsgwCqrMZ+NU
JTAGEqho8Q8VE5lU/TWorve9ZseAKWyQepz+X/RbkqF5+Y/M3VZIzOPz26wT3EhI1ie59wTJ0jIr
0cRk7+ENKFnhV7aHw+WnMa8HzU9QpBmHjn++T4AwNpBWybwmhSTgZDH3qyeQqmAfpYGdL6GBPFTb
gXAS65zHU6EGlliClGOg4MzUrqWif6O3HmC2RgYAJsSSsWn1/OHW6z+6poJT3WOchyB2OLvBF++C
6aWkpnr6X2ZuSDJP+uTzGzeVpzSmsYJTSL9HLWcOf1SsizXYHCJ3rN6mI9KanDTV14mQMDUDlkhz
92kpYZEuJ1gZmTP1JbkJqfdMIKMUabowKU1zQ/JztjzGLGma1SNS/VbUw1l+m36fC2a0bQJDlQ2P
ar6FA8jegWY06x2LH/WhoWfOFqdDI/C3WvN2wM6Cz3snQM7sm+wxoLFEjhsoWiB4RZICxHAYTf6w
VxOuWAX7emxlbJKYByE3bmU+kwEdEt2KK0rWt3YrtwSTzJm1LQCQHeNoqqyQdcZVjJAYQnAXaO9F
R0alPNMjek3n9AOnn1mJY5JGONqJlNymq8/bIWWMxJXTT05uZtwCyJepr4XctqblXZGsFwtzbwUb
3NlG8DNtwBD5A5oLqndLz+LyXAETdAo+yg97J9CD99/AO6m4JaRpAp8PG5MfdQCfnt0Izq19tclS
ThmdPbJ5lsN2fsDVV6E7JQxj7YB+Ha5EkoR9f6N9020jynibVmn14zja/pEv5p3pOYIXK7pxQ3xU
Rx7Gj3Zp04ADhiUTI7UtEU2MxRTOVB0ahhrVgZ3nHvrq8G07wiu2JFVcRMlqQa9H6XA2gBGSkFS6
lxMLDz3MnhK3a6yxNJBBOWXS9s+X7+/O4S2uQuZkyWjthyXx8mnTjmXpADW8OSigm3ViwHldwNv0
RjS3oKY2oA34GFcvb50p8VGnpgB6AKtkDwemeWuCjrLkPyDG2xJK02eNfkqvk9+935aYH5IA5141
ASWddi3Ng3G5lPFdsDnppVCS6AtTtIUk82XqrTXh3V795tNNB6q4w7knre+I49hf/s16Hc0c91lt
b2EnOgorIt1iMVc5//zgFheFt9g8VEfAt+q7Nyi98lFeLUFJL+NhR7MQFHwlxOmMnFZ8hC+uwowG
sUrlj6ZdiHEf+ULf7brxn8Pykd51f1mEpWoC311kvW/uH0hEbb4slb46VIepImkSLEhsIz4A2asV
cGZljkfGxBMFKEwY/sSjpsMDOiWZKZHPb6qBj5WjDj2m/TY+HnNxvXcJN4FuDiReb3ppL0knGX3n
phNQ5bQy9OIIdkFRHZdGaB7ihk4rPxGgDobNeTwVC3FFRm2XbClo8ivB428TMdQEl91fRaYWg8z3
gTJdIU7NF1z+Dq1b+YKWIEVhFCuH0fojr7xxLuWE315cws0HTKL9ekAZEMsddo25VZWh08BiUH0q
ju3aezLjucynXdRYPSU7MmEWYp2+f7TH8Mlt2V/qTVLFf6jjy8ty6bPbn7y8JTWmOOxQqnlt4Qzg
JgYnuRw+p03bxwBgLtJvKzoCt7TfRum/phzPUv460U/nHq5UyNuqJa2j7sO/wAgMKOFzk6JGAMvo
6w8kUhkn+kjNRqR/kbNwg7AFTpETkxHq6rg9sHuQD3lPqjyKRjz9WX+Bcu+MQ8WZBnwAwbwgCPo0
wQCOKgSA851lUAUQR5HhYYeLuelIypN4Umiy1/BjN3m0j6fkXaMWbmyQ4i5WuaRYJeH13LEGmMff
k/f2GBjyKvoNGMu6Ow/RxDirtauwmROEzCDK6PArMDL76CUX7zgespftLRdlG7fExKQ9U659V0Rp
Tb611JIsXelFV9rZOhBK2rXSFL0kL+QQ88Xbd16fVCjR07X89KldMCbbErQkEFizVs86dZB040NY
4phQ5rOrH7lk0Ij6jt2NWV8VxaZpY+Hr4t2r0xA13knEabIpZIcXESyNb/g/OcgDopp65LEOXmdU
txL7+feAd+55pI+9GaLg2vmp940b1gQ5gSCQ+H6T7Vip6nENcUgF6JKygezUHkBnd2qcFij0XRKZ
AbZ11igaoT7evpy0D80gyotDubXCpPavKA1w+O7Wzt1wTOY11aaon/53E+MOMhb+LgFN30SSjX1J
YsihJz0IYRc2z/RDWcCJF34q4IONjCKz+oajvwHMyr7zkYGzmc9wcVz7Nx5z7s+UHi8qVkgcggpU
GLxNGhyCVARyKuwLD55ow8Q69z7TZKTV2T9ZnB6rAr5uyPR5Q/30mIInNokb94uoUD1hehKdMxeD
OnsU8syCL6D5sQGiGJptcP+b/0jQwU8IWb9IOpmy3i5TwAcmPr8lFWwoGe831OuyvHLpnE6jiSHv
hIO49eWl2OhNRs10aiMQMcK0C6dd0jwEab+9NRTARfuUeRvpSwcaMi8wM9cqfiy43q1NPxlFVhdL
FyT+AysvT+rH/uzrhNJmYcaqgs/3k4R6DLDGZjGRnKiWEYOgZqQ1sRt39f+uk7XJeHa247fjVXZe
FkpuBG50grH0o5BTTr+juU/Tp2QLVvjjxgjO6Ry1nQ8ewwNEoc2Ec7Y/iBTEGAeFoUKP21Dzuu7/
SSrLhlf43/tMAEogova3Qusv0XJyeix5mdBcfqQx0qFh+muGLcp4ui3yDa622lnI3RfNNbvjM8au
egt5l02iBbiYAbQQC2xH9jgB+c9JFrHTWb/HailrqwrQnvEzfvlE9Dj3waqOeFRCyNvRowI3fHPl
ZwpfWwEmK7rEKUQHnRGzNmaJ2z6yjKByLTGrIff92n/Nwy5MUabJ2SoIH1k8ZPv0928WfJ+VvpNk
nek6GJTd4q6i1DPQi9vxNs+pRX733G0IQUMT/x82R4YJpIOixfy0639fpGgBpmhyW/7TRV5nR0RV
WFMHRnHLTWh0NPID5iRCAsMmu9Mcve+WA1ZIstAjMrCIrVyIhpiZznntmLKXNKDhicH3feBOdy3M
JT9J1+xSc78T923VgY+xqBEG/3JoNVlKUWbx4FlOImzPUM9XOQrUqykGTyA/Ssca1gC0zPEN0Utb
He4tK30ED04VJOpkqXyGSw6eOyyWuyPdjbn0FBCb5LHBw1nPbLa8xvfNgIx9+db2qOG/5Z+uDEeO
1gLQWWOPCZE7pasRax75c+zEsh6BU2+kIKDcNiwvriRr1xgGxCF4i5HOK2QF2H+2JPBKlo4v5VjT
tVYT/qFzn3wwRWRyUqtXyu/bsrQJQAXfCVgd/YSBbl1KuoPzepwHABd8VqRQX1KZkHWUzmFv/T04
Z8igP2xJDGd5UjrxFZroLeskhm9cVh3TIhMvdLMnbb6jYmS44w+RNzFs40pGVBrc3Tdm+xNPwN5V
0g0gQGEJrY04z3HijFO1btePYzgcWs/0/SAiU/guPNRbVSBsg79lq9sKe03uc+fRokDF6/BQBHAR
8gnwDOdUyaXWAhF9na5pWmt0z6UwEqlMyTrycWa3TU4+aY6x8hLpybauGI4mMCGURJgMB0rHE2GC
yntjW/G/myIKiFL2xT4ZMxLq319rvP4UYqSLrnMfcrmk6vI5i++0N6LPF5mTfLvYXGFijCODDlhi
xlT0VBq0gWUImdA0HeH4HF5SfaJi4qgUzFtwV4e3RSunKOKmGvcOu4DLCSrlGm/YbwduoozYUXkr
MLWz3tIF5c4b6fzSD2/A+i3tpwcw7cBtenqEkei5zyKBzqcmu9VAiIdTNSXEBVM1KF/jVB6mEdd4
eYKIJNMb3Rze/89qu9n/e5Rf6lcuPpMNvwxrKTJ3AEEE5NUh/rebGaCadhJQBdNAcrFCuQgaEV09
EjIio0M9o2iqNQ1cAwyo5NBzqe1HEChiURq8N6Ht4qUFxptGsVgh4iZ2eBqfBljk7T+kUn8wPoMk
R2jeCvrtdpeMAWiW8buuy+0dsWv+ZJL11PaUmF08hK8v3r0rs9omkbXRxUoQoZiNUc6K3V6QtrX6
48381uyYcRPbk5d7W7DwUFwnIm6nlGkIRa5Z3TMIksYyPjgDDWvO9SvkJwzGZQX3CQsHc+F1bzpn
sKSPoapbmVJZZaXzqW7cA4n71ds8xS6ZtqDaWZ3AblQDLx1tFcQao0xzLP4nVMHBOW+U1pf4dEfb
MtfL6AAtbMXvax2yce0TmQxoLGYhY3Hi+Rqsn6UN9e5xvNOjw//3wxZZgow8z7ryNEiADwfp/D98
Tr/ApnOh9+8ch8VdwlLvNYY8tbhsuKR6aeTWoUGUQYYhokm/fVEDvlyiadHUf8f52jKf7B0FL48h
rXtzosqD1lF7IMj0Lgf4+JhlkrIZ+X/bHyHVJR5tXjSRdPJF3q61CXskOg8qNq24NOJBc6X5bqmx
LMazsCIUfjB8dnhMNLPLy2iwK8893O3I14ALLo3UzQjYXfg02gyIcThpg1wjp4Dv4WpZuQsaiD8F
k0Mj+4wHvHMhKvR65iGHfJkzI5qiNnoIj3QYB1sc/Sr9f32UtJ/ol2iMoEc/DwvKDMMzEwXCLho1
U9hUaVcDoMGo03EhIMTo6xxanBElHI99OzomMkfDgbqcvgk2PGhGjk2Z4qaQLFtZgX5IL0iVoT5F
kN36HLxHqD6xfBY/R/Z+t1/OSLZ4nyQj2mb1SQBWYaqGksLxVvmh1QAFO3oQBTLNTfqBxB2OuPh2
H18gGIXGIY8ov904av5Z+Hf+QVRoj29blrXiTPkZlZuxOx12pBaNE4sRE89OabiNeGRFVqL+ucpZ
u3RC7ozvFKwmam+8usOmF7OEgcOFsEOjvO0FG+cASQoAIf7zCPlkdKyeSEF+EWB/8Z8K0UvlYyaf
PkPf9dkAKxsxBYe2X9XE93Qjl590hfMhu7L0rO0OJ9ITT4c28kxH3TRIQiHc8/X5tMGLldw1w2CF
pu1sQp1s8mFTsxK7xloSavfT8Jv0udzwwRniscv4QW+dOOg1G4pvbWR7kb4iZYaw6PNAQ5gLJqAZ
1tw9eAZF9YxSJkHapwb+oILNbek1LdYHQM6tKazqQv8HYaTiyNcU+G5FxqQV+Xkm2RDMdlxRXmhq
POvigANYzqqsDLLTKdBTx+DRTxQUqnqWj2sgmzeWWf/Mcpq9YUgMPWu1O4go98HZASGDTVNNlOmO
kcForbSKx8NzWvMo9aF6qHIjJxtkM10/yhYQ23jpxQwtsqo2poYlThobPLlJ01/E+GnW7eVYghV+
mUhgE0t0To7WtLhN5BPFlcuqDeZBY8rMcwIYsWAZX7pNLxOw7HiWbVd3frGeZ7v3GseD8cR035ZA
NoxPvXCu2kD1eyKmix0R+ya15o+zs005D1JQf673+p/aTD6uu2etXtC/hjxGLtdgyss1Kj08lMhz
sQICkSItI6BtqtP/Hiwg8QODswL8jetLw8NLwAUgXBHUWstPGdWH1MyQOA76gAb62dZbTS45Aguo
C5U/h4bHi+6rr4hHeKWjQfGPqJk+cIZ3y/U440dAqus77Z0IhR5X1Lopve4gSrfyXIY09FN4wzsC
p9aw/z4VbD8G2dF7uVHOweCSI+iNUn+cpzjFxAggM11B0K3E8ljqx5rNd3PDI2H3l9zDCUpIww7u
HnEcC+rPEvNWvC9+sJe9voscJXKECt2pfiMwf3JS79aNh/pPkU/E1yOluOv+FUn05pPRx7Zd6snM
4O//NYy1vp5ImaObVH6dAEFT3ceHRZKDztntVEBonMAm2l4GkhWkNYwXooHBl+OhoiMjXxczx/ez
7UzUWH4ZeZhHzxQNSsiPMoGZjubkft0YUprc+JFwfhaTvgtCW4HcPljNh3hoalj2+z983SV/Rb3v
779a5iUtbJboNNHrZQqHdIeCZreYjcWmJ/+mlkIKj0e2K56DCNFTB07RxHpd+HihsvivYUO7fSJu
lE1APNR3zHgWtDwnOpY4vbEqb7STsVFC+Gxt0dKCB0AAwaZ5c9+bp1vJF6MFanl3wZOXZ5+yEoF9
nkEEWnBQZg59/UQdqbMglIBvRcst5FOcW6tLraZTYprSbpmzulueQ9Iwznm1ysFfF/9fZjNyIf4y
0oYULsxv7jgT/bstLvpyVS87Qs8xhq3fDQktZ5I3pUXmWkXn5moOzaF0xh5DZxDwymqhDm8Nj8lQ
wfMr54wJ18XrhCaZRKXS4eZ4rgDiH4HI5BRE3R9YEx5Cw85E5aYQXeYhssiwrGUin3RBUL1yOZ/P
K8KUtzc+lR0Ca0rK4hJGugAvzlFeMLc0b+IMzofhJW18zqTZZ0EaSxfXQBEyX+Mp58MKn1Pn6et1
+WP4slEv4Ou5eien86heQ407q41GfDgbvt9XpFbEonzDAu5wXtUKdfz63lV5/rsOxt7k0mzkO1S2
cN277pR21Amz4FSG1QvZgj9jS3cowWxbxvopgyoDFIAxESp7HMMQIZIon3ks8Akz1riUQWZ3Jwm5
wwwl/sZH5txOZq2a4bbne+br7b45lK7I/LZKaadpJ6xA5992pd4LyrNKceYn+A7gD/p5Oo3swN3X
frjZa4IAPq6hb7rKxSins8M+uODeCOkK/ZWm51rCBKJ3oLWpjx5ngr1g5FumK3fn7PusKM9JJNpk
QEiSAcWFxx4U/fOLnVQVh/G/BwaNBF/nRimYrgynfu/VP6lqxATuqTjuaLWSrgfN2aHwVyDCzhrS
jinZJy4IbOCSzzplwxxXXo1XfoFy7wJFpenuUU9PcsQqe3MdasfABh7YgQWE5GzMAN8821y6zexq
mGrDnHqPGor/Pf2yyABWjnkYSgwao3vbaH3NjqSfJwTo3wp0brzdxi7zsZ5d7aKIuvgo+087bUDZ
4cakXssV/s3JffK0HREtR/HRV9gZjez7arzYOZuvLSoxgaXsPpq27goGOSJZoWvfIRKdpR5mAMnO
RU7hrJEJZx3gehoVLZjuEHUMrQCKJ50Ktvb5t7UI6Bg7GpFBdaI+Cwl3mpvRNZ0RV/vaBQNDNfQQ
m4XUEbqCpay54ntqapmpGVsdUSKSmCYLvvp5yyDRhsyWx0L5N6GOP6v57vWrKGvETLyFDsXnLFJ2
NHzmLRLMNm73NogEyurSdMui2uXGw93bsep6zVY4xPLAjAZgBBxtT6N1/C7/xJgUbJTngzPBHVXn
28xPomefTeKx+0yEdayFRE5ITF6buAGkBDnA28kIgRnBBpxEnjdxlXesiK99KY/54snFc25DR1P5
oy5h+zeja9aVUJCL0nXb8qplV/YY/yfvFNNrGyMH+Pk6M8DYawXfLbzD9KPmrCHAtDIkiOX/QCly
JI/TNSUC22+G66ZTVbmgcagfuFW3AKDf/WreIxWJzVA7rWqMKKS6Nw9mJZx8at/TL7rQSdKiATx4
2SRsCDP+xCUW/WPG89pWHpzgX3WI0W11pf2cbQseuZjTF1a4+vEOqtvWUWSNDZG5lA1MnA+8jPua
7Mt5k12ulDSJbKuLyRrODeKZjC1nZj7XhgTvRmEWeSQZ7uSDTHIFZt3t6NthrZxZu7mlLMroTpga
TMMd/ZlNaow0wyREEYHgSMVr47jX/D1aDTb0meSXobamTS6sqEdEgq3uiSWE/FNpL2e5hB2Iin4J
/xaRwVvg2mdoWoKlvb/Y7hYo8vRtweMH4lAcURX+nJHMyrEWARbPonwZrZvtWysB9fPdGlUGh0xs
exnSd4dPaQJxtbxeEFwE+SYQxyGMYSFaqJUSTQeKCKzwmbIP+BwKO1/nmF46dnHZtELECjqEHrVB
WJv/vO52OKsAjbqmY6ZLoEFdO2/Nck2N5e9YBkszh+NtXs5cLBW+6gFUFJNk7C4ChChp7OX/gFBz
ZqaGcwdkLlIpLmO89tA8h/nvqg3YVQE4czXGoeNr16A0ZHe/c9H1C3oLYXazUtgGf4Y3o38fP3Mk
IbkZ+00qT1gDAw/hkbvfJFj1H6KJCHjhO4ef9kyQJt5JUS7nA8QlIyGRYLTrhRY4TIgelWgCSiun
bQOlncy2GeKbSAvGX/BV3YpvKWnPRlt8QnwA4mbg+r4UU8s3tj66Too3ugd7EVlrABgyk5Mx80Kh
2bOgLWWDFSRgtT+Za32IIDPOaPhfpjvS2oLzkCwS2RBJR5ZM2IbYEKoqfRlkLzxzys/BEgiIuRSA
dVL1D+NHEnNSf0MhrynLe1ZfnApyE1/QEqtYJRx6KKWw8zwHzDqLrmNIhft8MHHfVn2tAmkmb1to
pEf104V2D6k+0xo+FMliwnjvvqy91wyI9iXvW5Ti9AS2+FSMAbrWpZHXuF43y5lFVpxbRlwydI3/
e/A7WtliZEUp/QmqbRMSpjHJ45G6IrvffcCsheFGYd4zknuOp6WBu0NJsa87r3ruwHHAMJHnJPot
j2YvWv0DGSXgiWJL+8tbII/Vmu9x1WTSfndJIK75Xn2f1vb4wBaQ9ILmAf+LlbCYnYQn8v62YXQp
MKGnGFsyA2kVahN86M5Kz3UmwLBe0e8gzP3chVEvtw9OBG341qiYqne8e7sgjriZ+iwypQa+LlLE
LCKI461J/g4PWD3U+UHkgaXQYVGHUWnlvJT8Rj6s/cxy2eSgilJg9hyJg5Mx0Ig3M+q+qUuTEn1Y
dOM/U7MzICq635K4Q+JZ1XhjEc/z/IeoXTNZ8NgS0PeB7F0LoJEzGxsf/77C2T8J27J0lXRygYO2
hXnE90oyPXhsPubDerWu6j2AO65SsYnC0pr0hlX9C9wgRzRte3jTnPOXV59wzyKDAQ9IC0pvRTbp
95FHOO7wsX1IU0vvudbmYOYyAgnbUFBWbhSQdggPJo0sF0lOVwoICcE0itJZb+Do6TksCUesDkAI
BV85zO2iRf8HBlskDW5GBVQk80EsHuKFAuQPuWPglBjr+C1PGDvm/ofBBfTN8PO70X3sYyxskRLW
Oz6v5Itn8pN8eAqw++NxTRZ89b1VRLhFBllFREjQbpTI/LJ1DVMwBI3Gih60cn/UOgPvMgxoek+0
GyY4tnQFMLJF7kX43KS4UKj3mprPdWYrQ0nGWr5JEqdqQV+UP7RMhhhfCjs34eDOUAE6/edOo74G
kDs9XRLY131heXqDyAKonAuvwxrHnAWPGDLcqbZ+q5Xqiw9L3+QOgk/tQBWQyf8YNE5AzL3u796/
bm5G0X5Y6J08t+YSnd65/ZMAqRi7kz/c5hln1r5eWfqcy4MXKUHnIQA9RQYG9Oo5o2W5XGutQr7S
omMCfWtBERoOGaZ37GacT000eWo3aH9H4Dnh48joZ7jZJ2zjqTichW7tc9AnprR7uR3tEq4tPdwE
oz+vlsnFSIDHb0UrP+8qM4R6uvfRHDENQEQDo5V/BFxKtZ2F94J7kxAN51MJdfm+n5/3KU47yd6S
UXwoRhqCAW6x/eoFAGfyCh4NehaDmpfHtuzIQls9hPOzCPAiBh4cvdL6OvHrrz8eSlZvrDAHtYqm
hGasEpaMwGO9WaamHNmsWpmrWBVRVyx0t67gJBz5tzpvF0Cag73Y2Vj/JgqGbNIRCK44FsiOEtEV
PmRNDEFAAK6gvUVVqWEGzWT94JRFkWzDWyVM/SUnV6Mtvh1Zlt3S4AjzaBF9Grd3ZwPd2l2x/fxw
66Gkg5umD494sZJD4kk4HqswFgQ8bFeLmgy+C+0qUGlpWWEU452KdqM2NBdH8a/3SPZQCPtCZknE
9nvANm2tm0MUk9Kuzx/TCKG5ghg6wU6ZdzGVG/NZYrmC0YZvgFrXK4Lnj9b8+0SSEhu3/6pUy439
Vh6cHN1v3IkGYYeBKM7yr6kK3SajlcL4Eh0JiT9UWRMEf9URWWMEfF12+b6L+bl0IT01NxCdcNOH
QCBEWsFT05cRhRDci69aynBB24fN7YlgPH9DCntrkFlrRc5NDr3IGtjqUZBwm2gnTKYTjL7TmLAL
W4okoe2G/I3lX2SfvWFnWFwXaUjgvsQ/K9hxMtc9NYo+K+zkBG+wdiM2PK3xFk57/tynLas7bqBl
n3Sstv3EIYnHg++LQV0vfnMNPm0Oa0JYNMiyQ/fNCon41t2dWCJTFNHVbbd+tLtUMQ1K6YPTT57g
APaT9dQUZ7NCeywLkAUIt+YF8eL3r+Pb2fQfnJH/mDIsizfjmSfCWoBAQRBnNcXDZ4gqpR2QLGpN
FiI02vknr9b1J88jKMqULUjTCj5ScmAI+CEJT30DpfBfTHWPoOmNa/Oer/w1jxlar8zMMoWEyGlV
ZO3WVR6Ftkwf3j+CRBmlTUFiNp1bMCUcnEHxkgkCmZdptZA7UqbM2MCiy/JB12yNccF8kVabFXd3
43dO/7/gt5g+fFUxKyJFKwveiix/O5xWZecPaSbkiKpNL+XBpOxfE/wJu/udR/UpZUNiHAKzqk+Q
hRrt9NuCvB+n3HyhOF4zWNanyduNIvR7tvifAmSZK6DA7DzhQoc6k5m8aFLtc4MQogcQeDrGI7kn
awH0BPouoagawP914ihB1DiL/XmFkAZAG578DLAwSmvoOewoerHP2RjRAKh+ZAF+ZYOOX+uWB4n9
p5faIPeGMf3TIacnQFZho/20uEEC/jOSTqhXE+QnP0rCBPlavQ5LZyRf+XAUHBpaxCwpvx/atIks
D+lnX5b7ROC6SEKjMgQYi5kltwQvoBjggsmMUeLPe6GRe/+qvCTPleIHR9+zFR93m2ICBBgLhvzU
b6Wlt7qth/QN7UGKk066NtavPqDZIKizW99fyrIBZY+9E2hj4zvgS0ChAFJN5v+0js+vsnHN4b/O
EiuHSSOQnBZ31eOfg6exKB6hma3OVgWKYn9SoTJRuS+kk2AVqxdgiNpAHRyOODhC9nK0VOEfEQWD
QW+JaizgePBzJgDqKwiFwSg5mJdKtbduNJsOzwWhfe+X8myKCZLcenAeZqQKY+gCQFyGFUnINSZn
rkP9BMzGoP0QMJHovS373gyMzdb8qfyKzb2YVv5ANKUACGyx8s6OvMrM5PhLyTvv2MJxjqfY4RRZ
S5Mef/VIhWdWwtdzWr6xAOPLnD5M2jC9fvBY8/ZrV1OKpxPhp6V788MVjjUPs/5MPXx2kyC/Uf7h
GuAduPyQooA3K9YIQE2swX5ip4+tQ5dQxeyee4m6RzNeSuhCdUN938+60bXMdHrOpmhIJSXqOeb3
7DqXzdzMk/5wQdQVuAB44f6gq5JhGctMtYB1kEvnRmZRfksC9jPlLivWtuG8n+v58VRxaeZdSUsJ
neUlAhHRRblZNuMDJblT588yIGsqiUpRWKYCOr+0K2xnquN0woFMgkFSXq6cb9Dx78Tq+PRcEFqJ
p02BkI7AQUfyfKh0BC3JTMAe19mNytutkIn1XZfASOAWj8sasc2JsSdS5x3nTig68TjQI6cE0q4o
U+vfbj3myeNsB2l/GEPHNDfndBOUvxmSgEEoDDm0UOiy3n0HX1nTj1zjAhV9Ul1NcozHZH+HXhjh
wXx80zdUoZRM8zr1NxUfgPqmNRrcuQBryyVFFcZYEiqWCJiaY0M8+qdeQ3gyx/NaBuAfgSZjAIXr
uZjkum/x4u7KV3z9sBh0hewhlrhgdJzr0C7+5P+q8VMwSFYtvVKOfZrEgDNkpIAEYwWZ83PENqqP
GooNFQeAmZH4R/J3/KNgGEHe4/NVbLnoicdoURwl8NDUBqRCqx4RlFe/8vR4G4s04ZLl1UTUiMc4
2Ec0dgi8rcOvlvLcqqQGVT8f8FeqQ8O9a0ecJXUbXPvWGMMJufcGl6b5/qabPjJYtqV0+jk7kjKd
U1yq9kWfCw6UmVeLqgZ/HKphZMH258TUrwJXcs0Bpp/wSoxUHzaRn1k15PpTr8vUKQFh2oZemdw8
YJJGtUcV19Hta664Mg4CB7dexfVTqbgs9Fo07iR/XkSFNpiKksXPC2K/IfUVQHQWMw18zB4DO1Vs
NQ+d7HI9NDRCbPOwaRlFIJyCvtzBmHeyEG6BfEPC2V8jTTQZNg99xl6DI9JWa76JYMxboYuVGAmq
qs6cRky5KKJzRT51MAbeQFUN9uKY4xWWD61JZ28aHg5yW5rMNAmOL+5gc0gU30GFQFw8ACvvBdOv
VW1U1JSjAe4NzEHOZEueuv9OPnNYo2aO+lVM3VDaKkZ3kzCVtWoOzwwKHlCdH8xR+x5Ub1AMfSYS
cQiRuqAqsdA8mmKtfbtDH3sBuNjqQRrxg6SMhfg1ln3kMUONY5mbEyo01feVtkSruHKj6NrQmDRu
ykGrDGUsV1kafOXAaU4kI7S3lfFFlpsXSJUAHClLNOBQ1t2CLohwMzBlf9ERtetUaMEwzTORRyl1
N9ZITDDsLZLd+tCH7qQHSye3zcPMBIEFnZUHvm/P0JHX/DWLerX3lyDA2MLZmGfNqHgEZ6Qtj+5a
LiimYqzzncH8eqwgouK07DuI83xyBF0B8YLRgcFUvUWNAt3CvcBeMFtjXzxi7wS/XFNV70vc9Mne
Aspqoc8oBG/Uqfug/QUSNi28klQO/HYcTmRDUT9RP4SO2d3sYSsmTUqdvfAeNp5l9iCjLvXrsX0I
s9bFGHCC10m39JxGVO1WMwdVd0oT6h81JB1JiYzSFEFwz5bUuIvNJ6lxS7H3AygjSjdEjKUnOGBG
nAs1HhmWT5RHbHPIetGiZy7aI76sUrDOVbXozif+6CECi2j8X3FnSMtTT8s7RyDH6e2Ru0XpZTPW
mQUAka9OZ7CCqSyibl+s2PqnDVbZfF8+LLK4KpMvK84mo7s+CIRjn2QoDInyddIMUCCB6mbibwVU
I6x2gZIWLOIdwSupesMdqay1J1Wl3ipvy0UT5IJ7VBqF+S6Kt2ZZMlZUpPXVPP3HoYwdQgNU4WWe
ZXauYQ+kE7DAqZS38ypM/k10J8p67ueucFgYb+dh+hoECzw3sMP6CNrPUmpwQFqjQp1aKi408Q0O
UZcImYB27ErZVeNPhWoZIeqdaz13mw2ROiQX1vfYp0pJDcNZC8r994OEMYFFWI1Ph7gryr6Ht9kF
seOAkjJLoA8YtnX/cfe4HRycL4JwPk+6muumIDkj4Aur6WQ7U+ajYr8MquoJJ6FdzS7ep3KBEZLB
+r4QUkiRtjse5czRbMKjUWFE1pcTVkgemkvUgdMZLPz1vm3Zh2UBDWrCci72P7LCzmh2WArtIpyc
SNwLNZ05H4APvRs8JP9FZ5oJyd5kJ4Dujx7M6g8XV2/4NaeFFg930/vqaldaouERQxXR87FT24bs
KmMxRpYCuUmSqGVcCarWKnJu2cPuVhp0fmP7watn2qmCFIG+4vB5JVO/beYs/ZmtejHQs1RbmpCP
0kNiLs3JVMBl+vJyJr8zsgKPEdyYjqUvGZIngYV/tYyjkc96utw1lyko09dugwnov33ayGRtI8fl
9hvDRnqeDsrUFdyhm0RaD+evIsVuxikujH2jyZ4R+kxSveobt+BNionsJfGzi6YjqwJ3S46MVtWg
65a3ONySNvc2foMglJZY+vTGVk5awKldjIgWFxfWqW+Nn6L+jbdJoBqA2uqi0jMLh09RTevP5h3h
6sHNVDLIctmP6Wx/H6q4uumo6Dek5tEspDUOkzajX/0L7IZEKGN1nKu/R42/eYe3cKV+tUHctGlz
UOBxYip4mTNfomiPJJthBtM6g4CP2iM/gEenutuWs8deVTGTskR0eV97TXupX9Ii/iTYfAOG9tNl
3a34f5GavSo0OLlj2q/XP/+Vs8OLwIswtwz3gyhL88/tYvYXC9pOVTt87bX8CKt237MD07H4NqhR
I/XCCRgHAQkLphxRj3QpQH/gSkrTa5Yb7/qlAEAqh9FhYhvOf0Y1mPIXHEzGb/Nvi1SwFigAg07o
cCc+teQum2NKNqwHcVzycazOz1w5BP1436DsHo2EbdE5RQXSKuhUnotf9pSLdAfzKELIuwqosEVZ
HPBCIyokJEG1J7596/FDyyeRRcipKThR1BMHfhnPeH3QqfWehIyNF46WG4R65Zjz/6W02+ucY3RZ
BBYUusKQOzEvODZ1RtzPTU1MwhqiUVHKxcuPI3mfDX8sFOqxIPPyiMFCNjiQZMiUMwnKJKqac/gz
zhd50bZZJqtdLgCWAwK4QClDtZZDFscpWJcVd8PBDavbk9xpOkF1sld8DhJ6Nrx50LScUuG4BIm/
ko7WaVORMtWfpE3zwZeSTj/Axi6kbhoX/fDe4da5H5Mn65b192aaFmipZTkbRIVOoddI+YVts7bF
XPnnbXe3pAS2s//revQxCAtZB7jF8CzG40/Wa7UuM+4DBbzJDePsbdOSLa6HnlihFWmFJqlSXmud
fKeCmL3hBK0NxIAo2bcRcur8fRAoP2EIZR36pa3hz5qnAMe33J2zLMoF+3aqXBGYR2kLvFxj9of+
ZOzpUC0rvPNys//7CSNHonuuKYiX3pCOm37RvIs5xy9CJyaqWh/HB8xPGb4j+I9215WhzXnyEMqY
tJj+Yfc2ePINsRPoUiUHPELjEdbKL4xI4ebzAG9f5fD2mvzsIFDKLhWAGW3lv6mCKSIV3wBeDL9o
t0saTfPtncmfrjW9Uctr6z8BMKKtIEA5A1u69vUv/Llp434c2BY/NuzuyUII+B5G/5gSwm047E5u
bLfDkbjouI/hHJ5o56IHi0Akpz2p8FZR8DT93NdxtSk3ufzbULkjwPkMSO3LlqSS9KlPJVySkzTa
fLZUnEb8MfB42HpMTdnkZCMdi06IQrGsSWb3RGmEeMnizEQxBrTyKsAAJzjivqBmZxNDsqqTKgtp
N4cv9BZmi/QwsnHijshai70seIiduDwlMgBDrf8XSdEiPMYNmD9Pj0U9o0XW4iqdnA/iER174MFn
M5/YZRjySzWwZt2Nu6tKuknbnGPAaenp+nsi6Ud5pLKPgOQeiOOJ8PXpHytIKSEF58o4HG0nnYjl
AXjvsor8UTvhY4+aMhAOgiTOxqAgj8ps5avC+JDY+hhUyUN1yYvzVlAdrLFy44R3cZRRiW45arK3
0NkKdI3V9ql/NAHih27FBZrE+JiCoDxmj/Le7P5Qrytky99MHbB9A/LTTftT59Hoy9hO//i40uA8
zZN2aESrHLmy4JuKxVsuDdr5bpYnFXJHGG5XNt5bz5vExJ7EinzXYlhIm9LREb86TwxEwj/eHm9h
lLzXiPnAE2K8jswz2B0N5rc2+bR86DoA302lpy0gk32FL/jSpO0GO2xkpDgIiKNGeArF71zEwQAR
gcBbz1AdNtUU5T5kLqX+9DUm+HxwkXRgp0Ax+J48S+BKNUG2eDokXyT3TwGEhpRTcUN1xzaRYMOG
yettPV+sWvZyVAum6B2QoT+d1p6qZEAIXyABVy+RDYigboXE+lc7bNgMPgGx3vfodyD2fhlThlnS
NuuUdwm9DxJtj7feNqL53CoOwmPeqMhrmbEpL1eZrtY6zL8wgy24cfUZOfZKupcKpXDxSk4SAUCl
PSsAOJ0UP/Bjr7BQzct6akDUBdxqEMcsMNN9eq/GDvmHTtTSe0443s70Y67C5EeQKPsiPd70o2gy
EvCuC61Ji6OQedNDNxB95O2luxqP5W4kc9raciufAmI1oYrtEnZyMv00bqJPWGzcTukQytON1+VG
ivJHXkRwXzqU+nv9wxsyXiAv1rzjoteMOJZRmer+o2IQzWiEwRe8xMVXbVSl6AR3tm72uctGNDXl
3F5VZfzbFm4eSpxVzYhrPFjiTuG1hMrzUSO5J5DNiZ8Ityoc4/3ObCG6Lb05ldTIcF0GVS8Cpkdm
5GEOPCenP+j38M1mRkFVEUbfHfSZagoCH5Qr6l0ct/O3QPWHCIZ8EQRxDphxQKbvBnPwJVvK/v1v
Clem31Uwy7zBXwkq2RytnhNoR92SFg/KECe1wLIZ8O9dja30dLTtopgDQo1kDVsTKyhVuq8r1wdh
IDiqSvFVCZViiSf69UKOohZjFThwBvvfvJUa6x97Y5OfbW/2fhBaeNemHa7SRBRpFveBcPi5ENJO
sgb4Smhyrle6UbOCF7qPDV952WTgvtPmW9n7e8yXOKf4MeDRiQTsgePngRe8222I630hZnZoXVeQ
RM5LB6rAHwB81fPN1sVMMBheycFX9THrPwXvHHQYjsCV/bYCOCwLzaUjkuTd8asrdROXaCL7kAxW
fYXUQvX3jlzD/woZAG5HfbYdeWZiex7h8KHZZcTOipbWMr5NITCYSbPg0cj45aUwsXZFVofZ7eho
ptkaQg85JBwXso6JfgHKbfSjctaSIJBxZKjRmUwAlMF6AJv0qbfQtg7MwAB/OD2vIrByqTaE6E8M
qzvWXO6YANsABQSFWdpN1RQEiusBPbYh/bGpa1XDi52ntGqrQGKI0LLlsIyRyD9SlwCSg/jDtKKr
pzgK9zKTqG6kTxiD5hf5flTPc3VSFhx4mWmmt/oEpXOajqGGsVDzeNxSmtxhcn+sK0rdZuC1yRP7
opM0pB8xr8YYjU91i/Qzmz+8YVvXS5r39jh1o67Ht1+wtXww4URMB2bq4+L/UKNS9yUI8ZPYGbdO
nBO4sIUxvugsf7wNXSEsdb+n9e9lIGgN50zS4LUbYH8/dkFVsdrgfh5sY6gQIfmcf1PwEAr/jjHv
6KRN3rO/Ek13G+r0VcOh2SGa8M6CiCRSIaffBSBrm30E1x026UWqCWvVZJUQBCNZ7a8ludoC2AxI
VCmrBO1AJGGGNvQ/hQWSRfgGGelAhP/R+KMbOidJNft5MCbo57SKpOvSkD0TwjzOn1ILRzD+yhpt
S1ECkkUqnDlssu893rx1TvTFIR7kRJJ3qRkxH2sLl8fOaYnQsK3KY9NFtdJNp/ERsvSzqWvGZM2w
hmeVvQ5S7VAmb02+1VskCe0DBSUHuS5TfXkisPZ1D2pksWzH3NPnast5pirk3Y3d+tREeECEfH4L
mHDmWNhwa9dtFahj3sfBG7igqxhfYFr6Ro3QnK77t7/Gb4Ht4JGX8P4aAgg7iIjXiU+MnGRF4YW6
8WbGpQjoc+t1yxSvRH2ZR9PTzNcRiTdR8gc91enoKTROS+Ytj/2sZ6m5Iuent7xogw3xo6pzirla
s1F0pp5SE5o3YBo89ps/GmS29Yx5PpJkteFywMvPfz9r0PCVjPFQiXwkZuYod2FBg2LewpCF6mRM
f5uTNXWvA/1PE+HKZQLvJJJ6JFOhImMsyJ8Sp81r026CasA0WOf3cs3TyepX98+3O/sNuiVFBLu+
0xR6h6d7eX3B/oCAclGqsTWnbunmSkCjlSW8HFme7V9miUslq+fxCLlkNUKiLgFN9yXQyt8w9f0P
ja1kjbAV5JhIHcBPKRfraWWeTRBEhfFLYwpdCyiMOFCw37NNyqeK1VefpcG/gvIEiKnUS7Q9l91E
GZcf4ZLYoy0A26EhWZEiln277BwaaxU5JG+jGSkf2KLQ2N73ByNzKjjU/EVPmYL4nw2MJ0w1D9UR
rj9pWJp+rFbjonkggD8kYBpHbM477QLdXtyNHjXtUg0xhkotSKAlGyhcWBc+65XgJqsv/FJPcX5M
O1Vcf2OJ4L6RYD2vMtPvbrfvcKfDJ+sr9Z/6iadq/9mouLibXMG7hR/orXDzleCkOHeDEFZYNe0I
8TrcUnZ8s+SyJpHy+kXNCxQ3rgJkOjh+5LvTgDv+rUIDUtqSbYzgW9yuKZtJB2aBiqSjbrlIdewG
P/5BSQbE+9injfGWWEC+L0vKGWTe3suyFWxPBs3VCNCDJcRt0K0SrM1piUTlyopQutCzldgh3q+W
RUg+subn8hQHbhJ1vxt0r1n73Xl1PV7GBfuLRP98dNH6wTNnqy32GYEfrCmGBPvBXShTa7geg0KU
iU4/UjHMp6SGISIlTV+psTniNRpTaf02+6aqudFac5KtwZXPyqhDalbgSFHiQRzSFANneWQU3rOV
ZPpiGEnwSkKfZa9LrECDO4ZNT8XtcuvaGJ69kYRLiCqEym2tMax4iWcfZ0/Zi0jMLPa8qVcPphy1
DHFZcKg1sNoNXY4Wv/QgXp6dObzXu3NmgSjOccDUAQM+dr5Y5xtdvi4WytddGU5cfAKbmk8tX9WF
9RHPH6P9xzx1YlNsv9AvhgFzLJwx7L16qH4rbFTySzxIubtvUGtYudJWgjYXAgGNdSy5gexRRII+
Ub0j7YXYwlTJ2lSG/1FRoqKcEt3xLnciNi1XhKPCZYGSxyko8mNB+m7MS/LSL8NuwBD/L5SfLIiO
M7R0ZTuhvKxgVrv/mIUOu1ZCZtuJX6wtzKQKmwk0odH9I4uPTHxxaSk9nu4pxPEwpvLUA9UrsYlM
rB27pFH8Jg3c0wTBK3ENFfTFkXSnQMRzLirpUf6ouWfYcov3FaB+C4PnaSpuh2I1kkqjb16keLiP
xGaAEPS3nf0SdizZLSHu5ErJWvPEvpDIVLUN0r4cLzB2P+zE97p0G6DGP3eyiy8kZJiFqus64z1F
ocDqILMHtCqs0BeXzvv+nXQ8vfev+Tb5qTobqO07HJmNEWxUHAVukOia45BQoKlkGb33pXcmz/n7
g6ypgvlgtr6JpP9pjW1tM9VAcnFUYFhjyt3IhuphCK8a0H7wlI2qlhz+WdwRFGUTuuX5JN211voK
PU5gymNrCvcPMChK4tx2AHV0YtPwoY5JW4bkmE5QuXdGAMxucmxvv6MOjd33Xs++kolaVDtrt7cq
JBT/HSv/K7JLTqq5t29tBXsUCLilE0K58lNGKCCKfjUCfV/6NinyBHYMm9UeWdvxY/epVMNerLUu
FmnKPsYA/ZrUXDPWoM4bE2uTqHF2anXh8Ac9phu2bKhubFyPdliN+wxM5tfR+IhNB0nwF6XZv8cZ
7lvQLJv037IQvtEafSN8p2HF3ij7N5X3ggzS+Sl6ErQnJlpQ1gIwLGTGrqnIECl0uXIQ1oueLKjY
1Zws3T89jxkTFJ93/BmAZLgq+21fRSKXX94cOMScFX7AjEsO9aABRXOSGGqrYiwR/MuT0/v2s35b
xvIioyL2UbV9MWW/LShQUJXEd2JhmKopSU8qLoJxxDHyicXO3PeoRHAPLsV40LfQUr3Vs1S1IEZG
O4NX/5gD8BMbVJW2T3mMDffhrV/XfXylWHQUXs6tVlhMgtZzzQvfqeBTSdGqgcysVX+4d3fe/kxH
z/qY/PjFw/TRE7XJ0Q3ziHDwyrxCMyQJqbQjkMURtQIiN5ELBN7tCBHl8kVSgQR/LTfmjG0QbFpL
xnRZRDxBTAoBWhfUAf/7z+a27ymWyAHH4iL/Ag/GmC1vA2kuVaXJbM6gn3BcfPNPm4A+/H6a/r+5
T627lEaavci6v+cgyV4B/58ZhwUhafvvNVPHtRmPP+Foj9pcNpyMm0eRO82gQzZBZgn8fef4TtrH
s3GwUSS6fWSiNuLOXGHnGCaKvXYlYao98HWjJ0TvyzX4nnsn29D/SP+9jrEpcqKDz9j5S+vzi4Wv
VTznVVGkzJPvwL/dh9Yy1OnqnU6b9azfPD9b291ua/mjc2MPrBRHj3E+8xk+OFJfQktd51T/lQ+7
FCfQZTWyUD1u75HGhbJStnaoUS/Acr7UebwfnRXtT0mpmdsGudO5vOK1nN0UzLO/7nhpLz6CX9KW
Fa5+k3OMhNemasA01tKsDlNYORxF6vgPgkI96S0xDkTMbewx5jOLxdnFrSPdu9YffaQfCFhuGr0h
PQsEDNl2r2/lfpGJIsdbfHiT4XWAPL8TcspKss9XbGK2FuBmhZsUlJy4fZ5oz1VjkpYbmcJPhhet
43UqafVI9LPCs8tTc2KzYn2MfXYdEUSO1+nBH4k5d7VN272p4V56Ukk3YbSqXpr+Ct/+5lvJGBRc
9sYW1bKQYZqqewsQYo7Qm+/AjvRtZjDrm5mMZpSpknvauQf7/k2ktnn+EzLP6NeaZUZMpt8OMQJ2
oakEEjygWgrF2OUSdjiJq+TCRa99v9rRGSa9NkcLwF/5NfSkd4nCvigopnQu0LLueTDqkhcXlLlM
k+D43UDzCOn4nYE3XEKq22wvLVmw9vSdD7u2PetwDPwnIlOkjFl/Cnq/OG4+WXs6u669O7AjEPoi
KWXd4ozzJHatS1B7ue/kkEKGY47V4MlUH0ywOeBnPeX5FFNRbwXU0DcNP29exze0wApLgxFQQ7ks
0XStjv1ttFygIz5/d3q9dDsbKeINoW/OvcnYv0CxHqXpIERefFWYYyrjws3BFMfk0UMnHcc4G7Ew
eqnxGN+wXVmqseYM0TS2KSI2sU7IkdPX+Pu34YKNtzYQZPXvkw6JdkQLrSyNt0/MeqsWdAklXHUv
FMR67HQ8WjAbTb51sFzxNsuPwwpPlbgrP1CLW1WQeFL6LHlLjpzzw3XwC6W4expR+y1TGI03+ArO
+1qIRFZx7NElNztXnzzB/9NipSSSu5kwANU8fvCIK/cGgSgbrQPdjHa8fBaGrYfdsiqWeYqMuvef
iHEV5EKN59IBVE9QLh8G0zgzMCBN9Y+nt8wHsts4aHAKAWxmYB1GW3TfZb8j8q/Jo+is5+TVhymY
S9tmz60o3MablPFWgxUkjCEcYJBZ03EqkBH7OxNoWZ5wvafRC0MACwPCrgV8/Bhi05he5553J3j5
p8mxsZ1ois3x5LO7PJ/CFekQtJruqnSlR81gMBWc1PzHHFvGfYrOm6ipzXNWaoU50wJD3hJ/eaYp
mP+osaxayyWtTsyHQPUtnpsUIqz9f6kxiweXO9e7FXrD7btQNdjaVn3ES7wJanjr4bZxnE83/+ZE
IR7zunpLrdS6orrMmqEHe08RBrDXM1/ViICYe2osf453pIMVbRMzSqvSUFh53YWQHgVrP4wINosw
M9olU43sM7Na1uXHgaNuQDpBJtpbv5XZLMggzOOJo06GNCA9NzYd0Mqx/qmHEYYgpSB4RC5Wr5bh
pvtn+rH8IXVu3Go5rKPtWiqij+od8ngYfmP2A/pFqjIO52zkFexxDksnfUYOzfowbNimA22JhM/H
k21R4Dk3pbDArfUVgYviZKlwZvZn5gDeZOBddJN0LfqAflKK0Fw5fim/UdtwHcYTeV4pvA7lhcQW
RSCs/RAZTXKz7xM1wHxne+NKazgHjgshf18OgcnH++Twihyc27AkRY9lwFrm01pn1DR6bbXi2ilp
8gKobx208DiXDa632SUnTjrP59jdPXGzRQ1EE9IHyQbMmj6/HdsMUh4DEl/h42ua+1qSy0X150mz
2SdtRjP1GO88JX6/rttOPass6xf3BIJ8AszHaOlucDf0hFVbgV7ZMcKfBvXXy4HraRMZ8uvVDc+i
bYaMmK0OA3CFvVuBomaN05PLIrypG12x3lDc34VRPQcOx9/gqIf+7dVKf35xFun1r6jd/8m2fBel
zEMhf4Qw/bWIsC+qH8SUdii261Rf/kBaHNSxGk0uGsC32ckrwCO9pLMy+WFxxDS7n312Wa2dVOnm
ZQFkUBzqdG3MsTy+3o9oR3e7XkfOUox3C9Xrjkh/XOaycypeYe1GKLbP12PePJmYKwkKc8KuuNjI
J4KjzKlq3gOYSFIOWjWIfAR/LxmsoSrtI+9k3ZnJGOypFe6L472jff4mn9ZXEU59259jv5INduOD
4+TSljRbySCIam2kLWMivXBtUndA1M2Nd1AMtjAp74xZ9qa/hjkAmjQdSivNZS5jGIBofJmOw6pc
lOZYu1HPcHBOGHtD44E5zl6Ly5yD6O7KCJPJxg9RYLmb6X9ER14pa89lxMbFd0Nk6bi6sjxdGdLz
4ORIB2IhxR/WqG/Vkbls7Zn84pCQ0riO2ilPKCbJu4RhLTKLmRg7aedVEfR+M9ifnIVfPdxE3Uc1
IpD5ebtVehbicbrP9JTAlTkL++VGDAZP0BMPMNBrjvD4EYav+INw6900GhmrjewfETE5JGWF8N+O
dbHx0ZQE/e2iiyFSQQGFGcnk/JB/oD7r6r+HLofdZK4N8H4D3qfF0eupq2dPWzWtXezS630xJAIM
/jpeDvPsHhGv/EmriN54X8DKgVs/KvXRUE569BZHaHZkTDbjpBrOhqMXVkCHXqIRWhx32GwBrnld
WkyUbp4rCgEplJGg64tXUOJDmF0HZLIeulNXsKNol1/FhjCvrQUFNpurhQLS42FGNQnm/pH9aZ7N
8mSLdduKs3VP+LPGuKyVMqOWctijI5X8ymPEaEsLimvJM4/MQvgk18o6r82R1FnayeelcMje2zPv
RZslkYVlYTaX2R5/8T5EyGWPLm4lb2u/NFM6l//E8fggQoY53SSRgqymmCv33VQX6V330xoza/cl
sAPkXiycInh9A5eppd0BExfSZ+o0P31qBWNxcJvdt+RgBJBK0tB0Hdivvof/uNn+zKIoC9gPSOJz
bT2sIJohpJZGHkLMN92Hb23tqg2/m4+APL54hv9KEV7webfoEV821dDA7UMphKWDC5Av2HnGHL4F
BOrSVtCyzbzJ8wivNe0lW7AvIyAoi/G0IPo7n3J6Srv7tBhvyMv1HQzn9N+RJezx/OS5BQlSAPpd
NNXZpWhdaTBMvy4GBgpeaAnoYqWhTgebwoudtuce8yMwqVA1o5haQ/dNsV+OVIC8bQwPZyhOUIDb
RmUXoAgVQahUzQedRvuIBkqjaYDWGwpXwr4AIfIKBDLNZnufmAZP+ww5HtsRRyL9RL1aL3TuOW+P
QKhVENvLlW2JKEVBWubzPQsN38mpOUtg4wqRScML7J2o7momghl+uPBRYDACaoxQoNEi3H0vNcet
n3gPU019VHGwLUxvpWLlaecI0FeuumoAeFbqIoMS+glE/DNfMWIAt4YjqrPnTkMNTgs93zjOAKVM
PEgURxUvW7jk6YkW1iwe73UawzvCUftYOSiC6wswQE1O/UIxQDI3rExTL4R5eHIrz+mh4qdf1cR/
rXBUOsl/xfrkDYz8mo4+mZrjo9yVCPu9T9Gw4oiqZOtSKaWafz3kVkKuyZuPYU1y51c6Q9sPz1W4
vEzPDQF/8nds4WdEKi9lX3GDC3R0BFv/naK6FonCLu9ed2sqtcvJw8X/WOf63kyCDjA6QGsr9q7J
jYv4fL+pNnNQlX1NhLeeI8NzSZ8sRcOZds/Xk1YglVCxaVnW/qq4B7QNq7Waz15y2xRX57778S7J
334a6OOvREnyTyQ6RHaN85OJ4/6DMwZ+v7sWT6ONWWXbuWj0F/afuVDjupyEr1AGPmPOjfRrAyW2
oSEIi4Z9GqTDryOegZp9Td+ge49X/dGOLOkiouXzhfwPOkQIorn9jW01vMtlb0wuaEBYc2sqasPf
Syicx0MTWBouiL/SO/2kHtHR2gzpYIEITVATh4ZPXLCQeUScnAYTDyyfLatNJNMPKamr3Wwdn/rU
Tiu5qusgpwJeIKZAshjkGTXGSdy+tW/pdhd3r4WTnOIjk8H02Lu95+e4imVbB3e6uXa1TPnOpC3O
IyE7TBrjZoHNbmBGFVsXBnxWYboVIapNDfQVNip57fdsdldO1nt2GyQjVTYlLYUDy/OZXJbAXBWO
7y3rXSkh4HDv5Fc8NFBs6pR9361OTcLjWXreRq88KOJoXpiAOfNbweV5voSnXJw6iG4qoafw/ld+
zeJmzBf06g8wMaOhHycng4EbyU9RL0p8Q8reuN+BGp6Itv5qnpPAKmyQaBog0detmPaGefq+KC6I
A+q+dp9atSwPVF08wFkipJSHkARoL0U580Pq3msiyxfqRT1M4dXAyW4+kMeVrbRpBiUUkaDmFIbH
bd+3gWJi4zFtKffJWIDkBtZmQhhw34T2I4Qz+1TKea2zUrUiFE/7ijSwAbZ8NsrCzQByrCB8xYK4
4HvCBDpy0/LiLNW+SvxalwbFh89u1QPBz8JlJtkMlmpbmw4D+RBFoMRsdO/XNpTwgk1SyEFR8hlG
Cbf3Ww37fK61UId7a0UOWV/Wtt49zpdwgAyetuTveQqGerO3WQQC5RenTL3rInEJBIGQls2cNGFm
x4uK/Db7fTx6jopV9CA4PVjOMSGyYa3ktr0+7cYwT7+QgJNs1Ig7zAnbJeGeJqXgUB8kt2xLLggF
CoaIVyYa7z1vO11C93m+SzP7VlAuaW12f3lMYcPzdpmBRmWEBle7dYbQQw4WRIAkhbpzEeFvfWzk
DpYmq0JHMr2/JU6H6DT0XvOzRGqQLohjmXTde4W/QdXYj60eXLnWE8GX1b87/xWbhyn/MMWOblyj
nQL/Wxn+t0TBJIdwKms177eHr5MaoDHzWqsH0FVP2d5aPtUQllvBmYTTynYaLx8jZnhyd92914pC
P3rG/Dnz4U/cm5Hc87bdRbDEtAVOVHc4POTh5Z4nNwsxpdUfGwmc5G6jP9EqoQ0b0IcPTQVGvQpC
U4aG2wirLWCJqhmV9GHfNydTo/2ZmsiAHKxRBLjunfiEFfSq1mqhLnvFcXYdAsGAza5QTwIBd/JU
5Xv6RWhRYT5bIwXbHByq2s37P49FRjHWrUarxpc14rI9N2U/CcCClfzNhjES5DT3srwxVaJVdfiv
yo0ux/zA38djUYAGZy7obulvUB/0QeQTAHruaHzUFvqIcxSfJk5AO79EOeYhu5jbKFko0vmwYepK
mxDhivwbgKPGYQIOcdoqJr0MDcDxk0erOzF2c9PROMIjbWWCaIX5It5rCzZGgMbpMnqBfDqWSpHY
wxcPOL07ZAB0S1jFIw3Xwm7Z2ALs8Ep1WYjgpTAgdyqGgQBzpe+/n0PPMudxMj8BaQ6jag2LRQFv
c2wkVxKoUgd0cKG9VjIouFQbiglT2eqhbiaq9OcJdB9jLuBpzfdo1s7C3qJSBN0G512F70wkreFA
JMJqqdn18ZQkgqBsIoIZKP9R2SFqNrcaGGAaWms4iV/nQQsYoXhSwsXfqe5hKw3wTywHrBrtSVUZ
H/1Ual4OFESbBlvBcikUu+0xuuvvItlZNZ3G/ans7z/t4bk7qzV37JCVmBtu7VsNK/1dhKll2osn
8Llo640niiLByiu1g1c2yNZjAmKnUoYD3/XdiKUV6sYLK/QitfUXSFpc87VReEc+TKmV6YVqLQh6
xZ0sISbelys8AyfJP3sqUF2X8VGtgm5ShSe5EXrou8kDiuqeffvD1jGU7E1h/rH2HVITseaaDirK
av7VIuOFRf5Rr+CXBz0zDGmdcYuX/gzhNSdxASmiod6X9kbH1uhfe9Mk+GJk7w67nisChD9u0fKR
V3+0mXYquq2s7oDr9Xt982u4n7AovcE7Lu+B1ju+4QsL0yNmL8rFuDFm59RtKU96nRTUq7URrnuQ
N25eHIbvdtn/mUyzhv+1Pul8FlhCRa0Bc149f25N+4D7daqmPukfLIetCWgTIA7fU+I3tTkOYEyt
q45THgA84pGc6qF3ordeCN5tFbW0JSdOAIyjXo97oDvgexkYEy9kbOEOhQGi89N3xw0Ek9xljOSr
p8x4eaAyjzp4UALvNxQUE4WFETDVGvG7N7do1OXfQM84+V7gInkusXf2RTRnt5LNHU1ofFV2n1ie
LxWqqxES5dJIytxDMW6h++3G5fcimIybATFmecuHGvZdpTtTgK2P+0dx/dY76EZN64x+h5XmBatP
Ri7eWkrdLVM9sYjhLvTp24o9Y9VR0MC0V7TMFUu6fKWOKSODRfeydPQvqGFrCrjPX/GZqxTt8WtR
W7DQy/gon6R4XB2alHzqDU/x0DMI4WYGCix9L+IK+3KfsUbaPz0yHIc/5pBPCKD1jR8dsU1Nxx4A
g2I2hCnyzS4a+FLFRYrgJcIufvdrWhiZeiDLzmHR5brlKjqgAinRfeei3GlaeiMaObIbNlCqaaWv
3D8i0Hp7lqtRZBBp8toOANDtcotAPBL0U2rG25+nJAuAo3TPxT1GHBpdwPl3lpu3m3XY+mHLvMrn
5gE8emoLQ64ojRULED8btz7I6/NJ1z25fYRWUiWqIYkmZC3qvgaOTBTsSNL0O9M86yNFrLZJGxW6
KP2ut0W/fNhVPaHqerN8cEiJ2av1wCy+JnI9E1nwcmUH7J1UcggwLj61uo/wHA9sg2waQearKnFv
OEbsqhh+RTn7tKpGFPaneMz8UyFeTxlUYM6vHVxUkyRMsqlebFnOKhCM3uIaM2WM5e1BONJJdlqr
b5OAzPZdR1xTRqUi4nN/NEGCvn7E9+p//SThJ7HRcmn4qAVLXdKmfoQDvSkSNGIori0dTzEpl7aQ
T6ZYo18IvVkMavkcCX9OGCp7tF48nveywu4M34xt91ddUb39inxIrs+BeR1sI7UYWO7QpO5cUgk8
Zfnu1Q3KglgR+7A1mDxJUvXuhMhlNuMnGCgXU1G69lXNm2CDnfteDFmOgSMtidBgFUafhDqbX69j
7a2h63fLCyOX0qAKXfeD6dG7quvThKv0h5gO98J/UqQ7rjFNjpWHKGgZg5QffDMqZAJHypwYa8oy
lFRu4P5nyknGPjOsTp3CkGUv4JKifob4aUW8LEfBmOWNSl4ZdmJsYFNPws+G614gjk/td54CXm4L
gAEQppbJBT9PdjB166u1Www+sfatVhcP5bSXstfL4dKvYw+8a/oOHsV8R1iWF3E86HnOAx34kJp/
nZERCblF4Q9HuTedEaQNZyrZbnsyK0M7WYugdpmIR/4LXGuqqZV33gkj7y5RKyu9Wh/OPJzal6iC
9z2KaWRkMr3Ov18D5tQWXiPNtNYys7EqpwUxvQOR9SZSe/TYADdKpMJhIhrUCQDsbMUNlN/sn1/k
/dUnCLkQjyDSfxFPhSMiuJST63+GfyF3IcaedcKTFmxjrGnxumSpBc0NTFo6/wwdvk6Evj77ahXo
PMqJFMZskevCPFlzYnNicEtcFdDBHBog+BkXKCxl69ew9Rn2XZZ2MEjZVF9OsCOfSIX47G9hPrla
kMnu8VL2gtOXJbDa1zL9BnkIVG5rjSHzTEClMBG4NVkiYrTMCiWtwPYgXsnKnn3zlSV9aA88js5V
Wz5m8rpp8edvt5J7CNC53vjIJXgkhwamkI0kSPAiVaz5ZBRGdDxcQWJqt90hx3ACdVnMOoUiyQ0z
WH/BaY15+5QZyD3AIJ168oz4pgengQw+plMIQwTZzY2tDkT1LNRzEYzQK7O9Brt0Jo/kaZYWPRu4
fa5tMmkfRBAo83Ix6SXBZVVAAT8qCt8LBXc9ivo13s23djJskECslxX1YB6mmNK3HXoDmNQwvuQK
X+qpVrog2F2O0XFrynYf+IgL4g3d1IPDAkOoIh7VRWA3W+wLQ9TpTWU+7AuVB2FaBUIge9obnTz1
pQC8zaXwMqaP8j6haOS+YYbY8QcNzdvlnOUAqaZBUC9sqwAQVeCOlBHzm9IEnhdRSXSZmDqYwRGb
aQYLNANZAEdHYN/1gyEJOXRF8kyymAoS7DjdL9i88B4rotq9yG397u3j66AeCUe04Lf8fYXoWTg9
McQ24+BUH5SEItiFV1kBJ2Hd1UZrG7U5csiOQ2/A39FVcZb63GfgrhW8EfEtunVS6F8DTld8sC0I
tl0MSTSFbCLELrCYi3/K7pApVluaYupSt9x8Wu+j4wpZOhEeu7Ii4DyB4yU+ZSfKX++CNUp+zUnh
n+X5m0xfFKVkXxhHKt1Ub1p9JJMzdtqf/aY15zBaiZdsonelLLSyVF7KnzkRE9bTcGk7OBw9g22T
9CI96Ha6g/jUa8TjfWOWoJN8I77Cjh3XqaqDWSf/z2sm9F98e9ix/rg6FX5/0wTGIdOo1jf6qq94
NVxvpi874hi2l56JKGQ/c0IXxz0XkoMDqEuBP44hv3pn/DnJLFFGJ22+3X/jB42fN0jJj37/3t7u
WwL8vMRhuoy80Oa7zXcFrBybTYAiVdUmQh7x22fpneuZWOA9x4bNMpT/2rxzZPR9x76d8UlOevV1
xvbWkclGdcRtsbYdOEjs2a0OajdkHMjgmLnLvEC75sez1CNoA3nUqnetEwxpJHeKzeb/aVylw0s6
Qj2+kI2X8dUyV4UQq+VVsXc1t/gt3dM4oQGeRL+eeDb1yZtTRfWtleJpVHxTUw5S4cusySTcXcMJ
xVMKONr5rU66v7U95rpVc1gpB+zKXEGFLhyBW6FALmNWbLSq1BOSBWxGuGbzE6uaRZ7+aZfP9BqH
X5yAaXwhQ3sZtdEsDZlPF2UpPpp2ZCX6hK5aML1WQ2WiohiC7EFc91as1o774GEh9sANYhCPxaKo
WbUnvamRRJ1hTxNdoBmvic569VjTklM9G2b4yG8ILcSvhTkwWPKz8E1jaafeBQ32HwPqLlsM8K2F
+HaaLAiisTmAezqNB1Y/7pYjLT/xWpsckR4dM7WdjQ5sHJGWqdxXB0O9eEmsK/Tg726VYcnyNWo6
dAuZiRm7+0Q4qOp6TN/Trl6RqzVw7c6idUuz2xyDk/uuxPbVRYCRS5svBByfNRN7wfj6Ot42il7F
XBf6l2mZ075/kIglaBtpjDnwMUqx7MC2tpF2+bvkd/b17c+HUm7nxwmOgWVeTgrZRd6pMPAWghiP
w+Gt+VGttPAv5gsLiu0EVpX/r91eqeM/F4z7oYVbcxRsDZfipqbOyUZuQsEvCR1WOSesyxOUFZnJ
tGOtNQFlG0rJxMYtRF6jEGCa0V6JsiGHhcZoilN+TShng8gEO0ZC2B7WkaqaGWggUnwac848BBfw
R2Svmj39HvhBdGDYub15ZRa3hwTItCs7rtuhcKW3ac3QbEPNYAMRb3rivX2GX0UfKN9l6rCiP29w
0o1vvGgwgzL7MYwVbnSAAWywqTJHOpfsftwrpF9sZU+mo9inhHIPZrfd/Ybu3oXCRX9FXRs0EbCd
aBwjUNiK6t6u4WeyqeQBS3by1GzPSC2MaBETqzflJmtVGD47LGFojxWFgPFNjr+no6SxU1qjhfVp
i7RMCN58G8rCPeuVEZpfQcWL/t+RkjAaN5symsE1q52KRHJi6isxYuUFT4aZ9AUP+QWN85M6n1v1
9zKNEJehwntH0U0C3FTLbVtBF/ML2lV6JLH8wRLFB8GmqwpbwuPIX3E3vIaVk2gKX4ZVQZy4JTRo
2zsb49VK70QLMv3YNvPD7LjtQV1+ALThb/vC/WBEb36nnLxslB5h3M0aK9c0/t3RV/rYFEXX22aL
F34vqJbQpG8LOL/zS9Cb+BCzA/YjqUZsyBqgtWKKKtpjjsh1PcxSI/iRjdfBK/P+ALeaQx6jHnOt
6n5z2wQ7WzMVyW0TCS/OCjowYPKUaVWoKt4Hhs9SAqmULSX7g9fIkYzXmidklnCC0DTAf4TE6IOu
TvyYBwPBAk8fsI7eNJMa6tQRiyc1YSiTToe0AnvMvaHyh+5hFDPg7jbDYnb2oXhtXyw72Nd+2ffs
uMU3EoclkFiN5EO4kJ6jwnnh5M+mTPpmh/8XTjD3O2fdUCdVaYN/mfMT87/JfT6VU96gbm0r58b/
KxcVH+9fpnzkr1sscqwXD9Qz4VOcAUvxE805PCmPYRV5kbMclYrFvJhgttJA3FrBbCaGR3UJ6393
RZTfoy+nj/GYHV6VOzBJLr7WYYq7SS8igS5JzHCuKty9Arcvf2vtpK4gZhAvKBlWPDKv6l/Amsfo
VqD1GvWg92zs9PzGNnTxR9vpR/xYlPvDzGhoJQrDwhxkt4BI8Epc5RX6WLLaynWZUHDCvr9RFg9r
vjIRdvTvHNN6C/azoyp9Nec8zKLY+eOju1M8tk7ckKozPfy2poTuzM2L3Hxglz2zEs3lgYibxZvX
fcgHKBqDMJrVvKcKISoSmDYsnaxxK2sPI1Q9Wvp0BgT9yA6BfyUJKdPnQ7rpiZdPyHY3O1yXm22+
DCom0lcB/PaTxm26lHXji0vzezbWfRSdij4ItYHGZWT7kNZJucAug/cUWkW8pHK+EJfw7bGh+Dgk
BV4CWkGvv3mMjB7t2mCHJcb1Y8TAvpYR9ueiAighH0sLEyVoYOeeexrXswYLxicaq8WLp8fCFe6W
9ucfpvSR/SIiTAyOu9NqWnzhQwrV3GEyrhrXv2fJnTTYNihtkCqNNUxitNNbzQuFq8WU9liD0Rin
w1xxCrxLIAq3HMMl2TSceiTPFl37rvz7oMXlUQ7FGSmtnor2fvafVB0f62UM/1auAQE+5Osw4CDl
t8gW2NXcfQQQTTJvxCRIQuRyFr1VM0KcXmiWbBku5UkM83Az4UPGiV1A6MyEHESv+sw4MWhOhkX3
CdKhyONlBNumkn3TtZXMVbg4jhuE7WnItiXLGKv+X4/sppr2+MFhRMP9qQN2CxIMH0Ru5Wn2I6/R
xXc3nR9S1RAljQDueYMG072Bkm4tHVFPX1PIJZFMRzQgQvtsNvb9AIeN8Hs09dmmgIXANYp/csny
L4QRsD79tgkaH7jatlfBEhX2KW4aucfUfhv0f0ODV149PF+iOMVlC3Ydob17TafU32MNpFMCvkdq
rKqD/wKSn57hLcbXI5KZM0v6lZfJ9rXGGF6CWfV+HJ0b0km6+6cCg1MN5z70Zv59nFa7zrNM5IuW
0WocLv6RsLzd3c0rd1TjvyzPJ9ALDGfCOzYucQLzKKVRyIbEa1ayTzgSpo88mOLMUa9MS0nxzTb7
xgRGFRkpi0+taxieqGB9Uc1tXRei90FHUE6tt0XgCNcYeu7nZXch/oVqZbeLSPWjsHZ7GmmNtwB2
bEZwuzZkX3xrmTcS9qTRado0FqxlUXeR9aNAz5z44CtPu0T5SjtnaWppz6jslaIJVShmSdnWU17i
FOwKzu3vUJIEPCP3kAukIfoBBP33iRFq2LB/sn9mYZa1vJli/a1QeLDBGnbuc6hq++bKmAQjub29
P4i8VxwzqwXP00ghvY5GtBg4J/WKoaOlgz5e9HEV7dIn6f/baJnYjN3aSyHVcVV8yZdgV/5C5T//
b8StdjwDa/W1zF2iu7+x/dIk6abdvbdlBTYOTpEnn58X9Zvg/K6UEpjnLtNMxtmNDV9QQXgSdJIQ
pNfJW3+Cc9PYHF6siRdQ3Xh3LZP4miDq3rvV+1wY0v4IshWfidydYeJck0eCe9qUqmGJXP5UcupX
gpGPxOh0ZFOESEdu+3zczJX6pf7w7ITxVDzo1HrEYXJxaH/2sDrbFyz68thmMyq2uFLcDF6xx2nb
z1SXWKC8S12ySz+18hfZJTXqPqdpYqZttG/n3QrdTV8wQqnr+Kkcam9ivciWTn7DshULCMZPbNh0
9pZHwe+gbtJVdH1jk13+JzQq9QF2E2UMQZZ3qrCPzgM3NdRhn/SgmKdepJLPfSWhPKNJsgsl52bc
B4jq2ymVtRlMmuR8MNE1F+s4UYH6Ab5M4r3uGnYwpl8tXNhlqt9KWqrcRCqGpjS3Db0pIA238ZrM
ApdYOqdrHcdLKKMj53BnUIWDYhczyGNOue4v+YcEsmA2P0Dx3IfaQKv6r6MLFpmpDueqg58vV8Tr
LzaRO9pIITcN8Lw+wZTKV6inwgQUkNrPhycxJmKI/xdT9J8WIXhEra44wsT0reZMQUJ26NjDYuo+
6a4ue2DrU2d/O0QDngxUUYku8CKUfKac0Ilqc609dNhJ40XJoqszXToFf4i+8GPFXEdLJBza8PYM
dfeymIwRPt0OD8D4+/7aHlR8kiujdFbV0Bo1w7DuvYNvMmoJusgRjvTWloSRPXgyxYVrTQuhxXc9
TDqjB7bG3zrLelnlsNEIZZyQNOpxbpPe4SylWQp8oQLRjmshT0CNeaXf2M0N//VGDAipDhcvZI+Y
JLpyTG2sVgdHhAVUr0kBgBxFktsyt9scf64LoB5F4Je68kgo6SxVNc0qvnn5BNUx0db/D5zYydVB
E0BaAswOR1k9Ou060D8F9Aaksfvj+0ghZF+tmW/pG9CsiskzxpwuUppQvXruN9QguN3XeiJlK2Wn
nziJmACDzc+KykPMthQDSKkrAGNLNj89XD2m8BY8nsf80ua88Zv5GxG0IEvftrM5ryhn67rejF9K
kLZLwtTdjvWcE+udCfbCwFNskYHiLV8Mn48lMp3kQB2iSX+xWlEjN5pThWIH+E+NbMx13gVfLw1b
U1/uy0xfkutVSN/1wzCIynTwMeqWoP5Ie/BfoHOY+UM36KR23K31grEs/fiSuK5DsSPhKXuaEyz1
Xle//eHKbz3CkXn0fPhd7dsfyMMHd3/roxhR3AzmuvG7ZxxVJBA3xY6I16kIbXzDkSNcU4G+8NVN
B4Eiw8Ekm46FZc4QnAQzwwkn/xAp0pvLlls366kGXli59sOTpDVmqjDIRtvv2i3EKRI6uy1cg2lW
hokJB+/h+gpRwMeYJsx5tf/v/xZK2KKM/JQXKdlTdtt+0IERYIs3po9/yDt0NU2ggp0P/uI1mK3s
k8hdqwu49yas1JCEZOuEIKI8niddJX0hrTGFL+pgn82SF8Zw4wIDLNam2MS4nt9lkok/T01F0T/1
zvCvurs6NABXaFM+JH1gjsRoIFiEg+xJYK8retJ1gme+FuLl9n91csRXM0RgUV4QQWnkqlWcDqux
NsOz271c/zr4u3J1cVfFxX3U3iFipWHqyt4hsQVz7P4g9qoI1SjZGfGpeqEO3qeP3tVDKsRt6SRu
rPpw/JyMUZFhfzeju4Odp5H6uQPqIKRVvLMeEpppSJGVgO0VJEESY+Ru4mp3AZg2DbdBgX3XUzXK
mAccnkaObo3OemEFuRUCBtuYoWI9l9BM98AFTN82XCIiA9sVWqa4zSCOM1pI03NofVg4hId4JLw2
w/rz8ufe05Kh/L8Z6/kihZfRaGryVHL+g8B3kfnvPC03BF6tO86gRsWOOmAjzbUYrLEI63G9mRNJ
dMRu00CVvdjb2xkIWhgcrE9OyMYBJ93/p+DjgowZ46gbvhTs1D6xNrAC6IAn6U9+K1bbPnKFpGTg
3s6ZdRpHJyN0X5klLwMHjRmoBBIsh2/C/CZinT7Q5gM/0mfl9RgRNCg1fvbL9SaroBoQbYmqqNBZ
eCL6+UNdbVb4Q7++z5e60B6Av9Q9gvxSyax/KxglUvCDjtYDStw6r/r2wwORCpbieAlYbCDCs7Bk
Ef169oit4PbC1c0xz87teEa1R//9/8W2VxqyHqE0ag8fo8V+MB6UPGOIXdQ0XmXpMLx70QUziHyk
95mtuIZyl4ma6thoYSCT9lbm5LxbZxfFZrksG2ZDGit6Fd46UAVh9o/daM6S6tdvkoo1Cyp+bXRo
q8t2a0AARLQYu+k55LYDJLnPp3EMJwvQWuvsJxYIFGmINNL0P6jK9fNuYT3ItZnykZ920kzVdWYV
EWatjee0OiVbqweTQkc4QxEO7P4ub6q2NnAgZQ+sJoupgisv4TQLz1NA8MyTXToNcZda4iv/ERSf
hFU/r6oZh/lZO/DCBigwf1Dba9hmXr08K4RUr02FxXJCHW90JFZu9uqi6Bymlumeo2h3MHkR7qIX
f6IPK1JxixFjjlsj2nifm2xsxm0XNI4JFNG0bb9ZujBHz5v/agPKZ1phSQzQsKsCGIPcwHjpxpiW
IAPfG1q1V0g7T9gnTdVlBl90k7Jjs0TCuP7J+NTo6eZ7TKjiTzH7SoWQ2vBsLMdbLgqc5XJytWZX
gPz4xrgQXa3W0YqzYmziiB1kB4c9j+1XpbYFcExfSzE4mu6Bden3fwuVueFFaRZWqPMB0T1vNSn3
p3fTiM4rUT+p3FyD1Hl99JUkpFgRY3yW16XaBDzkY2ve0RrFlYmZuZv/qDSnqopQV7OT3pilgehj
pvnVFYPEnVEYpVZH7urD4losmzjE4cW9FRIF0qCG8DRXKakIr2Gq6ICEt4/CBNLxrmPVJdBPEork
Ueq16751/KTIUbYCYtHPLlftuWyU3Gpvgih7PIolLQc2BUi4lIuFjhqkgep/8iYu9xbbEz6t+3aW
8qcvpGBTPXN+7kTYMLWqh3NTte9wsZxF3sgJjWn+y4dkVU6o0RivrafT+MTtI+kg6bdsnliRUnQF
2Qw5Hz5xGNIJxM4EjRiL/o+ZkkQBIfXQAWbjApl78oMp//C4zLYUVW9v3SvW48se3zuseNfps7vQ
Zr56E6wBgWMCS4bgPh/aMHCt3NVv+xcNpiN6KL/36xGxcXIUzVGGjJVGiXx3y8ZUiFaad3XEAK4b
3439udsg33JHmXQ3bhetj60YETWrONg8Ts25c9LG7ZZNTnN/N4DLo6W1OD+2xKvDJ3Lf+ijau37Y
ui3SK7Vk1wWn/fsJEkRP+Bth1+frmd4sGWj3jfWgf5rgAZj+2NpftYpbp7rfghI7zwBENvrLwX0n
f5RAlsbcE3cAObU/VHFx+M4SQZojXycUWrIEg9DWfFX6Z2M/pGMhNvT4w7jOxz5UoK9nkbkZiewe
8ywwKVWrzeZdm/ISGSduSX6iWQ9QOGU2cv1KSy7QpQVmFjtcPcO/trWMU64QXJ2A5ePdiv5+msi8
z8h744fM6MzYACWpxKOGjzbfDt+bNaLKTjoIrrT/or6QxcAtIwss7nfZoqA/H2udftVaXsjdIQWf
XSpiu1frpvzrGQ7/dx2/7CrX20ROozac/+1lPcfk4Om0p1h3tDwqHHMc7VMkakAEgy/8PGyZDbNb
BM0dPM1G80fVLgEdC04t2Tv5y646uJVsHa5J0Ai8M8x2+p+csz3RdVordg2kKAVf9+dhn2FbAvaC
F0xPn3F7CFrr6MtxRCFmniTce+vtZF8hzyVoj8rb7zX9tW9sYClI/2ZKMri6UFOb95uLi2pKM6i5
n6nnzpDxGOnlzagwJiX6jhb2PS49IWY+EKWRS3PWUKDUt7Tbzjd92LnrnbN067IxBR7jOpRZdeTY
9j9HptBCSHSWx6OFb2Rl00X+sehPqfzzX7UTIVnN/QAvWEW4lHNH70bCN/bj14VRkeCDG97Pul2M
qc2jvTxoZhxrzJ9EmAUVS6tr2hKQ1ZowFqjBZQM6vzuSzM+aAUGZJUlaIj8Mo4y3pnhBt9OjoMP/
wzGKCvnBDqn37nAV41KUEfvwYsX4ZPrknzwsO0IOmJ3/wioHFs84fMYpJpQDohlB45sJv280bTCQ
CciOtznY54i6QHD1G2LDYJinarfKa9VpQCWoTObA+c7+D8H+0o80XHfhbN+1o8TIws8SFyrIdTAE
aNP88Pc2A2MrGHgeHoTrGCnxcOriblvtUrn9sUkX4e7Q7UBKs8yRMZE7muVwVHl4UTT70lVeb4VP
m0PyNCgAQRmv7vuj+ModpL+GpsQTJBUZsemyDA0C5HOgJ/GpsPEuNR9jgCwdFdQJ23lhB0Mc/Ql0
dTC4rjlqu43PvBKKoSG24BsxP5rHvAqAtBzRCIQV+WdVZz1juDATZe/DD+7MVM3ee2uH8b8wO3cG
RJ/3zsa2djeTGOP1c6uxdof9sTYD+fGmH/dKcFQ9rbhhmbYVbGPswfaaVULVZCiWojPLdZHGYJB6
kZEmIbg7b1GDTw8A8j3Fteb/pBsymf4iX3MfF3y4a3aKThi2RFqlkIvEiQI221gX/K64PKX6ks6x
yR9F/3MBH1eMN0GF55/X2G2VBmuYxSxrIF817tyG5F7qjUtoRGO1Rk3IVTRACo+Gej93YVmZhGNi
XRkXIcJ2qA6c/O4VR6NNXQvwbkON4aqmeNnGuHXIs8Yp1XcJJmCzHt48/a8rflSGxozDYyfzConz
JmRvgAJ7EkD1sqFRxJbrA8yOZZaleJnMQZPRUByalD8cj7GGYG0HaSC/oBEj7OFFDzUzZUjxFto5
c14HAUaGT4wCtnE9FKrg7itHEJGDPJDWaPJIuRWOM0xkjVGaMaNsADgbUlWBCdc0fo8WfhIh0xII
vO0SqeSM2Pt04MLoOIJAfZ6/FFRR+D/RyNxZk9LzZckBEcn5hIX7JjZUhFrW0ZpZPOHoO/BUn+zP
VqgQOtEKmUAe/+cSiAXCkfmRvg2Zp+oSjbL9zNg0dIGvWW3fYJMfXn60F47WUd1ZMRvzV9QiGZWM
70vLGV44vYAbnSHL8raG2rL7Wmgcb5WTu2GF0UvIVlMy4XqO7bd+nRl5wwSAs5DRDy2j/xGvY09w
w5orDuOArWE5dELsrCXwbo5JRj6M+eP0mHo30+cgM8AVME8ow4XBuAUiwOXh3Wc0JvHxDEJhEiZa
cUSgT+WTuTqcuvUEQm9GWLFb/XxuNPlt3al8UIFuv9uDRIIZi+gQOFQm3WwsoOt3Yno95v3Mn2/U
OSX2TklrmcAU/jJ3Si/nhjXr5w9OJfrvSIJ3Z8oelbKkDuTxyS/dhiSKPLuELmtLlH13mbwoLDTm
J5LeQ7UJz9/ETiwVuKTTl+eHAloB6Epew3n2WabNI0g021FRr7n5CJbpyKNYFBQwOfqURLG1IO3B
FIo8mZDu9uJbWOGv6pSvcuxWLWHIrpyzXjRFXa8HCinP5x6zf53qaFE4woG4rx3kbSCdGkLUcRdh
1vGSB8d9d6sxuxRuK8pNf5LzecCLMzx2EZ8nUCXVzM4Fh9EAyUhc+Qb4Gb02bAqXt2QNEXyoO6r1
hR+0MelV8WIIlr7kNeSOT9LLZoXlhbnKCfT/BZ62FvG2Mskk3FCts0krosydgepB/3uutZU2PF4V
lnoMxSiBZiihz71WJ/1FcDYwLB87HLTujQTl51yr6jTsujNOcw7lAW3IMy6L8XsdgHXUFs/KmtGw
yBVK0tiHTSsGVC2Qm4wgsdldXWDES2iqBU2o742wEx1TTUMT4qopEYb1BeWRr92rDQ5CVLr5gY/e
HLK8DRBkBiyEUbCvnFzyuj0xnY1Og7iWiGtrAcH9CzdloE2jvkSSC4Vtjf2kMONpaS/enFZHH4nP
2WuWFYMU1ehpfyIAN/89aH0lpZZ0DQlGhaeCBrJOdvnlug8Jwgek2a0uTJG7UVPP+jxQrhXOqEJ6
0kZgQYiDu/HONpFGzFaYDZflGLY0FVGXKq4ci1SeyKWxDuWjtsblMmVZxJN7NbZM4n5sljcOBrN9
AaU/9+wpysa8Rcj9DFvCJ/ddxR7W91bLze9zatOBflW+ASV6wWrO13h3jvK/F6LmBYetuTe9DmW8
KNgHc7+l4wUXc7O/204iAhBceCKtixeHrNGibMZEYXPqQZkQJcr4zulXlxrXyhkRaourNN227edP
+EejJy4/8HoDG9K4tMptPhl7WQNEFZhsMjUcKHmJaJQwV3EUwiXlOQHCkaMYGwyM7PvMQZdsJiAg
EPb1QWO14QMw+Rw6S4BY/aDA5Rm2sqNf9rEmsZz1bhKXBLN2IWVQ/dO9ULl6J2s+oBfZIvwI4dPL
7klfKZHvMWtn75zfIi3LnB3wFDckl9yPaqjHKYtGWkSLlPMcri3aA1oPnGB5CVSr6c4JErY/CvJ3
ddBd7LLfD3nMiDH1SCpsOi1clawMVGeNj1dpw1iXegmLlBC6cz1HM6j9YxbdsPm/ZPm/nNaPnBok
gOj1wJ7ut9A/gf9mYlgjk23JDMZWL9tLSXIwliCDhgfEj89pTc9nVBFJ8ybPeLDpnoLI/mni9TUV
hQDyEvQCxmS42eswd8kEA/fu6XztufSO/iZD8MFRD4YMPFS6XY9oWDNcfCJNYsPtuUc4agLfcv+u
JI+ehgyMDkNfgd/CS+Z3eFb7F46btijY1OZDU21CBoK5JsMndHnch6lNFRYtGI3vSqwFXd++GMUm
Rw0MetcBwNeJHeHQeAw9K/+asY4/w7hyQuJH6MXvla+dKb6l6zZ3vndhLs3b3qGWkORrZEf1EN9g
pHX6c0PNsh4Or31r47iDaYeAGCKUKHaXPiz3choNOI3dDK4G0hoGL+wT5ZmMoLGuba0JWruPkCPt
GJIZewiACZhivHEnz/satif29kFpJiFb/7/ymTdxe8atLbLSLwksiBIXIkZnljkDpMNN9y1odIpR
o9msP1iD00H2GTcFEExo2EG9CwL2CZg9v5MbekVzmMojbgo7RM5FjBoCRfUJYWtVdZF3K/FdtAG9
XGxTKwrB7FqfLoHL9HvB+YfwlWaE57U1rWLP+yu6bpLEs4k1DgGkEZ/5Sl4/VlP6b4R79ohOWg2X
jMjTg9s7yB6HGJ7PYwmWjH6trsWfcE5x0hwTc8npH2ZQ5S40eO6JEMXRT3XuvoTrlgSpRiF2uCGx
g72YM8PCEvlt/iovaDXB1kvPbB+lwx87m936o4indDdg4upjC97andAEk1kNN/xWGho2mlY23+UM
abSXeXtqiKK6U/ydLd1vawWN5sPVMWYQytljMDKYJozUO+2HzztH2psXEfrsUWkJW2F0PmrR79WK
/pS/NwwnrBmw8Av1c7uT+FrmU5/RQa0qItEwpqptN9vSHnhTH2KWJT+LeBE7bztSbxf+vN1VHKI3
smJkR4hiphexvyEwMUDe0LR2OcQYjZBXS07nTI91l3/pktYrPVjWOEqYuAdpaq3qyeMhylK3FPYn
q+6lYmm8Ek3IKRGOroRGyC+bbPuRWZFtpjSypHtIuxN2icaobow7BUZ69NxNFZHd3UyRgNx4X7fp
RuiIACy/Uj8HJ56g9vVdB2BApBWWnSAsvbnPdMZYjs6kK2x1CWwLKd9GvPfLh0c1hBm1ufdRiMil
NQoCTIBex3vAMx+vUMQwcT4z7zcyx1Rh9F/jIYAwbc1Krbf8Z0RA67oz9McaQ9qnASgjZWFWtxcs
2ntsdXzI2Iq+C9ht/WuKg2y/0avIz1f1/lAh6GfSVJN5CoRg82czGNq1fjz7bgbswX4L8xDyJI/9
tk6fgXChGySebOW4CCs47UciDy433YeqPnywguYW5rlDQLFh9jIuzgaLllDJp13+LqheadAIqRzv
lPgoLhmt1hJhifsWdCJtLE9PI8TXsCGbuzUv56cAlfse0eNHJBr0SkD9ZGhGrsbIELkOJeoQZ96E
ExXsgOqYDJGeY0vF61CMBI8IhO8v/dHIElZ1Cam/wODy+VKP7VxAp0ddXofKeupiXZUWz7I6x1Md
A4hTc9rKMXtPhuAseZAlW9XbztOmpSqrg03c99dO6LYz8i+qBJOtzy9ebZd1Cf7SoRYoUEU9P8oW
Pn9uV1WrqrGTZpC52RImRNVmLExptMa+Tq4kB8dZmP94syG9+3cmOEQv9WWv2224Wn2wEaG6jeQr
wzolNlnipcslCwXJJruzQfSRrd9EqIhihAwoyutyNZJh6zXZYiwGFEjuO7PAotM4Mfp+A+jC96Kj
+KpYYh0DFEj0XurfuOrBxCR+nqjGqcD8nJXG3PWv2VaDw+qIlpkWk6IacRFgr/RNYf0alvIFDnKb
bVQ42kuacC4EGthm1JXr4QJMhnedB7HwgQySIkfCQa+SR9h/On16b3RbwKhJ/83mhAtlJcnRvFxx
rFRePeUqL8Ho42GJz51jN4URxCj4x/D9QjUn5yXoqCX5Ud88x5TJVBNdIu9TlYcOz1wQJxvjkSO+
1RsVRi101sjRws00HSupebH/4QsDrGQ4CwtnaMJP0oROU09h9IJgHsE6K3maA1rK1GLadddL0Xrh
8jMAmHe3yeCxfhENXaq0JM5di9ygtSix287vBSO8j14Cw8yjqcw40KUkPi8IO8b3bDezh5jV+Usx
v23M6HWN4VcJQl8u3qEsa2WxKFNF+R00+82VvNFZE8RC3rxVZVmFltKKiZlJflOMk6xWJOjhTb9z
NI/CelaKsgJ6e4duK80mL7Mfv1GhhiCQOIwV7t65GN6w0IU1dTzJ2dQ5sVpBOOFJXqSQbviL9ywE
3Mf+JYEbY8TDulsDbqLsmVSwEKrWWPoYGtgwcVCNOqD2gCm5XsocxxQ0cKjhLAEDB9tJjy8nBzfC
5mbxBDFXqcTGiUeuegvWSG+yhXmkn7XMiMnl/aLhFnF3eBHB0L4rgRJNNNUHGAuuCaamfoyYPKyn
oeaD6z0Jj1ZLq0woqEY+TjAKRWoNomO5XXgFuf27p1bJSGRoRX4APZe+PQ8zpIH0j+8ppYFBmvV4
HW0xjHBxlCiTWhpq0XYX/bLpWWJxgtLc4WQHlnkiBwpVZa9yrJBm9zkOCErsQQ6XCMCoANFkzGJd
PWTmlwL/fjpxfYZq8KNRCLeL4nK4bpu3vGSY7xkXOEqpyX9N2vqL0IQSyzWMIn9JZjMvv3cT+fap
N5GsqceAHd9hZ7dOsbpHTRJSt23CrJbcPGp/dLr5DwelXGV4cyB7GnOP30g4V0QjA4fY3bhfiId0
I5TLFJnK+2pkZwk49NuerumaMnkaE3NMvY4rlHVEi8MNThe/GK1sjkzbrrnpPOwJQ7v/eGox5jD5
xTdStpNciBxbTfG1T+/jHABL/3APxbBoXQZnjIsWO9gDKQRBtoByPMayXmZTDfk0VoskJm2BiX51
FsFaykNmLbgwepbjE81HigfAMcqvMj2N8kvKQvhXmw1ffH81YxshCM/nkOoqR8z/shU/scL/w1NZ
NNuQkLK7sa7ezY9CiY3E3iIpdMVHBkGqNFbONT7S1PdM6UAHTu4vrLYPTDIBpd3a5T1CPDqR7RG0
wCf5SSE9VoIY83dnM7mLVRdwlBtG416IooNXcgRs+zNj5xj4MX4gAXK25uM898dLOKeoj2tT86SC
RZCa6b8ZeAyEKPKsxwutuqnpOX6YFkuW2/v7dMHxpAuy5JpxMxOvfgbEJN2IbTlWX7p9m7/PZjzJ
viWfzwHjt1j7zQm1J9t+Ofj2n47qqdlyTBwhzTkz9nC34NUIGNE8Brx0gkTtz3Pgs1RQjaVtSlLA
+at5us/qA9/xblYYblSZxh1Z0T1xm5p/OjpYgGqH9RSvtNIZk7OxnaEiGMIyFwZy0nsFIzd1mLHY
cIwNrCOlJLTKi36pMCPhZVgLUlJHPPilAnx2ne78Qz00IQ8BvggsGFtI6WbnOQPMrydNJTS69P8Z
q2WKDoHP9E1k1YXn9XAJqVt0dqKGP+3PjlpDNGvl9YntfYlP/9oDWjkJrjlk05+QKXPIdreZ+0jg
MHzC6RLIRErN81qyQ87Hu4nNbQWFqcUSB3mXj6LWFo/zzJq8HNN7SY155DO9RvtXsln2n1S17usG
hQTNUhAWyuY522vr5tyAq/HgnIMTpwButHAvhwkLHBnoeywcWdV/xn4gsCVZGtsEyI0WbGOr1Y28
DSU62SeYHoxHqJK2jHZaVW7ymSKe/kFpTeaQej747U8jPLW6x/QwjPPrHqmMxR65xn6lmxrQPDcH
uG7aaYzQPYZRrg7C5hjnH4cebrkq22PZldqiLH2Y4pvyDZsZwqbPQpNbL+UhIH0qsZk91SbUUnQ1
M/JJfFtrJU0SgX32ubetzyth07IYCU8xL/03YHPHpUA7xCrYIuqE1hVdpesuegXTqPCSyh7kv1t1
+vMMZO+tXJZYdHiBY/9PCLQVC0z5Ie0ftiOw37hRekrM540vW/VQghLbhxbZj1M+aiIXqrVhpGRO
hMzZC2bB7vB8RhsnBVeoTcyq0Rh6flhzQ2gNtkRvuC+lFGuABegRyhS00B6M4HS/iyu4/1WVtKc8
MgNfyqZpbiYcmbVmmGJjRR5cy+1nXmRGhKfA3lodMM9Dg6vHUOGbO77msscH8+lILgxeGQ6r4Y+S
x8RBqcxDlwVA7h/aJKssohAsBNiJYlg24AOhvSvhaLa52EPALehzAotQugJMXior9ot4qFj/xQsE
u4S4A0i4OOcJrJAellkKYcy/oEgpjwb/OIYtxJP2dGFsPBbWqmzFS4QYaqNnZgHXtJThyM07zkFu
AWPfAvDlXaulce8OVUyptagf2bfkjf9SJUQeAuyrjytxcJwlGjo+I9TapMDsQbPhyhH+Dd1BGIrn
AkB2DJBSdgVZUJp1pn6rCBRbgd4ofuq1Y/OgQlssypFR3dVR9o5C0q+Dl4DJOtlEYbCwVTP2Uz6m
efIDvh5adeYTBmhjq5C1CT7Sp/+aZ9MqZWUO7PVyB4gWc1vzFfB49EsYMxzANa6hbrUYrE5Em6eq
exHa61qr0Z9KGSPpMAnXH2/U/jDmIT2UNmrULNi2CrEYY51s21ubic4VkI7812LOKl8Q8fgVjeDJ
3COTlZe+JBnJVfvuKCoFiitWQKcwvg0C2oQ1FvSV9sLzMe9iC4PcZB+/3jOeOO43qp6ElHYIgPgh
vOywMSft/qbh7WeNIRnZVCve2KxfVTY+6zFfdVZk7tCAchOBpkZk7lKKVmKjkS8XG5vR8SnB57kQ
qiK+0WwAR5+cSNlXt6ymvD0AFxNWaMvdxqsPHMZQ34Gnm70MigLNm9++GjEfHfYUm3xGQycKt6dq
bNIMtwNleU1dubN0EVxqt4+brufsLS4B5jU5u4FaftNkqCkQgZnf6FQzbrfJaHG1OoBRK1hifZGi
fCY27tEr9CvhIkEH7AwX3FF8Ve6q3BbTu0qrzpFDvgoIptjXMWC5SGocx4KgPsVpG+3RE2ZS76jB
T1kVvb7sw2m2DyN2K+5lgEc93rTWTs59pm0mXjNoZ6KlZjurmmvHumdkareZ76cn0kXXNgTROT5l
iA3jj4c2+z9dHMYIbXV0eh6IacVuPfvzzJmAz943a1x70wnEfVLW2WxPBtY8k/jcqX9wGdReTu/C
APGMeqvSnPC+MOf2gJfslOT7MV6zIZE+ZBAZ3zdUceuiOFdM6AuaZwdxneVdrGZGoDFJTUSpJr9V
DJmoZQa874VJciqIqdgD2JcpLR6EypHWd3b86ZcjWdCgMuz7qT7cIiog+Pei94SoRUyqmMA2LBUM
w8H7Suy8rFB+7MKCtqrEpUSLYdiZW4wtN6CphnpgY6/UJy6ULl1jK+sOTAMPqwncru3LJECjWcPO
X66Odsxnh3KilrTea5mjnTp+UixCNoqRdNJTjpWSxdw7wd8ZdFXlQJox5ZinguBYnNoGayluP02L
YCnVt1MxvsODyjpMPoURc0DTsgrSzfikvPKwYcCtOYkh7aoB8YuATUbQIke+lwMOGA8XwGEUvQfL
5UwFTb9G60xzYN/gKkSX/GhIPYzLdZFFFA2Tps4jN9AmKmizZLV0SJYr5RJQh6/QMNN2vb4OS/m+
2z0TkoL9k5o9yxnrgulJO2taWTGCSiWu1TmoGz18ilxCYFY0Ut3B8vW9sxAZWne2cXT4MWVca83C
X4FTD4e/D6AKwTqavmYYi4DWfq+LZz7ZMTqaeJ2MTt0vOMO3XTNXVs6TWup2YC5UVnv8kLq4Nnmn
CG03TxxS1gXkVYuHLyJcE43KIPJc0a4U0sCEXtOeN7CTXq+HS7Ye/M/L5zK2nU69NhZ2lCoHJS9k
HGyFKXkoxqL1QtrGafc6OR1ypYadBU1AOXl34ybT5o9OGKA0SOUvdUNja+eKCRogrA5Fio2GOkQs
J3cvxmfLOE7yBqY3F/XTObq8TdBVNjq0AewKw8U2JKUt/aKwX4+eNjSthKU9GwLwbfriRjGyruNX
k3fHApFnOgne2rSdFJm9PYjnTswENIG7KY28pSxICKqhvJtnyU4InYRw3jXv0m2SffC7A0Lsp7mU
2RpnJAyyUkVRniN33HC3WoV08Jw3NBFPmFl/hmWFfWAI+5/763UzUghaaho5lo3ycWSH6ItPk71e
DHQwCVby/Q93dMdGy6xwEADwfTWqJlGDyGP4rN2jK12IwmKnPZjsUN4dHCqSEldGEcWz516MeYQ6
gJ9i2vLkp9hChOR1c36Sh4phXXlfoh8OC/i5ip5IAt7As9+AMAtgphEr3u+oyA0ciYM2cEk6r2ew
e04xJk37rRkSCcRgMn2BUQELwGO5LieLrNA4fz3P1k8kZ6u1/T7j9shJ4wb/ScyC3i9ZRopQfCU1
8cvgfD+P2VFG03bHoqAaNklJlbylzUt0Im3HDzrPcdIEtmk92Y3bspzC121rFon15M+YLujtxY2w
e+U6LQfarQvYjFdASEtVyfJe4TCHLSLq0GLGuzV1EeJia0/RkkEWOQ6TKB89Ym79HRUAw4e4ZYvz
IFO+sTHAddD8Wx0m4EB2W8cLmrLGvTp6WIruIjWMULxM2QfNqUgnnXvtfJd572AkszVDFZfjwESQ
7XYJCOqFYDWwgcCLF83AkLILP0KrNBeT+cNp17hqB4fklfC/XchN8vClcO4pdyy0TLS+EQD8qhe+
WmQQ9lChjxqCA6WssTIU0do4anrmvLcTJeEJkuUiEwvpXG2ImDvrMEz3BSfQL5arFOJaYQ3WJnf2
Vsvomv+ENjU1sAiRBg6N47btaWsjNvCSRQ4AjKW5EtwrGGbQOf56RX0T4PUiIOEYtcGEQp62NUg4
7MGexvRVkNgT4wITD6nfTgQdKNS/vlj4aWzbxLYHLaB9NSs3nV9F6OW981DUXJVUEeKyuR4TqxmV
68cBR0Q5wmNMZqjXkl1+xYmJ1cCRjsxMZ7eaO+z3S0cCxy1qgXMa/lnGhdXNA6hJVPj4hduDAKtS
MiaZ1NChNzakJySKJocj5C6K7X/cryhV60Gqjm84eheDOG5407ojWPwKlSegjs3t60MOtZe9eWoI
LUyHoLmvWMOEuWhEjI3t+rAdsSofYM+H2Rx/Muqx/jgmLXqXpAwoGNZgCYJgCCE4zk0Jdv2l0vXd
yyUfaTal10Vc2mZ1g/zZ8qI8mBdMhzLNJVO8aWZdPDqHhbMpv1xKkdSlrtix/FRkgw1RkX8JDAU1
Xwp8YWMbu5xBpB8V83Iiykcg5I3stw6QceDKicYRPrnGdA7/XLGwiMfC1HnYrQ0IvlBrIXvLGDl0
hKEUb2hSypfSUnQbDFI6zfmhZ/9/uVsJ3+t+EF/XwQ2zERK5hqrxLWzcqtRWIQrseV8L2Cu4/IkY
KzH2hJ7w/P4lJD5gpVzMLi5toWoTaniqrvL+8rToTytHD7UqwBt2aVRGwGuUJsCRQcppPpZ/hv/F
lXBxuQ23Ju0lfGdg/jl/V/dFTkW2F+DLlFY6Rw57oZWmPlTL2CXLg3OtYOhgStuNhhh22EZDGdLz
dmwCjZ3AxL+9ewN3XFfcGiUmKGbyx5oI2BmanGUODCnjGfha9luRZw4wOx08k5yaPS8LXmUyB9I0
vRZC/yT9kOG2/Sa34dINLg5TAWjYXX5yFgUe0/WjQstlHdZGqYyshFguJGMWtYdr7NSDmic2mq0N
hnBCBiNR2LLAqpfUniKtME63/ZH0pfLoQ6/S8rT8YGHIR2Iukwzhch/AUK4fD+2ABViPh2cDaeQN
dAGaRiA4TYm/f2PhRsqT1Yp51FcLEMBjgRtVror7tLWFPx6ON1bHwA4gRVId1adqOQeu8vWBCfEo
wslotM30YEVH8rsx1sj8soSLEBMx+DSy/CvHsG086T094RFoQiZpwsDCrSBnKWpHQSz6GKKgFtsW
f/hN70q0HeRZzY8HhCaZYH3UdK1P8ghkFMP+uHHRBukiNSNUE3BdkXv915HdvK+fAzJXA7w870Hq
yd+h6DAJb+7u8F9UYA24wukih6ppPivxD4GnF/55StTKhOQwcr99lYW2iln3J96F1jrg91Z+adAv
bBU3BJcdFxP6OPh97vjbvISUmBibwtviJ9vIQmfTW2mPRPRJms/IuYzbB0foJ2wqYid0ANRZ8n8d
BTcrZto8FCY6w2sYlsXMPk6UiEWoOaPxjiCPCNjMC42mo1J55/2CiPJLS+3mbHiPUcVU94puFkV6
8y98hEjk/dMoRwQUhvVQeVS10Ve3nR9ylJMGOy2nn6J6xydlPW1rWqgFBNkZk1F1oQFfjuQYHJnX
7Fuf7JNNUVb6zSngLw/ieS1xGyYnYxyGwiuH5ssTPgw92TdwNjxpAXuLD6LZ8kRLlgrkfwbXon5N
ssSUJj0OmJQy/TQIOARLL5CTKwp87tQvL+mqvk7ZjKprUftXBWq6jHRVBZngARuYBDcaEXz5tRsJ
BKEgjJ+LUxZURv3KA/Y097xo+J4EmQ9w70TZuMdBtNUtigDPPy/2vxPWJug+/lNkLIxEwsd02iOi
lTyPkB6YzfsN6QSAScZaVJRQsnGj21+MtJMW2K/tQnkQvocXecAsUMbcUakIR9v0/TuybaJ3Ji9k
Xs8SavZQ1pKL6zBEaTlfBm4pfWu0TpuCqkOdiC3yk+lbSPP6L/pHChSf8Pg0808bHgHKegRPp6lC
dgZ82P3emK2uC7ZvFya2w3PURvZvudmo1/T6VtkXlIKf47B6bGyn2YHcJGfprmhGJLxJA32lTxSe
Y0B4EyJyBrCnrAHgC+fiPySe9Bn7S6vqTRa9lVMNDMOhmVF1vf/UUmPiWbVsK96YGYx2h1lUZs6v
20bV37tKO90qpFvMlrVUbnG715H4UOClLziig6ZRs0EfMC/B9AN6KGSPR4hKg274FnHGWK1HyzZ8
ruEhqxr12CgJ3KZUgGkA0TZqhVQRpQAGjlOelEDb/3Txm3lO33Pmk6PTL/7P+SjzFgeJiz5rCbar
gTj7AXZrBEgM3vl3rdjs7oG0qC6sygnHkot31XDHBzWZtwpVACaYcVTE7P1hz0LqKHyE/4fy6n8N
iRYpjPGNI3Jla3xUMAKOdDLtJgBYwCrbkxp+67yIUc/q3mXISzyPanmtJDWIU6n8B2pOEjkajDBt
ASRaDZ7nqWcp3sSRiEQrSQTYi7RhTu4aQdOGZ5e8w8RgCZCXXQKbtaYgPtG5mcIfWYyQCl+15BqZ
7WQcSSNAcUE1Fw3O0O3g7eHEADQed/34QAAuCT8Nxk4+CxNKlL4VqU2mrviCOvKSHSMJqQsbqqyi
lMuOHNvLo1XpHD3aZdMdyhtiBiu5D0W9wl1KfHj718II4FQ3h4Uy3u3cKIwUAeOgq9BZp7dkg+Ef
opGWkJQjPoJqUve2Ymft4bIARM6tkIW5cXYTnZapvBccJnmGIOYpPybP+NvPvnHhIcQZ5JYeOfW5
PzeuqW5yQ58DcDXesuwWsEQaFNhvNYWAzqwdQEMkcT9DaNRqTitndOsnMzJgTkwK2wonyHPTF9F8
KEk5OEOLNDfPRdWXxhR7IgkKVj/j6vzieH7LP8NvphHr76FT4Mwg5Ak8BjOt4aRMMcoaoqRuWqhF
3p4n/xc0hy52kRGdNfs3UovKrwJTW416DCH4tIyzLOBtPF+Si3cdZ0zeg6uWSX0hHzV4D/drO8S2
izt5GiEpcFQRgFPGSpgIKwmiOqUHidh8o3N/ijBXFWkGwiTStjOtLSJ/3vKc2ymyx7sHQimo8jla
epo5/HMYaS7lfW0kfkxVht5zW+4bFBIetriYQyWyl211xN0CyuMb6jgZTmGWV3nLtahC/O0y1axj
6CSJ99QJr1VG9tWKMGRbdJ23LaEyVZPtwFtWd++vo+NZjkEJcUOSj3lWaIrAIvEQ7nLftPWLal5+
FAx4P/s6V0SrWUl56QWBBJ++4qQIv2KPvyCfO7HIuqDkqOMaFpTZg0rx2iECJUBhH8QauqASH9XJ
RNIYA5g38hwnX9+dri5sXWzTJAMzn3ZTgY5zXOWVdbN4kgMLJ/1gh3QmqqqeNjubM8AzDg2oEgCJ
Qy0DhJRxBQPeNlxUb58cjTCcDnm1oEcPYA4UFqTnBfOPfhNYcY7X5pDSlygDSC0W4pfDpMBaxORI
IWM0BrvnZTsSis/w1E1u5LoGWiK8jW7dqnsqF9S1xm+D6ixTILrIHhDUVAAEdW+9MUdQL/sQNBk6
42PvwEMp2nLEwQX/CuwNKCmZkXcbcJ1ghD7WNQDscdFU09yJe4f86K4HCsEr1NJCF7ZoCsf95/Yl
1tY2BPEv8lFRl1ca7igClcOD+yKQj/J35TVErP0MPoHRhTSNGwXAgNZEj7svD7rmySlQkAFLs/i6
+kIjABtrnaPErRXZQPBAxmqCGDrv9OjBXxmf5XugMsKnRIaWo/fZQVHjzPQTCdFPO0+ailc4F0OE
etvRAQ2HPF9Zwm/GmMQEey2o+e8yX+VnpEJMZMzca/CPIO9eyoSMJK6DsmzfG0F/4lljD3dZoNZX
EIT7YkCioR6DcHiQKhUy2kKuT90fr6alpsYV2GQQhUe4iS1jbHzWlGJxbf7beAUDOLy0irIZWPU/
ebaVvKDKdcNgCBqPjDeH72YIExAlNzUTE647EBeMu5zsnobGQgZOr3wZA26EIMtnkVBb7kgKZsdJ
83P6fge2+Ncup7YuHi7mmzBWycd3BnCyaxv10AOmP4bM8k4O9psMpEM4wb3tsF1tla40/rPXNjm1
Pv0wEkPEjBs8JInz06XzgyvPP3MLbfM1VZZvuyTsF7+ADSJPOITW/6dYcZZzd+Sh/vlOFwU2vvKx
JjgSvM1TVMr2v4NB2KSRfbse3Jr6l/LXxsqPhMi3VhIWQ6yyqdo+mtfWNcC0/hDDNUPHo0ki1a+O
bVyZyZNWATVSoUF5lQsNX+LKvlBfv5iUkBDYOLd1lzJAkImzFPU8quYvU9tFMSM1fvoE4Cc3aKnR
O6+0ulx6NYttdPnN2vhnA97xZYr5KCk5BvwDC3/MvAFZkvTylGf6ggL2DtA7VrYwf46Ex3MxiY8d
CDH69w32FsM8+Q0M/PdGGs0hKZiWlHfCQT3sdNJoOi5LFjWSMyWWrGgRYRFjd0IDGhCwDmUmm00I
5M4VwMYLGGiI/MW6ZNkhM4y/vX6u8z6OmWrWbigMrHR2tLzlKH43MbyH6NEJAM/YO+OcMobx0Heq
OyCSf6RqN/44EILN0S2++Po5/a/19pjSS3InGBkDQYQgyAGOUtdhoCoKWU56fsltu0rnKOO7/4DO
nj0aEfGEVO8A7MdVURrxCNUBhIEmifFJwnZf1SRTHrNQxn4MO+PvSTvStXp7oXgD0HP1EpZrpszO
vU3Mer8OPbnx2v1fssOtU3Mp2AAA1+/mxRCaPzO8537iFaP97dLsKGA99AVU9r/ZrDWXp68XAtf+
U390k7Y42C8OXIk5xvaQyUqNIlIX0RDIw659saYYocYrgm421BTVowiema11WSDC9Sx6wcRGXwBD
Cgxg/emePa4jElPxG5nPwQVjJ5RChI4rC4us2a2XKgIbZdYtrct2luI+Flxc1ckqPRKPT5vMGGeO
RjnZ8/5vbUnk0g75SQveedTe/ZgOf1ecWF/jOiczK+GF1yrYhdk8exKLx/4HtsvQ0LlwYjle/T5c
//xa1CToj1ViKq2mNhpmzHBBQJx/XZgipWUiy86lBNnp9UJ5wbjeRj0QzNuVYxMzyZImkxYQzY+V
G72Wq7+G8opn8KF6Rus6zXuuDXSXeI/9WE74ik9LBdc9P9G+XBDjJtShP4TlmZCCEQOkmjrPIKJx
+SeOTV20oIpA8ivny6tLpMUfIGopz4DfPnnVaj2QUm5PLNHHYTj3nx/WGE03fRE+ejp7HAFUTWq+
SFEZtYhzeOtR78Vr9xSU1BJNPG6z1axhKMMjRaKQBooRszim/vGXMyrMtlQn+WzeHlnRBETxF7Es
JyY4PmFnmj3updafd/lvjLhcXowBeMb0zscLrNG8WeDkC/y//gzyRkxM+oGL3PcIHzZ2jmJUSzvt
kPsyT4npzUmP3Puvhb7E9pcoFoUueLbw08tgNQaGSm9YYzJJysmNbHaZfXWBlq7DEaHpEyjLsp/d
/GM5GUQ74/azu97WQ63W+R5L8vOzAE34H7Evb2IaOdVU9t3aD4W+OyIggLJZR7xnXKP+InwUfSZC
oWH598L2k+DWpc71al+BDObhzwByQ0cq/MWQzdbW0hBRAiLb66yb1cmu3RCtoy9G89xySGj5YxYM
gedYMR2Td7VBS+68rp3z//xPpo57ujyh+ub93NDoByc7pdY6pQyNcMSW1dVNM6huOvFAZp9z8/NF
NUBdGhZKbOqCvHEXcOO3uRyOdjpakjXMORgTQWLFby1ru7HMb2RpkMH43wL1t3O4WaGOH/DWUoTy
W/D+li4ARCX1iKyn5njqJdI42UgJ6wQMc5vvEWVEIUtaDTCthryGPt0nSTx63naHqEVs/BPDoPul
Q3HJvhgN1rsomva+COQbWrZCDQwyCTEkcUDVmH8TR1XjKCFrOQ/GNotf6AqqEKOL6ii+I9SNn7uU
tNeXyyk4WZ36qr1fGk8oKfI8iVkGD1zxNBCCm9ZBI/nfDMr9e1NgqkottdWZ1foTqMdJ2nJz7Wy7
7EC2r3kXnkAwQcXTuOYlGeO+S8oszCtA8UfsLvYfMRCOJ/INXmupkvYz8PQK9q1vRueVPHFphblV
nkPrC7cgsdu+TAi9qyE/efIxq/n6eYV/addn62pXi85nTbETjMwb7aXw5wdkP47hBp1GQFuuZFqz
62HbStjRSTHZ2AYan5Lnu37oI+rxvQr73re4Tpi7WmZ/UKBzdCtg8kQteScYZI14FPH6JadAsjBC
obwYf13ZVZMATCM7r39mKGQrbg+Xa+JljlAUdkDc/Du5wccSDHN28JttUAUpyNyXkv//Yhq4DS+0
QiU8bySGlHkQuoO0KxwK3w1zjP1K2vH1AVdGkrpgaH+IyUhQmA4YRwr1HaI93yxu/9rq1UDEMNl4
kreufvW9Yja5pOVj0EC867mM6KBHFOucQRVM8aU99CTXuONckWywGYX3nDDjBoIvxvdsN+wkJOG7
4i/hcWe9kfMW6+MRQmwIaBSAFyLQL2KT10JU1amPsWUS4P+Pg5mzR5k+HFCJz0aB/zyqkmUsjtAz
9+NVAjLNX7ZKVOP28j0vdUi23t6FeLhip2M3RpNrUloDFdhHH1pOoty79AoE81T1VFyd6FNvufwt
In1h6RU/3Pll6HZsqOs97K4rWfYM7U+i7zuQ1vXndZNGMvyqDCzJa1ucdFlF4d3DNofIsKZ6Y3bh
VI2AFFP62yO8AAOweOlqQDAV08iCm4JDy3eqZPKcWqVNAQRKMPYC7lJzqNw104rB8LrV/No+7XJv
XvqYFPaV4QpEmNqGxNhcSxDBX8h0Mdeu1vl24C1SCv0h0Kh2iUlPEcNjMY9Wt58evrKD7htTzzDF
vBBAj0meT0U92e7ebeyoGZ/Jb0DGWUEyQVdyXQmGTgD/CSSpDP/BaOBCIROsNUB6O2Ey4H8uU845
rMxUIl2dioAAHnWqXjbkpSL04SRbmMPBgm73jvL0dHZ20r9xNtICQmtS/so0lw34Ax/l+LupEavr
Gov+DrHS3GgwBvAV/jykgHKEKG6nfzmmMVBV+mxeujRYsiBat2qfMHT/czA78vJrdCkCAjXEwtLT
OfDvYRCKEOJfQt6aL8r4dDgvcr4dix8D4JxTlOtZMXRgNgT/G0BjYiaP/gtWHbhf4XTZmlvK141J
BPbRSRBB26PwMkzCHKXzEnNn5RxXJJA3GYva4sEVkXv3L+J8/1ExLQJlBHJKYhZjcvElhbOk1YwS
B5DKKR0DzBPgBPq6PR9JIKUgIk+Ge8H7pq9HY+SF1J8xNrtv+MBnGI22IpXeRdCItv2vzv5BBtAl
A95uX+iFv3UMUQTVR9EH/6vAZUlmHH+2WObBekNsZNW1ZR3hiEr5C+jWR7FgXtvr/RqDI18Au1ZJ
TWKoo9o+RdJluTWqbBIx2w4SYYLCh/GFVTqu0tdhari97nAdIbIQFC8JkRIDzH2GJOXXgxwvDfbN
TTBqb7zq9G3ZiK+hvGo9fFzuzbMynBVMrpxz5A5OPHsI1Nc2BFjupGdzjYIBwJ7bMERuwWtCQ7xq
2pSTm9QQCyGvvB61jOOJLlU8WEutJBXzRWW8BuAcSYTpKe9vpSI0axi9WJEmKHvdi7rbi23aXxSV
ryQsRFmnwQcdt9G9E3fkRiPfRbqpRMEQGQWOVHHAtoudt9U60i2riTXR/+jeKOkgFnN3Fmnck/xn
iOqUZHFQvXnJH7inn8CJoXcmZLgzW8nejQ23V4Aq808ZEXUyda/n41Qaiw8N1LJYHfGDSIIntpGX
181ibU3+Ow+R7Nj+2i6RVHBDaaS5BwGAHXicvDFAk4g6XGXexOMV1cHigMWccfwV1p/oW+UJefFm
SzklhG6Yo/Cv6C+5hpbQjEF1AngIaKLXcGdq3YWRA9LHgpSBXKh9IamY/Vgl1eicc6sAHUx2Fadf
lJMgd/KAMcZhZ9r8GkX1TXcTfqC5HNk44IZCpnsR3r9qlyZqcbcVttjTvJphdZiCXxYptrwoptin
/2eNM9MSUgbGbzkiQBT/FW8P9AxJmn+Ummt80JWVFfcOUEd44ECMBPeh2/44cw/27BpHX3VidUB7
/IQscp/7C8ccydaK6WxUwYPmtgYsFXW/oh/qckrVnt4+CN6mZbayQtB3hg6NdbcTxVB1M0IhL6Eq
Grov28dBBsC8FaUBGlHjafHQJRSRXD+NcEjevy7lub3s109jZeyBAkY1P4lc+KCUzNGG2hKuiM/S
iJIgD1IiqF3MzR31JlFuKrVgh24rNc0ZUw5D2tN/EwbnGjaod1VsOzrw5p+ib/YEbMnVSI2jFyMc
ChX4l1XNpUNq506bQtSZpqKt35RRm3pI8Gj6p2se2dYQ13y34PGA/Y3e633A6M8VldVCg5UDgeKY
5qxw30rU8VFvFspbFgAxV+P3g4P45LfgmYl00K9gnY0pxXrN+POItmMeiW/TPGq6S7Dgko8T9x8p
iijV3cf23M3WZP/yAVypxG8YO5/ZkFs3wDOZkZqGKrrsrVdSLAhJEGALwWv6NVbMZ5yu2uFaLOqs
Pv2bWVbA0EFJY2zuJMs9HUUNVP85IglXay8L3Q53ETOxk4mFiEux48tAnwxf1DGeY307KLSGK7Hg
v5tEnmvZKq4r+SputD16otjQ0SvK4CIXTdk59vQzwV27PyuEWQli9f6ApRk5m3ohN6UH2hUpqX/T
4xsbdFfYY8m6RlyRL7o8v1kV2vdrN4T7rHVxi+pyLUov1PVQJKsPeZlVJn2K6Q59jzUIW4EKAmW7
cXhdhz0wetXf74+a83U3aR2oWl5rDWRqkrtQLX+u1OxhoUGy9YzXgaigigyEugVJEDoicm4uxFnL
6Hq2ftDFNNGr9BCmjFpJI907TUDJLgMOcTLQVLx7rdtb2H8LeYe9VMwMHuD6gIIhrklGBHLSWMZU
sllIMLpKJ3SU9/m7i4ZWezoAM+HFIaOn1zJd47eE3//ApJcx2dPjUwqDoOynJLDrWVZgIwId34Ch
V64Ykpcz8/PLTub7EgWTp0PyJBZv0yBXnJ+qLCyH/KEavW7QXXdVT1oivsnUH88SgWj2Z4xiHjjp
pO/ZV2aFI1T0I3NozAlAf223NewNBe7FFbsjISvn9p7ff/VR13QspiJXDub2tKpyAZl6NhjJy4h3
xdQMkfed3xWTTV3+9JI6QrypaO71v3ruwCo3sEsdiMl3MTz5xp5leBYL+bgCeX88z8cNZdsy7CzE
UjPM57Pxtzht/7poOzn6YU6y3Vtwxq4ns+x1U4BrmehHwTyyIo4tfQbWqqwAE0N4sRAF3SgJXbl9
hSwPpTo3UH14BVSIQIviV3q6DhJQxNx7iiDv8TrCNByhSs30TBakUyCnoQuZqpNL7C0M70Jkjv9u
KtEgugRSQte1kPHHKE+7RCXyu0gqc7hCcs4a6k0Lc2Irvcz1wt0nYTLtKF9PR9Bmk7Lr+DWdVx0G
f/BRdy3MnHqnTPzuRXPteagC9QRWR1jAU2lqKzBesHhdmCLZESwi7uh97llXPrzV/lfvJlXchyVj
WEc9I1wcOOwxvP+i9zI65nz0rWgreGt9wcA02SYFn4PFF0hZRM1H0O7il54152G48LabGVaNEzZT
Y/wi4dTwZIxEzgxFKh5oE+GB5diOqEArrni9Xii3pguuAd1tYssGbeB+A7Cn2XklkyXmZVe2365k
1tSBaGYAEr2hTAEzeRHbuuOYHroNV0LqhvbueQ6axTwcsC3HMsP9CbWtTlCOYNjlwr8Elnq7bWs1
kNzkM6iOH+Svox17oolPy51Ty+asyk/j5HMXDxnSr271cn7YzTnvYqjkQKnp7LdKFmI+9yCzMw+c
UhpRMbaOQs9gN/Sv+2kwbrtMxsuqkmod4uPcs9x22PLtDCnKL57QJfDkroOdttrhVH9tG1Og2Uh0
zP0CmqUljgBB7EWvbTkGJt2Z5ypEYlRPN2qNQOnVtzYZcR/QV4w2xarkASEdWbZ+VaWeES66qruc
IxB9+PvM4S6CDPMFDkCe+UEUzqUIksSIesINFjq36rZrfeF3iWfHHcPsGmT4Ue9BkGSFy6oDgriv
/GjktNd4NPoKwQaAD/M3ULt0G0nkp9I2C1FBZ4EFQw1hn6zcaFRbZXndWe31eeWEdm3bZS1KYL2P
K4z13DyKkt7aHy2v5YLkZvO/sghRb16mtCVcT/2jcg7BJavVhqfFjWcG7WPYLTzRWYrGpBnm9iPZ
dlGJnT0D+Z+BwQ6QB+PPGXlb3cxHGxIgVB5xCmp6ylom4WORVf78Er+oJDdQ609ozRLQwvDrpvtq
SfcSWdj0Ypgg964elYCnhusUsfJJ+Zkq5EPi+vl0Fo6aLNrP8D6tViGm8+KHP8U9el/g9STl6dUS
SBeHfV4pg7EXXdh9POhrYzQOQ67pxhbQycXAXSwAvaFT/kY1iRnS6IRstPb6FlncfhHU/fwfR4gu
o9OxfJs3d2bU2iQXvmN33FYgifBdls+J9ZNLlOewHM41xlUtPHJsz37mYHBL0Y6loPw0ru+2Tzf+
stRXjvOEEbvvXKIN6SbA5A+5DAHaaa8htY2YvQ73xvqQOdbn1YfbxZabiJo+m48ox66bg8NBvVh9
ffaQOKA7iIfV7LTOHTb27ciigMJwE9/WeYpLIQXc11B5N9VMTBLUWnZJ95iegfjRlgcQzJLjyuUY
bHvOfnSGAspBLql+SmSIEqPt0jbiMN4qtZb0LqFY27fWQ0ZIMoQ24Yc21mzywu+wamIzoC0b5vsu
13CTKobWZlsBD+aub3O5EvZVwkhXUU2brFoXzCYBx3a1MobU2mCrtKzjwMsta6bQc9j8CYQGO1XO
xZuP+f18txlrR502LQ2o06ovA0DryicoREIJRzK9GlPUiysM4aizdL5pK1/u5D0g7tWefvdnauP7
mEwcBUHmHV0rcYpQgW74yPo35v5+TeG0rYDyoRHGCt6ZCq29CdiNI4ViG08b7vM9alx6EljiQS4S
wBbNyusApPbkQV2h5XE1t+hmSRVZjvBxk7LJ5h5kgD9ZRLhz1jx2jHtqYS61uV/9PFTLCtBDdrRH
K2X9zVVmdM2+Ky3Y7l7po64coiPXR1ovVxMoG8scfqO+mvKFfy8kto0xKTMF/BFs9wFIpxwo/dnd
79IAgAOXyiw7G72NPsYkygUKd2m4bM9VFpvYITUQb27rS5/uLjkczD0xxbhnE4ool+CvuJ5pC32u
Q4aD3By2GKtlM/608rDNPBt1sMGKOL1jSAfib9cr8sAkhEh4TC8Ds7Z0wbPSVUlHglNCWewRakwy
yiq+Z2ti7irG4HnPNivYWPR9IWGKkLSuA2VVPiMksvs3P5EIhDKmLYmHblCa7xWIeZtuDn95VzvV
ywm6PNQVbTWIZrDte6JGgOn72J6ztGKRpQIi1aiJlHLvgF+gsp6O4SaUlxlK0M9yFVr03Ih5+VHR
rfxYLZxe9lafvdWhTBf2SyTmd81jIMhlrfRSuChJuTiQi4HP8WkWfGimZmKUmohfCBsLWuvhkky7
wBLYOCARBKCMSCMY7UQyzmd9Wd7Sx30+XdgiE3NEQn5tU38ceJh+Cv52ApHVJrGuYPc4NB9ZNEYM
mTfFQbYuiB8/XTHrhgZvvr4zouRGQCwsr8LTB1tz2d/k9dp0EUeRfM4Y1+Ukn9QnpAe0mca2Kl9t
zUqNQCIrsOXxHemGEhl/L2ARVk1MMyYxzKPdflQWE9zEVyP7N51siepnNK6nUeXsrmx21uR1vL3H
UNKdND8va4D6DXdHpVmz4EWNd4E21G1ECTgALwSDsuB/MIBxK5Bvrbkb/s6W+zQwI33q59TMB21B
wjFP2NOCtJBt7gptUTWSvJmmMdANdZBfNP+J7upC/fChbk7xegH7kBAzTq8rBqhQb421Xt4NmgEC
Sfw6rVJ2+6V9syY14ALrIaSz0ByI0j/1CMbwnH0HljSN4sIE3qX5h/pCmwTLLgbtLlrYL+5fK9Q7
yyF7gsUtquqG+J7s+8GI57VUgipinZwRchHcMOzPGd0wuB7I4m3cCxlRqMqyZLD+yH8B7Whk8axP
TPpPFPF4d3qx3FYTohX8YuLDXU2n2EGtwhLuzhUNUhbdJm+stPlr6qOa6N8QlUoYqCwF1czegt79
PMD/SQtka/FfXVB1qBvyrhcKpxLoctgQYPzXB+de9fhD+LLBAEpN8Rh5SkXcFrwQI5cH3NDj+7gS
mqf+eE1rQ4UyDfXQIfP3v2pwAte9wIvWmGqeuT0R0MKG0uHsbPQAcw9PX7HPaHRG47kZ2AAfHWRW
OuHf5zw7vhjEaAp0giUkwcPTu5Lh6fuKMHquhkHgFDAsbavFLucj1qelcUpDXsZiPC9ugKxO3/Ad
kU3Snbig73gn85LG/fmFtJ500+NsPSaAu1Tg9ht6QraB2zbW5BY6E7tjRWfnkt1HGHNVktjxVO0e
GebSzBie+tzUlo4407n0YhG0xUdLRjHLPes/CQ4JJtziCJ7H+VZRQFNMhdGxBSiK5MwOabQmlvdu
20IbsDqbhpGPHfzS8kHlmD6289TcBZapLXZUR/EweZ2YU9C2wqRhvNtVwlyraPqyAuMNi/dMuyHJ
pUO3Z3gC7N+CgLQDNhSR783NNXIkSz4kxMnjWswRQAw+DJ9z0Yl+Dr/iw2jviqWJAf4sIF9ftGLh
SlMVoJmB+EbJEM9SCRVxmlHa9pEaqkQZF3TS22DU3muuVi41P7TWT0hbXHvvS8Nw+Mgtlzwrevuq
37gdk8Cer1+BJNIFQhNvNJ0cfsAepeMG/vp1qXmKXjaH2Zt4YZhA53D8zuGIUqv5N2W2e0v+jzdW
J0grvgZBgP/B1zGoCxEUEnUgEmJdwJ1v3od78TtyIYEk6D2ZDyXUJwYlkbVMsRf95nMkInSG2QI6
YinxcZZPjEsroRpCT0CBYxG20PA0gfm+k2/uJRpC6Fdd6D4dmfJw1w0SiEVcbGU/pWpqQNBFMWEm
8WKQZh6WQY5pv5cFh9HKMwCP2sjC0BeLdU0r8XK0B0VEbOVmfDHuzEnEgi+QReThJ2jrwubl6gEJ
ymH2gDfPP5G4JnzV0Eyidcr9i3Ulv3MNBDfMguhEVyObxNyC6SrgigEln5bp+d+1CB91/yM2sGvM
WtmIslWZUdFfWWylz0x5rQ1GgLoj5z+DhC5CrjMGcINoCE6MucofS3ASaSgsONSk9N1p10aaVhOy
siEZDuSTAmEO+PwztKXkn5Mg25iSlx7IDFma0e8Igh1FemxSzQyUQSF3bAtnUtxKgAcesFK8+gqI
jONkxIB/WuBvZ41jP8MfDpFsA1fQrhazqxRLzvL5d4jsEvQ6/DATY3KlwoFWdWX4oQ+F81tjv4NL
2wClaCIF/G69my15P5gWjZREe9RQw/yiqtelMSH+CrmNUI1cafMRRLfGtBBqQiOX1pr5+3BLymNl
3PDaeEo+PGl/xLKaLRcaiIHxMZGIx1HazAS+ffg/ta4T6VOGyBwC2v4NPgDCI3Pvr0tQ3xHjQ7lb
tzIHph1sYibZ54BMZXlPpwqV11T+u26OHIDo3DAI6yLcl9WNLY+2v8pFdCdgM0GrGbBr1Qd6ii6p
4G/ZvoyHSGLXXKMp5R7y8UrJ0Qzwb6DaB6kUDd4SLdZuu66tF9ng1ghbWwZ4vDA4ZneqEuptaa5U
ERDMGktxcFWWFQZOklBA2/lXpfVg01Jg5mL2piYDxDGCxriowe1NSwyG6CqO3TD0oiwS77NZPy+D
1WAC6BrmBk/XyZcQBqW8QQ8mreKlVJm5jtAnqjg0fB7oXKvPRM1IOXKGqdu/M7ERwg3ryYnwWJXn
z4ekxVmxvri2UCCcrYtwQETkTVOC6sBVqPzNrKzMuRWJ1WaTihXmMWTm3llccYc6uDnVA0gt5qv2
bi6NrLt+o1iTzkJYpsCPZjKs8CcQ+yPeUOQZmEf8TjvQ4+xAgNVfSm4NKWq2JMd6vgVSxoEuzzZk
0OxPj8FB9S3Xg3Lro68AdHhTpijW25xqmJBrfTVBMPzHAEPU7B3y+xsUQ+OB7/J6D+eH2sBSB12l
g+W0dH56NgfgIYpSVQ5jooO5i837u0GOzfBmv+JttbVA4CqSlB7GvnOQC4CEJXf151iw8Rv7+6jO
bpBWK0xg6sclgaH8x/KM4/t4NP+YLNlCuRjJQulD6syaXLqtRvRz04nh3iuNX6v2xJ28e5nvnOy9
dUoGFApzzUL/OMx5gJrLgijy8dBURcBgD/GOVoicVYWU9iYar13lyhkiIf/V2jo6bJzFfSBSuHBU
hNwXIdT/IQKurjzGWuFE9TZ967QmcjhWXiM+nIrxo9X2A09kNQ1Hf20tRjYRmU6N/6yChbycNHpy
vL4AQSBK7po8NRVUk3jS/MAV1MCkht2h1zVqZ/KRy+dUkjX+M/CSP7R58h4Ake9bWz8dVdq9BbQ3
+Ys+26PEDaG+uFVOpuO+8/xnJHcTnGlwQ2fwwbCkZ0vDq0onr/3hqmy8POSL9y4lM56Y5W/8VX6g
019sV7P1qpe6hlEXZmnEpmBLhVEHXwtIL+AmN46+EZ/QkGb5Qa7LH4wBInskVnqlfGk7gtuVnfQ7
7NoqHSwvCwTK6fQtO2CH7gGwmrM4gsRMPbiejd6tffczH1R5bdp2N4bIje6A3V7eUUPQHvYZzJNu
RwLf8Skbm/nq2dwsk1X+hHq7l6T/91HxyxCw/wQAl+EKGmGpo7+awqx1JFbFBwyicsRuAZHjNdXp
3Mm38Sz3srU6wBMsgT/LAv++mSZxbmNdmb2Qt/56U0jA4tcRoqFcIG5vaNCbsNlHLuwTxGt8ZAog
kIDi8IZsDDP+G930aaH5u6wer1mrIfkeEan635G0+LIUBm3yZZ3VpyRMjtLFVOJRgM8AegOjkmb/
25bOVku1A89UeBhMZ+mfHm04bb9w2AeUWId3iAH3pwDHqrLfv11amx0wZXbeG/98NYx610Gb7WI6
vCQYjJH7rKhfngqqeqh4RTLR8bD7ghwqoqDZNvf03cLPJ6IixviTxZ7PolMBOrVWDxQEwXMH/wok
HU7DIp4lQSVLCvwn8oRm8VivO5pV/rtJUOIIl1KEYldh2y0cKC0SpHXjBJd+uDe/EqvEC6IhQEYA
5eeTHO5e05gf9sdEv/dXe1OBnE1bad+iqoVF3Ig5S2EumbpWvivCBcz0qbDG1nbgIwyOAecKQuNj
9OOA/1Co46XWhWGbywJupm9HwTP4XkMf2PwBEq525EbJxC+5QNYfbAZl1sH5QmK/ZJWy/o4pME+M
BlFYd8uJa3I25bOhTRxcqqfAT8nz8qzCSQkWM9zEZjSRWeRoOPSbyPoW9j8s5fWX7l0PO6yApzaj
dz3o9jEgXVc7MqxmcV3KfRmgY3XdDPoBhh2fuYGROCcnsC4y1CXmj60ATz5UrHwU0TGlt1creJtw
lYvT7cd4gSSD4i4hYDXjh9y4HSaX1eOeqO9Jx1tL2mlFiamdeJFkAuFzhvDDQCvcnOTCN/3ZcoIs
ebO6aLPXhYFCddHUM55w6rHnrOEwJsnaHydOpQwKjCxFbG5xmxVABsbs4rJccHR8tfESono87nuU
xcGo2fKgJYQO/Q/OeMdYqOk1yAThjENX4yFWURENPbx2yqIy+0eEJF3NQPBUdVSlKbxCQ8zgkRa0
ZA1oyLQhe/3iqstezYkm2ecQgjAz9ZOOJu/3PxihdR/6zRuGRdFXwaIUQC5KvXc/erHUtrMGF8jL
QZ5PPDo8W9XgMpaLYQOdlAt6mW9nZSFsHhYEJFDNTJuVegLN8N6TscNNDL/mkQf4oKyg5pEN4w5M
X9SZqVBZxYqcIaOqzK6Tquhm7KeE/kiayCPbFduNiE5XyTNJFPPYQ1Za0LL/Gt08PdsScY5NFSJ+
8Zmr8Yw1IvO8oooVuMy1oPaZkhQoZZSgy4AB+YdIkSOKXXkXqw8HqSUfcTYehfJuneyoVLpP5d+l
50TqRkwv0klKV3eCMDx5WNiN+LGca+ASmi/k5j/SJMQ9mgeCtQHa69/66gQ/RlYVcpC2QCULMF8p
km4vTAkAm6oKuf9sPkWYj7yjvL4ckGvYxwcaKbobrtXgiAaWO5OU3XosCIEY9hlHZLwmz14bTZ92
yys5ITzZZk8/AXS38IPKumAOd1zOkwuBPWZXHTpCjjvvnNeqYyNoIh3WQH8W62OPbC1QP44V6zH1
XcRbmCCBefSXgG/1fYO0e+Pf/rpzWYWzA23oMJiOjhLmzvQFZ+eIrMDTtcXP2VETOMG2n9Odli7j
5uxU4R4v+qAEzUMjUlh4niyThlZUSebyFPLBUdty2BT5T6elIQ2+e4tQAwgUFQDc1mGKnDQYGa6P
utBXkvat4bAC2vH1lpDnBsXNXN4Gv5ObAGl4qfBAMtKTCsDPvCKZQvq9MZOQDnzoLhV5Lqf2tKac
q4DOLIDKI0H/2yZvSLpXuo7rmq8PX+xe9pxnFtmTzWMG7SB1vHOtMnohNwMtR84x6PjTHGYr2TZL
IVeYuZiOXNhcQRHmApBCtyeacNbh3r6+VE5HFDCzctERPsXW6IJMRv9j+XAZJ4cRqFFs7kUbQe4Z
PTItDcsi3znH4eqvJjo4RR5rpBFINFt7BdQMzxH6PGGyEVkj2qzrjQvupsG+6jaWPlQa38AdYXvX
X9oXnR4rrcQaxO5DIfLVStk7hx9miD5ziQLoSujB4xv6SohgGTVQSQNoRBSvryqXujBREGtIaX8N
qoOEQaG7vRSBePP3dfjsh0+G+D5hZtSMsyvZZsXp8JgDrYTH790sRYMehrGQhs59tDLmI0tRgAHK
SaCUG79KZ/FFvpFS3NBCvlkdlnci1mNlqMO2mpgJDpoZglixqAhAecnvZoMOP0HyMBks2uCAOatm
Hn5ZYswZqv+XAJDPmTgHMwfrPw2RIdXSpLcRaW6tCBxp+eM8OV8xCw6Vh3ip7cgz8oJ1guOsvQNF
oNC7Bs+lsoCTbLUQ/uKDvc+KFtRqmAscZhrdfuZTJLzB5CNEDfRgCip2KUFR4vNmuPU2imoqzrEQ
73mZpfIMj3v8KAHsVljjbWMuUH/0/Ry2eRWvDaluHwAFE6dMXiHIHwfIQ23xNvgDQXWALLUrTiJB
Hkcc2qdgFbTmGLxUQtTiCGGC3M2QfRqyrEDIaoN3ZHF2HeLVSTnMZRfRdr94tWa653keXLyXu6d6
fUQoxvufNK19Vdi9otwTpxnxetl83HBdgv4E1+oKPessA1O+QyuxPjILyImCifzAld9n0MT/KLb5
2PwToEI4cY53FJHISo0eeCJTiw3Q59Af0sBGuHopQlQeq3REIvjXDpO3U/ZpDBgbbXXllhpnZ3qw
WA8jkuY8vWs6UgkTvsFSiwaIDxPJpUYEvkWnLjzo46Kn20rtyqiyJe3L/PUxxanRRA2ar/tZ97cn
BJVfBoFlMCKfl+fCE20Wv5yQrn1UnMDAeZpa0vbemTshN9KGbtIBGAqFy5fl9Nj1KUbgVZPx3BDm
p3gx+TdFnfbuNc5fRA6UWychmiCRL092OoeMIvec78Nkbd9nAtq2BjWx3PxETW9IpglbfmIjMRFY
My1jDIExyJMNYi4YtpeT73VLrFY7751U2bBNZJd3CB+HNn+g0BGN8UzH0gVKId4sPFKnhBk7zXDj
KK7rE7CRcWUzGVGyE2Rvfh6wc0A/rbeDGQdDRd32UNAxteKVVPKCGTj71t2OfXKsT4Ge3hSsHQm+
QIsEY9jfUE77Qn0eGxM6oe0EI2A9Nm37K+6TpJZ5ds5uD63ZqLKPczzVad8agFkyO164dYqis2is
Y+LD0fyeSVCsztlS1rC/HwwP4Kwr6dsEP0vx9zIUk8eJonZCdDQAwVzesRufu1KX/umKaFdRnzxa
JgdJ1cLlz8kmWBFUxxivDxObsA0Wad3rDJDQBbHkxJAU+npizbtkFP/Sr29zbNVqnjdJpW4KkkJ/
NFcYpoTiyZ0AWP8cBY9mcE27ERAXGr6BCsgOaeZxCrAO+qHSvMq3YtMeUrUhrcYT/0wi2K9UEmwj
Xr+jJIJnnt/6Rd1cJnDLHUaQhj4jaBEcBGVMghgrH2edJMuYbWJssyl8GzT0vbQSqeQ1M45z99P2
E90S9PJ6g5m1J7ljoTLWo+JwvEodaNa5e8M9qr3hhfw+FiS36RBU09fqtroxIPGDGb8Ut/+5z5Db
W0u12XZ30+ct2f3hYbGQ5eVYHffASFaO7QFAQUPPDnNEhRvagz/GIzwrqnZEuwrxZnOauJDQqlbo
OWWtlsnaeXuwyqo8kaUSYEm0a/J++MerW5Ds3XiuzLVYzAJcW5wuiHqJebg7qak6f9OkkP0nlygy
zEGe7J6z10CIb+lYp1Vk9EN/V9jdtCd8Muqz0YejgmA0TKJdnUJc01aiM3IpFkXiZncnmNBok0kB
MOET6i6BWDz11WIExXKOoCAr0hd8Q6NQ6URIIRDxKPgOR+Pj1CQGaKbOY91EfTVovUseuZAWHUpG
oxTXw4ogKfemhZ8XhH3hszuc0TijE7x6UWcNONsOhKoCcfmkoomN/MAibFsdvcfvVN9X1MneKFdt
nxx+I5VEwZq8a0pkXFubgD72qlMiRKoj/xIguLJwOAPHLObZJUOg4updYMQPj8Ghk3FCWhFbtddC
itgBEkkEO7XpVg/K2JFmUckI4owqaPprFXBL0sFnx+AKfdA2wc6qW2RhtygGBZHCTTvNq+azhjE3
Ac3l96jMw1I/K3aM6PPpjDnAMLHQNX33h46X7kjOMuRMYh1Ux0++Eal4q6WSiS1jSUcODamNAdDs
pYgwdjcJHLGmtgqKeDXupj048S7DAVSe0RFVKAWSem7+xurr9pZFNpasqutA3/25VIfvB27w3NP9
hw3bN920aXi2AeyfC7PeKZZwb/zWXmBfP1MOU3Gzcuup7lIi3M6RrdeIopd0o1rl3pOLJTCMaL2h
3kHYGqzkRqssCsciDMTF52CsgRpqtI3ZeSeghB24gOzwdAJS70QFPVbm9cA0wrIR2LnIX9zBipQn
AFRmG5yVVfGREEF/vNoPq3CUxwaCePbsVpOO1TsUOx6kY2NTupFUYI1vARPf6L5X/TROhXKKdQiU
EKsHs6jtBLcCirvQRAMHOkEu0MzzwkveH/cN3juUnjEbo0oLV7RrHyZToUJET4Jk+rfGO41Anb71
osg7Sdc3qZnxMDrAAajKAp/PfO3IrRChhOMEa+NHrxsGyTV6Xkd5VRqv14k109GnWfQhStxUHTOu
KiyhDYsCmdM1Aw0O06eJK1GjrCEZDnsevpC6KJWUi2xzXzu0AoYcNhLd5GF7lEGZpArN53BudwWr
Aiiev3A/p8+KC1X3RMYBTZIg+4P2i8RR3V+qZua/Wdz0pAqcHdXY6KsXPgAZ0Nq0XuNaABF7Cd8t
pUbRS587Mh7CmevKdfP7cbJ/85/OgND1buPngKyIXxvt2jphB3pyTcDVms3uhz9xbrLa3a9b1sl9
Z8cfWXUWixUZvUB8BpD0mkoW1kt8UFbMk9SKK3l0UvfkOPSQpwWntcyhCYLPXq/E0lzkcrQIdJDy
RJ1PNuCgZpQ0L03js9KVTn7XF0IYSgtg6kplLw8NjLaUPvH7n7kYYi+aEkafSZDjEs+LclDBJcIr
lAQYL3IGqLpXrj3AVKSc69tjvplE5Ofyz0VdVpiWOvvZkFLjR+3G7bEBlfFcccDClD9RUxgrbM++
yeaGn6u52Vo4KjrAAkO0tOIxF3TqwbU3/iVS2VQl2SBAEwytf1z53sa2xXqD9vDMFTBeR5qYarpY
/5iBkzTMBz2hlK4DAtxjdT1bfHheE1m2Tr4s5t91uo7sEazluMnnZBuB80ngwbzFaJxed0qw75Fq
dDSoOHWbNnOovuiw6L2d765ssHcMY2gtgiNbYv42p7orLZ5xGA3Aws6JFKg0IQpJOebxMLTjgmyb
tYiDqKtGEeUuOfnMNWieLvLBrSPQpOnfORxqUMBSu8PH7pJRYskwiNuoApAgitjYB4nIg92qcJcX
LtXcazguhGMFDzfY8rAy4LyGZTHvanTvZZgLOYOjbdSNtNDdibHmmynl0XmpyeS7Xka/Hl1PblnO
6IwA/FfHBjsBeok1mySVN1s+v7JjVgbkb+MpA4phY/zOZDn/ua9VG73m1GL87EBUnbcxDekkCIqz
EnkZbMbh3CMGkz23PgCA/wIHH7lF6iMOssP5DcAP7evLOVdrVpSOUTuTUCLsX0IuzWnqrXfQhSBS
QxwnXS3ZPAqs2tFEot9ui/OmVkCSLYE6rW0fmd2/HGab73eCpLLr/OJwD6/3b86dtSaSpB7NB35r
HzPnZZ6A2hgjBfl3z9PrBgoX8QssT/xaiW3lI7yVDN4rCRzVbNj1okv7EypIlJNH8Z1RqEnkLCHB
UIIYh0hqWcC7SJBJx6/DB3AOVXN6D8+586NWkv0PENjkK3xkmgpMHJRBzUjhz6KcoW0qUKmzDsnF
53wHFZ7CMXwAH3YMoexVsnEgoM+SKPPwWeGVQ0C6SMVxK7ysRC0TYZ0quED4ENIVApnTf1VW7gqG
x5zRHEqJuQBcIaK0hTkmn4Cud5lwIn+BybGXTe7k/yfC53Z3qES1YKbLlvZsH5l3HxproDekLfkl
aDRj4pwf5JKltJ+NW9aN6ZilJQgPtE9hclclQbmXTl1Gfw4HBBvCI6N9eIi4GDuHh4Cmwk2ikqkA
MkzEb4/dbS1p1oYDt+XL59dXrS2VdPSGf/HaVkIM+RNPt+fLoIt6+bAcPdnGsqSAYsUwzZ10LZy6
wmt22eLKOFwXP8m4MCmh5oNKknuOteptPQwdrRm/FaYLABFi2dlaImobtvm5utgHZeHvlIaxsfS2
ga5QNjzWOYN01MCB3dOSGwE1D7cA3kUZO37nLY7X3z/gkCImDlDgtu64vV3iolZ1AAhRBjOKsinD
YsU5g0ateBhiHeG5fWrbEa+MYkhAQ8WiDMTWuXGbyqiyG081SYlY22SbdD0E2tfz58TFBDwNLx25
DVUCWYlqJ3dwnHVcEEGfZY/EEKRu2lb1qpEFWOsc+8pQJB71BAmprLF3NVTZbfp2LrIvwOSpzmkX
yV+CnEw52ITPcWopiWOqmYRmU9uCfedmHWNFOaDsOdI9V+IbwJpR65SSj4AgdHs0AcJS0cnq72C0
Aq5dskAeoJ28dPdUcqwgITuhOqZ3nNQKR1P7TdLD0PDGfJg6XLSUw1v4YX5m93ItJ0y044j71p4t
Ap9pHH5MlX9VPce2zpJUxyPQQ1SbKOs92xQiY5dxiLx3am22RKyUqewnY7uZ9ckfyECO2B2RtLPw
n1540xl0frfrkVp12hpHWeqNDotRZeFsVww12TCclyX+uY/aBUQtItbFu1ht9dxjcRCnur46Zj9a
12kctWbIDhqe3tWlSDcugreUBdxPmMaNbZu+FKvY1U4mfQqtnGmnF/Hf/Y8SuX8gdylSc2mjWSp5
jZPJT7BsakzIF8AJKuNeX7UM9DbLewkgnClVuBbD2Qk2SMUDt60NslrprQx77wv9tAGkWafZXWwi
RKRxyiRb+R2QLusXjcd8lTeNLVnBYYzCbUGpnxgGsF49Do1JYftqUIGGJWIJgS3wSsVtWlsebh7H
mdF2AJSIWzEzbuLwo3F8j8ZKx1ylmOssBVR/JUw8Yq1NfI5twX9ZyI6IgHpKzh80byf94iW16/Os
+meQ3EU+ESRJFBak0iqDULHdcvjHQzr1PSYDpYqkP1RGx/cS4IXfKoSII3ptSQJRnjWRBZ2ts2jX
NcOjm3WOvo7+TMrYUIemoaiOjoHD4MgfrGK+A80dn/l6B3TjKP1x8lmO5/v/Z4n9u4nqPx0tshFS
OUNkiY4Zq61DNQdpnj0/vkprTfK173aAh4GECbij9dRVSFCNmZ3nZlEXp3/wicTogtWzyxnpedga
wjGsJmG2UfRDWrL4tAK32W5RWU3LIk6CKlD7SST9h2WRhJpPyKyOZH41f8x6ZKw4kn0UtzACTIe8
2fvmq4bdB0OqlmNHokGAld+/2w2T7JqPIt/eqmfGQO1ANWDyJ/bazXCQwvXa9yI+/OLijX/Q4Ah2
DncVhMKmUufN/uPCeePcq/V7wQ6JjnVnX0u/0lOyrqGqS1YKczLXuAb9Bo2FjoyQbpwxI+JnLxwR
xHY4QSIpSv8ZETfQ2qJ74loTQLG96jqCr78xA3I9N4HOTq6m8l+KrCx85CrukZtzA/6SsDhltNz8
sJNe9PlRuaBKebLxalKu5eaDdgn5glV1E6bmktJjo5g782VA3biNNBtYX08kSSgipM7ADh0EWPQd
KCZlO1toGJAIYz5X9gpv1zAOLrLW7ZJ/pMN9ylFHyaT3B2wvZmPYEF5z2ATvQi3ITDjyQFmKwPGC
urrJfrIbBiMDs6D1Gw1S5NVjdzPLxptdokgiH+0C8Ww5ths69RvL/mCHmQKL8ywd1aHKJty2g0bD
U4b/QpF7qzbf/DLoDQ74liFuNlM1bV2RC+cl9q7jS0F4vG84UpJcZKOO6k73UZd5KwrHqVXmIYHD
M06KCzjCfmGh6yM6/IiyFQKBEtB2QC85lr6+aLJJVxCuu2PyjNwK3BhsqxRTmT0UFIUI3g8Is6DD
Vnno5XQ/Wc9A0ZOzRgnwd3wonjimfyIdEhHCxEhFK5vu1glk+8jZ9Cy3BKmqsyGI6Ecj37z78T3f
vZiOppkFkByL6RieRrZLDX4+nucLh1dyhaAHe+6iFRtIHRZl3QSHbkO3A+DzhUPi4DqlbJulJckK
z3zSBSCrZ0QEDPWpy+i72OJSjoqq181eHu6k0P7RKukQODKTXPCbPuMOFRNSAqscWs001qeiJlm4
j6kawulGfNGgcMMCbmqmXk9A5cvv/x8180ljVttfOTWI3rhNIlFS+LO72TE9ta9yNaxVBI+E1X3G
zMoY1sLgo+JDYw/nY/shwAe2aYs8Pm0hFqH/aECV4GW9k8aRA6ap9tcJPpNWmmgOXm1ggB5zORZh
UB1/8kBwzkEmkxd/9jS9uTex+2ZyNUl4im/G3vkG1+5SuSUsSH322XYE7iZe4zYjsuqM8k+4Vws4
0uZmlxpogPR/xos25iFGqtE7ZiiT3e43ggxdwxj340rOJTg7BJovYUjxv5U0Y1t7Uevj5o7xpPFq
5ZVOKMyD+T08xxn2l0mcDljWRkr2E2xQQnnYYzyNHlczBuzS7FRh9jNfes5yICXNaUXe+oQZaVYQ
gYu0L1eWmoqN4TJGYBEnbYZEDICvAT5AD6R3vB7fxZzgY2mVPVKH2/VesYjBtzzCX63d/ThWIz04
uf+Gd5VvqglcXyrNcmL5eF5MvX83xsXpI1ArWd2+slYk0eHAeQefKpRLVGGz4uziK2qjjIY2LOkv
BhhHPX/m5zA31+emOKRhdH1PAMXLPcjvBWGdzsXcaj6YxAFENgqWYTdMJqJbniHte90aYwvOVN3k
HSLmprEGqtMlz3LIpottDgcPdNzasukZ6ZgggNc6h/6iNK66KmoBUksKfat/LdgNhl1CS1yABozx
0s1iaOZlRn6c0VGOWwuzBuK+1EYVfu1kl3onYKlfJwbJR0i4BqczEWb9VHl7+0UcAmeJZsF6TFHE
3a5dJ+zCfJgNmqNFUhxwcwFNTl8T2lYvIRK+pdy5JreNSGISsujtU5bsbPXoqYV9hbI9UMmgofeD
VqlmwULnOmzMzCM/UAJaXgZOAiVwQjl6K7aYSVxxX6ZQbGxNRpY8+222sJtWk9J4EESL25Dq48W/
WY4LvDEECPh1yLOspjjoPQZrWByjoW412RaNAlSE9Xnhg6AZhlUVy/2tilNeGzLS88QGh9SLrq5T
XR+5zhS5gbPgyggVLXyBzMJWAsKXNBUT6ck+OGzqDu5PpfTidzi96GIie3GCeGaB0jOGtILk1AqL
gQVWNoKRKd2MKVBOdeV4zfjr0fLH7UMWKkQvYaezd/Fa+N1fQlWsGZrNzUdV3Iy/bcmuMekK/tAU
Zn+M036s6Wp3HUDGoIDzZBkmFysLJbz+Zh3ZkqD30s9X214S0dK0DF+04279qmWXrmMlZjepf+2g
LFJetX5cjiQEUtNvcGL3KXmEOjyxtUc7XA45Va9BbPVkBCmPmEMBD5nKFd1pnCZSDTMsp5CBNcLu
wPh0Non3sMc3wPNUIqUhhTgbKSe7hXcfYKM5usu/NXqV+85OteDnetGlpCdJQBjfplN9XPVJM3wz
q2b2jUOhS0tJBuRTerP27GQL/YyRrp5n0yuonwbTFQZ3G7I0zI9OwIw1QnRw/msJC86lDVcz0j7M
KCojGb66E/J8bkjPWqizzqi9xmFVW42TbKOUiAxxNoc+Jno3JQX7QcAVYqMubmGiS7UgRS+m9X9x
2kTJ2fBqXNuG2Yr6YMbQHULlMwAmEBIWaGxoi3/6b6QnF3gxkVso64EvtnEk+pOLJgYzOKHE+iZP
DgrFJE+mR/UPKiC04Ofx9Dc2H7HFtu/aTmNO6hfAKxT7BdIFyLQCZbkauleV/heSGUZyWnVvDL4a
knrS3D0uQ1RV8Saei9wbVeqr/j14K24IcWLoO/AsCDUQ+LOUksSib9YUKt40W4c9+IpPWbEsqvDA
qY8AfI9+l7F79NDKJSefPhGaN/DqlhKGBARywUMxJ+bgKhZDNmorLWbxsOAz10mUHSYrMpmlVu9E
SBetxL8/LV9wngx9ivzvXf43XFHtJ88YkurZ4oK8ND4XdQhTCAKpbX3TapzwRbNCXGE62yMmqftf
QodXQvOKgir9fcNbBZ4y3j3bojaHozc0sg0O94jsqSJUGYFSW9hGM5bLZv9q55cXpcChXA69DEtp
rOqtR7bHFdKiEdls6LTBXKVTxJlrSA62QyirzyPkNAxKslVHtEstgP2lEwLw2aaaCi7AAxoTKjPB
iVAWnmWJwYmgRcSUUEfOjdl0Hhk4xACNhuxtttWRE+UN9EeAszYI3RLdAO2LMlS7VaYnKWT0dfvs
7H7B3D6CDNaeEvYoI5JskjO/9CJPbrzo1gUvjOqXFDkM85pohOsDTrVWL2tAiuXUSEJKF1QFMbBZ
8hZS+QMmSxwEf20FxZx1GVn0kLt8sz7wJ0IprTUe/jcmXrLaKNDjev014zzIFXkxxjYjNlk6WaWt
3qn1M/vTUwyNvxWd0mzINz8h9dGtcFKL+4LAxhsd1q6EjOz8ulWdiOWismIGwMJ0jgnlwmha7CD0
5BspoxwYXaOigZ0pU2VgyAdAjqWzFd92W3I3vFWw5GzMcWd2mOtf755HnTwM4AmMOFU83TMSlacQ
TNDX5pw34566PC+IPvPdIO2DT+bmMu6TK0az5Q1+0wsuSxsKJmsbafCW/0VsshAYb71d5/WuKVNX
0HP5HEYo0kZ4++n/GUXHDASD6vZdiAMIFXMBabIMJHkP3AwohfeHeHaiv7UMwq/Ltxs9LiSwTWP6
jMm93PuDYGol013cRsIgKVjYeiSEaquBL6ppoAa6C6rY/qgJnjBA8/njpScTMSVV/GkOAPAnXc0h
l13D7+7DEcXHOnq4N0yBlTqwo/shMHdOVWqDiVarfsGRBqWq2d5oLQY9HXJNwoVEpNHj4YT/KorT
QlNravwPfHri8jWU+ekFYiDqxaF4V9LSqrAH/+7gAaH4vrRnhf8g0khswxnXgVMcjlK+CjI8NDNB
Qbm+iY/y/7kDYiBCa05717yqxLXASSJwVgAR23E7FPyxUiGxx+VkanPOHwcP5pvD1o4/3FfDPp83
tOyhT1l/37jEY/XO7sC4NyyIe+Oon+H6DDumifWwIm/PvKFsxbyINZk589h/RxiK4OuSgAe43DhH
XAgEuNmDFecDQAtdZSbh90XfGmGjzDQdTH2aIwONtdj48tIuJyIyU4YbRKGrtErvkXWLxSolNpIG
xGT6OeSSA2kWpDuMMR+R9xodoAWwEY+9/UCjz8y/O0n8AMpxwhVYNjl/5Zldzbq++zEPvjCGOCn6
eSk3a4QeNa9wfX5jkUUalv2ueu2mmcaoS97DuilFeObZP8qU/7F5ros/rKyF8ItBUYEWw9XsPIhg
KDajjqiYJL3hXJMtUxETEz2BhjZ24LO+z343j3DRc8rMJTirWrpcxKsznnh5emY2jzLhKEThidsT
thCL0At81V7LcTkKdc7eCDqgiSJByCHgDV4J8TSp9kJ5DIGBlPJGVT9AXZIF+aao3hG9gaYDi59v
WZEO9cin1FAiURMHr9CVDy45apJ+FZWCCfs35vg670tcFTSexCJtMserg1Y11Qs6FGcVquR9YMpG
V68lxWBsaS962cZifjAN2lTLv2e9B1CEVycl2wuGcoJgmgxeTWKiGv1UfM/MisaVxRnVCk48VgSB
MgOPzOp2aveuYCCCVb3aAWRekKQdJwExEoDCDeRfza5JivGoZUW3zPxrzOuENCPS+nKJCGYZ6ZjP
Up880G7VtwsLY1hQQiwmviPBygd9rwkhlBM+Q0/Q4ehyCXPIGVYD5ojqC3iwKht4WArcO+dixqdN
LK8nJLUj0PsJ1CXQaKi6/YmEmlIYT2x80pm9rC67VB6YVMix7Wc3DbrS8elTJ+hjPP813kQgdk0B
N1Adn3VBnSSrXIBqxVHZy6IqdWbYtNUPuSMJC8Zd3m5lhK084Mnz74NtMO9TWLHjJxZdDKpAHpS7
i9RA23BHGd26pTDankcl1jfET2VFqZnr3UueZ1Hvr3T7ilsJdHs/6HArf7rjJjVspd14rEU842W/
m/RVMIN0mCGvkDDynDLVJe/AIBdG7MgkDJk/eMleYmQJFGNf1ZSm6IQg+1hiHFvTeB4+wq7NMgaa
FRqscoZaO5fZKW+J9bDu301OuXW43hmNo8bj8UvA7TRYy3lMsPnZ297xMP70zfeEm17g4bVC1Huc
JvshM1kvmnuE1E+nPTGWX5aY3D+UH+WZCLj25Fgar+JsB6Nl6x0lTtJiKT6V8xQDkKdicP+IFDBX
q1HBvcA0Smhlbif6pqqSFpM3+TES9e8Y4ztjIz/Vt0G+QD2rzEl5M48f6EwS13W0nloaIDk8rI/Q
AQIt0Md6K+iiK7Gyh26cfXakEtXeBjj6wo47cwXWhSnrEhZPeeEiClEj81eP9QZvSaq1f2LfyOyS
sdsdMcG8DYQT7TCCLllYNcR965zgdeqGi9odMBy/vzRRjLCkIBd78CXF30Nii5Pdr/DMefgGg5ZW
jwmu9hDzlGt4dSGibsV9+9jZevjR+FkHvmzUo9j/+LfzhKMAe7BPQurHSUk4Cg8+00CeM4RZve6l
HDPM+qm85wA5obPI2Q66N0v1rkajDqmmHHfEtIWGseEm4Jiwy6ml7VKb+mBy2FMl9Ue+V4oZHh4T
CyJzsj6/T+mT8p761jSE3kmampMtJhgr2R/85aOtxAxmUIH1UieB9t+K/A9fE/sfqWm6hl1WcOd7
X14IyBNGdGuQcce+IwJIk59izl9JSuIh5KH6LWLaT8KkfOnBPi2oXbRDJNcynuF75CV+bqw47nnT
nPkI0bfI24uEmZmpNPOMBsLsyw69pRc8uMGL11HkyF+RL7pxvtZVY76b5k6gHgYUoShth1Q9z/rL
R2+OgUrYMCy0olShRjkwAM9adkZW0ND2HTqnshorWrdQiAEKvZTrmuufgKZxPZXkwV8b6E6/1ouW
1qoOiMgChtw+9fBwxGGt94FkC8XqrDgwEoJU3qLkLfo0ueFvZOb32H/EZ0cVn6mFmSFwJgk/a3fF
GDB0zZwigBwHxN6RzAF9z1QAbrPGrAWZtnT2tuRkpVq8GhaGGnBoNgtEVWe7RvSWSWN2rqDEiRY2
3KhNHGslig7fCcMdtvDTlj0I8fuvrkajx62vITszbmgKxjKRpOSTwo+jjzlEnOBxjr4cHL0KhmeW
0kG0Nz+yKol5KPddKTwsRHrjckmc1ukg1TM/UtDHN0I0MHGmu4Fiqv3g2Wj3HAIs+rdC7Eu5U0Zm
TDBARj6nIlIVK18R3cXszURlRkC7oLlB2v10ieQgVX9enrLPfsIRZBEAYU4UDtvbQ3BdPEjEeOSc
Shr1cDXoRNTynCXuUVfXXfUI0rq+LTlf/BcUGiDs94fRLGP1dtFgCbHM9XlyNGM+xDdU0OvGAl5R
k3RyiAqhNL9I9QA6CTbkUaTypNMRcFXHsl/8HOTmmRRz7ZyFtLMjAo8UH2XZb3PC/XgjPrEXESmF
hIDHKpDE3SE9wTAPwOEUZWF33NJMfVhhTsKaPlQFHxbZH9oH03CzN319MME8yFy5qh4Z0uu72J+I
sIo2mFPVvfqKauAVwf8CEt6YMWNH3Ky87zSe08X7M+A9/oAMfIONsIYgg+H89QIUdqLRvm2zD6PC
gWjICP0GF1RRD7Twc2/LFLfXmXhfN/qBTtqkcHgaHJcqvRTvgzq8ausPnUrz1msOWFDmCfJp/+NA
IdSyEfxJ1s023lx13d/9cIjAUB3QVl+J66yHm83s+QjufXnWA1MyOwUQwsubgL9v0bOoZcD4hkIs
pKxX4vLKSlTQCScFYbsJYsDeygUvgFL9eMPWmhwXf3+V3t/Q9e4NRfCpXxvj15suCd7s5nB7G/G4
5yIspIa5iiopzWE2EeL2WO+NI1oaPWj6i5viLUgFflPR/ajHRMHyZrDbCw4Ddu955jMpuheQlMwA
4rwUdlaEXyn+qx+EQ9S4fElC33aPJJQUxAC/gCcjnclJrDUPeHz2BHmGTJNBj3evsrqrvYZX4YkE
2pkWhJu4QCRdDuFXPNxv2pdSxhtgvYtnWFKPULls89gurJv62SydBhFsjuVmkHjG8YjqGodowNji
8K5umpuuYHdKcCJYBSZiAsTDmbG6N6Bnk7X4LGC/vYxznIkpBgn4Jg0V/W0geYEnKIGI5TCUsdnu
k7BMyw/8WpDoOgCvojsZdTWVuBdbGYss8m7ms6WODfE7Sd1ZlaMP1xwSduAh4Gi/NeDA8mNKX7AY
8GSg8CSHSUI1cgFH1W5Wud3N3/fqYKHa7iQl54K8yn3QSr9HJJUuZeQepFynPkzzfyabsMrX+kgN
wIWgVgT0guWjXJPMD24korVuHW3I2cNW4G7cdk3JDLyPb2/EFQk/8QCX2aBCICnZ9Ju6mkFidLt+
jyUc1b5h/DAekiGfb+dgha0QJ8IT8YvMjk9rTRNnXhDwxlkrSY9xjaTSUPMYEzh4fJTQFIxlkx9B
7ngRLENSpYx+Gzp4h476qJOda9p3tSdXttM4Q6EvFKtDLOjhXgv/7Z7QcF3rk22uPQ+tl0IkKX39
pd54iBNnsanXj5fJ/rhzJEB3Ql2uvu16/5cWHjCkJXOooXqyzPiHGwvvSY5GceaxljiRjeYWuq3H
jPWJDlC6XCInmGBy6Moe+lMPelepbcn3IC/VI298jxS07MHMAgAmu0XnTGqc0aPsrtjUzb40GdsT
Kq3nGQKsj0ncHnlKqgFyOV+79xhETIyos5GY0lbUGuV0HzKBpKpPaDakNBVU6Xb7M7SiAnWhvU0I
xnz5VLJUIASg/H9FAEW0xG6y3AJG46jlY2B7kKni5Bw4lMwJOYWBPQjh1Z9MMOWcplAIc7HwekKN
UCQvWEcuKqyNWpdadwz/SX7MkERmgsxNElLx/F1U0Pi10ff+QNeqwkjyuEoqVEUHogfLNGnuj49u
28XQHsW5ty1saiG0SgxCmt+9IdNpO7w0MJa1nnGtW72kQkPBzLVFACgu695F5N/w6QrEl2RNTjeA
5l+yPbd/ElKEZh1lAQvwyH6jPrFomG/Pn6hjyC/AvLJaziUmKUXhdKKxikwzfHIgwAdpkH9S10Z/
7gV/qrrfA9zzuH6U4N18wewXl2OYhvBVgzQuEIyVsnG+OOMrT9j2e0aiFyZcv84yuW6u7h24cmsY
wdeJcCl7u5zGVvZLOeOPEzEY5aSAneKyzBmOiNG1U/v+ZniwOK8xyTrUnx5xVVcSI7opnvBlfPyA
eYRjom5x/0JYzAXJ+DM5iqQZz7pASWTcr8v68Grim0id/YMh1Sp9/Vhi74/1Fc1GPLIW0/EKoIlg
mtkXPHYxqI4IGYGL88pA8nSair802nJOwwpVL/wo+N7JIXqb4rajB71mLUNvXteTBro5efNgNgiT
BmRWRnhPcGpdpIjjZ2eh8oML0dPSIJ1BO1zG1+0NZfa+xAM1i7qguFQ1cXKeWJSRMOQN+nZ57Pn0
kCott1jk8GQunPYF/o4HbKRl11eA5Z3/rtEfqfn6l6cF3WXgwcFygLzSYxyJC1F/sEMUGG/Xm7Ih
6D9mDFILvcQicmGkMupaLBmZpji0ayvEQhAydAOuKooGggdwtWIVg5+LWiQJZZzFgmuTp6uI0Rmo
EjltcfnRs4HDBvQdlfJy1dPKBYe8nDBCcQXDyq617ljEt5nHidj1N7jUlEPGOkqkq4Ben6Ul8xQb
R2aMt59IGvWXUZUU5Mp7QhvapywpBfCj8bpVEn5JeG86gAXrpdTh37VMnC4zf9wsFJnZ18rICfWM
BnDz0gvEgAgQ9cKKPOjA7bbc9vxAcXkxbPd9YE7r5JkpE/3vESJaskRs47nSB+S1QoW564GBGg5T
9y5QIZN6dFD6BwC2ZCA1LDkAVvPXJ1DHmM0mRcLup0SjxsGcaRhiLFtbtJqnm8nM7amYo0+66ODu
cIQXhV4JEM03uO/aGV9KUDku83F0E0NdBqPTDXKgRwAETgjo6I70OZghZGgKwfNh6DtCvEMdOg6R
d+AuakltX2TIAZzdzwcj9sAqzVUCpKSPxvwSKPbeMR4FjVk0GADy1N53F1Ispj4L8lqvZ2hcVEc8
k0S4/calJMU0AWCIydoUr6jiBE9VXS2P45FNEA0zLnZJo7C6U4fjc8dch7t73AL/9KjOSTLFUegm
nb+vS81lq9kTvlEJid0vTZXF+5V7+Qgpy0dEng3uuxRQQYOhfDn7GZdKmpVJDpYVYteb90zcc0U2
Pi86ELfJO6GF4dX6rUCv4fAmTCoj1BZ2A83g0fUXCECvwAgDFkkEM7FVLugnZ8vLuuDwhwZF6+9V
n3Mryu21q/fWP1CFkTbyJ7kU94sUglSSGWYPbxIN9p8XhYbw9inv9z+5m0wjJlvXXjuNyezwgGXt
72FPc/0/8yKa8DbrNBRPbxJtd3uCxC1R78jMe2boyH1HyaW1scAjfOHjI4I6DTZxSZTsjZTLLPJw
0yPoMjMG7TFlSH0l709eHoa9g+N74czIboFagT4nzzNijdRunFZpZ3lMwM+Fa/uzXiT8gTYgfO3F
5Q5havZ8TCYJf9d6mRomRnXgu4HQKwN9zxYQPrCRwT+6wI9cw7ikOc70iiwIiHJYs3mbgF1VcVqq
g4ihQuykmTMp01xsMvxUQg8j1ktjmr6hPs269HwHkoxm4bxjjLWwZdL3DHU5vSFoZij8hclj639O
eCqpPzvMlrgbVPNmDQBIcVkmcvQRo6Q43Y1/t+1FVGiHvF1qWIPl74e8SylUhh18eDmnDWhjFAuc
Gny7+2G85bHEilXF1spHLwkXZP3uz9UwHCxrHFF3rV1n+i6Np762EW9e6G3iANM2+kh1H/bY1T6K
ZGEmJfPvoBmtGtpsKYokkFuQ9YvJ6ZWwSYg00Bwe+saT3aED/u67W3ucbt1N2FBxcCgGCbB0KmUr
Y1lpw4lRi3mqqW6YghYVlBqhRoRyQkEKLtI9RubyVMRv67Sa7CNvNlA+mBmvYmp0GrfkYQKwkDaV
JXh7TFsid0fW0nN9evpHjGmf33xjthgKfenDEPw/M4GmgM22f0ipHSj/xq+kdO1EyuZ5IgHkILOL
0IYfleM6xC4jm8TyuVSzEZ9pu+OeFjus0sIM4PKm59a3OPjP7g2HQYbHRzIccmd8tnzBCB0q5nPk
HbACN/mKClvp00KZKhVE3/UZvJbQsWgLI0ZzJLJ6TIC0UwSQGI9YANKRSFzDWIcDN5WNaUG1Jp1W
q7l/UAoXciMR9yj+Eux5HBziIF9XWdGXFqwByb2huzamtSt2CVQ/Yf8Kxu2KHVyADBaN6r5USGIc
z8GogIc5pXVRGd9THWlJtITiT+5+dqUddn1jFK45mf85Jyy9pq4HL3Z/aHwlQyh/PqzaLHc8b493
Mjt67OOPOxCmhUBxvQ8E1EzjyQIpbYIaJ/YVfsCfzv5Jt3VyJW5oipiXUXGyHKOU8zvLejX7xEaJ
KszxTYvAxDSQeeuZfv9x2kPylSHLbzYNL3NfmAPOqZ7KSVddIXwJ8lf2EF2JZEr+2auj4erdZP3C
SAikHvk7LLFy08F2ihyKUJk42jwcyY3vbORFxTm1hrQAOQzwgdaKeebETgbu9hd4h1VBSNokB3Zx
A5UOdQVjZfWBqMvInnCIwYMWQKctqk44wtelaRyjEgu161xPYEW7E3BRjwqcI96LVhvKGjOY9s71
vEg3uNi8FA0ACfe0Yy1Ls3IDuDvKWQzxPSbYQ1foVRiTD97Q41ZWENxxnzFm59F6pWdUA8rueCmt
Id3uTCKgU1C9aGNVmkKMyOgnvjhrohrofH2PsMLXTUakYTwfNx5Fly7V/wBhU9DVpcMeLoLr77Rt
rtwrcOgNOrTbr8IVF2EDodlB9UlCSU9j1d34Zeu51K5y7pBlU1uM2V+Pk++00sK4Xh8DtkemQjbN
2MVp2LbLhHXgpGP/D/QBZkHkIK73mPvG0okUyKwiPhhGW9BRc4SnjYPYxh6MyHlqEcTuANnD34dQ
4qystq4dHRSSfryX4AhUm+yAa8EIvsAS+h7aljFfC4hTJ/iSupwFRQR132GnNGD5FqLQh/XqAyuE
e0FDXHYij0Y2SBVWIjvUoZ0d7PlIzfvT7RX5ElJy9tXZ40wUz39Hx50J+DxFrwLbSpIYEx64F1em
iRzIb90AFVz4KphkHM8sFEa0jXUFTI0qTLkULiMCWzfAiPJarvFQYmtRBVtJ8dJxBQelauEbT9tP
/xbS7HmqdiugEwZNT9iCsOwdZgUymSJxPlnRxyvlFrChH48Vqz5rnxSvtIjHSrl5pWwYwq6OfFYp
80B+OUoiGdBohtU0CPVeXG2fef4CJAbXPdPGTFUX3SE0ftgmBzvfTVgKghk6mwWFFNLYAR5hZENU
pBtzEQfNMfe+VwidlGY6Lffbg9acpAl4o7wR2f+MTuK6CfcdsysDZAuGxG7m8fDGTyHbah9GsxzN
8Z7C9s1Q6sRDS8wE1o7z/Kkk18zRFm5o8B/UuqMP28YBDvqabGjoaeIqwsTmaoM3gsJvWQpsj9oA
Fp305Zcd9CFNQeg8XO8TGXtrNBpfavaVMAmrKAxwMMRywBupKpkqVci86qLpCqMBJO0TMiOJu2A+
HEqc3BGJKjsUIBkMfm82uhzpJVlHblIAk7JkjRA0WdiRoookLsSJTe30MUOtdidMs4nkMyk5x7wW
kPWPU+azs9BtuAxZPSfH/ogKjltKv5AcoVSkjMltELA6fqqN1wQtgf9Ivxw8EnvUhJ1up2GvHXhc
r/v9QOGAGRORAp0SmhLMjkaFzgWEti26HE0Log/JQ0Xb7C+ZWZcr7/YDTuuY1rECNU/QVgqPrA5C
DzRyG/0AWyhJzSNwX0IbUuhnmC7tn7+Gjn143LCSCLJz6QKg97s+elitSJ9gkvFqWkioKLVS8Cnj
dmwk+CcU3cYca8J5stNM4RyYtQNVlFd6JFMDv+S+l71iEsUxbwbl+5+B/M7imk2Z7LZrnAYgGYTG
7w5gHstvOfvEPYdeilAO9hCc7CB6ptTcpI5MNkkeRbCg7ZvUMZrA/0MnPWqX0JAqJ7Te3fYU7wmR
j/VB3tfpGA0xYHgt1ZM4lrsaJzcgh9Z2NDnVjaJ+Id19v9zGDt8n4cpFFpSaaVsLupNWk5BkxDHG
+KOnXBHB4Df84M7XUR6vXJwutM2rx1GAlR77hWrESbOzn5qAvp6WtExFkbmg/shK0LRwEKCRZRSn
9NbPoRfkXfH+ly6A1kowOQuUZL2xblsroXUrnqnaJE63HOXHIwe1BgUe1SsKcBQk3p58eR9MmXIz
X/EdytD16mxpNmuy0yFARvtvOK6cuVW8C4drAyuTN6uqtyhU9MVDZr9Uan3o0mK4C3X715BmpoF8
q/R6pvBe28o140s7LT8u77AgviVTDV4c4EEeI41u9PZUFMiisibEtitrMckecWTMUrX4dUJgmGYJ
mxTvMbXR4bUO6yiQdlMNs/LSy0uD5QY030Ql+ng29haPotZoHikB/e55ANlz6LqJQwrRPVu98bLk
JpdQ/CbkXGeoTdzQIEBrvKUHyB5f+hGPITgWzdU6BVvQVnKkVWsEEwItmPT7NwBqO6SD1PV9YtPx
d8Br1k+IzGeyuqEiSdJdNsm6OTNIvVBhQ1K5rdyrCGbIu8nNm34FY1Ph1RbYs7fwXA4C2a1WblqC
O/GTrDv9o6X8DStDpLyiO9F0NgFF5e2bD9a3SYX2tGZOx47hyNTZyrbXYg40iPZJinsAO9h/pWZb
DfXGm8hRh+U153QSJPyapygARjRY49M7SfCigNHUj/new7saWGaQkZwYY+zw7JPh2p94BB1o3frh
nH+6hzH4VpEgjZa3wN/uDUkK6xe0eiOPACKK/sYhhmh4RQSE27apajZCyXcPWSjbG5HcJdacroer
bgs8dN3HeKuFHARnBCXGIbQV4WZFQU5cgZqlbANTU4zo8o3KJwaP5W9NTMgy9+4Drv0OUw9iBsW5
1XHpRef+WOq/lO/qn6s65P/Lf6OmgfsrhQZ+cY007rQ/AygxA9uubclwu0iAx1LFPBA6wC5oZWZr
WI+1c1rBtSVR6xgNfeVQn9IKDdIRp/Ol10KNHe0tGktUbdsYy8+ecMjTVtFIzPA796igfdT7AXBV
jFGLHynoOzBs3gJST1D6hJGCTFJeVI2QkThSRKqbjPijjGmVeyBeLvHAG1xjOsi5lM1m0pGXyx5O
AFIE/uq52JrD6aVCgW1T6yDrSroaFXKKqVdQFopyEB24mPCv61cH4xOVz3S+eiKaGhKha/3hnR3C
lt9g5Vq8WKphnhtWWZoyz+p8FZA+DDmUGXo4Zy7bXkeIpqwlQf8on/JTna63ZLITqL5eBVHqj9Ur
Vv6IvUFRecSnyfMFKcKzwytwwrMKQ8CPETyxDGV8YdRNqik4eqddq9x3bcyZXe+rO/xBUTXj5i+Y
uZ4HdwtT9c8oMKD5n0xe9vfEEbChaDf+hYRxfnXWsswTwV3Wwc0KSN08HVn0NzFuYBbxgOY7MjEk
RqkpEbROnIkV2NKBkI4dNL2+IluIm1p7sjBWztSDRGS7aNe8YOX+NUI8f0g3XGtdW+HbQz2dc3Fj
P6z9lMlpA2vm0coFRBkplJ0gVthSrWS/V+h9EEm9f9QBR7+Crd/HiOBoujtnvWxyUVV5nSLvi8zm
3FO7JticeajyvYGKJ7PpzHXwaHOMO4UYP6cuNsUxd0LoEpKEun8CM4fVBED5rzmGyl/39qT1/K5n
1plZ4HorWea2qCo09/7yDApv5bx/JKpG+F7qwHfB18WjKvtQZGhvNMQAM9P0lAaa1on45ugr3aD0
wknDB5qQ6ALl/icTKv2EEybDS3Xjg84z11hTP+uI3FkIkQzxOSRoSz+6gxvYwnqRlWo8+AanwzQ3
6X2uhIE4d8i9X/Ja+YOIkDqwvk+eAwWPa32MmhAEUGEZ6gkAJR5ljLgG1RxTORpn1a7qXq0oASIN
KIkUBebOscD+yI/SYfxv8cqXfkKBVd++BQ3D0GhGg/LT0ywS9/JmwMxTVX3XcDUigw/qbEWuUDCr
EF1ZeJDr6z2khf9q3SR8gWzysz3Ciu1cBm9/a1trtWuiH6z52BUl967hHJchifo8WCMZv+Ow9moa
1rMVzT9ztSwS1MD0TFoiJpzvgH1A4/X0bQyup95oA3/JB6kQ0ladSib2js3RWSOgeQ4PTXYKpW35
t88z4dCoAUdkGvcW2h4+b+9IjJblfm9r1qyQbm6P7zVRmv7TXyC2foeKCk2HkuHwonlhq47EXYQS
XAlVReSfpDhlGvYM+uRwVh08OpzB61DkyVAot7/FAe1lZocTDx8oPkAaQTOYHh2pORnKcd49vHg+
rK+3qZsdXSU4EfYRDtOncbzaZ132wGoY6VFadvz8FJSTHgNWBI1xn6YHKJREqOYJhjlfycUTiEJr
M16L1kzUSI+uFlllqM9mu/PYTv5G3MIvSmDbTcOeyCrH0UTf7QPp2Gm/7sJQole3gaDBFqxgBFcl
YkSVKtVX1ltFA99kHv7OBl+MZw8KNU2TnpdhSM+6WuAl0apJjkceIl+rW05T8x6fk+XBxGKnP0+2
rkq6nGuAe/qXKDlpaEJh963TsmzizUkjgPxnRsn45dhmF/D4l+n6qu388BcF/X3MMvICcW2TtGLe
sXKQ4jsdXEUvs5d8CQ/5bZEfnxfUVyi0JJok7kfxTYZtwV5N0ZfNkZNQ7LLXWgWsbjZpjJCKRh5I
Zt4elGFLpUc4BLimUSTVpUOnHRz5lUclGu6sRA1TcvVJcd5gSE/g8RFIkesvJoGUIku0H+9hzrG3
4MBfa2y8Ljcd78ngiO/LsTvkC163v3bII31H2u/I/436C6ZmR7BcbqYPKCxEeJ7m1ddxM0YlUY1Z
h4MsbV/VvB5zCWRfLjxMWbKwJQcAT3XRqmMgwpkgTPIIfszv1yst9UnaNiatqHfyLZWRDvl/KmD5
1YycId/t2Kkl7yN+2Nt+b+4b1JAa7+k3HQp0OIt1DnqJ9SZZXg7Dn2iAOu6x9weCnRmGZLic0A+J
bBsmie6HpOIdYtKlguMhBDyB/Edlxe6LJPrJZTQxYwDynJ81Uy5EVNGj/nJ3Z3sNGgv7157qGXaR
ASTJadoGBDCztrkbCojuVIbRxyw4YYG80MvDYdZIsqTx0iLExLSUQ3CoZ92Z301TlByzR54DiIAB
wV+EjBrc+pnbRh1qVrxLenxZ1yHJQ8k9wQfa8Qn0msX+09gf/Yb33TMvVh4eieAjfA0uA2tXgdOl
JF4VTvu7lMkAR2tX0B5KWqcIMmYqyvOBWeDQvtDj30rk/C446In+NB2rwZJxeq8XtqIxXK9472jT
LYZ8VOa1rgZG39jVJHErzsm4IoeOErKUcly7WgMuosv1BpPsfO3o6sa3F2wcVZv0ATEiBU8Y2brd
ukmy53zGXi4HyUgKvy28D3cnm/96uytGnPPLJVnYFEa8zrhw7PLs1Kb2pqFBA2FbVUJkcPqFoWWq
W+OdP2qF+m3F9X/j6vZVXy+Km18R+xeCDUKrPrSKyhZF8kEGfCyUNfes3ysQSOJ1HCtaCa95N/9c
owxq2SGQp8lsA5HZOijINBf1QRxqtCjoDOlBJUatBNoz7+vsyVyKYYU/N8sb+WRkZgcVZAadHxON
AcrlUAqzUU7yG0S9xsURIAAB17gApt0M+ZFgcTHJXxmm4tEmjHdmrKI/NL+j2ItNRH5M1rAg4S2m
f0a3qLShpLz6ivNXCnJ0k+mn1C5LbXGsZQ0cb5Z3J5SUoOALgODoualo/+y2/S9CFa2tphZBNT2O
hWhGtzkanujUa8Z9ZUvGpNjx9FRVcAy/P3wnjLswMA581MqF2jo8sbIb4IjcJBeNOZvwzN4UMZhn
NV6ZNQowH62lP9YfBfr+KxJ1y1eC6inyUJ7Gui4Jr0nrMYBPELoYKifDLJjZkfh/0qhWbR0OdOS5
LmsooHKgUq5MdeU3q1Qw6cEkLJwVx5jzck3Srf5VtZ0oQFTA5FF4AVrb1UZrczq15T1uO8c6Yusl
9jmn+riyayC1SBJ9xLpdP3XkvJAYt6vGqzvTepzmJsB/M5sZgy8wmzHE8K5qiRil0F/l0J5Iyw/p
QOixdD+5wtyzlaZAi2xDYxk582Pd6b4NEJh25LpnX6EguVrHKaQvdoo08kz//gC3y7Sn01H7dp50
h1WXgCOBnFdnR2SAAG58dBKZed+FUz4IzhsWyS1gmkf+LETpYJUSIpU+u1brcMzEWdC0DUaGNaSF
SGnfiHCcVgfPA2cqnW/qs62EllU9It5pclC52qwYxHud2iL4MLMtO2WoBwaLw79s+i7mp8t4fPUF
dG32+eTvHg8COFvgOScZW8dVuywNHrpER3ra9YZEdfV7RL1FlqvdN6OZAvykHbZ7Lx8RHGmVX7Kz
6kMQtEW9WCNNPzjhV7F8zEIDa76aL9zKFW0bxVjNMG3eRltsgquPvc3IYulYl91LwszSSqigUVeD
R+IfmRztaeeNrGdvl6PNCeiH0zlmELb23dt/ctVP/vVAt397xKAVsZ9s4poqBgqVZpDI6zmbFO7l
8Z1D3iar9aKWad/FL9naObeYDrdqpNfjeC+qb0sqTczTXo+GTwFOoZUyn7NGi5GkbcjV0BWN+MoL
gEkIUtE5XmS/7Q+Y9gh0p+BV15bnNiPT2kYvC6UBU56f4grtbmTgtr3Di7LpOoTx7jFbH8KxHVT5
JMYQHuNH2fapjOuMiyPg2PJ2iouA/ti5j7bFFASX4U6TZpIQChtBkvHG8B2FL6O6OuDVJtmqc3qK
KDwuAtrlKdBU06uc6WfXKz2ShO/7bZpyd7nD9r2rsNwHM7ypnVwtQ757dKSvRKx+YAx3gc3NgsZO
VA6xnleZTSOqV+zw/2yAYCt48Gmo2Hz+bNB9uZBZd9Ki2JsqZciXg745F/VOteWxAnCVcqy9lyRe
I8NB1F3At4IQp+zHjAVzTBAP9gjc6G5cs2WbmddRTcn2BOVjrMQnLIV71jNMt51uXQbZFl86cIrT
La5+RmkxpPvrWYIMmQZZrd7ybylitlhjTihlotk6ksC/sf6aE9KCp+88ysgCOyi2wZfm9IqghS6C
yDUnb0m7yeYrz+GPdQnV9oYKgq8NyDPXa4ATNI+DFYSc2QR1pHHSuXxouOkLWtvkOfi1PildoSlJ
7hnTob1IwpDXPtTIr/eAT+QdQANAnbyiDKHw+3uRKrbHrIYBLdktfLdBvB43ZLOJtWAfu70bDhNa
EGD8sePJmVA2R/5mk4Zr5V96ZiUreTWrv5gteK59pG6mPgtqIS3leGuTM2ZPReJC8xJRy+lVvWAc
W/kZGYJUL+H4QKnG+pAt3cFlu1v2Ye9t4q1Oaj/Z400K7Q9AZWSSxl9ubjYgA5UKJtiSGOYZ2tpE
DgMGcNdoHvwTOm1Q71zHpqjdbBZkN+NFSi1NMKblQ2051cBRHicLQ+sxyiyc+EvBHrCgQ6YCETp8
3PsU2KZU33L0uobS+9Xsrf7zp089Q5hna/SFsAFYXgoStd+VHml5KZ5U6fjNKGQWBhnAvPMC/B7z
KTmjOd/OSyjdUfGufOeVgs6BMCitMmE8+XUfy1VTEPqgsM7CctKFTZguLLs8zursZYR0ZTDlVSJG
jYGjWIVS1/l+tIRM1E3XAGZsEDlfI1LWTxazjekfdQJiMBpS69g8G4Ke1IcIBIcWDAWvkE19HshE
UYoYHVldFXc6W5aXfR/gt+eUuD/pLzgOs4lWNaU4EerBDkhM5OWMXaIQjDJimmfG9wmT+93O4hV1
bIVak5ZovXXn+xf6AoIToEcxx+tK9wGFbbzUGJ8QUa+kmoDZC1zPerBDRkvs1sXtpcLJS76TB3aj
rZMlJBGhYc7JAl0uCj+IAHfWZ7WoMe2Zw4r6OhJBgQN0RKXQP+QC36UmCUYkL807UfRnup1E9zI3
i5UcrkzXIE8NUsGclGoLNr6kwGKgTPaRe0w7c/5bXjaxCtgm+lRsx0A8EXsyenfyzeQw2OUP5M2C
1eO5EH8HaF2sv+gqCU0XJRq94nMGUXgWM5RQVzjbfonp/BxoXT1DoVhsgTX1DaNwJVkZjXmCsZQ8
f/7SKGGDjnbaM2muUglnMaHkP69KaDRnijxAhk8qOwk3dQFgdTqA86n+9wKHLJZF3rB9WI7EhvuR
IVpJPU+58ToQxNBcU+5LgTYMVTgNBFwk0s7dyqUIG7g2jB6ldA1AqEHvrtvQQekVpXTzJLyEZD7c
sqstVTHyMFbmwznzrtdvrISZjOO89z1bFvrnxT3kS0zfloEhu4FFhknK0JTb4ka+ufhKXXNCUx5H
ZioWQlnJRKGxOG3D319oCWzFOqtU1m8BxOEusYNe1wnds9qrhLIR9KLD+WjPQX3Q9bvEJTG5xsm5
jikh0XWMqcpJnvchGe3V5Sjkwy/NYEGrTV1Y8LrJBGojLr87EBzatMrdaMXjjxh2tWHc+RJAu6oQ
1M5som9mlCsTn5U1k3xCMB0qXbHSEcFgC/al/UGLlovF89T8j+DevUUL99FDUv/EbsaGkXXTAvGB
6+G4RwyZrCGPMe04NPB/Uro64wicn62Jp+SP8kJy/6e9ouAofG5G2RF/HjOd2kZsMnPIvegCqas4
NVK1u/Re9PTd5jdBIjXDDOV+SYnvC5+N1lHV20auxrHWPyoXm+n2TYa15kg2biniafEJ3RP8Eh9V
8L9Mv1QiEKMiWpH3oXEBjVRqOMaGuEtB/eo2wyPNayfPYnXGhoWyhx7XDd03mJE8SROqPygINUWU
1sogzpv8F2MNArWyQfSCHNb+hcsh98uEmRBygXzg4bGoQ37GeL/KCwebJY70WiOd7AlyxZ6gzG3U
Ph4ylDAgIviItfxhEpePzcODCuzmbt1BF6y1Awbyu8Jt2++EByBevBkhWb9dgnYg/F/UPZI+k0G3
hdlUFSYD2YgdVh4X/1erhvknqVdDqpWxMFXfQW89UOvqU3YZortPYIhrh+QHPLPfLUM0OHmYMbKB
2xsSgmP2XMC/Aie5a/+QCBxXwGHrwa8W7NkmQQ9QWZnSBZuXs1ZI+SFmD3QX5IEEX3N1rA4OcFkO
oIK3SzJg73rQYKOqfMUm5a7OiD8dJNglqe9vsJdA+dXaqzjrYEspDahcgxkEL6cv6D2e9fcQyKo2
5AYJHO9YBziqaB5C8gzJs/VHIq+qi1Z2mQYBscAHj833LXADLsApNuA5ONDFY9eHd8X8HIaqZTUB
+ejvHiBfwgMfBiQs7VaehIHKd4acfi2xJ46OLaG157eogAaqEUNQC2/83E1Jfb9LteVez5v9hLqQ
Tv7VLglVDmELf4PEG10B8fiaXmtiLxbgGQedHanF9XYZYY3YTOoUYW0pIk2surKoWXuxVKCtHCmx
jTmwvuAM5C5c0dMDdtWdNhR8xwuqjPaImP/Zj1YReegrIpgwcdjPY02mqJu+1WZfAOxjcbwL9Hl7
wc8zjikcNUia57avUKLVezVC3ikmiMebAGKMx3Jf/ZgHjcEelRFHp0GjcXdI1GmPvptVRQoU7by5
jzFTQ+uRLLz3QR6iT/ubZHpa31OsOPKjpZIAU7h5UbNDokoOJCWkhnsrKMSUYpkArff6r+hYLqH9
mnrEYp7plhashzrbOUx4rQQy90AZR+sDMLqQQOppx6PKD66v7aCXXFv9vn3Esg2ovZxCx/qobFY6
fvBY+ZAPNAiv68FGWvX7yn9m+YVr5Pevx217A+b1ov0NxzEohj3xDXxtKfQxV++loyyZLCbTtFkE
vVOP6lCkSnz4WITLullcBIzLtUjqfBTn311YbYOUF/w2PbXorwjfrRuPAsBtflRa6I4uinDUypvb
RXeknz0d+v9bCo3+s3a8Fih4un64yva+nRnomQs3XpQJXvHgORr4FnGrjwnQzOchLCYLvKXFu4Z9
HMTHh3Pr6L9/yScua5/VpNa6B3NGIWzu6FDaQxw8HE3zTuOi16WDvk/zyI4VnPjEOH7b3hmmbeZQ
PTTtybnrri7i+lMDvj14K6koWrSfb229Lj+ZpJak8HNEsTb5whynx67E8reT9OoiWF2y8O9K2/Xl
ezb1mGzTftjORAMssvPIXpCWiDiHdZOvYG0qR9U4UKQtETjPFqJ49hS3iCXgmCGTmuldblvMPqJl
2mlVbFgBiejRWheodiz12Oo8qCHP8UCI6mB6z5jftgLUZ6MDlvKjIkJN7uaDRy6/1iGv+J15WZCp
KZ6PfYlc6mBJYpjtETYpHGhoZPfeVg7rkdfJT/16yPlttsAUkaozncUJN4yq0DMjB9efpV2M4S4g
9Tp7tYVSnh0SnFyfsduM/e/NUv0Zqyz68ymhoYohlTKn45Vixtr/TYQEzaekEz7gXrhAr7AbDfFp
Eu9G4kThzgRajYZOToBJ+LdPnyTQPIe/qKwIiC/zbG36TMRVlRiKLz/hA1qW8gs/9ISKjrAQaIPZ
l/k6Gj5sM2niLwV7nyk/VWRR/8AmpdR6oPE9ORatAWsR7L0nqd8GuRHVITLokpYbrnPnuyc0nixL
zjeomfnYTd7HOkLyRdPdkZmhqhWk3ia9/KXMK/sb+C4eVkp4I34ni6+2PVv+ngU0cuY7z3NGfuDy
QSUw/AEa0x32xnXrteULjQTphDMvYTz/4/LBydCdEY4GXZ4T2bjtqxVULdWepMHZWyIeyWfft+dM
EXOptNCs9Qn0uXI8nCGYL+rU30pRCdqwtR0/l6tzG2HSVnPXyilgF/5dXHrnThTetS+VrgmLHdHY
4HUbWjQTwq99HwYOGuSynCaeNz1W3CzT5EoVRhvV/cpXzun/6MrwlifIuUu+r2ik+JPdzQJaT/Ef
18d9qDvci8H2KG4Z7+hYypw488kZCc/ZaTlRmFzy7gZz3hAeaaJszqI8kS6E8GPNuOwd4JCA6X2g
PIi5U8eobW1ojIRUENxjhp4YxXdxIjHhX5Cx9FHeCJYTS/akwJ99ABBSMKg8QIT5EIzzcXJcC9qd
YtCuJap38OaqxW5K2zWdcM5eoBf3c+2neSuOIJoNia8WNJ/ppJVE9bLuv2acO4LMuAUW2D6K+NUP
rVnaf33tI8SApGzITli2aeC7akaQuKoCmoB6TI9Jw05WiONP/x0Ub4jY3g2yP4yUZCRUpKZo8W3P
B/cK+041sb8DT9kDq/J2rgKhBYdnLkI75wFwpyl66tsURFDcmPqo3+7+us1QDjOsA4S0rLL3U7ne
Jiv23R36oMVyiW+tXg7eCi+pYBNpiO9jruqLIxLb6gbOxHns+HWSZk3ItVMB7jJu/ajTi0DmjJ1x
qOaTQap+/BC8NU5WN6PZ5Jw+Rj3StC1UUKst506qm98epQUkOgebOteWqwNyzxnXaAKocojEEbWg
/DME333ZjeHMgJVmOYLR75tqig8Q/fmbvphN+NyDtmFeTsjtQo47bs6KD4LeS3MscyPCOhnCouiL
djxt3w7mco0d80zOUE2ssir/EzUWdODQ1w/hHZZbGBNtRZImEqVG1F0VlXCpEtTkLLGuikAClNlH
RJmVwTULzFoUxKc0M5y4LqI/l5P+LAtws0NxtHhZh576nOC/zktovm2ipI4ijMkneh9qTRTnGEFt
H5PSGaqX6TrCD9yBk2CU5JbxZKuTgW2krxsure7ruSTQrlOavVKZCKsg5pKNChzPVYz1ZAcCEw9+
FT3+x4PqQCO9EbqUoUlFBrrdb56f1geQyImkOdTCLMsSSbEeRnMyJZCj9meh7okuEfr4NvXK8/lV
MdHCzkygzALmScaAmN2Tyht9RSmt7jZUoHkBL0Dp5WSNcqaFtmLMlA5omenti2Nei8hjoeLd2Cjz
H+9MCPr3uZBRp3iaH9/xOHF6EJ+ECsLaSxcfNanOfBp03OIe1jfW9cSpfP+gGxUUbVFslVl+QNxf
7EKL1MiQRV8PnA1vPJkB0GnmvVlcnscIdLDhpnJ+GiRq+Zit1WaWsT4YQgZB0dXAnXr9N+hZODcy
JOiPTN1yJXX9NR1LA+9ou3QmLEyZVcpx49WL8JcRW+uO/q+cg9UbvGiaOOKWW/BWau7YlTj3Fz2U
lAF5FdzdFks3JpwmW6CHwZvXzOGnnXKuNJKsLT9UtogDG7qa9659rqMzZ7Dv2nYaWgEUZO6lU7fG
fE9Z+OEBXVOdSsnrR08qKS9xRZyqyxEdO5ZAFSW0X/0sCWcNCg8lh3DzUC3Fq4mQgluwBTb4wNlU
ZcsF5Q8hNh7uIkQq75aVQVZTC5PCJ46kNNBYuXUxd2S6NWdsUBSJcM+ICn1rosWlHYgBuafsiqjB
UjBB38Vl7+qu1UPVb4FnQMnwKYRuzyoqecGScvLCGhgYWCz9JiczKD1xkjL68rxPmHxO5rJ4dloT
dl8lWBoopR5RCG2sGb8+ESwNnc0TnXl71+H5XCqAhN600tcxTZ3UrP+8P6J4yqYo0NEazGdLHdns
wcZE4GBl/dG/OxkisvrmCTrUCK16QICPAVm+a4k+4e92hF6gWhQMsduJmIBgGQeLk4RhnrUfSkLt
nIoUyb+lYiQv2v7Z//KJPDEDNHZdGLtLoIOwOoMMBmlltMpfV0LiYaq+B69HNN7QpUMXmPhvufdJ
zvNy/6hZeSB1C8g2Qq9qwgbo+/CfFgDBcudXC/Mb/CecSakiJEUhyiWSkUSVrubEe9n3ZCKuIo/+
t0VDX7AAi9fg1qO7PLyKXNcZjmC/9lJ4QmNlsRlfjVzGoPi8y+PBrR09pEEIXLjXogL7AtmOyvPO
PrIVka7/y+jTTK+AGsM76xhel5F7Nc4riC5MDTkQ+KCYlNwVOQyF8GbvIob6JFjtJsRv2T+6gFt0
p01Ce7z3fxOj5VEv6Hm0pTdUwfA8C+I/XuK76dxS9bmtZkLyYkREkWVpeXmFqboyZScTUaIZTkBI
3lo0DU3Loo4JhKsx/0QRgO0ZLqUGpcsRfQb7+nVHX/rJfxTgtzBbNZhejZ1+x36fA5boJ+t8NnNb
P5GSJc3gyt6yyiIEAtc9d1RV6pdFqf94GgaeNU9K3NK7UYUL1/wJcdJwe+4h+2UixRG8ibvJNExj
fpeCFAs7Xw6qFv7mBGQXmAZvBbBqtzCTDuaZcNc8J8wJxm0Muv/qeyvqAk9auBKbDH4ci1yW4JDd
xLjJcGM2U34JTnjj/+Kx8I4Ez2FWVIMla4PW5h33IWoQqQ5wY/XdT5ovoOJbVpXSvuTtfkwyslVq
NBaFaRlypdIx5H0B2QNVFLo08irCuqj1zXTwWE++0S/WuP2Ft4E0hnxMG+uRjTIoy8OJ9skplsZX
jqLo1CvzRiB+4G5w9F3B1+T81Rn+1uMQLJN289QQwwinjis7Gsu1aOVC1g6RncWF32ZCjQY7u8Rm
LZG/GInFpNX8fQ3rmkNXMRbXzLUxMw2owvcNqzT2bvmU3HNHQ4HSaN8gcA3Enz8vJTmaFN4bCJxe
mjifFB0fNxL4/iolT/8KORODyCDfzDYpFHLAiFs7TS23svzGcRaEOBFYIIEqMYC2oabA7KZZxUgP
ZHp+PNGtKFyqbwOEeRCOvlm0VJMvC4hVe/chpzBQ09QIajGn1JRwgXmtvH9Bs6ehLEKXAQ9aMqui
76Cjja/EnAv0gWHWuspsrStCuWVXqLZ5P9rNuh54PwijjUwC8PgXdaakZojvb9KYeILzejxRxyPd
6ZSPhv2IR/M4fPsF4PzwiESbiSfKbVAi0BWOrom+9afqVeCBpLogA8IYDiIRfVnDvOSCLTH9Cca2
eHd03ui2PyEzRhZnGoenzZFsJGQxKlQZo8JqIUjZJJf+QCxr2CSlCRmgJrH3QYeL1cKgPUNkZxPY
VLNrplgDxh7rNnaEVaZlcvlbt+9+jbVot/+aOHuuh1gyNCfr/Biza4sWJXhwhzAFQeBhRzqo7fUL
lknbYsRbebvTKqgrXXkVyx8U6vKaQIvHxPnmxdZ1BydgoVZRz7qYpAl8/vaCfBLr1OfNgxLNx9Cs
I1eAm+YwI1QnKbeQy9++r8wWWkA4UE447dj0e1H97y0cjGozYi5HkPR/rK23gyfQ1hYKq+y2/aXu
+AUwQPaDeFXvi1q9SyjAy8a8+htTQALHncjPkGCyPsw16UWxD21s6m3ZIFq+NaLqUrEKuFKxTt0c
QTT/0RjPccXt4c9MWBdesiSEu3Nf5eqQp0sjtkkm7h36WqXR6yOnBJvHHjFrU6hIR4Iv2olXfjOA
3o4TEvQT1Tg7Oo/aLM5MGldJ/nuHwpjBdXk80DTFHjjX+U5+5wBTGCGVQgywvgCUX3BCIiryp5Eq
xmHRo2/eIGexS77S6khiNZZC2N7c31kj4gU3Hgba5p5hsYxt8GXXe70JiCetR7+j+iA/PEAWwGbq
5i06dKhrwXHEe49IsRyFp63vTxdCRyTRURVBUMMlIpuDwuoobCvDhUBTgAdI+ICidLcdoLFgJgQB
pYEH+t0DlJIxjKvyL59lChTZ6KpktSjqFgrf1FHIAZXsVQ7KTHYD1e8VFB0b/v5jytkVc3yTs6Ts
jgKn6brIwcivumHq4llxnTQxwxIrmWQRr+MZ8n7vZQJQOf5aDNACIzaY+AEhZhaLkb/RDBqNPIsV
niV443sZx7MDUWNYv4PpYcerSihO3ZoMStbsPVnMi9CdN976UVWpHUuTcUujZE2cFzYaBZRJ9PLf
bEjWA8fvoaMO7pMeQ5FPzm8W273GYfrCiuZjf2yRg/ZMWkRW3o3BX1ybnL+0F3GJ2W1IcGddsB07
khUNUUImjf+dudN8H5M8fN71j2uIpJ49zl/ahlhVqz7hvYPZhoFmOntqgk/zWHVZYw9ffDHm2g09
dwjI0pTvyAZsxQ0jRfn/6LQ3xAlq7l6f5fOvmd0rIvB1mpugzVigqmlCBzCK6lzIXDXCnvrFrqL3
M5e13nRxMg/rEW6KzNL/AmB4MKrZkAI666zwfBOobuCm/FCSVDWhzxz9veRs/Os2cMCagrnFduH9
xU9a3xyOGbjcMPmBd3L1AA4NTLBFXzCkBGIoCtiRgppS4zrXtA/kxKyF4vzGjyw9EOJjATejq6kP
Y21xLSrGOx1xIMjIMaxQjUipZoVXhqsWktx6OJlPO5e1hYGddyMQguknMMWILkFXmRTthF/7quMv
pW7BhlB3BypHE/tG0wwYtnzZ9sh/fxokz7J9C2tYRnrFLED7lnUhw1KI5FjlRnMS9u0XXLMVCHKi
DU7vB1fcpuPMmhS/MDNexMu9LLp6SKpnXf1vQrHCB+mW1Q/7R7KQcGyF8+8BHpXten+I03iF8cpI
NgvMgD9KbDOpu/gtYF5We1U93OQPQA5OYSOE/O8QhGjpIFQ33j2DpU9MxUW+859Fc+LoRdBCyoTA
5dyHZNw69Gy39mCxjy7zDXXjiQiPftJi695Zr4sUcJ7Nttw3rXATolg+1IQxGwfB8R8vg7OutSVT
iMbPoop3VY7jC62vV1ECrZP4fZmLyGBmhpBJrmR77IAbb0uKvhOahkRAtZLsmfgtaXymfLg+ukA0
Xn1+fNa8ch4gaEdMC3QNmlILdAXd6/JdJzgunT8rf6d4Cwcmm5Ke/kE9v0J18V5vF5RSWMuEOkRK
rO02ETV7dMSSDzsZCraAMgYl668TQbMi1yqyINR7xzsABwmQOb32UpYxk5L1nHzAY3MWxnFaoG0r
Z26KTNMNfvpo+yDcsN8elduk725+249bMK4Hz9GqdFmmxeiFFUZV4dXYwvbdKLaz4Fowx0AXVsfT
81Ab9+jKQgCEdRHSW2ncmxWHv/QiW8fCmS3CBHiK3c3Wdw8nFV3f6/FXEIh7w/nHN5SBXKHl6835
MVG0Ai9RmikcKklcAH7l1iqT948+F8TjySGzRGXnizTjG+anAzntZtmyCVg4uYyg9VaS14Qr6a0g
ANf59SAoxXaNXcdQl+ehbMEjQ2uosZZQIDbYB2PECiDKVkN41BOG+whLEyy+IzihXlIJ5h5RbSIr
DKfFeOz1jUwUZIYx6GJPOG0aoUPMIQe5ELUQeqG+NPBUtsmENU01qqszx1bM6PFVZAlg1ZkK04lQ
gGpmhWgX86D/z3dmQ+YXpIDHrB4S/9g0gYoEN2ZT7uyJEWPLYat/3uNK5FOWEflts119poHUHeVj
PlPAzTNkZKz+9MUqgEwoxS2oxEni5tZDFVmkriuycI9YmXesBb43Rho9hwNyOlZxNrp3MM4BN9mW
ZAFKi0/y1zsqO5Mdm5qXeP/YD9yplMKiGtZMVt+I0PYqSkGp48d9JSwe7lO73jqU2nIswlof703I
nStmfy3mZBsglF+dPmewnJhpqyi2hSHiE+Pm3wqQV7QesuhjZ6NucXlKvZfYWiKw5H6duqvCy0yc
+IKC8bFanWkLsIEvynTEx+YoUvQo+n1zLhwm/01VntESIxkE2SoHo2QA71yLo6/h+M8xmbfjXw+A
1Yv89i+QYh6d2E+vFoQvXKUIzYnA42XjnGTbjxJ7/kx6T1C3civW3O3onqNTcnPc2bCozPAI2b4I
w82ghIlDxTriwIjn/bi8Vpdu/nIr/5NMka0lUgDIFUpnOUiScQ/d+Y7vhGluZZz81MY2jSFIvubr
eJer0A81immjvhgSrCN1lLKTiEZdgDxVam3O6dQiwGkdrYb91QybZwmVMOnvYhAc+B55OVNDA1Vb
t6IPA8Pfu5Mh6NXXDtwVIgqCb94i8eUWKZtB1fuOF08UagoH+omFSVuplmV5/cqDkpUVsNTVaDXo
675E0yPfRPgt31I9swKoEQ6hal6e9lO3PNc8iT2MYFCBdn5qW2qVpkfBTUOChiHxdYU26bBMS/5e
mez6OVb/2ajGSQ3JOSIZpEWUdxT8w7j7xDKDzGL1hpS+nMhiHt3CjnCfMuyUfBv9/k4CFb0Gvjg2
ze3lWsLk9+VsU4aeWnM/sPUTmIhrSijuNOPW0WkIE25CN5hYm7zFo2Z4IRIGRrC0WhJVbmkmJWQr
+JLEUHoqkzPvt3tqP4nC/G6XQPSrfB401rSgxwiiHg0PrcMovNBIk7YUL1SY9AJKSj9nAhhNABt1
88EiEFr3ipmZyAF+kxYGILZNxsFctzPFLM3RCOqCiv8tbD5EL+fzV1h3aEktIIV5cDJoO6bTbpxr
u4M2M4JY5rGhQzmJS5lBYNBly+di8vJpCFATg33p7GUmJVYk0QFr3JOuPOng5c+AJpDvdXBh9zKX
IhXPHkKR8eDbCDusxikQaCTY5znWUrQ4v0lN9W66lP62nV1W1qbiLPE9p5YKK8vTH+F1YsruuMIf
GFJMFwSez4aL54SRwxveWdCqIwDqaYDCCu28scHj7/+9ON31RqOvqlA1Dv0c+I0xu/H+rF/KWNtW
dmg3GmjDpv4VUPD0urKrGiyMyi6rDzlZYKUO1yXSvt3Kgbbs7mMjq0H92u5hUmdgDhOc1eYF+hfd
KcHO9V1fu0TnligXpqtLO3ppXSANui4CGmlV5DFwD6UoUm+BJq8tVc0uqcECPhMoDvfKL69/q11J
CRNnJ/Osf1b9hDGREYIYfCFheUoAoV+EwElS9LvjICP/eWhtfsjQY4+0pJMOrt/aeqASiJwgqTJi
q0X4BvjS9VyA/MR4tM2SQIagd/vInPiBWoT8wvzZwUw/1xmc7SSBwrqWmiSxkMp1cG9S0aBzNITB
AlGRcoN9TtsksJSRNsCA9tsa2qYfQysgQrXF2DfD06XpZAPR4YCSfW0AHkAMqIBuI48jqDE8SCik
JZ+Ns+mLKruoWTMgpHdEfC22NiilfkkLFeVxDR4xwQcrNAgLLNVr0YQ2mPcSdf3ARyPG8SY8v+2G
3wgAiUSVD1txLxipbVSSJhIBWlFlCbgLf+ukVDvEylBSkspnvHlgNteMijUbGADcogVYQOYSCeTz
P1ZvKnjaRM8/YMlSj/6EAYKSFC/5pMPzSu2ao5bZCRu/bqAMr5WPAHBjgSzZOu3nU+UNtL6a/W1Q
JOTcFRnhwALkF1G96+sxOrikgk5EL5mT5cD9MFGvrAZjnurahrsYtQ7I17hunpc//2s5c+P1TECl
wntA/PcPJsKZsZH/5+Jw8q0i7IYJ6c3l5yjQyoRaN+/na53jyZDGBBmM7FGX+s5ym4ETKBF0lLAx
i1xw8rcjljNGKTY/8yKfUW72ezgMsfJeISnhrjSyGb4mPo9pay8Xc6yeOmUl6M3zG5NQL1W2QBFx
DEz9icIOHd63hqEPL5UuUQ+k6b31H0gzvEJvT+ZTqD0fK2P6QO1rMIKD4FjtvoLxTyafA27OtDYd
0XhH77kMAJAl5ZoOwW+G/cbrs8VHRysemEmCFemTifJrtgEw8bxpPlupIWeS6p235S3s/A9A42pk
efAPH+RQLNycvpSx03juhHp3poA/fnzF+/D2sx5+o3t3PlQB3kPbc0mD7waNE6iS0CnSjpsyg2E0
uBRZ6lu+DjmeqhfeMB2YCXyHgqJxfKiXaLmULdm2vAgVerS/KDEZrbQ2nQ67/La9lykWmHHabFcX
OIEDU2m94MQiitehiXuicxg8mjkkuLazR/GRi93qvesxFM5xGSJ/ksLgyMX6N3Taq6GOFj4ZQVBd
YfeKHOj2p6AakADNTkQnTArymSf0q71o89i60j+l7urEoEEsWiODpILuTykWdHy1lQOwyKxg7+du
NmvfO7M7PYVb++h6FNlmK3m51/f2nKpBvz/+3GFnqdIGgXaaHWYND/Q7CPBchXuGAjoJh+W+FW+L
1u+qRJCrJH3ZbBLQjxx5zw3DvEfPZCRL2IrGB8yt1WzcIH2HTeq2MTy+9StV8ZlWGL0u+0va/aAH
oKsd8DXlUuJvjlhNae2EKsedctwZeEqoA1X9YHumEmS7xbddFTVc56VgTGUMbHfi3yAE8fOiAGTx
746cQbSa0MrnxsTl87y641H86T3JDzuPy4f7s3K1qW/MNQQMdBQRazttjHaTgZZF/akGl2OKNoS4
GiK3ME/1ZwCt7DBxEkM+ODCBfejlaKqww4rRUwtb8m+Yc2wl4b+sSJmlCcW00YsocKJoxaJcsvdf
tvYQ41CKxhyPMaGl+y9lgH1AmTetKmNQYwCMJnCGUSTRFFfV/IZbr1zCQLj2BwETNmyRgVhC0A0b
ZiJinGsUqTTvcuo5LKOGqoSTgILELRE/4Fk2EoOEUnpsntXGJ26/R4gf4Ut4ZL8iWzwon/oQg57H
5fTT00zox9RZQiSN6bf7scjGS/RqYi7loinPHOcfHa3+pbULZY6qs+cvYTxqprCwxtBmdBDes3v6
HZrnJTFCBW0UTlsPTVTKV2c4PK28YOqVHcDGkOc56ZPYS3+Jmf1VcJKNuusNOdZWTsrBDC2zIpu3
/FDpKnM9F7wYOLBrcJWW3nopdn6sE4hDSY8/NcyCwpypU4ocD0dDYwWyilW/5nsg++qsfoB5IPcO
OZGsKsHczbfAusQUZRiOXPOkkAiq1pf7tr5k5aqsheuHYMvES5y84kr96LZeCHZt/qx6He5o0d8j
CSfNEPDss0naipg5P+xgkqqcws4FgnLam7RYG8URNVoocMVgyrjbnixyVkvIriPhSvYO3tbJ50U2
3C4FBLPbtRR3TRrOhzd6I4WmfOplnULxn2ThuXzuaw13vp1s1X+m0B+Z6MOPq/nRfSqKxvftJGUO
+EvWHSccYcOvH9G2sbnjNxuvy0AEBPih6FuiCJoxAek3NE7uo3bYCXRE/rWBzO8zXg/DzShu9cLd
v3Ku2OOvJknLHmHo/hEzSwLbqLVzAsKhoFCQ22mDf4qiyTbrvnWyP/ZlSlLC27bXCiwAsoH4VcTC
2qs58xSI0gjJs8oBkR/JtvHwiRTU7nMhzwqU1SKBeYG5T44rvG6BKQIrpLOg7i2kAQ5xgEGyumTr
Onx+0Su/FbVcU4s4BEZ8Fx+V+Ezl4Jsgwha5zIe6dr1ryXRj+QxMUeZimjvTzeIOulGQqiViDxiW
BmiJs2dJ0i/ItuezYEHD9CZFySemt+iZa4YL2BRvJZzKA8dysRKsv9ewKOshSkZnweZ3I+alqtnW
E6hbb5Jb4RtAEZ/T4k+0uLSWp8kMQzGSaVyLpNB/8g8PtMaR37sIxj9NpP5QfKxqIzfl7eKbaWyT
KENirvDKVjq12rA3Glm/5uieJY/3bBH3CAxGSt1kYYoUJgQueVmY9mj7t0AAuab0VyIPGeFzfmRE
wkVM5ioQUDOk/sWBU0VWvg/SwkRebrVwqcecCE6hrHTVKA0mUxfAf2RbYfvpqky8TSl4yjuzvwki
5vD8PLjvH85YBq5pZmEzOol753yrW8KeTW3fWyLQoYCqVre4lC9WQ3ulrdlMYGkodN5A7LFIyTni
Wn7sbOhkoEKClZ7JNG1Of1w2p5/Sjtfoz2QQtvVs3qs3Z1C8xnoN3cdsdTles82pItvshT+HVjsD
MJ/dl1wqAPNKiaOv2iowkZ6lmMiot/VLe7iu6ruM7cqe+KK43MRw+8K4KcsT8H0qG3Xz7u6Zelzn
+4AdgUEG9wXi5Jsyr8XmEF9gkW7FgdKtJkfRz7lK4LYGLGG8ngaXQwlb56DsNeU7g4oFNDfQG1zf
LFthMZiJdEXwCXbC6I8kFsC0o78JUa8tXtiJrh+3DAK77Y4cnfP86PPvsuOu1gFYUhsHKfA+6Oif
2wofTZC9UIFwGW56u6GLQGvNjA5zWYlX3b+GYHRZufmm1PoT1TJWWQTcMkSGLc3OmB+2qit3hq2i
PM2921rVVrd3XUTICg4rx2RO0KXX4KV79cqc0EoGncGPiG7ijyQK0Oz5rKVjBZWTH9LAgJGDcfkO
bus7j+qeIySVT1zIFwM+BCUozEkSJtRFI1XWm+mqyiTF9fttU4k3zKXq2qUS5p9UwzTq0rWTc07g
WBWBGTDINKqN98iUqZE3DyKudCczkmlzqEQPBb4gbrD7mbLAQHfwUOCawz5FO31N0qggXj2XYnxC
zd3ToSCvKbPNSUdKUX28rPgG0v0k40DXV37k4vhJIZm2siy4XFKx/cvyeiaya8O+EB/5B7ksxTTj
Q/8lG9a3k/LakmrJgJaptE0lsGUgkfOnoovYLYHpVaQid6+bZIC6ejT4E/Cp57XZEySNRVUjvNVp
qimHiCJicMbpz/hps0Niz4o1ulQPEiyUZCSOA5dub7KxzAxbKZRUBDDlDxTwS+/v9VtNzzKEFKoT
5TVZ0FWOVs7xgocY2H+BeC7P5dtadY8uPJHD43tMQnyq12I1YbBn9LI9Pl7v2pyTPRhAlxuN5WnW
ReH8P4l9t/rORbCgem2pciwiJpsBYB/MoX3U/lHVwfI2gRMFLtbzJjUJghEL42UvvvgkHGzqZ4DA
GpCN5Qpi9D8tBIvm7P6qENdUnCV9m+pjAEs0QDfCJbwMIO0kbz82IVSGxT8JNBpfpfg434GxMYWq
2xCWbl3vcwsh2c4f0S5jB3lF1elwR9YSq66Ifb1mYSI8zxDeV2pyyLeJyH2s070F1Sco1yFrUbta
sVYs4/nXgf6y2dhYX0nFoBLJ6sNsCooUWQlQOnrC7HdvRMB3Nyn4KYSJ5z5L1XPjykWGGzK3ECsK
9xb29VJ+ileJ2QKJWlw9FJu62Rpmv6h4m4aOBbgBSCe3bBRuBJWOgCCsLxVO08Wr0dt1/WuYI9NC
o5TtGic45T0abwus2meMZGkBxQiq+W8M1+/fUMKe3F/Rxg1Y0q1Pfsqs8mKgflwXpOm9miYJPxzB
93LESkFltepeRoS3HrR726FbQKehq/R8gi9ihSz/ID76gynsv+6kV7va7FOs5JykTk2adn2aXrEb
9nldv9u1G8CDBg8i2BukLXKc4PYkCW+pjgbqBdMbKwBaflPH6laYSt41vSwBPKpis8YoE3StYDXB
NofF9C+oR4xj/UZ9BJOyk97fBTJi9YDjOlMkX4LX7E/WkLN2yiiXg91SZH/3l9HqaVCgb1+YVUpA
G5V/xrc0lAMMDfkb5Fa0LzJcTBDwvO3FWKP3yaJMb5Dxl72V9AyesJYtDWrlTzLXy0uMg5Qb0Qmj
dyfldi1IorI2uimL7wjELOJGE2mphmveNFW6CiO4ayJhx7fB+hPR2ATfa+6x2BsCvYcDX4EaV/+0
RlkAgY/+wm19AvJd8IG6Gw+w6kekE8NkEVNAlccuyXlWoQwJzssHu+T+i96I8XX+xK9nBrtw7Mow
QIiU1LA0vT8aJM/GwJzo8tvh2K8T4YypcPIPMcyDc1NWKLPVJDai97KoxGdcmYuu9wOdcIY8vmpp
4buQedGNSyPH2WovVL5a4+wYqQ8nTmmzTUFcY45qbDluvQUqg5K3BafBG+s2gflDQu1eZ9D3u9xE
6/HzdZHNcH5N/Ar//WWM3qSyl+tp8jr5NxHhwfOVv0K+YADq62VKLaVzfvULxWRh7gLn7VZtRaIp
VjOws7sxnzKUsIBk4EnpLZsjyws1F0C8Qa4qmDBXqKxnq08CQbuIv1ZZXzX6C5OAB6ToHDeIMGqm
9nurS1ElfEfd/aWwgPO7BJuJBMooEpZlMtMHYgOIkAx7HkTOt0g1REGhztyIBn3gbBN8XeqI/sS6
Sg32H5zbu3Ds6Z8CDeCDVXnIgH+Hwpqc2HVRV2LpVBfnD5zdXcipAQAgWfxVF1M02yzjwMQTBEah
p92N46vGjGRyKpVr7j62u8zbgaBqUN5U4Bi1AbigjcPZnjbH9BsHsVugVH4GfqW+Ciz8KgZ1UpTZ
FBm+ubBN8arghnY0K2EsclLrqADCU5+P61nIrZxJGhySPx6Yt1csk03hZj/MKWvYK2etZwwU+0bc
Ho8EUW6mHiCgnJYQdaUPk902ZW1wU0sIKpCXDB37FQYt27JqZHcKrZE+2egezRKP1AoSU+XMKtxB
ot4nctqXI9HM/LJ93ke6YQ/8gB0mK09Mw2DIg6zAUs7Orxs/W8DWaDLftPevPKG43sIDOBmhe1u2
7Hb+Vxvc3glFTRtS6O/KrSQTamFjAKMkNFxrWXO+kyzcCi4Bs8X3gdTPGQdKPNzbRPONvow7S+R6
XK0RlpmWOaqJkHxDzSACFl+5HZ3u5VHPj2Yi32gleJfpg9MZ+63dn17EAWmN3UZgt8VcBser2c9I
9Jn2odmsp54dSPTgc3AUEcua1J6/z4FzmUxS8bS+TJ48VPgWHwhOE63kI+2eDUr2nkuczz23H9sT
0WrEN0Trj7wWbsCPncW6RJ3NkliU6az7Frq/c/8IJNAMQWN+NrM2+v6OHWq/6FUdVXIUysgyJO+u
EXNrNvi4TOzdke9/bdG72RI+MsvdVc69TpFej/5f1MzUvXkdkeETBLgrl3VY3ukrQwWI+h5hikku
8XIYtnHYGAE9sAhIsECVK9A77B22YioDvjcEh2hk9ZCl8tpQJlv8PONCYU8NhFmM3ePR4TXMoSCy
xxSl1ok7B8lByxbAIfmPrAz9KFdFYs/gViPhz40aPDVKn0xKBUYH09Fav+9+P17X8VNldMDXUNdq
mzjUlPclHeDbk6ACw28GTJcqso6JW45dndjMke1CAr0qoQ/nZQFhTkaV21voB6yb/P8bpXbW2zxI
6diBZqJCNS2XEFBb0dIV2gGf52P8ljML1U3xiTV+/fmhfG7BQ2WPRZdVE41U3rhYAKqSxL76Os3x
82WLpqVo4IqQCwaeEzYZM1TI+nl7l2aioP/S+wl+CYc7EvZpgo7xEFBnxy9Z5rNNplO1WfR7jlrG
laWM3xpJSgK4v3+U1DWtDRCfGDfs55fy/XMUJ8c8mXwLoHuyvDATcOQ0TecfaxCf3vk2EhLk3f5C
s0ZkBtghn9yjcAVZ6CcmjHMCj0iEscaymYpSPCD4HnPtqL9OjHfL9zygrsvfNQza7JBQVAg6Nhqb
88enz6x0epL8FO1zQEkV5BvQtOBy+N9BardpO4PVLgStOEqbn6mYCipl+Tj8eCTcCMfiwJ/S1g6Z
mGnEAtg7QPmDKSib3seYsgvmTMb+ZD/BsOHVNuUPrrzYEAVMPldPNKpCdkLdX4TOaydvaXFHlZo5
slqWgyXuO6cKFuG8yOuIQgsogedJfW//jQK1kavA4FBiM3nmYftFKNIUy/sBVRJFOdnG7XUHhxMj
uSkFZesoI3Xj/b9J6HfI6yM5HVTWyb9nelNYkQUh8oeySnndF8+r9BmRe7gMlNuFBQFXooAFViLw
u6UCz+v6kBZFoG4dLAOXrrZMkPs8Hoo5SCOBSLDu8yYiD1WuAI0WqkyTnt3EV1Cq4czwYKTCaPOe
jS+CiK2E6ONgoTVo4CytLMppJOkY0zcRKfMYPwEX0c8jgsAe9gKx2XHWdJ6uCVYy8yFNQXykdWPY
wOZM5S3tNaMkkBNB3+eBgRxTwSD5ss5/rigj5zPWup+zZSjTPZ/0K9HuAREch4mqb7CAw6XwwXae
272krmfGLtbepIhQkEAmpSDXm+deNSs/tKNQPYVk7J4nY+twOkaJ62pSZw9nVBnXchIY5ZTB41wz
nK3YHicXj1FJkkmGWewcUSj2konyTZOjM3WJF2sJBlF1VstTuoaDRBgekpQn9st5xaK8QVtrqDZq
sNFnvJjoUrCtwlQ2S5R7JtfWw8hlA2McDUBftPT37yNuCvc9e4/FlU2pr7xKC3KHHdpOGXYD7+ac
R6c95+XbyZGWFLDemPC1bTW/2JbGioCNTgMt9D4IS5QNMUqJWugVepu8h1e0mJm2I6sQKzO/njXp
TT8N+exfC/TsgBZUomLHX5SMDug3Vf013eUvsfv5x3zuswYvK3z7JlRkq6SVgRbl1hZ8i1Afjd9C
UIIWWskX6VoioFm6Zezr49t4RJ3gmIHBEl0LyDotdtfPK2KL8b4NGAyS4dBzxPtfRz7CqxTuL+r9
6SCec1YLjKrefJPesOtD4UeiO33jeCkWJqDlFAKsoMyFVOi5XD3cBTGecyHrct9/HMRUCmYdnoyi
mvf24a/kXGaX3YMtN+VhwTIzwj8ei7Zz+rEs0fXM7s4hJzriY7gvyaZl7nrSe0VIhNslaD8IFjxt
OkgjAEvXTUo+Dp1/0GYCvPSChsj242UHa9sS4qOE2PlXAVE4O0mqT78+YpNDpbnsMkutWMQ6cZkn
Noh806IJ5ejxu21xpBh6VmvtJhkmGu0sd/5FnTeMYglpBhLNRWMS4NEnUTZYEsjvnk2RP/xgBS+Q
lDkNdxqu956VNhuR2LGg+wx2XX4T98D+0GB429Ve29Cl8spjNYKltVRIrVDZfac5ACWP7dVnsmQb
plt/vfjBdb0GHUwy+dD00jDFmBQPE5OIUt10mlnE79vecDUWU/6azhlwixrTK3+Q0nwBlkK13o4i
COaC6n9YahiYkN0BlBNqIMJApY45DJkyD8l9uy1vK10YLAbJ4njWLG4IHcoamNNw/Td6/7kM6j8S
4QOxEXh/asOwSelkwIZo5NSVePZhJcND6SrX3sDqFuVms19rdpD5PT/bRyUbMppuFv4qtx0nQnvv
3c3t4Vc/T9NkEymOX6foYheAD+UNFdalpUAt2Kc3fI9CboYACk3WDVj9tZNzSU1EJe6A9Tv+i8/M
2pokjqWXmHQCurpXUE9M67q8DigC4zKpm1dBxx3tJAaQVQiprzU+oGrEevRgJrF02TtI/ni5wo/x
XN7825STeaO/8Wjd3ibMOnML0DrxL9BjCHf/BoGllq1Lb1unLvfE8ucDqZ7xzn7Mwh3IEgVs3hIP
7Pq9Wvn0Jc9pgZL2bX8qInPbVrGGCKKG1i7uD+D5GhXTZCganluteZBin+jzjort+yAP69XqDPl/
Ox3WN+4W2Zk7Tw6YF4yaXofQVsEvlwP7f48S4aRxYDRoz5ELKwJa52INHJ/MBqxv2czZc7X/EaCO
yt1nDnH8wD1oQ4vqCeoXpfH23vAzsWvjFrL8t1oZxYIcvhsIknVITnBUZcjiWigrkEy2/j7EWO6t
TdEjM3iRI5uiLqCTukbyT8ZZtVcR+D0GKbVfG+VwAhV3tGsQk6H84dJGr+DOT+i0BSvWDodPT6NQ
rnRm+ADbtQs2BYKtfP9hCCLNP6UqDWhtCouSF9RJE8LYQAA2TW33PmM/G+ke7ZUPzNwKjBEW1ld6
8JBFt+uC8crr9GITBu2lh2BS8CW2qhREfA98yLyLjCMB6usM4OzUqMkLQZyLMCbt6w2miHI7cEpi
jNjvn5QgFqR5w61glCm9WgF9NumAcZOPN2TFOwIebBO77EWItVhCMg5saCfUWO86HC7VzhiSgmqo
x3tRudSAXqFG3G+eX/CwCgP43Pg2XdQju/mL3g+VPQiRuyXftAj+2JytakADwDt+VzTJrPbBfpHB
CN3rm6YkmPiqLcP5Vdt8DYjyTWB1hsydEvplTZMnv7XSgyCN6lJ/RzFH08QrJLUSrEo+4a+2uISu
8Y19LT3q6GTXKZepHnWDWBVbIOXxvbhzqgd2V/ppVmiJXjvbfvk/hbaL9Ma3mUfC3XbLhrsbE+rT
45YExv9JhWZkWSXdMmfClv4m2SaGrraPLOvzr6IRy+YZ9GqSvA4z7HMp6aYpjzmE7WPNNyRq1j5n
aXN/NPih7fcce/he/XqXKXu2eJ5TK5mokHqgpe+ORKY1Ds1BSh6YMKGGRI6nNfxhhp4qCD4jrCUR
UBGMaAFAEHBB2VTRwBM3Lw9u8owJgL5KUvn4r/Wr2sUqcZMz8ApGfWHYKrNbJhO7/pXdb7RzAtOG
nuP264MCih6me4HBfU/du0pR1e8j94ZWG9UYVr+Vcq9C/2MGS9Z/kMdG3hc2TlRXANRLpbBbf9mj
38HL+FNQ/cHms7GzWMlOxIWmSXkEKeXm8HDfEvtxnzlWQ6XFpHjx1FKvj6bJOTAnx+0lk3SJ177W
dxsD0woBctHS1cySTaP6JxW06iTgpcdmjv4kmSlevHgSz94yGHi/8cES+KFSok23359AMctRkxfr
AAeW0FEFtgLuXCT3/amWf+wxq8MhBCuA0x5FfOLJx6DAODjELJ0mNwlEkfbxxEUCNOHhntNBAldB
d6hCEKHIhf5nqpHaO75vsbsUq+oYCS8Vo0Wy+vy74oT4mA0rbc06IatqTVZIqtY5hCvluIypsR6t
EJPoiZWNImvDzn0hXamC6J+9W9+8zP6xDVO0h4V7uWddjmPi/ySWQTXHKhhUC3iA1YFJYZPxHESO
a0SDiyCzY4M5J+p2Znm4uzqavDDz1joTE1A0vilnbp9Q57llw7Stud5JbhWGzWh2zM/YY8/RZ9Od
hTp47P0LZx+2W1HXXwJQkAPD/SPEdNgw0/MWPIX9e7NiY/RQLKa/H+bceQZ5VKdL48Aypz4vR7eW
nwcyTTZehFDfhMxeADAQFFUFYVUHlrtID0fxptEtWCAxcBw0buxRo+rvVQ4SGIy5p39saPHNxhaq
j431ZcYy+ROPVPXfYVF07GX/y0UeRZ7+Mxe9HHeRrWtRyOATycPEmBVdt90JJwV4Jfj0lmltc6NO
J1XmWdsuPPDXSEvvMuvHpSbCNYo3QANFJRrxj3Y5nzw7uA78s/f5Pw0XHdW7mlHmp6dKdEBUARi8
Xwx/WNeHX7FGEAQlZlHNnkquNvSor3HO/8slB1u2vIAYCwh/4P56VYbkgy7M8vM0UbVNL/1gIsd6
+swQgqCPCg1E1hxEFA5ZSK4KLXRQnw6S0rAcyl87qs8sErXaVckkfqIib0rJRSlX8J7OxLTYpSHl
UbtOYq7MExgTsY76penzvyYJKiyZci/w0nGwasrtJjFqRTzXqaZq2sQ4dOXFE9Bc6OKSUgfpICm5
FK/KNOlTiZ+iYrRmu9e14WuwBcttrLlWGm5z3Hk+2qHN5oXdWspoEY1x2MMIW5DMAG8BZ7v50+Tu
ymIvKpxGbMm2HbzaCQKgwM+9VT/auAZou7xLGZRpFbMUNUZ0YjBh+6s2JEF9nZOaEPxw363C4VYF
7VIoC2l2SA01G7NRPhEbIgquO312jxKLVZTrWixx0EqAP3vMMherY7wK+KREXYcY0vS6wVnBlNaY
4t0yZLQq2t5DHi4NW+A2j+zKre3Q8HSq9HqcWirEYHYvnyEKduGoWSCUm2ogpBJ0AQNiYmthFHBu
bG50DfytPBqgNmZhRovyrnR2+4FFgvt5LSTjE/vXnJ5MGASZgHZsRGr/+j9tsg0NyFqjJaRqFToR
oqsszI43tuo8YmGEU5sBFvWE8IHsh+mJVKgPLQjzdHm8m0YeVSb46Y0EmRFdKYaCKRSwLiS93be4
QHAKPjzbNNI0URROJx6BcsRWMXFz3EsmIJWtjReWmF5HQmXuw16tWCROi/zhBxfVUtDSnM6d22Ot
13vvSKsZkANujaxtRKp0FSX03xDfmGynzqJTqQvVex4cpQQ6Dr0NCUtKkARbVwzF2O8b9YQ2F7Ap
Il4d8b72dNCy7Uku5KlSs6EzOVqxVnNZ5RY34BKvfFCRr//t0ZrkOqVtphuCHdt4oqSXMd8Fdv6j
Z6DiqKkFPSWPo/zz6uu1L3CxbXFpgRHw6IxxlE9mixvQGFpt5n3r1lz9Lwxe2G0oDjlAVEN9/9bx
b5TZhA4EJES9ADoPfa9zyMfcAQzW5pfI2Ns/UogzfbfYme7WLyVI87PGwpUXLVlg6XgxGyAZ1H7r
WWJymS2upGJjhNQCLi8HHPdMI68MTMg/ad/2Lgsu/VS/qJa37FWdYUjCIRfSnP0xNaUsqT9DYuJK
ez6tAvF4NqQTTrmqUKN4ATKEtFx2VVTMFXUyaxlB5uxdKpOzbzmlXc4Ix3ynVZ1yupx7fuHiZso9
nfTAw+QHUHMu/NkjLJ26OHTpyI9LdPFKW/qW9BvmlkckYL60hWi7WgdhLZEaWFtRjIQkna+kim+W
xRDrSJ4JFf5Wa4hnmWlCuoR3N++YveFBzLXWa0zMEOH9/6Jl2rQUHNGSfUR7fi4exlHew+6kgMuo
9knAkWlku+meArpyY1xCClhQA6mHHRlQms9vsJluDkE32BYmEBAq+QG4zR83GQ9ohd9p2fR70HwJ
1zkq8Ux07Qnl0uLZ+Wum27uAFTSZQ1WaRA/6diQgVw24guYIT4SNKSPboGYBbBr6N6unyL8rKKkF
w1IJjem3SxDDkdmKU6uX4JJmEfN7tQyxtOhKpziM9zVeCll6Y8XGCh20my0pfypIXCy1yFU64NQD
ngAe4meeuQkXGIuVgDlqcWSCD6Tak/aFEUCymZsF6q6BNp7BB5ppVVB/4vGPn3fPGehNZEDEMwtd
xSPlTuLr3Rq/v3JgoRm/+FxhVEekyQloIG9qKhdcSNcwD2DBp45WrAQojbeZxzQvBOPj2DvqyTDG
iaIs7rAAL5g1U/uuIDHcPqRqckq7/MYrTJoQbW1hFyInhwbE9ZrezJnGi+tn0INyOTQeYzXPKG0R
/YB5g+ZvaUx6gGveaciPdbx5OlUG8J9x6pkrSbieieZcFtoOYjobeQtqnCo+YqPGm1g3uPvYVENj
/l6YamVRzQ5ue7H36h1Ugkqwk4xBOip9OQf1dRIsc3U9jlgN5WYF0Mjx/fJEjMSclVBdolSngcO2
b5DqC2AoiI3VDUht1JV8fAXbXqY3t7dNSOXNcZNkWVY3hTbx7iVzF40V9mLfyGygXqV8DGCHQmwy
52didLU/kALaItIX5pRXf7OociKAHh9Njtxm/2enqAbBuyWlEQOwO7Lh8sX/LQEQk8qIHam2PI+v
2uIgF84v73I5m+kXjBQ7NEqkymlMKqEE02KQU6WwB8cnVkzEC/RdTsLVUuHXp1FI6dQLhSufWVEb
c1oF5nQuTC0fX95ujMJXtcettfA99PvxQjsE2+A3OyE0EMPxoUbJEcHgLZPdGJ37vMEmWYjmDsUt
iBodZHGpmSYUmsfhy/df0CA/M69Rl2pvLpDNUzv800x7J/5vR8YTmSa6BLQzGFyeCAUlXxyRwNi5
7Sa+TE7SpAfghRMvECMRxX4ounTJWAfbUvnFl4VPvNuzRWqTwAgRJuW+D9nJBW/9whIXAhPt3oce
41uqVjCvtWWCmgfRAzAvZcpxYtx2DqGNRyQE83DtRospA7nS+iKOEJjqVFt8UG4UuCCtTABmh5tB
cVYKnPIvRe6/j+5KPPZpHfLtbU9Lfgsgp9PB8Dq11QeobtAinMjixSCvU+20O+Nf9Vmjv3iHMN+o
oe0rANDxAnID6oHCRX+3/Pij61fMmLmU+GmqldQhUzYbWdYpZOzYfNtGCsmj9mzKVlzFMO18xThQ
Ms2Upvx88Twm+xuFbihF8S2ZDMwREZXIgMpk5knIJ3AGvft+3lolftmhyk6JniPbS6TozS9l96B7
ePtyCbeIr5re2XBjGNCn1WF9aELtNMjvA031ZoAmfpui5aCAiLAHwY+H2sr9XU1miaGCQ/C8076I
7as/X8+5JdchXxWgR5BLj8IDLLw177fpEQK6yJpXUJ0AlShC3yMFw+QEv3KoJ/P/DYysOf/Y3vav
8XGgyIQZmKkS25P4gUfECJEdDq6ESizhUdKXMmUZZG3dmppVoefR3qcj0nvPqYma9OW46CsJxM+h
1bg3AKUa7CyBbrctBOCw9sQbYxqpT8sTOe1NMiE1/KcTn6NHXr7jujyFI8Gihm/5PShpQ7eEjkZP
FeOCtGrF0a6mVUMFYnqtbFMnksA2lhz9/P5TD3ckB6/bWzPG8aSmtGlG487yTjquIkW2xjNmDzxN
mFcJhk55dQPfMKdm+w2eD8Fu6c7WFtXTwxGBgjByt/j7PixwWm9ZLVqMSBogVAY2z3jFQKV516gE
clH3j92AqBgy91C0YrXAgAXAf6EkuUVjUfVgKbdFhENZ22V72MDRh2IKr2Me6P3sPLYk1lImP03Z
WmZ645K2nndfjfepI6QYfK0ZVrcaog3T/fhtXT1jc8SXuR3ZPtA7Jtu/nL+rFRltAtdMXQ6rvPpn
cilGGMsrZ96JhwRhqLmXcUFx3XmtluR/nPm23n5eMA5EL5Cx/h5555ZyjYhDDsFMq3aXXnLQYNXx
j/+hr2dX4GJ0SCZALIjuXPSEmuI+hY1Prh/EdeGfxcPokstWbGbRMSBBxwNTQ3vXRPTaHG4OWxOO
ZH0RGvD5hb8ooRAWzPVz5L05ocasqG/+9UjgX1SSx8IHS0hpl3yQ+7HW32M0ITX0u4W+90BIXLWW
OAncTI6/K1ZgCAY7V3G4fJlQQA1GSlDWTG1VenNNogpRN+Ye8If8vA/0Zk8atsyQnPDfaBDhjsp9
D472DO6DEpvgWtMIMXWNQ8QwtzoR5bcqi3UZvUzbq35e0mcreMPpsfKY+TMjzVm2S7fIsrWc8Ns5
UPCzYYXj0qDfCjXl9j/6ppSy4st3QhbhAegpziZjB6Lyl3q6EUGNiAgLqld9NOGBCMDLD0tnbcBK
mharB4sPFzulwi33nEXEgklqpUtz/HXKy/1Lu8QalJZbHb05LfEUjXzjbfaMEIYjqoGpe3zo0KtM
yyeAjMxxzmsRsBoel8jP2bY8jRO+jeDpQZNLsY8WTZIwORL3YyvvWxkQl2sRnyuH04mFwJyar8M7
2dJ3C710RjdDaJ95/Wa1F+jhSoi/fr9YV+xm45fFFI9wquY1TZI7iDEzjJhMN1+xCkKXBT167m6s
/aVk3JK70dzLUYaYgq/0bbbd7SNVG+x7ExIVRtQyn5p41AhH4iiPvsvEhujmb+eETdAUsr9miPmm
/nghQa12NGlig5MVpFZm8gpHC4ENySC8uCFYwjnXcD67lrXpA7Kei4QGqumZ7gWxaDc4QTabBV2x
0bHQlM/To06kB2qAXo2ADGbUitXh0488xyMV2EhY3f83NSouKMvLZjVWcEjp2g9yO2JmkFaRqgFk
bnsb53tvvVzLWDvwByJ8J2kK6NOO5tL1lZsUgbpFO1tnmOylz1asIyApaRFW6joqkY1fSM+i6H/m
WnexAuWlFfeHvb+IT5m6rJGbanrNHAo2txQZZTwrD1uJkbV4FmR9Fio3Lo+478P3hR6I8gAindgB
mEy2zCxPZXArW3lpLsx2akSfcsrmA6/CkIBJqueNCRV4CwmMqORcUxF6IAsyBVBayn3TGdHCctC2
Ism2N5Rb4Hl6JYVZGPwXJoaiokNngly4b64ewa6YRjJaLfIkXaRrfK2odGQAX10NARLZqw3VxkDl
8al5N8RSuB7Y4cTRm/GPv+FIxB4myo7uHKmrr7f0tCfMGLX7RFBybe3bR5WNYUE7dqSbKAvaNfmX
2XizCkLsTELcprvvctCP1ddI3+MWk394G7cYIovYVOBx3bLcjzbQejYdVZPptUIIkzf5+NowSc/N
43OeY6zDVUD2uYjjxIf24TmPYm02KMV8gvqZxSLq5RVu0RBtjtKuXJJ0Q+uZ6F/ZyPz5BFhEOyM9
R634wUcrtpfWuUFELVGi/jKHszlp+8bSpiuId8xaO724AgHXZclEiIuBrwRQbdVFZl6O7+oOZRTS
WGgXCotuki6gp0BSYwgNlmpdPAkcZtz3PIDes4qCXQ9/vgdF34DAcVdWATe2epKuA4/IJOhMkNNj
MPrU+f9jzqwvEpdWMFvY40kgdbuAf9dheR2F/y+hWCYsuI/8yMW+JOKPFHyP2fDFyabfnG6FwHoX
PS6Rie6RxSPT/BbvV+gurygUHUAWT5zkuUe+vpLCrraWmBs73zqffFY2WlKYNAiODdoxQIOUlFFs
PY12zdaYJ5od5i4EBwJAEPl1S1+OwL41ZTSuw0RS7sqOisQ0AmD1rK3puKbxvp7vqUiBE8ZVwmgT
audGReNvng4064rR/Drq3B+h70AO/N7R/J/aGrQMrC86LMq/vsgTO/LKVhDZvg1DFcG5px+XhUV6
4TxbZH59ej6fEkIXEsDtUuX4GD4faA2VwRvrokPQyTvdZgUcwGrnfSmpQmC0A9OgFPZ9eqhFtTUl
pSddsYf6llggg0NuVCL5rlpL6yRN9dO+pTx3RuF2EvYIsdkPgcb0l0YXsHcRbD0j5+0wczkbKVOX
I4H7vCSI/kgOsHYzuB2Yc/pA8fpQCgGGBtxW9iWaJhvYi083qVxMqVVtTbiB0Gd+UH3f47UgkDR9
i9KaVn6IaPsbFSPJYtiD4KNdOFRIgpS+Yx3xcZk3raeZfo/yRBzxD1lJcqX38oRb8R2wvwLqDSgD
GkeNLujuperKNoSu0eT7d7H9GZKLmIU1dqqHNFSpsTA4vlNxZ2RzNLgohPTkYrP4OBhZna00S8R8
G69WVw7TgXUanXBr1vqgPAWsJlpT07VaaLuJrWZWyO+RLXudMtzUJzZqchrdktAlaE8sMmPrfEvY
H8DXS4fGJWSVRPxDBeVYbrNnMGovjXx3QUCOtnLbFMh5CL9wiNiLPz9sd9C7lCOz5TX/goS8bkzk
0O2tLn9fshuuHkIg1GG5+Vt/RqRBRZZwQHytcjL1f3e0L31BdhsdGNxnRaLbjDI/BBVxIeSqQ8BS
Usv37ljjBGICQPOwUBnE65f+MvlU1lBApj10sbtSO6sq3DDeRGTrYcd8MbhryMmIRxE6fDhiJCb7
B8L+APqdZE9PypFy0Pd1u3U6rzBnp+8VIEQj8Ctay8lrDRZ6dlBjej0hFkHmyXmQGCTmqk0HxMWk
wuXwxovRkgjd0xjNGxtjXpWjLjzrZgIGnnOLoaFNkY+7p5wtGy2H/x6UtBgDKf/h/d57S+ELjbb2
qTt+FbL/FdfYa7DGb65b9qZq/To+zyWUfzsyhPgOCZX5Clct8dqoe4YF6ljLpA7JDuJIOcrLWQby
Cr2qhWUIXy9SilpxdpHlN5CZH8IRm6MsVG7+T+4yr6BgfHAXKSNn/vz3S4HBE3qNtM5+18K5OE2C
ac9FP4siNrsuOjeLv+LHK8kAd5JJJiqiPEEezPSL5YVe/j+hkn8dqt0eqFAHURwECCF3fwnym7UT
4860u64ty29qkWmElDBi/lgM7kR+ULFa1D6+ihO/3nm+Uyj7sQ0BZm3V/ubiPfZgQwVJ3vyKtXRN
xMxb7flQeonRIlT9Go70xgIHFWQKamE91d6aS48yxmhqx6ztBqLWay/adOOD8+z+yh67bUH+UBYF
3HLfTCFYj6GFZ3Qda6JdSQ8+ieGp7NOtrzoCH4JBeAodxoB9yXNP5gv4ie3nftNwAt7oGlZxx/5p
8fyj8ge9VxKrksKBPpgHEhe/qLWNfuJ3hPgckGMuZZeQMEXRvoqOUi+ElhRGiZsQxOOrqXA79b8h
JJPQiINN5PhjIzj6ztirSDW61Htk3F4oXZqhzfSdWojOzXxbfKSTPYK4vUf+ZhJSZ0CKTnBSfBix
vFGnWCcHP4FLyKlq28cuormPBe754Ab+c2s+ntVVfxTKPdoON8/NP2vrgeiKGKkh+PGMTvktbL19
tsohBNX9KMtc+jYTua73IYn074hNs1il+OFKGefEdmSxTIrYFpYApcHx7VnLXgTtZdl6iSi1xEe/
qBiebXpEmg0aK/lELwnorChh8TRFqBcr8umWt61ZBbYIV0dRJGutCXrPp9gmAL1Dkw3/BeRezfZu
GrC36Pe674hVDBqFhZS1sn1FD/5MBjyo4jfV1MEkBHZeIuJwL3zRJwgOqN+deOz7+IIy9uSKhgT7
ev2JzCCrhVyXcThaHOZMypwtyeVRzkBKnORXH0TmMroGVVvef5EWY1PHgu1zkvZIsadTgrVxXfbT
Wo3q/HcAIZKxMYOoJucvibLEcpl70OpOz3C+uptKWvDqr9AqtzcLs6dqf6Oll7DeRxfC9wHVDVx9
gxPsPyYlVgtEiAKJFH2x5hxJBNkPpPZM/vSkSD1iLVSfKSlalGfjoEPbvw1+cNLxx6AcI/6+Swkn
w8oZ7Yzccb8BfWBzj5o6cI4s2CQf9sW0s2IxMgKo1xzSjDCkmUiXTmgAHabTqXlOrNk4Gf40lB9b
LkfkjBlcr8CJXCFcCKJgq5dfpGkKmYTvsRcvcVu9Zx5pVbGR/e55QYVHZ5tc6W3zHauZ6KfBFRor
nplk+jmFCJE5Gf4zkejuVmA8hVAn8ODQ3a4nkoXLM/3vkM2fcogTxby+3Jwy1YWUFBeaPJNxDvAC
6zQyav0aik3LETh5uwBetttp4E2BacxuSACQCSXFYjAtFhCr1k381PLulZtCpj6WLoJ6IdDxQhlT
DQmi1Zf6whl/78gyABh7KlRQ36pSjJKwOjUwQknX5AXLocw1PnxWGzszc88iSHdpk9+8vsZbwczI
o87/s2meQtQZF6kwh7TFMihE6DmfQ8O/ebQ59uwkflWdj+GC3KnCkkhdJxaBE15utKSQnhI4yIl3
mYYX7OmeJBBUhrEd6Z/DJxfM2mIKSiXAol7r6tu1KY+EImI1Sz9UKt1aZg4lGPnawUxP4ciINw+K
Amr8ZwIqj9Xd0rhI6O7Oo2GyI6bB/863e3uvW26GTHaunYbm/Lc5txKIyJKeI3W6v30k8J7marFS
Wu0kkOD7Q3wgRIlIjg/dFdAQQ/3TgPBGEaZ5Ix14eqpTN3/XgCixpfHTDDv8JwLOJeuQmZqQmL9O
r9z/KMoGGSNuv/39V/ZlHp3uS5zbPcpn7MOsmEQ3eyeRVM/Z1K80klIh5zo3HhgqWNypBX+mtvT8
q6xxFEhT2cXeYmJpYkl2fCvTZR+FU1YeAjMgkN9QnNG0Z3NEcAEDQCscdCOl5YBDN0EQu4lKSVm3
oUtQ/1dn+aOWwqjG1O/uN89EbsbT2UF3Uut0KAEROB9zCJMv8NZkU/mcniVMJgQw2Y9++j64GIP0
MiwoimMdpmEepbR2vvvZeRZjPOzuZ/wuqr0xRl0+lwyq3QKsy90GrCWmjoz/xBNnw1Imt9FdQAQN
W1GbEMltLTyn6xtMVgpa4zK/8gQUtlzi2xJW6bh9kLCOpRBBBAZ+ThECeZ/uvGRlqmtVs0HB2Yhj
U4ce2tRw7X9GKI63C1Vzonz61N7Q2dX6JAdZJlIhhj75eJPdJMOTi42BLg3SY1Bj7q759dYnTjDZ
LfCWS8Gu6/zdBIH8K9DSeDcq6dE9q9o2GM3nsJ4oe1JR2gbNw10xYWt/qi3Z1KSzOBO1OOaFy8bg
e6WqYc4/tmbM6Jc2NIIhDlePV8Ij5RX9ri+cpgi1+7IZwcxJGnbb0FOjWzqt4TSs0r2eJG3FRcTw
D8yfCYvx9bNfycgV5xqcgCMWX+rzpdvsiOWLOOr9BMpkCz/ZchpRnBbYqYbR6/BfBfngbVilTxmM
68593spocM+Fa93DwyB0A7I6RufyOu3bEQPil24AkgABHlMghzNiapwhfqSHy22I3OQiaeCBXewb
DcFM0JqbahHBtqz2aZZ04maONYKc1KESPJf+DgXuQCnp30dYxhqxV5BcCfR5H1Si+CKRQ5PUa4Of
OnuQXK9/P/RupK3SbJMzjzokES2NNAfLsvrTCP6mtaZh2qI8X9XLJV8PFnuZDp31dhqBrT184O5C
VNfJ+Sh91fnDnbRJr7HfsI0cbOCafHIp8GGNDbXsVE78JqFdHd73j7YUEkCmTydviSW/ZZLvdEf7
tWZjfw3CfTgfLlSmisd05u0ovIDG7U4ZLtpUNjE9lfc4aB1T20oOqEdQT2o56zhcdV/ob440q95i
LyoWOC2R5lv0OGBT1kglCspmzdTC/7Gp3zw97OTL4wnQHLc02HNm6mHJITDGz5MF2t3KLz4jIfWI
D9k56pn4wyPlV4GAjMAI3VRTBaIXBqB0jEQPGX6zhPuL5B0EV33U8GGw9csjtneZJyrNAKRuAEbw
bIa5Kl73Li356aUuDLFopK2d3XZFaPsk6skin3n8zzrSIR+jOdaA9M4QZf2kNjEpUw9APfAF8FiO
8z9C26bZCEprPG3J0a1dT+rPzU2iFe4q9uaDhq+HCknmTRc2dEVkUK1GZVNePDvcW5x6yILqlIzM
iJTC5eCUvIKvoZZWcu4mt/k7QrZZ50UmI+ETY2MmvX+bYAWDmAuptXOYFDh+ynU2OhMAhhL7XHB7
SQcZ87sbWD8U1cuivWsvuCaw16mDx6NhC/aBgr3+xPmSeQoyhIiKrR+NVqdQ8XnuQ+RHPD7jwTti
dr7jTLqGTuoxd8KsDbEHUHQ1vScdjGjeFstdChNovhdp5aD24dLpFpr0Dv+N7X0GVQaw7A+jUmbT
Y08v/MJI+vgEDLvAMFSlZWPoYPj2uX64W0Mq/8EJSgIcn5QD4E5PMD8B7v1w4nteqx2Vk72/urDb
EQMWuw1AmVpB+vPPXH5fl6cEiMaAxVn2k4Eox28tRo3fOGL52MQKcPPdkn5HUjEP/eNJmWB7BYMZ
3JBuKx7nQ+Ai+OqGOrMUkg39PTCeLif4As6F6faRcVYdePxzis1Ich7ZV1BsspzRXMq2VvnNmNfJ
SFKfnXgnET93yPYCL0VQhkJvRHKP2uO8NUlf9FKck+6JiRy0p0MnpRcTdKZ5DKejZrDoM1X8kLpy
mtks9LFTitATTnf7Ixr8UPbyqlgvgNtNYV9gkca/W2IE/CuOWqyVc36dofI9qJM0DLoYbn31KEBr
fw8At0wpM1DKzgH3wjay3/wgjC217hXakcvxQkpdiQeQj16zTiFTeo9k033RRWhyVxiJlM1jHyv8
xI5dx+1+O3gRyN3JXDAhbhdP/ZSNZhzJFxi2WMwV9KwkOCMuytpa62zcSs7vkiPggATludC40vjQ
zeq1PFEwiWkv0FMIKMAAwkE2aSsI2TH2ekVX7ziB1u1jyKXSie6H9eNiALzGOsUIY5XldVTx7PVt
6t2+UpCan9KbcC6DXRWLCKBGCz0Gl/Q91kJndiUDdIbOB6q7K41A2mekNSrvSQjIm3sMY9XVmCUM
2+mB4abHhsOP+RWkHDSQ/VEDUeZMLD86byx2ZaDNzisqAv/H/TDgvTig9txXF7BCisrO21bwXDBF
CC1S9ZEaDNjT6GjLIo+fbdjZ36lW+TN4KLxtJ/v7lVyrvvIVHJ0E1zSmAi10aka7vQYQuzjIjfFV
lfY0usL8Lc63sfKFHuiMyafJgVXG9ffOqk0e7KfQrjmZxezEadU2ptqkLVgwtzIAhuh4vU8lg/V0
/PwGOxjXy+EvAoB4RxWzqsywFAPJOsLZKqvjt7jtqEmkTLgrBDl2Mwm+riVkdra2AwXaAg5qRd5b
fflu1vMskFJw7S7AhNmt4ewVZNGfyaV6NoSWCZBJETzo/VfrOkgsTbvfHw1Cb9BR8PTI3Gqm2f23
rRLtATvHucx7uf8djC7Bzu87/25qNGdF5cRnAYA0wOwnmkpBu6rY0+rB5rHCWmb08muUy/uxm9qr
3LMljHG2+97bsB3QFYjHj2N1TraFxm6lXg6KBsY8u9Sly+anuXXRmTse1vL9frtXNiXUs1z4WtcV
mmf966Gl8Uh6D1zMtQHPjTKKprLEqjp6PzSpVpQ5T6uEGNWM3R92tzabM64PYtbrLnrxJ/5e2EXJ
+5zp1VVKeJBirPa916p3yJuBAtOpuC9EaFPtR4f/799P3sh6jxMQ5GwpEV02wXqq66ufpAtBqjg9
ceTJO+w+bliAvLu6eHNBnN3Ng5gA6JTnQvI8t7yDHAA4BFXLsfVW4OGx/ccZtfTr2PcOH0/BmOK3
LMRErlbn8GAnKDtGJ+azeeocVKfnDpA3LZ8AB1js8vLi83EMFYCDb+ajOfCqB0BZL2K0aPtSRzco
ezQScpbwHlPMYtn1FgOwnAC2G7xERO9rYY5MJO+IG2WdpjuEkkzO8lNA0xU7FYtdctAT7IHnbirJ
X2NKqlOzcwih2aEAgw6ObClXw9e1ATH2tzVr9OnG8+KsVutOW1JFFogDptkErtakufCP4uNUika5
K1jxMiQpWHezgXK53gXALUQrb4V3yOgzaJLKrQHg+UcF45qn8Bkruk4f1z5Q8a6P1QbuVQsQSkQY
eGY/Tk5aoGCJGGz7Ao7n1h2QPIlPaby8OtNaWhfmzQD5nr/AQ11B+nLfYqJ2tDXMHtgjanqf38o/
WCT4NjH7vUzBAg7xkxf/9q5a4Zleg7jSoZUEiwSdK933CsQzDsJMvYwyMwdE5gEnoqJhsVeXJ2wM
uIVNKmu7Dbgaz+5aPpQBotbXEwrPBmD69OvWj5NGNvPaO0lSv0KUCppxLx8Ixdevr0YfbC6sIXXW
cwkMMneMwZfqcuniCpS1aYLaiStIOjns5ZmbgS3+PY1FcBDN+EYn7v0WHECC1s4ZSyEb4qybsAcC
yBSpYPQxAS6+D4eyl75KyE72jpz43YkD8B/hM1MxYlXCZVKiPBIU6aY2PwUzh06pu24R/VhbiPMF
vCbuyIfrxXqHxxJtwvQmgfOZB7sP/dbUr+P/55VMXOnwk1A3BxMcPNU6r3PFR3v4o80o3W7Bzm1n
wJmNSpRGgcxoTq+s82RjoXoNk03QrQddw5+aubjDw5ssKbnRT8VAdHjIFzvdIM2AonrqBM/UVxDr
ltKw+7Gbb8vqUKZfKHW6fbR7pq/6F3/DVii1vnElhyTtxcImuwubwiOcLKwXja/5N8R0DVbOf22a
8OSMckSRDFBiAHa9ivSOz41KfGPPQ9gCh9gRNnFSbEkLrQy47mX5tjzCTO//I11J7EoziWf8Z790
yceqp8JFByLPB4069DA72u8M0bbbPgUQosfgrZn8Ac8k51Lk6S8EizaslfzPsbpKzQGUVljzi7B8
a3cF7ccFgZ3IkZO3J87p1FVn17nGwUXNYjFYPQXrDcKP7fdM3dZJNBsth0wCytuER43tjjkz4SD+
DSQ+gjkyKK3oKi81jRjNhI8aFCFLE+fqoR48ViBepTN46rnS6m4IBywP5C3dr0l85Tpo/hwAuSOQ
v07fNT/MC07+jiX8mNqwQk8bHj6Paz8UosqvX6roMtA33Or/zEmC5HTvOc5thliLYPT3TbVL1MFj
6kN8iyRW+2934qHOn8ghPc5KOrdVN1nkXk1SMb5iEbrDGTxSe9uhcBKwx9ikgvQIZpQBzmNWCaYM
69NRv6fVxqcxJwClsIL1NXabDO4KhBp9WaM6kJ6BnkE8r7Vp4xaGBbub1p+XU3V+ZuTZnPdouJxT
l7+bjryZIXVw1uIG28XNidc0OGGr4D5ANdL9UPS2AjpJRrhevFoUfn4o3nMHAwcVi+Q+HySiHxUN
K7mjoc/d9867sqCrYncCJydCnuy5UYdtX9dRGH5kGViAxP/6s0AIFKBmU1wNNEMEJIULZOuGIgt1
QmK22VF826hd1WSgFvcn5uPtr+gWPuYTRoiSxebZjECqZEIydU7PT7H+viCGaganZ/lVGX1I7IK1
ljGZvWkqdhTrNhPDw4lWo+lKp8EbD+uKoEsFLBfJ1fcbBgUGrryk4wDavs+PE0BQWm1+RufmwZZA
3rIC4osqGZYLw85MA7uKa3GapeSs2OUAFUEu9esBrzVM11eK1zg66u0oVKs+6aanR4cJDPDF18HK
4/Q/mI97SJWfNrT2qveHZwxwG1xQ+5+CWOJI9gmgaQ8rsU1zGhV29hZON2mLhmW8TORQCBBNtjWG
NpSJ5+BEujarGCHG4wAAF2HHXM4ximpvc/v0Ne9l5PqCgw7IKAzElvSQxH9KlTgN8Jip+Aggkq+P
hTM2yTdrDr0adWWPL638mgcYC8kIFhKLE/MGPduR1eq+nI2pv3oyk2PTNtJJLKTY38vsnGoHQGAc
8heDiM+8Q2JvqTtLCAvx/4ElMBHY4VUUO2QWsn+yEA5HePd5tav/vNd4s++3iIAswviwNV1mI0VQ
8elhMyLHQrDGZVMLH5IXCn2j/7JYY5i0vO+v72ZzAN3WZJOQWpbhiBsyksuJ44qREhw9XnfUnipP
JlbHu+XI8c7PPcjIA5mJltBo6rdqaJWyqbtz2ZnD3N7pEAsbkHZmOZC86NSbHSAe5yjkbLw+HSk2
PF67Dz8WufmWB0eYz9Ng3BFsL2mJHdp9yj/pq+5hNj/50Ht8o8OowW8yqUVIYp2G1m8kkuZnXN4t
ofWfAP27fvU0sy3jO2ftk1IjXk4T4j0SdccEYpZM/B893+Aa/qaGPlaSPkLc+ouVAWEhKjTOqItu
o3Eghrucbx8J4MPTRdzEjbsLPYltO5U9hZ7hIeZcnzg03Ni1WxF3BPvEJb+nTMGh6mfRjtlgpOdr
xuxyRKk61i2b5AgLpnUe1NPqxt8xbF82+Yk/SSsH5HdCCA1UQpTit1W/y9H1U/Or4DxC2Wy2FP9G
D8zfHCfnHQA33sG5UalkYWw8If00heZYRrqR/9ICHvc9d+YbshVFQReAA9tQ7WOKmS6+TH7RcG/V
UYPn2uvKTX2Ml4DihzveuMalNai7mXLuYWOOzGkjYARgF6tVEZ3YTSjFq/OtU1p2lSBK5yWWWtVp
aA8sBb5kXW9X5GTNf9eK7rZF2LQwgfZHiQ3/uFAJfxfDgtLG+FJkPXOTyEoCYqCtxGrPrVloS/zl
l1LooebsefxbesVsuLpAjAS7Auu3ba5bW4myVgKeZiZASiuTjNkdyGobOopEFMq11HaoI/8sahDT
8lH3uZfK9nnJFNYC7zFxYJxueULiJLd0CEvAvOClc0ta9jbWigdbZLle1LK3hMai/xORtIl1VuYw
GfyjtVLyyWCu6oEzuN/UX4t/MVLWES0rfvuTAadtyv8oIt/N5km5ahUBpcs3n3XiGgrs/OzNz9pX
bpxTj9TnFkJwfz8tOZPe+19Lj5uwFW9SkGEbWjZyaX/SL6rOUfhmMub7WS5bp+tsuqV3/pB+1Fxo
QvEiYV8psTawSOrRRgIbVQlE6tjGVcqZ+UugqWZfZeGEP0RV00UcFA3Iy6NKdeiPx0P/HwJnZN1i
smgAWxgcxhBjSgpClp94ju2id4K8xF8vG6geRyCJjuQ/23Gxw6y4xx3IcovsprbjuY2w4DTiVLee
08PiAF8LlXgdxqJ8dVlcL1NoR2XGP3aLgBDOAdDp4IEcE+htJr5K6c7CDCwgJhIwYy2m+NElVdSl
FqYKnpdFCTuOeDpm6NkVm++Lj30TY+/2qwBis4tRtqvy4fPCA8/MbQEolo4/QXlZT+krZAVKq3+Y
oUCve9opO4A88T+p/jV6UwjW4SWK5tzO1OEDD8r0bT6zAtsdGbt7GxKLdg5djzdISfn1m9tqpWL2
qiCgZKBI/Z9D/7oF0SwDz98NwzoLyeq1RS2glnB7uOqNaF2IiG9QCCggwzFghW1IbiFIFMYhCU5U
Ga0PzkgQZZEfH9VrCZgZwx54GSP48aplFlIbcGSKsWVR48JqwviZeBcClCu3aTtJY4T8lKbpZdO3
JjfDniTKxmfZ1ZrJl0hgkaqM5FPc9yEi80eToUl4BgcuD8r3dFtneH9d8c2Hclr6LzmMo9Plf/hT
OA/Fbmtnyb+xAneDUdEyH9DiKAhCIHtRmQZc6e7oYIAELE8FaMQmJJLupaDat1V4q+SsfvXZ6UIw
XVX1UbbwJYuLL6IaVPCxqYb7Ownt7CjvYk65/K5titIzpaAw5Kqonf6fn4pjhTuevGT1ww3/VP5O
A/MRlaWuQDpuXmyxwss7zt5BLxjf21Bxr8WCFTfdBVXoDMsWmSwh8IY9U0P8PeAxx9NmgWaaTqHj
dGfoeUYR5R0pl6DwD90xcooilFMGkdMdAbYTCmVQFoCz+Hyo/PbgKsij1UpEhhUZKfjHldYpb/l9
rPQ4pu1LdMwVSbyYk4Jdh6lwciKgrEMtIjCVDB7QIVfkGobA6M7ynQic6TA4eu5inXqKluijR+77
DNp9uUaoyXjtlnbSj28hm5ds9W6CDK+idGEgKvBAqe+/fU9FPbNsReeFeulfCv6iS7QS3F5fH6aM
GHEk/zTkktxXGSm14poQ3Gslggru8qb4OQz73Ydee5RdB6PmVpISvmQeRJmZGPaY3NeFzHuShmt8
C9OVvnrsVVlvCOALtVAZ0zXeCQnqkll2kkHR1nXotFVz+ohyH0hDrh13oQYFEZa9bu3En0UJNMdY
9IvTxkyQYlCpHywjZo5HGvQKNH8p5lhePXTYKRdwHjiMUJYpNgO1NCX5Q/GuNky55Nv6nmYo8ajI
P8cmY8h+qxXRw7v4VBbHOZoSanxRrb/8/DZrUZpz9/+9/zvkUeC4lvJdPoGaNcE9x2BsYWxxJriO
c9a6ST4p33LDQrlPqigyeoAfYTIjStmXtxwemXySjswfr92ysvG0SJ0YLrWcrI2IOM24GhU8r+CF
U3dp8A9HtKytztCbQm/35g9XeUGaQO98wjVaz6CEaqRQxxyNLipzAnj5Zkmoze7cYWoo6u2gnkF3
dAXtHYar/ktGaSeZJ0m7Uoc77r2KkMQAs4E8l0SKZv3UtKwR7YFMc9yy2hM7qVpFtmngL6Xj5uZg
MzHeH4gqoJcBLPbL/liQjhRLhMn6MvwdHrFKY4GLHwlmnTH6SKcXnQy/aeTl/TZGPhZcVTeUc3ia
COILRYncb6P9LDX/BPcY+2YxXNjXKcgMojfipJn2mCBHJf8i6mJK8RIP0dNoXlsx5RgNOg2mSct0
kn58rePQ0ySbyJ10nhiMQ9SK/QKfx++w2hawFUxArpq2MbZhvlOR4/VqrESpuRzAVEIQhIme88iu
FtTpkUh/UIDcgy7MUb52KI+Bl0dfwktB6U21PuEgUKhWqVwRICneszb+4wnlVTN3YXBN8veggDG3
FtvneDlH5zGY94h9T4EeOdXECNgEwS+rAa5YTW0YXpYx5/jYJAL1+M8POJyEEJzwi7IE4jHgnxRd
fWGCkhyylwi94ERvPM3ymFUqF0dmmT1tcJJuW7p4M4SfYA+q+ZIsTJf0GDnbt4rDv4EkWrOrcFec
PdELfMQ12MyDdQ2nwirl8ShcdfajHMvdGpKcJtQ6t1FksE8WcryKqDU8oG+IiiZStRxYqv2eRQoO
cVkib6xfy7u93HzgBp8FaI5LeEQR6kJOMx1qcLu+oUkvDa/TJf9jJ1Nc10XbN+1iGdsUhaNNIQJH
/WbxGUM2104IOqtJNNExEmQ9AOKdkDrLNqX9hPIMzHwDecMFrd9zGhSwAuudOL3GRC6JGh53ghX6
ceHB5gsDkTb6LFl/9RHhCaHPg+xskZ8kDhjh3hb2Pjnp7/mzuPFc2+pY0FPUzDAQCsiD0bszkOW1
uBs6mULqGULCyPdNzxIchJS/gyIPJW6OQ7dFaldNUrpsgzACqDBf1EUHSLcIegZRFcZmyWYTzHEr
5oSZ/+jKI9AwKOfN80An2Rnl+Su9hiMt0eAdJPJT8hxVaDG+MXx+cVYRG1fxCREqy7UgpFfFkJuL
Gf0ZPhatymhRpRkqzlrsXD7ZTMVAjJOuUg6UBv63ThWMa5C5VehTANcs7Zp6tbt0C186YvpL/hDK
rFR/AzSJYNOp9U/OVOGA4lchzDy5qjbg+r9COlJmdDsITHZSz97UvBdx0jCbJ+SiNw3ZsN2Rn0a4
eS4Xc5DUcxTw3Z1FNKYAR7HaljLxN2he/KD/RwYM58UdXQM/Te95et9/xo1VkFryLEMaQnONSfMe
Moa7R2qY3dDbV9hcXROU/mHinzUe0cS38+TaHO1gfu8dZrnfN4fNxgIxTOcAfN1/puyKmF20tuXr
mFfaxVYt8YA69OClGt/dxYrP06JcsFZidoWZmv7grl4XGPBoPHqx4XqWteporqwajlCzj0qoAmpK
lp2VMFsOZWBoc6NVKEiMONLtedyXCP0xpBYP5B6NNL2mjTJsVrlfPUkju822BIP5ilQiRnbWoTiu
br21Bd9XKhWdTK7EiVoAaptkErzMm31L3QbGUaMNC0RV7Z2CJTRO3fjqAgbtbxMS/lb5Ss0uFle/
tkpYXfil/1wtaoH5xwWY94fEbqWX1bvWKcAs+GpPEEUCm+5hb1Z2252AS2f2+6K7zf4KybQoekDc
/B2JC9gBH35/jXeu/GdXjP2Qc0RakNI9geZmh5wikS0ZAMO6OTVRjoOr9pC4NspQKDWttfJk4c4w
2VZO9iLloV4yuCyiqn+M38dEvHp+Xxb+Y+EiBFVHeta6M4z3oC+YGjkXVRFnR1tePkDMKLKb5ezX
8rXjHQs2wo6iJ+xl9D1rtcIgDAOC11UENPJ/FAyyZC62MbLvBAdj6iXtsVyBXZO2Xbej5hUTmY70
yQ+egU+kRdKYAF8W+yZpfZJLmcmbzOPoqX6M5midIYFVXhCZHL5K7ruBOcL1SGw/xfB63dRirT5p
qsMM0ts/oTrLtb4Tt8eeS7VDsn2SqHSTU+nfzVGNNfsgTZ0UO4RNWQG4poL0W8KiyY7Pv/F2X/Mv
EAEcemHO/OX1ZvRhUY/1PZ20NVSesK51P3SroDlr6FWobLcW3zEF+i/QpHwHWf3fchyFbL6YRD6I
7L2bLMfSYmuNEDUQq5QO7pETA9kW+5gIUl5/cjP+zqblP4m0YafIORrjq3c4Jar8KVSyCMXVWD2j
8LuW6t+G64R91QVQmFQrUa92GMBjXwes399O+W7VrPb26g66irICi5fwwrsK1x2vPtj4I1u9aYEP
1UrHx65qpOh0ltaM7kHEbx8FCgeEbyM6fCwL38fdymOGsGbEqpWpzgFCqGwzmwrB3CGYiwZ6XdEN
NWyP7oiHjyLjx0QINEOmWcp+jQ2tgEIRVUXxTI1NYs1LE8TRefWCAc/ciHSOqQx8Xxi/Qvel14fZ
iv/DyvjPUeM9xLugtaYEmiVhXXMzmO7BqDRvdJGed60w2rLbLM1q5G0NqtPNvlPccPi6+y11IfVw
a06vDteUJJ4bgF74Db9Pqe5wj1ws4RVcjEUnyvxws97bReYJRaCCpcz1IcJsGEZpC3DJNsfiRp3a
KyoEZ3nxLlZbTg8GFzcB+vyeQQyLycbn6w+D4IcI/8gbmOBcl4T7iDFqSmCr0Dj6qlttjTAriMpR
QvxuZ71Mky007tb8SspaPLcObHeqKEz2iSK4CR5U18rz0Ore0ZhoqAONDYqln1eVeyieeCeRcwUU
qFbl7FNtctyCP4zha5NrUJvT7oepyimCCHrjNeqVIubm+/uiWzerp7Sx1W6vtXVC2VtWa6KIGsTO
S/TzuBXqk08bvBMeaSon67TcEIqEdygxOjeVM8Ojz9Cjk/PVYoGkfAdMjVIoKT5nQ7s2wrRmqEQG
nxXdGMJetg+yuWcVkHzJ/D6sLtQZ+jVP0Gyw8VSKscB4VJyprrBlMvbt3BMmCG995zq4k5xQltjM
ZczZA2YACa4UeASSEw34h1c8REr2u3JGDePUBYqynVsNYmMyOGBMOTUYe7IgNuVEW9hjTH9YbGAY
4IIRp/Wjfdvob5uYqmpA/NUOYn8CByFish9b/fprFQw0g7aMdBWFgOG4mKttFilgoAu8i23ckYBz
9FOziSLd0alVcXalk8Tfm2yoci2iGnIv9sFsDb6ffA66XOZOuSj+xP80nKOCr5vWOF3+fM07eWgN
omSXiqaMWL8JeyKrzFhiCKJbOpX0Sss1XntzRuZyG9fkIMPqLAhFFbEzrjwFn+R7WzHzHEjRNh82
YNwliN+kpJI5u3tdQI8UBgv9uZAfIosaBfo6f5QCbyza6L/2nvi5wQ/TY588u2i2g9c5H6mx3TOm
o/b5G4XitDs+1EQ4+icIw14C9toWslnfTm2J/+IDdmbLhtiIDY5RhhQleVjWBePJfsRffceBZY2N
66LaU2u4Ruc7VpDUGdmHym+y/Ru1KHxnhJTlsjGdAuBh5gUEYn1WKHWTSPBrQMsb5PtDNuJXZJoR
3SsP8SOY+nmcALYEi/+ERAv5uPgzMAgRlLlTSrX3LGj6KdHwQ8LKsjOsziS0oMuXUCbs20uEcWcz
mdLOL22aV6Qr6XuLX/peZM4If6qjMgijWCV8J8Gav6X/QCyeDopoXy+F0HAchhIM5GOaVpfx8+LN
7VshqAde/U1f6EZxruffZSXyx3yW/OKxhPKq9sQ4PeJYQeHUz7p6+kLNtS9nu/2EVU24h5wNViS5
FUefNpHK6DXK66AMN7rX93Y12xGALJEqUbgvmCFb3m1KHlxHo5PJLc71opVOp2CNXH5uO27ZOjA0
WKe7ZBPpreiVNrt7OTwteuTy0DRQZxNVsAwIdAEV/hyIH6bzXGeW7BcOLXscEDi3Q6Tgw/TDQCnD
qm+ZN7VPxFxshZZpjq2csJbK4BuWCcBvoBL7D1Gq7ugXkN+WSiWAzNqeWQ+FN94o6EnDU8VqpQVA
P1jVu72i7jVMub3Nq/BXPyO04SimH2nH9Wj5L68blMejxHPL49Wk1N/nyQR2ffMcBf3rLLrJBlRj
0qVmrKPUuL/zVFgcWjsShco/fFKrlyrNHGpr7VxpU9sHQCiAY01w2Rfd6KrsOhHV90MVS1lD+w5F
WgbBp0VUel5TIA2DWLi8ug2LSJNmHWPPrxHIDe6dE/nRaoCVSCCbwIFtr71tbwDKcWoWrU9UC1X/
Qo+JIvANp842effy/AejiN6+t8oQclmS/86Cz6ZUNPRGHv1EizBTLRwmvMV6/Dv065/K1PnwYaaK
O4/OxydNP87c3KCaE1QstFI+Hky6r9N9BsvO2eBC4PICTGQCe6rwplbnNp5Y65lfqXRkNLUTKArL
wziSFV2E0mrb92q5cu/kaMkUTY2IYQQtWOgk51pZMqAdvEsnYIgqM920Pe5/QU/HrINDy6Ot4b+j
QGt+SrGjs/qNVQQgzirAiIwj8K0asPyNaRcwJq91oXT5Zt6xhpASusrr+2h1C1Q/MFBiOyONN4I3
wjKrV9MdJxwn0dyfCYH0uqmCNNnmXLsSpeZswHoPtuGIsYSzo6A2TvRRT/xWy2WeFWTJVlLriCyR
CBU5oW/3tv66uAl4qY1VbEMFZfhccTHsHmHdyk7WP9WGfhGg5Hu72zEQcUaiWQSgfzGb4jxQGSw2
QBrv80bQIdW1c//Dnh0ZDOk947u/98o+ElaAzeN/eE7JcwfAMaoyJi2xqCkrCiGXrKcj/u+BZYZV
doDICFJe9PZRxh1Cw+6geO6jk71Vj12W2U87HNFI4LzsdTTFRvN0mgio2tzmia04jHcRcA1aXFNL
S8ZbDK07cx8Vqch3TFsnm/+JO1Sdovi8f1xZrTczNS9zzfPM+5bA0f5nKezi3VLKZiUzudEAwnPa
BrLSjmmqMRw5ZpFDwtZsF21V2vsRl10CLHy99UDtE67RpDbI++7McNzTBqc861OB1ZfdrKIpPCum
AoULzEoEOIHr+YpeBgSlFs6b47unkWAyWcd+E5Gv7HR6C+KS4D6STcdzmp5qmgcg5POkkzesrVXe
AZo4Fc8cgGYnBIdM4tEuKJDyOWBvlUDNQOefrIJslICAmYT+MAR9BRc0XW4zayuSOzvMQyIdUKZe
H5FCyuqoIuKHZzi55rFEb3mOlQljXmoekwyhRxBReEjbneWvGw/5JDvEzNEJvZRhzw1bQGpOcbU2
M8Uk3zmHHKmU7B+LNUQZFqNdfB6oYdfsvoz0HbECBvhoYU1LA4WtPxhcQQ5LY3kWYJar3vSYmSa1
zUEpx8hk56TvzFVBl2bJomWm91+L2pil/gJ5N4OXgj1s00DRDsypcSil6j2y1xr/w/Uth6jRsykZ
My1O6erT5GqEEYcRvYF6aWnPX/HF7EEha7PyLNR59eg1J/TyRQL0NoR5ewcw+/40DIHP+rDc9S5r
0LGKp+Sr1RFdj9EBS1lYF8WFxWzuqYYszGY5D4VUfwKtfw76asg4u7yd4rOTdO6I44epyqaukb2b
BHpzn83IMqwM7WdeLnRPX/uAC3gUUN68lUzzzSPXE7Yj/hxsja6DhAIvhAE2Gc8dWwQetQeyz83c
SDyT84SnfvI4iUw58cT0KHNpDc+S0kEWSSE8eGba4nJK87fPAfE4Tmdi3WSu4UnPbTiOGdSDDiG+
U8GlBk45lfQ4ZHxPZcAp0T7QEKe66oATD7Rxs3bV6NDWRXPytGSR7njEyf2nb4qqhjwWlHfipXf5
Rt51R2pWPFJBZZtwDDFbMfJdR6HD7hmxlKGrWbWI07JvCf6fYD41KDdGXwD0/HhIBJTffbk3hibo
tYV4o4ascaZ0XOpGWmHC5W0SVLBG+ypzPOSIVwv15N9zYVU21zD9wJFAz3/ortkmpm54el2xbamn
2l9hr+yegyzidg7kM2FN6x0lCIyRvh3Wjqr3CaFQ5psHf1LMZ0hDKoD+sUscxwx58ZmqOmEJq1j2
C4YNzRrylWASpVSHdoXuUx0stdkt4gfPwf3KHjM1++ieFS8l1CfEO+z8ZQ9rDYDOXdcROx9gmQfx
zdLCSm4Gy1Y+bB59/0IfqGvF1lQVac353jsrhSPB6n2s0RnY0UVkWNffZWZX8JFaOTQ0enYjIk6s
iZC7YpOVhXrNjEDTRfRuq5L8Ji9Nv9nZ3HYwOJIPS4UII6i7SPT74GPuCGVWLqdCz/BCCS81RhBM
xZd/Q2uNUpP1Wskbbl2lbYAw5cvo4CCxFNzcYRn45jzb8LvAIhKqW4/eOffVl270L5UEKBDScHlg
biKrXiH8Z/Q7cj7fWuUAsjwqPuKvQZMMUVNIfuaICuHdu9O2yIphBJqvqb39lLlDO9ICLlLvaHxm
hkjahwJAsv/H8Bkd2p7UJ49uWEr+Sonh6W+VczMzz08NKMKCSG0j+kZD/bVH07CvbfDe4E26dine
akCLH+65zmuKLPne2R9DtbegvTOG3Jb6dqUp9Hq98E5GA/19XMMjejBkIxJwIcrszI14CfvWatf3
wR+KLtmdrNOlBmTQySBDrvJ6g93Vawg73ZZlxNUOzr7zlGUzLxKm5FOJg10SWWkk+GkLvgXOej5k
+F81Gr3qUDLVeHKOxfJ+3uYehClIoaF61C0fV8iaBZANB5cxjRHNrmBxOzsWl2j8I6+g/q4bh4dV
zfreQs8YopuET9inVg8pLj+AUfBz9CamfJG9PqX6D2g4D/0H/53LlErQv7bHivXSXHX10h6JjXWc
cWKUu6N0pcANYLwqALayIAV70xqjMof9nF1svsqpZyX/DJpHe7BnkdWiwO1gfMI2WNakLy8stFig
mSh5Tspx9ERBZswoP/3sOGwyiM0Le6LZsHE4Djj1ISxswNwiqpiCj5T6eqKUJaqf58+a44M1hyVY
89h/1oXwst3p5UOrFvtUNfU8QsNx652DGMDPOtngW2wcFtWMB7nrM3ld3kJCz7EWJ32YfvRfeJyo
TUhxzakoVdU5PJtegw670D+RIyLFJluISJsQWP4WihqFuTVHzMkdQxiVBtxxztN82cTxwPtYksZS
T0HT35zx8ueSlTLvm9vzJMzdBkf/JEJ6WVwe6ZnJkUGj1UMfMck9rpIdcLUori0IAS9MKoR0QbAU
siDzxzjbRU1b+PyKSOTtRQI4pRJXX1Ip4zACBl+4sgvg5w2MqmJxOYJ0Mq1UDrQh2/gKW0Ztcon7
dQcG1+gwd3RCJPQ2h6js5RqQzohIF+leo4o4fuktJcld1v4Mq3sFGyXBgJwT2FdsPRWhtrWuc0/Z
xTtaDEXco15l04SvOUrubzp46CCPrdZXrPuqLqIRlzBbVYhaF3A1ixz5bnjVrhTuRKHpoUNlkMHm
RCFCinFM2yznt+fsDJHYeZ9P1L4bIZeP02lMdin/1nltc0Amh8RsSsbV88E4aHm4DgR71PQVoF9W
a1OmC0NHWiym2mVGDatRMMjOGD1NqDjjSVMrLqRyQR1pleNj15B3ORcyMzupTotrZij+fhSGoqlp
9tbdt90Af/gEE9UWk7Kqeuh9YvEvvgy7WLOF+0kq4vSs4yPuOUD/jMBVbcGAtK1AUxQWgvQM2fam
2/MilRMXq+M2fpkSw6Z6zVqLyb72TGbsXZO93vhVQlfYyyJ0R1H0bYshae1BNIiu5LXqXKGLFY9t
wWrWfkRwP5PE2wZ8ko/Fbm9a0EMA8aKLxQL9iWbhoeb1M2ho5hn3D3wSfTxC1y1ooofenEMOQQ73
Qj9yKwGaEHaDARvG3n0YVkRGxVzIesaE2UoKUpp+JqKUWarxlRZL/Xv9EQEsjQKcV4Va33tY37HR
I5fnLJpBYuhZ2OIs7X0ieEGYGaD7prT6KJQ75JZYjsGNUjFg49PiWwyhkKsf1FzgW69HeUy34DeG
Ju7nTBwJPJCwxteM61VivOdJN0ljSRHLJqvl09xOoYasPPrEVtme/QpdWni+ndQBwz2eaNvxKaud
4n2dRTx2ah5ie9sPoAcEdGkE5Ky5eUwfplG4WCGF66bhKu1aRUHeWQG6bgkrsFLWkPTSmmx0Bcph
Ye085R9aonz7MAk5hoebjF38sAihqr5nvEOylwlBbPlgCzka/rEKimg3aQHv7ZpRpY1gOqeQ5mpc
Ki3Y5FYKLFamA9yeEuzfmXf9fLkLnRcy0WqIe1Zkrlux3huAt8EVNJ/P2ZtUzRP/kQsAKC4iGToh
5aB3GbDdhGgn9+tFlCpOflJ6CmV5+iDYbZwxSC6deTiKD8LxfGTfCKDcK7Zi58elLHep48lHey4g
B1b9BwGEHGOSmAOeTJrWqpsRWZgEB8b6apTG8OZzoAEGn+95zEG9gdtR8QXWtxRO7CzaOmuBbCav
tymWgaFTs/YU+gBGMa5E67teKfW5l8wb28ogQ/aa8J/67uSaYns5g8lF+gn2UtEu5QAnxDO9nNRg
xglGnme9GvpnJIzNQBwtcOTrLmrj+lSNvyfyNzfTlyw9za9EJzA3HRX481afdLPrSsmRgGtvI/aY
pISN8sW6xeCCR7OnS36b6OJpqkSRKCYDAMeQnRsbXBITTA2LY4HkdKZAjiEbh4i7K0GncHLJpD/2
jqaHPwy3O+rXF45SnDA1+DlSZ5eRN5N+uLZ6ym//iCkXpTl5PhBoyV7b9Md9JWBkHIdwsDDFmSJT
vO9IkaSgxIwIq6DtcghUJ3oxJ7qK8QRlEF+d+20rRH3YHzF8/h1lSKPlP7YjZNdws0zTy6EmyFHF
SQxSpOS7amiQ0h9xqJDPltC9YZqQIhMinCrxWcfLPwhwFLLEUtYtGmuCCRLNd+Ht/aMT5De9NSlA
ay8QFWVuKII+3AfQuWdxYCrTD3qeM8uW/eLFbmDklT9gT31/mIPs2ocvZer2rWgKLrCIYQE9g0lo
mnJRRYQqIFeQ+VxfCJ1ysleJykhshSC48RnG+l78Kqhy2RkMjqA/Ctr9jBmBXri0b0+I09OfspLe
w4lRVtqdvkDMqsPD4reaFbGr70KJPeVA+KgC4QZ2a1ZYWljM/5cOh2XL6Lrg+5wFOe3oPXVlo/yO
MJAIaItf8Df8QD5YyN6o1egXF46oo/4v1I83KM4VsWNcu7VgGwnJGgk082SxHOCsnodHhh4dbSD5
aDF1jDMN68bj+PoRYiOECMVDEAXomuDqaAIQ4WCn4AMWzZ6nkZCjGvtVf3y2qL6WYEXvmIy2HG5a
nMeWTpAp/FzglnE4qPdTU+aeQkiZK9y7fwYgHDl/qBgAt8lfegrX0/usTTKT3/kX9ahLBhWEIji/
Ee7UzXetoWlfNt/CuqWSljdiqDGqZhqI4tbIiWT34EZpy0uS0SdbVAncNcET4cy9UfF9hVext4Jb
1p82wxTHpHyGfWx1iwN9A8r/QLw9IlrzV/OYh287GMo9gvQ4I8dJuItcjo3E+ul+f1ZPi6gjthJ8
CNdzzFGRa19sQ6ZEOqUNN1tnQy0Fb4O9AAoCqrRJlGJ32sOYGwbpl2OENjzYR4bOekj8kYPR8hc8
fCGF+oyEJcQvkQPJH0Tl2Wn3zmNOdxvbK5RjVfkX8O8V2c1Gv1oE1Gtb78/mLVluuk6IaOtsfRxR
WYIknzcSUIe1XSJq3+RPxdM8NxmDX/CBSbt6KWO1rBXF+0r043D8ZusAKSyvHNyW+lKnbBBe0Gep
jSi6+R4oFM4h70Lx9dvNtwl32RYZhqbrPRNLcmfNqfV5oKOjL/ILEJQqI/JCjv6PcSDHmGqqUGXX
3cVVvN0t87t3chiElizo3ZEXElBs/rd/pWEJItORblVvgDD8hAcu7yD3fVJ5IgSo0jw2YUj5CAs8
BQbBznEYw8ka5wQgh+dz068x1tOL/63xvlPqK4VtRmUsnIMT87we+ZgSynQbEa7VFD6WOpWCzwKd
WYNcrtQ0jVlhmd7PzbrXoE02cXimPz4QzGPr7dQxMNSwtm413Kakl+BdhJB9bj2EiBmsVTNy93mm
SmBQ2Io4ARYCI5baztHzOaApxYKDw68zi49DxX1ObMuT7R/H5n9eWNYjgMUSXnVp9h7vtJYtIFjq
1tbUr73Q7p7SdBx3BmN8hiyF7u+IMvTaZButtCnQJ3/7JKe7r51yN3P+ckQMPjmfyQ1+VlxSOpYU
AcWLv48Q/Q1pom6LkVZjGoIBrTmhGvkKiPdY7NnWGXkjJqlY6mxEalbqsue2gx56ofce/1CaMdpl
aUJQn9qzP5uFzLBoaMZqPHP0Sr8gruzpT4CBUx+SGBfzJ02KzAQl+cYSkWZ6XWrXlKSJfVQFVUYO
uMj3wOrmncDZXXB/+l9ptnhS6IfuJcwM9x3LVF1rDCLBSNkN69l76ZN9HDbQlT4QzDMnWF+L55S3
bCgGMs5wqSX6/fvwMLxWAmfpYZm9bfBUMkOkoAlM0CYjvpzGTo6tno0zQVAk86Sbjh+5w2ihp18T
VH2vUFwID/8QImge5RY/PrVQyS+fCcKR4hn9HYdxVDtny9R6HMG6Wa6LJEjRfQL1gAfsJXkVQo+9
L14ROfkLrClLhA2RRLoay7aq1JLhULkGkG2oobkCZfzVxrMH43g7P/BUYxzaWoEUMWtLCvKrYHlj
JOknNETiITdIIbqUuACZ84qQQ0okBvHB/jtKlsCNgyKNq+dQHVQNrZuLd4KSTt0paRH+hZvoNZV4
ODIzLDcurRE7Akjt/rXMTW9hdDxIuEZGJslx4mbXgJalDFWLPA0vXusgNBFgAy4eZTmpsUIcHzz7
4YSAn2Sq34JTbySFdjylg3J/tKRNeDz9q3AB0KUom3BqWrUJ6HLe2cH6jJzEl92pSjlwc/Oij/N4
OHLrVfB28I+YuFjpkkI2f33tQz3zg35trp6rbr20HG4GXBnkbAmYpfA/dzGMl1H7wX5GYREyPUXx
9y6wH+rBeRuspyLjA03pUSscOIV+/sLEtYFql4S0RzWYoC/6qnSWAf1s0+6e60nmpO/LZrNw9lbk
CCroosmbrfoXQ+bTJCJfzREsbNi11XND4ZQwyHi0DZSNppr2KERusVclukl7Frt+ctG1zoboHN0a
NMDeLmqvSHzEC2plgbBotyKGh9JCNLNCGnvrC1za7ggQD7b3aABapt4itS1wOwjN1JcDeH19kZGu
EijvDXoK3BnL/gcRy7tFO9S8a+AipyUCDSv4GupZCzr51+nlBTbiSKlOqNgPmNlmIDDFwHOmnUHb
r+XQg34tZGV3ZgjJXtenQjvWWV7ncqcdjSnc0ajw+BjcjzB6/igcDvLU0EBaDaLep7xNLNVZVM4M
TJeE9g22G1P8u3RxxiX6/ZCEoM1LN6IDBiOKhmSHa4VvUmIOafXlib8cSaf4vO32IdljCxCBwQV0
jyCvQkB71Vutfi0CPjmJcAT59kFhGPs99mbdh6ys3+TEV/O+wInZr1t4FRwLhxYtvvSkicyuhJnI
bUniCvDj9oqf/dVlmbrrF5gDmGBcWJRDWLtbeo3aqvU0lECS724M87bFunaTE0XfPjyynm5cY9vT
e7UA4FXOYXGHT+drUSdDO9pHGZKjFEhP1vqfyXKNKGFQDEgpa9cgZkfPaa3e3Z8zgPmQMMN01i80
YJlrlGXvFucf0Vp+eIgD+lppxpx3cHPragMm3dVpaO5NX0KaN/LEz/rf/qtrCmwNmpk/cSuQ1Awr
N4AB+P/SOnNoRQ5pWnxod1FrWZ4sbfbB8r8xI4MYwSN6CIr8uqJ2a3WnwnHadpCCemPs+YbhAYlc
uAmPTdeRABgXxT6N9FwRphCCHmLWJQ5BFWNrrBlEizgRFmXocb+mgVhTgmdsYbLCO0K22zlASwWI
KPjUIuR9gZ3Z+Ddrc9x+mKAHmjxEAKh4yY/MKz04KDCqhZYsyIslHV4QgdKTYgdOIjUB4fCy/BoV
gloDipgTz0kPRraipUCFrUG4W0CYpAf9wLyQe+Zm7EMNKH7TXL0ouJeVxNRuBzTjuCF1CniLcGrK
r8dykiEyfxiPFjydL/qIjNlIfcnyE2HYYiXyk9YRtHrcuLdDxoAk1F8cHEEb85vm7KcvGB+E0OjU
oyZvOjq2lJ4iHUMrzRJAax6ay4JD8/GwJdSvdinukARM/vtzXkomxzjkFqgAADUVodoIz9qX0Ahf
akDK8PpUI99+gz82i84QouoEXq7R9FZZgMUSnwYhSN/PuG2ZGXecsjkg/ctNifZaV40JqJ+JmvtI
jIoPZkBoalc+fKpwCS4Pu1MMOb6LXSEzZMenfBAu6o7ryLO/M2R2KbjjJQj3d6ATuy8Lw5W4rmky
3PHzN0C9vviTKVOqH4dRjF4vyA4V1TVk86Dt7M3kkHeVMs+8+aJxTDE6OxmbL/AYNMMLI2X0STu4
2MRGzrRYa8KCXDwcGpf4ap5tuFJYBcrgsEXb+MmB7lF2YuB++TF+lI8F8twZa8QwLbgdloRGAwj/
1p/ZukMr1iKz+JO8J/sC2lWtfiS0m/cQwlt8biJSC6uEATE2Wi703LW7K33CcNqYW7WVWKTeSS9T
DP2Hkxf4cmdzy+Ferd3ZeO3AhAKPUKNQakzJxI9ejrDsj49VdsddyVU+3GiR696JQawN3R3a7PjD
W2cH0ggNikkiBHWwfmpWsiwwQOOUpXKjRzyXrpUAFgXoq9rZ65iYx7JWFjbc9GRk49TUJfc5eoKZ
idpM5EHylrlliS5UWR6hjLLILiKP0CDX7ltncoSt3CKBOpjygpOqxP3HUapoy530sBbTiuiyt50V
gB1aEWArrYSbMF1cOaTRrccdN+ZKxZzzvE59UdwU58kABRR/62C+hxunQE+K0ZYwQbp/yRScpv0H
zTKHzhYwGD5OtuOyrMmg/KQ0lBR84xTGl6gPR2j43dX4e87bZKzAvJK8SWG9754pOWFlC5RbmRJN
B+sADcHRfBbpXWhnSSgFY54tEn8Sp2Kmv81KyMJNQh8h/w/1XHsuCvbsvioNFRULOADyGdBAqJef
Zje4ISt1S6fgUTFvnRoJPpAmyCA88v7UX2ZsBeORECdUdXInsiIHuKrTog1XVWT6lkOujFcQbcsN
MG18H7Sq8vLUO28BZ2+qGDQglusYOsWQCkF1GeLtbQgdiTefNfijjPf4uROY78ixwQV2WehcfYZm
VHeQ2b1FfPfmQ3r5tRn9TEs1v/BlNbIBQdQUNggvPMeWqHGl/x6xXoSK4OM1Gibu5Y4tcXadqE26
C0aA2juodXcYwoy2FyxJI7EL1gjc944Kph7I8x7BmXRjRS3ZH2EzmBYZC2a5dNr9mZoQg3Cf7Ldw
s924xd0+RUx1PmswFxanHCd1n9+JP7Io4oBPGNMVJ9D/vbMhewPYozaQxHTo5byI2xllkqF1tV+M
iMbqI1x37NNr0WyFScSDFiAroP8kkjthxkQfps0nw6750r+k/EVjb1WSu0T6TayI5av6PsLemQhz
Wdteu6sFhngvDFxr1h8nWF4ASCW5UR6xmplsio9Q+4ECHqB9MgGrZTvfZ8vHwYJjmsc0n5GTcfqs
pjgMd7lOBI8DQU6aFEp4+FM3xA/hSyX7dwwb9/ZPV5AfexVhVfxI4BW8bS2fBi1EdCxlXbUXqDEL
lMQitwCJDxf9JWLehButbw4BNyrMd1T1U0gT/06X1G+CekS9W0dtd7aa4NAGCzn0ssl0jPFX8C7E
kpx5okC8H4pzkls/ImNEHH4z0M+j2veBD95Dsdd60dXB7DVQSfUBr4mLy0sd4v7tdJSmMw3ryUIj
2V9tyKiGyQjWAfIWtW4wv0xQXD4T1NsRs/ZqqtsOZiwjrmnu0Z93enjPtLx8K2yQ0NS1DciQDAuz
m8AMVHilTMRCGHfHVLJUtJOfu8P0Irv0gNsqT/VlcwfcnOSfLT0nWSwKyIjlvZW4WO1+lCToHVDG
1grp/ySfJCl2GhSwYGXPlSPbhwPTU1GS0jIovukQmeVjAGZ94mMezoBXQkKVbt+euNzulVXjsjDw
556MZSbBrDhdI2AU4jn6BpwwBosDMC6MZMtretJEtbmIrPBe4XYRVH3ULionZbRhok3XzpXkv8Yk
mUhCpT1j1E362LVADDnCW7gAjpX+50ZhFrRAi3FbUSvIjEZOJTpjPLKyvXwnt3d7d9VfMdZG61dR
acD7YqZWjGwZYz78j1crUr6QqXBNrsFt5T14T5f5ERikqiRIYXPUBaMBhd8nweOiDYPOdldKrCko
eqKNaFdGHuoEIaqL6VStULAIXcAe6Vye/Mi/8pPWFwuPpfYVAauF6IU5o6g5k9CJxZ4E+7Ug/DO3
ZmbDyyyf/aWOruZj3mAnOlxSpF7vb9jFngxfQHeLMCQNHt5NOuBBwmLZjG/JfVfLXwYRsnntlZeR
QzidpVQLBHcWD8x3WOqyxYVEwKrDvc2uFfpDC3+m2AQ6WZ96trdldI5LClkkXtpJdoyHXYOy5FcR
CROQB1AHNceiPlQzVoEsgwN5cExj3VGihU5RYQpNFRn8YiX022ZGW92N5WNBhMwrEIazGy7ZDEWZ
/4stt/Jyv6R+wUjcjXBDmuJf425U30/tNnj7W8xhIGnuqJ001swCA61UcNlr9W0GSXwKKiJmX0OW
CDQb0ax7/ynXv8MgJ3V6oz5k3wLrbR5BjLFa6NiXUpQd2FYnXvndppDKJy5PyHlAOYQFS6SRP0My
VdMk8Sosl3Tj6ypHYJ8YlszkwzqDhkBWwOf4cfVX/6+QY/eH43JyVZV0TRnIhAcl5j3PIaXjnwCN
bpgFRdcAK83TDzsyMbC/dHsgdyL48jkFNOgLfTW6K3jCdN7jWJ8OEP+CpPEEZsfuQzENN37vQ9Lw
STZWArl8B+xyOCKY73wkJGD5tx4S+uBf9ifV4vGE8nSko5LCrWbSbltOiWX0U15l7q3AHIoCx1XV
wF8gpfbrYtFco44UFPgLIhk4zRtm3QcsfPa3uOKYtnEGqgoC4YQ6qqLdlb6mV+cJ+tEjBwhUeU8D
FWHuy+UxVDoS6OCiiKxa+kjWgPWrpqzcGvVCjBEx42AVSM/4lL2FwwLmt9LfWfyiPEpnTJwCBfb2
Loxd/in6oFOxO2VfZONQ7FFUkWa5CQFf55R3hWGRUyubJLKm2wdU3vsafGtXwnx8kmZ3eoCBcKs+
AL40uyEY8F/Nkk4/4cd2Gzaved3pRTKyOhoDnHWJZABEXMEKGuDo2MxjZpM2ZmvbOTs2l+s+DL0N
8Wj6/GJifLWZnYJUIx8C93GS/gjK4VB6IBVe276tvhsRNsgP8FjlmEikyIhsTQer+E5btIL91KT1
oGQCokZMEKyZ21xrbul8voSJjBQTjjdQtj+hNcy0TVuiaprBB/ThZ6fcrCurfGo4fSdP2ftovVS6
VagbnicAsuqDiHuB7l0tdIadFs462Tzw7g4r4zFbP8utO8WSp5z6Jz+II1aP5ZyadiyvsOb5yVJS
y4FASf8OYwqh0cUg+Z7d91MdAxaQ0wllqTdjIe8jFDsTlWpkTJDtnE9Uprqa9Q8NT6u2tjT02DaR
gBu073kSiNUnDcSDbYlqDFq1dW5MWJC/6fGm7b+Sk0pA2uYpleEmj8Io2/Y9zuijTPKnVru9xS6x
jMP8SlQn5WJgwr5KYnbjZ3j5m0/vwUM8JJCC+RAsds32C1RuGNiGb4E418mF706Iz8adzqoqTaaY
rrtnYUhqhfnDwTyJdEdDxFoZEOskt+R5uSPdBFe6h1i3thqnYRm3vJuE23Cl5YZurP785FboOpZ4
11v+G77/6eioIEf8SPArxv5+4F2W/TyfflgqCQiUUOAos10QPDzwlGGDNOfGPR6WKiKQ7+CNSlD7
tEkTE6OK7rtMcGSs7C2cFsC7N5iE234wzos6U5Iohv8V1o7aTjzJHeYLyuOrVd+Fy+cLazb1iWhR
nLpmbS4fxBQHEcK4W04M9ZdRsfJojKAyCyUZ5fnQIj/Q3lNlMuBYO9HhwZAwMOUo/wXuoVid3Z6W
jGOgqGvBgP8DEPYxH81yFl0w5uiGT1nFQVtmd+3jEjh6hOMGU89i/7qS8guPO7baZJOjtQ/MLQ4v
rMK0qgbjQ8SAwHynSZI5FDFdHaHBOuGubJRlPAUFaBgwNc0sR1rtDkgW9ei5COFYo+Tm9C6g6F/Q
ZNmIMefdPNoFKQZBwxYnXax7r16oM+NqlLHn/ICS+WqMSyfwc2R1SeP/lk64AjeCRlpr21aMfbXN
Jfddfzu07mKa6UXMCLpYfZKhJVBCrXKlaS8k/QYhoL1swz0DZN1XBcgU032x7rH7n95aQar0N764
n3z7ZNXuxZcq2GGxWMDXzEJ9WtTaY5MTb8c3zL5H2NeHKT4GpZLtbIN9uBuRy7n/2fgakBL4Ti2s
J7DZwDaDLu/VrB/VxYqZvdrGJTewaHmh1UHwQTfGfRCFz4Gpx3Rpp3TdDoXbrfToowabKkmx1u0l
RAJcGFfDdaZLBJcesbXPYJYifk8kUhm4itBjxi93k4Wz+Ok9+/3SjqAeNXaWvhmio35zaASMnsug
7eA5vKquBFjBGOX3MUVfR94X6I+KPHymrR88hAG5xWdnHnEBhwEVWRHHQHnYGhfWPyy8Kmbzl52n
U5fCLrwXPsy7fD4Zy/snsvt7ngiAsKoSVwrQD2ClBCIpjhepEsxZQxoRyiwAI3FRPBB/RA+pE8P2
oVoen+kXJsNGYEDXy3VdER8S9a9jXYT+QFlb17nT2lR9Ii6Nbs5cdQLlqQnwOTwT1hBDOrVPYHmB
Szfw+8PMUA+2JEQ72mgnzp4WnPRavHsJaAe1jwD5CP9r+Ra89CAnaPK7eqXg8ox/OdwQ8gxBBKIT
rCqNRS1oCN7eKNWXj/mYj+6978XDkMVDC9HtQxLwBDoC57fY/x4iANyswSk8bp9ldZaYFbN90pbN
fDJEcCEVpOKmyfdH1aXkZE5FCf8wAmdqb1IdHus3l3IrFcMjZRnbH4nSfIvPqNpQiaZPi8F5Q6zt
WFylFr2OupsQaUoDxsEfCixOTC9J80BwGc1hE1zLxL0aAYIYbL3kyDKW7FyuWpP6k9z4FN/AoA5x
KEdmgR31jp+QzIM4aTDk1tg/mOB+3EUiv3a0QjU/K4Uz+9Bjif6cFuztgbyEblDWVL23BD/jmIqe
jVnPe3FyAnhFIUXMe7OkI8eurY4d54hQ7QK3BNG8uIpR1mi7eoxBRqSqbTURRvjDK7DzEUmqCUOU
aYGgIDplpS8eqaSpvvZhhp8tz2EKIZkipY0BvYNwH4gU6Le5MuxbyIGz3g/G2oVzbVCYWjCfXwMD
SzSnuhwzJIRAR5K2urFI3QWvw8y0ctNe5gGnx7D9p+4OGBRnKqYIw/SMXjOXN03656TjJsCab3mM
FvCHuwmnB8ubyhggmeP+Cjd+j2rIPdeH7V9+F7UyxAKiH68zdEVegy7b5/FF3YrqZWO0zIkav5o4
kpW0NAu5sHrarQKmd6diyCA3bMQ58Uf+UJMwcCY85aQYAdnL1ZB1NM8jNp8JPxLa2sN2vslau9da
tjelC3zykVhf1DHcQvsU0/y/mTNXBiIGjqT6tcHAKh03/2SGIFQ4VzGA9CvssD5vJtfDIqMB3dGI
TajP6kTmDg9IdiPN/47elx+i48wJS5UEczjCkQqWbIB2X4fOVsKid85p1PzCxMJJpWliI/bFTKLD
aU8/T20uJMdFerCucV6L3tyGriGoi9blXhcL/bKX2BmlG/Yug/hUBgkOAM7f5TgUkCA4mvTIV8bj
EDtF2U+kXriiWLZClK0pE6wpGtqOSHTJADs9xaj7kDpJ6p3PRBYPdFHYqhg7x55RGCPQZw9EoOv6
2ysRyiAlsd5welLUb6hjy77t/L0frsGd9WXWnYeWM1lsM4eQLcz7cTYQiD5l4G2IdDgMHBpff6l7
Vogf2ucBP8E9FPK608XGRib9B0uhJeZeE36VAWyX0kXoK0es/tGxpVIRTQ4epx7H+7K6pXol9dg9
IztPQdg825REpiukCbp9JwX24D4RrIuYUfJERv0zO3RP2W4m+90sDTNDHNoWOjft3W40K7YZgQAW
6xxIjVFakT6T6WNjCBIt3dPgtUF4h6wT6PzWxSKETMiV0tscsq6FMfVllOCj+/BMAs3p3fWhCw7v
PNy5RjqMn2rjhc7FCJ0SFKY+S0WAp00KyOlVRGUPXRFhUL6RGt9RaVBuHtQVMTCbwm1SQxC6gJ8/
mzWNjkbW6bEArVRv/gB5PlW2Y7Y2+phfNv/tO0FagyuSiQWFkkMA/u6ZLUBd6HGouxN4WVDYQmw4
qCddrqwgHwgMiOsPfnHWQedZNKtt05fRuUPy+E/OmUSuEXbt/MhHzLMbG6dZrwbeDANbh76mj/CL
r5izmPLBC18cbtjm9jd5MeNGilXGwIYGYx6QB3/lUYZgWbscG5gnfvMgGjg/uX/vM2WNKwEcSLxR
/HEslIVbU80wQuuTfXzswhGILQX0231Waw/wQD2AKDG/yGTbykFiEPS0oKas0i3SBly8/pP0XW0m
f0/srtzDysFG2ZBLfwg4sleDldUy30+KBgqNihEefAJM0We3X+xcOBPyIerChnOg1VqCTulcnpfd
w0rr47LeiAc2aKl1xlBuRINpeqwSuG6WFc3n71dqv1q2JgCwooTOz1/RW8g4giWv4azvzN5Wy7SJ
lyYD/JRMeAlROHLCQCNNbo5rsn0ua2O9nYOpAMzvRjZ8PPbBqNmTrWXNHLt9BxZXpUOneHUsFcre
izG48ozzzNRLjSx4Th2v4DQb+Q7r6/RGnTXAbQ0/LwS55Ttexpm1sM+JtwRW7Not7cIy5FKJixGd
rNz8aDEBqK+ISUtf+IbvDiNxDqJbK0N/dXjN1Ellcg93YaX40vdYmS04o/ABmaTQcSJFTKbaqJrF
CySTsiE1GKl9PSdOZOCa4Q8ZYpxGgeshLGqF7y+4EniNHlUJyAN3BmOq5YauEHdWD/YEBZMiEQCk
H2vAlEKAv/23q9aExFCrBwfwDGeOEILHt7wOlWocDbB/jUn934mrdSUmKMUAZFfXVYPTpl8a8dlc
el5woZgJv7KwdR7x/0Bhh/H7HwKWqC65MsfjJLHT7lGMXfvj1lNrdNkY2M5J8XJ4qW06e3TJNKlA
z076Vabq5nx1Dr+6Dscc1+hrHGuQaoF3DaCQR01KbVnDbaPhhC7HjMVgadwxgBol/ZlsBxFIDAl/
qxOQvlxsZdHyd2orzDZWFfzj7gAMWMCw+8Z+Mlu4zA2BRBNzX+E83IkyJLH0tlOvtoFaByV0RYno
FSaWBvuJnkI6qJI8j32e6CdtOhhlhNuJTghURI2DJojajJJ/F+Yp/UbJA9w8c/qO/WneEYj74w1s
x0xfu0Alh6oWszqkIibJiBPEMK9btxPOsoLJSZ8DeHGNYKw5U25PIIj0m3krCQ4iR3urwDsXw//V
B15He/4RKGRi0z+2Hx3hhsaLRoOnMoWbkcvd56M1lZ1YK1BGzjN7C8yq6vOY60y8C2KiKOCL7eIp
U8j/VHXd6SiObYrCP97eW5nU6NZChybZuz9BRAkN/X0jHS4PYI0tw95GyN8+3GXZSjBSf9To99oJ
RJKphN6pjgZibBkCWac/l5HgtRYMJm1XB447nua7tRtmNQB+ncHzi6kNtFPRqceDJMpP/6Oy+yvZ
X1JSSPeu1uLepnfzNn6ZRPVsywOSCpfmJjJiOEw1YuHccEdGfT1z7l1M2h3rJLugbwJ5D813NBSe
HL8V9XMtcTb8WrVbIRC9xP6Cc6N123DhtFzbU+DSXJ48ZzmmkoMv1hA2n4ZrL0eqAr256JnMHzaZ
igdB2Ulu0RMjYEqcRgrMj7BOM11asFBUyYKQwy072PACORYAgnxn0QXA9KhFCRtZN+oEPWrfzBxK
95sTwFH8FbTr21ObdJxbytxB+FiYb69hEsLu+gp5gIynQFvyvOgT6CYoUkQum7PvwltinIzrMj/T
7pa5yQCK9qQBHwPrEuhqn9y81ASG7kq9dKkCgBwwOFF7y6U5Kqz9g4+dAC25Qj05GN3eQhn8J7Ay
uk4ODooyTtu5wwyyHNu12v10KaoLdGL/2ysWMgmFoVaj+XsU9cCiagoVLrsG5vhl8kNSPy+EaZzM
7N9MPOmRqafsCW86HufaRr8WmMTUgJnj+24waOuOinIKcEVSjMTookrxnmgvEKR6X+Ckrk9DCTo2
sWZZ+4eMVN2/0MEANcV7rj7gcbCjMIvTU4tZ+BpZvxta2hUqsRp9uSexG6jAaAKOzqhSCM1V94xo
EVIJg74P4dkxPEVAZsKsEwbuXw6g6/RtqS98oKYUVCecAlgib6S++1qCeVyPFja9BJoGM4Ypx4kq
76pYGFptXfuazcD+EpMrpxWgwxRkWI2E6ub2gF0zgLBSjUmSbLg8hXI3aUOV63lTCwfFpAyL4raJ
a/avB+AUxgYpx86QUW6vaIgpofxiDVW8C7HmeQd1wl9n7XTPf6b2k/xWyAvRtXRz4bvVfVohLI8V
7QVjmRwDh/gjrh+bRjVdC9Vm4ihGJfLR59ZT4EPRS32TI64hqyvkqpac4u7m/AO+H7ZxaTzZd21v
g1+izRjiWQ4sexupepAPkAe79we44I3HzmH3Sscq0OjPMC7laLMSevPmSsxFJiRCSb0L4FmAQB/2
wK8CaG9vblmnQYtcwjhoazrZOb0GmSYpipvQpRl6wCopWW//mIR2zhap4Eg1dM7JpegTd5c4L4FU
ZHdFIerxyS4SIRas/yzs51tddVJ6FE+0EtYCKA5DMInwOqh4C4Kdoks3En3BRwaHIAeMwnp7xEj4
x8JT7B3/XLvLihXeWr9t3lPw9lrxC4qGInCgS/NtqIk2haUpZsh09Kwd5kn/knEQhMUqX7B6UO6I
vkx9ZDlTSgGiGrBSs3x2WYR1UPKFiiRxAHHR7hmO/QYPZZX+xcQEawKnuVZl2QE4VVtjKwBMREfB
5ucMCwdDO9JCUYVN05xPZXpzEqanudup3qUKwA3MkG1ubqjlu2sANjZrn/Dc1+dfBQDW3JRWvLv9
bpVA5B0T48cru0XYHD3xUzPdnp8yLH4lkY/kcjkUgKfviJuRe5qIc2AAcdaLBFnHJsueFQIJBDbx
+Dk1g5FZ7vh1F1sc9TP3tvqYPdbvnV/ocSCDN5F6rbgvqrn61qqvFo+4jDtFzk09aER+jD5jpHA7
d1qKW+Ofv6uAc4zuEhtaPkNcfmtKeWn8KJQnIJPmNn6XxM9wqfEbktsXUBqPG0rSDuJ/R42V9xOV
0vkoJ5PpMhoGwnIDmOl/yFuk3vV2wqDYsW+Xn7KsuNl4fW35LUn3Zaer7WyLIheOxVY8Besa9pVs
XzN5eNZjif3rADZi3swWMLhhAX9Hg1Aw0X1HA4dc4iyjcLsWIQi4vNitAPLz9yfIYCOeyniJBXLu
htxIWwYQKXp52qzn0D0GrBbTNju6fMZJ4xy2/X3RluZnfTAmaipzzr6vXi1FkTeW9yduBDpkIW/3
cvfAdK6bP+7tgmMWxp4DtR62L6/5I2WOFQsTjKmB6GN9REO1dGYkmuFL3fOYUP15ouU6of/9ILI6
n79mC9mjaPYEcmBFhQOuTmq7WPRBB2fadtVm1zCsvbHOkeDt29+e9GDqgy+a1yk90RFKmiawzO8e
WH4SJQ83CwEK30RlFRPCqtFKHnSUpgQf1vgNJtEUNo15b2aWEykXgLkqkDvNQYmg4VDa+zGeH3b2
eXO78dW4ZRTPa9rqyp1fpxV+CEk7bDyLPfqwGEu34X6f2F3tl9EoStlB3ZZCRfuWPhsyKGSo2xcF
3r8owwpkZB+U7id4nkA4SjXF2XPsW1LkJO647GCFrLn8eYdD2nRzbVU1NunlC04psB02NWlqVrqE
eTInKKpucnuA6B2zmP5tk1yva5gv591sWvX7tRDYy/SfVGCBaGGnUYu8lHbkKUxI6soYKrgwa4rv
Sm0IhXyqw3Js4ypeWPWDTatxFYKQ6I4r0WoZ+AjUptZYhSiOGpM9yVs+gf/693K6+OsK7bcpltWG
dmxt68oa4izzrtFUJdfQ3u1Y3qgbBpNddQqh9gUSeKmGEynVwz9DD1N4Pec0MUiHzABPMmweeyvG
78E9wGdT7l3KXhGANOpr6lhQJqbF+UDUndbRBjN3v9PpU6/qXIH3bF9TC1f3f+A0NVUceVUFrv3G
S84JbtQMk/ls/kIcqdOLg2jEFLcxwrn++PdzPKI5EWGQQaMlbT2s40gdPsld9LzQTljT6n7m0jQg
ZThu1LQ5nxHlc6EXWdT4NrucyDM5SLX4Ue9TgiPZJ8rEkxF3apbDzy6ZEVdLvs/vW6m2OYXbd+QH
/PkZNi1rEMxaEt00rigVBb7CicHYERyfUOruMHgi+hqaskjQFJTqsk1gynKN5qJADrfiP2cAwfHP
z9JRMCYMT7YCaEy7vTMbFRKQ5QB6jt91l7WJ66ia03kZoB6Ng8xYUVbsqnVTOqtxWVzlx+PGcNVw
6iv/QcNv/TSuzdeJkqB/qCTzYEWXAJXA2SO7N8QZRrBcLc7vjWjiB+Tg6uIfUhPnzQ8P00ilXQuh
BzXfcERHLtGKV76ni82bO2h6De978R0eyTjeq295UrsuBreC7Ckprw6FsL8FgIg6sS/4QvXds0JL
d88pVp5+ZlSc9uNiviUdjZZ3QZ4NTYq8nbt7BJ6LMPL/Mdt8cSPbNNfQQBObvDv+5TdUlqziRrDr
SjSmDeKc69h8APlCF68+NiV/MjOaG+bNvBKIYSQqMdn1u+XJlwKoCeWfDOjdFFRNXTleRZneQDWu
hJOTg4jyVbH37VUAqCuvzuvx6R4G3rpQsgnc0NPra8VGPsXdo2k+KPAOaUIIijCw6//U4rPmrmtY
itDuRlBuP6WtxfIT2wHDc2SOo9szxopykFqAxPY/CO+pzTl1VwK6AYPlvzI5g/prbgE04sPpl+9h
Zfje4EAV87JZD++ae+4GT/rr40YkvwiCOsB/7bDy4tb8JY2rYBIP0fupdFHobaVCdNXDVKQTafVq
VYWn/Bih3U0i9pY1hnDAoU4Tpv42FOpZ7SwohY1LOBvw7+LtlSe3ihQQpNEpLWfazLQtthtIDpvN
wbwiCxF45NqruzF+uJUklPdIsLq2aqdggtDPQsPL80OdseStQzy3+tPoZoVVIjrhXxfiddCAKXdy
sRHSrTX3yO1NPRWi1KtVNOOxIcoas05UGLbVJ8aNqt6FZxoenJFjQ7kj7nNEQJndAkW1rg8NPsMd
X8p9q9cni2gUUxIczrp9Hdn88ueGAQfaHjR5e45Tw4Ho2Xr34rRcVOpOY4MzlvXrAKETj+rhrGXK
t/Qr/XdWAzUHP/8wafZkLOz1hdEAL/QMRnbj4iT82ETsIiklzgHSOEjhhCRvZaPWmr2bwXVLctcO
hVcH0ZxurxlMxl1G2VVqc0QPEzJr4IuUgm3WTzSUk8TXFYSuCiXejlSygH9FPUTFuqaaGCTWnfFM
InCvIpSYG7vNaTiqVsWAXw4Q8UVWc7Hf9x93Xyztr+LVlcocKCaPSERjoRRIHr0jekCuh62gQi1j
ZorL3GQaWwsZmYPprfa4vt2MKlNIXN2RmtxXNbSdYjJbgLxCKSuc/rbLuJtWNpfJes9duljLscBv
kYiOaR81bXcQ190XRq3U+wmn/ntZ2eEjF7uaCEdkFavRhc+D2PKh2A2fSxZdto+pzUpslESxvTxk
hisUMgt+SJmh8a2CLoF9KTU4v/8CoyEVTSbK8L0Yqi+VCUTFyve8KZ7/9Xyl8NkwNo1lv7i/nx8k
YiEMkavPAFA/ogjFlcUhK3kcclZBU9g14KuIiKyovYfN83JmCW1+053gI0xRh1mZ+B38WHpKOI9E
SHdToChOg1yl57rpkVCoT6qQnbm7WMHdKgIb/lgLLrlPcXTQfS58ggx1iLSpbOMrqv/fhCjJHIGd
DWvye7vWFfrPVf5mI3Dkn1VGZ7kT/K4Tu6wpwUt0OlEvvbhn00avFZf20g/RdYnu/o+L4K6Affds
+aMPG2UkXcJppVSZSxPMPvI4KOWyixV9WvKq5vWdPIYgLq1GnhkmnAEytyFDQIjoEC+BsYIwlg1M
3kY0mgOjNeZHKJiw1BeAmkGT+SCklrzMm/sRwA47GIBc1ZZ8WgHxP+LPzMuX9cNyyqEK5Ob22YI2
C6BoLzboRQSlL8hzZxAM3xll7WGxG9vovoL75l/1d3WYIkIKeSUScKwwbu0HZes1n74e8v4srqsH
nIwa+JRSzp/KuAVrBR/2H7yyG7uSwD4nFMs5Ah0DgCTX81gqF/k8AxLWRcsjbKhYAtHXzCoFNrJ9
XvjHMWN9SOfW+MrJ2HpsKTMxGDrqgwHQgOaQolPJLLXLqOCI1XiTvKikHunc/rHFPwtwqgUJmB7Z
DWB7i2BSW5g52UwsqdkQwVugN5V0vF+x0z0Slwt5LCdJRXJutQfx4SbB4SnEZkrXx6O4M55+i/A9
/YRTbHNGtW04nhNwxQmDCFw/H9rVVhC/uGUfxpf3OUmBHS+2eLE7iYETMdbZdpYQodZQ9HPS1Ihw
xpardCN9NZ9q78q4AUhnBKRaaXvDCI9SdKZ4mMUtvra+qQ4YcFSwb61eXlwNNHnuPMbRTmd0mBXn
/tsiTba/FL9i2Q/x0rPYR2XMCfNWbYu06LfqFC0//yNnWZLrVfS2G0hW9ZIozdcHNN7zLQrdDra+
MxcS6/N5RwJgMqCIlDDvWn83LgCq9GPfiIZgqcwS95yjAI2+e5t8iMWqiOt0AZ3Cc504Pyo9Giro
kKD3vtvwuQgg3ELb9ltQmtXRvEfAP+VKLE0LVNGgoTcGcRGT0HbSlRBYWhhIRme6CUTZ7G3tPe8G
KhrgteGOvMFYQD4rHsSHqIRsSyMUJvf9XI1wTkQhzHYchCocwZErLmdG7SNtuESutFwXzzOBmjS8
tYvlU2rOBP/b73pa29wIHksFTQqSuu5HtDVf6cyugqM4hN+n6NZjNz04uAGOUGaYcRPuppSa1JtK
+aDg05BCi22ztfiaqV/H/sMl6ogaVISC0eG9ziAnuulqxSjv2StiNncrS2kK9QiqKnC2cKv/uBpI
YNI8aExMniDgHrboaPU+INoJAc9yOSpsUSvvrGmnIbLMDLTOV7kzdMTtXNWQrzySaXi3LGHLljD5
qLN4z3an2odmGBkWDUC/5tX/aL6V3RUlJ/slcKYqIOe9YPcFeuZ0G4lrfnTnFpJyWQ8bH8CD90nb
DPrSDK8wFMl4CffqWMr9AWkEungm3S0CZGDFeLqKslpsStqOQxPq4C1xLoRlrRRb2Xv72uKJrfxj
H+mqpdXxiT6Adj37z4f7Z5yzAxrqYwzcPdw0tRsyqepu8y0+rhe5iuVH1VR8PI8rOkm/8TE1yhqQ
3kI0+vuwtnx6I1xi2LhDmr29ZN4E55y9iae8QBbfTXjWRpRQHAmgavm9tKJDV7h/BHvE42WZHEZe
ndL9TLp4mlr1ICiPNuj+3bJTDsbc7f9E1vzbtOUuo3f2/JYohiFbzDK01EJSGHddTeuMJOu77kba
sEg8Js8M2luKqrFM7y7k58gbJdS2fqo/+GytE+hIXc3h7AW6MWma3du1ODX2KCUnRc6spFvyYHIw
3CoM6kfCOOe5Pr+MtgZ4swp3Woz6t6H37Wcyg1wHF2fuKJygGWLoAfb4ttiVvadWZ3ZkO0mxifGs
Sd1VU1ly6EflvGXDmWmNR30J4lqY+tYr/PQVdOq/T0l33iUr4UK6nkC890ATf6gioX/NkU5bcHG0
MnSRqExhrU/mPxDxOIryXZOzkzvweogtTzEYloCem8WIssy9wo3Eh0Ys6j+hUqUM3d0OkKP50+bz
OloXZlzkeYzX2p63C7rUDbAo0RzJ7Rti1rzrGPG2q7VFPvQ0uT/4ov8Z5DUX4zZ+c4JTl9pWBitB
o6p5OAiCUjUu8FEGX8Nj5eMvCg4osYU6TysWDlaNaNV01w02mS++ypCqIhdeNmrWON5HN7BLzqZH
ZhryJY2P0/T/wOOfuinfqozRaMhYB1HGClQ1nbjYElYuuoyxQysxNGODEW8I1lv2AmXIoN8YSc2t
SE3xGJqZ3D7rQUTGWTegAl5wyVhsGgoZeew37SyFNMH9vzX13tLxPxroydnXGLu2t4D028TBRgFP
Kd3KzTURlUilFrvYUQ2dd7TAP5G1+1Hf1heBGkZYo/VZgDIDCAvKdtpYs2LrsUF77p55vzN2gvtI
RsclXgLDCghkJ1lnmO2hnXwIfKI2xfUTmSQToovlPK+D0q00KWs4QRGhkSUSX3deU1MjIdEdbsyK
QmwvOCVGLHydPmreEyWW6Iiq4hCba3rLp6ZfBlh4KiHjPxxlGiIxCT3EGd77XoUbx6uJLFX92+tt
MlKX7uGmK0YFyGSrpHOuP8ZQnOvn+AShInlC7X6gxP+o3GALYqeTtsl75vCIXJ01Br80pOmvP4WW
wFOC9nYw+7PBf/4hVRbKGLp6xLcwiyPxVYIk0G1fKaiIxHZvKEa5WSKs6ATz2vKJgC8LOKG3pMDZ
aRkDtT8WrU6NEvA/E3b6pAiUKGmhQWs1RNu0KdJIermnDSNww4qPtEyzz3SCYGjMbpwX2iH9byT7
gJhnyo4yhI9DMkuwx8I7JBg+Trh7CMnTBUsMreVdtSJtQ9DXctIQorNPmYS5IS6z8ybKB8V7f2Qp
unHgcp55DwZRNIsAvsPIicUHGV+aCJzKEmXBa+9FQEp7dSzUGielG1a9I9Em1imfAjBzIcSySi1z
MxS1t9nwlRyG4DVF0YWYZJyJbOuryb6CNPc0JfZECPbM19b66okYnCBIzz1SHKYAnPqf+ru+Vkpq
/ljUbBGxfk9RaC7wG903w1sPb2j0L+tN6BHTpFZFGxLhdfbaba+Rwl23oRV0bR/iHMltvyopQjGd
g4g35h3wGucFZqe3EWnE3HGRiGdp/Tf2rDnmYxmV6eJNN9Kgg03icvmG79tnZNNC1ZMA5xDeIUqr
0T3opAeXvnf4h71T8qyaUyEe+xz6qxLIqimOVfg+j8zNh1gcxvda//GGhx6OKG4s16IM76WN0Jz6
quZtCGq0h7MeB8BAXR3sD8y6OCRRfV644/fif+mxaY9+MzoZt8ujZnmIxGvIr0T/p5GcqNDdTJdv
mlbwF8kmEzEO95XGFdLIbOHQc/jsGmWt1X67oU6l5dZfkbiypegCjSmYC4DIEaSBdZfIf+BIrjyX
/NFnSoNjWFsdak6rbGv+IJwiNj36ksJiI2H/P2nAkzAPkyEHqTdUcpnDRme9yhGJShMttX0dbdhU
9E5zOhb/TSFBzzDRwYNJx6hJ1qfIZOHvoCwl5XiiV3IMkDPX3N2mJDFlfE4TBlhg+1HrSKqQh0bt
zTp2k/7VLNgwz20YKR2fu8aTjm7kfiW1HbAvbA86qUs6EWGiUNVA6v7th1+l5NnnGA+CRAxhIw2j
2INNSicILZSBhAQeb2dOI2QqXgEWhlfgCcMxKKQDUIQDDxhEbdL2QYkJJCAAhHuOOAMw39UIM7wg
dcrTTSVjgJb1nvpwT9A9gq14ezH+72GH32W3eveiMnaEoGVonpNQYx++KqH6+VUZ5PHf6yr3IW0u
aGSPYQ1aIcu47h7FOt2JQtdEdg2OnrA2hsi/802GLuD4SFLW4JS7aRinGsFfPty1XL6Oo3bLe+3n
Ab6L1OD4nAbOPq4t2N3oHk1dfE1saGbhcWjtbJ8VzbpRfDGf34rV1QQhgC8GSdlX/UW2ywp/uy0e
DRB2yys9Uwj5/2FihTasrBw1yyGf2pV6aO/CAy5ecItzKS+NdBf3MfZCoBXTKs7slxMPQFIA8Vxq
uVaFRV/2bWRfU92zejR1jC9ovTt42fo/9qB/zJOQR8X+hi3IT8OMOfEw8fHP0meKD/ReEIpLllYB
9BlZcWVSOSWkAt86Yb+3MVb4TgiTZoHH3682m9TRHNc7CxLG3Htq9ex/LsiZAMqeZjo+a7Q2b29L
/rb1tN7ilX7Imy6gE3AWvcP0lrNEhz58PuDT2fJgnOnBSvh3dQdjSPQjzqAcPcP+MKNFiEvBlyYY
yBZWmtSzCpSvsxZD/dr5Ric5gDz5iOEcrVOIofj/TatT+7FGZ5Tljfpqj8zxuUhJPBm+NhC+UYIF
WDJhP2diM6M3ciKtDN91QS9R7rWRML3nA4ZtSE62yGUhHl0FjYAS7Y9lmhXcEk6QWlauoIPJVPa/
I82BXsxLW8yw1odOEH1aibpEa9QfqMQvrA8L4an0OXJsI/trkV98D7iP4+dcs9r/+5qusbhuXdU/
GHKeisiM+5hwEL46IOw6jLBJJuFFN30VL4sSgw4kmpRoxpiXBOZRfxxoPX6I4P3kKePCQxIaQ38Y
Y3u/arvv5RJOLAowNbgd9bWOCGIUcv3PNqob331TxPAEyaQpB9wftfq+VxfSSnEtvE9yc4Ri58Tn
0Qd3SW6QqlRA9ZuNJQasacD1Mb5DlCoVYQdFosjBVr1xEHsZkwVdDuysIKVVQCHX3DgSm8i9KQQ9
5URE4SVh+ASeygj22SWC+EiMs0ENi/Ya7l8qIaA50RhRhxqjEvDZHW9UfG4a4tUVSByTbPId35RG
kSM2CT1af7H0VQfzZoUU+ItDqMhLl10xWD5JT3FOBgxWBg7xZj10B90nXgeLSPErSzyvSu9OZdz8
L6nQS6dv6Kn0dqe+f5xb6YnSOGw5aKW28lghgiFmTKwnEHJIkZKIfKfKpSPU7hW4GaZpdcG0gSws
Irp1Om2wUKmGjUsxKL7/nDuPV9gLQFAepEOFHdXjnk0b7ujc4cpfyF80XWEBYLV+rY9uMBsEbXl+
D4Lpa6FJUUez2H3Wx3zL9kDy67ZlcGPoS87XMIBatk4iNX7+VzkNPl5o+JiXyHkVh3oW/SOglK1r
jrbUCQOhNFmjj26SBD6lpb0OGTf1Lzux/32rOiAFimgfLl7CAUgFWsiwzj2Vnstt5AXcJBiIKQg5
tL5FS0txz5oapcwdCynLjFFjW9Oo71Pty7w4jVlcx1rnr3+6UtLjnxHwAyZnsFi20ybMTHCZE05V
rEh6Xns/rlwU1rJ22wL61DDH053xLJgM8ik6EPmjuMJnUQrgqgNVtn9p5d+CT/CsXjV7WMUTw8a5
HHrTVQW0PL/04YZHicV2QjBj4iV+iXKQoHQofsmGPHLNsPsw1XWB8otZiMEOx9SYXeKqE1X6QnRK
6laa0oyVSat/lkaBrQ+D5gV+CvdevGPBIttLtgtbOXfZ8FxkGCoOWlvoMnP/PJL2pl+40pcezxli
ITT0N2/AbIBKXY+nJLgVHH5w5jRCUPW/FBco6FWEVblufgRDRcRv73F1z0aTTXQLtFXWWYyeyevn
eWa2SQ2gw2MJYlQW/cmdoanIIqrqgDajMJaquxKnFAlhrHbuxW/c1oBgOV9C0q3YSJQyTfh+mGHL
3fveUNTnEE2hMjYRC83m1TziahkFnYQTWa+/c0pr2mPUiEHBIHW4YVnuSIvvYhl378Jy2ogLfb0w
KRJ10PA9Fpau0T/m5q1wNvHMTKB7hGaykpn7N85eacmZjj51BZx9SXA1IPWTa68Lu3hdH4DvalMe
YEGik7WN6WdiGbbfUpEu5N5446b1oCYo7wJnIjEShqvT60S0q3fERpmOYzxB8eLak+IAzgvZHG+L
EEbSoC0TuOXHpjhXChNo+Z87FJFbGTys1TkpOSTqPGdjv4vugcIOA1+w9zBgItNfi2dOk1ptlICT
1ERC+ey7nlrLq9pqWttidYbBkdCxCZZs4h1wDPMaLBcBcGBTmcPcGlvjyQElLGDXbdjwgbQ3UHUC
hRtLjiy7gOCL1EzkF6+6dYx2cjvhIqsboT8LJ3AMHjiF8N+izTUGKELk93oTIBIZJbF1iVyQvns8
ESqQYwfgN3WBtGZLEGYBCOCP4/54daK/sG8khXQ5sOo/ShhPYjp2AgJqVQP7FH9Qa1KvNxGSJiK0
Y+JK+1XXS5vya8/vXyzERtJ7jaSr46FyeUWlcR8AzHVSMpsUe2HaAVBAWHQO34DAWAyGWUPF8yD/
bt+cvFFNuKWEQ5L8WmHoLzRW7MpYbyfvcD4KCzOcKVgVmvzNrfVnPXi2KBWGISZmukILO3C2HuKL
13k6xN6lGf1uRCmQVRk/s6Z6r9YTFNhXGfBAuKa9ueMAIfon5waMEfkSsg9H8SgWiVlW33EVZLns
fkqjIJd58MGlegUGB0FPlc1UpgTSmNy+f7ANKVELiGZ+nTn+Sz3Vf3MZdV2MC1MUxGlmLI6smKM5
mj66lGsuYlh6ebAmQ+yfZ32BHuMGRLNUTrBQzX6LBoh46wmIiQSfq4c+/xGZPUwFrhz/vIRH3c7D
kX4R35rMTOkQtGgABSXKS4JiG4wppI6SkRklJ7bu4o2r4wwOThHIYLCXCyb7oCZJL54reQBjUN1l
1f840pGSWr5ZaOrKQTvFUing1LCPIQM1MzkeZ+R8BaIeSYyZ+BqAbjEu41OFkN9J65p8Y93E5eXt
G3Hu5BMKORsHnx8gLlSTpWXgQ4FVV9A/L0tuATA71IbZNsN+cxty+tfPb61YOopzVftjYNO7y2fp
Yuy7BMXihtxMQ0ubXaY8C5YSUa6hUEHgRwHHgJlmrphyH0ixKIO0BnYVs2XxnGJZEoOvLQ3v5a+O
N8bsuHnYlj5mlDIrJczdC4yFE1Oc/Pc7dq8UQRDStEtiAfw/Owx2cU4eTbv6+YCN3+4Co7Nlk7YA
QPmpcVgrGtkKWn1osdxFd1NT4YNSHElA+0uelu3Zs8wZJwGGbpDasm4yJ0If1V2LeN/jQJdJkZs3
c8UsBZskBHX1HLMtGj1lypqZrv/bjLh6cV0+0i72P7nSVJhJ54ctHfS3aNDSTkmj0Uv2IXjGrFDy
0xHN5HnqiigHxWWYuXfOerJ/uZCGYznCc3CVg6PaOPaZ8tVaGcmPubZ5zbrIHUmWhaYu6CUGHxAl
x9+XHGJzd4t8dy3gmdixrHD8V2cb/7BBFDDcjUKDp/yyESNyTITVNOSiza9szSFHqrx7NaiuxVpA
rq63obKFJzRkNSuHwWxEpyxXr5SlgFt298P9tc8inifw+6GFS6uEe8eQ+ZfkV+h9RPFrjOwf/cfk
zkP5fAIQGa4xHdW1s0iHSMVIC/B8Igf4qZal3Fss7TlNXg97jmezIsDjCsFgUa85rmJtTiCH86OU
wXagrW0yG2xMBi4C+WUir1bNQHBiFJsqZHcBCaPH/FTv6FnmOKexRN1IjUkz3/yDwnGmA5Yf4qpD
99INdbAATvSINueBrNhdGEk9rBsOqTWDaC3bOt+sljzeWsKU+qoDQaRrm8eTOqh5EOX6KHEvmQz5
/QggqEAehBfWBx/U+6aaICdaXX+O4Fuu+g0l3P+Tchlk9SQWJCL6T7DkMKro4EYs1VbRIxuTaGCg
EmjSumeLC1S9t6zkbC0pqekeZQO23J8NL16UTSjQ3WE3CYswouS6sQQfraJRTcJAuuCis+k9oCs0
S2sgFgCCSFu984OuOpPLcmmYfo3tNYRE3UZOMt11Ji8NsdAO91cpCL1GE1uX6ls96o0P7EZxwHsO
DDmV6ALK+QtkjdYGfve3s9png5HT0pFQcUNYOcAZ+JCpQg2xmwJo2wAmoIZVFBpD1Dm+i7biRk3i
jdg6H5PwZYMP1mP/yxblLuCA/0pbN2mqYEqDimNjXEQ5bljt925ULkiA7yP9C7HnQDjOfFEssgIe
550upTkTyETAD0BEwgGRn9SJNq9sA9so+GNwdvdsQXI2eT1EIBB5dtYrmPiKg1rw5wXvSXBrN1OT
J2Y2QdoQW0ifq+H/Jha7gVRudqAkS3psYSfjKU7eEPjL+lmXPG4DANuTEbW9wsgNBQgJBls14BW3
7BRQ5TQ9qNqPokvfwYfkQPAf0wu0R/smsvo8r/AW3/6fs5HpOVX3jTbhe0YkI8R8aCD5Jo4BQbpO
8LOkK+H2I00a5HFxgK+RAcQd9ABNDcPwCrZMfhe1CqKf599Fvz4GK+HED/U2Rln4uXL2Xkb5kVjP
loLw2e4Q8lccyQFaKIHvWCTK4feiueAUrkM9/gY1IlBUe2zSXPrIcpBfZPMjdTeuNykDhaX/cWk/
qW3Sf8xhSV+TWMbSrsrx7TMax8F0HjZsFJv3sUPdOlQeE4IPMk8IO8jfv+N+I8oYbxBwKwtlFA7J
FhL/04RvjA/9OVRh4jpu61c/EfkDmr0M82I+WcaMNJv2zmka9ql8SRqyFI9FGANr8bHPXjge1MWN
v6TefeysxF7EMPhCfvgGUB3/uIbwhspdIswVXlWZODr/iv0oqzhiTimh/SQO12XT1WCXv5BW0Hc3
hP9yJ++zN8Dy4o64uqSqgqpe7Eb+pK0sJREp2+jOAUxHNdLb9OvOxnI1ZsmFn+gP7k2Fj8YcFiNf
OlqJFdcyr+Qde+ZETPTHVcMRHwDXO7qux2of91a5QG1nyPzLSh7cZI3tCegUNb1EWSiocuiZEswy
Cb0S9Q3CLQUm2hb3neIcd+AWU4J4pAgkHuzFVEypKLHRBorqTzjgOuqxLDti1E5AqQrH1etA5gf1
dxM2WUz0POH3VnjvoFViuYZ+62NCvTQ+BSzzSbUuz8fNGU5NJfqhJH6Zr215pWmY3PUNpo0BMkN9
9JbORPxjmpltRLv82GKMYJmJpSmE1WZuu1ykcvCnKn7pFm0tBtHC8JY8HihmGAVn2yTgNOjtx7xa
Z5EmV48LouoRl2LLs3w7QMxxlmbXiDQEV/dFV7cVfsJPydMuTxvRU1wNWUqGHqK1aPpK4QFWF9pH
C/Pm3TnrALlTlqX7TDtEwV6nk9v+AC2aHBtCaomeO2of4Qj8KLlBpFfBdKnCiGc082mDaltqFOKE
U4sa8HM9BjVk6rIbfv2jpgY+kvBUmuZo5ekafvXh9PG9QmrbGO0uG3M1OsdsIkjGoViuwswSghqW
Om+ldCcQUNmFValDnNikerhY8veymA19ubXD/wICE1momPOl53ug4UmiuiWVey5NxiomGBQpx7zi
bxkYkzZvVhBPOvdpDf2QKpoSvf17q8sx/JPfp1NMndvGhq8Ytq5b+MjP7E5PgMHLEVHo7+UfAaBU
QCbl3hO2GNOVUZtEnzTe4+scE54L9rO6r997pgiQL7ix86rmzB65K+l9V0xa5KYYF0wg/xZYRr+z
tW6M5+EwnyfNv1XR2g4KK6U1MxKqZlVVzJ7Wli7IaX6GmeD5snZ1lCpdl15MYUBkzSDBDU4hgbmj
Gx9KY7cIBLR/adQTMvYK/pPaurvCg5x8WZRAPvjTCBomxaKTqv+30dAbDKTaNs9obJP6aF4jKo2I
xxC7rH8mfd7tJvGEHozxj7m5jyII14PJPbD3NWBvl7r4L2OdtsmbYCsphbmHrwQ1v7idkNYHO2kp
HDJipfYUA2EZcaT0ndSp/Q0BIiIHkvKaEy4wAuEQQUQC9+z60A07gYhLubON5HOqCVLFT94NHEbC
VGV2nlblSaAjx6ITFWFCI/ZCEb7OeyDe+nwx2GpK0Mx2oFwuj+ylaN6vpt/9Gx14v45S5lgj3Bp2
D5XD7J/7zgt8eXVk8amx06QFSLr4yZWXk4qoMeDPtRxI21lZXamsuf5mc5QMy2wQszXnYw5+/qWG
Qh5BiB0TjXp4cpse3wF8ooKdTXGQUo7kiH4VcaSaJe1StWbRL/pZpfSkVgwUDvNkwdlq7Jhn+rFb
ewtogfF7Rt63cqs4vG0iRLWBYiVwQvtEVHCy+CoXfrY2ZS3tvg7EnebGqNxQ358GxdYAUSeGgO9o
Fa0BTF/E9i0bXg5O0tWErNOzAUNeOHSpAbfthg7hxsM/oxWO2uG9vqtc/wIARuYxewAzkMHcGnqr
eOy/IHL12Mhi4wBUXGi1VxkRb2B2Ul7FpUu1H92m0sI1DdIkvL+0jbIMwMsr41pViK8Vc+oyOSuE
lkG5jYKE9e/llDsSb5PFT1bJTshDwx0+soKH/tAeVB0gPvRnzAxKQnamxCmNhApvVpMYFDWPmGoZ
OsKJhX5LDaiK119dkO+cYeJ0RQ6ajMNrS9e72z6vwM98ljxcyS1N5jJH03Oco3lQYVh7pTd+/3ze
I28UlVY8hKTJp1LAt0nQQE+NJBmRdZSgs7z5qzyK+gTUIAetwi0cNiUMIlZteiiOCTmBsVgw5mAQ
/cXuTY/BZEerMRaYLJHB+Q57t5NMawUYzQ5wY3CtoVU/E1UF9hrdU/0oY5Or1vdBqX8SFYHSu31C
4TxbV+ZehmGvMfAmyHbfOM1/xh9Q3C8VdTXqwHEIA9+1JtrbPnNsR8+erRPUVw50DcumPS6MHVrS
b/23fa9qqz9tF93rqBRXu/lEQBTwi2CAoF/PpwO2WSEliQhUA2yGTeRcPcpZSUM4EE/vYaspo6rA
ssXmV9RSyD/+rR73AcFWq+bwnCQGM2ItRKlMYQgH3gPy0SBu+HGQFSM7p2JV9nkkW1DEX+5oUHqq
ULkC+oZfdOYf6btHp/Emnj4wkEYBOaiQmX5O5o8AyAfWEPszHxH9/l3wDbnIL7RDlEx83/eXii7n
CceUwTJ17/i6+3kLd3DEMFQxhrJvvH30hvaTOFhmwzSw+XdpBWjt2HhhlfW7aUDjeA9ToMghkdQC
GnPD97HoijJsvcOW9+W3lHzgV83iVPXbcORd0VJCz13L81MWkehtMCMD+LEfnKipxyU7kI/WULcY
UYxDDsJFSX4y6Qj37kuh2P87uWsgVNUoT01eAQAlFQEzNLKGOYrzHFkYl84x1EF3a5lM5h1bHRGI
NuZNEwTJr1qvdJN+O+/jE3Eu2W+xZ7zlxYBHoGfLHQcpLnJREpMdWN4sEwsZ2zql9cR/rZjz/2j1
+vRIuj0YuIj+NiJUTYCQuYDA6ngwBj+W8Pz5zQ64GZ7rDBDk/N14A7sfo9AqhsqweR38Vmo/Xn9q
KWDx9FMo7wQtWrEEUtKgiSdBqzbl1O6z6BjKA37ecO6Qr8zIHfQBT8LtHqok3REYx4HByMyDGhgt
fAnXWTiHRnGsizb8rtJ61JKwyKhF7Sx8/AOOto5+fsgV5KQJ94n6hGiZyRl77pXlkn/yz4v9roWX
MjKZnihb2aPodB9AtvSBl1jODYasftJpgywbyLoXeWoRLIlzaqRMMgqpS83HKSnnktp0t8OTkznt
1zG9M8PQCOqbohOqPUNJfjnrU6ZaGSkrkTs4XkS3l3OI5uwR/kAUXFeatBEFh6SIpNsW3R1kqpzb
fw+mmozQ8yqezhELobQHghKHNauI2hjBQHo99hRKROqOzJxWR00B5xrFus9/Dzgejr+nSAKD/iqm
vDvkOitb79NpEw5qef33tWfFcubtb7LgNZ068/U2EaNahZoEK5YoH0/tUbs7jyagbtutJpMHSfg2
0TBtonuevA0PUvaQEfPYi6zmNLLd9Puj2InQ1Bu23qGrZNMRlbzvkSECy9DL3RbSySFzui9xlva0
aLAtYmHjvx/7Ic1EKHtQWd/qZFftdxdzxslLeVkxJ+uun9YAhBgJ8jooviCpNDrL5BuGYSW0+Amv
W3H5d/4GxZ4KLyStUC0+pPemkt+WUkcgfg/yIvzANidD2Kxw4F8XPinNtxWYeeuEKEsEC0JoRZmY
8eQz+UkixtUZQgfNysQho7XMinA2a0qoQAMq/BkRdNdQ/axJpR6s0k1NhBx8mnEF/EWZ0+PfJ6YS
uE5qmVdTGR7BOh1nSzICrUs3bnIowai0zzl7T6tvpznn7eFabkG42mcJGd2+pluVt3A5yipkuH5c
Cvit3wOX87hzc1yYBQb638fOL9A7C4BRIcj+4sLCA1zJhR45QBtIMY+OVVkSKKkmidjBGBJXiShJ
NoQ8x05PRDDxwzp0pN2zco4IE8VeX/4Vo8b2RZ20QOxOGlwoIygWFm2Y29tGN5dp6ocRKnauVbmq
9eiddDHgUDH/lbQPG7QH5M/Xan5bMlu73Wbn6b06dJFBY9C2YFfgJlMOtMSVWyAcVziDvepnfsov
RRMUy2YfttudrSozmjLtEMytgvizw4AV65YUMX4S4adUasQ9kfdyFaLHpT/g0nJd1NjE4+1Qb0Lp
AxOXzIbRkvLUOFC4JuCNPp+XhqFStTr5lt+/Po34P6I3IRurORra9QyMOuDttl61oOmTWJZNPLw0
cKsxgfTVxLD1n86gZ6OQI/wWqZTf3zasp26UTQDn1X/FjJtwYZKE8y0m/CTeQoKRfiCig379+glh
oSMilM6ZW+KLabpFnl/hFIfgVAvCiVdNCAX2CPh8CEt0X/QsT5HPQsTSVulWpFOpBGgJxBEtZRvR
SH2O81FGsC2XEZoMPwASngMGcrPWEN9XagiAq8VZcVUQwyVbmf8jI+XojBkOOaHzBIcQA9CaHIlr
oNeWaFZ8fsfoJoMlRTSlbupZyVN/781ZZAINv8BReBnpNqh/pVUfWUuLb3EJY6Revstdjbs3ATUp
zquf76jux9nnq+MphK8oB4f/dbXo3Y/13F2BdM/eDIyeVgo8+/MFZMCg8HADWLk3KQ1NZJ0Vwnqk
eLQexkSJii/hMMR8dsNU0ijFoCeAGCe+oEE3bOu87nF9ZAIeciVqCSB+JXJ0TTxITmJL50gR65Jv
lN+/bXTp2FNBXawPeDPzr8wh5A0nLSR+Bk+U4ks6l7xzq+Sr0Uw7/+44Q/oLzKgEL/ViWnjhrCww
SV6nU5yp+dOdaOd7ulpZgtDfyZT480cxss5drfIYTYd5oFSJ21SqSTWGFUcGVLvIPhL41mJV7xsM
mGmc2U4+DOluLEyfVeTgq+lqFIpobs4YYhts3rUI5LvR3J85aprv/T5zlkILdLzMzOlPFD7LjqBF
GMLnT2wt9w9bfVnETX14micjhAWZT9usQlNEpfW8KlvO2nr/JUNZm6TrxsqsB59SrcmYKDse9gMH
GcY/ifJgsgr7/LTZyWNo9XFAJPHMoocLCT3CAMm6W4LNG3p+avbdGw1d87/bYHywE7K6mdSGW5Ej
v+whxfQ4MBI6iN3OE6RYMxr+ekO7niGMiSQao70ykau+zOYYDtU4i8elMGuZv3w/Hlhitb+EZtVy
vwdYIwvFrTwH+XH/n5PlFCXxwNCajTkLVO0wMYpSQQ+KgIEbaAtHTVN3TTP/wJx+hZlDDYyfKBS3
SjWRRbyg8PfcXvJ555iDDaQShxwPFhU7+DchtaxJMrhbYo9Ci0fNvtZVXgB4DymraBOy+wNT6QXj
VA/DfXLAozRb/ByaXs59RMWC+Yu6G+MDFq5mn0jko1cXQb3fvPtWRmrKkfnIqa7iCYWhbfWdkrn0
HTzp1eiXxf2D3tQQiii8+HHyqnCN8ErDGOSRMAWpCP5yA3AdXvHB2WAaTJxkSO817COIJNreNuD5
iiFe2viQW7HkNPhEu3i8vcl9+U63qPjZLBaxH+jKLl3iyS9jrKwjdzp9Qq8PdVrV8riQJIbKHr/p
Rk3oCNycP5q86mW4VPsIP1fhU/SiBz7jIsF3mzlMLXSeTt4a543duD3bGxrhXzdljth5LlzRH2Wu
umFtOoNBQrX87KDWJ+1NlLkxhOwZICrqG9+L/q3pC3iDJF61rkOvQ8m7VcfmMfhUOEry+9CV3OEh
dX+m0eyK9nxqsS+VFY3p/Z76S6jwhiTjgqvEsfXot4Ll6PYUa1B7jzE5u14r2e4EJwG+Sj3/7t2z
GSa9WO/EdxAW5LRAp7byFhScONPvaKun5C/vW78HxOonsBFFeke5SGUClY56jW1SNbm+ju/KBT+x
i2TEGVegHMtjbjM63CpeRutfOiWdhKCg0Gjh7sELm1QQFgeQ/AxPGAXjWwzYzfKfS2HlnZby5xLg
2aajazpBXb4QuC4QCRAfCeUD9K6OX/iPpuGG9AzCADMoWZSck2zZoY5eSiAQ1XG/WbgokOvmD/xd
n7CnHfxWJi+pVNTFvP+DqAl0qe5kX9VJdSXw1Xqap2TQ0KNgETfCmyjhimuvQEee+vJQIHxaGB4t
+HosT5P8MnBIJfemMwJoMdkH4hURHZiS/hJZyFYYPkFBcxmlKmXVa0o14s7wfN1TWXQnRfwMwFjj
+Fca2iGOH6K49KsZGrComGjPSY12H2CDX0n3P3uD28zcykmgVRwKrsQ6npLoMNPDs4ZB2VXJy18K
dGOOxKRdpCA7n+vWvz0hqtSJjoKZuusI4E7kQpSTJQkT9RxAoIP/nfPhF6lmxpX3BsGg/jyNSlNo
ahjsivjRqpVu4w5FJ39hEzA/EtvxVpywtTH9p0L3+1U/jMR/j+9zJF2hDdoT8IaKg7RNN7R/MM23
bRBRmmjrrb03POHQdQmZig4VHQqjINc0Q/moWBry5+eW0BTrtWY8X02Z+9mfVOU1bdRj1U6GV0gC
Y28JwBwbzSCDU3RdoA98jInoEfmP896q+YTYDWDRNIKS8Po5Xe5Hv1JcWHecJMFzX4wExhx7stG3
Tzozi20D8hklgsal/uztWkHhu3hey3MjUU/u6IjsGfJpxlX1ESGF+EtExrpAv6ytqFCVgopqnwpc
bvuqlAa1tAkbUJsH5Csb75ijDrxqQtxSL7kGQPK9N+GyV1QvH7u1DwMqgvUwXwtrd5L5CgSJfBGo
fs0yRhuiqbQRutyMYpdpwKEgkOr+5drgg81pXvA5AmkfDRvK6XZQ38KLKivHx802J5xn3p+vHcH3
S/WyIBc1BsUv627ZgRcch2aOTo35mpQsvULYgoZ7i/8oUa7Nye/S7EE2Isxfb2JH0O4LAaEEFaUQ
JQp0npNQtBRIIEE3zFKsbXyQy704h+6RyV6YlTHruP5DQhb5kiA+hRoH29a4vH8LXm1F5QdWOuKu
4wyY3aNmgbkpbUhJ4U4spx/2kLPSJtjEPY0aWXIJLyBKnIfpzvOR/8SxoCqRQ5/z95chZLrLBqBm
S0agmAyoWaUN0fOiL4AiD/W4VHE7YoP2GCn32n9ArEJD3CvnnbiSqXtZO46XQgZltmwAzEjZfmkS
Sb/FoLyUk/cT8Qf8UqNCGQj1APelpoWUGfcI+Xl0p8RI61seRer2LEqI23lP9MCnwbWCUV3W0vy8
XSo3ZFBItc+ggujF4STb1sFPhlvqfUWxG3V/S8+6EUFLnd7hIS7uXuQ9KI7wYcBQzSqsoGJGqNcY
iHVu246TySxRfsxY16ZAR/+nozmtumd0mLLmXabqkyoQ2EYAsLBalS5pvnm679zeqGJQz9FESYf/
+Jy7iZcu03Yg2CzSg3StfhkgbBAghKeVcJ8nD8cczSaaj7kKV1hQplHMl61FahKC5C/20CxUbf4w
DU4VgYdr+F8lpcIfjaSbaOP8t9Z2E9QizA+118AlGq5AjGhPwzZ/PsYKV5wQJNRnIDFSzWjE9M3R
HsBlqs2I7NQLayrMMHaIk6uiuSzclz4TZHFeQ8ACe8iwlES9wMzgpfsujfSXc/xJpEhVbOxsqZa2
LymBf9Q/+VY9CP/sf+CZVP7WTbaiUPlQ0AGl+jdWKaoZm4YdM7l2KzmYf02wbSCOZi8JoRuHm9U2
t6WRc2di9xmTA8fQWNiDCWkNdATj8C446nU9OdzYnz0g+b8nb68li6fGCl2GVODx2XVsPZJAyHGD
kTxnaHBUW1da25wWLq34Y+kvMwOXoBqnlwqbS6bCvSPTTYv8fjNN5vxuD0NWEeatz48U65/iiSPl
4tVnjgvdxvibg1GbGgvCk4uzIfqMZ77N0G0kvWOCuqlrXQIXyPiIqOC1KCV+9AOlXBsGvZjqUq58
nBjAvnAoAxJrs4RdFnEENncrUfU5Dpq95q+A17tGwJwtDEYytMODCMM7EBnksnulYyl/voMo1NwU
/8BcPNB3Y3k/fUmMM+o1OCBgWNYI9lFZXIPC5/1VpIM8HdkeCRAufQT2G0fT/NDgPiwOzelXxXa6
1HryORsqJOTfPdUO2CK2CcSGgT0eDOsnmZQBdLMkqCqw+NsiCFP6TmIvG9x97fdMk0Xos2EXyHze
dkAOMbIDXhTpOUtnj6boaMVnHhBrBnJ7D5UOoqrXsGM6Yk8mWJ63x8xXC+8PgEvSOXTTbt8I82P/
IvwTsuuM+CN4tDYvFHxfUXFjo1PUDNDoMCX/N2CM6ONpxiy+xF14UsfE9FfQetK/6G+WkVVPUqoo
R2fWqCh8qTZrzHbqv2Vy3PYbC40fzAEx5OOlX6bc9SoBh21sTcctVGk71+hJyzW+W71iXnF2T92f
Yzvd1DdvUumjBfPmVbk1qqv3fGKGabOoiSxfN/xqsVVzIpB2hV4XYLpJYpf7a1aaf4aFKxneAKp8
OQKuuYIdRIDzs+88yYuGnIMbYC0dZ+OGfifelBO8oQCSvE68srRSQNf7hxo4cL9dsQl2qO2mZaHN
0ELZrOuTYClX48V26WHE4goZpuk1L0PXD3Qus4ggn1638WtxJ5wfhZLfAguitlVIvQMV5K8Ad+LZ
O6VF8hW745yUjYwDvVz2mL+G+CibtqvIC/eGx6bfgWtn2azngOnOZep2W+Y8bmoDl1TsCHpu2LQe
QAXoqikzPyHrK/8vYzqbHbLuis3BauVb3OSnhKRFZLK0UYBRtEskXA0ZOHS4Q2ZhyCAWA6Pi2jyF
fMWbLjoVpJ6ewwJ8iMQb9r62kFR/vK75WDsgWizoaf2Tm3lPtzL2L8kerr9UelyYS0aFa4u8f7NC
ZuaVlYmlfQYCQpvvs6/RWiZZwIjAd/NKmgIBV48W0nyUm0IJbgRzNB1/n3WEh2Go/3t946U2vo2w
VqxK1Oc7iJMTlCQ38dXllCVCkBhitI1l4yZyXhtgzQxtsbsd2MFO0kv0mIaJEu6AQEUdWj+SI9dz
W/5H5tBMfXBx3nwN2137Fu0ZP3z04N97UE3NfjQDyeSl2RzVP6jmFkobuyviPNHkPXts08REjJ7S
FgCBedShb2Kr5IgQ30v23ChFkX1i+kk8jVF+Ybg9qSdiaKqFDvmU9jVG4rz57MvaGpq8iTfRvHsL
BxZ1oYXNtkDabvVtRfla7Gl8THAfANUA92RKTKaUMbikcwt0LNPIvkNRDpt9UJIg97aOQpEOoftk
wyPwuALIwLP9y6EnSOqf2BwGl+QCjT8yrqr9vhgJ3l52+XYNKrmHh99ysWhG54nUNX6aBsxBAPI2
LuXZoerYxTiLzc2/jNeFfTENZSdPyiq/4+MD7smPBZggQPCVcfQC9dAbyQl95MhQ+yPX8xReV8e6
9WheFmc+7W6PvC5KxVM4rAcMNc+yB0is9GiCQc7UUdsJvYesyvBrfnI+niayzb5SXrzGpZLa3vWU
ZHdNsRtAqhzDTucjxxrq9uBjGhqmvibt2q+VA4jCNpeP+pSXAhkKxe1YvN/vp3AncyebIZxeCg8n
KV1b+g3fP3moJkAj0YKClxcQ8GhGBfvWFgDGqZRuJrZir1Iz05Wfh0uxLTYMGegpmZIih5X1myOJ
oymqr2kbEwEOJx8vwHmz9AFL6hFuquRgvtqzIufUrZ6qB6U9FQITlfDu6F+gFC/hsrxLjenF5lRc
Jsy82CIneSFmcYGyiauZKlTFProvxyRNK9FC0CC3usLAGqQNEEJEzh830T6bH0v82R2vsetUIyWq
Y3cnOPTl2edPDp42TrSnHPyjx6O3c3/xcrxO4f75diNjKfJcvOWRpXnRepIsj9IyFALemJd30nyH
eS1O2TnQqx1uJvAggwfwDpA4WkzCxrgyujfQUmOF80Vpld4nynXyLZHKQTIOvJkQgt/gjHdL/+GS
1hMxPCBEjKkfhBbq3xYA+Bx9kOvtQwjeUb1ct+UE4ub/f52YuYGydo3Plv0uVuVVB9LmyseCwuRp
9bGER4qMFKFUikBRreksoV8NPotHy0MyyEp4ZY0K3viEsgiVN39yAMZlstDFwWlLgUVhol2dU+CD
T0CMVQlyyvd3vyG0oDFsyjZu3aNh7Dq3yex7dRaG75S1jpAikrqOwqSdkY+NEw9G9U16fdONm94T
aGivZr1gBsmEQNUlxRrbh0uGL5tFlbM1e2PyDd/yERqmWtRv3IE0RJA8jlE9BC9yGWh0bZHZ/mRm
ygqhFJ/yl2IAWLbHcIul1KytW0C0xejx5GxzxYvQ9xqN4iQA58GZIjGg/xnBNJgVQ2xxd4sf92JO
DaOwlxPGTRFz7IRIZS0n7/5nnUoBEKu5LzZ0e54hdXENbphMC3/8DvtNEaLbGi3CdavJw1/oHkmZ
7l8QVpW7jRQfMufISYZ3GWQWea8yTHlSR5gxhMUrq7nSbq22KX5SGkHXamQ7ki0RDzHlp8i04Wi/
xjwxTe3hWuMPDIQK1HhU9S9/+NVC/siyWsmx6h6nzBqyrpIyMoeXssE4NmBwjEMBNFXbGahbdoXV
SX3ggstVXgcT7egshEU3OmR0h7LkGHjuLK8Er3MRHtO1zQfx1iwEUYNOwtTeORsVefv379D7Y4YE
eec428kAQIeiUV9glRjgVDJJqEkoX465i9XNMBU4Ko2/WvtJTuYzZDVT11lOokwU+W2/cIaAkWhH
fKw7ZmT4WMnV4ObE/zyQ7jMRSXLVyZe6D2jEnnZgkFRtKZzOKdeyhEFvRqeQpP2bO2+EO0APOnqD
/wi9x0F4XafmCF5DNWbji5HdzHin78TH0wVZFVxHE6+yRqapaHQT6uQEX6CSwp6xrK99Km64wfYh
vRPYpi6HGDy5w3OzdujX2+ypl6cB2Ek5sXHxZ/w3Jp+aaG3Y5l6hdDxmHM3GLSjlzZUBijE7yW7x
8aaCzD6kEAueoeGKeO/QzUNzLGboApx+VjlmjygjoHByMkhYGhiumFBoScEtC/iFhXTblDTjfrUR
L6YNNMUIbgU/0dygh+Ob9kQ7JRjOqfgl0N/ItarJF9bxqsZAca7kBtFtrZ6dEddCuQ59GKv5qECH
MO3CVPTNdpVj7MGm/8f1ZjD5VnpoCYVNkIyxComhfX21/uDLjX+nM3MM1HceQOgWAc5igSL7lJ6r
AfE4n49sFA7ESWO+1ZhXPr7X9O4Ke1xlEVN3m4rYs/IAU4bTmdBUbca+UeIV7uGIaLCrLogTv3IZ
322DnmqWbuccvTfRwhg9zfv9R1rqmkLmY2KCLDQaeqMPtNKomT3SPo5hYTUnSeq5q/MYNAi9iGDk
CMzDAyOyi58wPfDQO1tX6+an/f36+OUb/S4f2/ydly0JSKQeEdQCJc9ynmq5EShUtwDhWwIEh52M
pB9TtLHAY9E49gpcYgvf4uBAHEngKhh+qSCruwwt2tZgYkIBWmlyvOWLnog2fjZp2vR161OeCcnx
InqR8RzpcWOAs2sf2V1HXxmB2IELLIy1msteU7iyppsDjayBHeN82HPAUpb20Sh0BUnZzi8/gUpq
VUICJLyhj+8SpeXzvBOJDPbgLLV08p3ZPOZMzurbHdLq6JrBc4F4UWRvFUkF9wj9eOUB3tq5LAHC
JCxUSUshpdgFcREcnrTbcXRZ4QwOFfjXPD6p8pXgT4K80bIMd584BsqJaWFNUh4SY5ivT1MjaMJv
Jnj/Dr19/12U/MDTrn8JSbdPRkIMCe7SLjbu1XD/ns0/zA74JXDCR41lN31+dCrHGzPByng20Sts
sZQkxgcU+fAiB4+QxhPB6OfZvCLykrZFwhCCOUt8TamLFBajpkbYDpYcGVHEcpKXxUY6Bn6gn+U2
Z0c6V38Y3rxEWLRQYO1Hj/HP+dg9O83L9LlwiDdIq5QDMO4gqJtpp5XQm9du4JCyRe/NiYlxP7jZ
AEGkd9o0LG6xAhh6VxE7ZAb6p9IX75elwhQUdqyDfhzo3+nFApvGzs/N/9KngjgmCOiaN2voB8O0
mqlBdwVdVaKtp2Ei3LAMm9HCnOqrKV4XsG0f0UlyCTjHRGpjld7SS3++xGmLiEHQCVWJUwx8pRKF
pvWZgKE0kh3CbtZ5BoCbEpxqz2ZFMWPJ0Pe1RtLNyHEsHChRTfMfba7uqCa0AVhc9z42YK2TwkOj
hIIpGWk97IC0dGmPE8rPLp1v6tBhUNaWmM5pgZ5eb1eKpVCWnroQFtxMiOqAma8Oqe1jnFDcwRXb
0BWeVsy5WD3QGJiHwLa5vktYcD6HWYmP8gF8CvmUUiwy0IPuclCGrnXSNOCnnQz60W9Y+waNQiNn
RqPCgLeLFjxuASDNgAw3wipvz47t6PmJlZ2N2awQgtwnO8ukRbl0UXIVGr3PStlyGBHbvJdC71S2
rC/nQfV2ZJBAemqCOta++gDI25Fuf1orX+hpagS/+lugjvRY5qpFCa5FfM6Fgsp5Qrul7SVYe+iT
x1xfDOzm+p+MXLx9isSJ4552AFXJwd4xaGrHdIgFkjSOyYWmcr6X/amS2MTX9FBcv6C3tnnrV0C4
GFK3e0Trnuy/MR9zTU9ElO6TOs1PO4ztnu1r2u11LIhE4swQB0oUmpQCIxsGN5FEWVvU7DPLLYhJ
xM1b2bETXe/Itrcbf42CX4nRQKDRhBCSUxZZYRY5FqDwqlRuVkd5vUUwPlJdHh2SlQFm9CeIqIT/
3VPxyc+rEYT9wXVQZznPp/1D8ccE5yKa40se1njlfbXpk+rAOPBz5fRyoWWLgiPRSXlaHfIO0FzQ
NuzsIhgfEhCDlpDWdgkmOihZNkAyFUVCCNc8pD/YMu14/SXLw8DgCnApbkeEH3mq+J52JIdILHXj
O2OeGWHoB7tp6gYXustSa2Kvu0IGlsSpLl/xmOC+gBRZWVayToVLMjI5kAOORnTkn5OHqUuotbfy
lEsvYp/ccCPmuwbPZF3B59ywJ7VOPqf531noI9MY+20POLUBXitfDYFOymkbHTeIxebigEv9uTyN
bLhQtcBLBObnhCkb28EnCp3oLtBkr/3qxchY7Y4OTO20yNbpSfzn8OLyVc2zxQKe6S4w4nni2QCv
DjuTeNLbHMOh/cDtBXxxKFqHpTWb47I+kz+F8nzxbtMYvK6k+iVESi0RPscen7egxjtSRrZa/ZHu
AY9D6cJ0DH5EkOm8beJSxJi5aQv2wWoh3vLswdHK4mhXDktKPYk1FbbINd3GmgDNzzQSivtLTfZL
MOyPkr8zkFKsPjdAJF5cD2ZIUk67Xhe9Idq8lN+xzsSFwl7fMeCOq2SrOk0adeXFuH4Dm0Vt4yWS
2DAZrUxPWclN44Dxqupce/A2uA4Gune+0BlsD1z7ldt8K+HGQplzT6eO18RJ3IToomT79hkcT8YX
rAv7IQxeaTKpVM4bSLl1V1dFIArw466+OkWjyrHlF4yx0wkIWdYiJYTMJy1IVqjgLKaV+7CFqhQw
foGTBe1hAojaSYT//MfdHUMXuXQFYDeqXso2JU6eI+dQaaQxjWTkNJATd1UXUVpyXjyWeu8TEGSD
i9Y2fo/dNSbnRHI34a5NYoby070tFB8tvZVNanvz1d+At4jHs8Iv5qvPG9ntNNhaNtax6Kq/I0Wg
Y+s/nUIKjJYM2QwC85V1beWZ3cwxiYqYz0oeFxC5vtXl8og/X4GQzD0EhwRQumLS65mJ5ngRKqyM
ZYkMH4imy6uJzy4hSTjuaHqbaDtW7JwNlOqw7jhavuLKIcW0z8yyfgtcS/v/71yBR5fd9h3sSPOr
LQohgl/ivsYZiZGWI75YAeHuyTm1KL/I9slDA83hggvFp5GVESU3CuR/DAYkD8uNF1hVGIVcHbDb
06b5vOWRG/4mUnIkG9CIzIm+K8obNPkZtJMdj8hfahMFHDZIeutXN3U+tKhtOkThWkmvZD9cpwhx
+epWMJdg0zrGjf6fzbDhCBY9u+a9GrRGSjkz1HkJGelDtALZvrsTlK6OT5jA6q0qLpC5DxYDgadU
Dyg3wXyTdVZMj4c2+Gt1U0Fh+OBdr/ZJyznFVaNL28YPjyGYBnu4ZB9Ti+Hvg9dpD0yBcHnBPdNF
bxTeHBI76i1jDtdsoerrp+L1FbvUc9GepJHYxMnutNc60pfwCIeeprr4MMUeTpfVTENPm/QWhBsb
24wSR0Z/qZ4+WL5la+nfr5oVrXEbKu5yqBtAxKz2y3aDz/f+T5FP6tSPfekm7yJRM5rbTDe+IlZq
3Hj1NvfXN1Y7QE8rCXb0h2uM5nDmwvP51Vpt/aIMCw9whqnI6hdIkjU7+hcRKD5l4cKSdFBT1UcI
CukUaQZ6b+kg2fa+nYAFXkjTaU/lirQLQsmbHZ9toBm8/nyf6cxynyCxSEcD4SowIYLWhbbd3YF0
V/vxjaWaR1d1FoLLGAtenpcae6dohCwaooWYeMU6cITbAu1UYMXdBVNRdS5t4Cv7xuDsJe3uOxlV
Z4EoCP9O7k5jYShPTbWwLgW/zTAW+180uDNYik1ug3SDG3/1TWhAWFSxGbAK85v3YZi14rswSb0F
4r4gzdNMTGA+Xr9A7uo/p7uG29fo3sTT9bun+sEx5uoH4p6MHU7p/y7tT2qGZQQyssBF1JGXqqq7
PwbTz6MAM6PX9/fc5tmJiIeauAr59uoX2T1HF1j9IZuJDSAnLk7gp9CwebXWD6Ol/ebPckMkvk9V
MrRXjWBvVU58Eix0U+I2Llom+1vzSZwrUpKnpkto5KnxI56wgphM9xCfXKtTdg/hUQc9AzTLjVUS
IlqxDx6FS8JJxSjZ3sZyQP3akMLb6yJbxmPl+Ac6qv+hnOIqZWSrdZIeUnvVgqbeiU5HxhsYiYzG
gDLbKLe9QzPdtTneDVGmlhaxjzWYY5RunUmVaYNkwvrtCjbIMTUNO/5TZp5Gego2DldS/GrAPjMJ
gA0NBubs1fKrJtoagMUms3fGHNs9XzhqaHFRFyLIE1aZn8qj3gAopvRHxcplNFVghZDIPj8J/j4c
ygGkjysOWAj3+dEEYOC7xCeHa2LU2Lg8pIrzh4nOq9R3PZLpyzxfL2bCYQbeT0Ouae1VH7IwlKxU
b5uzT+/0H890725ADY8fyNhlpfrNZYRXoQpjZ7bHCYz22116eNSlRmWnbiLuMAlzcMMtKNSoYHpg
vX0XIjjfbrEFBxfP8oq592Oq1IJQvtvJcFDxuGUoCNohZZfblp48seX6BfOQ407QeSmTBOh5KNCW
6RQizWe2CpQf50xrECU2tTQJq4Jl9WsJOi49/3F8JD/Mq2QIEqO34JQQQJAc13pJZo/UwZ8s5wX+
hs/HpTAML0H7Xqy8cL0/sS2UJjpUnH4Rp+1ZuS6tuXQduy7WEaWeSkEub3JmJB3UokdbHIRUQlhB
Z4Pz/KuXbEV53i7buGLNGEVNPDtoeYG9104TawPLTf4teNwclWgp2G7tOZSwy+6nXikpsKQEMCyT
49KX55xFJvBr8zDUyhdgVi8VURBzFw1DSsQylIOQoUdnSwhsNzyla9T4UWqS+gdiBXCWCsCLJWm7
Hgf48yUI4OB2o62Y9W+Z3Xr85cWxlyZLswULv5GBVu7+/kc19laUXPcH/EdrK2egfWcOPtm9y6BJ
nFgQQ9jdRnk5bnwIW8k5RhkrjRTk50zH2e6ZeKFMEHcacOLJz/juXxEliESeLX81cHqnTogrES94
NSaZNNydZIKZ9pf8CbBtNbs5oBzQhqyYgK/XiLf2INAAceAdeQeXyR35OeN0cLqyd3XZ1lFhyvvu
vfZfO0NsX2V5CHQhu9ONlZcLQL7pnNdbCkYg+GeKH8IpkEUW9aXoSpu8U++MzowruqMYJyXeb6dF
OkgK+CaZIbd2AHzlCRjeFbhbB2BbJRKVc6sK1OWoQfo8dsbXumntTz9CBNFD/qV6kPAlvSN+F8dQ
4Gb1AVy7EtGVmToD466YBlwzj0/pvuDeinosH80iYcx9Nd5NF/4BCn86EJ5CjBH4TInfudgtgzNt
99l1SM8lBkg/hLrn5guhZylGpgmCMt1tjw0mTO1FilXqwyf6UODjW5T1lePdP8qzUemYHWulEJbH
cWsc0pnptqKAwVpQx3/S8Q7/uUklZHyKj+l+VPZpeKi1BPZpvfODlf2vqOPAarwMRpa1e4G36xPY
OU0DSIzYZB8OD8UJGqNSXpDZx2H159i3CPYvYtQEhr2IpkZxtnsqQp9nixU+w2X11os1UyjHb1qc
3w14606J4x+QC7Oxm63gY7krmngVzBN9zkyNd6LPqIVdhcVLuZPZUvuID/n3t7Iftj+L/DTbvvE9
/CppNadNjangVLan2nlOuMxa7nN05bkAtf/KTmCUnbHVL1AkTgCzrz07Y5tWgrbsVlPnqXN85Vnt
ofSXz4plqBfijntzxznSs8itFmbsn2qHwtBklpmIMxivvgq11AB7cFuK0kkRho9XptthhB8Y58DV
SeQOqrQs9q084zUz+hHv25LJJ4dRB/ckUfKtMPaF/Ll2CNFsdyq1/Uz3RdmfmDGlqnUbhPEFnOnb
NrU49BUCnX8qXExaF3EZLyf+beH8OnkLtqjwssJzR3VO71UJyNUYd1oMB05fx1nPnnikLfCb8OFL
JoHX5yR8HxS92b5hq0LCt8pOWAH5kUY2TcgYjuZMCNENWNJ2KfH8iEjXIZs+wc/zIioklL2YBvuY
yJd2MPp0LCbWOl/ybgtgweplSbvo8KCiDu+W9aDZzrNwmSBR9UE9Q1FL5NBQ/7IMWB7g+nT4jFrr
NsaK9PNNcPanSQpMzzxfHNdgsPGcAEic9EXlHH+2m9Y/7qVcSnPgS6xhZeKyZHyrb7wdi6iV25yD
IkGj8LlUWfDga3T5159BjOtmzcxxI3RQw6pONAeolNCI8RtJ5C/Kc6MXgVOpEA8lpjho3b60Zd/e
L5N2ihasSY62K1Sp6Qew2wfA3t7k68Xa6uomTiMI8/zzAtm/DrxgRRwYDti1nFOJQbDImct8f2YA
XXOxThZHw7s+5sDGgVKByu8S1yHiaLEIuUf+2nIYphPKN5ZUwPG9hw1FNmt45QAr26ehKMhxKbir
wvriDXsoPu9rIVDlvu5gocl2bT3GAYJdtZREa+URu/s86lScEtgZpGPTmflfS0malabnwzGc1SYL
hJghR0S5ij0G1fDzEmg+0aorUPih04JO8yoPgOR58o10HAJOx00/KurDGcCNGh4HDErv8ge2IfWO
QbGS7jHkRUCHjSr4dxQpsGo/PTYXggWKhLMU7WpLZdIwvepXAQQoiuLtW8Q09wKZfdAvwt4caosp
4OFDgLMYlrf8tFSsp7Nh6xqwMNsCRJjrpTacybBJHh30KQ5IGe8uOM1ksyvIpCwhfH4zozaZNfgo
HlnALDhd5c/J4t9Rvtk1X0uyAVxZtQCS9KLOHx6oFHEQIQE0g9u8Sp49nlKA7q/sgUE9hj4OuK8g
3IotmcbSXgiNfsX/t50BlIul/0mtHKAoFIfDKR1Pty6Q6QseRetUoQ3gp2zM7gv9pNU3ltFs4PtM
WY7BBH5sR9G7iqO0lUR8DKHdOl/0XeDu0f+KtCEyOaeS8Hw318ivQTc5n8cOnbaFRc79kfePOYWj
k4drJKygIVbT7EbrfAllzuF3d1Nefn1GEsMb8CXlRs/lEbZ5azjG5QXRfGswSkONR5XFxzKSHNUb
w42PAdPFIv2l4f66UtV8SOManh2W+en0o1gqGBXrkpTuxviUsgCAXHH8cNKjczEBl1QPU6fKz2Zd
xs1hGdRC0fwuaaL6wYvVlH42TGLQCrFumWtM9x4dYMF+FHj1SoBE1vk7kQDUrazKQpp+ej+dyV1W
i2BNz7t5i9kSIn2hJjpxx2320/LXqKkx+TtszJE6L0inTo72Qui8mxVeRzZiE+ImcqvTd7Pk9u1K
eGeFX+7dDP7cNEz95GSTDYL2Vz5qr884WNHI25j1aH3JeHyR8QF6IvSQtXXEOhsFd6y3fhosWDq+
Cu9O1FTanqAyCIfJ8ngdMMk9+zyNwhjwKKk+Z1i7/OeZwBOeHs5hTylj5qAcVRZJTPVUWGalc0we
OBzxnnQyWV42JGFisaM+TlUE6pag1hFQpoGuKy5tNM4UPxjkByPrGQX6LIsgUqwhSTrQBws2538d
J7tW8WfsKLD8kiRZ+grjCburRisubjIAcoWFzBR4H1lfgbFvGeRjxZ8NhazKBqU+uu1mwX4b4Gq6
UCDtYONv/nDATXOZuOHiL4CqhATAsrT4TwZop41jj7UahJtkNUYyPByCcD3fIP5eOglO2n+Fywju
MDjWOi0mqr6kCdGFxLr6ATCY/jvkMQI8LfCVJS4kGbOWzFcvbTbqnxOV9OjVHowa68CeA6l6P7c2
8QUqbu8H/Rzv0TBrsO+MGdFn1r7Lmf76vu9fCf6cEXit58NVPNZwScq4OrWe2MkOi0DhXqOLWQ9G
qp7BycVGCoJQFOyipf5jqIFvYPKps7RoDAgTR7Yz5KkKmhxLiJ35uRNLnVSwjZWTYLhNLE+Yzn+7
1bIiOKyOXzwQRCjakXIQQ9yksl45FMvVYpT0Mm6rEtjPg4PAOzBTw6qtXT9I0KEPFQ9SDL4yDzag
VPOPRDB3xJGToSPp17ZMmBUUSwNRvvFmRlkT6T4eYzvN/BlK+EN3MKIUaisYEMvwot/FcMcToSay
99HxUWeyotg4wuCCy2SPLBOlOk+IYnIXLNcrNLuIHzJsUFqRz+ArdcfaxoO4n/jj9fWasJpWG1zG
4L3vQ/dWwtDi0pDcIa1YQJ5Fje0hICYcMV48MjPJCzF13VPkNdRbLADFyKaJqL/+qh8I3TM9Qk3m
0CSqwE8OKsSQunZZxE+XhoWWzqeBqOjZqZj68fXi0XFtl2xBQsF81Jg/xyKktgXwDer8fHcSfqu6
QCsaIG6Kc7IroXI7uIQEegnAS/R4OMROyG6nRnHmDZNVxC5XSh5qzMTy63Cu+n7Y91LRm7lHLrA+
KJp+c4gnWxLcPz23uSG5WVL2zE6R57y9ONR+8UfPuebP2m++l0N6LZvxzmC27mtxHlvxQ/8tEN56
DBEZbycW0akey/feGuhhG93ZRP8v0lqexpY9rgLVivJBR1bMoc7OtT84/qUAS1oeay/+y4M5OnsK
OmKkywPVNPREBuvzH6WwYW5jFazRWo24T5CVUcCnRB1bQ2Qasl8v+ZHRnBYDPKfbsFZOe55YQhvU
ELnbcgNW2d8Y/w1Nhw4blXtJupxB0E0Kf5isJWetO8hOjCvzpEOiNgYXTCMnDR2H8ingBwLcbabT
uEu6Jq5Cf464naJl8X+ERmWB3eA8TwmzzKe7rOK480VieffxqQuLltw8iI9Itzz7Q5F1E7fC/e+J
attgBB8SDcBv5zmGHjmSe8/u6OWSZomiYidvzmPMYO5SLudp7LzRQeFF2zsffE8t/HGuzGhY83gb
HVnga9exm4J1nsIaCOf6wH4L9KaT1rDR9p9Z3i9YlFHSHs+m/rUXtw7cgd9ZaZuVoMqBFLznwg4U
gtwjLP/3BLCFmmLU/dmBySRRyDfZaVzBUDSKn7lhf1wZWvHWROlzMU+WMKvO0KXXPTq81dvTiyAN
q222Wn0caxhqnpNhGLkBDj8LkAmaGVrkmSTWMqDy604Rj91xzIwv614h4/tnVE75JQF8z0L4xUea
XiK7O0HqZx11rFewzpUb6jN1j0MfvDh0TDjgcfRFHUB31rQSoh+TVICbEUq0oRqZeuslmRRcw5G2
yYWg1XiNYkpfcUGQeoBotNdg6bOlPoGXan1GBwpDMGk/VEXIESoLvq8kNzc2CCUFLhOXWUgJcxNN
2XgYBp4qf2UyA6VV+LAv6pUjuEIbCo82WzbzS9cFhGRopeKeHuxkp99YB07eM0nwx/8Lv0NFVLfX
QTQulilDL7oe0EtZeb9EDXh6BsLALkskUnICB0nwCbjgFrj4s4EMtD8r9c+MSHk5HB0a5HM3TZ45
GBl73utldBh2CEGTrfPbieJUkpX90NsgyW6DqRyvJmEVTgUvRcNlVbAABGDgm8CadYsU/rs4OltM
PeOnexYib/2H7OapyKW8pqnS329ZZWc9o+i8WAqOxw85ka99Yk0yu7PxQnEWKRS1UxTEf2o44PgM
VraN2XnKsrzJNWZBwozSKhG8hYAWsEouimqHEZYze8irKMkWe8Sy4uNpTplCuoNBp4oFb3PtMbFw
SccK9tBmEXGmkhFWh/iDF8vavm+tTdyDxJStEJzV432dKt/StO5oquFpGfAoKLW4GPKgFC4MSyGz
PGgbK/53lQFF+LvbiAce3MJLS8PgNtzDa1aYsmtD8aOj9VkqUl+QFr/O5XW4HJOfXXLijcDziIR5
EXBucILd28HEDU2jcOvuDG9I5CM1fg8749OvIOO8/Vdb0NwttT8+3WJMRQkccsmN1nxhfbF9daqv
5U4/kuOPWtx1yp1Fz7JGjJj7jRq9obH2qhjSr+y53PXlbqPUvsu7N8FR7XEFjKZ/cGGlJmHNdWJu
XHIhZAe6a5k8uCc400vmzd6mMLGDu2aQ0wbcscjLk+dePTdcwUr9gJYNADzgr9mCnYmEGnmIM8iY
9Bekkp42W50h5ey4ne6BvNtkyl/LEWthYrCMNtRMR0s3vNgCQsnFyk9fgGrMZTMra3t0D4V25pP2
RORiFJM45DVP6LSmwD/J/7POK7OAPzN1empBQ+dyUUDWk1TwoYXrzmd9d/h7y7sDviSo8AeBqJkA
nRt5QSJGM4BsHwAi7fTc/uuC2euGGD19/pJLWwdINfA8DzY0luoqovYCtDzNcLGuBq52u43kfgVD
ilVmy5qsV9gXzsTPIQhQ/yYU6v/ExhloNR4FrJxBI5XMoXefDz53BY0FiTDTJ/p+YoHCZC3myK+o
GiWoRkbOvRkhT2jcDJgWJvCUu3s5CUKlZRTrP5a5IGZZNgMtzXK+tmJjqS/o9Gu7Cf9muQqEm4O2
jQXDF1l548aWCS3JVbPvPB3JnS8+R/m4X5P27xbYN1fY+DLefSlBBKqcgfQxkOAjXFSxmMgfsU9E
jqEzBrWbnSNXd2SrRH0GANQDL8Rah3whUZZr4R0TsB77mpN2xP8/qpo0KCHjopa0A6Eaxjd0jwth
2z+3wQFXJUt2AY+P5bg9m67A/1FvYXq0P0FFczl8Y0PLkofr6lcJIujzKSR/zi0Y7ZAcX0yC13d2
jTBQAWFDx/0ceZ5W1AUDfz9Kts3P9aECFsGqSg5pgMHBWM0X44A71rGOE24eSzClP8fGsWhMiCCC
mPNsz0wJNvMEW/vqO/aezGL3/gWQMN9H3jRmm5sX7SRzEkxIQqx5i8FFlYoR9cEpTGN4l5bUtfFQ
MGQQPOmIgW8lEeqnPy1Jn/WCNavcSShleS8y58RKiJEd4z/1/Nb/NEvHwVCKzoG76JGPqdMIsB3K
tnxyfe4EmFOGaLVratsWfVJqU7lUICKfH+G46KNKMbsao+uqqhTArMyLmn2Z0kLZPn7XqhEA2r5m
FN36Ucp49JQSsk9gFJu7Ax0YARrzCRlN4A/SEGFlleKgGir+mc2vaIfkl1bngPO37n3lm8FmNIMl
QYpa35mhVPkiFmEFbZnw/cqmnzxemEdg3o3bS+eq10F0lPgCjowZLQU97OtE2YOkXyx70GmJJlPH
7LuvkbciAMhxro9TB6uNcmnQkmfm538xu/cTgnAfXbywfq73UJcyWpX6VmwZkQ9YiyIU/rbuFunx
HNeMCfrVtdFodIIfcMGTfVhv2PCCvFwtRoQWBUP1lzrthiGhDWlkVvm8RSIgY+UgswQvQl+mZow2
gsCIlrt9bPfO1MbPx8spBFoNSlA2LlHvKYTv7Jjk/zBgvlXCS2StuQgf/6z5wQooWxLtoHyaxXvp
YHoTRolI4k54RB59aVcoZ78u7FU+0me/skNpDOz1X5OKJGacRX/NUBrcQjoqQC/I3uzWq5zt3Eip
Qpkpz/0gGELjblu65m/8yrwrTGZk/TVdJZDlgJ71Rn9ie33RiUWyrktHoL1Zckim9WTG9Xnmy7VS
XfT4by6qGTZk9PJp0R2xROBVqOahVgpL5uhrqEtV/ZtPFWkl1j2JiPxt02+D9WawL919UiUBNGPd
jZBVF4LXlS5PIaffeZVbmnHtMbz8mpnAKZC/lWUOezoe6uy3fOXpYWPJtlepi9Oy0o554dKeStq3
jvw46yidVv+2fDj0MiiVW+XS1V7048c7msYNXhCR/OSenFtiJWV5KMXrQFVF/1PLfCC/n+WZypY4
debUoQCpH0ACA0jursjGHgJi9By6vy2UZv/ix3GSkLzXCcZ8nz3vQzy2+eMCpD5JqGPBNrZzH/Yu
aGO+lQGDvrKWZsyLzoEJPQjlSQo2BZMDlLA+rapsfHGceYSSlKYI5+9sLwZTF9I8ncaCgZhNlypk
ETVVPEzSavhnwqfohD3318wjzFjq9QWH4yG5GWlBf7kaRmd5gP2susKUO5GKATgEYwkmA6OPeoR/
ky1mGdBswexpmYlSS7NgP/J2wEZrlgRhHXqm7ZeZmAZhYhMh+QQODxnprk/uvXky9GsQgNW0EGa6
I+GsJQnfqvYpaNXTDPELMXy2agFt8xIKLr8oHHXml0a1lge7ZVGipwkNnziR84m3P+DjfOwheK7O
bshqiEIOtHzFUv70TRyFuWxioEB7We67/NGWptlUsQI8/Ya1EHzRtUaxyEw5RH3eIp8JcrUrd9tz
qSQJN/rUXEecECA6lVYJNq/wmrVWYyBmCUL/ME7N9JssFkReaGYGiVns5LChHwfqzjkI1kEoGKkn
pbynVYEAuDpjk7LuE12lNhwt/wSN3ARsq5J+qoM8ql/vPditXOCG+zHH7W4JthKaEfVHBhaTeMUp
HsY4LkphSP/g3KQ3bOJ9IDD/OUxVJxVExj2p2d4DgZnLAYb03oaE6JDjdFaBo9MB1+IMNEYTwtIa
jN/w+8HdMkjqZvrLG4O6+2TWzqsnmMhl0vo0dvHyOlOuLZVdfTF46SD8FvqTwHpqMleHt8QcC6zC
XVt9N875HASqz5nx2YlongvNkEaQNPPsbxgidXhwk5efl+rYQgjolTodUXSYYuo1/XhY3FVZLqQJ
DFq0F6s7dzxOC1zpNNEDFnnlVah+9J4ZES367MidwomMkDyKU3pJq1+TbQEV5o9sGkj3yqA6auMY
XlDUkzGdB/JzD43KWa4SpEuZ3MPCnyuIo62JQsfTKdeumCoM/vAJuqSAEwd/8vchAhxHXDoZZiyE
hsWJcrb4lPGKNiU6JluT+2lARU0td8eUAFFV25KLl5XOaKZQAUtsXJjlP36oHguMRA/mNW8Z9Dt3
OKzlUQArggQqgZzI0wFdyaoolAxow4HBasJVaPcXw8qoL5vyuQmuuGuWEjBopfAfzg1qWc9CNYji
yUlqxlZhdQM9ZZwO/HWtfmAnEWjo9TQQVN5KXB6tJ8QFmtZ515OOr+Jyz16MMmW4RIfhn++2JKZO
SM9dCjpO5Zn6nCWXGppvthNuVuJ1Ki/tlWQydYSqnMADh5JjitsE0r0TK+x2erjXa60PkYbhdww4
DOpyGRDGWwuOyjX1xG/pYuW49L4Wwl1qr635vGOMy4UTad38UUxMXqUTvTZrzjZYJDglvnzdWG2I
goFbD9g04HYGE7uBqfXorP02pdRQmHaN68llUYjBwKAGREmBvFmeN55cbZ4VdOTByDqdLzUI8km6
Um1PXg6181ytrrBdNtoaFRAijkTUlrV6anaptRUYXiQF+8oou8yxLTscMlhRcd7kmSyjgukedv6u
52Ls4FTmpqogbEBPLsR8WfR/EvMe7fCFH/yy11xt7GyNQB5ZJLBESXBHhrQiVFVINvNK7tvymFHf
4JiSdiYcADvMcrBNV6MWjrqtnQVe/K+TKPZOXWr3rWcCUlgJ2gyGkrC8o8VjhGac8jH7ERvpDPEM
2ognttctEX0RCqfbhUM+EsD4IhpM7YWCq/apw10mMWf0rdjAvFVqMzsEjYLDXSQqp+9NyLF9xGl0
FZmwQFT4/PdflxZD0jtbAgtKi2kWVf8TSValBrQdhA4Zva8N62ZcY7LQMuxMlGu3qE4eqduAtFav
80j/YBmSk6wcD27cLpk3Vfw2VxbT7hIUlvOTNZxSj7v8IO5/SAARdefxBuu349u+OfU98qiYj8jQ
Lu92Ik+WqUhyQEIujCxf7tfRln3u6F1924SrfqEDgX02eh/147YEgOAgmgrQHV5hcC4/HC1WZoRv
erGAAZIjMr5lnUmIk06fjpVzhhFV+ztamufO4v21yYEpDHp67cX3fKBiGl4MFe2k+6Tk3sqHDvuJ
PfcVvfmo12dHq0k0NcT3SiyNhNu9qpgfzWqoi/wIyToCUttrq4R3X33Zy2GxsEUYOWeUfioQvEto
MV0miiI3/x9A4OeDlEMBnvot6X9EII0jYLBZSGnENsWllAJkY2hlSmUPuRzYmdtZi7DPA4IPZbLX
zHZpShCPo39BFCCrFZzmU+M7pZhNxoA8j20w+MrThdWDUmJ8XF6Y02bFLeXs2La26VJ6SaVTzpmH
OFhihobZfLuPCz6CJ+SBU9esbUpdJoUIWV5h9AcQOa/36EIlH7E1M4L2nI3jUu13zjt5EYpTO9Vt
DKHK2lfW9TyQ3PE1RG5bFQ4nv6ChicUDq7cnVEJAlKyMBUjwyo/9fMQmMqYViyIBmTzrgY6E874L
ocpuk26XVMg/PSzIzJ1YOyBN0HnJ6XItGnLu8Z89d70by5/qWQWRE3aRmPfAvn7gy3PZL/clloDN
VOsC3l7FcUHxxCoMubQPPmpF5qTzquNxOq0uEVTZ6IgapystbtDWPiIsNRULLjf3VeoDCbWIeQBk
rdxXrMtu0uq1cncVeRZOhGwxqWMxUm9et55Kg+9bZfRIgK1WSYtpCtL8gu8Ofk09baHvjZgz2LTT
oFDWE2flf370XbgCXBP/u9Mw+mEg8b0iPyrjkyhM/MMyiLX+xwwq7y1tX275Bqx6U4Du0EwIY69X
nv9RsHtr7ez/l0i42KSPXBmJ8jGdo/gBQDnsBLGs/iSzG1Ie7OATijOK5WsjYw7PeVfxlgmESk1O
9x9bW7rO66+kCDayqPJvCA+1FM8Q/jgwIH1R8fD+dumLIEIwAYH/kjcQLNr92NrLzK8+PnAocuJB
x2et7Ic5/YZkMeP1v3advS5EuGM032H3+lehF+TIOSr3ExJMAUzfHQw+d/9L2r+q2lep8qjdMF78
XT8IKiXA78iDzkA15ZYqN2Ubnkk2GN75TH3mRbCbcdlIwM/eGpkSTyBaRjVE2n3kEm0PUUGvxguM
bEkjac1P+tlAhbTOeUc1iywOxVk9bstGyQayVhiNi4rVspeX8EMVjGFW9FJwlWH95dfKA0xWVEeY
Khe6gKTVYA7/ENJWOpYgfFqCEZPiPYoDzl/MNN+lJ/BKRlglqCpSGadc0efocaDBaspkzF8IxDBg
6pBKrFPRuUrfB9jWpu/LGWftpq5UweFH3CT7eghtQaWpXHPE9QTjx6WliNQsUExgFzmOlRz4eOeY
GbWI0Y6DyR/xzc3WZ8TCju1CpZvi3FvoZSnHC1YKYM6sQrbSyGMoYYY6ngM/CBN4cc1cmF+uZBM7
NMZY28hNrftGpecuO+1750T9R8hNvguYcZCF6F1YlWvol8pZvIaeW9lLx4gOLKCd4wnQM9E5FVPd
fWps48gfHSEAyD+SuRXppRquSeaOTV+1ImNY1n8Jla1uzSKaiz3XUb1/8IPLbeehc1Xx2y0TK6hx
AEs942eYuSF/W6YVL/ioACJ5Ovf777hL0yUywFf6g8eK/mQvtBS3ciZGdhgLOtAl0IWlqKz1Fkbm
khyK5uFaT2ga2Z7EEfu6qEAR2ND4xxnXJootvLcybpBmHd96lG4OKbk7CaXkBYRXYhk+7W2r+Avq
hmcW5IegaGbxr4352rkXDbN0df0G2GWFaXMSOkRCu70poK0SWpxjhkJsU/4sgOzZq1B3yadaPuJv
/VyOMx4UToMvVmmi1F1i/XfVWxEk/0cHT0fyr94cDRAGtjTETnsZVEWwKIxAHSNJ5srblYMUcmOA
ScbJ8wo6mdaMG8V4yslVlG4jyrcHOkTIuvi99hcOS8kE1itwdlcZLcTHH4QkbEYE4LK+rJEnfu9A
Q1PrcvK3Q7HGVFDjxQpq3dUJlZSUF+3yfJ/DvOlfWTjLrIfwlB/KgZggWypXCUlbtAzUbuI5+iYh
9Hz+6PVgGYF5cAO4+iUIszoPnN6pmxzak/ybg6nKxx8tKOtupvSdA5k3WZXDDq4BpTu0LXFL/cvq
7XNKbk90AHwF0mBOFWiR3nQp0TurUWxTnb2pNJ6MGf1nPr5alko8Dh1TLorSw4b0DA40/zXmn+Bx
UW56Ytww6MMXt3YRInJK3fOOylYQlivm8EEb1y/HozMq4KaOTRipcKU266YQUnzXLvZEnn+dMIiD
ozv0QogFIm180L9y7LtLYzwa6rhQ0loGiuxYUu2v1G7ofsvEUT9twJPVtU2pPQ7bSCINpt+mCAKF
VtncCZ/4lU1Tq1AsJRUMOurBYqHx3Kq0Fwdlu4nrwnBO2OLFxRHpx2d46sVENGy/bOgbT8e8wcAe
CL2caEpXntBpIfwIvajbqMDwGsdbu2XvXErAx8f/4DIdXWQ/uo+Tplf4bdge2kaG3I+YkVm+kSPs
9XknFmfS6wAaMv/Vr2bfwmT99eoAWcd0ed39IH45bTIMTNx00dKX/2bJH6E8GpT5K9aJeWYFD8y8
AVFLVbYhQdeFa3wzrgwP9+gzaoHQ+jTzReiDGBWwGMFdJgYkSEB3z/6G8qdbMxBaZWQbCiC1LWMc
zBBvs3ED8t4RA4c2L1I8aNlxhi/mLOgrysduEh3HsfelPFFOz9J66QVy6oJwCjaIxG7wUOGRit30
nlJSVbHlEpcVIIc9+GWSIULT+uSMv5oLP30jMc4Q80DnseNXnUXLmZefIZEuOf6kRASO8saBRg5f
PKhierrCJeX0AcZZcJ4GI57qZwEd47A+/vX+giXoEas/rDT9G8c5/PbTJ/IvLFQQzocsXJ/aLjjt
C3jWWxHCaLOzWs2y1z13ddw+vwnUpnolt+AtjTkQ9QJTs9rP3cCanKhQSk7m+wXF0hxkVLQ/nFVB
t/qsiF199MRbFOSvpNxWFhdVojURgz+2Mdu25nCW9oXT9Lw5NLIugnn1YI6KgX0h6RDOqltpi/XI
ct4CQNXU2RtXG1ghhFN5B64UUH2AYcwfjmcsBJBSm1AugFsBFE0BSIUfgscOWbaoiI3QJcRvGMfn
0DdwAYWwiRtKhdi5PzktQ6qitB3pHGW4iokA6uvQ+a/NqjP6isrb40hkrU0QBz6wAoK6AC9MKkaS
6S3boZiOSKuVpgvoGGE5xSzoHCgNmUhMbO550r8oJyWINKjpw4HPq8IlZnLgNrexspvZCiVYANzH
KSUC8M/EOEh++YRN/C/nc+6tJ0n/M0m+ZJXSLZTYVaIkvdbkBJt8CU57LlLpRq8L0n6LXArxAxh0
iHlLS0cwXifXef7KibC9eI9L6nmWErxwfbzJxo1/Kly4isb2GQudMIB7s65zdcokR+NPPftRP4pL
u9LQUsjcaWs7mtaKVGTjnbTZlp+fIIg1LFggZdsOyBBPGVezgW9vtJihK+RinCNBa5Y07kE8sKvL
wUtlegoOv0eOg7nsg84jm/FB2GN5V0BH20MyzlYUo9lC+6KQBI0Hu1kUzjfayPr/UAi6TbQ0LBop
hUTCXn5dW9exbJHojNPK5BvQBCCDlg3o5zYAxxaLgJYvcerjceYMmtqTyUDx3VKuxvgW+5U4/tuE
FSFkOjRK4WxGsx1jyzzD4wn2+ax8L9bfTJVkaVxYK89o08N0sNB0tUcNd0Eh//UEe8jwUjLYtir8
r4lFaIRCtePfuldo48bjJEnHtSjIafW9qLeciNYhzQd5btbtWPit6bGmRLWpN2sLNUXIJMY11vUA
KOMKW+BR1W1O6yigwVFbrv6BlqMv4rdVFDi8iToH110gAGwHG5NyXN7Rmo99uvSPsbvrpPM8bVvr
QLluaHC3Wqf6IDeKqmPaCOAdOjAG876+xp1/RV2OsL9hS4zcFl14x5fWJXaJIDeES3NmMHX3LqIM
xAgZjl2uJM8TVrWqiLGwNZ0CFzLzA1ppiOrFqR8cnfpzfG7QUpMnN6PBsWA+hMqXdzCo9IFG48xm
4HvE58d9K9ch9kuigmIN5NbkGBlHY27Pk9pAUCBiqLh+qLGv3egB4jLA0b6Y8kiX4bRdDw3O8FMW
/y1FljpdtPlKHRsnwfxoSfaSmzY6u9uCddegMnz1DG+AmOnMGPEnoApUaGzhqBAzzB//Jdj0EfSK
xuFVDarNqs/Dd9rRz8R8Uf0z9j/hz7nwBWl+0ftU5m0pqhNxB6sjJUxEsxI8tlFMMg44NKcjLdZd
DLA/BwqNdGDc8qu2emdyRl/QhvSm3q7WRmI7cRaW4iVzxTyMRQ7uCzcvou5jNnGbcJdaNqri/LkM
bApzvXlFH1hWGYqC2Qgse2EmsjM0jJqT8Z90Fj35gzfEbqN+UXI1cqqK9NlVKXcK9g1T+O9v2fEw
WihHjsYo4EIHKIJibvtyKx/zc6NifGcA/Kquxc1d7qXlW9pa6gB3R16tcAUG3Gc57ysW8kwzwt6f
fJ2pEDPmBwohKZKaeNgucNDm8WLziyWRiitgya/K3W5n6yBnCDsmOL9fItxnvpHu+iSbDNAI050e
ppmBwyC7K7xS3+vwkiZjOPf5k3WaJCMt50G7Bqcvq/TF9LUMyw3A5EVNMwJ2vJPhMOLiEKmVArUX
Mxd7mpmmq456oSRiBX+QYdcOwqoKnGburx6WOw5we9rYeaQ+djtSCYNn9jNxo4CIhRBSx5sccz71
5pF5X4LuX5M6CoQeOOzku+UmX2XTdCOzPmUyGvTgfAs13KCMjrs2FTGM/qitqyJmr0wjx/rfYHPF
tnfO7IrmDAsMWLDfvmH7hH0J3Mwl8ESvm6a6z7lyubEu0564YKkegtmNv6fI//ruA81p1e7KAvq9
vn+ykeBUEcC/qlWguA2osHDRK5f9czzokz2WHVh/dkn3TRpW9EMTZ41PIG8tXSHVWISKknnJCXfD
NJEaA+y961b+zUXsyC6wdnf71nTdAUgMy+Rdkx4WnmkwE3amzmWhOP17Z89sN233GgDr64cWAPQF
A30fvPsIQCUnt0ZC9vFcyv7oIdzzwhE2U4L2J1ebK0dHnGerDe/MfAbu4mNQpBOMuzkqkhYCyV2u
LiTxDCgDCSKGp1JouDeWJthNXzTZeO5Cv7jMMc9gU+mYrufVwxVWCFJ6N8UvxzRLWn+RD7wM88qt
Uz125Fc5no4E39SH2oNerW6XYhJ7d26bWMFan6rwtypP85SPbv5T5QXHymf9rwPUbcnDiVYUqfCS
Zj/aONv6v8A+soHFcVMNGVRKQN/KXea3U5FuaZRBSFUif3g0XEFd6nXNl/7jbd6XoUJwILgjxEWZ
G0tzeie/YYaj+ueOXTeDUDbE99/hZl+2O9yRInivMI+wer/eHOevER3mkhkFIMezDne6URoY2w1b
7tZOmEC9/QJ5yERN9hYYEiL/vvbHpPYubqb9Jknms9HHxgW4zzN0vqgUn3kZa26dSpoUlfIzRPTV
kLsYxtgvCQmjAcv+6qujNdoJE2jH4Xf1jH6RINLh8bo8peuyFISA3RTxOtDQt2s/4XsowderQ37d
aUTouFjHQ5gbOOoN8dcFFAD6oQDwxQz9IXnlM2bENUE0SheUtQZ20qaOtVup3VJTU+9KSLWAn+PD
qdgWxp3eJMZfqHrbMUiG+h7j+gORpgfhvhj3ASqLBHvqMaTkW3rum6M9fJw8+PsgBIcNb3aD6x7Z
7PLcL1Wl1XCJcdCxontvfgfUEmlB6MD0xvw76NYpJjtZNYe6ZINv+BnUO3xcurMmZg1TY2cGTpE4
mLE+hJiuVpBUHp1qZH91TOq0H7J5H089syBUcXabT0gcdqMqJTtf4bupIjfU+a6KL0NOzksgJs1K
YA1TBpR+Yp7X20jxZgSyo1M53TF0Yx0JlVNmunA6TK8GN3FUW2kxJRwsxNtpQOWsjLIm53IpW6vx
+kxga+z9go9i0QkKoB0JsToptppxH0b60QoFibla60Xl9JMXIS5YaFdWrH/QRvuIZJWq9wVedXH6
xtRxwAW43+YgsYN95bc+V8AEZZzfQEFc7yZOfH0RPYNNFmo1QDqHF5oO48Rvh8V30zlLFQ9ld9u6
MMFPkubf2FotVZIsnpLgT4IQW8WNZt+WS0do0JnJlVZffKiPZ/AGes6cyJdTL3tVMl5VzBPkJ9FY
zyoNocFCp5zSyRr6fDl1Lp4R6nicROaRLC77ab1kG3iDbC+UNSgNdysDlow+jyXrQyRZmQ0omdJJ
MOT1VVKbeT2AcOCL0Xnf3/7xDCknQb+E43eNVQuJpq9GTk+QHh8lfy3kT9TH9UGq/RpOmGSNQaR2
o5K1A0iy1B6cT6jfudI8lU6+NfkMuOwUtGzsVs/fB/aOY9QPOePDlrrz/ieKE6BJgAkEwWL5Maul
I2rot51MsidGgS1mfVrZCGWj/5VKXUo50whDb8BTGXNraJEbmyqM1XzTCNaI4X7GrCVhZ+z+li8o
lWBVO5kJ9LQTIWuOrwk7X8aRSoUWR5u+cMTPi61iO1oEIco3mhTEi6NfGtGpKRRKa8fGXx4oYy79
CgwZJAb0PQCtAhe7NAhe5lRc6THDJCYA3dgzjNQG5rtfGzQVMGvPg8S4h0owvTnowGhdubNU3AS3
7UYqLgxWWzT0eBykbnJnxEzml3hJvBvaHBi08F/Be0NolsJSrXEC5cCAHl4m46NdmMbCVYuXrJmU
9CJkUpra9x5EfJej0ciSiN+BNzuVXeEqX9Omelgz0pyRDBIzzTQkrYQzQ/ixfK4wg1OgB5rHXCjt
UGx6SNKE8Vg2+tZMiAJniQfDjuXikFGKrra+qTY7EaAIVTBQpwWhcg0NIQ0LZ/P66QIzvJxqkJ+A
XL9v23bWstXSyjg4nBA/rNnyDAWIUysUrXby/7A83hdNbGqzs6zILJkllTaWj4VVbmaSkcxyOcA/
bMCIdPqkS0hL5aCjwQiczxZYRiRX2HJDY7BctRy9Fo3/dg1dZ9TfYo+q3LiEjD/7P+if7U+raGB/
xk+Mo09aSgSVp+iZQeTLVTbM0WBwU9Jh1cOHI+ZgdcZFOULM4yib1NedDetMcSWsKe7qOJmny5CJ
YKrSJ/A2b0Bqxhz6Vw78ROdXO7dKt6q+nWnTK/0mWIObzvsVdOXuZw3owzudt9au39qpoS7g3CGX
iM2z6sG6khp6v3Bb4oYnsbkcLATv8jBreZNSpO7VHXdFCi9SbMsTUrL8lp6hUP2omh3Ydeu6x+LO
grEXPGChP0MYBJVKJo+1OB/PIH9eYFk1e5CdtxIrfFWBEFR7xBohSEX9WEMjpNuIIG3sFqeAkZBZ
mVUYArzmKfYpwYVbCmiqo9bWrRuHw6r8tt1hl/sXtk2nEm4/8sUF+osU9zHXYOaQD2dU9M6Y1+ra
nJlGtzvCkKLptjS4/oFz2cxQi2aeDh2xZ0JTTiDvrckxx+/GLlaTcnYpuvle/PaBjSp9NlSIN5uY
22c+JMBoANHrwJPEAxpVjOQpmPfsZHljFX7Ujk7mejdocPPorRJhVz/xbqpwZdlUGg4vyFrta+cr
kJFWFU5DUDAZJwsfQkpuE9KdSrYrdOsYmVTRP1tt9ES8cdbhVRBgTH3/y/VPC608hCuJH5x9xXsb
MSEyzTYsqiPO24HwAneiKJGpSHo/WShBEVIOQkoT+PJNXPLPmszj2n1bUQ8e0JtDjQvNEJCyiWAf
cVazvy2P0ggazYoJkFm8f4QFAFpbq2pw1tLCj/WDFS6Di8HaAM48QXvc9MqW7BH4qD/bknT5nNzO
Xwp87K11h159XL1CACXpIbrBMAVreGdrkLtuJ+GTW5W87LoD6C0WaFN3C2y1CfbxaYi2bu/P77aZ
o8nBOl4hOD4xiD8382rbeoZwPIT3RHdZo8lLItwU7Bl9nP57HM6nC2BaC0PjwAB8nb6jKdH5l/xe
25FK504Ks/nRPsiZ8Edud2+V+NZjU3YOJOE22nWEDuue6xNHm0+lqDdr7m5TZ8RyKq2411uIEmjx
+6643sEuMnptTR6riwuPUo6xnHgkw0R12NqB2HImF6PU8xkvWrglO5sxdEddIXWkgRPAuNugFS8d
g3vwDOs8ng7VpO4TPY+VfJ9seT2UJYx69i8JFLsLMs87pCJbC1G2Dg3vlM0YWNpOAqvOP6u5Mab+
tEW9UEixXwIlBzmCKsXRHg2driN2Xaa0FgeB5QmE8e3HCR5l3xC0tWjtomBJNvVqtIcD3yZ220+Z
WwApXQI5vqTTPPyvuyQ6ZhNBLsXzEcKk/NcIa4QAzCK9NnFSaHhUE2A8E1H38qWz9GHzXbVvRJCC
FaIaN7LjC8pPUYq5hS8F3HAW9RHtdkxFCoW0eKBdE21Mx1EyuA2cf1qFY3lah8E8Qxa/6W0zt+wD
jC28gBBupDkIdoti87D5zCMGAkRZ6IrbLgGzl2hJ6i2HjT5r2GSpFY2VIo4juuzztvmR17RMz7HX
OhYiSVKneceRkoH4c22YhJxYW1hufdbLc6QUkNcEyljxGytSqLcE/4ihu+bnuuGRr+ypFAJbRkOn
/oIQdYslD2AwRlL0zD0bQdKe+HWjIzM69c5rFf9jSJncQEKss1gFldKRDG/x4IUR3+hLiW8sexhW
fzWb14+kkfEeuyeNAuQbar/QWOBoREztftZFHML8/gROPorzSThg1Nj+VrFpypXzS0KSkHQxWpBm
fdXBmDAoL/voSqH3MhJ//k9pR/vPrhiiqWJLWn9mK4u1RntGz32LR2RR7OhQ1fd4dmfKUDyRv7Db
nFABZI1/hrk/FBbN3j1tpDn4mcvC5j5uZRaUN2TaMxuw9TevHrV9o5F/1vSBuL5BYp/E/3DJq/1j
ln+8PncdOMq5nSC+C9vC+tsf1/PEJzLkC6QO3rjSL28JUNkViPxMW5xNUBXOJN4pnqYrlHL5qohh
RenhG8K8PzKy1G4hrHbXbDeg7oD68/mctvho41iLrNuZEEzRfaIbxEpBBPwKRJ/Iedqga/YgDMrF
pKToDtINMwCL1m1bNlVGFqaagVapm/Z/KGsTyvL1w/Txf/MQvx0+YHlkV4ptlvrQbmO93xcNKoqV
SaN9Z9bC+kvX+thddlafqc+u1+Omvuuorf6uxjYRm866ZlgjGHi9CXBdBDzwr0ZRm/s6QI9xscmc
XQCx5OYWCnvOkeEx1ArPp1IaG215yAeb4+y1xiVnFf36yJ9etUviL2yknpw3rY56Fhn2Ni2CZfLC
Pi7pDrpkscWm3/oMDJAX7c+wIr1z/x1IebAtulfp+ihbkJ317cHzExlkmrPYC/VsCuPYe6rHqkjy
X9BiCgyahPD9SQWMjbvo//Si0CxBVZhGNCWi3Ou59zzDUL3THJdK01Izys4zKRP3sBpj8PKYb3ax
q8+3Nr4wRg9PF0QgNsCV9QFKTirJuR64ocxoyAwJKXShTNA3Iok2BbD69gOciBMK8TEuGARf//Bk
bkbdTM+B/+sniqOlQ1EmWJGnojwmeaEDvmzZHZMRcDLrscqBNrsXAvHDhutBjxGou7u723SL3Pgz
HP+LnCJ55XTH+HXgEV4DfDra0tlJJKzZ+iRg/m5wlSCbjahCFMBKynDM7vy73Cn4fKXxBgfGseGN
eRJW5UiI3DgT7qBlgHc0VqE4I7H/lPR0QEyox2AcuD8iQXI2ZrjfL9ps4aUe0eCqmddhgYT9gonM
5IqQk+GPUT8/X2RVYqtUTMbTDFYSq7R6q3LkOrcO8y+TfWxXjWcRO8LXpkB7UmZo/RxMp6pM/j0P
dK7QYCr1MVQcSqvGSdtsv1ZGhfWlN8+VN2/7LXsFiq82ozcBa/hk0IpIN3poAAHppnOLX0UyU+Na
FkQlQXOwYZ2ZUmipBQ35aJ1NkO8F/twM/udkL+Ii6nYiTpRr1rhlzvzerw2+iYAYWYW7VJwjepIE
yHXkecAK7fkHrmlAcpb/iEc9+qt7bPYM6ClPQzL830QBsxblDqj83g18bXMk2zF8a3rDSLGRNjnz
WI1HXePW540gY8Mk+NgS237TW09O5BqMhX6+ykEF5XjYs/Xj22OLwNsGIm4fNKuJxwjQP9SejBLq
7zMCQZ2UDyS6X2qK+MvVDqZx1dXSBVVmb5UFVTreRRCgcERrLOM8aA+hSSbYyAEa5H8dWBE7vlX+
sQFPyRQwpOaRREQhQ93I/1QOfedRTAn/vuyDmHeLYzAUdQlyTvFcU/+ULVpBapvHJCyxCIX6b8Cq
t97lIHrD4TFyVXIjdY4adjWGKPVkebeFO9YLpfvCJcJku22/lnhca6CMVDBSxx0F9GxmRmUPlPqC
BjPD88CfDiEAxffGHdupL+16z2xICrKtKfmUsBUXPGsy0dIa7SHOv6ZZZv9aVpoKARVo+7bzEGNa
9TxnEmaKYVPuYm/9raHJgVim8j1L0PENgYYtVKA6SrkYukjIrPF6ZvVI9OKgH7YLyJvTs2cvXW8c
kGhEZ7eqdpXqUoQ+J+PUDp15pIE6PVOcEoSWhcL9N9tOLtcpnti8xw0xgu5LnbWpUixvPRsHo+Ru
9qtbldArHbSQucY5Fj6Bbj9iuXYqlDJNqAQHNnvvzN+d08zmowwkjt5Z2nnmP6VDhutYITyVi30Z
cY9U7O59i8d9FbXkgMxTr50czlsEX6IwgH/i/BCZJfLb6my6Pqc+tg7lX1PCP9E/7iC/O31kZ9VK
629ttk+LIbSXLRyTJsoIsPAfFhd+lh7PvdH1m/LMSOgpf/JFgNEEbYhSewmqaOToqij3GS++Nk/H
AfDH5khGsYowxrx4Zl3jvdLpprrIY4ZGOjnRmI7CyNG5iS6yFC0VVo1C60gmRGUCO+Oy3f/3/dXG
pqZGTFmWugttvjkHANxeqyzMcF2ebq44mawETuuFthCGHF7V7ZeCA4QowyokJFJvFC4qM6kJVTp9
mu+X66ISdYaeTBijXdauNG4QUAtXmOfFvtspMA2+oGX01CC9zQN1qdfJVxZfEFqNJN19oYKMjIeq
UZo+GufIRRmfURk3hY9kdc2OiHovR6PCykn1WcVETbBp4NJWq3CHsBP5qfSleJYgf3yHR9v4z61C
QAYaMsqNaaq59HrbytSaFWv6HiBB6suJY/vhn4sg60PxbMq12INeCrKLosvwN4knFyFctq7qDkpE
AnwKflgyYTUOFKB+ClH8lpUiqvIgyvKBO5W5umvOiGaPOWCrIriJqJ8iT0ineu3h1V7cFRPXFpfa
BQoT17a9dKLlwNSmzs5boN0UHn91SpAzr7LpE/FSaPinLNvmcz80DbiDUmN/IAPdipzieNFYg89u
0BvwgENufRFnvifSB1SOfv7StGw6ome6T43tpDeY7uceNB9/fDepMyUFyq8p9sjT5Vw0uRN4++eo
vSJepEehXYqE9gNGLofpadJjRHVFBwpcMM+fsPZCA+97rec37IiH7WG08YFDOvw97EbUC6oVvSI1
r6wljGp/rMIP33u/Z3G5C3838I79QLXlKZh31zvF97V7j97sKxwYhkpsn7Olf0YPJdbCUJ1rgf0d
UiYsqxlofG3HweY3GfSo9GoYC9cJmm6PJ3f2dc+JYevVA7jC/vqT79QKR5TpBG05byLiKlKM4aej
K2qFeKmNRtmnyYsO5yngErE6ivjT6rY7q8C4iK3VgilJKo4D8d0HA0d2UMOL94LFhchy0PC/berJ
y5FZ67mFc1AuvUQcW+RVXVicNOW0+cwrM41RlmVH9QSUjHENR37dqximQJszeglhWDiQomB/QOlt
tIx3l3tbP9s8LCXZQYc60bLslf0whZEaAIoamFabYukVOULMLNIoYBiRA4kOu0IMYfD8dMZnqJ6D
lWWJhcfyy78HzDMLObAP2pq6VFfWaSgMbU9WjfgBQCS59haMluDivQqmrDPEwJECrTy0T+9z+MPU
DGunDeqzt1qYo5avA1QsND64r2Ii0bGFe+h318xY2yGXWHqczO6BNvm3GTfkTsrSmvJ139FL+fzQ
SATPW5IQ8yIQ7INz+0f5nJYnFlrtyzitEeq4f8fVQlmflF/5sPpap6IQspSPvNemlyHGh6MqVJIB
hAfhGXFGl/N+bgdTq6sFS5nSoUmTwHJpkOPI17IDqf/GXbZzcAAIFMDAO+H0NaPYIXlMFPAj5Pc1
LoIcz4ohAuxERol4/0Y690RdHS95Ba7L8SRXePKUAmz6sl5QpfAYuS/H4cmd6uMPMwfgSWnE7hBk
0ZUx+YflADtHST+cyX5JWS3TIvz+JNo7QGcppcHMeO0TYF5jefLmOoKRwuxEjwMXox9g6vm9PusV
3S58rLNPw3qtut3ULIeGg38emvL/IwPeTJDdRmXENInrQ7+4v8fBfG1D9LrwxxYzJ+1NgxllrhSx
OicuBcHLCbJ2IIzVi7imOE4+RnpuDcOFkRqhj2wNY4dmYjYMnLZHp4DLbw3YloQgOCl6tosTSF8j
HD3HerFRBbJEyWlmQfy5/K/Cb5AogW+lAHuU2UCZ/1NjqpivrqdPDCKENSECpGtluhU6/DVBbf9e
R5o5n4Bpt5oQN0X552zByxgXpg9GqeBGUTCIK3gGljshN1Yum2IrweUJNR4Ymzfw6BW7V3Ok5RHN
G7XBdSYAwkfsO/sArLIaDu7tSVJc2yU26/aa3J11KHCdpUFvbwWpqEDiIhtMH5qV4PyYc+D8ABZv
/62a42PKtuEHQMWgR+eT6seGhJ54t22rmT7ILUB8bYpN21zmaagE9djmIYhmCK4PddLSWQMopFWZ
bIqOYDCMzSWSowQghLWuWzT8OA6UM08YWxRpoBcgP3bnRvzPevAG6edSeMzAufvSmVBPhzzND+R5
6ULrmlylsuqwiCS749YSys9857+XXZc5+zVpCMhx5IyDcyKJZutKKUX9yrWTl5oc1NX7UCzOCHGp
NBJQVBKm4IPz/rxtTOdSc9Yw2oWdHLtR/JieSXatAh+uPOQz4mDjTweiB+o8xwGGwIkK/5BQYDOx
3ckh8gp90/TNUWiy/M0xbxkQ2HCx7Y86qolhWmDaBLPACTZFfkhWqUJSHOJ5KDt0wSBZqHTJ9Hhu
ixBciHImgPjWckqg98U7JjOQ7mIBDeRsRJ72E8+ie88xQdlLa2NGAPgwBRpT/iaHoass/rLU90Wt
2IDJYeVxEEjiXHzFy8YZbz+rTtozvqzyvAa1c9vOimccWgytfQkBWpH5gsC9KFaJBqXwnSKJZuNn
HSqk9Y9gK3X/32Gj7qRYkM2vCk527WZDomBLk1tF5zSmNMsN6zSC8Oo3LlEUzw89/6nLVqJPZWxG
CD0Os5vsoSerySzYfHL8tWiSITgVjZ7I8nM11/DHsPyMDCBGKj0rUCByQVScW0dQi5iAFlwXaPsi
tsPw9h2xmBYJRp529KJc7MHuKwSfAuiuEXH0oQM4NapvVhqU2X5rYczl4yZ0Y1/GSaKfqryWN0+N
WsXlJyGCjzoOhF3bIDv6zwoJ3YqBEvj8MJZC88Tvni28oyWj2hpnzRQeLEqo3li6EicI1okK4G39
5KKM3F/BSWDQTEoIAJswjQcVzGThEL9/gqeaC5CXuVgEQOZisnUnrUhaCEzleJBbEnfS0l12XfFL
HKxwFffy3LdxfycrwIFUH6VXIGVBI7hTY9ryh5KHYPYt9cmprQjbFf/yDi5LSr0Dp810uzL89VtV
nIaX4LoB9NLZSx/LFRDuJzl2nZOOuESY1T0KDpeEtVb0Bj1kiPkEB6UQHPdAjxbbIrSwS9sCE+y1
p9TnXD2xBqTn8pE3CC7PROelw3/PWkSpkQvBSAIw0GOyd2wMPS0FGP8WWSApmema5zek5c+M4RyV
MufEwy6SZWmajUGEizgu0Gvo/uSDRomKiZjXZcg6t69tnWc2/xUx/3lwXj1js0tBynp+nxsmm0y5
Hlb5t9V7kGYMhsJzpqV2BMVcgj0fpFD8dVwTYGP4RkwPsT0jChTAur4Xj7k9GaUtnEI+627ZGbmp
lddnfi7KOlbX9jQQPEEGibEkwNrxcyl+hSqAIS1wYWWooOa3U11jyUEt/TW3FupGe3yAlOLoVppL
7ZbBRiOswhQGYmI5dokWz5JQm1q8vvOFhESnXR1nVU+8yBScqfdvnsJ2QIdAQQg70EEdHT9azkz1
zTZPtdIbgc2M8o78jaFaCmCehnfgFLK5b06FiwUk2tu2SmNc2NTBg8EO6pr76khReXMhNllKjV+x
2a5GXQJrQAa4cf1WvArQpiTAwG/UOvIPSNO7uSeX1ozxj40fj7jxU3FG2b9JXA7bJHSrKAFLa+eN
fBZ69z6Fcx3z2CG1qG6ycIxrWWegPVq0WqXku4Z+55H1IDHyXpD0RIQ9VBiSXRORCavznm6ShjzA
D8OScKrYJAnG7s+hL5CSlHaAsl9zV9EqyHYHCrOTOfV5SpU8x/ygxikEgKAyDVrZPw5dt4xfcVCk
7K1SO+ZjsUx14HbaS5z+BQJVoungSwUbjCk356zp1DSg/lh1uqI3gSAuEFIam20JtzjOuGvlxweX
pJiWccHHKfzTghIxqf7wFNoPDBwquF9OtbgaFjefSujR54fWaadc694XC9K7osxvMkfDSuizHq3L
oVjsNAy9H8inGU45D7tneS3yPO3pwzGy3TCWyMUo7Y/fyBNhawzOmECnXPIfG+QakqFHabtXEhE7
MkvmILV/28gJknWrAwKh34n7PMQxqk7WJELbuBEEwYVoy6DzbqoHayjJcq+7ClpuSRWRSKhewylm
8FU357fBCR72dSg1t5AA9LMxBeZrc94V15X7EcmzEC/3DohcZdktuWiguOr/iJswY2RoOu4MKC6o
HB1MhKrgaeEP6KgpxxFbK5rDI4geT6hYCA0/V8p0J1jMv1Qb1vudnHlJt28GKDup8v1HJndQvuRv
mvucTHiR2aG9KHDYXYn/XJulpokIC4SZiCb+6w6FRFbCwWp/wwHBeRkciqkrbtx2SCSUNnNMJ9Rq
5UL1SVqEXYbppxZKUoK4o/GnESw9FTl23IDSMuWbR+x7Fwxe30BcbHXKueUWEn3P3d4vu/mEv0qj
c92GPo6feoxDuU4CmnZ+ciUDznHMkLmLlwX+fhzoYFRGHvZybr2EOlEh0un21piaLDcyW8IoTE3o
ZOI3USCUD9xkZqjE7S0Ln3QqJ4my4kBBa5HXYEauuJIrnEVrlD99vi4bos6aAvP7EKeKnKPn9hkw
NECGnAHv+YyWRDQeHg5Ye5vlytoqGQJ4sgHex5jYoZcLfRbCcvVrOxHLfhlMjnzV14vJTBKEam6v
vhyEi8Pm2bhNxaOd+MZ/PF7lh7800K7bt+lgJK3XxL20bm6E3h9V1bsy3E0nBIrv8jD8Wu+KjNFq
WBXhqmX7hALH3TBQQZoGIfp2f1sgtG4TxVM7YnWcEoT0jsu242D0lKSrsev8X+dMguuc7qt/+v6W
xC/2e5bxxuvqIHcnioN0Mp6zBf1KLvQrFO42coVmL5z4u5zpP+fsH7eMWXXYB8bcrb8UoIFvtkpM
uc/YyluW3w3pcpGaOT5LOah/vuvuGjKMuQWFzTCDFpW+a1zp0s8Gd6+nNyXNT6Dm2+gwJqYXk73Q
uKtm0GcwEv5H/25TP34ndcVfMiFmgXv30p29cdz4LDqy+DPD0bjFHEo/fbG+PaxQVJRNHhp0mpmB
6CCPyRn0UTMtNPOtN6zG2eNwQ8Fn5ILzEYv/a8kyMqj/o/iHinIpXkjY6DzQUvX1reFpoCIyk3nB
UsiK66QRT3By9zpBEbj1zMtykenILfACeYkjwd8qczP1Aa/h+ElGlyDXlPS683qHSiMTVa8OPylO
bP6u2PGkCGXExKrApfuVSrqfpF5e20aDN2uLdDLB2TwElP9r60OwnAzrEkdqTaTpU1l2jGOpnS+f
rZLpaaZzgqRkHewoxrEgG6Z1e+xyCXn1SlX8Ls+yf2gYVLYamGZrWiIO9WnjZAQz31B7xqVDOCSd
X59PIllZnzWRjOTxRtNejo4evyjQq4uEgsKwqj7st8nSwf+kKZO6kbGpi0YKS4SU1kdGghU8lyEe
GkRX9ERqapzddCmpkRmES7+A4H8N22you2jro+yj/ymHhvrG9f0Ryq8BiaBR8158sBM55l6Hieqd
YYiadldwMIO24aW5N5cc4cdu9pqf1skRhbz08HNttev0dTTEx+/kUIlBBp/+3jMbZSRqPzhZ3vac
7URm+456LM2ZuDNVxaOZ04lRrSnt2rPecjjjcEX3O5vu8u5ODY/NGlLcyHbuO4oUHIoC3M/FmR0o
3/RT0qrShbZ2D8z+HP++rkRAN79bHzrja2eyBa/qFcFlKSNpLRkKUUWRllMo45KTI3q/0z9JEXdl
bPl45mC2fCovt7hE0Ww2X7MEIK90sC9zQt/XVoNqJLk1roLe4a57TGMqav/tZTBS0nr4s395jmKs
YhLF1nDr2+eDHAaOcvq4B8Gf2G8+BYXpIPh3wCyCX4dXFgRs666bRMDRPGbz3cSm7NF+75stFHBo
8CZcVoEP+I+nc/92imRzA9SC4gikKfPLTdWFu1qbkg0Js9AQWO0Xvg9mjX4ngO8XkiBgetlYCReX
TTdIxs2oxx1I0UxLmcCOnyKRiBgEZHy97gfJRlqktMBVAP6ZX9vD3KpdwWmTlnEQsdsfP9NUkL2s
AxWdwPNOpSq85H7ZzHEHMofkH2Mbu2u6Qc+/TtpfnouK1x+anJJV+z1kHYM64+/arqA4PJLXYM/L
gDetS3tqD3MOczAo4pN38RMocd+8QPznRY1A7kVWFq8aryyHpRPBXZn/zhVsU+WyXyEooBF69Ii1
xDiyW1ObIoxGeN2ryktPgDzbABncFFETMgY1+pRlmNNuW6FbQXupMsXGLPpLPxWTntmypE+9oLN3
R4W3IzkdHH3Z09wQSmyGt/+M9AmkOa3v/y6OmJYp4oVRLmMl0rzIS4VUqiFqLLKkKviRA6tFJzaT
tk0TPN5MMnSS1ceWtohLxhRCNiz3qI1X7mxIu+kfl57nRtQHsfujKD7zW8GWBZK3160gvosdEyim
8p4mz2VqGHncdmT30ymkQIo6b3yu6rEH3Uh/COcv7n41S0q3onCIi8a0ENsk4NAuMuAGoK2bbxCp
gWEjtoOYDOQWXHA8wISsoNPGtHxXwYaxalWeG7+ZOLWTkj7st97c8uml8+1ZENwImLeyVFEGcVbM
SkJAnX2I5NRYic1iRHVE2sgklye3jbqtjlP8PCPSWCzhmsWYuIMDGI1vxjVp5eIC7GsrSXsufo6i
HTFj/GgQ718ZntmWtWTU+P1g+QJeUSnEOpLwgS9W4Thhi0SLu5Fufd+SlX1NBb6geJ8woU/B+JvS
3OVaBvE/RaqT7FtSZPMOc/ioatFiRg8tNwCtl1uRMXXuGYBfa+Takn+IQZUlumHeghsX0LDeI+H/
CrMv0Ay9legZMvkxHuLFw+8s3N2gaYwYUNwaZ2j9rlmTZLY3TgR98qL5Y4yR+kkkNa9cfI6hMc1o
T4eQ8kFUXPND8MBwnrFwro8Rt3zGpJUU6iIZzMOAWLGwiezOVRvzyXxkKVQg4Y8i2Jeyys98/yol
UuK7c8L8nodYANGZmzv/qy3lPXbKKQJUpd4ssU83izhF5gmlB3DzM9Zt/5i2ssqvirZdqPbyIcOq
tL/V8NnpaL9BNixjvD5oWAB+v+oQY/sOb3Pmc+QuOCBzT+DGOH2t1TMCjJF3DlvhwttAAlmfabfv
PE2jlYncmT85V05D9vwOIx9t0mKto81u/6AIbRB6g3uyLmbhEzSavN0lVJ2yeAds+uJtSJ53aWWV
BSHo/vL6tM7KS9jNn3TDhZ4WdggBlyTym115kg1Df+fpN5nNjAe/p4DAF+kXHfIb9HzU4hmlBpWT
kUDy6p3HG/koaam/3q/G47QxW5NeubOBWx34WSZM4h+BIay8/qADeolfwGKP+4+W7kn8d0WaXGwg
emUwQDsV8zV0e9irAw1sOlBW2AKh6XCjX7nd5Am70F0bUUow2GN5RUhS/fheDekXWVaHl7MAwup/
TjloRrNFASGlOyfITGzwAGLMZbL8W72On+VomjYTNwXnVw6OBK3JtrH0CHMzTPNx+Mrop5HuhiX1
1UvNfQyhV4nzLwGn24g28TBmj5c3h8kLLJ1X/iARdWpj8+lhHZ5aSHLq1/H8VEAj4jCaLwa0przH
gWa4NXyB8TZcq1j0JAnYHBZUf4Ai3KqTVzM8m7LhJOaKRfDn7//U3qtsRSp1w0Z9LfdgaVQTUX7t
nusG1oTLaBEazLPpU33vsZpE7Q5mK3JFtkxabxyQILYg7/vkVtgRXsXIRyq60dZbdvphoqmPe9vU
d2Syj6v2z6xZmgcfTj8u6KmO+ExrmIPh2554odEjzYgtiWWd68+meA9kF1f/8A8jbZ7anIxitBEQ
pu4/kJla58TBm8ByJkmJuvkUTVs9+bwuh8YBslCFp9+RTXLttYASNnF92t35oytmr8tN6eHQ/g++
N7aZC9ePySdzjglyoHE+kEuzD8cG3eK6I+Ua3kNoj2p6j3IKfjCRUjwx4IY4XeS4Dh01iR5a8XET
8Wdnjj7Dz+GzQSQG/pxwPJIL5s/I13DE3fMA73GZXRlBj30QMQEWzGh9i5RLsL5uGAxQB6VpQIIj
W+qDmBSKEhaQ8WyMprunrUWsF3Rym8io10m23H3M2gjIGeZAuVTp81ftLWsRtGATbPO8pJ7KLfh7
o8w6srxeuNkIpUonAMeTFgFMNuICyRCBzXmMl05H7uPhdMa+mO0nT01e3kRORIalcbFrYbMY8Vns
KPl6S/RrvvfWgKav4cUUfnJwt194DWmuHloxij3Emmpg0EBrLPBdR5ON5gv1QtqsCHGgkJImxGYz
qKQc+IxH3Ftsm8A2Cmd/oUpn37j4Fu6fwsecZowLzBSqwTakiWxCbIR3af4TYrYpAE7xZMpw61uC
LErXqdMr4BvXBWw/fUBZNCxrB5evZFPP1zbHpHkKuu65753TQTbaUQrzFvnq0lKZ2QGwSQnSrsYR
9p+K8BchA2cdUp7OK5ZOEiwi/HJ93Q6PYSPlspA/NsPTt/7O/HNvrdbSzwjguylz1ge+20CbYxCb
B82TuDEv5rp7E+0KHChqEBjGFwCDBAiK3qnhhYsp9qwAMKh2x38CNPoKqRW3KGns/szbIo/px3TJ
qkmEtybE/H16rYgozAgdXd61JaAnCJGEZhEiAB39gaVUew5Vtk/hi1X443G5kvL3IPat2xIrnqV9
Pd33FCqvz+6XaPhLd9JrYu76zHATSloKKiwh7OFPascXPq3JqxDNA6unuw48CfBh4QkJV6ebDU0P
Vr4b0KJbF1wnR5G756g1jPQWx6sE3eYpVgh46caUQpj5itc8W+t04yTsKzEQxz3NyZlmHrHb1G3k
GpiONQeZeE+jQMd5dfbQyxKmu3SO//vlOhFHJ2Lv1MIS+JosT25BDRsG8CLoTUMpRWe3esVsGJJ4
A3Vtzh7fKah9s0D0BUj4FGAwx7+ys+o31B8mRxS1KSuBu4Q2j9G8beHdwztQBxPNjt/LDWxkUt7x
IzjXhEJ6hxdVI9yt4TD5Vsb5PrM/qMq5kEwRKZPwYLnY7T1VBslRm8h+zGm46Dt7t8bdAVUenaFS
egeE6MERKgqM5Cfn9AHxJJQ0PLTrmWDPU4Z6LvZoZAQXLU+3zfGXKoGvKSuQyH0njAKHK/mHw0F9
UvkBjZSBzKfrhMLZGusS9oC0Z/wHfuDKcYxjD86nPfC0QCAmQ/s+GAzQ/4rMarUMVGmcPv5l1d+K
HILz4wCCm7ADFLPOfrHjPsZX8/Qs03Yo5TQ+XCOENPfVecTuHsxyFI9RBk2HA84FmpKqWzXQKVXy
9BrNwOIzeUU6qRkWLjaJBPTxqbxh5CyNTdmrvMgqwc0PBfDbwfpN6cwv7gpVMTyEfT8I+tXXioYK
l2Whal7WMB90aARqDKrx5AGUNpyihxwXuQmuStt814lra7MOQ6S54fftweE8TuyD+mEDp+nfH0E0
SfqY0U6nyNPdVtZlPFPMNX8q+d82XpvsS9xyp19ywf48s9pP/qYsrT4bJxsBYphbQdAZchCYLHhm
nAn9gztHy69dplzjSt/NTFoS0oij7s2/zidjpG85hubTmuXJ806x5pZG6uVLyykkUOyEmqTpVbYf
qlDRTUghLJ/gZY37MuKsV8OhShRRyo69csA9xk4mAoYC3Z0rO4+/RhYDJdCV/wwHVpEJ39imp2Dh
hnp2MllxeaEVO3Oz+KAuHrbqEn+SPoFP7KY42X+zlv8Z+PCbXqHlS6zweAomQuPjBXB6xbGuQR35
3Sw5vKeIx5a+VarVwG0mCvPVMLny/QlNKu7WRtsLZ3JQ2ZCC/FGeb4Ifbtx+r6xxN+ujXXFvJnnT
iUoZX1xlUkkmqy9jbPDhgyxbNwXnLs36G7CcTBdvOSvS0RivcDEur4s2NLlVBlr3ZyaNjitBPWXb
R2xuWboV0hmQXjQBOV8blJIGHuCSGCBdtafNcMG9mGxjndTLjRncaRBHNNqTtr3Z8eRe7AqYWMwt
czRwKWhkE4VW33seIJqNxD6eBeZlPvNyDjhe1ick8OKhAu1jznRsuoDYYYz8gapI7LyZZXR8Vzu6
TAaqRiKcm19JwgG+ZRVOaMzGWux1ywLBNNd4XYo4K/ysy48qMJr2Ly9Ouw5IYc3n00VM9Bwzm2I0
E4cjysUv6Zrl0EMTLhATvAB6ruX+L4uV6ufXpJY+x2b7thsJW1qdPTfQacsUs3Sbbn6nDPMHiAWo
Hw28biIenxzYaxDY8dB3/TDXcgBQ8dTLM2woAqM/WUMuVZEI+Y8q8G6aDdb+SZf/38a559KgL2yj
CmbuIsxKZuHdBvjd0KP5J9fErN7ShLSybNZqy66KZWvR2DtEIwzlpFP0WpRJIErtsrN/wx3z1KTc
1wTKnNmi6jg2zFTsdZOzn6XsmhSZu64NVwGEaNglDZ69jSChI7kK8U1VLjivzL3bUp3QTItbiNBo
X3GsdBcBnyDu9HW+YS44++wNwdO2h4PmdJfBNs+qcFLoLB9jvpkeRDKmdDTPTCUlcg1k+WcysmcV
WO/bxSi3PbVEP4u+Z/Pa1cwOKrxE/kcX+6yjM/kjUN69cOn11n8V7iqRUsqihP/M64+I7+sbNa1o
GyfILrip2UhBFsvoKETHzWjKfv/pWxfKltqMBqdlf7LiwaqlWK9hmt78Wbd9vK9E4UQxERvr/PSC
MuERlveOEzF1FIKtbbZ5aHWbeKnPf3FP+LF3T5mQ0p3Y0IOC5gp2ipOm6L7eXe36hv4+XiL6UfSg
tIc/uaezPOz7Ue2cGhmCwb2wXHu+3suqHfLZ9KceJO+MRn8FCbqTrFJwgzXPbtz6jK6xeF/SNFwe
/dixIEoFXrwpWSre/R16tt98ISW/ZHRKWZmgCK277FF0I+Yxojp8E2OZtVlN60g4d4vyYf2sqBiY
N3ME+HOkqb24Q3kqNX3/9qOSUb5Wk2AMgmDT6BHY93ad5/QygADN3NJsnA8jbObOKP94zalI6+hd
5cpHJmcjjbIm6QQ9dmT4ghE44dG3VzlmuVesIWyRnydG3dsdMlVsHLiUv29u38PtL7P0aVMvhymJ
vjQMsGtyXrSK1BgCzqDywya3fWX084D2nRTrHBoK5VBq5Gmf6sueLLLaFcj9DDgpUhIfL9nmNMOU
VjRr1GFOvYm7pD9xD6qI9JGi0yyQp4mdwWpGZWKZB1M/96AISrD3OpCNdbWyvHUHrKItrnY1RoEX
9NM3KzXjyAT7ebZiUmxJNPbPQ5NdYMYPH2oQutzY+kF4Xdnz3PVWTmORTw5Ehcd1V8/Dch2dQr+G
pYoSd5IVQEim8DTXOoi5nrpyL2bPFmLuIXtEgJ/0GXFunfCebn48djO1x6ldQ1iPshfet8UATVCs
sQbZ1CqWAGQm4NysDymwgF2Z+wUyr0oRGW6Y/Q7vjLPiiwaApm7wNyGEVgyMxdkeRTGA14vMNkjT
S//Uln6Flylvl7yWEVOQWf37lge4jgKc1oMW44JC6/cnCA06mm/CKe5SQmRFnfgKQHaYupVwa90W
kaTfN23AJ5YVQNv7tro7tQejdihfmg2A4+gU8rocEQHCF37QzPdN9s/YiG4+Y4PSIeVjxKniVWI4
PrYbtqGVcTw99tYMbvZ6SbxFGKQCdXayhyXMMIZcHiQr1nV6DxouhZHbbNjI5CL8G6Gq/shaFQ8r
mqBknbq31FDtJkn2oUniEoJjyohrbgqrhFbms/FaHdc5hFwDzfJu4MZyFvljnUEHYuJgrblZ3sT5
WW37e8aw79lWRf/ow+LW/oQxsaghnDL+muv8tmY5x6tCuLs7xcicoOzM6nMjmgO44XK3deElSA2C
Z0oCDdrGByQK5omUiTImBv5W78BYj5vbP1D69TtFW6z5YCYquqrFMvE7lnrFtz5xBuqAKKPv2CIv
PRvOl2q1jqICsViuUQ+r3Rvn1CglEY5eRce0Tq6G+ReW2iPwcCImipirrp1gclavU/9D89DJicXj
Jm1ARGjF9iBFlmUDpeEkxczz92Z33UV0/R6tndfE09xix+5yZ/DG/Jl/9wL5CXGd8pJi3NEnjy00
8YhE9TXraFypuCGvKHR0hyyzshLDklgK80WxgzTzmZL2nQ0i1IwAg9qim2chJU5wazIkfQ3EHE83
xS1ouwYpM7aoDIgwfgg+FYxY4cgSyzB2C3jWhMPp0aIi07PF7cv/r9lgRJOJ/RkHNVALml3wwDvE
EUHmRm6nWCHETy38mSEb04f+UIEdA3/0GN/CXVREaTb+CXY+Sg3iMfJyyYKUBIBMJJ1nkIqd3SBi
qQoC0eP3SUUHGqUR+CRfIQ41YwRkXb8VQ7vFDi0TaIYp3E7Fxhn/I6dehi0dhVA7aJqiR5ssBmyH
i62g3N40sH2zVCuGxUnTXY7NwmJYG3NXc8BaU/4Szgrczh/p5NY4kB8dJetyeIsKAqICHlng5YMp
hczCU85LYF9qi5g/PDviTbgfDga311lld7Qvfs8HMCn1vB2Tnz3u4tpCzWWvmd3rKicP6WP5jEeh
2tHt9+pqXxprQa1F5JLzWrMpzDSG9bz0tleJJBkd3nPX+4SKkdUWY9TTtbShALGXgCMQkJc1rzmZ
R2SUR7gQ685S3blUGYF6vFj8Ewp8PkwUMOtEnx+NDz4Blzp4SFCG4w3qffTtLJEWadhC8mzNSgRo
byjaTZYLSfc8BOJRiHAiUzMKCKLp8ZCAZl/PmM5PadxkXedu6mlUHVcpmXEEa/AUIGjYw7bSJuLg
BsHsCbmXRrmoHb2gJJuj6rw7aE1gqO3r2ok7lCf8vSqNwnhWmD3+uAP7D1cQ35i46pXF4Tsl9n8H
tC3kxvcxVXhCNBfQ9L+114Dfd6pcT8ZQXWj/DSRRpgc+EtFUhGlw8aeeX5BK74Bv37EPYV+m3/t2
vUppb0lL+FYrQ55cioo6dzuIdUulVHs5BnlCnYV7F8o9ZvnR6UTiB0mPT5twcYyo2fW/LCIzjpM6
JpKMAG068uw/Og/a1a403Fw0AMO66Mxo1f9N4zPfOQYrVVfWcs/1spB45bhKjK+HntM50XldTNIg
oiTM2v1cPA6C9bgWxjhrFbTojA0kQ3SV4R57wYyNAca0axcvhMYIotQTK+/wXT58kkcVz8BVjBqc
8+shf0O+mkJew06YjsLlVuxWFGB/dfWh7OXwg5pPaIwMovSucCQUWZQWlMH8KGG8n8TnL3S+be9K
x1t5j/XVeZ3tMB9IYBuqbC+yGuVGCnjPBz54nIafN8dwmJ1bzW8ngJJYeXOdX7M2G458kkwgybMv
SIMzfAo74idqx6Brk1/CBm926+1YRdyEY3wxO+Ap0Mxu7hxGCYiyZJq3B5FWeHB7og6IrfPT0gNO
3VTjqChogeLpURB/xU7H7k/V6Gambhp+nTW1O3T13nVx2tC8GJ3X+Q9Z2GqCS5wGNkDsl3Y1bSpV
9deErBfAFABAERD1XPGn4sZqsdFjNTqDnD1/AcYDN4CAjPOR1quELXEAf8Qa5mjVs0BM9KpK5Ycv
ZaHoj/hrpEen+uYY6ubDW+zv1cSLKrfVjHaWArudXiu9fFCdYqmFlPe8fmNOyyaXroea1bjDBLav
hoCCEB5ymR0drOy8aEeI07qpYF1e/K545+q1c+lewfQMBnY3kxeL3huanoxK4V5RxfS15E3SYFAU
GziOfOjSVw7kDNhs/3Z+CdUAaeQLJTQB2l/zxr04StIglhLMoXgh5RDRPjVhuV+nFLBhkB3R2RR8
ZYPR+4oU/uuFnxHNDb/zEypFvMpCqIuzHk6R8wa9ueeJqiaR2omchNvPpDiLTZVaJqV4sRt7SRjp
CxlRxVFzc2z0F3nqmUCrwFBIDmRPqBuvIqpNBkWCiJ2UWz8r31A9PJM58xIDK4gfyuVsY9YC/jQW
LjQARc17JPeGF8cnjkdmabwawaLxVyfb/VIlEJr6aymTj5IcoN55yb8V31jkfFHdJq0Hej+jDFgJ
Klp1EqHRgOVid7Fmx2z1AaNOuHttBogxOedN4TxJf7/DII6oF48M80g2TKrUHyj3XMpdZiwxanp4
cv3sRouApzhbru1ShATGIW70VNk2PVHWT/CtzIY4Wz/F3XkhsIaUosQTkD3MZr55BUsuWAKMEHRf
JdixGVDKIGUoKi/5Sal8CVdhejCf0BKskqE9x2CpTtVnx1QTU9Cqcyt/zSqvydnkHOy6YaSCS+Ch
R7M0UOk3v5rTj56DfW7H3Mmu6zzKIZ7xuhdpVlLvqfKqFw3xTmLn8OmyWCtOVKbaSRbenBkiX2+6
YeFiaT9WRZghhmqpLmJiY4UXkFPiPJWnTuB2QtEk+J66C+k2FkzRsI6iwWR7V9pBPB2e6bXN6oLU
M3XVfUpL+KBFKY33MDa0AD/Unk8wBHOdkXTIgI6lBT3Y4gC1uDfHc3k1mPWu51fCGRAJVmvGK3nM
X1Y8+vXF0gumdXLj8EZMVZrqhtN+nsAGsclYBEBUQEmztgRO57P0Us8d9W6rYhBw0Kq309eYHN9r
VMfXcoa9Fwv5njb970+0c8kIAgG/1T8L9Jd5PHtnBpT/W7GhHSKVN9l4q3wZ2T6w9a3feBzD6rdG
PGmv1miucfInRvvuIrE35/f2OprcYnKP8qfr5NSGWCyADJO9pEM5HrsqvA/x6JdNIXMOMN68Yw7D
ZvOi90D87QhYcIJ6TzyBHgctL9HyS6K3KQwYBFxzlbp8/XlsbAt2dC/ZiOl8p5SpWYmAk5BggsEg
yqXEAinkO4l83+rjQl0kTQ0ICoyR2eGm4N7Qj8LSPLDn0VLlhttgQPRJ2XNSq0+6oJoEfV5pas0c
cGWHn7G+O029QTR0KYYOO4aAafAQmHv9zEhmBadOZnQyu1rAboMAUGhSTAyIbKldaQolRQIPIqZ5
k9xIbqZRDmi18SsHOZ1e5z/lSCkSbxFHAfEX+lslOKqbzJ1qSqTc3gGoSb5NFWWVlHihwZmWzoZJ
8UN3KlIkO/0mAJIx5m3fPLuSKnrNWcFE9g/Iy25F/cWfn5rlsgzni0WmbsQL8gIIZCqkf57BwVHV
xDyHYLI7J+qRUMpmTfnenexdKvfxaePoi3lodLtAiA8AiSerfZ5KWUFORhWZsGz8z8kP9Cxlifj7
J9xN3yOc/59SENxMXbjKyGpsaMJvoMJ2Yx2gQU2H0qNgwrOdsM75NDQa0GrEiIyVV66f/EHQiBs2
MhoKvZkdMQC1eRcU8QqqYLKsjzL+ru/Lu6zii25oIxlzdth9WvOXgnLya3ThzsaUwG1Yx4cceRLp
hUXllCQ15rRS4XdPS/McjpSYGM0xUwKUCq8JdaR1jHT6NjB8lot9VYz4dO90LcR56uq2frZkYLeZ
qNv/hla19z5biAqmwSnzaznHuzA9nziJJiIhWmBLl+wW4SJ/D8u1cEqnq7ncmVX+CVGmSa81FVDY
WdA9u/TpnQqBw+unmedNTOHnR5U0GOzr9tXP32uSVWaet32jbu3dyiqfhd1Lq6tpf20qGrc2nJRg
dgdRBn5qK3yBrm7in7LfS8YnY6IT3uhLNy6EqPY3dIi16BdejVoPL7SMgOIWhacay2jVMoSSMqO7
iSKpKEJSXS6ZUhMGgfcyxkB63m/Up2J6dIi4G6biiAArNAyQnKGJcNyqGk+6TDhkepB7JrWRsPcM
4pO799gIYxiV9kPNuyABvdEg34bOqB2GwA9yGqGPIQqTsuVlaOxd2jW8BXvxwYLtW4LSavGfvjes
i8mTGtuRUnzg3qrbef9zAliusRvbEUbIG5P48h9S5BOymWnbkkqsJw3Tk5sW3eLC9O0IDQ9R2hX5
lpYUAZdgFD5OIbhLR+bzVs4TclGY49gSOxIASwR7qlbHI8tmnFzdqx6Uur8XZ+0ZkAAnxMUEE2pP
pXy7WkVNFUc/+x7fvvRwFPJhwq2AHdUYwglBLoo3iOMTpNWazxazzQmxs8/Dmu95nCLruWqvY8PW
ufJdthKwh2i609rlc/7K+KPb+/fPrfvJrsHEPaXd4zavBm1vYOKGOlXQ8zyrMWiseMVZFYzRQfUB
yeNv5gADXxmYE62ZKIzpRaWiS3tsoXgIxFdmYmtTZtCmwnJnsmB1uLJ9+ehwqogU3k44P9+VwllX
QYFxaT/MsNgU6KVT1PTBEfgj9DjwFHzCB7mhcUC/BVwYNej5zbiWFL2ibffwiqSKjNv3pPjbWmEc
0qDaqn/Tc5j5jwUDIiZxegBYZV0IjUuJeMnGs+YlkjAgRWYLu80DYRLQTV7VUp9nNiLp3tu6qZVl
KcfX+YaX+fsSvyJqvN+Yt9CPi9wdTZSRKZyze9FNdAhSUGxV5+5ePJEO9dk3s0QYzQzW3xi3oMeG
e8jwxGuguOgc7RGUr9oNYDT5vCM23b5SQAe2RLiigurwa1icFleZz21dlI7NHDPBEVdUlXM13Lad
oNG3//q0/y9OHsHWyW1u6wJrVb/ki1s9ymG2yHFDOqyZb6idXwF2EqiDSotukTllq0XA8BG+M+ed
mTfsDVgcr+Ew8tzQOlsV+hkOz9GyteJv+ycDE4MpuUGrsAX0KnzwjpysBmwzvkf6U8J3yCJzoi7y
XoCMEzaeSmMOhyE3ZmkoV4mlHHLBirftF0lIYuPp0+/ZWc+qrqB6+/K0YtOaj9PHKWSnIVGGs2uc
p7/zF6vrITOMgJR7iPmTnaEfFItir/K2+F53PR8GUfa1iHj5J65wm71bOrOgXhTE/c/E0V7ajImw
mJ7oEjAGGccMuERAvtbknIOrn3WYVhyYZ0SW+v2aK/H7jSmKwQ75BkW7zKGUuCBSY736Cl/46aA+
ipPRG6jDh3tsLU6+IYXr4AMZ7mRJUuwn2IPfaEME9t2FAqV0iJ3FoLWBIJvXV7eh2R36lHYw028d
Pgp3TqYbav0qJMpfQaxYgSvHTjFetIUMOrUzN64KYYSz09leVga65HsD8Hfm5mvwrAGcTb4l2Bt7
BgBWMUJAHF9+8wei3g7pUTkALjYIhdXkWiogbgqKJQ8bhBwRJ3vLAW552aweHNvE9/JrGW4+81vf
7xBkWM6B4LMtRv6JhL1gePohyMWWH9CN2XcwHqwHOgThbrxXhLlDxkWGz36SrcwZY5hvttlzPej8
dAZHbgOGJNBnFEjix+y76AnAYzJQXGRYroIm+v3GEN8IXj/kTFpsX+zG7oRAEkIs879dFCzsDxTS
hHRQFTDNpvgNb23ktD+Lw0NiVegJXOq94/o0fliEWyoLBPWCGASQqgnnCMTbSRYjXR0gZYScS3MJ
LpJe0nr6N+fzHt4wPonI8+4A41EnIsygiWuYqwJocPwey6/g/59KfhQSWrbqP16I/cQP94oAkHtq
sBS9dRr8JoSFr5MvF5ouLJbgomIjJEPr+m4L6e+uRCy6RkmewXeSUrq7QiXIdrUQl96dZK9t9cHi
QiE4DYSP1VkziJMSF16Uu4FQ9Van0NvwPIEWI1+fRUtd2QhDSsCBgsnMq7qpfhSjtsCtXNyD2p7s
L9ykg1UqovKR1zE+c8zu7X5ZKDnXdRrhRJlJnJE4H66Ndfb8rkqIuwAJZ90Cq/+6w7QRpBm4R5OG
DFxWXttysBEO5FTvlx9Ly3IwHQiGJQpBiOuOKp34ABG6As53vRktikOimWJISUYTzMcBzRaZajqe
Z86W5c9M3k7/EQZ/mv9v0PrUCTc/QEDv+K7fzziwUaFZqy2BvXadNVqFdpdowd+dUzt8a1PdAgMT
6xmjsGXKZMU2BU/cijWnL//ioitBuOTvq9sm36Iu5LK9Wmro2K8uF7HlgUDBLN3HvliN8+GCRZJI
sb4BztmqgThwW2gQL2TjFJkhsi+ywQBcVJXo9Rz/UJjjYOFmwNOJjlzD2ke9mKhGifazxfBa0Ku7
gtGnqocaMhuBm+ZAD3ZpIfiWFn2tIPiPIMthKJQmPmhb7DvMaQ/X/rrmUY191JM5N5HQI9DCmhan
3WSkPw7f4ZZlhbu1UNuowprv5P3Lz5r6pQJCvIAgtMwzUSOcribk09b1NsYPDQdV2U8M6GzeKcw3
bwFFpENOjQfL4pcebKV7ZE3lkozXagFuqVFkkQay5DweKHNu6Zyq0Zy/qMYtsUE04FygQrHfLNQt
2T5TdtHVlJLnOjAAVmWAP/pl4/JdcP6+OCClIEWoo2Ih2eut3sHlgKCdIkl1brfPidJMtGd+5Ufy
cFLxdV0BLT8Tp9LuxjNeJnAERqawR9Wz3UN8qaOyr8U3HOCqo7zSrR9oQ0MJbziy9uCtG16fo/xa
qhHqfDkvZTg9lCCCMBzMKO78UcDcSpq56SQ8PqR9kC+2u9d2K3AZA2tM4zmeWJLWjtE+VYuDtErm
7phSCWh7h9wTLa+o75MnkPkQBqj93wljqzLb4I+qWiADyAUU6Vy/G3IdyANJgw0H2EcZNl3P4mg5
SLyx7ILwZZ+rt3jk9o/lmZ2o6kWlj/7mZNJSpXVw5llypljTM7TXw91dR5B/HKnvjlNjQR/nxJ0h
jsMeUoTHGBquV83Z9WFTPfFRKmGK1VFmdvX8v1A/GV0HXxqeHBfPzZbDBKcmseRcsjCvySn+hpG6
gOQcY9xRwoaRuV+ypirLTpg74swM+EiBzgGbhofDzGG+CG3KAhiNUbQydqM2nq3Nf0unRuV7u9BP
8nQDjYZjWCfnVdeOl/MKRaMA4au5RXa+C1MQXKJ0ZgEHOvET46zjOLHpTlJN1trSW7UWhVoaGE/p
OvJ26Qj6mBAHeGN/lR1Os/RbkX+n3FYuDGHRdb/k/xRZPjJ35uOh3ECkkBYef8nKiHF5CHbDjNkk
7hYZapzE6yvIFAvvRMNcgwbh3Q6o/FnOVMqXRw55t/cwTUHoZ6wumwLldyIgFWFNJJM4463+sOMF
lwPIDDgTPC3MOW4n9g2+j6bmyjRbMRn/AWpy5VxbmUAQ1ZpJ5B9QJRIDbtdl64fHOTK0DkxZKAIC
XPbtaRSywEOn3+0076lnvGg5g18iw0YlyTH6LmuSVaA2zHD5zsPT+cPK5P7qBbwjRUxirCD7LO2a
3hr3+wSqrbJbc+UOolSEVG1UC7uo145ALn6A0LJN4nwXbf+ex2I9hOAgLMZm58ZAbkSx28zsnHGF
W3qRf4nZ14fw2tUCYXR84u1VLyESJTxnXXOVXM7qCU05YPAeLHxp/k9AAZqN/c00duw2LoDDYWoL
KsggJSu45ND3RD1HMo5mILaHcrtNAQQBXtRZRE9VfNLPVKgQiSoCYJkB0BVFxo+0OOhtaHx5m/mR
NmqApo7EHyZq4titVLAhdbuCJGqg2Jj5sr0AVJvauqXATBhL/SggQn+gVAO2yd6AriObipYYzi10
Un5FOCv9C4YxFT7JAzua7YfazI7toZZZohcLwacUmoTJvbrUk6uCqEvLFwwiuRMX2kg65sQ9y8ub
qIo6sNw7Dhyx+6QhT0EyJztuC4wx4idiJR9M1m6xLTfkQzzbuqete3zAjXbPGcnhBXxQz9bBrf4o
StKSCNkC4Lgh9XTLEaPCAeRZy4oWRHjmDut7yXogzWuyssGIBtE9psy2GuKNKia6PL0dLexrLodq
VCVLRIUM9tbffmjxoajbUeK3XtoEi1Ss+bzXFCGqbpxOHxrydWiNlhLKXAxELpKGwXZzUg6kroaA
2o8ZCTmXONSkIMp+bc2kK55WNaZHWYh6ahOZXajPlRVlyoCKqc1FBm3R3ahJi47V+0r5KMyab21x
agWT/r0aclGqkzcvzfI/yu6WizPM6YpOIiTIlAT/G7Itq/FmYdRAvKzMEJeWbiIMvmsbdjaf2QqH
y4KAIeJVspelFxhHIgpTebd9rwK42oAlDRvjS4yy7F6vuykhptKbO62JdSPM/dj8GpP5ujU2sQoI
7zmbzsQm57BNI9tlECWpSrb4RiVwBXSxEoFu8VewDHP3h41u8W1jTOcbl084gBydnCJKd1FCeGlF
ljxRQNB37ntnVVJO2oTUfQpOPVbQlXd5KUIsB3mMCnhtoEbDPFgBNCfPiuiUoZ/0sp+7BIg2rcS5
BgJfIHKfVpUCuh6GC/+EPYzP05zp1hWyU9xFPVNVJrpaD7+pEN2LsnevqIR8k2P4n6Yx9dUFVGnS
jfc0aZNKnmotjgf38Q94xddKvL6CHRFoV6BTJWUw7UuedhEUCLLIuhPKMublf79+GSVIsdF5qVtT
Zd63B+E7yo/FF4gX+tgxvBi+il4Yd0jB69YJtKWRsEkfVIjYsE9j1JUkgNEk+iEngugxmKoJOl1D
vnOVs0OvyxuK/pl7JNxsCuAl9KvLywhbvt/Mi68fQUZjHphswpgGPNjfGL/rmkwRTLtCqKXMG5H9
dkPZjRwzdPU0/AK1qO58PQXqrj8VlM5P6aWhJSDaFLAeKWY/3uHhekEPX0/Zf5Fv4RMGaM+vJzey
jIzX+6YHaKtDJxqGq1BZo3VPl4OTsabwLOOuyqznSkSH7UiT/u3tlG6zF2MP8095R74vA4Mllc+g
wgBaDybD68NwkZD4XvR1q4RzHAOd0QfsnYXxQzUsSn86LTVsiUhriPG3yG3I3WoRIVqJYc2BJo4i
Lb8+GvyfmIinKqGMwXGdLEDB46ybW4nsKko/M0jd5leViih0BhwnrqcOiGHSaYNG62puw/h2NFXi
qhuCnCSGFQEGel3YoJ7I6cBtUPeTWBCspSI464huyctCckFsDOU3s+LU35hIvvprv9ZtVIv7SpP2
sSrjPCGErFhpqiIYItbS7xIN5YnPgodaHm4FU8cD+R7qFQdnb29jJPS/sSMJhp4PEFwBJA+4nNY4
XdKIWCx+QxzrLCrhgtoj8kgt4T5jRWFn580N4RoYzkqEHCutbzbmqKI6icZgaw9X2KjorRqhtH4B
cYwggwu51k7OSFNo0aCHszH7t990uWFku3nMJIzX5Qh/xbrhxjj5TCqSnXBrNP0CjQttdrA1VxXd
PhmzFcdY2q/bvjEh1+fRTgfZt0QxLkkjOThlBzCwD4pWlf3p2kiLA6JkzC+6h3y9wbMIj1k7zjwf
Ic/lAsV0kh4Dw3/PjFLzASpYiB8kHWJbaY5xNUD+ayujuSA195mrQEoEplkPyhkx7Z+SO3snFyA+
Chc/lGfEvGgNf6Exzt/XlBNvBqUXmi1WJGzgll5C49xFV1AVuUtS0j1qgHGZEx3D8rjvm0NVs598
JBRrqZDQ3/+B0oKSepdR0IJJv7Pytp7f6VBMXvmRAOWOwfnROmNsWvM4dNo8/RSKtYjG7gHAB1rW
+zTUzRH+8xgSQ+xGqYwn+wAjFifKAxnI47+njPkHv9IhzCVdxgql6nSLjHx2XYVkHlBR/lyjnLI4
cs9X4dxy8AAuFWblDTfji4M7VMPylXo9QJejXlKepZ69DUu9axLPDnEcly+N+An3kloofgW02PcB
WQqOpPTnBIYYOs7VzKef8STYBltjvTWsuwpv2VGZYpvGbrZbwKyN9z2W7/fLgRKknnbcic2EE6Ey
um5fIYJ4Dd4JO5it29e617Izw2goT/gJ1LRMgrFinCCF4bUIBXEa5QVdTQIMOELZAD4KKFCrfErH
1G8gX1YSBo1phA02y2HGloJ8/Z5JsVvxHR2DBjWJYvqPtmSh8Ap5T4rG216v7DYZMcmNNbnTrOtd
72DAcpu9hiyEzD2HJ0UH8Gtck6x/+NtOBcp1xfc12zyNdoR68iuTi8xPQ4umCdrxrVdb8bbandF2
fqZ7Xab/AdDr6juAyVo8oZ46ds8t+nqZwFAyPbq8KlXrf+NYC7bPNjuIpGmZe4uqdAwSoxVymIVk
Oin+47N8XmOCO6poisjo4EwrVIyqd+IZXoiq3L7YBoTyxVWSGfpbifU2fidoIc/b+41FohxmupNG
cXMtPK01nope0E1ijSLD7WYn8w1Bqy9oMSxmMNxXQdGlSZ0bJ6TU4fL5vItkRqR8MPszY83syZiP
aVb2H1F03NkKu17CalZ46j9zVBacbVKqwAhvD27Jl9m7DlK3G7jx644Ny/ezMjWKLWa+mIPKPnt5
u3FnKuiQpBNDGlpvyBDN//3n8SwRJgJSpQJ5/EQBO5FdqNysebv2aoFY4JoCfwaQYbX3xiLJtbJg
rPIE+kOuLcsrLYhEZLVFzT+MJ16eYTRXhq1mQTnHFzCEemDY7HzCmgQc5jt9awj6GQKUm9/p5clA
eOzpxBjQJnFD+xlX8IgVlIvpDRgZjXwiRrx12p0VHGH93pTFyORc0YBW2nhZzu1qHMWqSxWiaZ6M
LcjKrTbSYGGHSJmdp/tN8sHfk4V+wXiybT98FZhWJZXBvoJZPFMkWvEPn4nZULuFr5co4kZvQOi/
0aZwx7N7vEUVLtS7bVn10CW4JEuy/a0FIND3D4axj32oI7EOUJNtiN1fugkhRO/g2vPb+FSj6i71
OyqG/vSq5KaDnv58LuS3GChWG1SnEhY12aRdd+CRtcBdFsoxpXIMuVaP51v6b4g2Wkt0Kp4I0+q4
iSF7WgU6nu8DiNBvL7XX6rU+w13mYAa1dZqm3EtxUwadCxXQrzFkp/YfnCd8Qz8IQDiN03J80pzr
F3RalWJPoBTbETXuaSc2LHTS2XXyh78tTqwRhLQsk32FWvlGFQ6NQiRPpjF2DY4woD1BU6ipszlb
BORZwAK00OPiXbQwC7vupO/LqRvT0aRKJpOIfe/mcQezFezH4LdnS7dVZ+fWBIYo0RiycXiUHf0E
ybeYQ8kzC6drckId7j7X2x4YDcwUiKYHa+lD/hdBO5UvcqaVkUxr9IvXztrW9pjhBED4ZGXIWV25
2HwBgtEoPEnnqPY9NkJQtXq4bGd1cKH1Y+kn1XRgOpAaZNXVORjKeXd/9KlAYGN58+UxoFUtbbfH
wX18Rtg3Eicn9msJU3sRkU7MXCeCCKZtJsyubwxf3mgfh/tlFEjBxZzRMlYpnix2+eLMaEP4zcHD
p0icNR+GcL+hnmM4Ehicbacc90W4Kyqqrf5LjnpvGgJdSQL/xnZe5Wslgq23CqqjiedK5n5FxiHH
Wo6dTPR0KUdxlkrbvpc0qstKzwhJGoUbF1N6vhHxtc0pFuHCxq5CA4UrBTLkLIHtCtWIxZzXcN+e
0yUZLGO68SUsXRSZnpasysZzaLnJPrHDTJlu/vGw4O4ia4tqya1GUGOUzRTgIp8MtaopE+ciBZL4
iaRzjED/lm4tKP3toZgncmNohiVK+J48+2yMUR3zEUIieSZmNBAHRByZ1aaC6m+RSMpl+wDh2pOZ
VhufHpt3fPHsGQY6X7EDrugNmDzyxB4d3wAqSHi0yW5DlC5wCC7vqam+rkl5hIcxpJdjN7jQBw6Q
eVluaAyJ/w4lHI/URjheNiY/f/etj7HTu5EpjdJrG/L+NbNOXMcojXD6y7B+al3e0TJPEiVUW6av
CVtb0EXV9XAAsR3qjq9n/FaGWpePDpBi7lJcKm8Is3PUZB+5Z8htWMnHUVfN1nlZ9H046QJ1nsPc
N+1wgkw6I3XjUkrditaJQksg3FWp1DEuSPKn1+4q41GF8ThCBPx3QPG9KuRsFuHB4rYYmTVuMv5Z
RdnKl4y5Dgmpa38c26xAsziUIR2rbFtnIFjrHDO9BVtbGpAVqNNNvnRhoZGC/ebPmxVGkMnJwwX7
6V/wM6gxBo99/cT/iWBkm4hYYEXQTOZSlcpcjJzc2U5pVf47AMSYPj0dsXtejzCv9z/wnZH5Qslr
keSLPcjh2wnOGqDO5yx7T4ht0MADeSTJp1sKHWGTOZTw1/P51uh5BinqW0fXf4+4NiEA/yt825vu
xa3IS3O1rk2jaCWqCR/ZxBihQWfQ7l/5gzZFE7vOdlvIGkUXSM+JjLrE0HhYxZYQvUafLg/uYWj+
8JiTlwd/DEC7D5mf7/LBvvaxepzP7Nr0Mdxrw2NE4DyTLgIiHuEnOD+aWwv29M3IxLl0c9LHqkPY
kIUP9OtNNvILEJvOZ2nBi8wyaGPOdNGQCyT7VU4QopX6YCD3cxGbAspgiIVZVj9IOlwTHkTYfQ2P
fX7rCh5Gy+ebsZPTt6Pv3ngi5W3vubLpR/IuFP/R19LusoSfxWfi5GkaC+BpdiyjNu+XnGV3niZ/
DFbj3B5ih7GYfnPariG0ui0SgvVqqvTx1mlOJW2rpKTr3iz5t4oUOMIh9WGDu5cFt3sri35qDk66
dgJFVu86f5mZUI19iWeOV6CAXGzJOGJXjpkc+w2RhOYC0WUA98XEqJt2pYQB/wv13VW5HCFymsSC
d4pfX+YLuZEd95o+swrFx7lPsFIrJQjV3wqOZdNNFbGmbpUL0L6IQmfqi4Za7eDHW/z0ljGdk/VB
4wYaLL7TE1a1Dg2HQDNhKGK0qg+Y5GWH8KzCjyJDAUOL/I1WGKBfYGycokUSkzV/yHUcOdGzwNFq
35Cn51bs5XLkiJlTLeGeCPuQ81l3DIZjLN34xnJHBOiIZkjjeSCxV/DuwSQqwrXPC9IkO2Nop4IP
wu+UvW1jqYsY6QLVP6pr1zTjFalYuRFeSjlCl08qKR62cIyKeZpk5uYyWHq0h15zf7U2f4TLHx8m
hhLsMzly1GWoTPu5DhPejk9VinCnOIpdk2d0S7V3z5+SMB7SpI5+16ANr6ON1oqyIDws3io8IPGJ
N6toySpXUEv2GOg8wY9FjuJ66prOgH72wgLvB3zoLRAzOmWZeJBbbnEfwSRilnDABPzIoso1+1Fs
FBfnJiIgLHyw5zd5D8St8RsKU6Cgn04KCjp4ob7JBngO4MzW5bbQk1PS6+CBE74uPXAuT/v4WANP
imZxqwH5rb9K3mKuBtzX20crKi4Q+3P72Me1OYKwSo1qEehdk89FLuSSZj489Iez/GHa7aZeYIn4
w94874GNMxZCp4cUiZvDlbEcYc/HQ+bzTSWgOouqTUIPlZnNG9SgnLiGiggKIHGGjGG5XzeNZzAD
04dljl4JDiSW7F6clUiqv8y0WIe4uA6Ae28cAaeKaZfOGGuVlh96rk58KjerRFH9ZenkhN84LiEo
w/YtkzVQI4YCq9v0gE0rkZzmjfOfTpxC6jU1naV9RJAbafuNyb4+dziA878cHGnsxiONHjp8nwmJ
qg8UQDv9+CkkGDnjUra2fgW5PcAhHfrNhmKz3GKOtKS7XDN2qF19mRGnUXRPNFoNF7ryW0aAMC7o
br7Up+0tHkalKW3cuVXQBR3MUE6Dk4lwwT2Lm/z6IXlMjiyC1asDBJNi3GjIpyHDcdurAyMjXVlz
96aT9vbM576dQhxNLJnQi4osonDUbBZG70juGPBc9hYLHICkq44Ay++QP6i7Fj2I710hT7NFE1Rr
cMfXBglCdxmT8lnVUw39CAT8URG8p1PGyA5QHN3cZBlqOsRxPEGwD7fbCX21kuGTMTmaeCGUHzKI
ivsl+hdsWTI15rA4WfpKl2pygK0sCzh8t62wXlcCimCqh3PDMM9ROOx4Zddl+5gbxIN/6mAShSCM
wNbHWafVecKquANL+t1otD0YpZduW8enPjpIdMMHWLLzmG/tov7sGW/XPsmyluuWDj4A2xaHgA1C
dhl22jrCdOXnLSdLprdbynHqZknTlmsTsw6KzVFACq2QiQPcnvePRQsTx6oj8wAa4vWeZsXB836o
3AkPacIV4ZRX8Ne3Z41aOJ5MEBdz7v5nfe4lTxjssNHzZ9STMQvcq1GvqYbV5pgD/zkCFba5Nw4X
Gr6dBqzknrxphT3pdqw52grUiqYfixeRj00dGG+AekUJqBQnlj0Axa3EpiiOlQg6GOFuv8pH4iGu
hbraG/38xFl6gEhg7puI63UhdUcz6C3UVnqy99Iy5XBNdHuGIf7HiS5P9Jtm8FGtFkiUzkYPY+yg
a0qixWwhZT87qtORKGfpQz0wTsM1ZlxXBCMa9uK/2ACZOTFiPEvA/uzq2vU0slQ1pkuDaVIegaMr
lTT1iOV/E/90MasPNzvA43LcTiI9HbxSTEV0mUk0D+MlUKSu8tQaN6RuWFCK7a6cV+6smkOuqI3O
AZ51VKnC5rfToAH2JacEY020oDsvOdnWa+aNncy7clFV5NDSWMcqA5nZPTaVkA5I0IDINdE2BAhq
hWIxhNg+QWDVS23Zc5GcUyxxGomFQDpqbiq3TJ0nJMJegIxsBtSXgVNAKblUgVFgm+9NWAj60KS/
UYh5FZeA7p1AZkLpBaPGV3FII3dLE6Vnohbu3TgKlfMnhHBAdyfUw4ndQxwEH6uq6VDowjzVEzj0
GI/Qvn5885mT0fEG3n+BHQ0Il3R08uLAluogMpcAmsTK3bixIUMK5c/uLdKZaJ/uLjK3FCbJ/p+8
IYOQ/h7xN248E1XL659STxa7A/C33FcTWx29SDdYidlktC3x0OClKrjYD5lnuyUPaP7VbBeg+K2S
IskleqifPV+Xxx+gy/yAYm6Vq92xc4ONjHZVC7iqU5ui6if4zU/rt1iY5xftfHZgbbSswVYzwCbg
mKkYI73ZsYZ4pJ/56+g398neH2VVlTYzn92FrfIX0uviEhJd+bfJy7/vs7EoZgotVX0ISZmA/kCS
XJsckA3WnUGICg3qlX0crnlV9zBVPB5XpZwC8V/nu3ncElF0vZd4FyUGZTfmhgCSCT5fxdCF4XFT
T7Y8CkYur7l29ouxJt+tNnDptAIO14M0z7+spLl1vQWsITsRnTFDppxVu6hVsNUMdcamTMAj0qp0
vIrFpVmC84Qm+4uP8wr03OIyHLXlEkrA22HSWJfYSDU9LV/kW5QXi7AoJZ0HKr3kZEiB6qI9Vzf5
Qdb5w8DX/76pdp6IK1sR2oN3veFcoOD++NBZPVYe2QaqBDyPSF/V1GmAuLp820yXvlGFDf5jMFF5
zlWoskH2GOWJ8nn3dsb30TJOkgqJpYpVPyR2+B498lFuS4Ryu5a64zP+KKDwKR/DZoxAeyVPHwlV
LKBf8ceHyKXtVAB1MbtZbi0sf//M42Dfhw8d0Lma8AtWW+h3GcZP8i4p2yYjODuQwp2bsq08UWv4
9LUzlGeeT5AU66AuUmDqdfulXLruS0slQsrzgNR81df3bdp7RbC2ukAIAxcU4SM8+sWNVSHm3J12
CfOX7NPHOw0X/KBuPgWH9TePN/4bBOavWnAeo7kDg1v4xepEbSt6pO60IfYf/yzs2YB7FCONqRY2
EjFa+mcC+10EXjPcvp+kr0SUUlmqvtdGN+TPIC36DW43kQ3pN3tzxD/oJGsrAL9U1pDG4mEYwJoz
qaLKq9+zNnUxcDXmBQLjjERnHxeD7A25yUOKNeV3J+QMJCHVyJMmenZC43F+tecUg0qYp/r3PBG+
H03xh6/DB4D/PSmiqchd/k/Jzfvex+HhbrzjbwcBPU4rM/zkHCnfgnbRBS1UbMT3oCP/a4oOPnCh
/QizrAqJz4f2oQ9tcaNC0pSFKKjRE0ExeUaMc3gc5gLwuBEQ+GISGJFrZN8hn5gnHkKf8y0aGGgz
Hs+1vCcVvU6y9942vq6+15Ei8HAenjwsdiB4EiRxW09TSJltOfGnVRJT3TEiBb1e4yIgerQKTn+B
U1PyR0cK2pskR5zunKa8clv9jV7e8nLY/ut5zuS7zR+12rSCRN5kQuGNPX/yxlHtlqrAFkPNjNj0
tchiAffWNFpp5cHdQV0W50Z/h49N3xjHpnfYMIbj4of7EVBvosi271ds3kTXZb+cRHebLVyjbIIE
VuCAageuwt38ZlfkbLU6iuB5nPgwJIpg7QELJuTMMYB4FhANZDsHyud8iyFjfYrw7TIEWmoiCrNT
vHpS+VeyWbXvwPYwNQOuDDd2Smxtsnl1yTkqhoF5lO7RGd0WMzXF+iAcs/dVckYOSJNyFIt/KPov
M+MbfyZCv6h6W+XTutXiQnZUfVZcZUddGxPhbg8KiEBwDaUDbLB8ZZ/R+UcefM0z96fstRW/YbYy
PNqXxBz2/6FlPKQLS1sLPHG/rjFknOlYjCcgt1lxcbMYPYix7eL1mpQ2h80vR0m/XvBEC2NirFHw
wIkRbODkAonKNGPF/n9MD+eaLmAn5ub+2BAeplpVVppN6oQ4E+9TdgFhFju8f6PQpOA+SgFXLYr6
NtMSMyEPNAP7VqkkM6o+eEbYE9xjv291NsTl9Q7eOgrzK/AlZ7H4uhqviOYzxCxqYj+HYz1KfLof
sRSW79DWFB8clsSNagKeHRO5tPBdW/oshAN5TLbYm34MfAWS76kqUl2rd23aJYWwdBXLqoyeeQD0
76fIlr1P3OqzxnLE00mtR37/6dvuCn8Lutu5JzwLRdAZ5dQRo+071AKk04gPVYM+Mu0sKzALrMcz
FwhtWtL554eg75QKBkSVavltFtCDXJVbStU4VUdnPYF25wcD+vxVHPriQXs/qdc4SADgsbXLPXdW
DhEGZMlvMhQfXtOB0jMSOX91/bf2NUyASgz7JkmlajzRmw76RtkekVeCCGqw2+nryb8Q02Ago4aR
EtUhCi8dGyv33CpIaCJP6v56svaiRaKU1fToCITRvveuGsPYEa7DHv4FGRvVeke1FZOxTAFd8lhl
cKVdHnyrBUokpzctMutZgnfitfyAiolybAvMWo93009gS7tQ0JeduhwhNHh3jb95/NciG1HFO+K9
7jt/dLq+uf6y3lNNmvs1vgL0SB758D/ueUS7shy9BUoh/bFJDZLznpnumXGwG1jLX292TOoj7/A/
JagglQFNBGgBv79qHIbpMMc1X9QfpQgzU9+Eg8kHmaILLM/PLfEPd3SAOrSHSXI3B4Vz5VUa+AyY
Z/tzEGOWN6bL3GG+tiKsNAob+MTx8ETybSKxRGJ86L/Oqxj1CyEGbf4vLQXkfiuufDwRHKo9BIqU
0cgWQecwPHLMLVHUtil3VM5RCFaBJEOvoXkM6gjSiEF9HFvLVIhNBVojT3SLKuOykOEV6iBVZNT1
LBNqw/iIIdnt5KDSwtmFzYzJpzLtEI/Q7BDZkSp3GYuVQcpwiG6Fxuu115a79R57HN42HW3VODj3
vYn5Xdy4N7H5zenlE3D7SucK2+3jaH4ltY8fmdjB7VuMQ8GCilLHcDQEZM2TxmJtXxO+43RRXfXY
+hFOTMaLN8T0tsMCShk9xuZtlBumv/Q8FF/99Q6AGh2TsbXPqs4l7Z6wnMrdaNxbVHrWhH4595iZ
EcZc6ZO9asvuZTSvXGTWEMKc0sjUioj3Fpw+ptLJuhv1y2kTSNbe/BivXywrxRmmomCbJfjxKUYZ
SP9jf9e4RzM/osFH+SRTHVqmQEijFfChjpI/PL/Zqge7tFtkwbxB1dFHZdBi04TCU6MgY7xnaO9l
t4KuwIBxThetIeH5GqriRRl4RtY0uObikirFjSlrA79PYcg/eR7B/hlZTfF3xYMpOtwBHnZlUYj7
oNnt6frIitvScVoTxS5MmUDuViWXRDMNX4tZ5YrHcqDnEeT7dYP+/Bk92SJOe+ss8G8yy4pyXO6B
hopUb4JAAo78BMYp4CpAyxzImcghNnSB7TLKiK6JbqneUHbX+BYEht80onzrDoiJUhWuv6x4yjMa
3tFkmfx4UJWGUsW7JKs1bqaB7V/K/uzbMv42XTqo2GfotrGa4pmonqA67dnE4JDlBXJTdRSDMK1z
/l6evhio5bbkm/s3+qZQJWG9zV+LSCE+3tajMGZ62VQmzHPu6Br0GcL7Mmd/E9ATBMl63qaUy5iR
t42aok0o9+ouet6pfgpPSlmNY4ccYwpuD/xu1l9YtkE8UjACVGJjZfqVPseRrRjL0qXFXpab1MP2
X+O23yzQVPFvc1R2WbPgGuREVFKoCMHphmd7jk2x7d47KAA2wJjvrEFL4T0Kor//fvqxvbQ1M42t
BT+jubiCOwk3l+fRmf0os+paXlbbi3887PyqPTVq4Ts8RpQH2F7VctJL8r+SjNZ/ahRlMqrunMJY
Ar5ao2Os7z2pEO6rdUglvgTFAWxlh9D4tAvcQZlsL75AFOJBs2dMZme6B6U5dRJDiLeNuIcVcMmx
7agqk37GW++F/9HUBcR5NExBML8y0LkGq82n5yVsAXyhWbXIDxZTxW2Mdg9Wg0dEqBJk8Mv0pPSR
umjlH9v+ZD9IZRRsqnoBsavT98Alx+mBRUdmjyz36jXZEykGne0XnAELdPnwGP1vZsPJUcBqwq4W
cAk2AOST9IO6CZfKd7cw15EtVm5W04c4mPrhULrGdVl+hDEcuzhGOQ6l9fDqsQNDQztPVwG/4A9g
FMG/UO+kWQb4Q+jZdPHdNXp9af8rsIwN7br0dDOnrM2SQInEd37ybhjZc3EZbcZ+Hwh6h+zYlr1j
BVE4/VEiGNAGlOK8F0CaW8xKCPhm80DUF8MIp99FsRbSmUkxTmuKe1pINVkT0TZ2+l9Onr1crAz/
gm3TJ6H3L2yA5YI1h5dyRpLupl5JK4mIeppPOYl6inde98Vc8GqjJgnE+vD05ooPH7If7NZXPRFi
3u8Cd4XimN7X/j28dK0uremrM44OKbNJJ102NTAj2rY39f2dSAG9RiMDXHYZvxkq2xhxS5pwxOMf
CKW0iTjBlRz55t2Gxuouq924BmQtRNVytpucF4bz/vSqqOEy1uPBX62SF/WfpxKiVX2VqgiUhr5/
sJOi4FPf7h8USmF5RZc7rSOBj6CVVPDE/FZ4N6Hxd60updaySORTQeJp4QG2VyA/MZ+uRHM25eNp
WH8caY6SZI+ZgXo+PxclBZUxnlE1BwrMzF5snXaHupLcyx3d5hOyUst/l/0bo7gR6UroaI9MNebi
IXDq3pJXXxjWpt8lVy77fkDuem6PQYbjwFBleqHXQlY8NOdE4vmIS5oNReU5ttW1OEEuQYW55nix
l0E9rXNrf/F6xaoOlt0GllrtuuV98kDnHyh1C8ozNyFyzWYQQMu92NR2cHnz7VV6CSD7kA1JHOhT
m/wzTVMSxHUbdhbiLmrGTEkIHavJCt7p1GO2VhnoBMUg7fJCxBmq2CFJ0EfrSEUAEx3Q9BL6FIln
Rzjo+26hhUjS3hpg6uNQCdVnmXhxoe1gQP+4l9rf360xn8Lr8SxbB6OKHEUXcFy2N08pjb6OLso2
UuajAFdXRMKK8flhWAd2h5m/iY5FpmE6K2pY9CPmlF0vPf21ASbMspb7cFExwBKNISE/dCneYNhh
/OjSY08V6rFl53KD0sZoAvug/r0/b4H4TiXrf+rktfICdbysFqmB7wq008av/5mk41LZIgl0B5GT
VZhMIpmyIksbenC4utA6btei9oYxYwO34+w1MHlrV/IeM3BOHZYmgcRreCaKQdATIxNgyKraUIYG
LhGyWxki4ItUcoOPTRjtPmPy2/7qYPH0l3VQL05vc8i68z1cdoTj627rZLgUNg9f3R+xFT00+yX1
5iGc+/81oYzCDcBmXLxX7Cbz/cMmymQTtkBbuck7tz41lkoKK6NDhcf5oeREo1uJTVIUHShQj8Fz
7w09cAL1135h+cVtDzua1QHqMRbAbWDCvli1bxh17Cptqi3HRs1BgfTr1c6ySEPgqFgyY+dXw7FD
L4EljEZFPqPoV2TRhP/GOB6qPXw1Ujsz0iz53raeAax1uUposkLDRr9d7cYarNj7MeUb2E9ONwIG
mnG4m8vzvDJBhlxIcTZ7r6zPKNhMxKvxhrKmtpfljuM+Q6l53wbU1JdjjgauDR8AENrwJYmrWuXs
68HJIKiL2rMpxawmWLj63OOgaTOyup8K3E0t3FgESKj1IruHxtKQezjdr3A+dsyT1VpqdKkuHeVO
MgvcOfQtFNXSt1eXV/PQmfOj/xlTf+UVPXjzvREDKfTYLNVnGzXu0eisHaukX5m0y+WGEeec94tf
gtMKf26Ysvw0ZpaTOQFDFgngnPlphPujyxnnWE8IBaYPEc32rJShBOvwzDtg2BNK+XaacRuVWzls
x3uZr/opxcavXH0MVltI4sq2JIFrIHKN33ELIQtioRV2iWQVmBiakFhTBqMezJF6k0xQw0+mK2G3
DiaeJ1BTG5l4JOoWsw2iTOZ/dFW4odOw1GpP+/Ke/pJ86qH1dwtp0OXdiW+0fmq7YtgPe+jr2KHH
HYgssNDVubozHxvpkpdF1UBs2TCKb1XsLGXOdpG55D2HJnSgQrP3ogr2gC9yWPLQeuXYDKaUYd2N
do4LT5P7j5NJbgYLri7ljStJ/SG4+7YALyIO2IOUruiUsG7BOqV2T+9UbzAHlQrW8kQ2bU2+r2HK
j9RUiLVjN9IMpCDSNfCGeGT9mrBpw3xa9EmAeVsTCEF9mmoQ1mkdtjPNID7PSxAa6eNTs8Jolc21
AEnubSkZK1PdE2y+GakmmklHQdWr4XHv8UTmpD4pHARdjlGwfjt0W3jqRHlVNjUW0tEzV5fpuU45
hvqsjQ99mbVw9sKbwZPvDNfropupvPIVAUsJVXRuk8Kcans2sXhdXVDx8jZue/npT+zrB0Y+9iwv
A4jRz9NTGqczAuFI49JM8MZr4iW9nASsNdO73ZyFSeHAcy01vNDtC3nZwamwmGVKbn3DrEKzTWa8
NbrxUO64nMP3N65SNG0t/gYdbcHRp3c9d5Idfctr3uGyD/opH06Qf1/dvMjxyhwguGJMZ1Rtte3M
Zcw2oqToXa48Zb3sUySzA1WKHkE+/CDVh1xfblVu7c3B/H9R93L5ZSCfVw7D5SY5c3CsQOGvByIR
pfNoFwgcrh1YAse6Ut0bi3FC58+GTW0suDZdbe147IeQL6kO9UIac5vnXE9IffPEHIbj3Oy1HuTQ
lieqlPigVrpfxxc1co1wES2yOsaYU9Q+Y/ne2CD3mrkUUMwFQNDusANB11ZER8dADxorKnztjndh
cLiHaYyJbO6kwxwwFKP4uEnH3Hdd8JtsVIeVM41QeNdh/acXWhxlQ/nFr3PhAk9RegFqgXd3btIU
pPHijb8z2gTUKBys5DcbsEmt47rjptpxoQVp6G7HJ7qvuPl5H53rKOZWwropi2ao5R2wLFLoyN+I
Eunw0ygnWlixXvhUnV+37eqDPGMHeHITSlg5NN4mop1miD+aUIcBwSfHjzFy0/yVL5qqLdb1UyFg
zJzLa+z5uTqRy9wj4eG2r2H8C91PlyLcuNlxxYNZKyvnnpSrVr4uJ/qPpFEydO5Tg8Y65F78MffP
oY1SsrJzlsgJAZF3lYnIllAVJxDcv3FxbpxdICZUJiQJ3MMiWVBeqSunkKN4ZkWgkVxjZdFhhRbR
jO1EQICMkLbYw1MhyNmDJXFdER8+1OXeQTFWNRvYCk21UF19/hepj4/20b6tW8XO5VMTjvSeoO1g
wjMX/WfhI14vqlhAodbyEP8owj2h7JEjxLDqJ2c//4n1yoqk/GPMnF8t8hopp8JvWodqMpV5zk4v
GiABEFtXHl35d+Dq5ySqHkNwly7ma+XqQawixe59HBODejPe4La5zJ5x/eDegKTRkzRC3HseEtm2
G57z3/85nmA+E7340Hkjdfz2IwFvFtOLqXps6o5rsb2cS7inPBj0aJjwdBJA1WBcZSC8+1xP2z1p
+pS9N5SwcpCX143ngq4IUwB5j4vtiku062tLy+dLQ7caqHutlMOWgqgjL0VGbT4Qjp1BWkJxmvQA
ccVYUlRBWqwcpx8Ktyb+uUO0QNJg+RVj5uJ/q8bDQ4UOBHpYooubkWaQxz0+DHsjEGtyylqwxoL2
n7Km0p4A15Xqfsn9usoeHo5xsNOq+jzg90kk7jOI7enFEkcFuLXlF6f4yv8ID+JXXT7U3D4h8CZ5
3Oo5cEz1QMBxYWSraWh8TBG/Qmq2j0BSJ7DIhKk+hXhLUqBgz8GbZT8AK09pUm/BppsVqIOBnfb3
1UqMNPBfwL5b/sZ6ca2sKQ2pods92DG8M82vAtXecj2uW6KSswwhq1FR7N7s8syyDRtGvCQWOFd/
thZRydy1dkT0YnHhQ67LpR0ZJ3e3HfAOpPwxEoFdSIuC9yu3AeQVkRKpsfy25AvbCwyRNGKvNUlE
tY4DpZyyN4gLtUX1GRpiIicBUI7RdrSWDAUopnR6NR4TZdDVuikzau4b1glYiPdLgB4wf3ylSoft
IVrUv8cVEIMoiHzBrtm65BxyJxFs1mw0FkrzGwOhCqW8i7f5Rvoan6RwA9lW2ImhU41E2EmJ+kqx
Il7LpODiROkkSTxW2Et54dN1o28SBz94EyC1qVrWICqJAee5g/5ix02nay6HE6tmb4TYpd82uq/L
3UOre9jbtU1WlfmNf29CbH7/UcSPJH/YKURDVt4aRavSLKqpdCWK2soYvUUlL/UudQiWDrS1me+V
QJsYGDABvH8kXJ61LKDRDSxnjgxtFbvWLEbZjLYqRIkxibAr/LKJAlW2cz5EvAP+tqP5n28LH1ty
rFbtNoHUs0gZVi8RhYcnEu6ZtmvHgjrlzqEHe28IRJrxpa0hTUzlfpHdFWs91wYZqGct4JHyUHmN
cOZx2Xj5ezDyTw2M4mKKFHoCOHcI++rCpvZW6YMFmT8fKnQ4Q+rU5EL1TXTQ32N7jpgU7nYD2C/Q
5maoyDpwuv/Od/i92Yq1NcrcjOm00QcEmv2Q8k4jGzGoh3n+d4YsqY98YllqNvfOqlo7B+U8n9ng
lxmL0UFgBwQOuetXQRZbX7hYrU/P//mTUyjBS/f8zF844n6kw31HiuQxkNZMF3MDt+PhiKsOSyTF
WV79Jr/1fNKgyZ5swJ940IhUBZQ94S8PJQ+NwqUVh+be8orRDDPzlO6MYFAoIQGNYRolxQm26z8x
+d/nEHP920GykPy4PQXwzjFd3GYLD98fxhWVDV9Dyllp0opbj5g4K7V3QuzmWyljMVq2n4Vj3NXv
fJOsJVRnCS6I9ldq5nVvg8JWa5+soXRV2D56QZZa7ArJZx9Rk7nS3BjglzRKOeOxLBUzKZQNufiN
y3+IAUSLUYHe0tlMLrXnigygqkFuQQvOnwRnxQI3BDuEzpUtw9oxO9iLxVaJ9o+HMaiZjwtFaiaM
f9KxG6eDAYdMcoNnddo3IuSk9/q/XvqAnxr8t66Q5TfbiB2RT8x11JSftNBib95Ex2iKBLpgvQ2Z
K9nywK4rT+NVsX3GHpyEUU0+RzdiRbeeeoD/ToyhOBl/8chK10mqTRFrnH5HNGYcB7aZtTVUxw3O
gas89ADEm9ipT81WB7fAWVF9OK+LqntgXkwQ5z4G3cXYu2veLIusHXfbcZkju3HN2zy6307ZHpzS
DGPpVLDqUcVQhucTjND84Y0Ur3/RYFYRvfRRRjc7hTgW5fRMZUzrU+mIS+xa2rtm1uapJIvcC/Tv
5iUG99xQg8uAzlkuocx9x2C/HnJ1wiFngq/ybgy4e4xoi8duO0PG3Lc2svyfGnKe8FPa1BdnC8dX
UUUASNiNKRy/mAURML6z0DMLvVa5kGBMW9Gi+XpMm5gZaTCOwrGPtYkCQqcUb7l6G+KKRA5m0MbW
02vUV57tPiFDhAYNZ2orr4HUvtQGFz8MN9ld7NTs76FBvOydvvkzuAUMtcMqJlNgTdkcwKwYfbXR
yJ4hkquyJOQ/q8wp8H/J2fbmgtoIdotQ/KjJjlIbqe+BZesNM5M4iYgqhy7OmLM3c6edw5Z0/CaR
AZsCwSBEVU0++mV7FHsqO/+JBqFqZoNs36L1+/4mukK5SBYOX4CkbmNprxo9ChU60bsuUQZH3UKX
Oqf1jwgWtlNCb+L1diSPAQGUyFTBXlbtQuHlx8IqD/P+LFouxlGtkHzAwIlJnLUTFwX+drVTbFio
ScJhZdkJ/0JzXRbFP7OL6Q2seX4XeS3Gp8XAx9Nl2/s4TPAkhPMhTH0U04L1mPSJc+JyPFMHzOYE
FMOhmexmA0Ag3w8y3pAk+WSWiOTteBpHfDtAg4ZDuojZcJpDlQtkcjmh83HQHsX9Ff3M7uYauVjT
jK9ad8RRegQiBLC3aGXqzDh1sLY3tMhUgUDAnFNILcH/7FeDSgrAIMXU442GJDZ7n5mUgS3HkUFH
JlqbDBdhc+q1Fi9GREOKfOJJmhawHwUoICeL20oeU436BSsM6Dohno2R145giu68A2XhQAvToh5d
3shBZzHb2X6/3Yr0m3Ta62N25HUjnwkuYqHhjv+c8d46NK6Hx/4f8ocB6xF/9gAURcOfXoiQi4Nk
qQxfULF86PIB9g8rIdIB8KvNquVXhgTat63fRME3/MWgAa2sNJ82JroRkVM7QPmAgYJABQBJQIfB
gtD2MGjDtmJhX/V0+cz9SWYC/ufsXJKBKT1QTKBkPePRXsTEQk6toa8njecwp/5NkFVwLfgH659l
qETi9ysYqSoASvHJR7xtCt+UBf2zjtMtSekubsBRt2dVowOUHDm1ciJ5mZ8P+6gg9MVPSSkgwjWa
xmNJoBa4rRZqAIV+El3Pra3Qu9CkVW7ozs75wLNTB2i6OlTCosmahRq6ai5wx7xQ8uUJKchjxuC0
83nNOTAJ44AOWloXcJoaJw1ugINuLT/sUR7KZEsppYIiIvGU/GszzdIcFczU5romQaNlmgUKck1P
Vv3n4gDBGo5qpZjRoW7ATGBSsH0E56K6gvH2I41cbhl7/aXPAzoiVn6SpnxFPibuK0JKFp6NlVp0
/NftS8D1TDqwvCs1B8Om92RvSzk3pa27m90WvBlgnDNnXuLqfI36PjbwDHHDwJ08osR3ENHiZ76C
8ieZDp5i2HAqLcQXML6JLaMz9X0iHmqqo25UlrGW4UfPSq2Z1Us2O/wDARNOPaZOnkml+h/0SFce
bWFMU65eih1B5UVorus9sJQL5jYSB+wEh9Yw0RV3KsQ0gjb+nu63kLz0TWzmlG1yAMa4Nf1fXGVQ
OBZVUSDQRRqJuk5Ye+RZf3aUaM2RkO5Lj3WKVQgSJrJPcLLZ9e9YpbKkgXO/m581Sxbr1AecNSYx
EHiDfLcybLRGA2XRlXrvDdh86n3/DAmoL/nf/5SNMQpnZCRysALgzr1Cf53XodAenVtZoLNR1gqo
j0O0LVBTEANVpJhsACpjvWXZXsW55rjnZJZoASfqT1gPKoocr+X15NRureMHTiMEYtUHfsckEkKg
x3I8212f00MTHU+MvRIFyODbhn9H50y91GHH67uf3rXtpL/QyRiRkRZ5lTwEuxhM7Sl56ghEumfs
s9AwiSKxgX1RIyaWcxaiOKGASPztcflRzCWad/ICFOY5c6wqki6/QWKW2nT/WvNlKiBEKd6v8wFD
9EWlHwCprbKZBXwIxICJx+fKjmgxjWMNklIxeEzDyXxJYaNkAsfbYIBiVSpcIOLJ10/k1fWYGYe+
vpxjqLhVmfv4Hnhyj/SrX8saW/KU5S/+npZrUJQQmDNJG3tTD2V5TP+qNgdM9VxtrPFLSlpXSWN7
nRhy8f/eyzIQO7TY52+tVJC6WmZvSpjq0fC30mJAAbzO7rsQ/eaCWKOL46ioPaihXEQ4ILGZ95VT
O45FutupjGD0qZZXV2BlBJa3poctr8GinnmxzHpwG1wvEVg0Qy0A/OPsKfZ0cLtLzIlqapNch7LH
DX8BilrhqF+WMrXO0zLMuSWUpqksKuBiyLqm872eqTnqhU7uzFYfChBMeUoRZstcT/ipwBLJRTgb
lRLRNDZEYj92OLvmUufusdwNsHd0LYlrNK/iR7DkaCth6dItdgkMScYGeUmyvmwrSdqyx2FRki4C
VXlKX04Dbzw+fUaM15hc2q87iV+ksMRbsqHoK6PLireQ8E0o2smph+MtVODkzZ0e2TBE3X9YdVWj
4DdAYhhG+e8BO0Px4wJ67UPLUxKP4+foLICGhIq67TdRsRu6XqsbxLpU8jF4D++YG4NptBYaUKrV
72RRqS2GqqFUNZ1C2gw+RzNJIMXq/mx0NUTq8FXcl7nEhIrzJfFVzC+EeJwtd8vOxmK2cwEuwErJ
PJozcL+ii70s0Fsmt+qbVQqbFoID6/wCqArcgpJp/5dWgHz6sLe4bEontabaoBoq9GX8zo/6P7ST
tebGIDb+Gy58nAvNt7qHs4n6+47assnHy+3C/7ba4R5sOPW8Fy4iHbmmNCOe2wJrG/+Icf8btyS2
Gi61TlcOwfbf9vnV0AMZ2ouqQ1CoXCHwsxVafVP1GHn+Z4zpps1GONuBOagYIYjdlRkgNjfXduD+
eokqdJAkmR7M8gw6ntQP3WYD5Iu6GAJy1nR3wFCwsUvGplC2WXRtcJNTl7QaAsEy4qO4FQB88jaP
AN+0C4lub3b1TwjXW6xH1GdEGZNHG7Six6Hp8erxvevx+H2ZWZFimTSJ6n7jdcoi762b74W0Nh3g
8XlT1JHp1gqoUZFKkW+c9wSFUi4CW/5xlHOgmHP/dOF3FpsWiN9agf2fXDKXL8/eCMcJdtpS0eZd
tGONMo7uJmJlr40po2Q3SbRygPGlqLuLLvTrdPBpeCjv7GtTW5MCmQv7Furq2MAJz4rMtV1FxXrh
loNzyyVq5wnRjH/8gZQTdGYE93XpeqUa8IX0Nj/ksrQ1M8oHYRAgD7G5pWKIUF6Ld5X3dMFCcCcv
etfyLyHBhewZA1RwrCTv7OmbQZWemkjjLYJRUA03sJUiN0y3Y+a83vH3WE/Mq51uontwJw4kp2rz
mAfXNG5gns6SyH5jT0HIBRcIKp8NkO84A7hfSod2I3IKVGEajyRCcCe1ba8R6tnhR9apZSOt1eXs
G3LKw3fb7CY4v4CCj5FBCljw+bD8oU3mpORpSIy3PFemSWhPPg+84wPBQM7wLdlSCBkIza+tZyh5
od0j6NTmE18hOK51mG3DGQnPShCyRvBe/JdzRLzJNpXvCWVXvDTKIz+vS6JkIWvcPcLj22k0Y67M
KVGcMkDhh0vOQlF0Pbnbag2RbHO7hAg8Qn7w7eEr91KsM9f5sTYMMDkBVkQXZ2uMZTbjnmegMlXr
3dWgotQZl3M/iDY5EKmIx0Q74wSHF/MFhB8mJPQ1TsUlg92NVFmAFWzk37zF6ph9SiSQzH+8ZuhD
HQFlZTPLSobMX9lgI4yvNgTT9hHx+iIlhUJD/I3ncNbNu56dVPMtvnevmkJiKTQi15oD707zztMG
zto4A9jgefW7uIzKKW27T2K0l7Pkut2IWiE/JEfOnCvH0FZxGEBd4BtiZiEKPvndYJQBSBqsLN77
6+JmqXbKJqgRT+jTv8jw0CI6sztdwR8SVxEvqz+97E+UpEudNt4HNHWEt9f/muRXIABrTZFqfvk4
5I+YxLarRN9ibINSVLmSxSS0PiRDi+ZmX+HjAuWE7p37J1fEYxoZG+wRLhNsdy9zLlmLDPDkFQ1y
KzVeORIA7BpuuCMBdwCq9kOtuF37qdOV/5/xQhNg6j8V/10W8L5+Mono04LGUnoad1fURhHzuFBU
N47+WAOwjbzwX2NnBa+NHG/KTUpH0AbBCtKVgYlxYLx69Y314I/Etx8GZl/p4Q15zZR7T0DG1C1h
yUyr9jpceVfDvR+oZ7PIiZ84/EMvIm+N743EqFLoNKHTA6gamB67YAfrW37Q+QECp7DlbAtVY6q+
/rwKFAAsXVhV2nd0QOyK9QqrNTvOOvozlMseiDphihWnLn5ggZO9gjjWHIEVRwRQ7WN+okdB0qGW
Qr1+UWeYnhefKvaC95x6v1JoDA/jA6Bn1IjwoZSPqbc1uHcHeoo1QrL2BY22VJ9nujZ6la56Ry6C
UvWlqF+KEjt7u/zq7cRdOOvpKwGvDexJIh4M4dsTYoNtcD2yOGGSlQsj8aTfoCydSSYnEwpFThwy
sSujMLg8wH2PVXijBy4XAvK1bNZ4OSNCDb7X6uYDi/g7y2cUG2RKay4SYEfjp1MzxjMaUvAtEwbD
tQn3Ic5j3+3wW84HY9rr/dIjeladwChh5x4EI2dDfiI87YJo/6i8goFPVv+UvRTkjoiNKw3FFUaR
R8OKbHybHt4S5Bl1P4le+35ALgWvgeesF4dl/7M746wKQXSuJ8zi6jJabxKPOvW724bJEOxoncn6
E3jOmZdqduspwraWzjdwLiOsOz0mrjJbQxwNjRLIblu9DpXGdtsdhh/TbXhSSR2F59QYpPSyyIsT
lxY6MQ5m+C6Sa/VaaTTy9xcWou1aKVGBHn/PGB69tvrOd2zmP1UzCUf9+dGRn4y7OWPsvmYVqi9y
MhwkPHo1T8SICRKPARkjOePlowqbdUIW08cLQQbGfIyyIOAtniaAXIjrV3YxXSx9AfK8S+7zxlis
ECSYOjEyjTVJPnH0+2QzoPY594VFoUp2/xL/PVrVXX4ok+mFbv9Wn44uuSwIAHAKN2/HY3anMk0x
xE029BgrtGZP/AkN3+hsqnH53FGXXsq7Jpm9Xh02K7RTQdhpqr18LDIQ3J7wZdt88W8paPl7w9t2
k/MFboIhPVd8pBgCefzXXvKpLxFs+ZERX3/bJCa+Q7vgSN5ZcjL8FXTRgOB0V3rI9gnMEB4iJJNP
4Bg6TC4PfT+hy4Dofegzk/eP4S/BzDdhyjKSBEOR0a9I/8GrG0ctrsSLAG0+kEVmNXy1lk6bCawW
SvN3RlJcVeKFsuGQV3sBTEyNlpxLWlPkc3PD+B3Slng+5UL2zw0VPhX3OyL+GIvIdN1VJd6YMRZ4
+SYH3YO/o/55JX6NagX7QUv7xL4heZNGHM4O34daRWpYWRuXeWor39eh5McPTl1sQplTBhkVObi0
iuIw13tC1Mfa9T6hSMqbEQqSLNPXw/okw8Rw+4aqkWy/VveRou2t1joEtS7YZlxoYwo2edBGp4N7
2vhEHZG3gTZqfAIpHl1xj/zqXREW9c3Ae8NPYLigKgBxkjSWe2ed/XnnU4W321SJidVw7J9KgpiD
BKrn7elhX4X1PX3IIrHLAN5kFymKz1C1/ecvadrRzgTl4IpQtGtOEUqf3kNYe+ZQ1hniwdHUhCJI
04fSwVPy5CwIhB9gfIjz7ZgUAmKUM2Qkpb8CBIWoIfoqbpfyemyl/fPROoYKV/IQgdlGAIZpmWjb
/Ryviir9JgMtbDuABDXx01BQIV754UiTczZoc0IvGZWvom2Zi+uCQOG2Z9C/neTS2qV8z5LFjVuI
mfUxFvQfLOQfjOgkemUion0r73wQ1MIU+vroXatmQZaKVa0jsHh6J1SBs71Z12K6OFPkpxmCYoE/
BPIKlMFUEH1voexFOWhvvDdOM20yntQV5kUOBmSuxkR+U6TB+meUddUK7MKsFNrZlpq6GXyl/cik
GKjtGxdkOb9SCU6sujpsRoiYvAYtJfuXVTyJhN0GtfJ6B7uelzxha8TGyVRGiG1loL0r07vsQ+GR
eezMM24zxZsRhP+bIvLs7S0i2+oGfYXGOMZxhX6ojNiDb/XkUC4q0VrNBWicW5V15EyDA1uiO/zC
OLUK+g9TPjOJ3S4Ow43IFBdN5Ms6F/QaQ3jXCScf8mbPXf3qD+STjph2SMTZHhr3qBnMbu8h5amk
5n5Z387j7gyzRDQHsw2TKus7B/RSW9ODCCrF9T4CfnIgdWjDpftU6mac1FFNC/kocYhlWYk8+Nh4
9FvA/r6jMhfnn9XoZAqcBYJCDQsAAfMowdmCCsqWSdF/k39LDUfb4jJHne6iQwWwTtaPLxjE0Tw/
av5OT28V5mWzF9FO55x7uCBHgjDhYtDrcgjTNN28ZADGrPZGns9wZMnzx6WzslGOiveNrukujWX9
hKjsiGGgflgsbrjLEfZBtp9UQQ0PbKRlm1/fG7xP+83o/OIQIHpad3967PgODHk/RmqI/BEXSs47
hmadVliaeGV/1fD/6CMlUyMbBxS6kCp0gbf6WRn8++4K8UFlN9JlxnK3utbP/uvxL81ScvXfi4Hz
7peezfBWl2LKMXfnRJUuhV7djo8nqxiz6byfF34ZsmzD3MHZdkukd3kTUzke+ImtZiW4Es6cN4iZ
jCNvndLMzLXKw4ShEgPBZtN3W/+FfJeGAbngOswsKZZMYvw7vAyWu7OWZm5dWyV4wFT3O9rtgrtf
rMTkxFOWiJZC+jaWytnMOv7Vt4w7aHSe7jMx/0WBJySeydTClM2Tvu8W3jOliQIhcNnCrhe76maW
2/Y4syXQi/VfC/RDCfnLQMOgt9sqFBY6n/7SQ/MZiolUdgcNipe3FplgZESCsuQqcHQgWpnm0aLg
qliC/4uISqnXunV8ZuCIWXPi7o8Nta3RucKS0lQAwDglTu7P8O+4LfL4xIAopxXYMSJc/hwVcD+x
RZv0/D16QGcu0w2Uh/+5BlRenSo06H43/kzcoDM1jAVDnyDq1So+QG1bVoA1r7IIQ/h8Q4E5M2Qc
0P8e/P6rfDYTsJL7XeE1CTCCi2uKThhyh4tfZ8fLe9OMvJ93+X/d2S9zfRv7t4YqHdIbOGueKBGQ
STv4JptuWYMwTGJZDGYcRR+4GUAJvRSQQV3GndQrYL8x4YdrqtTy7OM3pQiLPidqRG6g8twTns/h
YEiqzhaSvuAks5NlNRmoopVkDt3xyN3PE/gxPA+zn6h4TMUDWhP1RPanpfTchHVaf2FbjOH/Q3ah
p9fFwrQrxSSHeNXs1P7D3ZOQJp1a8Q/4dKqkZu5PIrQolBsThf0tEi7I/w2I4/ThFAwMM35gb267
KjIKL7jfGycfonZv6vYRjgdCTc+VTfTzXKqPUWiYEJbZ9geeMUQRChPfpPInlOvTUV8ubGo+9yxP
1sewDcnQIbsUr0FZMvKxr5Z39BBjGV++ItD9hOHnvGxi9SjURoRa37YGDWFYtEEhhqEPegf05P9y
QRlKbnPoyl866QbQCSBZ2v9WIhzcFEr1DnazjOs8mCwTlFg3vX/vCf1vQg4C9LBw3gGP0DKhN/Iy
T6zUaI8Kdgzp7RQy29VW91dJD6am9UfDnUP1eg48VPgfxiaQ2uwkveib5HmF/+KOBNlZzTCHHGDL
D5KRcYFB8Qd4LQP2muoxi9YE5oTSpxn9K99b0vSZ/MkyY8d2JuFd3fhulQFe7ld+iMQEMiQuuOpp
uqmKCyJqG4hP84H3H8fwFrinsqQq2EUbwmz+hmchFtQqab8dZP5WAlAZSvX8XKBIQ7ZNkgI4m8HM
LwGglW3cNgJzdZuI0KcoBllsa/p+1/bFcvAS3JxRMOcwYmzZKsFsD5wnBQpKkioNqaUDDWj93PNI
yb994Pqri0wMpJIPcjbMLdPFsdLIa/517Vf9D8/hqbN0VfRWsfwiJhHPL9yxPgB0NYkoZwoNePuX
V6wuZ8X3ZdBz9R8aguUlSiNJ7tifx9HdWS9+Q7AhPBo5XaFJqLWZcYb/BHN2dd2+hR0Za9OxJX5S
Ff20q31iZpMJFNTnYGQcNQg2hz7H5nLCqP4erMZ8g2YkbqC9eYgudEDJpw5bSrxkqVy4hUMH+Akj
GYOuIuSr4O0igkC8qBl3t389z2cAq9+sAk2hWp/f/dN6dVfCgEbXfHmpwAoOw8hixdIFrgsC906H
8VA4BP6KSCeSanhXZST53HsWFT5ps1j7pbl1gVn6+lCrtHX/6ouS10IDx0fSjgl7KgLdmgxQ2wWL
Ni2UbmY1NbaWTGhCVRPzLbtDTupHX0a923+K2YtmBcAMb/6vRJQZ8FwjirC6+HIHLP4Lzm75SleX
KLN8GnRnNJpMcZsFq4Z0mUp3kaKBEq3K4IkMxeJg0tHVA8riDw47/arWJhl3pt81o2nWo0Doe0wi
2MzJg3vFz3qwHBZYLNvyOikyqD5p2m9ninr033wjfJKvMRo9X+S3NjF+tA99QUj5y/VD92yezq92
zeiqtJtZzfceNTC7wcgf7FGpKe1mYu6cBZGWKZ2nJFfsY200d3FvUvn8NOdustTgG0quYhg8J1u8
0dhUCwoxYmXrcGBb51hQ99C1Q1B8EZNHKa/GQ/Ym1fDhTlJLy9jLZ4z1ofSuJ7ZlXeHY/vVtZIlp
j0aCzJq5zNEmIENIul9LxKEgIoEEa7ubXokdkFyxhisryuIN4X1MBg5GHff6CaxtUz6MXz8bsqPg
8BRV/UHibvAGGbsAaKbAXndknwAXCdC5XsDhYT0PIPqUN8+gbZafJlQfqI4GLUa2dua8b8K6vxu7
liSkdfRJL1PZAFcgPob58PmbchvEu09PuGrIZQussUR2Bf8p8l38XDooq6tS15MWCoUSFIWuGMn3
+iU0SCtwI4eBeqDhxYClexVFCF4+KhSaOC/v+WF7ECqY+/d5wKX8UaAhbh9kzf4D1i4Cfxs/oOp0
UwMVqAgJC2EC+PWJvaTZwfil5lAaECZ73hodaHFAiv7DN7/iTLKeio8UmgtFM2pH5T8pzR4mjnAv
kw3ZhswjqywZcoHEjXZalvfoCjxMGhRs4j3s9tVXnpmcds9DKeF9acR1o8UMuLTaA38S5cJePDtW
vMoGddemmhNknGsFnpfxHPiufuNwOgOdZkXq74ilsl94VQHiirLc2vSlbuSDLIWZjxq0ea0Px5Ld
FNlnxI6bAuLkohnOfDD7MoHAiSSw73TSlny9tE8ZmNFtL0j2KAVwFTYB3BDwJNoyZiFGsWyleOAJ
IXRy3yKxj9I4mWDblTV0rNzkJWjUahUZ+ao/xUy59OgbXzIGHMWFaSVilGvXKTBbGt2BCWa7J/lz
I2B2+u6l5bKvTV4AB2OA2uO/rgmuDka1MnHZvJ/aLR5skJ8ESWiWp07qZbNX2+H7Tg5hJ9GGlIY/
PRM2bKX6PIdmu3Kx5uKkQxgPSW9KBI05794KkaNSa4UWy2vOwKf7LPqH6R32OCNKM6J0GO2WfBCA
Fxj8I2PEIF2Fh/oYddCrR1dslSnlhKL6tX0ZbS+xILIwnZBx4L7xxALjOzumbfgR7ZnrjXUrzGPd
9Guy/0V3h0xSyYOI1SwRFKtXDBxHF+fPx5xzlyoZcipTBcFEjtcAvsot5wPbnrcBpqzTOkWt7x3a
O9i+qnNF/17u2kzP0sxK4xZS2ylGsmj7aIaOvn7ZTJaokMXAbH/qXZso3G1SWSLrCp81Aw6UhcXg
MBxhiohmTwhFWw/rnSe7pJ7YKfPD7x4dmCnkOqSBwMLkiPqpK/0W+NJG7kJxZsfFNkSY5r2i6BIy
fkWy4QBcsFrRBFZNN7Neydd+/i7DRFtI2mHE2qe6k4TxMEcBZmsq2jmOIIXCr9PG0zir9c3tZaWM
Wo6fwO9CCOd+eDExvuEFih8YjyDyH+PjHzBYm4Kw6XPmmGmoivGKDbXGVaIUoO96nqg5rBI+UIYo
ASd+vCvHtM9pp6TFcqA3dqHo1l1BXoRd+CJ0J40ZmyEtqwEW0HvlK4j7MC9xt58nm1PuM2Nf4z9Y
+3knB44p4K7im+rxjPvNHqOYjOgZ+1Itz9dm1EamS4fXoev1FF60NV9RKacgFGCFSq6V4z2R4XuC
1yiNCuhZcqx3MLm+Ehi9fzTSB1o8ak0iq1cgwOtKhNPhqaSj9JWDv/CFTHAKwE2QnhPkNFNs3XUO
UWVzFy/9hWtmp0+kMxfDfdOHB8m5YvqrlFdZaL+tk859IcvRr0QY0+rn1Z2YoVKwG6z+nlo4nyZU
wPgjNGfsncczV5pivzBlARtJjTSQjDK17mND9r0U1e9HtwIBupqwCxby0BXr2HlCnCpXDS2RtO9d
xJ30QuMUPkoYrzaHl79Ovl1nYnunh2s9L8+Zu/ZNBs2lCawiuThwb8DY3QTw5uQH/0EV0/eRibct
+Uj8b/CJ+3qujVh8FxfQ4kZp0U3AhswZ3erZeegaOaw+NNUlBHAzCpTOygWwDfBmGo7g6sPIgTx7
ZTjXGtQ8tLd/LerOkF3pllD/sNx0lAbNtDySlEN1hBfdqTndxgkt3xd3KWY9f2T31hCLCpLgyFLE
e8yOIoo7L1ukioSQNPW/ByveoynykG7E9SXsYiOj8knJuhDMqhmYFxfFnRNFQzjRAbSnaGHTZ+my
zAHpG+4hV2clX2zMqWkE4IiUg5djWeGV4kRj6zka42haLVTeUZrR1Pxr9UCSKQFM6GDoTkc776eP
2emdBWr6T/iKwVWh5BTAnzOYNtt7XLuCN8LISENAw3Ts37Bi5rVw775UDwT4qkjYfcctuzTa0j+V
QzXzPe4GB7+GNndnOsBR2YmnAF8c+k4pym3T9ewU78wXEBPFBvQsw90hLhUB+gU2Jbl4IdJVrp7a
dwY58f0DAgHvtQrjiH0gWtMIKhKX/wEh55s19NW/ajS/p+r8b8chw95CUhgddWSa5DNIbAbtOHE6
D3+ga1Pm/fCpseglbKA/40aBejhHbYQ3LfHTZOJ7OE3yx/Ohi/PRdhEWEXCz5pXT0ITJNyHHURq1
jVexmzukitHL+sNfcqbHh+2K5Spl45A0FoNBC3pf4XYqClkw9D4+o/iZA4FoVbSm/a1aMURij7DM
apwLDIuuYGtmQqOv9CN2PlIdkwD6wPzXl6r0cehuv/i5MXzeKXP3rnKwBjXuFF3oPxppawSNDbW2
usXZfkOu0MQ1g5kv3FMp6qnfoSegvDRgHCQ3C0tCk393tdK0RlKFFe+7Sh5c90vRokWWpqG9PlKL
guW837FIWcsvvxlRgUUdpIYP5OO+JuLr+PvlvSL6PtZtF3QO4k9vOFG7FBYKOsudivKeA73Dxi78
CNuxWSbetk9f4iJct+kXuImgNNefJ8/zVHhA9AmvKjFLzw6rKv2nZ0f1doITgP2FTzEQ8xZAWpWT
p1/W4XFDDptjxuDj0Vq+ZxyOZkrG3KodZRTIUBI3Ulf6Qer6ekJTdkDJErGWyjeCW6IpLeJohYJk
DAPjTN0SDjEq4igx376WzuiCt0ZTdPi/x/6PdLRSpWGykl5HSOTSgshJyDcEXWzEleh5g9h03+UB
QZlo6vJoSg6Q8FGxElwgUE34jtjCeR2fvOQkPI/lA5Sn/qOSJlbRUHQvraXNDc0x7JXqQEdFHLml
KSxpBV7/4sFjcDw8MtFZRunOe+vaNo06dDqHYb47P0c1Bqa0aWjq0E233Yzq7FYU3yEhid5cd6H9
v6A5EiLTWPV1+ob3UEluVtPo3jD6mHPKVVwh8/K1LTrpyerIh86ynlHVAJsglC8GYbOzMdvjSzbq
MTXjeg32jxMAnZApHo2S+PVXpCPR+VCfZwN2rNI7W/duhrQ2znc8isz3vrk3rX5xOF+XNAacBoaJ
g58zNq4coj0YWKcdW+9ZlX6ndtSu/FjxTddU5tXhP8RCVHizG8rIetc1Lj745OWusHxQ9Fohb8sT
HcQzpc0+f2NUkLcCC0tJhbkXTkh6/3tbPOPQUVVgC3WCtq0jsNHARlbOKGdJub5MU38KfhDrH8pP
y1ZkX6/Btf02naq+Ypt8UMTNDRCcbgpn7T5J5J5D7JfuVZxtqJaYHMcQll8Cra/lUAr9h7l4s3HE
AyuvcE+8Nkw12qUHjdF53yN68ZJzGl7YzSrbS56NNkMTn8Ha1M4VBAylI45YZRc+aiTfkjyjC0rU
J18C887NfwgaXCdf4YbTCW4TehVg+2fEMr+6kCcRmh0yTW/V5FV/hUGlOUp/4bvpF11z0vBdfuQz
1+2YV3Yh1jxpIvjuPUBTWjpPQNvHzgkToBSh6MvU6KZgacq6vrmkekP262k7uiokCkCxVG7w6Ry+
WdWehnmdBnhALkU5tVy1PuN29+RAXgW6SHL70BF3ZYFxMvi/f/UND51GNv4N8zM/PyBCSaTQdeah
8lY/v1ELFsw6lOaYB5OJ91n3FwmhN+j8Q62QH3ht8nGlm+HIfUjVWlRHAm53TSsFoRbXUeUVpRZi
WoLvo6GMgPEFNF3qO37Cm/EP2PBRBDF9kJkpBxpdYGPIX5BwokJL9OAJDb1ucdlabMUXz92l0YT2
R7OK+dJWVTfquYBFkgA67Lf2JO/NcS3rJGoLaG9R1oNN9xewK3qH60ICgJZkD3f0vBLiWU8O4E4G
fHOwV4KrD1+Job36gpcw5scbJ2QERdGgboUvYdEr0zomgddSRGvf5sMUEqd1RnYYiH7pePvfNqYo
LTClvMKGRR+Li07JNotuQ5LeBBjTHTGpriVh9Jk+A8u2bYj8fFDOg3i0AtMW5F5S8xGBbPoPlwku
f6okpuEPpfgOcnOVxsbhIx3iCqTL4BtC9hjIbc5s9ZN6SMOZnqsriJMiNaKn+Wta2uhfQ6sBxgG7
yxicRh5ZcnbRuCGNJDdPmtKgolDja1onrLLPswCP+vYxMNUgNyenU3vm7d+o2sUroL+4ooc8nQ9F
X4FZCk9/UpIAKCXzxcemeElkXsupzWo/CFYIeIRAELlbL0WvblYavEsKN+tkgYNnjN7dpv717xfg
IZPby5x2IW+uwtORaTZLg/02lMpO1S8iUt87gAwkksbvMfc/eFQk1y14v9wehcyQO5O692s4SRBS
ZOTfYNiB1CGgteqmHiB74YEQiRjp03LNQpdlzcX6J9725W24NcTaPAlXGl+yCpz1X7QOEQkgh0qQ
z2htdnkppJaQgSKh/7Gyj9LfGcLLI7xZFKYix5SmwgNilbPWe0wCTnccQwIbO5yMt7rbXCRp1ZHD
8HAAfsxKSH4bu958xWxOm6VT+sOKDVOAlYjcmWL+o4LlkYj0qu7PblEQaRXY3IoCHIG39lD9F+CC
Y7tuE8+EsRU6buZzgsOyAh0OnyVTFwO2HSgRjnrTIx2LRDOOYLDrUO8cMIJxnRXq7+tqx47usyW7
S2F8g5QoUOiKyzv7TVVoLYHc3vLraTVFVGC7dumZbS0pJ1e3gAhocoIdryQyzECbwTCV4LzV0c7P
pNNoHlw+AbM+eUEVKzVYkmUQ1tQXjVYgQeul/3rNvbeQwjawRaAogWSQiDRDKU7ah4DCW+Nx8hHQ
j57eMu+2dR4G6nvS03fzLxAZnChTdlzhTCFS0v+szyUk0kGPI4TBBCIXTo+MgrOSlG45lVyMeBrV
hHdoWpNkVOwh2Q5fKqaxuqgDL2ukDD2czBPrsyMPfmkrY38S940k2v5/0E4d5Mgo8ZbvkwwmAjIg
8mugakkQnKRZRpJ8SuajJWNDiviN++TxV5kUU0HFZfaLzpan4VHzATNE53WRWur9nixyQ2hdC1Hw
rP3wrKj9i0fYMknVuat9RTazAab3jo8F9Pi9N5lgU7x33AaqUHQCnKSJzvJhZNzDNqFGILBQGz+w
edqIKdJ6Bxo7bu3NFGVRQ/IwAYt/gcyssvXcaEh2d1Sosr55jAZTFP2nSQYHH0LaKj4QMP0b6O0A
zP9AFmUHOVTLzgMDTzGXCrpMI3wD8G3gcPnIvXVhelhOKbqHto3trzrrPqs0lC2k9aPj5oI1Weyt
6gOTNDcPed/kyd8VK8FIgQ8IyUEAO1vJIHzWbrkfStIRxMXSP9y0y9JC1OLZ38qQnJO7KZUVqN/p
8P/mjNmzzQnax5EGksw34Qg4XNSo5+ydLydlA4qx8R5pvCfPMVCC5bgEyh5CSi3peR+zhOKpWhWj
IgQmt0VZI5lTYbJnkpV6RgCxfHo32f1/uuPML8cNAFxOE/qdPNWomyqzY2uxsxp5DntLp9ibfVQL
yCfS+bMX3HrLQWnpmFQsBpUOLV2In6UT56O4iFqH/eUDpqvSDCdcOhheA31Zi/8dkbsJWVfBQad1
GqYOD/V5oOmZq+Dys71h4D+3mSrnlhllQzN4S9uQLcDVFxGOUFRerQDxxlnMpmQyPl8GRG0AtUYs
BRSd3BbTeXNQu4ghseWVZ/15MVhVyB8ji2bE+EtPU+qIhxw4cLGnCE2dG3UWKZq8CAq/sL7gRfYc
wQyNmYdRdUaddh+gyOoHEzujkx6S+mcTdjHHG7EqSFubLlAy6uBLQS6OIp7pEBIzBp/IazLDMDr/
QH07aH2eDGvaAOB6XysKPN3Ya2qvxMNPUlXTBzAeUgJ4GldJwkTBk548T5Sk304sJrryAYzKM4v4
qTXB16h7+bMDnbjHE+f6tLB8L4uvN9w14UQROCd76o3NvwhaieJlOGrKIRoJl1VuhXk+AVX+ysCW
4UUN4bK+2+jjAyQUJ6O1L9HHKW7HpjE8Bfmf3ExtXGlLCc5RZwzQFEYD0KgMADVfsbAEHFn5I20Q
pwwqiDzJJ3WMt/2dzWmZGkeJS130x0TUV72ABOUzxJvQkvzDAaBAs93TJezve68Vh9X5fYAiSS70
XvqdTr83XFU4EO5aqYu1/stIZqoVXgCoz5KNZ5ctRmfeiH9t0P9oTa8Zw6pmpPPDJ+Tj8k7cBaau
kEMm/r4U+UEeVClnlh56ZbPFKP5rS1A27ggrR1mUGsvga/M5mP2p11f3jOpL/Tz+3xDPNJBeQJnb
QLh2X0NcrRXy5FN6SwmmU7ShTb0tqEjAjcR2+Fx1rE3LrXmXu60hWoPlYJMUcolOgIVWSHWwukpt
mARU9yeKevk0UxvWC00equo5iItpOZDtm7hk8rXk7IKj/ng1Pg76nKta8tZxhWHvue7FUCKCozYK
xGO4eWtkI5SNdR40n4bf6FVUEnQLFupJs6dbfZuDa2hEJrO1hwmXPu2I+48AXP+YZxO77q4pMK0z
9ByDyZfUpeo7cs5APKr7CcHuS+hm9DTkJ7CDQI2rZ6Wy5sPqrlKdAoFjx/7wh8rlfTOmGlCL7BDx
jHrCLJrJSbr0dAIXTEWUawIXbCbAYOt01p3y4kpmSIZNLuHHzXiIoG7oilqGoB6jruZKTyGuxUn8
rOjL5QIGPREH8n0Vj+zRbV42BI/+S2bquIuO+huQ20i/Ohgzra9HXFpJyShg/8Vu2su4xD63lDJW
kZJEatZg9QKP6Aroz3pirlXwtGAbSQClz7UoKnrzWTcIYK/LHdIIQFdhqPhIl5G8dp599661JFIF
SDomRBYFqLzHl19doN1cGAcPHAVwipyAgJwyrKahlGT6KG8GWoMsuP8R54aVgfR89aiTCHQGX8SZ
6QvP4ZtJIPX7su5YVIsfOSEo1hbPA5Sqqkzxan67+3RpOTa4vRZ6FPbpPh/mBcnuN+cO5sTxdB94
fZug1MYgG1rnhwDlr7DW9qPO1RmGpGMm8QjwusROjcdSsglIbOppWFN7qE70yueb2Q5qaX8NOoRy
s6VXprbwu3zclPY9Bx2KJjmc3O15TjEtHD1uNy+o1Y2Wo9jxW7Uv7PY8gwt5yURlvXsYDNBaxEFR
Ysc3MuIgwU+JxaEgmQFB6JQwBeDR2LMh/nCToDPhoPucTA3CqwYrvQl/vgBfeJqNoONtvYI1J+Mn
+0PgYxofzu9YkTMBNCqk4m8+vvqF+ugYrqeOEXvj0vYQdAzhq/pf4D7KFZeMU8rdFdv3hsJnhAk7
k+8q2Laz+8JUfxg46G/iw0mPJ7dMF4dWUVxaVnGqwTyA0o1cgsj2MKyRKoa2rOOikkSvvowoUjzV
E3DFovhdaczwb/Kj4QwucMbggqtoxn5Ldkm0E0bZQ0YTxNP4fyKqBnvBYZZoI+uijKhHAR1s5O75
bgmMj5J9YtJRu2fNqftYt6+xDTk1mAoLh0xuwHoHxxNX7IMBJGrKxc17fswF0RSJh/0Q/m2akajw
1KaS2pme4bYORNKS82HnwMvxpL6WM/VQ0zFLiEHFTIFIq6rvtRAlcyk2Nb/wtgHyPx+so09ksVmf
gIaYorvYa82xKKaUuQtK6+rm1rqv82L/2UGzaO1MPXyT1Ye8Gp/Yyb3C/FEKo1vqqbYyl19H1OUI
ZM4anHSsv5eAZ7wFmpBM6CULLy86qOU+I7LPivtJt1jgrtE/mXVMVzCuoXKENRwITigIGux6Dxn2
Srjt2cPPJxOnFryIOebgvhFFU6JYjYo0kRlkY17ILaCb56fV2bBlEiEiw+81UaCGv5WTJzee70AJ
xOJf0vplcmuG5pRchToGIR+ICPwq0AS/qqc0I9rcqFGuMay43Oe4L8TtNNA/J/UsCw3mbLKO2EY3
EJJFEAlRIzilO+NEIKCEwOZibEVuOP4CcdrsWuD1WWuO9mkTxj3b/Y33Et+BgQsfXVL6ebC/C77g
/sala3e0KhTHLrxhTRnhNSk5ZlcgvuQtDMDB1Ztqxl+31rA59ESuDHEkc8otboSNF87zeIvVznAX
OF02nFwA9/7ySnC5GaOIvg/00XO4zxWqTmyQx3GXLU2Ka/UeTNaY6/B2TrEXDZuSXzDrxw5QDhY/
ScGIqRvBX9nmlXVWOLDuD0Fo6pP65FNdOW/8K9zXssLtBzsT/zwbuuL84/tOrmfhrC4qKxTMMB83
sc4eVX34BoS5t6gXVThizMGlZ/v/58hwKU2uWLtNxx2w2fRFtOVT7/K3F2UIh6JmkSvBwoyLzim2
DiHuF/+4HYEP4Rlx9wS8L+FHo6S5BZBwZ0yj6lElZQWxipCkNey9OLlX0Jtx4Qy2LVLfKnYqelpf
lVbqZR1lzhbZyUOr2P7o02S/x6HAqX1niSuhgs6S8KgTbBsZGGORf6aGTSCD4eVvbnvDJK4AZpl+
GKZ/IbU/yQa457fjJcOwn14eptSMkv9xcOlJVmlOhcIajv12Zc0QYPldaEEEJa2nTxFdbQ6HJPFP
oAleQewVoSyd539hMeAJ9yqzoK7bru7FIKWRbYhOlCedQA0WnyAVkqnfu2Qn692ybivzaGVOFxEK
21vuWkIoer/x3kA7D0lQ5OjKxZiFQIvFCaDbYRMuBGCpLQdotKIRAmftsZR2mSyb5ojIhJPhwqBA
/0X1jIWBWCiW3zgvEDh2drtBsc1Zuxd8wjxI6iETSX15XeUYA8r6DcmAkwZBAh3eqOXEhVy+I6Wa
uKWm1wsq/rD9ZQCs4pV7dxzmoLv0GBF0OneO+92G0zgtETnNki29i79zRRP4C/kdYWb5BBgwMRqT
E6Y20k+7+DDgLM03iZz69WhJnRkF3E/lQzMp692WKOuV62oVFR4DxX7qDE7ka2hojNW4RV0t4Y73
p+oUYyYNgoecMS7Gi55/kRZom0E/3syLIZTTEklWHDdAfUVKwNc8X7Lw0vC3hzQoQKxFqcKjT+Gg
sTgAeUoQ+WWTi4N+w6mqX6/bXNBzUXtDwj3lNfMcYI6eTMq+G62VUQqnBh4aRXGx7lumpvRojNz/
1puZok9C1RxBET1H9niQGFffO/FKXgRixl8BfbGjdyHRKqAGBh/BI7NfN1Qh7BbiGhl8PPmS8jaU
9zMOkVI3qyyixGjMCxEeEzOZtyAURTl1UEZTwqUXOInq3lyxBiesIFVoyJvi27u+35B8GOAWGike
Y33G8lVwE6xEegh6saGxUqBNXHGuKBTbc3psxct/swntEBSXl2mp6bi1AvvXNJXNDNoIIdHi8Uiu
COLIJ4fXL/F3NxUiCjf7k69NpJAsZQfp4tsutRXrbVZGDtUCS5QBfh3k4m9EBL18B6nTHUnpys9b
ED6VFEleVqv3AaD3GM9zDIyPdE3jIwtoDB1RqmvrL9gv/+fXXoAU0ZsOTA+AP1x7lpehOEBwC6NQ
3GFvqN4xoTKw+ouOu/0Oo38YlIYYFDHZ+psHE48roSLCrD0vwI/MfavOG/HcEq06wI6hMmY9UZSg
bT5NGxx+NXcKDWvDUwM4GIJysuj05Oc9+v630J8W9/4rE8wjMNEeKm+ZriOHnSVWrt0kScVgswEm
QAZCcEkyPlSlsf68F2nIfVBF/9J7xCLHF5+f2ThCHuGL0+VwW6pnVuQconRibdCQXHgbDwEW1PN6
PHYsgUVU1j0Wl+GFLWfdUFn/KcwEXvXh3NRTMHmIZwdbrJCIJ6EBbWUMDOygNB8Jld1A3VqCQYaD
91GqiJO19PDrkFQACzMvFMLdk6vCmYgvS0WnSa6vg2YgE8/WzUAsmKAjCgDg6cCO37QvhXpNmoAX
RgLqnB8eP/oqktLljPC0kGlBsa5qJNhea0mgdMO6AJA3cpGugt5cGnBfYpLHnrdVWJwDTVsJvu47
MGHeM5W7s2QLRc8eVfM0HcxbBKp327TZ1bNZr1+hetMBn3ehRYB/s43ydccy5G1T0M5Kl3RbXT6a
TObXfvTjQMsEpyPwzJGJ/XpGnAflpDsB6m+X0GMKVyRX2wWx87rgo4gCXBCgodSiq6u3+hZNuuHR
RVwa93/h1gH0Mt0+HL3esZusTFfQkylyHpTM3OX4+2iBgOcsVfte2upoh8VsAVb+ZvIW88ABezpw
HoWroOoNqNJkYuqDtmmxRvmlEd3vRl2opMxbN+VcuYBRzB13eCVeEKQzx+ff2Kh+DcJZvZXsJhZ9
rqCez/2/CWKxk5r4Rb3spxEhsTQVlbNp0TANzehPHSrgH3XKugJD2d2BJApPRreGXqR8HedV2gwN
1S3/VsD+g3us2ny4vvN7w2KOpIci4EArqoo7Wn67vyGx5HyS5wGMNnM46SZmdr90H9uYiRgYjUJP
Fxgv6GKOH/FYRDxupX3UJPdPkHBk0MsAzE2BeVdgHR1JBRYZIbLTlBY0K5UoYTcnKW5xJBHpCL87
8wHH1r7KpYmFSiGBNIoiGORzFDC3clCy+2oDVXveGDJ/Cf2Erj0/eRKqIUdmeO/EF53G8/pR8evw
DdTmH9Ldip9dyUoD4fAScP2eKyxAU3Uv6Kh5Zb4CN6u5vGXDnJVPHefMTZ04WNycFOqSGf18BPtF
3FPuw6B7d2RHUknlJEk8VmoHFCBnG4ur/ndbaggVMUEQvN4BOhPvl/MlzsE9uqm7j05r4oOtRUfZ
52/GTMMT6mXWPix/zUy+TpwHP/8PSB14wBprwgZ1Qe/6eXqvdBS8Fb4rvvKTQkMYPnraDRMbBbmq
iFIE4jwePX5rqQTXjFoam9k2BXS/UeGt+fCVVHHDwmCz+YcpP+B7HqcCbdXxWpWm9cK61Z7V0I9u
QGn3Go+tDbum7A19paZM+3Y3lbrxVnmTGRrlJuGeSMiwtctGMb8Q+wyJeU8sN6+Vy3vnRrXjXdWc
KJzA+rwPm/t2HRwya3D3OFLYe+M3D8oTB3GPjvg0ZNVValZ0pzmAyocwQ7pNh4/f6zdo6I+X8ZP3
xwRc6oZsr3PXu3WUC7T7MCkXlV5szrd+r1smkP2Tr6uQ1eEpY5ak0UaZBBT5hLVQnXBO0sxDhRX/
EC+cfN0kM0TWwLggBbOHBy7uYPzYtccgJTLVWlUqjq9r6+uAAtTg1YvRRd1VEUw9MvrK7Cu2lSl6
FtiFcl+Dbxwj06tnU9zhDXSjRaIbW10sOnmxWAKiAPBt32xmIBHdWAbBZ0zEVqhasq+fhVmbg5dU
eajRqUmmxn3+fgH5B1uZ6ws0xXsNFJ4QHjreGc7437SYRpDY70bjP7COIvFRZ9Gn69+OAQ/8MXLb
kvmAGJruUVTIgWQ+vNdEl0B4rMxCuY+SQahwSmYrYhWYawxEvKLnZnFS7MJ4MHVkktX5ZbDgy8eV
SIu6dlz4Jq1atAGQFYDsTjIsWtYnqJxcJx38RhCH25x++2PRIcrEl+5oCFAF/hKkc41hhtTy0Mvr
ruh8ygMru45Zk64Ly/c8FWmRxhb6iZlNi6PrpglyJGD+7JUYvhD+vNw/9hbK+mTN3YPG1sRkfibr
CzPWBzoQ5a/zyfcSS9SXfhdOenTUoNG8RZXREXQ14fdpVe2E6PRdq/Sv9vPRBjTfHJ3+kr6t3C4H
GCK5OKU17EwWH+iaMBuu8y7dy1oCMlvcknrUqzsp4FdPENbvpJRKrai1l8wuKzvOKzyt83DcTBqI
3YlqKecHABBOavOVV0co3FUWUGXyPe/qWakZIHNtuO2r1dSiCnRduFSLa02KZnkFxN3SI46jKJyG
XHTLX7ZrlD10QtuEb29945ERO04106B/povTzQkZO0ZtWHKLbQedDcGbtAwCWx90gigeQlXFVu9Z
0FnCJxaQXB+GAmpLFTz0x9TBHPrv4WxFbI6uDYUUjLxC56xY4qHU68Z8evpW6z+0CTcKHwZz38V9
nx7PHn9rvqvP0KeqcL3eJYL4XrJamq1HECOxXx+DrAYdhhlsDSMJ7a9NrgVI7ntNpb8tLKlU0QWq
NnXC8ZFLHVaMdXHqyEAyE2mNu+eEvcVnuDuB1SXUlWadQAxfoan7Rf+W8zCJqU1By3oNwF8pL5yG
aRJg5wTD904FFXrFd5Wv2Ng4XvJhEuiDK1/YG/Wqx6lMlekMGl/qNtxdvZI+etuPq4/oMdcAJeC7
L20SLIVZsLjKkwARsxbgqWUA9gj6oBbcB9u+fGTVtI07f/6ROQPTrDsYHwd2jRGCCSmf2Wfx7Slm
ldj1TbfmGdUYa/RMtE5iKUaA7iDd0Vm9LSNSqPqzQE8L4ZTnNvTdcBLuboV3SRqWWtL0Gz6pEpcC
Fs0vRgEPi9bw6Om8Gw8iWc8BgBFN8y6G1OfR3PkEBc0KE11Vy9vYikHUd5YjY3qFG1wvwCLUs5o5
EfVYL5wlaNqQEVjNOr6Z67aSPfYjxa118WDV8H7gwOvq0ovmscs3wIUC67y0dgqSM/2A2Ul881Dw
g+vUcE+AGmXwyqNiP4W+i3UORkmy3y4gBULpkPxBM2pefDAEy/eS34/E7bp93U7ixthGxBvPT2tc
tJmjSt70TxX1zPqngCjGXRvWmKD46N6WwPfkXiP0TyBA/5ayzHAuZEuPDuwyh8QiI+RM2rrGg88A
g7Be7OE1DYdhScYN/TCY4BSQWxOtCuBBmYMjtl/Cho+4NiIYFg5oQKu5NBuuTw1xnKosBHvlyzA4
n08C426FUuOBSABrB4D4t3KhFM+LdaqabM1P2i+pYgeJUDc/2qrc4aXrHqD+i5Q4X9FfXdgFl2RD
ODZHPqk5PQT8OzRYwAz5E+zTl7Sq7M5jbKnawp/xuSgLWSRt7b7LV+VU3V6pqidYcSeRQBKGtlYR
Iy623k1/MvVpG2GIZYjWNqOeRg6Nzv2DBNxoapS5XA3v5wmw76jY0jWTl5zvFr6lP+DJAybyK1qx
X/zRuziFGy4/qiuEo+EgeCf20lOxJ5Tg64M9ST/VtvjkYPH1t4WRv1jUlr8rZ8QMmTOOpDicVZfz
bna3H6MOmWHmUVxcCFsiyXii7uR4wB6XnN5FpQtnyi54FYbkHaQCvq7B5B7PjSBm1ZUs4j2vPrSq
dT8ylIGK7ORrBXDra2jkvP6/+QxnOkwgI3M+K0HcrMX3gPDxBoJc34pqh/0bwVOxW9KiafDi6Q/l
bnRwOXCR5f2sI/0ro2LqWAEfIrlmJ2N1V8O9uabfNbraUA0xAoMd3mGyqXH1bonbqey0yqLuxaSm
n+YJ8kspd5uqBN1+/V0aF7nUDfGPp6hOuRnCMOyXW5V9ZKP779/8o+tc7fSmzivaLvOIQzUyBkYE
pOnXS0Ust+UAj28vH7v2FyZQ4MvFDKdWpYziIv5fkDSuY2qh9hPo/c5mr70TOpCkKhKGhvsneGYD
vjbla3ZgpwMbeYtBp67w5RnDzIWnagzk+29+gbpnYEkTPynbj8kGn9dDfl25o8tbKL6k8U+72r+R
sxMbjabsvl0haCkQNyLKwhvNuu5PLAfshPAFN/kvolJzQL4gjm5H6ZFI0fWGVgWeTCfVwBqrnTM+
rovm/mlmpQqu9uq1FrjwIkaHEGRb06ZNBYfH0miq+Fm5YNeWiykLo3A+FswaW8Efli72GrvEN3nB
ANVqDe5rIH7dCyhMOLHFl4dpo5rSdnzXUpBRL29kO/Xxxcxb3zR6X0WEFTPZ+bIRcmVbRkZR5rvj
09tJBiO7MBpzGWwei6Vtdc+FGSki66jgJN7qKOCXXHpnncJ/i0rR84sPS3Lz3KFN2M4nSDzgZTBT
PY9TB2zY2vaJu+7wMOhtj4EgQ2YfVcNsOxaabtvMBFOKT87BzrK7V1Zo/cXv98sxbmwpQckmNQxR
2FJJ4YBMQUul3yclUnd/6Vy4/icVRvBE+CvamWP9++V6OQtkUM+ShZES6WY5LVjcjDGrxj5zHRvy
GbNeWvQ/LqfGt7Sn4LOXGZG6jLG5s50CHZrX095ir76FaP36PTm6rJDdGNFRFpvTe5qyqaGkF/dD
Chpoo1rLLMf8ja7bTphTKc4k9dLhdNmBzNTnhKJL1IgK4xIwfXPJFcG3b7muY9gdaKOoBn5HJP2r
hIMjbPj2rF5cdUR4gd+OgIFg5JYJ9I8JoHiRb8Iah1Co/jkQHHNf4zb/qxFmSY0VsAOkde4Q1RLL
n1j5D6UGc+R8Bhga+zlG0n65qKTpK2XQGC1bOGtSc2ja28GymoeZlwh7hQV8UKnALmB8A8b7k/Hr
Qk9S8eCnB0ujrYz+jRQo3b0ddIGJKLvMY9yOppBtGeZ1ADwfGwIJG66NweV1Lw4ESNcz1xBZn/4I
FLVm1O/+RkyFdFpYycyb5G23wHknc7TTIGriHSb9sE9jJ/2l6bOMO7B4P7wTaOy+NP5w6URgvr81
6WN+X5FNi2osLgnY0O7+jnWFXPbMxEI1ZKmPQFj1OBwsdcNoyOeaaFGhrjMlk7r8QHDenkmL2Ozn
is3RNRACyQy9Yqp4j6/rUF68lU6x94XWhcuqiUAuuxyk9eZxHfpqzmwyMGV+OA7NHMvhO2IZvLhX
A9h8sMwk/iMbqCsH6Xte5lJ9lPI1wnQd8I9tXMv70yB5ctn3ZYgNh3YM/9uXD/91UdDs+yxR3asB
nfmJ+A2wD6zfZTn7YOy/CL9bLBaRYVW7tFmVtj/qomPxlQyZZ5zlfytTDoOgE6QoP69/9QvkiA1x
lzyYIOeZU2wbSOZ4Z3p1xiZYkI9p6PskUWqECOBbOkUBx12pG9933Uvtsve9QvB8QzhUtuN9Upun
1KF2TbvPJfup+R3kpM720kf7GtDSODL94ihadueufRcOWy8KGSbFc8fUX7GiRup1Ow5sTPtYJFfM
X/+62JzRJ2RJbD7YdA+SRQOjV0Jk8OiD2p+xQFHTkQItdvCGRHUTVo5lbvCAQKI+93UCBHTky0Jf
OEuFOQ8NSo83C78pF0SLfbKedJ4o0xC1B9VlyyFWfLGiQxbBKOPO2dBgfxYfB7vHqL656JbKwzQM
5SJoLdBhB/Kud85wBHT6egKRI7qZz1gw4b9fXJByxjcHTrcrfzDwoeGI8tfPXS+4eghseq3R6Tdc
wm0v95rKryb7V5nFrhgOWBc97xB5EdXaKKDUQoL5IZBCJWCCuOWsL2vApttrlGKU6Q7y3JF3ebOL
cH0Ki4jh+c+s4Hk2cd2VTFbfvxSkRDMnlvDX48ZJVjrhnSHBsvTECFUX6X0Gaf7v8fFQgzxXMXnl
niXRsTB7t+OlTWo2Wf+iGFldAO0bkgTK+my0dfW21vP0W15q2hTFSvwXNjNmhatKezJTcMAnJv9t
5AJOyFgK9FSnizO5rUEtGegMLKzkiwv6MLE4VUZPB/6YYwMqKsiqi8jIVzm9P/GOwuwo6dyaT9gi
HIYBj0rVvDCNhos42gOJfBGmaM5KeBdL2XqTODzo+AfAxC/wGml0gC/PVNfbjYHqGN9Luf27xvEa
0sOP+ofH+AuFx9HemmBnXcHonxu9ijZmqYBuN0wrhVutEgmmGE3B0nq1CYji21QyVhaD1Ew87Yb1
QJ9tPzz5wkpH8oBfgk28e0xMoF8d7P1vTLgf1mhslwb/Da/kAsr8ppnlMlDRzp6pp+9nApMu3WCn
23QLExMeGfyiBjkh0YEsYAuuI+fwtjoXrKW4kdCap6+orKQGIO3nNR3n+ts0l59l44BxhiB13naj
7J21Pqezy0wfZo0c2cdBzW05k5pySgv96l3HV/WxLjK9tUvbrH8zrixPiDBvKJigPmm95UOJNMVu
35dvcKCVqhi3ng8SRcYx6RkNRCD4zjSaeg9aA9AtHCwuyesnsVzJ2pC7sWtE1Jq1XtZayIX7Eegd
kqRfI024geAIRFdeazB+AlgKPyg1yD/s0QjNu5mOusSnthXPSK9uZLXNsH4eymbU1dckZ2bDAXYs
g7Gj6Xx6btYkDxJBcvPvX6VcJOSrcsqxOrCY2en6F/FGHd1DGe7rvz8eUk7b1aMmLOffcbKm+EeU
aIFvPpxKsjGSyF2bpZZoZkBjYwYqw48JX7IUyNS1CuJ+Oq3gr+2LMMLMoL1Y7pePtY/k76A6fPwK
pM/tJp/aZ/TrhuSKwU2xxCR+jM6urHkcFrWkza97KMXd59va+qTMpNT2iXu5r4+60R+3PNXws4yQ
8eu9aKJBu8BfT7EwizPgiVO29C5A1R4+uBNd57HbBDts7rsKqWdjV/5GIP+3U0dQVK41lp0Koq2V
d6QAYaRSBy2xkGW9+KZ+w+U6FfV+9PzAc3qeTSTs+1oAbJEwuJg3n1mr4s/dNpoOPKHYPBbOQmrN
inaiVVZpdtqtoVVqrbGr5kVw73BcjLNolazxtop8Ifg2raJMgq9Vms7loQZSBPLuWtxsrajyhw61
pvQw+/S3SVvhbQwEqrT6w3oUEhYx9Kd8ehKKNQ30rEkey9XxQeSr13dbQlLXYtjfTwlWCJnEpLrQ
YHOdGgsfauYSpcAzRM21MLgdgBzzN7Umfk4DDayr2Gg/LR4j0PzF8YTmJtvsV00YTWT7fWjFXNnb
QjILWrYzzap7g/jNI6DSQZqD26GC3FH0F1cYnUTuFlj3OhfH7C+8KcDBhzcloxjLM0JaiQ6gK+/T
UkB4a6MTJo1MbB/dv3xfa9q68gOBBxnI1eFoE/GASDIy+2R0/zu8FFSd6+CmINVBC3Y/nS4yUnsS
osDGHvJrtf0aFikI9jEzZDJB1r+nE5iL8JEkpke7VUuGXylnMTNikoigLMMST4DbwRnctWX6Sa9q
pQSAwruCuZsoeXR5Rdwy1cN5nP8mXcRJdwsCYTBWhkfnxVKOcyu2ZlKJ6l2LLR8Q+CpVQ8Pb6WbX
BvNnXzDvQbb7fHjGYXp29QXhdMIxHTmhmlHTDqShWXTKuM7gsxaz8E6sKlJULE4S6TRHIyn50siW
2re+UJpjwT41wtN29AoK+uvSU2wdum6z9yDEUSdNI+c6Bb5jHFd9k8SeFmb3h0dBIKFi36FWu+Rf
gT9cCnT/cwYGkB5QNUQxRhBg76gVX30nmVLW7WFFMfRoFHXJRuDUZGOPAehxcfsILbASB7BG8FXA
gcdc1WDZxevkFyrvU6tsDoGV0UmXlLyYMisjjEpWbCvk8JFaP6tCN5i0doWqnX8GiB8ON9vK3WTA
AGRv3Hph6g6imX0icn9B4quqHPSo/3xntRZh3g7V+82L3YUgUd3ZfmIoZW2sC4chrVWXy7fDdY0r
fZDDd90ziWTDXQh1jPZtNb17vxsNtbksIrR3wYL2eHefUQAQDjuVE1jt8loU7xwEnMoLpVYeteFE
1i5ypokza56i/dVwoYvLs38kR4LvkQml8TEiJJ5QlFIsh+wQNz258BzhkFU23ZzXfY2EMHnhxZyN
q5pSq2iLswqzEyr6btUMSueDaTIxIBsoAuqK6y0Q5WZLagIOLGLqeP7wOxbIkqvA58wDKXUM1t2J
A8h8eijWZy1sLV+m5XMGCBJN2MK275rha0v5PCPouR/aVqnvF1fjrn0k+Ojc4no0niXxqG8Wq25A
I0DY+0ConCqDW/qxQxRbk5pgnYj1OSFX3AZMl6wxcowmNYcmj8efvdq046IfSS7wQwxDK6KOv9v+
1/TUmRewIHAIwmCnN4v5wn+5rNFJehAwTq4BHZ6RbJcRGVZ8r0E9TvtTaxB630F9q5L42Ca8qMBI
beU2m2XwVy0M1kA6J4qSUqUfDj7f0CwynusVH8OsRMKU49ItFOKImq3Mn7YazsWBrFoj5ys9+p9r
rnckkJxtIjBJyQgBug3BIO+Pl0r2qVNZLP9/rldXENApQLnkGRlUioiIzZ7VosMdQEcDf+k4rcVV
ikV22R+3OHE54IZY6P067gpDRZhiVAZkvmUABo+tlqEv5dRe/1k9YvRkNMhz2l8/5yrt0oGfSbQH
3rs+nHyr5DXPwldLgh8qKv62nTMv9cVSzCPNcXDlySLfSqoyhotIX4d3oKEcx/Z3z7cJIx/SdLtX
EmavRJh7DMykK2vMZKzmtLEmY3oeaIdenKpAqNS0Ofo3oXsWyt3WuR4sHRszcG/IGJw6+Xbx/IZQ
EqatlWyQoGS+cG0x2CVCrIbQHx/t6XkjrrfxnhjLD6xmvNDxhL+K+jcLMlqXgyZXiGk2A7Am3ubP
na7n/wDa6Ehu8VCHqi3zbXj1o1feu3HowGyyWpF1RQtOi3dPupvlxjoBogGUFCMiOX+uTGCTessV
4wAnhY+zw7mbrKmbXlr+KUbfEMvhpPw2h5U5++hcvUnphTP5UUO+iM1Rl3htyLHLRQnWNljVjKPH
nnWovRtquVDPeq37OHKC69GegV20MwcUXZ4HS6XaZQlOhZDsglG7sKUkJW31KXxEDfXyO3oZ1HGn
7emT4DUvKd6ba4e8eyvK1Txhwb8EMzapTIL1/SRYpRbEq8SQSx8bNbow41sM4kBvLsn+hgYKHeMA
iJ7dMyaUIrnNNmyzESVTS8v8sHWNpFDMGQVMi2RsQpKj7XImT6C2TuygudA/qPuxjftg/bZ33vpK
HN1+aGd9Wr5jy6XZ3wDLkEACQX4y5d/MxjLJOcWh50mUbGvyqY4xtJDCi8Gc760WcX4xMV96rpw4
6Sa43K5Sh28mt5qHwUfoNmow71v5NetuCP52XITGdZxKLkZ1cmfSlEjBRdSxx39n6OvRcujs6190
DZrnzgXDDgcl4ZVAPfJDtCxHVcl0v3Krg931dhVnjW44CKTD4oY0N+aUMqSHF/dwuhbwqfnTh8PQ
3aAFgPSSxzmMycXDkq60xqj/HhS6r7mAoSVBzAJ82k0QjY64ft04Xa8epvVMHJqiTJ3LSYIi4fw5
vG423/6pRcUrWVayc1N5n36Y59STIKf0F9Whqfvxahi3w3DdUOdbbvDu2E5JTvlA21XNQJmEfEdQ
vDk53cGcp0piDangey1lY92tc+0c4ZsoZ0LIFOmxxe4xRPh5mEjwO1cMPJ8qpkTACqIBEXGnvM6h
XgmKBjf8pufeeX2AP9PoQMGUkxg3VOdwBJHZ6wxoji7GCw1xl++O9ROepJbEKilTfNTcz9eWPgNs
zp9OsIdNku6kl5K9qTWFkLKGp9r4Gd9Fek+d8QpGEF2Kvu/vN2wENlbyWrtjPud9mCcsM9k5zZDd
si0FkAbIXEsH4FfcIpLAdukzldPzCH7W/W40+9Go4QrpR9WKAFejdXYxpADssBd6iTRcmo2JIoYK
k7Dy4la11P3RR3s9+PgqcCmgpFFhskmm7fpS0hy3tLIiqONHZcd2o3seqrvbHqpxwFQywCYLhgxz
Qri54bvU4jP6Tpojy0PGil9XOc19fkXsKtMSdkwCR+Uo51deO1XIn5QcnLHRHFQxbuovkGFYwaq1
LuczKk47NVCcCg7vQaFXr9tOmh3wRVCm6SvGHxi6pyaVggA0jmcVxi8MNKcvlsnmx1DA2M74PpPc
Q3xA8KC0/erBUwW1QqpMaM1vnOyeT9h8k3Cpn3PTO0lVhtCE8x6x8mwVKUP1OUo5IzRjGbWY3nLT
C8qloJ3THLZYHqE1Qhw/p2c5h5EmG6BmW8H9atQvDmQb7Jhgb3qFL5lKOYXv92XuYet2aR4qfUCG
BWtf6JoJODiH1l0mEo7i0pUGqfcPnSSQ96aguZ7ehXh6MguIaf562gsOZRx1yqWX7R2ZNzq1GUTS
1h67HTIP4PXX+sInoxGo6r90KocGbnSr9WRD/aamebpa5lNyyJ+aqK7FjSpgh0eLXnHagX7mJ1i4
9KisbrXTOUwhl7DRFG7dYKW9lXM9s25MAeVnnIOrBSKOYxSw10zViEL6booSJz3bEh0qzN3fcxft
96FKzqHh9Re19vdHx2oI7xjOLkph8IuKL5SA6Vnbp0bqb8ISTBOHudyn2dWSc3tBnNLwb/93i5mq
ZdfjHYCsyJvwAe+o9qSGi2oSUM5f78YbHCqfMNXwfKDWCn8ymEfV33G+4D3WRpTBxDlBRLSMFcBI
r6Np2IOEs5Qj8xCzMUF/G4BMkmVZZq3ndsDsc6GsfetYYDXKbbScmp/DxdJ0WbYpCrTfLVqQiJwJ
qt0VQXboUvhdrgIBhKyOAh0G2TGqemdyvXPgqa3COUKT45ZxMPOBKCIGrEOhOBcuIFTe5nMk7Zum
U5lGoc1xY/K+6xCjnH0YaJiL2D6RnNCRgBpLVB3/OoE3VtUKt6BgWZfUNVdIrcd3M0Rti4k0eT9z
5UgYT9Cd8vX0kM+kB+jENk95nW5ANfHVIP/98orymiJWb5jXUdFLPmwphbu2doCTck63h9wvaINt
yPIZ8f59Xj06DefAMCcONwnbSBTyyEu2+aooZ/HahdDMYLjD9BPiPoacytUTumRkSdmRSgzcMcPw
rp7Wpz+38IMenCyN1B3jb8gMZ4Sp4fvspT6vYt16C5/2AlOz7ZIWM3qPdQYpPLt8C83q6rhWffJl
KvJy01Gxi9WYm4iabbdxArOZ7Bdawu9NsmFY7hcW4mcu+8Xag+KXXx8dQ6fKhGI3B7JyFHVCKb6v
ie2zLCc7zUmDfwxocYexozfZpSPN6nSnDsfDHGrfAsJwIYC5vzET/TpMVBgNZoSNV+dQn8o590Ty
NV62v7LfMZzON4AoZev4oQp92F/7VbAxCPQ7U3WSpR0jn5S8Euxv69HDSYcc3Asi1SFO+r6yRlZE
NlTgkNuY08XNS8cgFFEB4Y8aHFFsEEHbAII1BQb/EAOFKoXGkHX1ACgiUcFvYw1LsDYB/yzVZGkw
rw3fm/1UR97sXcUEbtQrR1mKt5VyfBGRBhnV5nB3HIM0US3GJblpeFuA4vmV20owdEsGfYUIvFpu
95o92ejSp8ZBC/RP+SCK9kKB6opzSo0ItQa8TIE0yl2Fn9VVC96zQ1JHJI0qh3GYE0kYvc5DglZL
KrHQ9ypg3m7wcZOGl25tictVosK2dXe3HYrxtoF8lxHWJ1SqHVfOReYwk79B3KKJtlnqgLCaY2t/
fuS5OcanHFpjUexqVpXBX3Lk9nQ0a5dCI7HcZMhf94ZSKvx40sK9n10tBMnuqjx2Kh8pnY0AKp6x
aI3y8vFcbG+hoE5jEx8fcMInfy+biWF3Ab7pD8YLlGBBbP5swIjBDuptTJtWk+mx/1hif19JKMsD
4xTmkWk8paNpm6an6p7hUZEPLkkemQNm7LRWxIzpXChwwTpCxOknKBWcsVE+RaBCjpkRmPOybFfP
SbQ4d7I3p/wRnmmiusqQq5oCtuwJEZ4ZXUCRpOPHJifhqeEIdS2sWg9yjlluThM5CsmgxX3VRE96
HjIlWu5vRCFhYtYtKJNa19cF72SC5pl7oQysEqer+3/OiFzuJtxLjPkfTVxUJEUGY0f+9ZjL+YO2
xNDERG3yvJrKLoQde4JxINJj5wQNS5/5kSIs//q1Z7qsxkNrZ2dp56OMDRC0GYklZNHuylswg2iX
XSJZzZo2vBrp7hqbOQ5Mr1fCZsqMBnOfVrP/szxlTNhN3UKGDOtRNBjKMxPuJURiAjinsfGm85pd
JljruEz+/GCjHKu/a9DrkmgtuSWjKdiJqhLLEKABxB+z+YO3xrbnVtAAHMoiA6qX8zeSNqE3fjPF
xI6qG74eWtO6SuikE3/fFDo1CgPRmqlSY/HIyt+nb7HfpHxBXKPyws91sU/uhiYBQFeZNE8kqIgi
nBbW0h4pYtzrQQ1lNKaxGvyBIFT5VqMUz11qMVdVMpnGa5HLM13uuw3p3t9vIkWvAV4iuGrVpw84
J2bUvA+Sw5j6u5nDoK1P38EJ9uppshbs0v0tSqVZK5pxa11AFN3gK8xAHChEdu1BJorslj+W403h
8K3Hzx6IkMEPx0QukaSaGBvf4lTRo/Iu5DnxlPCl13G2j6wxwPASEIYl9SbJ8/ixjTEJGEzKWqbH
Aibq0uPHXkYZTXmVY5BnTSFsk9lqN38Jya9P2aMgzXPacrVUapyCzyj+h1DRfEeCDtXAjXkQZLbt
orFvKaGe7SqZ2m1I7/IDCwMZWv40BWbw2JxD8edL8T/UbSh8GBI3t3KFXd8QoaYVTIgca/ryVCiD
COip7qrwkZ3TvIPaWNsxy23Gyd85+03+O4NubbRIT+HTsAf0csK77Nx4+wXTrHCfeK2quiOuEnqp
DVnJH5wyblvghhbMWxcwvCUBVtkcWzm5J2sbtvCUDZqhzyv5c/rYvBIvShzUOQquCA+U7HUVkLS+
W1lBMUsI0WkWVL2zEoSPGzHOoG5lxGuFNRXv59PyyjbSzZq/SEXKpxboj7bO6gOkEs2X+dlJ20CT
K00dL6zfMJRvQRXAGdNm7rsd6hRKlS5x5hYkLOok2iLykjxO1794X7RcabFr2iEo86QOVyM9e0sy
rWnDevIMbycBmBcPHG6ldilutj2g1yuAK1tZrGfrhCKgwJMLx7gMTT5LmubVr3U9+kd3wZJOApzL
4/MENl5n/4BxxSI6D2wJveJ6vOcAKCS0cICafvswBvSuIpGbiYqwV8WB6QWUuEPVV7Na0umoYA0a
xazN3ubt5qVBzktM4vL+kKbUjPuGayukqVSw/K/M/I0gefQZ7WjtMeGpRKF1kWFrS57Wfqywou+g
aREXOzykGWPmD9ulBgmLFTmUegf1X7ZSz19hMztqelpotFI6kf0pnUcJfYglCgc57MZCZbaKWvZL
U8rQqLgUQDyeq6WxK4H9fypdCIsZfyETDiy7j6XVKc0yGLYPqBAOU2z6v0RJIbuNuWUwh/F7xKQr
ChfqdaRKlkeHtOTy+EFYMY/9RUMKA+jP/F9+unxuJVC1n6c2HVOT4at1TgfV8b8eOuhBNiVwNdt+
5bBPyoAX5Sooe52vmXe14++m8Ay/nF2UxWReGcS25W+JMhF0dqpz44/iu5oSt48d/4mfLGMk5y66
AjdPNrkJL8evxCzaXv3URsarFNsDEXN64urtbPLJdjHjpvhCdujEqtawIpmn3yLpFxte7Zx9JXbu
welfPlc38Bcvl0Pxqj83AUU/Y0OYBPQaEf74Qibd1K04YGNL02G1xwHiYYPI29iTsPoPZooRxyyH
frwfGuKa04+z1owxh3wtuw6Z43GrornjH9Jha3bbfHVRc4jdBEDD6q2TZc+jW2uWIHb/YJljDgwo
Iocdw8BJFHMnrffK7/LrdGGdydr6wV9L762N2Qhhn4iQHTrdVMIHnG6hIW3cRB2I4rs9lW8tOukI
AhSHr6L+b27v0CdLVdA610IB7rJwBhbgG1p6+pwc9h7f/dCCkgOObd6uECagE5Mr4X5kTf/6hTVd
CGjVECN9Jln1W8XgEUa/sNdiWhgX5BntDkjsK0TscJEKkgE9kjW3D9ialLjZlUPqDSnzhJTs5G2y
3HJvV3SXIc/UKeYYKmtKXSM+suQ7Wa1b1b/q3srx1PXvYaFfgSve+3GOhCbnsP81NnJBvPozvZOq
+ucdsp5K1l2YbKsWId0lTPgS3nnPKBGID0jJnHMyK/OuuvJyD5lvetJrJ5ukwRprdhF9uz3KS+TJ
Y6VRsEflyFEyaByP6Rge+MZ4hIx+pWdN3/zUFgwvTYDH0YSvzI7JOdYiugR+QDNlcTfWY5/7sfAN
fKxhitOn1eKrEaTWlhwANBK7nIUmxH1WeupZ6pTzrtfjGHVM+HX/LXj1A7Cv5qjRtvrOJUsKrgMU
yc2oOvqmrXQYkFc8HWulspjH1wPtCGR2yaIAbATcoAPNDrWetdl7TDQFSJkSPWu7BUpkl2/WNkGS
LOaJayVHjUa8ZYlIvI9+VtaAtwn45oTc8bjHUcZVIkiCexwUgAbha8CrreyzS9BjdVdE/Yc7pNdp
tvjQCvAbrazJ8KivLIXGz5QPssq903d9q+6X1R7yPmElN8nRZcUVIxBl6pTlMOhtG6wTWg1w6zI3
sn1IBafN4Vip9Dce3yqp9mS7TgCYdkX97M5f7eKfUtBcJDkOCe1kU0T/J/UZN0gb3+06uiRYS8Wb
tDYG87/vpXujU1hxP79cjlF6yC13vRCVMUupfHW5M5O5SvqORwbFnJJCq278vVwB9wTxCLeUOZYI
JMaU+PaQ/gXotr6DPt3kgqQivNIF1joJfji00KAHGQsNqCpnYBDh+h410oW5WCKxSIOtRR3/27DN
iDbUKeTEg4V8vN8qiL29Bl9tLY/isiKyVGv197cFi7LumR8eCZb4D+4aOzvFlM7pOVIUdqe8fxv4
U1glFh1uVIR5GZqcuJsw+2m1yx3mLhpKaRC+/gpMSvDhi6dfOYktKWddRULCnJY/2IPSUd8VPuVf
RbiBANizhrQfDKa9hn+R+6+o9/Nns+tVhEV5+6u2dBQjxqXcCDUehQ7POE4BPBYtZKNJS0HD35pH
y+pep4zyZGaIcBI6BQ+6o50fAqFGzz/VW+9TyPee6T6m1gMlojSxeb9iFr5+FoH2saYafoAESBe4
DqMmoWrIdKZ4z34RXPAFdDGvnrfFN72pGicYfZX7Bgvamc/xhqph5BbtPRXUOY8MijIsANHeoJo/
+gbOKZ2CXsC2LALiNMigrk6h6lgblaeCqNh/koHUrUxFvpaWWAH/e7sssl7pJmHY1v3MhNRAJSJt
BFeKpXSL+DESN7fUekFtmcl/T7ccU9nNldgYbFakveO2NbRcASQV8LhIQ8EXSYpNoElY8MbZJjOv
O+lgElacU3f7/Q7VOYwzYBAe/C0nGWTd2fhr/JBeVxCv1VjfOP61Ae4OXgMMKAtoZH/XLI49Wfj2
cnXObCw41s1GH07wfCAMyZKx/DfTp7VGmxngWFKJ/nUb6RUldst9gDyhWlpuoutkv/QtU5jTuG9p
84m8JQ23qpeCQjcYx8P59SEaSRqTIT8CmkYTYf4A2guvQ+0+OzmZ0W+QXXGK/0u6IC6pJTEisFe0
JC1ZJ/MtbveVWApMQzcpIC6pw4DhH/fdZa5dLw30ChKG61NnYJB9rVXJKw041L3U/qLGCpdWu8lH
Lg2J2b79AiDG36erk5EtlgvGPD8ZGiuQijV8Hfe47FP8Fcmj+zM6RadeECuzzmoPjBKRy4T0oMHk
vnHBSxenfMxx0sbyzsfs5JAVp9Pm7rxr2ocVO21CtaQjTIWKNaR51X7CzSugTNuPKYbjTqO2TkjZ
4fcA6PSKkCUtRORR2aDvOBz3f7jcWQ3R6kaIzQkW8Sk0sgdJ+vxd2sGf/J+KRuetFen5kBqW+Jhm
HVyR0N2TsZKenzgXgCZZgx8daFh2oT/AMo/0lCRnsbLrs2WtEJpL7CtzFZPW+az2kXZsCJV7gBvg
kYIKndWT8xSgDBSS+4GLdZTWOD6Mqhihq8N/xlNqLFsuO0BpKXM8A0DWRF25pP6dfkBv9m5vgsD/
J8djrUeDoIwKQhSRdN3jGVdRsP8GNMxpi0iiKZIEcotK3jTNI6cZy7oXw1ZAiDc+xwP2vKqagtgU
ZEh7VVVnCi6bJjkexIRO0apid2EWQ8ezXBptcbg7QHMS/Wr0xwfhzlfusnJQezL72pSc+iFsMQso
j+oqyB4P085KXlL/mp/1LuMZs29vUNfx6smk39HFadqGBeGkYQi8fL3qh871LknA6/GT3I519UO2
pA93Fxpdb1VLwNUIdickS+umkDsTElCb4YxAmIwPT3RECsElvfRRwvnKGYB+I0tOputrheiscaUE
ywVTptOlUmrX6Lq8mWtC5pFPEe7sqWEJuM4nbJGLnojBPc9SyHcN24PBkJBDhe2HraDehW4IgtDb
ddFpBlgLMbIb0E7zBRniLeoEtMCiPK8PXL5XNntC2d7XHPOgYX1EtAS996P3qncFE091+GPotDVX
C4TvaysjSnOSAe2uGoLEqkgZentj2EWzE2Iys4laWdq3LthE45XkqvilPWguNIW3KAxjelcLhYsH
8fooYz04c/DVsdeXQBNoyow520TMwvuZ2U2Qk6C11qFe38Zuq8R5PzTdIEzGIFQPH+VuucctA2cE
toTdclUFdkio2SyjjPyaar4u0KbaMOzuP3iO8BTBEe+AXNjECg65fb5J4neLmuacpkwILFEC+8M9
jHjA2JN3GG4toJtt08j3c8GPzXQxmudVVCfLFiZa+llodkKOiHIKKVca0x28Na6xVU5tvVQi946j
2B5IPRhb+i7r3v8353F7PnxI2VBvjEK0KWduqGyYlrV+3VCR6wtNtEiqMIgPQk22tD26BLzhSJyc
3PWJZ/JbcBPaHbTPZKBT6r7pcZQCgbipt/lDsig8SVv7twJMb3RmTBmhFZirq6fIT2UpNrV0660H
FuDAotht7Fp2lAU/ttSus01TObb0oazmwX59R8v1W9XnPc3iubtbjS2RY5cFd+UUikSWutBJ2Y50
OyNC53OROy3rYyM2RcdmxVnpMBTbkqpayA35jdBpJWkQOGwN90o/IecBwEDZnCFx/V0CmUEbz3pM
Psede3Zjj/b0RCHhAcopenyL9mEW6nIwUQm5e6mGXaDsU7KUSSM9HIxuDcZBiKzdk9y7lVBHalzr
djcM1FbBo2lzzbKC32Hc+ttMiKpQl05KB8o2jlOAPDxk5Rto1+wdl5FdJAb+3sq+EksUzt5zQaGt
FNKP3DNIX73DnqQA5pTnePmjfzTmflDkX3f+6zFhqiPQTNmF54bW1wZNaX6SaBY3r6CMUmSRNOCN
bSos/cwLBKqGzD7udYXJCcgEhUP6JtG0Q5PoTypQB7FgayZHsMhRYJE/l6mS9C2Ard0pvCvIzAQ5
VknylcNU6rU5rhLf17rnnwL5/s3Y545RUoZQ6QYYfM3phySlaOBBJrFG8IIcWp3rDXrZnna2Y8mF
iFwhAXcSqeoOZBqY/KgMG+diiPvkAVLGP6cPTheT4KRiXMC6d0rESzWqRWbpnLcll29B/0OkC+S7
wVX+dDKEAqK1uHCJBQsYlJwvysdkKYobicY5Kx6aIDggN7gzGq0h8DeSAq1IOEFYy9BLjOiSw0WI
fftJGJgviYRarfCsHuFJWu27R1e+hWrsOMgBZcpnE73aRQpGn1GyHtwnYxceggyqU6RkfvRH6zpm
frBvsrhZnn0Mn8CWrm+XooDgTNoVsnl6aIbGDrLP6OUHhCB/5YhlVqpo0ushFszqkh7DaIm2c9YC
PR2DvyTxmK5uZkqG6H80dNkX34lrel+7OZWRlPXEPBuu3ew2fqqHl8Jvcz2QlRtb/fDuBXIy78CL
6Mf0WUqK83rd7buwcHLKTwCH/U/BBRBnZ7+kdq+DhycGxJ7qdMny9mKRMcIlWpmFHUnBe88NCSuG
peC3orCEmyUAVBUBwQ3E3Y7CtVwXCaFmpfd02zEa2GVsRtOwnMSifw+xpQAnlaivAKxK/gU/v6mb
7kot0HpT18y3xByY6QYBSR5Tf+IIcFgFUe2NE1TBhr5d7MalYJv/c36MBldpJDL0aR6OarqMtWH7
dG3iLJUBYU0GnS8oZfUp0V+20+yytFADDhscggk6rFAK3I6zpE1mSf+xdk3y81GCOXdV+uLFjEwF
pd9MrXP/Czqq6kOfPX7V3+0Ii353AXpgDFLGd446cQM9xds2p40bG/SN1gMlIpyIl9HWpPIIMBGy
rTmSKiY9j02q7ivqXmLJ+JsGYI6CCZ3m5uXtugU1G0X0SFb1fWoW7obfSHKNpFujGDtOIXy7lAkt
nDYSZOuhmNkV5GH5EhjCr24lKBjaQm/r0OKytDBY5t+c3doNKpmWihDszzl8S0J8iRnAQdHva6jU
jfrSkgXJNGHlFrn69rjGpICKKnO36POLDe5JE+UOhph7Y3aSRj0V1j3ZYhRJkPKBp+HQZj4m30f/
krICYKmGIyMJiFKcIYft+zxXpIT7/3NQoTvw0ZPMAuRVtG2thMhDDluyrAxC3CbOUqWlZJ5wm703
8Gyocw9o4PVQzt5jPKgBKCVRHvNOdAfOC8mRKcJg9kCgGGV0L8JGd7ncbu+t2T59kSvozDPdWKu2
ZvYJ9CLL+xE0TPXJSXVxGqH7LAUIaTFupbGZNtwid5Lnf8drol6TfK2eXvzLNVcEOKXMDdKePPkq
YC8rn+Dt69k0Vc2sXeaIgeKAJUc0WhdBBnqATcXuoAsyG/YNFCs9WKY1RmAyur+JDrYmQaBz2fSO
WA8cO4v7/ft5hIq9A4BXhhkFKnggBmBUDSZO4hoZmqf1QmzbXR3sp51Tlwh7l/26fi8fGa1pbYQD
mdL6VFPaG7rJ1iHCdQ4fpBNjakyArJebD+5WbmHKOWIRHbVm+ju08rlv1kgTZeBRyCLsEEioUKux
+VHtXSdZDjag85ZE+ln5EyMbkH48mZnmnVDWGYGjqHBGm4D+fxYrBWIlvgp6e5z99xHIMpmhaq5V
avKqa1OL+6zb/r8KiIuiTkvMrFASp0cWvwxTha34qsLA7260B4/Kn9T/5CKGWlnuXrcGkILkIkMU
FL4g8aNCNmh4kgh7qJm6jayKfIjfIpS5nYi60IA1wNT15+eqdXHfCV8vtGccBdNp0hGrdJw/hFDt
duYiSMSN2sn/EifzRhChiD9CHemlYrDYVEi9qbzK+pjotV4a9wJssyvYSrS2b2geYBBSGIjetMUN
z/Afu1zaM4vw5ZaHR+5mOMf9lyknHnF/QS0/RwmapNk+71B0ASbX7Tpk3/2gHm+JT9U2MlHQcfms
kc4H3qVka6YiX1p6mJKD2TCGLM1I5xrb2U+HkTmR69/yzBgKJ6q2OSL++wDV+tO9ZvbHp56Djv54
OrTnA3LSgYu54gHOI0xdg9tnnZUAh4Y9GPEL2C3Yw/7sO9w8/L23t/cWpySD2hfiQiOJ0PVHYklV
RGLtHEo4Kf0Y0T5x8IkxZa454syI4Fni47PWAuLzRjLcdhgHqAfmtYAsul/UHF1NlXKgfMiVFRCp
rf6m0wQK/wMPZsnHWWIZ6d7cr0GZNrEZ5iWYIa3CPd7ykgg6J/Uf57pgn2GQJWS2u6Sxi1caXoE4
pHOvsr5xw/IZcZxFcv84/U7J1nZxbDJ3jKhYvVgnlQtdXDNI9KbNiwLmXZ+lheySFylBbzbMM98x
sIB890Gw7Jnhls7x4zboHY5W6KJGAawNpplgrbwjWiIi9M3Vtcm86qqGWonJQvMQR7JFnabN9M/y
Gxo5gTcL49cEr5872Uk/Uh4LQB0seP8jw21wOOvgwa1GoTIQcy5eewZo4uSd7wqtG7o7rE+4EPVL
BlNRxZFfeUq0tmTNsC7gg73gDv4bOzs70RWaOx9Z7AF48bCX5qyJLpRTu/OLCXwTw4t+x8Ysd2bX
lbjfXSodBXkg8pCi5jkQMPRr2jwcSCA7CtS6RbK0v39hVz3El3pIotgu1WJ1l29a8oYLDLuWXD14
mAz/rE4vJSVjEcZO0pnxNyDIjVD03TNseF52NX2z56CHCUIAazsHg6TrTtLL81aal2hpPTEx33sk
8hlyTgE8tu8CI0PIWTyPEHhZqkSMk7LG5AUxw9u9JBszUFnCOEkMDwtxqOgDPRRU9qDCXPlE/i2L
yTJ2ewl5060/yCjxYmljULiVFNGig2Ld6t9HTusEwenpCJgLdlBR16bdw7b4Uacqn5BTJCaqNXZa
1hox8NYAUILK+6PUX4LcMPElmyYOiWzpqjc6P/fooQ3LRJlQHl1VR+1tuy4js0wqqQBUi93mJuN1
XkJeAd4v/5+t5L8888ik+9dzz0u3ogufv9vpQVx9jr5zjDHuBFiD0kGK44Vg1SXhV0o70vez3T/a
YXX+syQyCd99XiBUoFq/oZ1xyT1wGNW33xhsnGZAMrxg4FQWCV1qXs4ZjVdk530yVS6yQHJyDMZk
XyRm83uL70dlFFxGU7KbnOtf/1FHjRslJf4XlCkoJ48NB0t1HmwZB8UI0KRw1gyMRXUgHFUyrRGM
fSAjW1x9sL+FHLu/Eh0H7BIMqNxXTZeqz10iDIvzuv3jMTtEHrKA3nY3i0OXEMKFx3W9Xcnzh1P4
jfvOQZhbm/mgCZsAn+EjC+nn+U8MAVkYtwrKuJsi1TiAnNGiyRs1ZNUgSUnHich3999v7Mh41iL7
Qrjo5afzIrQlskDNOLpVwZ8A627LRL8L7hlxqON8AhmzhYfBHoR5xSeVBR+nA+iZ4XE3Tcv+95tp
+FJ1tozestFL2MCm02AuatX8hM5ro+C5aDN6LLZmp+JUiw7Erko1r4x/+npnuktxcUhQG6jE4htC
0QQC6UfipyRoRmW1aoiNH1xfWLcA5qKB6QsFU+73orDhAWAG7LYPRRbkPfUAfl27hzIpuPcI6A1E
IK01BjiulEJyT1fQBztrN7O1xu0RWO2F0pslyd3tpgqPp2GB4BpoqYiKEiu8FuAc+sNprruTh1ct
qeJ1RyjkMFmMV4r4nwp9Wl3OtIep5eNCfBbaLgJLe5Fr4R3DoavBfCkJSDWdsFLOH8KO6y2OhAhZ
WUyFwB/53tP6/REaUtN9i4bRNXb1cSAKAt0NJa9CLAi34zu6Y1oyksWXyg5i4c59FzPzWk97d2rE
T01q8sh+ucHYSrR1bzfOUqERy2eIhOaPmiXACBw91nSDozkdyP5iN14d0iXlVrBMcMR8raxYywIG
8nAof8HnsIMba0LulTo8nt77ytV+UO6DjD/6lK5ZfWOcVFuHjLBzSp8IfswU+wfTx+HqZvoqQD25
1Q5Ku+hi24xpcO7K6qiiChwytmmBMrrpnLK0Y9YVdrrAJNK9ZLGpWse47UbZ8U7b67bH/kNqtVwg
ovJFxpxhZFVfp1lZ6/2oe7RQrk7PJ7yq2n7Woko1vy+vruCMWEy0DFqXZgBGESfhF/PSkhy926Qt
shlC1dV8xBIu5A5LFaXib9IIIoJcQSnt1UzmEqmZuJrOsWedF7gPPe8ddIf4ze/Cf90JCYTzRNsH
V7gvfO5z0Sqa0Khfn5v/NZUSTSim4Nt1eXhUjtmTICbNnVyP5Rtsx0ezcvZpX8RHZvntTXsyQ9/R
xWKvUyGv+7Aab3gUZq5AD84kn96K9FcKZsBjNgfxpYtxE3kp4U5LDM7zpc/5r10tLT8oXwyZyNvS
cZVVclfU9/+HHuuyJhsundM/SEIQvbrRMHu/EiDXcswK7flyw2WxQ29gbWkxqcCQnKopj+zAcZS8
x7sZ9WoqVujaXxoAXB1wtQn2jUjL2MRHYQajKIe7iSdTaMaavxYrj0nOGLmOg5/yDbpAX4K+XCud
YarlIrU+1PT5Q+24oIpWH4hMuEoji2VKNmkLS7FD2ymdEVdZURErer/zgoLVI2nny0Z1iuGKS9SM
LNeghPhU9mx49+bFxaKiz+x7WWZZgTWT8VsKrzVKExV0wVXJE2xwgECavZXzFnxyIr+ZGRD3AKAN
2WVwSmJF4rKaBnCdn6z8yQrcqeYdom5Jn85fRgnfKcAi7Qt7rs8VYbp6FNX02Rw8ZA2FLW9TN44M
C+XPg6pqsjDb+PVMYplZeexx31B724XZyO6jrnelpe+dS9CqOGgK1F90SMpGFb+HQbNxsDYZksga
dzoZhB/8vxYPPByRvtleze4fj7Qsb3eqzE1G8egjLEJhe5clxxJJRc1P8lMSueutH2Zi3hdu4K00
fBstWAbrkX3uBCsAgL/A6bLD3LgMAOEa67x48u/PdkFKFy8VyCaw29Fyv82yhXBy8fx4sOAxRoBt
BBMRcGUWJDpHoRB0EHsZHHfgRdpR0cBpjVzGC2hwKXMKkJ9QGmo6HkWnrF0SA4tkCQGVz4i8woIr
Rc2Cvwe/Hw6TRvoAMnAN3NU8yY949RU6A9kWjy6vtNECiUjwwmjPArnyio4mkrJXOKXyDpL7lPi7
+JyoIL+pRSCH7WKaIi4Kjk8yHZCP+xcfoFNfEDoFxIFv5bqpTfJ3+MLQtXA5imoPB3HZUpkV3cBt
6M4Jcq4pqHciVjQn/QHUalve/2+J/wVH7YlogM2Gy02RzC7GX4ymV0C1vud0ayiV0QcaNLuU05cH
31gXCkWfkB002yzGy34+6gKmenXrPWWGIY/t4PzaJHEXqCG8hj9GwFLLu+c+tRduLmziPQ1asgtR
sT+J7+yjFMY2yw6Y3VxRiXJc6A61cfjX7fY1bXlLkxLGCCG8o0IQZszid2hIyEOQ1f2zpl9TegGF
3MOVj99N1yiokE/IpakOd4fWnNeaFgfQnq41AZ57oIoHiVjKbyXO5XpeLTT+8+vAGiOUk3+O6DWF
165sToKM0jJ0V1rD3peymfafIAG6TsHEKjYj6cQ9FrPJG1Q/v7it8QwNNguFBm652z6RahZajth7
qO1KViY6r6Z8dmfs4v0RD0pItI6sQco0l+w5YWvfnWk0NxCOs4fGJf7pI/OJA/Zn+CwZA7LJwUIs
OT6mqobVFsRcw/VV7Y8yQJl3V+YgDS1onv162eu7f3EkdwG2jGInTNiMK8gHqA3/bYWvkLjbCdNr
v8wzYOvrvC4aZTmley/Vc159MKcXbUB3DfVtccNGi/FdylkLS0z3+Km7bqyGLp+3mG0b8HwquAsZ
iJjXvk3Yfq4DIRmy/U7YtdR304hYAZgztfWnxWlliT2u7xvfsC+Ry6qnH3hwMW/N0FSPR2IQfY2o
GdT+AYOFAkaXs4J1RejJDguFCb8wimhQd0L/4OHTNTvrNyFIJ/eslJs2G9Itiw4q9DrKrhSlJiGq
mQkqID6VI5KCmgRlA+R00AO2lC8/gCwrUPIzpca+lKNRuc1wISWCypH9fnjB6liLCPqK3wXcz+Vz
kqkCZr9ZCyQ0TErRdvDdb75JKiu4iABK0IIPB6hzX5lUcBBkBVqNY1a2JXOBAgLKzwjr50gHh67M
9tZnJ0YgA0hvjs8xajTa8Wtf4EQavNJIsSsOZaCZZSrZJW2i4c/MCYSz4WXzjZRMuOZcgwqopmHG
jLh8Q/Eebu5fH41CfKLLaX95nVhYKBKg/8ZXV5z4wpfENMm/foqJ74yRbBsIwYVqZ8op6ZcGgKbV
X23RFV5FtzmY16pdgvqkCzVPtpwByn0lyxczdMir9yo/fOzO/4iyPu2MiLRyYZCDqFsriE2oekz7
y0DNHvPdTY5e7hhT+V+69PiwAUQbWzJZLuQRWf1sW90B0epzPmVgCszPZRKNMAyibFMP4gY8QNfI
jBLTGjBZz1FKJauHTX80e/n8B3CnidHejmA2JAXbAspHkOyx3DlLVS3Yb5LfuzvVaBIde7nNbR54
BSESey4d5wRyC6TEL38OiCsnb43ON1kJxxUybPwy6RR1Uy3armehu2KFqxDL0bHcQvjCQH4n5F4w
/SC47HHLKMhT84jVcSOZGDiMotqCE4VmxORT/tZ7/dB0Tcf86UaZs2e0jEQOzQCYMVoqJkvwAfhs
etmD8uQArDJzVJVzp5NEZdlAXrb5uiGx7jgcHRH1Q3GUTO34IgzCWKfI8WCpD+P86VmcFAp/VQms
p0apOwvJU+Iix3Le+U6GYfe789qePkRgYl819SB3jijb9EuHqTEzcbpKMnMJsKq0oPSSHwOTdTBG
z+EuERbPsu+yaCuDZ5M9GqzeyK9MymbXgtWGxFL9yzsaLXJR1BElHwMNIQjE7TwycZtJJ+mSjaI1
nox5SV6SJfIv5MvFmaPRgKwY+5RZh5oisqx0wQhL/yT0e2HrYwAFO4dSd1CIHc2h4sDPVfhXPaLW
lYjcejOCR5cRwALs2nx9StBdMVCUfGlc3dck40IgHGAmf000+9Av9MURfUXpG/UzRi5kd41N5fCy
XlIXv3YRULYFaPw70aanL0p0/e9e9pcyldT74TW2jvKEGujyn9uKpXL6Wj9YowybN/Ols2seCjOY
qh2Gd81W0lVMObXrHO+RzyFpDitv+yatCZTUSA1a4X+F2MSg5ZscIR+tdYd//Z3Oa2/uWW8lwP4W
+46P/+K0MdpUu6VkaANf/o3nDXXot1eo4vj9KXPZkwhqZ7zM6xzELmtlNPezOgHWvDnldjmk7Du5
ymCNr4Bedt6kj9Scr1j0hzaRFeelQAmwk2XaRx4riosE7r8hqlmaNecIbu2sVD7WPpx7EGQHmYnZ
ijzuvqDKdiXaq8x1BFp3lyLUp+bgcKxJlWZRnmco3jj6Cd+R3f2zEs8gQvkdB/7sWI3e4B+8xe2q
r1TgsEJP9O4GHyXflUipCyt0GHA9Pe+JoVl+GXqFM6XX/amd0pV/ag8TrIy0qr1Ue6ICjW2ERoqH
p8HsE6EHZeOmFhbOs75vg6u/dLjNjQdYSSgZTxlBltBVlSE1l2EngqBIbPy2SQ75WGWcpOf38L4t
vrOHskfc3OZo3qkkY9T2qEzH4S7/JuYWWAd0+fUUQj2xduOJqbX/ejG8/9HJChQqcxPwOn10iQbh
Lfd5C+txJ6DU85m98HMTruPmC9E5/Wiuq2BCWen68T8yTAo/6ZAVYdH1OtrFNdea70KrVLV1HuXs
FtZBGLmsyqdMyQD5MLnVunsMnPci7QII1d3kecXOLUvJixyK3h3hqJmrEB0w1l4A+2NPOWX2T4dR
k4bPL1DtK8HvY4lZo7q4jC4sYLxlFvShKj+LCKSXE61rg+kmDY9+1L5V7UOvDrB9e/006uDlMBhZ
d/nFwffgNZ6oxyOAi//+LfIDF0WTnhhCjVRiiMAVQ4rs2kF+SZqbH3YPTV/4bgSy1rrRZlcgvhiv
wdDVcNdD9ieHPtDCpXy02DOEMVQMgXDECVMk5FCIYYsy5d7IqTp6HCRzc3H4G6WPltPGsgrxJKUu
xtZ1bc1tl0LzhjBZfUVLys+pEUXv7eUualOF7KEm/fwo0SgOOx6gvNldI9qJ2C9IWV+VJLJmB+/5
3LRB3qZfxsfZm7Ls12v2Y6vY3vSkuDZgEGhmI7B1UqidfrIvE7MY2sEc635uhZhhE4W7nIc5mMXT
fKoFyr0xEypGc8obOI9n+dgZ6sHZ2G9V1uwTZyOnU1vXMlEBDdZdptDfhSKGbWgDrJbczXu0nTac
BY3JGOceWYJWC2mFvO5Uq9UF6Y3sdnd+J8c0OSY+ms7T5goWqYeeFPv1mORgoaKYt4LAJZt7ybi0
6mN7JcL7j5kmito1CabtMJ5VARh1O0zOqi4PtQ2pzFu5BcuIi0OqqJ8Bgf1lhMKvG8IjNRXWnbjm
vqnOn+jNFbS6fG4aPBKlQ7E0jCjkBJUKOG62WKKxJoDU+cxR2Jand4nIefRf/lvRoB3fLWbN+QnQ
mSmZKPP3gvOEBPXZM1Kfax2ndtIWugNaZ4L+QqFcOrzhTOjzUwfiVlqbl7C9ARjRdKTumlrI6yGU
7GTfxiZvh2AEl5gJTwWvtUrTZ5+3LhCxs4BqXo96y3QI9IkCHP/Pwk25a0ptCOj77q0QoLHmI50R
rUoW3xY5u/ESuFTY721gJaZLAFV0Be8Mz+h3X7hGROoGj1q2kZ4olcXJMlG8gEg45pRo2jgbZZQk
HpvUk+hgn3XZWmP5EzmezD6vwjY2ftMDKshA/E/RlsH/g+NT/PgoGekomi3tYgbtPKghJueayzKe
lWcRXJgAJJ/1Xwh6lfoYwh5ErRkLSccJqpbvjy4y8iLlhXqvIU+7ePHO6RyVzGsNrTbVqoBV7gaH
PJeSaO9Xp/yf7kP4njuivmXPRLryHRbNp2yEClUVA9zsUl198EKfeY4JPrrJqgnb59eXA4C4eW7E
chV4wkbsiuABx3sK+759wdJwQ7VZ/ljhl5V8ynHnLcn77uhyANFNt7k5LncWZE6A+gHXGmxHfzaa
oMzbUzm8rD/nheXrfbx5wJVbsf3cfPt8VoSWWkQ/2OaPu54CZmbC4NZ3ES+pE7FOTYlwCPsv81FQ
DBnf2OIU2R6w5F/qEKuB+5oPNTCND5TSTJmx9eWFpSIzeYayGD/UAfS/HL67PO+CPR4MoKw31F95
bHSYDtTkhfCDpUq5J89KxEOQd5e54XoZDcgqbVYwjIkDubp3/iAwaZSfLnFEuzh9Y+RXdSankXWH
BNf42bXabZzsMwAUVpydvzV+667N4dc/bTqOMJmgsufRU/UGVqAfmPlT0nG/wROSX9et86zNFpqR
uavETWv4De9ZGlPJSG+b0gEhEXfyoja7XDzWwR5Fn4Qcdn+jPD5Fn1rVFY2/cGDOpDGb5i3HabCx
EvBxnqbbqGi8zsxCQdUn88GM4wt3xdVf0t99UlJuQGVkpbRC9gn9BDgfMarZcSyEqSABJl2wu/VX
myO5lRzi9aPaN520xdWXaEnsm37my+SQXDz83fKOL0U+HgM7aJSDc97EGE0pEKPOOxQFmrjpKoJb
c17b7w/V/G88z/5TzDiMwNWRboFzCXXJIbFQAHa6VF5vRqM9iH2Tfqk1t+rG5kpUY4duHOVsheuL
8+nxzawS8yZX+/JIEazaOL+Xm8PPM7gDh+fUvNuCtKkfAm7pS0YNyN9Nsa+hhJeK35TcV10rBBGq
ZeKrFc9X2+2q40cKJKRtzpPZBex6Y6B3JG336QvTrjtstaJN3J7D4nDK1ufyj0+rU4JqWpnYuIFP
6/TH9PsfxwHGZsEMbxvKw5tQIbtW76Jf/iyOxZqmWlXzuMMJFdxDTLRO962vM0b7msPK/EGlyWYi
sDFqynBrAagyuUlBKpPqNGjPZR7GPEaDMo05EEzD0e0ILWvUs3/0PmLcFSMamkLLTQeU/uJmBCVv
4kXz3fub3azplRYKj4Rxj+m5hn/xB+O5Lop4IeoNAqAKaCnpzJPKhNrZ95RpKFJhiZZVJEDrIBJp
vEnIae/fdDejx3gYW5FpGAv0k3d+/gWd0rcrzfYA0KSwbARA8ZMY5oriS8BJgoJeKRcDbdPZYSjV
n7FzcLFyQjFtZ7HdUMLLJopJbM38/cideuSQTjjlDu5bU1FaA3DqMN+zTTtP3bdNO8Due9D0g0Xi
K94tjIXs5UootqYqpSTkVQJ+4GatmqzBGkM+UGmJUIsisuqkb4N9xyWpkqtCqPhM9KI55KN1VGcI
08qFMoVvTWqjvUHHSfMVK9fBfEVEp8IR3iPTQkfgdhuKUws9hAB8wfIbYg2uBLbv1xC80Fk9N+ph
GwSmiLUUQtbIX/KcTIM6N8ApyVihGuB/DceLQgO4laTLwc5jF3+CS3dNX6uW97hEOAv1Ob55foln
Vu23qTIjtHMFaJ1lXuXZ3ADBJMkCF9lpLGyRVNTnz/kuJMglGFx6er6SqqaR3gCG51xQ6jb8BBCt
z793bgkrn6b5ntITkdOhmJcYba1Doe7XLC/sHNdHH4u/iyeHGZX79w0dbENR09TfbohWpC2sMxtR
eT0FxIghxJoLBFmStOjtaJGmUukcNM4OUrkDt8OFmmtalh2muMEqgtcFsIU8+zmHN5pTywB29FDf
W8sKqDW9thyb9raNpHTQ7MjyXjetNKRX6ojAiGIw5AQa+xWALugpLd5LlrIcYalfGtDlMSED8rs6
Q3tW3suqrq23LBGNotaDVELRJyS608TLoBnIi1W0u41ebQTBE+b/S3DB4UuBkCeDzzCult+NE9EE
HiUwb4z3uhoND+zPvVrVZJpwQmt5bSDLVCckWqXfE0nsw6xkeDnK+6U0mzibOjgqJunLPfXw3PRa
Xa39oeNNeQrLmbvKnqwiSa8fQT+GiJc18wnvplWtOTEzm//Mo1qexFZGJlMRVyJU8fhgCFTfJK9G
GJiZNfG9cPyzFwX5jWk9cv6wSfXtBA0yquSBeb5qyQ4SnQCeXTKMQbccQjZSN2uwEikHZ53UV+We
jCGdemfHEZmTVITc9jgDoieQlp7OLQ4JuukxjXzlVJyKNMByV2f2n91zwAssb5R5aHPGvzTfSjAV
rqCDkbn5r5XqgwmGi01Pp9hzmGWNLkNiOvH6wvOBNhXeB/LBKHtD+oU3g3bINK9/jnEnyc6Bmny7
ZCEFErT2ueUxPJyjztLGuD7v63DQLqAcFFKgXaA5tGXPvnathAtSMnM7uulmuBpuoOZRekfjBsQT
rIidzYUWxH6s0QrJGOHm7PrN4zl2lkKsXIX8J5sBzCd/jyH3XKFtPhjkbPa1/btJp76wTwZyVpjL
VZMJtf98PC7hR9ibABG+UIxevPAj63cq6RaMgh0uwqbqv+DzpShknikJiZu4PUe5dvRN6r5hz27H
OSf7SQKQeaKQG6YiiWwYHl+Y05IzB9jCEcNtD2d40j+Puv47BmRl49GALhN1ZS19zGaPJQKIi/ys
LoLW49LlPM5YG63VBM6M0T+1pxCWZT1tiz8WT1K34xmJh6SgphfxCgABUxLBXRRhMSg98aoDq25v
gbu3px+FJ9BEfPwa8O+7rUmeuVO3FwiUmgxEiE8103odOVFiXymE48YDbK40NaC1L4sV+SHwK6ai
UmHmkRXg5P4fRtQgya4U1c2OSXoJRhqAtVBPVo1Xb6B16tEfXrDDmDN7ZkoZ4eOCZGwk01ReCRCm
LfXw3qu8pjzvpX7UVepoHNZBlWLZJo7ky22oDlN+lI6ci4DUTdXj0EoqNnHztHyXmmAdCX0wsMWj
fnavsb416SHAGSi3I4E1LNbUGKCXQzVoNALfUKVR6UFOlwzURtufoDVxnevNFMXqStDnc3i8LLb2
GZ2nufV8v6PlRgOvQsdqIRf9HJWTWdWEPuBcSOLJ2VBXbQXWQy49weSqoyiXl1/v75o+qM0cBJWB
xgXu/qtDXLOFe6cYrPKgXtr5cu9F9pcMi/fIE7revDaJVUOfPX8Ew/NdQU9xgXP1gYwvrD6l91xo
N0FYsaHIBDdSfVVGv6uc5eQki9e2OzdPe5NQIdZHsnCnEyIY3dgRTSlseP0wA6bGZqSij9onEtOZ
wyhUhb4fQcfSdZv58AusLFGf5DoOGmr68D6y1EVAKUzIOyhjUmFNiY3CXZN365bMC85aUznMlkFH
IIBHhqFVI3izpgp2OEFin1BRvkvIE8Fz2HSFbQlkWgSysUWIcQwTNIpTLRHuwkFdZxkTniQIjWlT
R3UXJUPxQTlkmXoxlmddgL3K11UWaTtQoSTyqYPTsD65nqa+H/jN4bKnv4mJnSG26OoDmyiMGWXj
gxFy842bLi1sVyNK6oFJf6aTeVRtNTgxP4eRnb16WTX+Q1gYKVO/kKU4dyECJjzfPWhvZsBBxgTO
0E6ewYGv/BIlArPGoEmE14Pfx4kUy91uNKXZ85x4ByPG/HdaxJu9rzzVbd/r4RQuKw/wEUq+S4vd
dKEaM5ig/HMQzHfL69NuMKXCryDitUQADjDQEhIUo0+QzhrsDIMphn3lbTOvl2yol7nVS4PhoYr8
JAHPx+YwjbasQBwzrmN8pnIvLeicZ4JIjNFEqIpTLQsVgPd9usHeq+KRSfyEMcfepefRg5ly20zh
O68iVzpNB+ZmoY4LHaf4hWRaIKQuM/QC/zlBf6zN3JEThhCB/9J0qRYtS8fMtsnDEqjUzgPyf15V
CHpVRjGdmiY+r5f8IhcvQvR2v3l7g6HqyZGqxDJRWqiu2XV5IyaosKSkhG1J4VPPNrO6V7MGDek3
2CaGrr0XNvLqlE/eXhXV5QK3JWfTvUl4kDNtpL0sAXfopWPgRo6u4hH+XVOwDh1KwRlQnCMaMoK+
XPUIKT1+XhH+Jeh1vgnaCb38rZPI9vapTv6+lvdVRiGl1RlXCaHmYyM8Wx37AAbC2TlAMjPmtCwW
4Vwjeha1n/ACCMbU43eXkW3fkpJcXh7og+LFEiofVLcL9fS0zuL4jT4/gvVVveYXcmvt3hUSO5AT
x+UASHArn3VcGggQN9JGC1xfVM7dtbVsENYvfuSBi8977RzwmbhXQnFtcGo/T0nQXo/Gj9Q+usmi
K7Ef9F/VRJmCIXJyuP94DJvO116o0A2Tdl0boXjC6/XqFM0v0KJ5KLrGxqJkIEP9O8MyhXMBQ7by
wgDwKAezXnqyLIlHZIZTdBzz0wW2W0vO/Ert4h0sseUHEEk5Vlf/i0ZL6yJX4RO7LCxMVT9O4zgO
gHO5eTg/1tSdFLKkBeANa04vpS91XSveFx3iie63Zu27YwuKbI8jDox26Netp7WloqujEcx6ISSf
3hBYF24YUHc4UEm03rEZ3OwND3BecrJ+4K4v/1dxUeVY91Z1tkQ6ibHLQj4mk7WSXxiaudsQNjjO
QLYaZW/luqqPkFYou9GhbV9wLqx835s5hEOwqNrs+iGVn0Imr+fV1mN25MYcdI6aeKjodCAtexJ1
PDgzMQQg/MTphuZoNT/HwqGYHxVZ17wW7qNBkbl626/AGCuxXSzN8Sd4/5yvR8Fq9tKOoysyLpKO
cMFtSPuSP88YUUQXOPjfaA+OpkGMeTxM4O1M5ZRP/ULN+s3lAFzBywPWO9ULOKB60derTDsf74rK
IoZsm30hMTCvHkrGxiKBiRD82Y97kWHgespMUsH+ExRYx+GV2vkxAqW/fEuFe2ZEpYhZ6kmuPuL1
lyJ9GJKggefkKAzNNlSpYlI8QrBT3nMW/nmc5XhsVDvxxj1by0tUOrYRsfMhb/Cqjgr784WFORWg
AeqXX1zmLAkrIWN4a2rXhvncF6f2hbC4xKX2nTwDlqvWsmh+pJ/XSNdalRT0b9jYW5EuZVS46Rjg
13cz8qUBx2nu8IrwMHcsfTDhQ/S92o0tfdirniZYLI7r78dF7z0dcogHeO6kS21juhy8GhJdJKJL
SNqtO75PeQtlxO5fDmdWzPaSHRXr3DlfGSSZhthaFYGSKO0p8IBQasG9cPrGHffzTpyEsiW+GKi4
QGHZbehbmEi/Ccq9hCKmFWN0MFfIanKKK/aKrh2idMxL11LWbwI1s3yFwgSA1DxQqyc6ow/Crkum
HnvvTdkCMXKnHrXQ1t2tWC8ho+whpP0+enegKr0NiKsD6O0OHorsUo7Y1OF5NR3OGrF9R4hkJSnL
huq8jrtOmvQL393pDjwtO0iZmK4GKVn1jyCuSSFqlPe2kNUEsGjcYk4nQPHvjGhaSMvATa8aoXj5
XDXZWfkJo4krUtzv5YsEXgHpvfd8UXnpIZDgYqn1PFhlzHRO3OJ+lMPPxIFu/7WiMPcwGmO7IY39
gZNiiBS4ndLE+zRUY+lw6xJKUqeElqOO28t5iX8UV6aURswD0TkFH2LJJRDrrSvEh5MwnY+Qtq12
3Y9dPB9NdZ6XsmnE9SAR3cUsm/Nt+1ytPuGvwrCMc0iI5v1wlQ07zMIJmjR5bHPaQ5GbF3oZD4GS
IuR+7+74fYZdlNmBTpjxXS6RXJ7a/iSOOVxsUQpONJXpd1rCJIhKNempacCpcXdmT1syw0efqMco
VcIR5LZRSfzo0NT7MOxD+japXkTbOvCP2CwOtw4eq77K8h5l2qXpo2GTgBsTX81TZIHbQ0kyk0Xn
Hs7gtF3wUFfvsJsWUzp5ZQL21cQ7y9ZeQjNIiblnqVV2hqQV4XLstzh4848Acu8cbFhmEqmh3XRX
PhiY7wRNKuIygeNDYaj1Fv1z0jxBZzh62xuCcvQBxwwtNGAdL67g9pgxu3RQ9hdlXx1ri30GFw9K
RWCfoO6b/pjKjV4uQmrN24Q5iDx5aur3nd3l+Rygun8XNPvzQxGmofu+zpQNakO6FVnae6SEcW3K
a2RzixO18GCEp7qXQtdpAlgyaJjW/HypttKihF/U1VdxDVCrTJEyw5ouGCNObkjppEbaNxKkr7ul
vdeYYMEBcCUQIYxpe0YFpQtnDX/uu8joMaUYBIptmNUwCn8zQQ33+N84irSM6OcVJ/3ZzzfUikdc
qh/a4wuWelht1pqM+CFHPUlxWQOIhwUfxx8mqbEEX74a19fkfXu/a5TOwvm1R583mBM6MvD5Nati
7k0LrNwIpeE77fon2hvGNDFWZZTyfGRGicIuYCvgtRwRxNjo3jEAGXnfU6tnUd0av67rA1Qr3j4+
eMLoXVI1mCK8eKDDoJS8ryQquUn8F+KxI5eTs9WIEZfrFa5HnFfqVuXqrxN6YipxZ7GjClOjrM78
Ovtezi0CEo7e8vvh5nZEJSnu2l6kOd9lK+PkSMHTqwEzLu8oh2CAkH+LJKzO1+NiqzHsXCieLjzf
Jp6mSNxxxKxToJVj8Jfh3s/5IgIea1UEPgokTFwtlOXlwnNFwg9X18s0MsN0/SuFN4RVSqAeLkH/
pklbxgcY6AarKMLVRrkQjAdoa25hnxy7k52gMepxYUwS4Iy4Wv/MYEc3cgA9mLPSCbwcpHrV+tT6
WGE1ol+NdIkYuRQKVKhEfVSQfCy8EnRG9N96qQKITQSs0nLdu37zXC6DQe7HlvmzqaAORbecrAOv
QTFlumHIR/ykNABycMjMiQDuM8bRwI0Tj7wzXOPbitYiEkkXEzQX4fFNMRak5thfD9fQ4xQJRhd9
+RjqcT1uoiC6LDlB4L2qYb5BRN+tJInbwfESC8qWEjK4b9IAlW1KHOTCJamafP4ifjGQ6KuinsV6
ohSrgtIKfTBatOhkiwFGH/r0le7pLIywLu38v+SB4E8iDwV5vlH+d0kF14tDBuGQUUgvd/cUjcAR
yDooJKCqIV+SSZDSuECaLQwx5p98SboZJrP1QYmRjGUvSlPfEb2wqWpprY/2fzgJLPtqKwg8OqdC
M7sc6Ujt3Kxw7NfxoDqe854Ikmxtc+UqR1w6gRS8mPddULStSIK/JNZDCy9CU7nj1Lwhsd5UG+Gk
2l/gDm73r45ItAnQY90qrZZlO7VfuWPIzC02yV6WvOjc0Aj0E9w55MmskAShdCqufSpMUuAoYWWp
SmA6s12w1FOq9i1gzNt1CWtix8o/LAu3cCgym8hY/XwT2Fo/gms6WjDle5Uo2denR18wYHXWcsa8
6ScJmQhMlMWNbDNuSfi2/r0DeWkh+QxcCCExWPuk0P3dsR/GLdsPumCd+ZefpFGZl3Qs6j3DlYi+
y2xtXjzyUGF2afZBWtaP8evhMwL40qROZPW00KtugqyunNDowUpkpXf3WTn7jbLzxU68mEki8Eud
TVVxwnYUccu5/U1HUKRLgY6qZJ0unPvOGK8RW1T3AyQpMTZvTAJliK6Y2VjZ1ZK1Q7j6H90hdYGJ
dQ/eTKZ+EHuHtKXxu7t2VxGF9mNQP3ly+wEgSOF7R0RfNxQkFriJXUlGKQORl131ehIIVWnoFVcp
UgrQp3jN6XZLrMcRlzmCoX0NvzkDPR73NE5i4aNrEVf5QD12zlQLkdwQBL6Veeisot+s5Z4A4I4c
oi357lHq0ovbiXZf3G68ArBx2pbUcbobIeogLYTxhmpueIru5P5QkgagtK4vyXBY+IcpR9ZR/RnL
rO4gY6O9k1Ezvod+r66A02FfowYJo1cKj9hTcz5SDJHdObKwiHSRrpVD7JZBC0Vo9vVYJrCFls1C
+bBRMiBuLpuvCYswOksAxJctbYKBIFBj5IxwEsUqUUKc2wQhMPQntmMJ3HBVfX9MeBDT1MYDWUWw
zp9FRit0OT/e9C1rsk6Xpe6Fu8SymcgeC+7L24xtVf8ijJQndgyMGQgOx0WmIT9Nm64rBJmmAcBa
JoEmxvM7oZ3v//SJ+4PKUxvMjlAwOxGIUBlHNITByZZFwkNpBuUZDMgG75DC4yZ3LJuVaVVDFB4e
trEskpauPA0IZLs4U5Sj6o7nFMybtfcwN8Vow8tQUDLnaye+y1ESave4JS04JgPr4GW9NmpwlXmR
UfmJTh1m6Y9SR+JNBgIoCUkzsQ1L9/bv79Iu64cQ+eDMs2D4kn9JH+M40XTbw/bVBuvD+ljDjYDO
4ie7VVyG2hds4IEadfYfrtHLKYVUn+nijlyHOycI3tKJnZriMG2yjN8vOT4mOFO+tpEhXIFohYbc
Q38w18KgS6iFWaTIBYTB5kwVR5+mVam2SHAg+gN04RKj1HU6+CDjOL6SeK8sB4ro6bFln9Sm3ZBZ
IJMOya5RKE1z5STgI/n/7N7fUbBMgBKZYuppYkE/tBdvcov79sXEt6R8p/YLYe/0VMLGyJTQBejU
7a8mP8cmPKVqK3hQQOgOIOghdoPN1rD4D8JldqkBQVF2is8lcQjUFGRgkP3tdmgGNce+P7agjmPK
IOU6I3kmakFPTopUNfOO+/LsHYB+69JHIkjo3AtB59qHCP8Wcv1qk0rhl5z7GBSXKA3HOaA2790B
cWGjGzKcBr5XZRYxp7hNsN4Qn8/1nQpBj/yhOfCLD9bXdcpDyo5ja/9rPC8yZYP0jqRxG2rFQZZC
W9lcJau8h9w0iPNcKlD7f8m/YxZlrSj5wRmzHoslmDYUuV4JTksuG6JngWOpUVaazoa6/E5hwJgw
W+sa+XV92UDgaKaknzJ6w0utBnQ2f/svc2QNzkjH1APF4LQS1av8rI/QYnVJkSOcEVCKUI2yVhAP
i1H4mkJhh5WwCvh3joFwuLnAgratqlxCULB3UcBQLGekPquyA4euWuxdYbrVIXMkNJcBedtYdEar
Edi9a5mHrCBt+dGtTr5FsSpd0hwS3m+D5a1CvXJhDXSaOKhqzWDS8LdHozZSV+XIM+pqSJyn4YEK
C+Xjc3eEpH0oMUM5B97tlbnewXUCkpL8SNtDJF+1VxQ2NSvOQIU1YgL5ouZSdotVsN63YK9b8C37
oLt7KDR9/Y6aDditDDf5AjToO4u7Pqsky2rLNfzLXlt++06gz3WbCrI2mzZe9svvweYetsFqbcm8
oZoK76cXhtxBgWppz2eaK+tqR7ruEdBhPLQTHE/45AgeV8cauPURKbV33vyKCWw31tABi8sEKsMT
x8FhutNWLl/LG22UpEQbNvo1S3Ms5RGkyFIoDHETz9OVO6uMiyfHVkablSafU2Yj37z87WTCjrub
fMoPYpwQgkSGSOV5VIZ14uAYP18b3J/DxIRtLqnTLA6M/tzWJb3LSnfGAhEtbM6cqbznGe2hxD2c
03/sNrAC/3YtfjUDZb8RPg813gMp+XT0IwVWAbQpQu8IWxynD4UU2Wkpm6gCUWDsx6MM8akXyI3r
6WQ76FpEWNDTkuET4DrZVXzw8429BNhVyWsBljr7l/Gxisy1Yr92CIx9UaVbUMMNPyIs9U02Bued
nm/g+OgaZeJSDDRgBRwvpvT95escftRuyUmLXbCKXHcbxAlH3WA9JHMqRUgCEgbo83FIky5xOxjF
OzsMbTEsYste6RJ/zDytPGMlVWFV3diOW6A0voOpPXfUrOFue5EcTj6ftfEBR5ekU7BZJvFobBvb
vkIblFzd8jrZBAvF8vO1bfNRkekRUfcn8DGcbC9STyf6K8RWEcRHLdMTvcLCtP33cvYEUxGpDMBG
0AGlxusx64hVD1+h1/49osqos+8OuEIYEKFCR9DhZsGkzQ5y3RSbD/QtBTRUXt3eaivsmk9+sUjs
PIjY6IxSgjvxDly7CjJiBhBjrUWGkS7uOcz+O0hX1nJTmnFVI4iM2ADA/goU0UVkDrSTo45AUywY
zGtaFdRt8v1uLXNFxh1nWmZCG8i+J7v3/5csLNoRe/uJ+vOgw5Qs3imn7lnumLqBtiQAzg7N0wqm
vIXsXmLNeJDAX7ygxawvMJjWSmO8Ph4MtWZ15nIMAAymk3QcnBJNSnVnePKK864o0jKXH51ArDnQ
IuPMzgVKBSoBr8PuO0RJ1PVywMdiWhOJsDGjM52u9nrf2zZ7Yf9LRVmT76oL0X9uo0LpOCf3+Iox
o85PtQIo5pdgFJ90qWTnY2dB+WNGriZqTPXf0oAKGFYPrpEAdsVqpEXhYS+AcrvL3gLdF5AhwuSS
6k4Lyy8GVArXI6v8abZ93NPGbH2KRHcGAc2qNSIlU3rGSgV58sxE3okFgfSlXR7x5keJ648q+0t5
kfZkrAIYb7UeXIvKyfoc/k6z6iSK42X3CdsBcKJW3bQBHQiItaB+pzdGnP0N1iwOtxCJkR7IiqC4
stVdbpwnXt8EsC/wmAA+tCx3ZlzuDVy9WFYapzmhfdiZPySDPCC7XGHDPe1/pWi2w9oO1CD9e5HO
x5Nl4hAWECZr5LbID4RsbMWaVvzckwWV65wV8n2M3+/zwwEoGPmM3IKP+CUOzau+ZPEDqrIJaDTC
Fb9XhjHYyjdjVBRIbcO2k3d+KMvNlZT01h8qqn9D6hyR0bKYUhlfAEiMML/0Huaorz0Bx/EL33QI
8nmIMuQgOZ3smUTzoP/Wmbfely4T41xgsJHUFRrqSn+OSohveEGsd1e6BCCLlUN7yqfqIyAOr9ps
GeKYe/FTXpJFNMhB+q1rnOzQyao3Kb46dvwWyT1IGtAAny9MJY88+htSReHzav7UtVN5h723gwTQ
U5C6avUg2gXI9nAumOvO3nIhjiE+SBgdFwaMOLT7Uj8QO+gIklDRKWzTfsx9ZosgPfS2K2WDdsnR
Q3bOs22NnAN/z/A+3cAqRO4QdMxOeF0aWRRYtkkeGI5W+2yGgFupEXVsFIwRecNZ4/TgjNQH+od7
45V+cwjIGUS8/KG9oZoJ6gUlbSzk1k0P5oFusiOmFO8J/rR0YgJliCRM7dfkYqeCNTpiozjY3dID
DwT9EGQHE71lvlFNkk9IHISF9IGoOKPb6Kkqjiwvyb0OpBhqH9GEN2H3WGK6Dyjtjyaw/Z1P+rWn
6h+i0hILb5cQGUwOuu7+Uf24DFvBajz/ymFuanYoUiww6MJcgLpb3VXUSrOR0+CtGORChBj3fKAN
ri1n2lo9YsJGzUCLWYhtakMdDLsus0hxWYylPCvMBFpWRPUuj91NHokSjLeR4lv8zH5HKa+MYnfL
+BEk5lQKIW1vBf5mmIEv46DaOroRK3MwyhweN9xdKbgILjRYpwM6lNLDwb7536Ypuge20pLTw3XJ
0pLuYJyptJFWsQRk9dn6FfxbB/cKom64WbCZZXRyu8enFsaJCL5YDaywUN2s3wHOcbZV6tn8MR0Z
fUjA4+ME14mCMtI21PsZe1fO3xA8HffuQC6s4IvVKnLj4UZoX34Tcgo+IFJLgNleLBiEVXqlKumU
nMIoVeJBqzkjLn73rMGxAUjJ8rIAHZ8+zKTNTZwp8cMpzJ3YlTXgaBlpshdVuelB5QzwEtmtpMO0
sSg8V+DPMWTldpdYlyqg91/93h9VHthge8H3BPFLIo+/Zr54Ekqz5o8aSfgOYFThJ9IhL1ujK2Lq
KfoA6vmyUhKg47hR4+O/ufaIbWToF+IBBInNRXADGQ/9+VOTXUSUZF1xGn6Fa+mS0Dj+OwbgBaOC
zEyVtkQYlCjR+FPUBVt+vWlM2toRY1e39Y26g8D7W89Chi64DCjFUbKGWWeC+xGiOotK+JwTcbXi
AwWSgth6Vc0LTBMaiaXdbbYZ4JWKtpJoBcATjLyDNG+0IeyAJmbBuyuhLJICzrokSzvsPCkKqxek
fzlY9tiI82A0bUXybaJ16KwlIKyfA8NQrx29yxp99fp0/OX23eSt0N8oQdvRz5B+yLT3U/V4umgX
08MjZVEFI5ULZvU3BlTtaYTEw+2z/5KcMnNepNrJ7c5Wj9JyKtPJ0ygjyZMg0kyD0shl/rfZvDyo
m03l84vohaoW/uVNR5A39xm8ik5xcE+/Kz8slLAp6imVbgd0JRrSD3QZaYJ661AyqdFGYvkkFm6L
ZCutkddd+bBqPnsLyq8vgmdez3k3/6CBpYNbj3anKeerQIOXE8LkOdrAautiObjEwHGdItDC529N
WEGtg8orhr+j/tVoqbFUstXQewn8oN7SPyWhKXC381aCRCWjy4uoPI1cCPQd2dIvPOdhDHCUauSd
HPbctlazjLcMAkcz/hqb3TXJXTuhqgqWWXyJZ4ZnYRAgTJpovg5AzgxiaCIc1JRPetfWWl2wIdM9
eM2hQ6gDWcz2KDNWX/gyUuj/2arWvUeA+cysssc649+bp1KmXUixbsKkgw09Zr5jqXfzGL2ARLzj
R/OH878bTbH4GI7Gw3iSvI0Yv1ND/SaGOjmE/YXGpOZit764nONgJEhis9tjQwcIsA7ALJ7fmKQ3
92/wtXQZRAJf3hJYAGy58T64huRNzJ+cALByHGyT7iU4LqmvHWyyTm2EqLLkyld8sK1m4FOSnwWl
dG7Te+5KGNhH/Kc04uMRyz9Vjv90b0LR2slQY+LEdYK/Ngtyb6rCFLqgPtCqVw3LRRdxS4pyY5ic
vc1FKGi7uE9CvK9Gh0cN8QWRwpTWc8Vj3QXueInC9Vk30YLNwAOqY8jZfX3tpTJShPdcdsRR0bBk
sTc44rPwYtZGBr4mBwLlYAiFsJddmflBvpLbdlfNLd/Q4FVK7uPO2ivnG9wNS68daBCwWWOitu92
moDSdoy7kmlC9W2Ja7/W491Gj1vFPEef5snF3vSxw7Z54DLiOB95x/3wvMAeiWUfL4ETbM0ce9hd
Lw+emJuyCDlG1hk5SoQLAT1x8tKD8J+Fil+F62NgMxMCl6sy8IvhZsLz0DVZEA59FU7XYhmVdBvF
3f+gShzYAfP999/CyH4KEa+4IpXyPicD32CIHMenDpj2/diSUH2pH5oJC8ERu4z0pGJ/KH6mbE4Y
UsUtymXYpym7AYLpB7knvj+3LMyeFboNt0ZHB3aTuyjhM0hUzrjl6cTlByc036fqSYFneR5FlOj1
D8hyrOn7pJgDFNLWeG3N2B/snOvtwrUcU405B59OR+7IFvWhCXDSxl8RJ91+t153fhdn5J/oVpGu
ZqfZs8SU/v40RZpT8sclwQ+k2KnTXoQjl2L6Ljf4/Yua7dyf+e46UwMg2eMohpuIVaWDDXwLiiLG
5sn4H6RkRh5oZ/AXn9IWrtMSESa2e3PqMdBK2GiG9jcRx9fpICvyPigB9so5g5xLqBTvOPNSuQqZ
g0P3L0qyRmt7Y3/uLHCzI7aCZ3rnYPFnajmfbAg1tqX/H6Hdc2wuG46GTmfiZifvzxd8bGi7QRcX
9rX7HeXqCHazT93adwG3/EYSLXIW/0y/VbubXcjfBXwzRhqKEypnHUDPJOb0k5fIQOGP9DYmwjsV
l3AXoiTmo6zangEwapwLGYgtOpcgvPxP17bziNxPGFGqDqrUfxv8SEkHti+nLLh0CuAaLgmhCA1A
IBqD3TB7GMaBtEmLda+8eydh0jInz37ljpPi0t3o7Na2OlKnkQMA8BdiagLpUUAde2Ds+GlH9003
PaLPND3QDgtYcqyuyxra3DvjeEi+Y5SdF0+b1bhnthyMF65UgTEINdFZ/LpmoKkTOjo2pLBsPehy
NaPB/0v1G8vpFV0CfPWD+YYCyod2Xo+MlPu9CznBYclx9eN4P6eJUlTz6f0C8W3RAQ1Nh/wVXnNt
EbT7il+5PREKMHsFzCQNeFvuDXWxKnrqhthpL+ZfPmV34KLaGljfd0jAfV7n3k0uvlbcTailHl0n
XFTQl9pSyw4KkDUirL0EkAZZ057FYCc/I0Q0OhxJDU4oSgFKllv8CmoCM2s59FN4UyYhgvBskp07
6VkvH0T36CdlZH4usOD2AHDGbQkhLb7cAX0lhogLn4yeAmExwbFb553NzTNdKn9EA6RWH30/2G3s
OB71OlwNcC6smjLQTv/+RjqlTEPfwW5fyLbsLQM6IUcuc7guMvWduJAxyP34xz8AQLdQNfD7NIST
JkB6ePsAU8blRvjxAFvmhu7cDso6MTGv/Jq9JYfAzw4NPNja+Z0+OzvefGXU2D7zl5Y9Vs5Qvf/y
0gIAx1QQtEqO+xEt83hefH2iPuN2TjOg+sS7MGPZJBX+ctZaaD9W6y/g3KCnaNTE/PWQewkDy+BD
fu+fCXzXv7+Gqppl6HEPGVUeH0dYUbXaUPNiUGK0S/04HZK+5n14QTIVFmAsootK+rtwdkx95C0k
VXkZ4Eq254c+LSkD1n6Ihzaln7VB43IhHQk/fI6g+OOarSZb5HxdvrGptX+tzAGj7FOiYFVtb2AF
E8cTZ2iCXR0MFxGOx/sR9BmPXx0cHDKLYtM8/BH70cWUn/Mf1uecOZk7OM88BHGaxXfk3V7I0AQl
SXux+hAH904n9Alo61BDlKsA0zTmt1DyZljaU7ca4Ptw3xciQalBs68HFjy25D9BF8Pv+kMqISJh
2PzTVoPIaKRGNqwY+xEzzZeG4o4kURavZGF56PCQ8TWcg1uPDQsNgWB4q2Ka9Mq7zbB6K4Zwyl3+
hS1Mo8piOG4FicolsSCYuoIgy6taHsbzEXnUBNMiwZ4tWlPy+dg9eH6XKLPxBsa7d3VTYgFKjrnk
tyoemsOCyB/Vi2JNzfKiewyeCiNQn5Gx5+dEIqexlnj6/zXnlEPKfbdtcXsmrXw6vG8r3jxXu2Nd
cUeGtdqeYXlwHUcanZ2mgczOdBIh/P1Gj23OEKmlTWQW49Iz2RGQpugEIb0TMISC7lUde3PV35dq
Jgxb8tc2TS++CwAkLzzhcbly6WRPreNbDvtSi/EPnU6ar/7BBhKM4yvfWkaYIpif/S25ZFaPNAhV
LHKMn+HkAaeat0Rm+6qmfQglxbmIbwnAOOAEsZFp+dhpWuF6YYhomPBUTAByzXgQ0/aJZ1UOfgVB
Kipsd/rSLXdsDjgp4oLeJ294MsZsFdkzapZLarcEXMLWGrxUiDvy+cJe8Z40Ggrb9h6mTxB4xcYb
ejZtWJ4E3juMzIm64LCPYwUuZMwWrk9HPuKkwMCOBOZi9CdJFFM623GMw4taoDeIMKZOcq9m6rJm
6v1F6qqQYvigJcCXBF3RLqf6PXR5Pb8/45BqpcTUbZjsIQkJk+QfreZ2ahBW863e6EaNKKIiQBHt
+v4OwMzlemihGDLjIcncxJ1OOWT23/2l8LWzBEJl2rZEPjkXudbJgRoF+TuR20j7Weh8mn4qEm1S
OUu+9bjKg/I5KfEfMvHg3JHlgJA0JAOeY9WnrjPO5ncBtM4KFSpkhSoWg1lAWu6u4kZYW8KIEYiG
9iSWncObB6lbdsSELraX+gZdKzgSdYQDGBVjIRBgvKu/vhW3Gkj7Q/MBMe8KI4XmbcdibQrV7p64
6+MQmPUSSsJgt1cv4QF3w6rHD6Xjt2yTRy8RntLZDKzlsMDZQ7GDSXxqxuM3XelIpo11NU3VPIzk
hjXx8pCqQq0RBnwFWniXotS9se1TM4Zn/ZJ0TamR82Ge6lNn7Y1zXqpM5KSfM7vziCcLRQgDz33J
Lu7x3hUN4SCPlBK63yOCQNrcPkdFlLVALoYK/GCEgjSXw4Eb9XpZP7DOioHysu2qOq7eKvxkE2CX
JgMr3p/vM8UY61C9KcyPfmQs9gnKFQ98gKu2YzYuo9nlXtExXSugotjru2OoH/EEMeFvmkXrmWLs
1LcyLBis9rteibFwoYMATgDICOx7xfIRnH21fdGtYFVS6vJPV63pGQscHsM9KBMqWWPEQFb/VMFl
fRr1mokU5ANw5hQan/5XQ6mrt3uUE3aYNvmwJoOLl8jXAJCBMw8K0YuKyT1IfzRFvMadhNwp8ULL
r/KG0sN9fAXDNoE1ZGyvJRpQeqrHGO1pELrLMfcE22hE+RN91juOIIXiwkh8J+1JrYhHABI3v0qO
FQ1pa1+WShThEtQRZjZOvz07I39fiScZZmkLhZPwjSSJUJG/YMadlb/e+416iOwmBN4055XkOoIZ
q2zw0WrxtSvt9hMsrF4TbSTVofVcETBLcNby5aN7685v/Qb6mv4K1svwwxZwa4df8d7p/gBxZH6K
57Xe4Ky29XuPmY80cB3WYew/qqc2iUukcMbFRCXJA/4Pi7M4KpSO720JzKP9vgAVZJzivc6PJbW4
ChHjv4EVZbx4frCNXP3PC52zVDzXmrG7SO6jt0zP3QnrB2yEPxIR6nXsWXrnQShDJsVISp8McTP+
hQSc6/I9QW1uqYEB4Cp5ztJRgn7DYMZ3d/Oa1BcHItLt7fWH2RC4+y/0fHC7sJbXPrtd4oBns/+a
1qLOKz+Mh2twIJkAvyAepFiSRtYMGVbcddh2Nx6C7MczqQPPRvW55c4FNfNxxsXY5zl0DVRb3zaX
WCZ+DxCXJRMD7vNw+07iFH/j0eOGg4fTXV2lkwbZ9d6aZ6NftM3tc/CzJ/U89NOkdqRE6zLMqwea
D2wd9nHyS93D5f0qq0dS51cxX1O95hHS4NGBlUxCx8ym41YSBzB64eraNWNtvz8DQi6fPmC2dq2m
rSdQa+Pom7OdS6cOeXA8rbyN7zqGhtaJdrVx04ikMPdsnPLP9EXfr8iXK7hXsA32/h4Cqf4qMY+o
gHizfYI7CRhNzrPZgiIqInn6fYqmFxi2Ub7PHCzaJiWDmU80C6lcoClIoh4aXyv/I52JcRBujNMy
B1u7HgO9HsFZQ3TTCf4mc9pVOAZQfDY1uSyViBNvSYzsoQM10zVfAZotqAkycZn+Ft6yee7OEhc7
BJ4NuEk3N6SGxllr9FuE/X3Ied6N0CjGrKi+4Uzzbo0j58CM1Xz67GRqPm8gxDvXVk0DW0xIVp7u
+vWldvZ3y1SIufL6YqnNtFA4j7wt/dYcvxXwPuH9mmiV/TQUo9b5rpuV8Z0LKiRhDPqlgJQ0AHSv
s4rZuhqlp247l+/oqO6AmTQ3R5kAFzKK+KCw6sR4Wd/9i2nzwmXazUUKDNkkrS3NPEJWCC+UpU0w
V5UJbpVsP869lFaZdrLOIFPgRV89hLE2jORy4PYlQhc61E1W2Ydp9ylMCdj11wC8SzKriJi4sESi
syhkRYhf5G60NXcsHi9nxJ6d4mPd04c32ExZFxIbpvfI2K+oRPkPolqVU5LE3X011C2ka0QR9dQ+
rZDXKqt+tNb0b34N1ouYoQ677/4dWD7tILRGvOqasQ96kuS0Kbm7TeLlvd5abGC/HcNMCGK5mMfH
PMp3zAgH40NIik9y9e7WEjRIFtrIBOnKclhv3+gXms7oYia43PVju15vpccVbb2lNnEa+0xqT7ZK
dri98XTgXlJV9tfTnXyFVdJCkBJPzoZFL5uy67BJt8cSOJCQrG/Ra/5uCJZ6s0Mmxo4p/mrPu9Ji
n8uydRUAaQfs7jEn/BOLTfu4mnR298RXWFn+9qyFiydwYJu1K1AIDkUCzy2itZNY8bk1MSCpBebN
tnOgvJoXtzDyX382sVn3W3MypMZzFVP+S+YI3gzGHnDFl5fSGHb3QbjOZzFmalgFFOzsCDCaxzEC
ZDeCFtKwgZu+NwVoYwN0z0IC5kpl8wOWv/+w5KCbW11BNIF3JMR/r0fPGxDnPtmq+7+s6BJGB71k
ruL3JCag/7gPZgCwYsg8EPGZrlLNd0dAHFStT+ljV6vSRPPITOQbbIg4xNUnFO5D3lR4SsVhRMDf
cJeICRZ5G0uncJJKY+Sny5gAIF+wlVqhsXLJ5EuZ91o4lg8xw9OEH9FMqiqaLZwJBY/LYlSv44Oa
giXRDHgITprZaA6vlzYeIOZCBngaXyVAtevjF9G2G6TiqR7SDcQ8Vz93MhyNzxyNyNZXFae7jQM6
MXtJGkHX/QxDwlGI9Jr7rVqSYuHP8kd7Ck7itc6K7XC64/akuTxBuwHBaES/dPc+5CisxnWSX6MQ
J8kV5qK5mtZxH//W/r4E0W0OaGwiBtdS71hOt0c+2ifuSBgCSrAT5s9Y/Bzjn3TrKw9vAPHbxY39
JrMZNix44SCZ6tydBwsyPsxo3uemagn2hI15pdpXNaJK4v5j62BaEpqnvvKW/wMTKLT9SWTxZOeO
lCp/Sup608cG5Ujm0WkWVU6iCgTiQAxXvRwkKafXfZ3jgnQ/63v6flydsWcsxrBfVlKndNZ2iZHk
AYfd4TzqCgtNCjssTQB/9S/If/j/mgZNd/1Ophxf2FdNh8HTROXOatTCSNzKP6s6fcsu9BBbhI51
id+cQ1DUl3EP6iSPAOwaY3fJ7uxpoJsuXMKcSpluNNHfWNwHPkWxscoLUXXoQaacnYiDCMdoc11v
5J2UcCbu3Tm7sJ+9zzSABvwYOJqTdBh4+SJ6Irkoj8E/ErxRxYGJ3XGcL0toLIAVTf1uiw3+zjV0
ioaGjZeTNRp1u7jrsm1TK8MJ1LnRQJydiG5SBClMsN66NwQ1pkyI8jwc1c3XTyfn9dLNRHKegplj
1Gfo7/HbYwq6WWYIUiAUPE/K9AFFBgpuA4h9BTANbdvpKybb6QFRneFibnTjr+K87OjMTPRnbLXS
slp1t8h9lnib3c7VvlCqyW+yJQCFkzXf6RZU+9EHz3TOux0MgtQMJKTz4pN15g2RNAd1y5RrV70i
H268D98tivA4h0mFu6QIMJpITV46gQMyaOAuYruoMewS1yY9t0nVYtoHS5c5UTwczR9302EyC0Ll
rfoaS6mnXLvDmkmoMT2RWFrJpgSxU3Ie8M8xjfMLmq4bvICdum3Cuc6oQk01m0oBlE72TtVNyoBU
Ltk21QuqWIRYr7Xrej+p8qTh12Qzg6Y3juL5yB2xacnNzmZE/xvGmmCf9epPZ5vhudlI3Q2D+mM+
6Mm4pVAUT1EW7ZjYsFcJRsTY/d46RZBfOyHRQO9S+eMRsDo7vX+flwzPLC4IP/pv5OXAneAktz/1
bdNYCmJ4tmJ0ptUSgteZyWgMXUlRzoPvsealDQoobSJSMbi44/UDyxTvUXzgUs6LLaIVGBPFDlOf
5X4e7uwgINR+aiHbtiAghsbnZXuWeue2ZcJ9pKyLZXtAe80TAhHoPArZJrWG2Xj4xYM9hDNDH31K
nGksjuf4B/G1lD2RBoiwzqygom1/5oi3RFCMXnjoM2EPfRuwRpKwP/RHqnk7F1oi0tHCP+kqJXip
Ue62V9MeDRq3Y/O3y2kkwl45BwbmGjgyGDimlrDc7/x3idbwryTcv0jboMnPAX4YwDWKaopCPnbn
kJVIliv2hDWDHip4We/3XEZZi/RRQfw+rPDXwcNHPVKJwVAAnTtaPLek6bQ11an/ecdjRGNIntoK
0CF34omF+t6aK+8GYXLE4Qllwk8naMlWuTjJDuBwQHwGSIe8oCZQUt0QjbjA5WUHAZ+r6qC9JwpN
sNLUOFCLkg8Zzt/0uwE1QBI0MlDDE2B94eWFKPZvARjRfC0JKEI7+m7ckwkUQdeVBEQoiDN8HCn4
pVqnO8qVd02DGARO8dWG4TAJcbgAKGY0MTLHNH4H6czAmm1ji8H63vz56IRIZ6V8b/jmtSSk6X0Z
NZfSo2cA0qCY4J97otCQnketwcPbhUGGjEAdMQBaTraIlKb2Ry4KjbZCFEFuPjJ9HsgTRxotBdq8
Beh2zDjsktccxu44KlqHQV1vydXuXgtefiDJN9xVY4sPpowg34JW1pREU1IPxJ/TGRj9CKEYOv2w
RK6EPLFPgjxPluUurUmGA3kji5/wwtLHGLGCz7nlxhgQN+Qn5gDoxXVVeH/DJ2692TUnblyA/fkj
0prsduJckLtVn7ZE804P6dOmbQTucXi6fFk+QebnCoE6llEEOsPy6nIpNJxb3E+OLofh/PiHH4qM
+lTX2lFH2Z8lEG8W2ebBApIv5Ps3d/MGs8Bwqpnb3AotHQP/P5ghcl5nbHJKfVNYpb1d8mLC8iFM
+lcNZAxA3p7c0eLeCWARZ+hhSV0g9vTXTMETzkbxj/svw05V939hTB5Xtuuc/yU3BYCVKpfdSd6l
kC+VyRqi45isnclGiNFG5KafsC2IBVNnjxjlHabEC7Eg4uSP8bAjV5MrqOjO9CDbIkU7p9W3tiPv
ZYPFH7M/1h6UuDHoinokdAImw8Yb56fF2SgJLtKB+jzbVYQmZhMbgSXlEfzQH5zrdETFr1A9r1IT
R16Hn0aWwBt+LJ+P3vCquElpB9Cw+rmUNY5M5WpRmUwT7HMhWdwtRoDgCrliYw0apD87bcpfYkkR
Gs2mgxAfYezA7I/ZNPG2KBu7VKRig5egNDIc6O2vJwpfMn3UO5oh7Xe1xIxlNh4itantsijI5dQt
jLcLudSr4b2aEIi38/Z/GHXnqOs0uzEuajxxd4eZdBj1FWR2lDU/b+wXK4kCjOd6K8eX4VGuTFj/
dVrLDHvhbf48ZRU4JFdcu7MQb7V23TNsurmZTaoftZRZ9VrewZrvBlQTxmjA2GFZaY9QhtBuasgY
HhbScqkL4r0zWD2wEw7squPnZt8tCTj0lUt045lovH7NwjvuuJB1lyMSpcPptlBssKI3QuQJ7BOn
aBzu4Jodz9FF75ZxlVub/i5F8nGGGrj5k1cra2uo8muy9mavRq7RZRVr7Pt3Q37mlMvIhVFangxz
11wz8psAEnUfpW8acvu6ZXgQVjLaD6AH/5O+4ObO/XgvJfcKOl1/9gkNCqq7uFHiMAgzyE1Qm7uC
CNFj9Sjg2nFyURxoQ//sLa7O2uET0DxyX5DcsvK/RGEEPaozWaKOrfcLRyPhp83218wVLJ71IepM
hlK6Ef3B1plvfN5RMypHI5My20WtYE/B78lKGj76hHffJ1gb3eCpPlvHc5H6UvbSosCU4vl1sBQR
y4ggN44hCa2x/ZfgFJqt5yKUBlSmYanoSbCwC5wIqSo5M1mChZQLoB5pyqked7FvYHERuudh1qJu
e0HPs1wBnsTo++/aumunbkxrLXneRoxCRs5UM1zgPcMfpTFNqOvBRrSci46zzeUr5F0i83z0NqgM
YMc5KwE87y+MpOKRuQoet/FdSjdiSADKvkdaQeIpLyTA9uMzbKON5L1ri0jf22E25e/TFjICC5L4
s6wpnUDcrXf7bmqy4weYwEx9lnXmQifw99TJLoVSkl0sIJNGdVwSUe9ib/dpsegaNsd1gk7QXv4N
bYOfZbRI8vpnk8Y0KFIUDnUo4Xm6XVnAxvjpwiBi7jbw9OVyEXKn4k+5O7ZZK5YcPDHA07Q6dCha
qIx0w+IvOjlzsIX7OpiBM8Vh/sb7jJDPgyrVXkAyYMe7YT01fCtS4GBDBdesGgrLTDVcqfVa35rd
226df24QHmZOqcZF7Ju7sICDo5EGQqDengAiZSMwo8kWR5xeUxJPTNdabo1LSIG1F09o7kwwa5QS
kCT5iAT64XVmjTk/aRCYX68Poi8DJW0QJ5FGs2+YyKN0qvV8ICuPBt1K8tssWJoASNm3al3QxXRJ
EpE8Is1UnInH44ffNP1E86T8w9D5eBhvEcm7enJ8uT3K0XjTXOoOP5jKTCPfvuKMf5YeU80V/6Bt
NCdExzuZKSW8q9VnNp4PTr7xK64irpa3476hIcwdAZpiMIa0qpbFxqJ8OAmUwb1sa9fH9f/sPYXp
JXeQyFVbwlBd6ZuTv9SANaBWYxsGUfl08+CyRzMykDtP9hKiOMm0JqsFNARKYoep+EyMJoWwzpla
BKj84AwSPxLSV2ySf0+CM2wiJpwYxvlWg4R9wRRZwCwaNO92g7VJN9Z96SIQMtnxcLfcK9xqxOAx
x2UURWhg7GHvpF9HT4otO1tS4n3rBb42twPTbZrw6eKXSVc1+u1cEcaL8ViVI0R8QzoiyxBABQEC
8JyIreOo4Wb7Sz0bSjHkPORhqG2XVCSmyWZm+k8cK9t+lK5T2cIvS/0mTtW3bEfNaPnpVNkkqdWs
6VUy5+FnUzg1hIfiqWg7w5u9qOsZc3pRvMb7I3wddz60+rRUsOj+Ys8KK8pqXORc3jim4fw34U1t
17Z5jmFleDgRwJBMC3bjaR/J5LOgz/SqrHibXD10i86JZFSWQ2jMMfCgAsljtc2m9AN6+g26ptEL
jOkFy5sp2wV14IC+OMeLJ9uMIyusvDJbMNmhpEZgvBIwbzrvZgb5Jt7BuPqQi86FJGvNU3iz7P6e
rEWCfePGkJZBev0cans31AfzIJu0ttlSHlTXZC7ELrbEH0XebvN7XMVJ6gPXQFn+GRi4uWIt+r/u
j43oz7RRvp07zSZik+s2Ftyaq/ySwAe5IpFgNKpULb6qaiBubPh9SnySsrg9BgyquhckzhAHbKfY
ojzQS7/+sAqUKHlMrqcSwSpISnhdL1dNl4eUEwiHTICoekxy+74mtXPPX+ZZRqbOcE2W2kpH37nC
6mztKJ5Tgc0xnsT1vcfgcEbxM5RAMeUDJlOQL3JPn4vKY9b3awE4s63U1mi1kTkPGGjjTTkn7a4f
kZUraN1YtJpjbdnnWNAN4vIU4/15+Z/IvKf+Xu0R/kkj/MbY5T/HGdJlpmT5GEBe8qYp3Xq2GngX
EJDrKBLK6iX5I3XXq+7KMoMaEMGXjCxSFiXT3AIndZ6cHS6ieOtRcwuAFydSbaS3y4RKWEKX/F6p
E4laSTDssreYNYlO0rjRI8G7HE0vDRVEtnrzVoZecxrmhghQOlkJuHW7GtZAOEZEXuutuvx+yJGu
0p/jMZOqyCdRo3gcu2zV/ZgNzGclLeH4xnnqTYzqhpVzByfK46EmHRopTA0rZQZH/htae7YWdW76
z1IGJtLRn3ShO6TuWX9ys/S7HDGrYVFORPTAka0eH0aENkiYcAf11ys6qzytSdD6VIpk2+Cc2/pF
HVZCy03zYHuTocxgwKmJAwtpo/b+P8A6u94dwbAq0lkU9/U29zoBwZF8O6qFv5KbZgNULI+uJht3
ktUop21jpYaHePZL41IPV6gDyDG7Mz4WngnEoodrpryaScB5JTScaGP6E4WnTLs5LyehS4mnftm1
dT+3etHpZ8VUSaB6cCpLkjC6wL2QlZaWOH2nFl6aM8Pc4KGs1HpoStKjnkyQtmh3HDeyr6LcYKr+
fc1sLVaZz3ujH+uK0ERtssA69k6Kd5nSH8r6OUOBLX7DTC29Ziliz1EiAQHwQ0TK/7nkKHF2pb5+
su3rqGlfdvHezNwVcNlM4IJlOAz4/yDobhdI6ql1vxLH1sKzGMq6X0NXDArC3VxDtyGDdy/e/azx
7NY4eTuprBB0W5gwKIixYTQoCzCZn3TcWr0VuFOCssTd6B9Uq6Eqslu+4NoyBw7z9ltryXJN2RuV
AwzkKLb2S0sJHi6YYT2jGooHZYm5KbPdFqVehabNkgBh8ByhNwsbY4VvdNIXwO+ENElP4mUTSL8D
nqxPX1qARCyXZA/L8KNQUwIknM0iPPLdt9Z4ZqcrjFkg+d7b9XasknquNITJ3ZjLtdKJJCorSnAq
X7UoccsuXwZsaXdgKOpFD28/6aX3HrGfSIH98JOJwpoGHGo6phaii2O7rOvly3SKhzjiOekUN8zO
BTwAf2kpIdnhmoIHWD2gyR1RQHSOQQoRSlP9x1bpSJqWyCLgjDXWBJ30eGrnJua5GeFSHQrA00OC
BszoMD01uUAiutC4nzAZkkXU4RaQUMuvOZoaGSBYba/iGvV1EUQFpf7mK+bcUR9RXj8qkaKDb3Qp
YWxGTCP3HcOaZrehtfmLPJAB0yuJTnJRGpshk1emLUjoywVL2w9UKtmGCTSbfC1a5JQ5PQjMr51J
xs3C++Y4o3vxUJH9XpCZNqQn/SEmt5uslQDQpZWHNbYLS5idD/iDMu0G1+iSvDYWMZBBVua76l1G
GncBU6UfFSgBbu5XFtTEOw6zLqpLbTO8P4+fjEiNM0F52YPyGlMmTGOpJ2yTxjZZ8I/ER8+RxOeH
8x1gAe+fDXrM7T8Rf7rwUB5tpdOyX/rWH6dERhpEjkzBVXifPBQ/99GD5g7kWyIJQY3XFW0em2a0
eBr33HziRwsttwG7P7YwOZBrT0+NqEku8FcLpc7P1f0keFMg/hPM8tSme4XPIXVMBVgDRNv+5KZG
7R2/i1kkyev+LBwDOvCE0SZKIJBIpZ8P6MXln89oZcYBhGex5nY4MC0IeIDM7LqTOnogw5dExgB1
SwBTxtFrYCI1d4hD9uNNMRlSW2+zbxnY6bDabKx1amBJknzdtf/zZtoUBN07VIaloHgktyKWGLpl
L05eN1dVqMVEUI3aTE8tfIdWpMPr1bOuod2YvlfRE2LjLM7lv96Lh/VvVGH25RhDhbI7I87WmYaE
yQ7GSQOTHxaM81z2pzHX6IXzyko3XuYgD4mNBIMFP9ercQjJ1eTa2u/aBKkdX+fS/Dq97VWwsQdn
tI9/Oi2tep0sJBqG60mfexHZSd6gQEvNw4I6GWwN1Kaw4PlTUIKMjVYwPZcfQ0O9u19r5HjZxt4E
XC7wEYs+tMV2PH4fr5241PJmISF+D0/T11nwVMzDLh9I/UFZ8rGYGTx3CqDDKf2sGFqYMqiYbDuy
soF55wft7cysQrICwPUwM/lmcyjF+sgdjNoyCx9OGnb1cFQ1bZABNgQLJGrD4JvG1cT/8kPd/wYN
Za4RoJMHo1Rzvj8vYj6IVa7OEoWf8LC70s4XZFo1WFqDwY2YOqG5pLRjSRnCYWhkoQF0ph1falz/
6um/2r6cc1QUyED4hX4zGLDwayDT7flVFnunbde+T4E/N5G/dmD+6ZK4ZxwH/Xna0USdgJTs/Tcf
SdMssgkGym3eNRCIdtcm8z0P9fSMqewWbbkvXh3wtn9Iv4Wgywbwf4q8/rdUU/COgB30tTaXnJB9
CTDDVuHylR4gdI3SnZsqL7b8l/P19E5TejwcE9XVrkObayImLGHmA0CB235hti9I9TIxhoog2YXx
9z5CjKWaequ/jnHq5HXJbVRjptsUd5pgxL5qIAfh5K4RdBWhDwl7bmkkKiTeXYvt7vDzdPZxcxXp
1Y8JLKnxt0+Wp92w5iffBUNaCscIHfl3kUT6Sy9o4+mVbqHtd8JGfOZITVpG2dxzcgNZS7uAynGZ
UWu77iikX+dliRsIzZ7U38BVTNCsG+SCG1w8Tz37oo1SpgouvQ2njlLz71LYftFglglIZGqqtf36
ekQijjloiRFq+romuna6WA2f8kJ3roU6jKWFSyJhJCA4AZLUuIORqTzDvyTikYqkzRXJxedYYfZb
3aLYjjRPBMrfa7g7T5aG6gJGFKnqzgNAT7trTYuj86a4Nnz6lDEfN+ytyuA5xGEZCM44PFOMZAgk
XRc6jF73OzgcR6WdjQZzZQazecQ2kPCZG7k4fnGwJzgb1EXcHJB6bzVisVx6vijg8K1taGzuQwj4
ck72u/vGHW8nUbla4SoNYGFOqC9Nw+HmUKehqjhAG/UL1zjCy5mViTJkDu8R0kp9Httg4upbh/Dq
DBPOBNhtCSyR7iRdv9j7KMh9QFJAZA1iuaoZz+McntZqnysBcPMjyecLLPCi9cee33sdyMGmuscx
EeFozoy495vMxCBWVdNSR21L5/GXZglo3b5YMV5gHW9Mo2wxYTMn+W2lZpmy0gWZByaVHHWyrj3h
4rwq25GDyCVyPr4G5U6ZRkzsEqGdXb7kFjVedkjq4p98K0AXJUVrRey9Owt82hBtHFYJZIVynUrS
jRkfMGesAj8JHjFC9F6o/FgEv8Xyu/QQWSNP/puYToZkrsN+t6HScU4iOQusM+008Z6CwHEbRX+K
ypsgBYv/SsPW/PVRFMFjqNKSqZKOh53VEZlnm2RS8aoRZFrGr8oXhCsve09qLAIkjcIMS7mjSUjq
COjgQsYDwK2Mn17EI9YdgQmOuLKai9E0TeVHSG9liGAkFk7OZcRjo5+xFHKkvFnyJHwR/doxIvZX
EQsdNWDYIeXI6gz6vz2Sd7nDjAxWX1XheYKSIYsKv+K/hjhcFJEE+rbMZ3qAEsABqjx1JCSE/dy3
+L9wyq1jSISKsl6vx7z678UvKtyAJPOwHF7mlpDWD7LLPkssApcOry9oWpxzDSeEPRSGd3aA3dYt
GExE894BnOPnTSRIsJxsEoBJCLZ6n78Qsn+pX93cwmytSRXlWXbBy7ZnyIe+iR+oALtuxPq7wBVX
9AWPfEQ/GSsc7HFrHdpAY2KT0KdJzU4oNjGWkzWMLE5pR7+0Oh81969E3nK/MehxEgMLvspbdAoA
Zn88Gi2MtA90KFZCNAqjAanu4hG2WDRSON1lrAZjNH+bK/+kMOGO+cmDqtP/C2mKRbbyEvCzYgki
ZWBP2+5DWZ3go9fuRWvmapvtOwCMJLfwJD2HAwfdK4uJglcY6OaV5sW8AWvxpk+d/QbwyAUPGvKf
lzHfdoPErmRDgft+pojnjmrq4q+I4kRVez9ILpG4Owl5OBv+jPz4Bbc3qqBOmLoPJOvBR2kGlTb8
oolDtO6USHaQc1JbTwKTO11Bjd990TSdXAMb9i4myMFe3CxFS90Libm5rFdlMSCy6JloaaUQvtPa
TljRgJ9SgAJ+0KrsKKVA2rJBAAC7opk3nadqJgwsNtSm9MSSkUZtGmTcHuMAag8+80p8M4nFfC7O
WXlKm7+6ritgGYPGZsbbtkAXkmokt3tEDIm2WPihQQD+NAWmRc4aZJEJNq+TpA1PYP8z5Kj64tEq
DQ/8LYXdT0gy7gFaFdet594LuGdDnaWeJv3a2AeKX5iBNfbKKAeXuKoAbd29aTof/LovWmsab9Db
lqZcRwDWu0q09VZheKCA04iotrGIgU/iue6BIbTOo6YyNDonHuWoC6u7WZt7t8R/XHSFrMKSUliF
76rfq4lV3edcY+85lmi9Q+c87+sf+Nm4AgXjnkww/D8xCXGgnVyyHK6XEE73fxNrrwSCAjf5tqzv
yY+zFr6qZiHt5O3EzFQEpynQRu5L4cZimSf4xHg2q85qBHS9TkTEooElMZSNr+pcN47IrsJ4Gm9t
5zPX1o69WDpKNRV1Axz5e/4HkTUiUCBAivNgpdZo5i3DYC7O00p3fWs97/Gg0avKye/DaB38uG72
Nz9Ge5VPFmMNrV3r0dkSfHKE0d6OjEIyNlt70SNuCcOR297njR+8RfCaPnuuS9Zf9qnOD84ndFW2
HPRMSPmaG+ac7SexCJX+/LvvFISDBNHAlpG2ud2LYXIur5JFT8RMA9BJk6muuSq8vzQcOYmxRUgN
HSA/1TGsmy6B+jq6ziz4tQSO3axkSeAcqW/Z+eQd0mGvjofDKC0p9wABVcK/znpvTDi4UA8rEfRH
PMp2SalVXUeRzdOsWJRRxCdraG8qnjyP/IRxVqjnWfINoxXzzsKgpsJnknxopDR+F58rWFzo4KpX
8XxKliv69oK+bEp2gZ1YtlNbf2/9gjpTYyzjdUxpZIrB/wnyPXlbUGU2dnXVuobDi1bqTRqA7nyG
szWs3HYEfTC7mckaFVzERSB2KbzMFUksrX1q5Ev9/2w/tFQAov36EshQpJc8lmOc33j5zlnREGS4
DekpWeFQ1VmZeBPT5rdpkv8gYPJVS2QbZJ5mUwF6yZgVomoZHHvp1qw0EKtZcdUfXmDhNGulmvAm
kakjisYMSHRX8Aqmm045rWbwdsTwOgGKFnNrOcG0IgQRFMftN/tdPquHPgPvGbaat0eRBV5IBjCZ
+lkyuufjdZP0Qgcw11sOtJGuxOjjiqXYGMtPbOQWGOq1OmlH8/cmex98B2gobOCIr5gW5uCWT8GL
hJGewrJ20y6Gmb8Mynq9Kwm5wEku1FmEzEvsAo7tofsJ0WGPtoyNz3qmRaRkgFt+sfUo/cTjJ+jo
ppf+azHGnic1THScWtFs1T/XmISYi/VwuDnhr7jCDyFaA1WcJq014ntcgZYhos/IBJcZPOTOpWIL
RgjezVahha9a8rrjmeA5kkTTS6CeoL3/a+Td5yfw2EJttIqXT2uhzwp9nANlImB93fw/hD3TzleA
FOGSVT2zXitFnsj9i3SO8hboH5oQq/CtE9iWUf9U2dPPXgK2Qnxt5RHPf5Qup8aVKJk7rOsGsHgX
1BA7w8lwd3rW8ouSXm8r+sOeAB5rgQqUAuhfn7E0jwlhk8v6Gh3APN6lLLeL4pFg5RS85I/IFYSP
J2VIoW5GUJiwvtFnQFsRz4Vg0AOHfyDJB9rzw7+9BFl12mHpDw8UA6lWOR5CEOUjvKX1QlUpKGJX
hA98Zkhmj3vI4fgYPTLUBnBDAXP0CfmN1FtIU61ICD8XR+x1z1YYuPyZt8ISbOsXnKOtJtQeTKF8
cyEuSOBRtoekjyh/PzfN90wmd248+D0KZodMxHTbBPB26flceGFsNkmQALf30Cw43Wp/RUh7+6m5
sa8ONlzvKccBxj7y0qTWZ7jiOo0jQ/cd+fLBzExZbZxGBUJzDzxE73ZCc9JNDmc33OUFFY8PTOe1
UEpUA8QC7PkEu8tHY9q97TzLbSZKQVJzJb1Axj5G4yGU6ArNIusVR0qgr73WCevodPSH6+uxocTo
07Wy/HdI62tiHGsQ11TpQHNL3Yn2dPuFyvYtdBcRbblrN2ELfOZ/kj2M6Vnlse2zAN55PRboQFbr
e3MApilwC2lS5VL3x6H10C1Miu4OMYwxNuHoKxAoPq9tA/yH0ZV+Wdbhcm+lS2ONstwbZExpkN1C
4jsn5j70Pun8097cLPyQ0VZAey+ENmqyFpKG0RlqgkGoEdZfWGo286xZK32Apasq6rF96ymEWRKd
RY37QtY8r8ZrE0Y19/oUKUx6pooyMta8D9xs3hO/UuUCsgAZHAV3ikZIP/B5uTqpFFkJ4FHSQWzp
hW/ASbipXmDIYXWOFduQM/6UAM6UjXidA24Y/FbXAXjViN1r0Zl0RYaajEsTFYk65MwHgtW6GSzq
Fq4by8JnYOa5XOUSqeBWulmRvR9Ysig60zlT3Mgd1ZaiJAsaeGmDyLbTbcKEwg9kUXflCFNt48dS
5HEGK/A/hA2bsczEtJK9U2qJVxx5rwftJPol9q2RjZN0TL0pQShSByF/OyuHefk0aPXKqegsQIo3
YkW134QMdnkyqmlDu7KJM4QIBc6Jic6rJDEu5SR8coEpw+AEaG6zYmUghMhcL17mkKuUElJ2hReM
BsujxKNHHIAEIYCSrpUZYo6RpESA4u/jkv9SEAj7La/TcRomUnH3GNEXH0mIqfLNng0uUbZ0Qk1I
747KkLJRzK7VHrnkic4eQwT8ZyH4mNGJiq7CH1iyvgOLOqJjmIDv5HY6jrtVTJOuAz/155iOFWDT
szivvA3XY0WrxdNyEp6v3qEvsXYdIrCQ+qsxDqGLkEBE9xteQIHSU8snQ5pWvg+wRls9UwPEIVbf
voic3HQoWZ6wUy3YnJ74npF5Ol6Yn2otcgajksiCZSuM/0GJlfJjLhjU5rIdifIlnpaycs7uXyl7
4eUqofs+YDhJfyh9SYImYWnsJBrxcDJv2vI6nFMg+DRJDNcQ/TJfl4h22yPfsDgGI5T2YvGAnllN
+PrrD3LY2vTsUeikztuYyfmkyHsZHHcLtmIXC95E9gWGb7JEtVJ4Z+fNq9IVN8EdGnyJG9WQZ+DN
y4OmU4uwPEZk9DZwRMvkjwONrv14TtNb03bgXINjvnKpeu+x03v3l64a9ahZxKrORN3WMuFm+G5w
oE7IQDRR601n2AjsgQnDEUO0gGgEVnw+jwNCeM4KfsMZ/InrpuHvwYW1qdT9g1KyUHs9ijhZzeZa
vL/5yUz4BS311a+HFU6kzDlJjEM5FBVaakd86dBztT6dXJS0pH90L4i1YYnbCVTcZQq2XsG/zrMa
h5xCm1IrxQ1OUI4aRn/yUwisnfC+xHZQYIu7wRChExqj8gp4Pmz+ZeeY8dv6O7pZCkodDgUCMZJs
ojjpfFc9v+k37LzuYfFjJOsYlQQn4xjqpQDbUyMLZedZugioRe2AVUA/dWi0VBah8EK/dnNcw8SP
rbDqzWKUsq008rEVmAq5k5wD2L5dWgnhIIsK8joxeYOmjz7OICeb/IGg2j815XkY80YtO7B6Sza+
Rx0YcR22RVoGo49ScTYw/hyU+yVR8/TijBQzkTERvBFiwaTs915cR1fqwqpXoWCwNE+jBC6+rveM
vpxSIvgohIaPuIaRIEAkNy+tlOXQizFJyyYdbccFdQwyYAeIDZuI+9oL6l/aSYkq7KQT2vw/vffh
7knrP7UHxNMaJDRXM9Og4X0evWB3DOXbyO3mrJDPajXY5GaRFSPZgcuXzS7DFt0/iMimw7DtuPD3
v/YQIryqvmMos2bkvZuGu+cYC/VTLZHUQ1eWJnvTcDC0VDC32pLoeeg7Wl372vr+eoptpSO/SN5I
Xmh7+3pC9JweaHxVYcO3YWPnBl34EVT5WZj9B2MQKQSOWzXizEfofTFxu/tiy1rnCF4haYxPHEqf
KJwKGnI4hpIX1cI6f6+MuSW3kpG6mFpzUfveMIsnodjOjmE8l1S5lonOzrA0dihUPbPOQJwqnj+S
dfZ8GOwC4s12WIbGxbgSPFlCzTD5ZfO/OsVPtAj3uEDT8bxT/lnIUS1wyqKf4/7XzP4i48LqrcuF
I6qGon5UKtuGQUqnn73ma+oH4rwUmb40R/0xKquUtXvMShkyxOqInmJxYhHCBw6OSDQya8hKCgcI
xI1IWgCxp7YeyPTr4iH1l8RlcpxoTeORNknZY5DY1dBeN7Hd/WsJbUxAEdPAmFwMjykhEclARNKb
cTFWjKrA01TF3ZLF3gv9eE0yMBg14FFH6FmlrrP8B86SvrWJQk8rl4Ro3VB6UX+1qd4pvnAQQXE2
/AeS8PxndxooZg+FFomPdTxl4CNcvy/Z6xT6d5MHgXFBPQ1jpjLnBAAcUeJwl011ekCpNuemVJdi
3oKAPODFniVx63WCrUmfJvnkQMH1Hz3CM2w/sNNBw5dtkljSz+jt7GDrmmFpEw+dV1qeP278ZaGp
8654lqE9VWj42NcggQTxjUDwkuAVOOnNMXUYLaRsY+j5qrwVjAOJGJ2jBIOtxIDNcDYAlwZouiFf
5NB3WHh0rl1LMs77Z+F7+C8BOfcCXIaUqC35KAaw5Mkt/YWbV8Le/sCHwqlF6riLjmBv1zbC91r2
RCAdpvPMDeo9JKrTdKr5OZiO7t668lL+Cd6OvGebU4tfc2kijjCj06sN10pGjsLBH/1pe52htYBN
HSI/EipSGOe5VluTUtfxU6H8tr8mEM78715RLSdgTR7uUZgHmqAh7u68Zana3P+YrntEP92Q0/rr
Gs5z2A9ruL8Kz+B0RJq+hzWT9XGRWf5O8qg7LE/3RVHU/Hv5gddiHZxfRBdm38OaBGjOndkt7Old
hTLZgLX0tKaG5eYgMA4kwi6xpSHIPy58Y/6mFpQFH6WoGCFhYxD/iUTVatoJhuX/0sOgM5nJmhWq
K4p66aPFVcdn0BA4QP9WxxkuU1gHt1UwjGJnas184cLydvVX7/g0XHPxil9u3Pk4Q31E6FJ0jXSr
1lszmLmQTnvUFHLfZGJCiOb7er7T7XBF0TmzustxdhqMMvp+l/oPfdTkip1Ixcn+XwzJAsT0J5wo
G98JKGRCet2ua+lzd2BTdpuRPKkc2SWG7OBOcC+UGyEGr4MjQq9bcIkqthhK1sEyljbf8IVX0XlV
IjebZUyqXGmyakTvyw1C61nqCDbLo6cD8DJE7aWCQ0+YEbPqS3faAvZoZEeQgEFrLoFdVVYRdBdz
CJb+Z/II1OPFFXhT2bi+onYlUwXpr4dY9OKZL89/RAXhCziscnoS5eAvCmHZZW+I2N0Q0Jtq5rLG
fEk8maUzcYUztYtGptXEnmCQzIOLgmJFFKNZdtpuIjgvoQGVo7bvVwWwyBeRZd9jgM6Pyrej2tvj
HeiuBUckHSzgl8XMVazUhiN4eAsTG8OpsIAP+x1OqeXU++PslWcGZb4l2eh7xGdppJ/G2lMWKsiV
6ehVol6nnr18wrfiWskQmIixxgLKEuPweabqX3vE8Coh6XTA2b368I1Y+2nQcrHR9EG9qBTwD8EE
t/psN8NSFpYpTVsL4dlzvoYiKzOqOYAKZwixP1cNkUCnFFKBDOl4EdV6eqyT3eTA4jweCMfb9uef
yTP1SiDOzhkxxeR2FUPG11W17r4VwdPqVVWR9qm0G7vbycP1eCKPK2EvNcuUG6bUPPhArkkK7Y0t
2/e1y8lQ6tK/X5v6y12pnMjO+XBBJn0jWC9+AVKbDz/AF0detXspi6mz03GW21isPJgQ9IwNF44/
x3AyMBg9OuRrwsqb4gHQNJkfU9upWOj6D9WJvQPeick/1i/L5trXwLa+4imnwJkozgnuTG27dgP4
TTjyFZamH+ET6ByuoRi5FFMzZJmd7LVdSVu+fIqylUNM7MKblbEnOTJZ0cEjOLei3/R/Og1YeMiB
5E+ZS5gS7hJqOwbMb3TE/5HfIPVbw1YLmPseL+DizrZWd7Ewvy+0Cn0mc1/NgevBbyf38PEzik/X
mEnYqXSyyo6nuZjB2tZMqJuMJ3c1f7HQ9TH3qQ+bPr7ADvwhy1YlnLXIasiwQYyrMcxTlNldOxtI
oROjmwd7Mx39WRuv1elc6VfxIfmgEGxw4pFhx7JH/nthY2jDfdFNYwALkC0lb3Fp/vKAQA4g73+/
sLMuxu6p9GJK9lnz18efqHps/iMFY9ei/hBi1kZo17jwOHHTUrJ89AEtHAcCVdbT3fP9vAdqIxmq
dcQ33rVAU4DlxIuxCrGU3p/soDl61adZCEAD36w2tCwn70b66EP50qZ+0mh23YG4uWH7tqREJujB
fzEf+R2WGM+V6ac6jtZinVYQdsPX5fXA9j1YPfhLsm2eFbwMaBnNobnNZ/HIVIPr9bDRLFd9GWps
FT7R6LpHYtRXPjzROoQgZJbPd40Fw5rGDSVhKKw55tqVZYHC5+UVLlTm1f3BVEBOdrJUhCRPdtGF
Q/N/KWATAeZ962QA54RZJwdZ14H/mGXoooVmeqmS8N2FpMT21Ro1BLdQAe+kUdzR8e8Zl/yq7lKU
Vx2lcK5CZ7c47r566PEFByQ5ExIonNALhg/sW5LzRrBZXET8ADldV9Kf5lix67MbfLI1WLnnUhRd
1JdNncibH5OE/qGsIArh1CfOAh4jnIbAsQK/MIn3XFUobz2fK6bea5SXMLgkbb3hDuIurGJlUuZN
MaTtFfKDzDtRyd1xDUw5fAXherl1WhqkAWMoh9v2OO7GltkBTXTMn+CYq4lLAMOpi7Uxl8XBYNvx
Dyxt0XmKScpX7YyQcUdxxflh+Tr74WwMqi4Z0BbSfnQWyKvyCQlAtiNRQEkqsM6VQ0Aft5OKjzuS
Ijxo3SCL8GuNQhb5ZkeRcaCPGT7Jt2CcwPckOb2nFH2Bsrl48Yw568wiy3C3PbI7zpIgLBB2hInq
VEt1kYZoDnD+/eYRnmwgnAgZ9VyeyJzpXJPkrgK/W5TK/SCZU8fN9KsKHAwlx2/qICcotrR9raLz
R2HxVx1ZqGH0hTgsDyXoLJ25kF0/GFhroP7657jWy4C2wRDEpTLEl+tqoKLNGopkJweqii9jQqNS
etMpmkwyXF59egOwR2A+qfVkwwgctFZxPjOMGHApRzB4FSx2QGAcBsFGle2QhM+HTkhDNWj4EM1s
EBblQZN6YKdAk6sw07NDvEt5xAfFx+KRKnDJE0lSbdzbNzroLMFP7KWv59VnEYhmCR507ns1AAmQ
YFfeLxTCyG78qTFxGpgpVdpySD9QyXySeYQ2ltJp6ukWry/HpUwzndvzzCO6h9K1pFhywx6IUrc7
SsLxRdYHyCALalhSyhsgWNZLRxnlehjYmxAHl1QvvThWZ8RQUdhnUCcSQMspu7TXOa9oZFRBbqpc
K4J3H8Cc7XEm5FBnoA2L4WkBI3/+0Y6vWCGtQo6M99EljQZedBkBHboGVvIL6UUbdtGGMiaymMzh
Rc+NRYc5k1JKpj3lQ+dwOEt0nY6o43TaON0kRf7SDRODqUJw7wNc2CA0VBFXMBdI1FrKHZtEz5pA
dKYMujdetpsnFi/HzWIYjjSMRoNVl/HzWa3iVsqzH1a+EwYRhz06kOHDLfETalUW8VMkXQB2138b
Xo5NKmegaLnyd2rXXlwnR8As7TxTBl/eCxpP0+HceFsJ5TVGEbkcFrKiHQLFLRa4m09Rg+GrxTNH
GokITBHskO5b35lrTJf9iQudiiNVBUYOrjOd7w0bvT9JzlFyTZH3Dq8qZVESAlFWBvGIu8k1xGum
ZA2WXK1auFvOcjv4LF1Lh0J8StJi2dpM1kELiAv1dSmSasYy55hIILExbfNgkI1LrcfiEpCfM/jE
oy7rBHu6KYJxINE/HAYqRgqxaczFJKXqz9DyUK2mItXZ1mTUf/vAxBb97d6RDp059R/Nl72VS9RO
xZUZot+uui+mSrlqMHV6wty+H7vYr3mvEk3r881OLDks7er8EniLm/g1du7uobeXP8wO7ATeEW6K
AqzusKM4XuCNBLOepK+te+B5TjloDzwcoTvRoNfwSiEgNLqBuNJ0c/Avh3pSgnVBKGC7sZRthn0Y
M+IeVhlREUyEYgiIMAmPA6L0G3m2l33ncwzlpmCgPzVye2n4emvCncCmO/udwaaS7h5/3IK9gaxq
M2SUVLk+qsxf+F5xroBzEA3D2pt6MJeyu3WyGR58SKEZ57+6zORTtk0kDmBJvbaYQ+kBdYU92jNK
mwqEzg61vlSIhrEDzVkifTZf0hYvPufxmGEjyHOcCCeGkbdhORFjmBY7m+2YKfFjqPkmPhS1lU+W
Uuew49nzmznVdljiXiW2I4TtI9h+VOPY1mmxic6nJYy1YSjJAK2yP6HQV0wGc8oqJ3YCFyb9SK2v
Va88sfYt9i9LW+SjT6Djhei9+xdxCgKml4+r8WpBq+UrazNqUt5SRM5Bs3/QbZDXmvScmtdVNvSC
Lek7v3frbhX33848mtWEVv0CPOGcO8lGtVFzqvbC+Fdu4YLesO3zHrAw3fyaQXjSUAJMVlPA5ela
3Irgr+5Zw1clUFb+UIPIJ5PKzjV737vE4gipGu7niIe+zxdS7+spHRcVNaiEwWWIztyNqb+Q1Qnj
CG/a5nYkKwU6XLQVeA3gQielAbkSRVuLfa7UKpiKt4MnC1U4APHdmPpCDygyRKUeexY6haNLfWxW
u1aGilAlZsUvfTaQBxmgpdS9xi8UABB1WD6GUFHi7oXnXFbW0X4Jq3hkhigEbf6AQhlC9w9+na7f
K4FwTi2/xo+ka08I4FkTpRfr0EwsFKWq1acl191wMG6nNscOsHMgOJEMQW4EvVXj2H24DFnWUkr6
lonB9Gcc3anYwSQC3Vd5c/txdmF+M+szCZARCY5V6YwD68wVbyK1iCy+83CvMwrMAN88WG6zuVxp
dvjnXa/UC9VXup7QAi5oFFgLY0deXowh9LWe3MEslKXn+jBb4WOBv/LS+ypRnQ7ixbowcpDuu+2+
0MdhlpbCA3mBTSSHFxAP3Nhx/LvzOk0Y2P4VMS1EdTNgSJOK0jd245IZfwGGT+zyr9Ki49FhYJCU
KY4q1i/uXBEhZ+/it4VNqT99M73jlw4SiaLbvRWwtf7cuyDxLrte0TLDITfn1BVVqfK1nJvr8k3x
LvpUX09EmSRhJn9gLDiAG5VoG3wSlj5Kkr59pYkejvw088rgvXK2HelbkqnAZ6SAYKblLs4pDlWJ
sWUSMI59A+srEmTWYJfnFe4Ne0/VO+E9V5HYWJI4JzHf40rqfy9oFga6+AfgXNjW92PrcL0G+TsB
nV+fNGjGyzcj/C4psZnK9Tc/SCYEd7KkyTMC1d7wd0nq4CgdfsYeKzDlf0wIlRCjYRBzbhelfd/y
4vUpM5y6t7x8nhWCSTFhr+2tHmPvOnnWyYKhSR/cO1CDbBkvPthZ8/ePzWduvFMmFHeXJ6rwG5CH
eD40FQlwpNfl+wdFj0KmApHUbuYuVHmpf/hCLrz4HRv0NeWHLXTfxEPqFqogsIJsDrKGC/EDfLFF
O5tr8Tm1GiYHtnU+DyYOoz0yozbl1ofPC6Qt2BCsSESjp+ilvzVzSUnaghvmxqAtZxpErHbmWWXa
100gYnR39e56Rhy9zML7/iKOmip2AydgDEuPKJi4vlUQ5s4eqLD/xxKJWp4/pE9lwPHQY76YKIQx
dShedKLcQlwWuUlXMVafvavHFb7tJoRJZ0sR5H4QABum/EYlf6kFuxhSY7cko83HaxRbfDBTDJwR
byDajJ3Uq4bLFSHSf3+Gh9Y00rTXiEFc434F682jxEEmUmAkkEYFj4tkmnQELrXJRTGxjA129d2a
B39DRut2UTqIzJ7KN+g3B6lBQgzIvfGP1pLmqTJJMPhNQeiaWKYZZ/uVOZcdN1cFB8ZdX+0wYeq3
iCqzKvz/GXVVYzBs3XoU0kb8aWlUm3hRlmq9CXDi6DAX8YY4LrkE+McxaTzg2SrAMdI+Toeg5z7g
PAtJZm7N04mv1LJbeF5pWxPlw+lyZdSWdTEpSd9zGVqtbImjfwaKulwpWwezDEI3t1gG5f+JCvkU
wrjDkGEvnbk/oEkLcj/0AHvbilDlFrvbfY8cdpx4XbPr3A12UqaoD7rnoax8EyNSlVfSHsEsFcns
Gplp6ww+8X3nDd/ixcJsa33phjzjQVY0JJIpORev/3BuVscD8Qh2/fsZsNDljP3e3RR83s2CLQyR
cTecUOFsq7DqsH1G9mPht8BWpnsOPs0cJt2lVtfglHPFfTZlXsYZ6FqQEJ3Df7+4eLUxSddUsUoo
AfRLLDezm541gJhigMtBzZ0ROziQYRng+Bn00B5c74F5awbdE+IqUl4UKgxO1rd6EFS0z7XJpb4s
jpA4PuGiCIQ23WMQ0lOmlowwsA9wbOHnFjafdznUF/QgyLMOmvgbd3Sf7vKqfmv7iIUwDpU1gpEM
8UVFDE6qFm9JMcC062LnFNgd5k5htLE8L3Detl8+bG773+tLVvMgu8+kibbRNQoBP8HZI3cxNH08
ej39Vu1nwJAHhtTDBTTQrV4PVakPKvxu2reLukeo1smqSM/MEpJ3E87ioi0vN24p32qjNUJe6z/D
1Mu8fa0KUHe+aCrNzLKmA5UZJs3EswMXPDgWtOBXuHwOZNqo24PWgOu1QZ7gHs6M6DfHEpW55P5W
KisL19LasxLUWkhst5b0yoaI64DcPWXA4P/mqmyEIWvt7maU7Evn+b9gi6v1mSo2RD6s3hDhu7yd
CW+rztAtbURTO0J0x9+EujmJmJ9iryepbeJHh/BZzg+xOcf6iVcIjV0ZRMzlBDN3/Utai8J8gHyR
wC00Ej/VI5FZzuauX1NHOFVyNxQd57AYN8djXHVDEx4fTbjw3oBywtjL2XjKLUhbwf2Q7PBCCo0w
LT7RV7VCi0YHAZnt/NYpB7DXJZ8fwBPAkcM772KnD3fOSchTWWwLYkninzXsRwQIqWDVXeLo2vNO
YYuDUY3IFUYG4owy2zbWjkq+Pgy5z4PIw1QKi6qA4+pMHN2QVF1ZDgDMBaEcBebKaa5dhgRjz1gU
zFxMfwBbjOxsAbEIKoLQI2Zvvcb5uWc+sD/xq+w3RF5JP7M72CJQx1fMlG0QGR3v6NUIWaCmeUS+
rPJll5AlETfaA3YAolVVVCTI2xRqCuBP7XMYhEg7J0KDr3H2+09sip6TQu7YWCYkoPcCzOPj9SxO
mqXRgmfX/j9wR9LG0+YQzXraqjVbiE/doLj1uAtyJ7kSVvWIjN4Ai81XpG5piDw4eIybk9oI+XWn
h4flT2MefTS8103KtBQBg3KpTzj8xymT1r+v0vpysN2niDqJ6BBOMPO0BUfJ+XXjmbR9C6t0T3E8
QN0Qvf3pN2p67TbwFaWxRNc6Z2zZIWGqxEkw+Oboev646/fPi7pPjacEuf4P5jP1gdqld3MMTdPl
NYs2/RJs9v06nQgjiZbpa28NHQDIsTeaTo/YaUmhnb4lmcDerv879Ql13Fp8Ma6F7zKIRPzW7hih
vWvaIuwzliIerDG8o6E1YJWnBIKa87e2qSCFgCHEENyakP2pAlX2uQPtMqsnvm7c5sRvMMDUGvDE
cNqBqFMbL1kkX3z5tP7JQ35Ijs+j9d5ct2PIkc5Ya0vrbzeuketH6xa5kMZUABc3+YVeW/vecDFW
8kRPCKbRFKJI00cNAkqfPclrC0MYnSJI81nl4XWeDtddq863rh4lZiOanoM28TnJbdM8NwMb+mlB
PZpkdGXwKrPPNT3M/HIp/9clF1/jBagA6JqBEsAJkRMMMiGx+TgROa6F63FfgK6OjJiReFC85J6+
s5b5bKU+Dz6voR2s3KqY+yIVEqnrNu/BG/NZo2iq1Yp3Va9oMt0krXtAE5HxFont8MRua0qJgjUW
xtkVDDxqT19WZfqqaN4E/szpj4RjL5uy1Sb81mJewmiwuuxXUgwqhH18dstRYnT0rse7ppLXnC9v
Bz2brJ2xSDTFoQ9QloS4E9rxSzymF0QEHq8A2gJtsJW/XL0o3+qrtPZnD+og7J5Phb+KfY20a92y
kA8OWHEH0+t3/qYnOZhMy2pHScPrsVJr5fIzNFIIDVAX6hVwc5lI06dyT6l/eVFKIxsUp4MaXTYn
76W4qPTZoXRZeHEW0f0WGnUVA2dlCTVn+i2+oiOgeL4gOU5KDAXCIy5PiS9Bis2MFrsRigzE9TBR
cPGpFMFSEdFxAJhNrtlq8dUVbdBzM3zoteAstHTzSTRruxAbMWjLXQLEBhilyAIUcTmBUS4OE+Fd
pSW2jtZFEr1twZUUft9C/o7T4SyyH/m6JtXdC6tHkvsnD0P8dJjgMizzpDaTdP22RxAf98mB9ixn
pZcdGaJSlH8wibD1MwKBwiAgxUCdR2L/XiczSjMEOqLQ1Tx2URMIhYr3Bd+vSAVuVRF6N/FD/G5h
clwU3Y6S8nOKAhGf1zX0Xkt5bFcR2QeaXwnqnWeUHm0t4aH2EUuc3r3VoJElul0JpmOyzQ/Aao4t
D11p5HjqEdIaAWQ4qtcRsAdaTHKWutk5qg0l7420vPR7OmS0pYnrHNtmFBDpgpZ4yumX07WisLwR
ha9cPiSn21pO9WtTuew2v/ZOtUhnIRgupNM8vCi7D6Lu6+dB8/qYKKzxBTguLoLmB+D7X3MQWpqn
0gYcFxyw0fqbum0cOMqtIDbU9OWTrJO3v2Pu5tzhqtsAsPSseI7vcfjz0qfvIWUgn28k05DPxj+P
PWtNFHXOOcJHlaWS+QKeSFsnuJ6FdBK0yUzZ5Rpkjr06yMy58l3RX2Wo5Uj+WsgnEYowQvC59+VS
2A2eUbQofBpdcC0/XpI7QHLU1tXbmCMlT8Kp0OOQ70xkWVtX3AHk3DdF0Uu+1e1lsg25saiLOOMT
bKSQpPWNZ9UDx5hwRCO4w4BcgwvmPKu8vvpa49LgTGHjv4zQoNYQx76HQ5Tt4vHZt8lRXI5l4vVn
qM3F2jbp1YmQdYtlol4+voZyc1i3UmDz2fOMGA7GEwJusX9bBvIsKL9JWF0UK3qTAhLo4gaGexl7
fiG4tykKVP2ed8QR73Aaf0MenU1bwaX+usbk9FZj2F4x2R5yBENoSnIL0CKdpoUtjTJ1jDp3EKbC
utz4W8Pob8IIjh3xvLlxGpeaVsEEjFMOQAFG7mcKGU8Y0udWFyYaCP7O6fSl/WeGuREhkiut9qCi
1rry1VAn0fgdjNjcB9LI6NuDALywB+ZKMi6vaiALxElUyNhI/YEwhM6jWb7HEiPo5ndRQDb+G5jD
/pKLsEfRVERh7wk4om6G2darM7sEvkaRdEZeYvRuD0fsOPzXXn3C9OGaatY85M6IsbW/eF5aoL4t
GoP078PhJeW+cgBj52WissXQZ/CQCcVUZxAIrjGvY/IPjhHFRb+dF5XVVZl2EZFNI2+MhXtbFd1c
xSsCi0g1P+VGjpWv5w4LrLJfjHWhspJS3J0FqzjOk8HLqjVefzbZ4qqvaUPXq1CP3UWX3E/ajkVz
VR393JYfk+NRfmQ9ko2E87YzFvy4Nu850ylChMRwwb+sh251BRGnnSR0e+eUGSA8uS+b3XESUNs0
RpYFvqv3gN7U6aqqUE++XSaXHSJlOozApD8MdSC77oIv13u7LD+fmGGDFbzRd8C/WWRE+LY26LiO
lwsRgOACLVCzy63TPN1fz3MgHnG7i+rQ95eu/tGfJrXeXXhNS3NQQnePdSF1OE2gqi5bD9VpkVPx
SQRtDHrfVjHUr4JUHZ1m0rN7sgnGQ6c31Ma53+G/YcWY29lj3LtR7bYeEmkJ0KX7fAowSxeUsdEe
zP4z4GKshxvWyUmd/c8spiR/0pGc+gEwxeBAM0fUHq9ZNmOffb6UXzxplQLoPMuUGHYy7tvXLBQR
mgol/s5nu+OhbPrS1Pe6pNVackEwv/v2fiYhlkxy8hx8hm8Ca+tnR/bdAXM+meyg4qW4CTB4A7fE
OHbTRIS41sluT4VwHUbn3V48SoTYrgfZwmJD5xHM7aB5QT4dxcg0SCcXuLFOrH7hWxeic/UPZ19p
sHtmUA+PqltY0lEeoOHFS2yqd3uD8OakfOkFksrUQwXiWSnhk+piHHfamveUCWyUqE7woACj1S17
EHi7gx4OpX1ek5j0GrRISi/3l6hpzXrhXDtJCxMnyTdGmNHSqff/r19S0VUgNTRZJqMg5FDIFtoU
DdI/s/VsMj92KlmT55C13urLfUf1f4ksSTQeag1GnLRwhzQ7o1LhacqJXeQ/Cq2jh6VTGnmnIF+M
vqXX+ZnIguQd6ID1fJL8orCPqq42lhdlosJ08EQh3vb63+dPmN4wXi1Z5aikv1mn5S//7SGkOZqv
ZPPW0x9zHIZPY3zXis/pIO41KSAuJfkjJK/SdUfz+K6jtSc54Qutvi2x0V/u+yx9it1mMfr//ktv
IhaRDuhH+uslXMZYUxjTuv4VpCbv994s/fRh++KTDnw4EOqy5ysWPDHHnEPeWk+lpt1JT7/X4rX/
3Ie8/kRvLoSOE6r2kcJhjVq3V0nzkTN74Xie5zMkea5gpai6tLmD40KWe9WmiwUSUht7lGpaiO5e
09EJJtQKQ9nKtR0YCrytiiEk6ta4ceLQ6jWb8Um1dm9s61uuaR/gKwwAPo41wxMqporzEfYSJtIa
JOtczGrkMPiB0NEIxFIACPa29C3Ric52s7Qp4i9jFbZo4QyqrBYM9J4NUOZzcqW4deja/FwDXYNr
X0HacYaa5cNmoUowrVZFt7Urzw16I77OeayfV0BNdFvjho/aihv/sa3DfAtwouuBG/R2OQhSVRLQ
pJfj/YP734XD2ABDfgDPdJeLqysaLfx72Fyck7roH3cxTQQh5UaF/1rX6aCOMa3g7Fsejn6tQvit
G623XniUzGx26S/HsG3Cdb0HGun9Qo1Zv2gSwTuj4JZxuVuNeuOBLt4a0StM4o/J6qI1Rb36pMlj
rHf9v5B7WSI9YKC+28+AnbcMTXxnoP3mO8vHLHisgIf7x6+Oj9fbhUY4owGt622k3I0w89XuCSTK
BeH8CLcMCdbykugrCzT7HbWmA7hmHP3aV2SVw902WdYwRbrHu6BJtcLX4AkkOKCBFDgrkBVgYBYN
0QbHSCMbNVZ5B+v7y74FN6gU1LvePZ2uwYF9AtIov6L4lyympvkMxQ/dbsOE8NK3MsaVfREYYI+j
S0s4cIP9fvbhdRUSPLXKI6QxTsCo1TWHhNQzHHXTREvzYJmmIgPBdstZWyw/NS8Gnpyy+Z8BP3lU
35Ol4s58BGEhgIlvwQJ6rCKwVQZ48meQ0kTC9WA9GEXrPZzx853RIJZynpmRUiPv61LDj9fdeKjT
vCE2A2fAktDsQ0AVmjrusVY/8w6V0f74+NXAStSm+DdzJRvpbdDRuextxhkkjocH2yJjPW55bxqu
Dyu9Wog9jyIHjBvWXqmqgwuZitS/RMeEmzC8zCnOR1HoEZAI4C7uXrz9cZEx/VeNEyp3H4URRdxH
UmNDttj3eCDAPn4N2HVNclY9XCfjFb8y663RoTaPA8WNU9By0PxwkKdPhAVmd2+TjCBKJIdcu4xW
5VowxUTwk6G8yn5DHijjCvCNdQLFDPPYRHdOzD5TzIDBU4t0mnjJk6exmyu1VvndR/xALfcS+gJ5
84XnWnHcXYNudImwf6Lwxv63Z2ikC8tIkW7K5atuGfvo9ntBMaARhPgcMgQMi96iYpC0DYonIm3r
NzxsgZgZY84vBgiZWI7LKT2MMZLzf+hIPzhbyXZ+IhfGl89GhifYJcO3Imrf0q4+VhGylKyAhBb6
TCvxvFwKhGE3EL9UqaBkiQFSx/Max06WJcP5g7NYUWhBwZtJMNdzmUqi5I/DlmM4thoEF3Jr+AVe
mRz6oDOQOWC/P9wQETvfsyqzNPDVlR0LFnSXq+pwTxs+u8038rQzH1bi06U7z1kt1H7RQLloO1X0
imS8U7od/RWJ3uzeHJFh388CUZpl2GCpQHWGg6ccvlZyyG4v561nY4BX5xCN0WGJxqc3zDRKCiR4
RoPfauFz/fpGkcQwlt2Aq7ZnMMia1gUWI+zKsWpSBv8D7cILSzfR6tjJ7Ay9kXqsmblRQhcvhV21
GyQaWgvRyC0miAzOZaQS96h9VFjTW1wqETNHi+VM7OkvPsSytsDhHdtLEvQfZ0MAOZOnJQDd4a/v
UyvuXQ83P33r0La8DP022/tkLKqUlyRLO0xz+Zkkn/aKA3RqySRg0iGCTzxWfrVZFJsAjORQncQJ
ffX8zTCjzwUYFSEhD5vLOen3VIyXU83lQzsQITdhH82E1flXW0lj6Xa9vQIgfheQVzHe7WOVFWIe
1RDZmHS0G2pyEijN5nYQaaIofojjNlqAdySJ5D8pXaOCxBTfBByvD7pMPvRgbUZ8oPGpR031LPyx
VaIkhhxD8jMWk7zQetSnVx8V6lm8aEQbL4eHV7PCcS9GeCg25kOql7+Y1bY+5ymcoUIjhSrJbjh4
58fDxoXjri5qMtSsT8YzYF8OSWiRti1TvnT5R8rjBO0pTCX3LDUoADZGdoQ2HJP+H4Poc+aZ2vjJ
WqgLSwhsaZNVe2CrrIZZyE/T/2XgcWNeKqlM/hFLjZv3REn8ytN5qDBrBM8RslMoJa2WApjQA5If
WUfIAJ6UXMlWqxwgTnruhIgf5aq4mOHSaHgfmMrlHAKv2YQW0DSv6ivP+MNVh69e4iaVukQgyZxZ
Rf1qOiDHTIPLnY6lg8bZVaBYyAZ6CEFqqMMH9718feoLZ2KVZpNWjwQuC4BrUD9a6AeYrgXeIbB5
nk3c7nVbmWyFWakkuvAWBlxps8lW4GbbW3b+m4jM4b0reIv2WGj8/YeD/ElHkOyF9VZZYEVlY+eG
J7KEB/70fXrHi69vj2KZtgMOtT8PpKu5vQRkh/LqEuG6CO8V9O5lGPM2iZuX7QA+QCcDmRuPdYbi
MdPXhhmx4bkUYW08YXyCs3Saiq0p/4A1GpMHeucSt4zLMv+0ITjhmiOhQZzdI6jUGsOzCVc+KyMn
Z9vC6/Cc4DprpLt/jqh7CsKkxTabzO31oJ5KEV6l+KgYVD+ebb07PqeLex+RSJEiUqqvMIXody9R
QdDzQ385mhmyXEGfba12HpN6rhhY4zkSPWa6TegvR55tqITOFxa4YtVg+1sdPNJwOYvt1PvM2DbI
GhV9gJG7THYkGEzgUqktUU5JWe/jFvvtUAznGqDgr+0zRC9VwMFEVl7PH5kb0gsB0PQuV2EYo3gU
x5z9wI6sF8Q9Tjf8P/hNq6s+l7+9wgdIFrpSSMR/BQsCKlA0BpD+ZeC9Ub53ZxeMfediTJuG3ho3
Pg0uSAcZGOlrAZKL0N3NLIOaFJMCjYRvQi6YGvauAqyrdm1PJltMBeoAIKFxTYee16itNXDRDE9P
NwVEHE2YfvoK0R5wiAt9WQeeVkI7yiqOEGHfNS5ZumjXkgUQ0y4YBiqKU1ikyT3UGAKqO8DchP+0
St64NhJeJUIAPy5/lcSbOVAFCaA/hLHrh92mAXU4o0xvPUqGnNo0Ey30tZFsFrtUixLW2psD13UW
BgpG0gZa18ih/1GS1e6drBlngybQyijPpoUhUH+xBvzNA9C5no3sg+PyJofohZtorlkdGSdh+MBu
Dcrz+ncNFsR1Mmtvlm292VMbzCkDno698dhCsAqHUnSuUiM152SzGxVdd7TVvyUykYYBmiH0ZS5U
yBpAiu3d8fw+8OKmmbH+Wk5gfm5CJGHtbBuKt8UylMhjQhoCPPK5OrCnUx2NNZStGDr2aGR2wI1y
T+ZjpThlTOsksYbxHGc88bsuqtUuDiaHQZZ5Npol94cwt7nih806I7PT72L92I/g6CxoouGwp5yW
SwKBZROOW5Q8GqoO+QgQEbbupsA0bJfIDxS+fgpRkPdYyrkAKG0U+YwNzriGWNOADUDvsk++IGNx
wPgmYdPEsdC5NjId2XPRSCG7kwwS+2Zudtp+XLo5sZnO8+RZLpRlHudedm/7AUIYk/aicgBbhLxM
F84ZBKnx0ruhIE518MH1yMeZRjML7rASqoxUJwgcWJrlHz08LhGgMMQmpZYiGF7dPkD2CCd0O/r2
T29Es/pmIBLxDRjyBdWvqa8zJ8TW0MabWoTJgjsB2xyln4eLJy2oyuOuT2MZdl88KKn3XfY61MB+
oaLY/2yKM1Tat1+YbUGZ0XSCGxsjW0NL/cnCOT7uDppKlyOg0bgoUUhH2Oc879bPdzkwrzCSfbH/
mEM08EJFRY/+sFil185+keHJcVrvRKrjVN7AhvHkP9OKSOoQtI2iYZZ0K7o48g+ONpac4eVf0LUh
weIhj8IipHKC0MLF3RDV9z2rNxXS0QTbsNKNmH0jQScKVxq4AnwIkBYVs5bmqeRGPpaXVFnHgE7+
Tn1gZNssbLj85czcDmD/Hi8cQh2mDnW/eV5lEud+sVZDPy3u5miGvlVIzUgiOBdIoZoF29pMgaSG
n8S6yBjSZ9LqUbwQ88z1rWmQplOOHqK3D8UHNWFVhge4qiQ1kDT3SvhHMbGJyeuNZTS+GgnGfCf5
U3YKeW7UIKB599tIZZR+wYBKOQc3s9K95JotLDhu7NZe54Hc0NdqtJKQTVtujM7v6Xc/FmBd6Gqe
8u3hnl/ApF+ZE2rjz9lNQ4c4DjibSxDHnD4sQCkOkyuVBZA427xidgiDszgSJSR062jwsQDjK8Xn
4exIYC9zrW6TbmNPnMTBR3Wl+dWWRP46LRWDVDgtuHg0ZO8iLmKyKUxtSs+32xTE+01NckW+dpJY
sXJpxGWomG379au/T90iF9JFrdWKDw9h4RSbtScSlWQF7lUBsAyxn/1Vca+ZCHuHpTt5Yhb4odqw
gdOHNDIwXHUz4V7BYk5IImqPdNaqqVva2v1q0tV3r7lUfJiLztFf9A2rWHocVeIGpxP/4kb1TanX
rNs+3p4JxfnXTvlOVtrbLmfwH0HHXf1cinpwlKO3Uf+2uvldyP6Pul/IiY7opS0XebYaVF9JeW9Y
sGd0OAX5Zxu+s/g0epnEIUYIPvN4c9AUiNWg184mWtmamxgDyQF27/+EDzHtOqhTn7knwIrOZM59
f6ZXjwY7XxOVckR+7V7YJ0pnmQmGM3VM3muWuaRmcj1IKeO0Zb9u92zXDlnHlVxQGmvMjE4S4vN1
vPE7Wy85Xnt7Ip7pBQTXzW+vffJabXML1y/igZ1OTlI1BjzVQTJPWo7TbN5Ttl5WoRIl9j29P2CQ
t5I2g/22VWxnWiNLJanMTHttAvpDehLAZDmSGbATl56CcSlqj63PIzUc0nCnu2PJq2wyOSXHRgAI
2gmvUXVKN5MVNrlVO7vgaLnlUb8MFsKzjNODtTyrxQlhJWHaExFmJ4JeKFQzvjrIeIMtxUM0Ol9L
tuhdU/5gWnPcnq9Dylup8/EgulDxxRkY4FuyRhBhcsqsHJ1tDKpUUFEkZfsUN3U4qM6p/gyp35Y7
gMDMM4G8PH9k0E+Gu7yKOrGstzdf43vBzZMbgR9XKkvv6BWef1R3q9wbV8IrZh7qQ5FLOgIbZwZd
YcUECWotiN515xWFFn9iMGG0rJuN4wmvw3cLKflm7YeLIDDs3P6TBfaL76tAXDWqV/z6EHQlttam
jg91PBfF/WyWWCeKxX+kr7Y/OAODgoAqDQZD/RdJouyN0QQXCcwzmuIppWyfcyLJZYTE0nLhLe5J
PRq52s4c/6ISHfEm+Hsdi9U9k6zSNKMtcnIYTxIqB9wqDRO5SntLF2lB+FdkGZo2CJJJVGRujLF6
gussQY7rrr+/cGBYbUBHL85sbgCDdtHIelRpVvqfTF4BkY2lnYqeArdTwNKRdrRV2Iy63znvhs7n
3tfzR7aPslF4SeKmfF2gp5kNpgVZ7hpmd1IxEISeutlzYxyH62z1jwOXqlZq/f+qZa1PMoYSD/SQ
qqOcvQODVRLv4GnktnQyvkM5hXlmeofo06RXkILobm82wZ8/4MQpfzUV8NULQKECm04/cLh2UHoE
Z/Yp4KsYdW50W2jVtstnDIsz734pMazXhANE0rRUqkQAdCxyFjbPJozLp0hP3N6kyYVbt1boAmsZ
QaaZcJYLzSqa7LUp4yJTxaIFLlV8tRmYrjuhJpdPAhxLcHmL7jSWxHIx85suOP7bpTpaiaRdxMrK
05Cf3IXikDfNB0/Xz0nUCkRut3AKETnsPOvDBE5ILvIzuD0F9+P04z6KvL6aNBEK+CgrlQZtmGVm
BHhEk4/2FsL6Ur2Sgou+kiWxNb2UvnvzBk9cvjtt1qDb1x3CN4KYW3pCQHosxrP6/VNQYdK1a15f
0pNlg+CK8iRL7482osPt6N97BIIrVLtaNIBcbbDFG1cWThHeMeIJO5ym03E4ygOfKFEzLACoEUR/
7ex3pWWp7Oe7KS+A7ar1I4yn5anhNeHHinFhvdWQ6tlps4Q9wYdTlioUwgtM3J9t0cKMwGyc12oP
zhdS1hCJWf3j+/8++NBf2qFQIMQC4+VhYeik2kYiCnG9cgWnJx97plvr+kQykURVPnxENaAJCg1a
OUvBAhTJU1rhYpjBrDn4TT3o+IuP3p0iwoz6cZmr4wtjIp2gHuxPnOmNOus0wGF/qC6CA+aDDSEP
ye6hs7DHayK1Rf+9GJ3z3K+bIocQpdGVaHxVwv/rrMu4n32q3U8f1Iq8YsxaziCrGHWijO/Yqfk5
Mbgdf5TPP7DzmhMj2vgqW0mHHVyoMdwB+/RyQ8y0iAw/A+FX8BQP8xCpm5zfX3RcMnx1AqGWboYb
TBjjWJMCeb5wfST3bOK+iY7pVLJpODD6G2HDKOxwPOxtOlDr63mw6wfOBbH6ctQt1i4XMYgwMar9
MLNghl38Q4xutD7Fauktgm9c9tRCkXpW0SoajKvkzTcRqMJFgwym1a5MYwayiCLVFi5sljRrdmER
9hIg+CCPJIXo6fpyo1ndGh3UZF2x4oCm4MbSOTS12itvZnN7j/DmGQgseYodZClvgaWmfYlI0tPu
0k1KhSgrhGUhmqL6ONPtzwv9LreCkRC7yx9fBfqEj7CX5hBCfqt+vxTQCExmiqU7xKRtlA6m25Th
vEEGDuYklb7B12W6AgZ/gAi91WnentTKV2jeH68pGSxCQtlMW4C62hvcXSefLvvXgM6779vTBr32
xW/mnwf3bd/qzl64u1Q191JCNdBn+zb8ujSBhpbb5Nds47zzPkx6SA3Wwt3VLUsURAoi+tD2RpYA
0wrYnZ/alyiwOETqh/R7dXxX9CBlitUkSpJKwYD+Rj/SOSGc4I0p6eO9cj4ob7BAKp0FT1ndFaAB
5WyBLA/NnuBoKV3VG4JUubvmyHL782yTQ3s07ChJIFe61BBkqErBOreefiKL9kbeQSq7DyYJsNfQ
3YUcNhrSscABDyOlL+eiNhpY0TqPS1gVkvCTeMtB2C6cxoXyhWlenrPCLXQ9aHtB7Zj+WuvIyWhv
ZSTcBuph05JN2P7XIzwbTYYvdXa87fZh8z5VHRkOagqny/Lq+PCpgL4xUUWwVA0yYFR9J0AUTUxG
I5ssXg52ozXe1ueB7y8wT25dDdvJ/DkGsjtm13rvGO9MdurCdsyK3agfK/l+KnORsZ3GPF+Ku9OQ
tEyeoKdHYl4j8APQsNUbLL00h3RjnTJkk9d42Tc7bJ9zCJCKpdeJB6sQnvnDrBmupRjTtp7JPusM
HFRrbVRbze+lkNK8upqzFcX46CUgqz7suGAoNurYfLa5upIwKcaRA+FRfc6ujzLaJKw5TmtfbT7n
/U2sFQkX51UPFClZtxLKJ9Slpu0mnkX8+gwvjqpDjofMt/mnTb98HMOO7u/E8Q+5BPXfh1+jKrxH
GnMHOjGr7jqpFv4CF5eDduJWHIvzI0+gDgZgfPBEtIwvhpkUArwyjiA6E21DIU7Jsm7mIMD1dUuE
vdGOcdq6uX81Kgt+Lk3IzZRvGIz/BmDstwtC0HA0gvB4TW4SgQGVUlKk1dlMXj5VOaK2/Ksbx4nQ
6lEenHoyhOH1cHJA5v3XIQX1RRDsfrveqyctcd3zzSfzT5hYC/majov/NNyy0jf91pohqIc8PBQA
MtsFwoPOpRYXqytAxQaBsHMxtLNXMezZi97bc761a9Q00zE7+Z/kEZ4WuH81DgMI9pgEGT7QpY5R
jySsQTpBJHzldCLSUe+TJH2McCvIyhbuRwWwcGeMY937ph5zsFFLG1JeSAqRfiSdlLbDEeBcVXcp
bqLVgCyZaj9zYx8YSxOGC9gvdkLxkv3qf1i9ltJf5CzuAOoM7fZx+Jhun6jchdfot6u+I4nSd8dp
TGu9Ovhr78kxPoL/8u7ggv5gg1gvc811FwnrusFl/0D+qSrXsCeFXGk3LnxF8wkmMPUIghdFvNsW
F7B9oQW5WlBFLog+QV0r7fUxciDjNcczTvWUJJqPRvs0nnbHq5GSt9u3BoCMJW/4qDOmwNE2a5nT
gV2ktJbRiMf/uNWgyjB0ZDCtMsUwHcWFVLsKXJCPTA/YB8BhrYVehH/LxbGMdOT2VZ5Hp9CT+ga5
uGhQTvmNCnKGiBlc8kit9pvQBPCY8IkJ5OFVo0C/hm1J5I+Jv7HLWm8ukVrIBuxohjiv3Eb20HQ4
KLTi/5tpVF6sRaY8+qnXNYPdMaP0MYRH3KRhDEkjrH0olQoI6g4pBF+TF45g6u9PoDXKF3ZN5ygz
4xZOa6x40HfEMo6F1mBfvks2WnoZEgqOEg7a7UpIuhLGJ0lru2DroZgdveLJD+KRrUc1lT15EW5j
KBvvc3HsGzulscRlKOGGZu15vDIFnfdDAghwIf3NxH9/nPgfP0X+CvpPUNeaf3IJaGgkKLhznnMX
NJZfHdvV+g6m7UCmwQlihwSwwSL2JWzo4K/MxlWEkbPtWOFBPxUPsCqGMxJcu0ONziOiH48B/g7p
bFGBlY95WWQuvuFhHvdQ6WijvEu+EJ37oOz/pQBSnhVvpZAMcdcRrngmT2xsbr6NdUIlBGTe/m/8
zPawog9EFXDalYCG+lMPlslSjA9UD0kSrRQTjOTft3/9EV/svbUhhG7XOqiTWSzg/aToJyW6ZEcw
A1YwdiNqoo7PSzqr19ldSsxlzq2yBNc5mI2jl36T01APNXK/5aEuChNTXObhV5qZ6IGUkAB1IBu/
raVxQ8TbHu2qmxnCNR1ZDO6kflU9To468iIHoVE6pZNklE725LJ9M2kOts3BD7er49Aat45dSaa+
krHfohx7+o7NNjDCFQY3B6NPWNntH7H6P9gJDEq/+JJ9dxyQiwoKJ9ildSOJnhdic050i1mIZlTq
vGp6EjM2meyo1Cr416ir0EQkqYUfto3vwdHjjI/0ABgGjOI/uhE5tFjDlvcX2kfMzyMvYP0J0I7q
3KlztcjdAKTD9zPCgZxcbaGFQIf32JMw2ZWcIDNPcwJeqEFjBN+P9rKRL/d+w81LPUHSgS8xsgqW
fMJq3JGxC5KP5tR+VXeHj26hGggDPNe+xM7CWDAEkrc3MgrZnjXM9AWhptsEXbpMbmX3slUPR6bZ
5EcOlgVLdQnzBztumM03jCELCRGqWmnE19ELY+rP4pfG1D+oTzgy2f+6Wn+2UR4AicbuUKQRoXaD
AJNHe9xVPQPfP/gywRVs+Py/D7rWOl3Z0ul1oJt8DgmM2V6PC88Qkk5XlJvYjfeFAqRrpOnA/toE
RnDZwWbbXcUvA3ZHs5i4Ry+pusAkiqmOMw0wKvmrsXt+FceLipasdgQQjfYL8LSXJzH3r/RjYwez
wu9mJQWrGnAxx6Qq3y3HrLutX/ztwYU58HX+xM6eX+zVRLOYDNkudoeh5IstOYoSMXaKVjsJAwxK
XuASM2yjSP0k8NGI6XLEzquEb9yFIurd8z9yV32JHtrfWmynP7T7/QrXqwimvP0NF7eqg29CVuOz
BFKxbl+hiJHKr19vlpWmgwr5Izyrb6nTXe5ZZZ86vmRyUtjmKRp1WwitL2RJwJIyr7sYdzu1LQKx
WzrieGcTXLTVQhWbRNnxPlWHcHQyGnpZQXwfXdGgIaEUGzredLhUURE0Pgxqf35yiWVFwIFFAUZQ
W2yfgFue6hCaL/X2wsLmQzHf3qNhdP2U+x0aCi62ovo1AhK808swUue6PsAm235pO8k/1fU1X4LF
AaGmNaoqkxMNAt1redR5Hea/HP0KWgs58AyqFR0ioXG9H4yEITEbb5BsUKB2O+nWzh9VwdIu057/
PcukdNZbHf/BkCIVlbWFP0gWp6I/yM+fLkTc9cL23SRqPJISsgTFk8G8SH4YavEqbbYYqZG1+XTk
FHEX7Jg80xlUynRP3ndybIxrv36fXt3n+cLhinJCXyQ37qKuq9sKcN2FA98lwiFuBSFKp7+2CRoV
rUjZBnhDLcTBeDbq4x4/b+XqpxPxZPgS6OFtdvVpp+/MoXw+OwWjFBJ9IdtlRfLJkskQi2nDhj/g
GsH4wphzh+BUoo40LmOiTd75DjzyjtQYMmySvF2qan4W4SLKmuT+dXjiB7XScXHcpjoN2RgRVi2H
IYiwlCe+jqIOeqRv+E6XlL3EVjpM5yEaedM9MXL70kLUeKKp5B8H1nJfYH6bNZdn6Ol9fMLKX1PE
7H5UspWNkUPdp2km0pXE699XNowzpq+tf5xot12OUYo7oW7HSVjyZTXvrqtY7I5x4UB5XEAkjDXt
61riZ4XTpyqxMU61JSaWPH4RNN3YH++ZWarkWZrReNh2US/YRbb40PVWUBla0auJ1+eTI17gyUoZ
+cy/O+8GHCdNhRaIOCTJ4w9wao7s+mB3QbGwNOP9Pzs1+5TaDS5911nKmYBMWU3qVWf09ObG5fca
Vthibku9I6Lx1te7NbO6RXc4SSvq/GUcaW7wRXhtVGwotMAqm/go/jp3QU2ASwATVqVuUxNAOrpO
ferrexe02GDRMwGZWJwWZLJfw63+IOnoU4X0BYV8XK1BxSEKwKKrARN+Ph+DqoICHU7BzE3zUIbm
7caqcsK/Q7/OzamSqJR3cPk/taiLM11GcrV9cuWGVZEjcS5bmeTM2jFi5qlzroFVDO7LYS5xPhj4
3YL9I4dTjaLgJTCLeX2vzJ4xOQ3WaGw00q7Aw0VlOPaszNmHCAPZVqi/XWqMHa1xSPwWOuEPftZ7
1n++XsHKFcZ+yDLyXgy3u6NiktWxZPmWHwwsnSSRodn3KZKSCWmKDq4SetapKsTkNkbAQabjZknq
hqLVul/dlFr+ahX7Nw9z7E1H2rObRxh4zE137KKcLMu0zv7POvk//6MJbM5e6OD6RLvjbegyQVq2
yfLdiWjsb4TOAP7f8XmFSteD/Q8K9e08SOimNjc4pPo5S5TdAXhUVksxC4s4Wtp0FYdBWt8bTwkA
zGZ6nou0jrP8TDYwXSk5e+uqZaCaWi/Ilqt6PKwcjeXvJ5qUZ+CpTdj9erH6bgyU/UFtHdun2x+b
6+AFNbHGizq621675f2mAM+hsXkHQ9koHrBbUfK40wulLUyGH/epmFudtBhq70mpN0a+BQJ7FWQP
I8pcPWuEzlOpqzmfTDXvY3Qz7AFskYjEL54timkf34bmiaauC8r5HMDYvn4aHBynRcFDWGiqKOoX
2M6qrfsIkgPq8eg7JVyo8iBNPmDit7ZqTpXNBd5iglyTU5jqMBQ8K8tANz/vJZQcgMaTuKt09bMy
bfYsxtNj+9sAf/Fq2OqwwCluTh3B9rHJRWYagRP6g60IXOkDhniwWs1aiKu+Dr/aUC3y9xGBKg+q
wtOrWBAdV8OGu93hUidnX7pHJUbvbo6OX+xC5qXvezYh0GDqH1yxyYWrtiUSLsGxBaF4vq1ZwfLL
/ib9YqsjNF6eMRYLDZmLzDOQ6/z5gsv3axTLyGdAzl58eNOnBjPVVzRU/gQ29Ej0HGP/4ph3peWz
Qz3B1aDSWI9PQCJ03j6myrVbuvcBL/GuQAahGJ1XN0UVV60bjoqwJN/Crng/ZRSTNPNRk+ZH6y9n
V7miMSSDNPN+elDJNdQ2XJyNQMOe9vxRcsfe3rUw8mOUNzl6EX/0/9BiCRv/Wtqqn+DAodBf3NL0
RsQzwVxR1sYltPpCCGbUCNTvwv4ZwE5As9cUIHuFxMUURiNQkaDNXYMuU3vysusszFdGWsHwus73
8pCcMhFXXzwKYiC/kV3bJ0YJc5NeBXmT6EDS0kVXqFuBIJhYVAfez1dGZeACN90lz/Wg47uF2Goc
4MjefdOoJDDryYe/LuJ90JTRRGa4XoJXLw+QlJ06zP6XeDdmNRXt/unqZLGFScmuQZv01uBC5/fX
sgKwVjhl73laLBvftRn1/hPpR/TTrjwisxjXCMrGxwUVj9Czn/ZK/MrWH3FW14e/zHo7dcECzpiR
yAYrUIFdRLe039DkC+bQLtHMZJ7O7pCHUR8CmA8EvEnUDQMKozJnLLF17Vk0lNJ/44slDfWR/X4x
iKB0gPVxa+4SGvjFPTjpsB8egSkqI1uMcKJgYFEFKVlBYvQ+BqtvBcaZsuCq9poe6gjUPZdJ+9QA
EO21HfwznSmxHidakUGpjVsc+qw+ptaTyxYgbAKqdTV1LzeJ/R6O44p3KY65+MUKW3N32UBieAKy
jjn+3DqXNQ9GNQKlcIelc1pve0zQBz+5g1qAq0qJ4X0J2alVDKwulIrtfrCXQOxssISSMD3pP+9N
04PpMLODPOEH2IZCtYQWRV4abaguwYaaBWq2ns3b0WdioC4KiXaRvVb15DMg6kE6WSggf82NEsJ6
6wo/WlmBVlhtRqHyK1IP/Vv6NXgjEunu4lui1IH6xgSozqzzYH8h9oD53K8tYdUCCJdDK07qoqsQ
hLT0x3lGE/6a0Tm3u/NFojQ+0S+7CnPR6p/bxWErypDNTHwiRtdajZv9gIgHyhy7s8h2DOYN0suO
YB1Fk7XQhxrX+QW1XX2hKM++FcWNvXnhG3C79hwWSpyX6gbVwpaLE5UHpr9iWFVjfg9U1DqeYx3c
GQ+yq0Wl/dSmLpShRla1lDiGX3FlWH69UDK1gED/QDNlT+gKjh5Y6Nud9sLS+nSb6QPGIEPSyk5E
KTCNSJYMhIRNyDj/TzwbcwkW+IJba0gDkrkVE8+eVvkzKqjPX8tqI8if21z4smITqj/mPcEMB4uB
Yu/IIysK5EeWsbu8LTe7EG+FRHazLgpOw561JKlE1w7NgziKY4dpSara0XGyVN5TbvSmRUA68/C7
W4dgquHuB2wI9yqlO4rCqRCUvngXNODs5u+4Qa22JIgvckKn+BZBsr6CnOC30RCHDGuxDpgZUfqJ
1pFfL/IJT9ZuRTVTsUsULX9hoN5drPJI0wjuZSX5LFlbOiz339Z7OwgcwDhuiNz+bi2gKxkasBql
hA/+hOXBjKxL4mHDPiINYDc9/R7s8uIfyCdu9xhRAStPCGTPO++2RXK/eRS7CGkGroTAPaxAMbRp
tfij0NGPS4Wz2goanha6qCwnadFFDF6QzLc9fVJVLVt/0OKhN5pXBkyeySZ8gKZeJfyJEqniurul
IvtJd2SMZcsA6UNs3LUnhmwLA/hs2xHfiUtKuh8Ro/IwSMQIfJxxGwtKtqQunirksWqujQG16VhY
IkUrzw0p3IzlBDS6Jw+Ojf1/zPhq3N1ixkjQHMTYZZRD/60FHspXkkB8bb8oge+4o7v5qRwOet+N
nNubQ8yxYA95nidAWFcpaSl+6zuLR/ThC0FtfP81/3ToUW+L9ktzPlMqfGm3JL6BF3dttXnFpKVc
WaWTPoeWKKSqwr5GbaMRwBU/pC6VtRoNQBhAmr7Z9VW41zEgtyHedTc1m4fFOb0dDOrzrgLKMarp
CADvBfuZiLZixliHTxXfjciqcXqy7TQIW+Of0cndkaaL9XbXVUA0hACh7svw09Y/DtXnsQRoPtKf
d4xsxHbenXtxNuepN/icYBO5RjzFqIsLI1p3h4ocSXuG19mzduU6xdxcQXenhm+XLvOGqvA7kSsR
ws+10AefFw4k+b9FnouNDPxoRa+orS25WDp5fx5hspOA4JuJ9RKsL42UV5+05fHkFykZn762x74W
Q3UVq6lQj0eNt3f136FL+5Pm7QtRIsc8Bg1vWilvho9lz+wrxciAVvWN5QK2Kr1Yo3rv/KFh0VCL
+QnVkiObLIlpepW1ngsihIUbFEFnJCSIN3QjhDa37k3Oi2bD8oNagMx//jT62wuPjKnecZdY/vR3
cQ1w2VnBkP52teGsaE+IStEPejciOaC/bwM8Do289Y2Lv65iMj7FuuY72XtkOXyEelPT4iRSM2ij
ibECArJEdE2G58siUU9SnJwJEjG/zlCaBrpg8f0N0bcO17yaLTM51LVAht7BsmtjjUF1O+JbRZoA
To6MApaKuG9IyVCqixeQyQxxR17H2aIxXHvUWOp1KHsAbTEfIOCTlYonQBCH94h7cCBxEl96+3sp
E4F4kZQdLE8qwl2lP4nhQqtBQUjVcr6fM2SoOSn47UB8upYPnX9LN0pOlSeMQb/6NiKqMadEuz7m
EGB9t/p9IJwsNFcIVTQo15Z+cbWf0jiVIWNHL3SVVcnB1ndrYc8jRtnP0JKVN5Fx2fL2ULpHPLgc
kviHHqjOmz4Kv4CP7IuirPQoTxz+GQAkUk0ouLuZ7gGbxcpjhG6nE3gDhQk6TDx9V8zuvPO0Ec66
c7hePQWlMHKtS/BxbqquuTgLDRo0W6MlQC0yQH0AOi/Uud8LGnemDGHoez0QOx6AcC3H7zxfOcO0
PR199X3RrvHAvOqyiKOaOdrT1XZ+4l6Oalj3VyHduV65LZTrXpbhOd57zyw3IwzzHk2j5JitQdsM
ENrqnwoGCv2ElPutjJZvv8KrTAAvvgcwGrAK8c72PAbR4aHdPBi8IgxZSqW6Ztn9MdkQk/sxoxPK
Pr7q/JB8j68kOf0Mh1M/yg53q6v4eiYpErm9z7YF3twS7PtKMv6eVA/1epPxr1SHRmcHAKIOC8io
MFuWMu7Ony0YG9P6sHzZSAFYwIqY3BKRFTn7zwbMFGNL6M3YbKhNwJ3QosrQqDvb7iVMPZpaTZrI
nhAK5Bv/w5dnRJ/6i5cKJICXgmx7XQmA3RuiFQhWx3CXhd4cDIno7Owh87zAtimpbuQWU4/t5uC0
6JezHu/2oEqL43M1Vk58pQpWhT4MMvW3tjk7NAOEnygRPU282dC5vfzQTyluvgv17AKDCvlOYlu8
XmuO9FsF3aML+Scbf9BSmSo4mNSNXxlz9WKcBioxypEklB86n737AGyeYkHKf+Ssf4oyRQvMIRd/
U+9Um9pYNxhXVbW0WKVlxy63vdvEs6O+PTWrj0uO4Za7rPwKRAB1v/wNNvpcwzXw8R4yjO6bsf0n
UOAX6HyWLofTNJE1TxiyS1IiDkghkfnqB37RwW8Ml/Rc9xms8k0iuvnzCvInWOyLFVEiHfxpwvPC
0kIdlHSiHggtTUiNdMb5MgSOLTHUWQ/r5jNyGB/PMCA7K215+9Cb5fojL2MXfsBSRBKycAFpVsRJ
iqV6Kt25xKXv7dfdTRjawikzU5fOD63Q7EIbwymk8Cyu8xwj/iVcUEhRyhFM7sjSxjevILWLUSSr
2RwanlYEWp24SBSpZf+4QAdxbqmpt3SXystia7KT+JtO0P4CX+UIzcNyre3768Vms7AIT2JgbyhC
u7Y5jCjZbRGThfYGEJEag712FX3gPOhyPFVbR4lDwxjDFZdwl2Fk8wOIbpBgcICKwtJTthhxUgX4
Ql8Vvtz+FzAhocEGyonLv4a1RgnbvB87YuibRKIJ6GyOZgX+ehNDl+NRDwZ8LbI5q0+S9PLM3+ah
FXA3k9IwwusRWos3ph09Ok/kkJ10LSKmMAWonbA5su7gPPBWiIiqGc5DJTRAFDuxEyJWsbZby9+4
+ogpNUUUTOuo2h8qAlxoqzW/PqvZsolnM82KDbrwzATbr8EhAb9b3mA7Vut/U8aEdhU4NK9og+Rc
xa/guAqZ6GcCLe1gfVzjL0X+qiVvAT1Vhcqns+263j6/Gri8emsK+4ARBvDSZZjW8dY/q5V1EtgD
Koyn8gJUsPXKVuBjl5L6m2I2wXX6nQpgUd6x7iheE1srDRuDZ1PRY8Ppb4FdegdJ+Y3CSuA9bPHO
Qvuie5ATNrPpf15cbp3bfIsaQppVj39VSZK9kli3LaJLh7ydk4HJe6woZSi2//1VtITzCcU5eFly
LO1TwsD9+dA2wIs+4oKbcOuTqNYKpPWYU1n44u0NJ1FmnDcNqXXay7uln3o213dAeCz73ymKzZYd
pOy1PXv45QOdheXCIi9IdbVMGebk/7Sr4wWaRUaPJuLFCpz4bRJLfg3b+kcpi0BEiRCjHCBHWlaq
IGhxL3QtrAEeMAY6Uwk1hsXqvRhn4jGiYqufossJi9QktJIEXEEwKgDhkgdZHAgDBLaOWzYwARTv
ywWZdyZF64m5bu2oqmnfG2yolWIDetN1cmt36P+Joco42ef5C6aZzNMZffv0Wn5q5T0NSaeBT/oA
+1OXnu7I+blynxQ3VyWPFtZCEAC+SmRdkg5ITONwVSnZyRRh9Z2my+52ljkXMgTsfv7MsdPIImbk
7Rq8lph4Cqb5d3tcNvWPAuqjRODo2rdmQ8ib+eEl0X/8Fr71NDprtFyPBViETkZResYAFaxaRgfa
cJnp14S6j1/lCH9HDwv1fhSu8yCIidcDzraTBiIa0WrOserwyujSyZTxGnAdEEdtvHQl2sFnpwMY
q8lsPrcOZn4B+RU78JyutF+aBIHJ01C1KDIU3hZ5Gt5IrzNzFlGk792/+spc2cvefz6SRlLPTG4U
44l1tk+s8cDSlT0Yv78DBn0rtwnsdHBvhynma2oHgKxZ4nVQDL13YiiRyFvFXowXpf/oZtSDQM9R
p2ozjIO1Yn4pF+POvxTSkBLDs4BPYVj89esr+rAOfBLFRbE0PhbiZ3eOlufIfH4AdxIQXVwyF3xX
DoWbMfmPGDluFeSHLMJb6V8TSFTEDs/maqACw0f7QN0O9cvfG0oWYdGLAyJQVHGnPjNKrm+Hlizq
GpRQhbX4wUyML2v4gIPcqlb7uDMyOC9RFdXufFeDmXZnYyl9tV2wKUY+fzzKNyF/BYmRCbX5ezi6
4wT5F0FKAgw8Yz6goCnk12vVGoHrLr8wkG3zTCzpGq1PqQ8EdrWFZo0MEqzI4Qu07ZnEDBwn2XKP
lCHVZ6xHW/wyv1cy3RephDnUBaxr6EQoAyKHdNrtBhKqRT082NCCG7D9S9AjxIiDZa7Po2f134Ub
RdOSkfzBlvfiWM6G6bgyrd/fJjQcWvajN7XrW87EqrknS9r45Zo8QTAmA+m6f1ggMNjXTwybE2fz
xlmnkaS7uL9xPDiJBJhz25xc//uVXnERezh2mIsll77y53A115Tw4HYnCn5XCof4fWL3LuuItbHj
RvAZdwQhMl7OB9WhQ7gq/geOyYsZwTAvnT3iNrBc0w81CxEn+h2GuSM4dwDDnKUaOMEgIE+Zm9xv
+wH2MlrB4J6u8z3zY6kiKcFMUX/K7hfSC277Cuc4P6ZuqLIylAnny1AjvHfX0qgz4PL0JvO+OsnT
OkxNtrW4JQNtFzD+QRM9a02MgUcJb7vrzQznrJXHO6RwELdKWvsPg12+Ocr++/u20dRjZDXnDyN5
t33k5u3/CP0PfxBECgrF30smfYmkOtMuIiJuCnfIaEnlv2JgGdboh0rLo+TYzJkFNlCXRC9l8WAp
yvzOZ7Jx0OB5rWnbNjX9EWVOxpfI2K0PWIUth48N33czo6FGGgx5dgJPv69c2TheG9khzcPwzeKE
urbCLQYjtEz4AF2uuVe6GMa/X9CApZCa25HZZhLg6FvS3juqN1rB+CRL79XPaGXcRO8cVJIv81sW
l9IxIr9O8qcYPx/bcdQiFD8Jv2Rcqy8L3U1w1MKHcqBMNf0YACYkISlV/uxMdGsIvtxBZDlpXHqm
P912kM7NzGfqmwjFlGwo8ShHOht1yNibTvsGKKXeTX8bOyKpvjaXFKYV2wlVPNfoBm8w/c6n1y+/
RbPX9yJxvYpgPmZGM8LOe5TwidiT1klCIfdZVZMvZlJJgjKskTZpGCbK/1lfp9sxALngD4kJryJ3
sXoovQBDA8eIPieNwv+VMNeE2rbQKoK7ZW0PSisGw18k6BluNUWoFJIi8CYU3p5zO8E2Zv8MJg1D
gHtRMYTfdjqLonwNnzASPJNO7S/hPeMfsNGQ5nTjnuG2CpC/ri4RAyxNEPvMLz1HSf3QnnfNnMgn
QjwtV+Sq9xF3ZBuqbZV+QnxLOj5m4eUoV4nw1omVTdjkMG6q8zNjz0ZlPnNhztsKBaS9uPmkBOA0
SFgkPn6EoAXR9XUnuAD4Y+uODs8McknyZzdRVJPzhvTXIenXphUREW0r81F+FbqjsCT8vvftQe2i
a9N5mpKRptqrYBvsFf59YUSku9+yL0XgR99p6pm5nopvaXuZwhyUhk5aBjrw//PXe536pQLvyY+V
iGKOaVwyXxYaJEPFBfwEK2QKJv50n0m5PqxzH7J24/B/+gLIxOPIkCwydKTzJ1DyZAe7dX3fs+BK
Ocba7SBEkwG4yur/mINGgWAhJkqSUcgxWH2Rmdmnqhjc8tj0Sw8qse5iV4UOp69CjnJw55yXtc+B
IRkm6xLiTZuKc7cHz03uenszv/HLGpGv05H6R74JSY46k8qYDHiTpcQ7SYNvK4S0z+F6wqU9cJNq
Tg3fidJY1KGJSEkEQ9732QLqyYpf+9Iph3D99ncrigkJSR7wEG3XKnI97RStgHm+0iTW5bUTsEMm
heZDaO7LikrIVyWKpRvaSsHUYPQIf2hFCE8swWW2evsXvRg+86RUccNAjcTGaMLFYXeTdP3K0eJn
IYSCFi7UfRX0wJ15Nb727Lw+gGhv3Zg4z5umh8+7DynQwl8Eppf7auOeSvIXkUadCX2QW1jdwPyW
nv2HkXh78SW3APjtfAZRtFLeFW8o5JyazaDYrR51fcCPq5UyzfXgcM0T6r6s1Ls8ApQDgp5ig7mi
P6Z3ZDgogHwTcJhiXIuF10uUJWsAYPwyI4t5QChFmshzRbUY/VfzOtTpDqmHfAxwkajU14yMMWp3
BKnrd2EBwjEf1NDHgZBUkikMnjXQ15UcYICelMiBuycY2QNwVXB8vywGyv6tTsGjkFZsq9VeO8EO
QUhCyhKAl857EjTri14lvVN5tbrgL7/R+sbp88/S3PKTzM5J85NZiKPeG5EhUJm6wk1c4fGFUUTv
XXLVj3+r+Kp9oPwVMe9stlLPZlZ2sK3J0/SevhWw8KQa/PYuHKpHlci/t7JbF3+Z/vB7N3sxfD7X
qSByPI+csGyBq8UMOHvgk7aqQVmyuDuo6uogwHkOuv2Er5g6v8E42aOIqi4JDMn2xv/X5Bp65Onb
uCNQ/gqrqnftElBIQEzOgtfBkQYqDlMoHLbAPU9k8XIuDxUNH2Kxo8B+uX4rfgF5cE4YmsL4zB3s
BEABOMA5XQVsN3pm2MN0bl60kTFgjmq6sC5I/yeH2hLilSu8iMvhEX/mMmm4gIAJW4AHAHE4veH9
DQRnFqMWI8WSvb2kg9mN7tmc/CwUZ6hFopDw1rhBqgVUpSuLMxN6ttqIT/QS1Gfbiz+BPVvPekZx
XJ0HXIE3Y8Tg+dOYL7Lc+MgYu1Fv94GUhFaXoJcdCt1jPoaX7Ovh/1ntG0RSrC6rQjWOF8rNkKXz
5D47b09MsXAE64lWCuFXuzQZS8068V/oxPrAgyOWFxrM6VIyoxI/kOciu3ZyQZvEdFLdE5t8z/rN
s8O5FvD0XBYuPh6OvK9znbJmEvhTopgoivCKkS7NRXVuM56gV0fjQhKqfYAGoG0es8Segm4vM4JT
es2xE/OxoowU52ZhDw9WI0xVyYxrzNVB+V5u1cBaYJlWBCEkG4L8Cvwhiv18Ecaoj9PHNXCGTnrm
R1Y5I+q0HkNSVYMHv7AIIJnf2t0I+4M2eFaekR4lavRM8xSElFDJjIl9Qs8zFfQBKPnbx++ptb8W
X1YP9UkOQmK0FSbx3Uc98nvNb+EO47dHPXgGMDUnaoXHeGrG6fOIOI+WTEZdVU2rQhCToL0YNIy2
Ektab2q6g4u61Y8Ne0kegtMfvT3mtike9tkXPhoNn/hrBQA5alSfmBlPhFJdd5HNIPj028gWR5N6
VljFu8MEeFfaqnvMXqqzAJFcxF4tDGYfdOIKlUChq3sP/IIlFQ68rvYZgxYsrGs1nG57auXSM4NS
buyR29BRoxMkYXwkrAwZmoDnhPgDys4+T+s7Au0Jyjhgd18G+/Xq1MpdC9jBpZThcmmWd8rEu5l+
sodXO/x6NK3hOm+7a1eg7mq5uey5RKlHPlo6+HJn4epIXZink2pOnqQYxLZsn+kqwPX303Bzeig2
pjThQOxXfF8sKx1CYDp7PodrJN8LnznZPNVEIcGYtQAPRArfLo9or874hYO2ATef5udHlggZWaSY
mWiOkrzM6Ed6Zi9aT+vVJT90EixpmqTNNuWrqnLSFX1ziRHAbrvYh7K/3skxzFhIOtw9wc921L00
PmnuJATUJZ43hYfIG2yNwKPcLTP9X+JRmmvH98Obs7AmcNGao3Hxh5d98+WAqhEF4/ud8dIDX12Q
IWkqfJeWDja7dCdaRGXGTDJyAQjFezb3epvCPseUf4cKDtga7Ao3Wz61Cil95Nj9hcPDZzc+3Ssu
JtBGV5maBu+GnIXDNCMAPXVi5RBqXEg2SXZpOlvV2jH5K/wo3e3Y1Jj+8vYLOH7UfBChJldOdDWi
RBdGWc96qeLrkrvlqbF1KeMzFK207dcEnWvnaSu8UBObsZ7ZXjuanNW1nF5ei6O4Mw64tR32sojS
2YoPI87Vgh3uzSmlgKj3JEkKAIQynSuz7TzFfwipSZCbWJzGfMDSH730DcTbrkp7HjXYOsEs2Ctn
CVXmxv+j3XpgfIoYS3Ni8PTXOAOIXlS1wopYZTK8Iicz1fuoFPKDucabTPVONebGX/j2kMbHdkh2
FS7imt32zKfILDpSmQ30mP9tPKaYR74/V72BDt4W+jZM+Nik/x6xPXCon5e/rkGENT+F8KRjfklE
yi7VL4G2eQ81MS+j+5TJ9kFoiG5puJ3lTACoqDk5PFpN+NEAhrlIFfrcewPogb8T0sbJJx/2E539
dqVnvYnsVdsuxhlWgwHZv/ugbKKh91Kk1dHd1CPWy1g1sduZImcApTp4QCn1PbT56X4AcZAO+sML
pap2yQqNDN8QdQUYkkxboXRBi8Bw+SHuyhS/mQWSY4YjlF9KhSd7loJfrcih5QjzcmN7iO092l1V
76KXFrUjg2nzZlsba9RLfHKtYuWespgayO+BNfb82HJnrpaXyGajnndLXp0nExCT3nvh0qDFeNGA
wncx36rIgHP5rjSS5aOSFQ2uAnaig7CHHFFSQU5cpTaeFkeLes29r9xMuIjEFH7oE/rLHMiZ34jK
OyeZkFBdOEr6y5JR7/atJqRlSbdw4WzqhTD3QTVQsQEZjp1QGItDIJg6FLpd8LdXiy69FQeTPvj7
kzcCm5mz18HZ/xeBuWMPuZKrmJ6QFfFuPvupt0P4HPJeYlzxYkJmmFTLt6Rbr4Q0Si4nsN58FBNl
5HvARxTGkvP8bf9RL2dZVJmbSGtMFD6y16So0VPWrJbneH1gU8zUzfTtVJ1IlpQ5/rlmVD6VSw8K
HAV9sR4juTqXPxFkZ+mRORfMGZva/MReOLMF6BbQpop9Lz//0OezT/sqgvo+zet9We4PCM93pwmU
UqNAnL4VRU4742IY4atURBzhwYvTMHYfYAHxbM2JaZXrmtpY4m8y/oAf68TjxnHnThl2oPgQ/gBT
VZ8Ak8yFaQnfRp3F6VwL9ZzverPyhnmdnrLnu5mikQ5LQygcj+jwWDAY0uqKi1up/0NwERi/R3Ry
8IZxEFNMhMS6Kx6SYYSPFb+IWKQ2fieCCtO6AqfYgwkVe0jSYrcJCAG9jLNOQCQJwUWjQJN29Ad8
5QUSEtesS++WCR10Avkf8u1eu188lgXcr1rmxES1uqXZnlN1edR8nFAmD6GW2JL8lQAf+z6jUQ2s
Nm/tOLdlpNOqyEHjXeuwiUJWUSliMWCO0dr2uejFWpm/MWE+1LQ7dqM7DfrrcNTvyqTAEKEH5cR6
J2+72K8+CQVdR3gwCTi973Seq9KQ3OQCTBufHWc908wQKLFpfpaVHcZc5k6A9481evbBi/jZ2l9N
ps1kbCnOPNh2rGgBo0h0LCOnAR23fA211uKfkfLOOrFEdZPYv9CQmlqa+1BcSSn3mlDCwQfI90oe
yVYLUyACmqn/s7XKdolBknRpeAYVGe/Ws5hYE/py5ybl/1hvN6iT2Pyx6959bzqfzj3OfoY/l/n5
lnE861CynjG0psH+SZ2WS+8E4pANUlzw7fbT7YBlQotUdDorpJlCElWtm0mLl+MVs+iVczz6gsFO
ng57ZOfEFD1kfchz3Exy8tGb0u9dBZal8KRAMTD/i4PcTC2sfeyLXjTk0emtz/3d6jbZHoEyHdrg
dsf+uE99+Po4YEH6Cbz4OxkXjQ9Lvw04HJ6+lrYoV3eAmDMXYtTIFZtjshdIuIRBo+e7Pz6H5QKi
KCxK+ypZLsz5bPZt9y6Y5nlt0qY7sZ245HNYurSYvvq8gMOnlxFvGexHv0vUdKN33NNFHkU2ajOj
Fam+cm82l5cYF2gER+Sl355JgpfAljH4WLE6nmOtuTtIZ0YyPj1Du187sReIT5OQmLo6KKUoxRvg
xyRiqEsF2Qq/xdWUepbwZbpKL5b3VgRRm+cOohWtMwB5LCJp3nVjbDJToYhHSrOI2qWOXTE56tbP
rdIathYIbvy4w/EzVZoUPaf3BTPx5/X/AXciNQ6NpGKUqHzX1Ke1M7ywCIMTUKqcRTZctgH72lVC
w9DjaTDCVv4vh164fEp4mkGRm4B18t0K9cKCrEFwdV+4WduVC6MXu7hBC8Pxcz9qW+LLTiHlngRM
bv3ZldHvgVc0ceIB4pIOWyMAQME9JSxhgzqENwI5McHTbwdHYQEoEsSA8/iWs6aUvNEOhCWQO2gw
xiJhu2y25ijSG1iODEpgpTtp9+ZTYXEHO8BZB8cX/hNurD83aDWcYWoqe3DJZed2QTORwkGOwJRk
Q7uzY4lVVCkNoGdm74yK8QT64Xwpz0jwGJ48bKq6eMnVIB7aglIQn38yF9SkRFa4kcDafcyi0G4F
JvKeoAJg4oEUGEJllXAH9vzoxCQbsT7zKXEkwGgoDIBzXso9eLoGsJdDO8XcBbOVMI4vo2BBwCLs
QpTiSL4/PGQMWMKHLFgQ8lEVzbzan/YtfNRKKfaQQ/eTmYY9r+eMldixILVwF9npwAhA8frfldyX
SPI5H8sIzkcG5+OYIoctOy411PXHpHDohKBonDKfN2xLCi+T219jSglUhsd0d7Spgqm/Q54Zrv44
jiij6U5m4IWIihULOiUvOUbgk4E+7g8iSMtx1dcyp8rlU4p94UjLQJKi5IEm7wzqP/ouvZiZAaDJ
z15u07W8bHtYXwcNDQ8TSeqvB6cZ0IclYjl5+8RmgWNGRDXpbt1tRcotEze5PmuvLBa2yV0bpNH3
DHNO/RdgbV5IpAgfQ9SCNutV7/1bmOlUtrlncrM4AldwIyHSiHBvunN9fc5DPxxjzLWw9goF4T6K
kmnW29U0cqc2NwGkDybNCZBm7Mu89QrCXftYzukb0KnJoN9vM4P71xwnjr/Csjz8aF9/xLQ+EVS/
T+0fsAxzeqyQv3xBRcvBvU75OiuHfCKU5wXqfjH5SmV/jIKVba7/iQEzB9er5lL9kdlo/TDKF733
VPf8GK9zk9kC/l4gXpIq3fjcgqkTSI8BpWQPmtKRyWT41dKbN6GNAdKUVbCNHTb0dzVG0Ia1AfE4
UFbqo0KT3/Ov+tqz5MwUYhUjhG/UDvidfxiXx6BeL3KGDgCQxaq02BIputP5YeG2yuYOOC7QOLUv
YwnsiTfEodFPVhRmriItcHFQ1mMLaqv6bbMr2uThC/HY2pLt3ieFI4+B3URbTYoyFpGYJ2PZ5T6Y
Ipj6X6hq04IiH2eb0Kabj5Rhglh6PcIr0KqshGVK3XJ9KiDDZg1LXC4Xv6cxI53e0poNAPbZRXKJ
9UaBXRc1EAF1jLZqIvkKO+eyO4BTbK5MKgMbqlwe2nLRYTC1DCC7cHmFZrEIuG6ynE76iJ9SPY6s
U+mLpNi7/fyV7UC1L0w4TkALHk80/jAxJS7ur56al2L/mOu1OvaVkqSKOBDKIRJhjtgv/pm3iUFc
12GYd3WOYflRmdFxmUi1CzPsAazfSlEkMC2kwH127LYEn5k0XYSBYsFuDn8PsYXSJ1rGy2A36R74
q9lk2bbHNmokpf8V8SloboztUhTTLa3WNmZIZGlucNypM7uiSUE+EQlRvJiWVEuvlNjEKhzIYY2K
eKh8KCiyLdN/8NtK0uyBN4Kti9/RJQdBM1mbogS1fQ39IbqkN6pGGOBCNO17wfCX1vQJ4D5MPY/w
GORW8wELUwhcCcCBfXiqW43qAnfGL+zawex//FKeoNAkMLlUEKkAqBEI7pRPQH4T5XfNqYKwPAIW
x9r2m474pDqWmx1Cva/SkBJqFs8Rzi/6jodXK2svupQy7hQ0KQgnCB1COJvdgAgWAyNWDCjLMNgq
gwfiBQWSaJNK1EqvxheK/h2YvrjFaL2WHRkW0QFFPLz5PrlPLWm14MyrPEOnD/sii8go4Nbts+1X
oHjNhUkBXdoHD0od8g/RZDjKa3T71+YWS0GtuMxEFNE63gkhbm5XW0Tqcp0VJhLns173ufDiPyXx
ZGBzijFBqycd+5Z/cPRvrWYp//Zf9Plbu4jm2FHoWsyNhbpvaLm/uhzuMdH8BJPLbquAIQIOlqJY
6QndljGTyPXnKfryoMpi7e9a014x6EOPl/k/otTLwN7OAdzq9HFHS5+YnDhAh3w7xNPyG5VyjqZf
r622vxSrRI+axvKy4TLtRjKCGA84uL8DvwCYXjbBYfbV0cIiqCP/Z5VPbwSeHoy7NuA5ABDJ7uW7
C8PUR7ZSEEyCvGmfIgFSs7VRwKzm9Bs7h0fQDYJeibSqlBNkMoTGm21FGc3pWDVETSqa9ZnYTk+W
GjGSQXZCSHnuleguOT2eTLm9gSC9Ql3652sv0St3YIWsFt3ONJ27Mqg+2OoMrm1NjX3BP/z4wHQ+
zIAkizX5iy2pXa95F4j+Bt2fvIHGn9VA4S+eaSKzOSQba7rlavnDlKIjkatj5NO60TGPgwSgaogA
Yms3MLj/aaVEzxwOsJ3CEdBjS54RgAAsqcvzR8tyv83XvHMeYm5MyBrTAqGyr7RQXLs59c3NNj+Q
aBxAWfiHCOoQv2ATHZ7ZnjT0EDKLc7y/slTeX1GFGv7MCHzxBTuJtnYAevGN4oPywN1/iBNxGEye
enGqE6z5BD4dHYaqm90q9WR6JExbcibX2vGSRBd2NgqLv2pR5+FGeqv0afmQ3rl4oztEYN0in8yH
Mb/G+WyWqBGaZMACppV9f4MWOWESxGgc3Eoq4zjBCp4b33UM+sEyg+kkpc8jx5Fw+koOxP/FuXpq
qQDvOzSvG01iS/vKu4o71zF+v/bnni4dHYZhSjN4uw8wIpe3dppwViVxbWBmR/6TrOU7Rys3czuO
uPjjzNgYBwHhlILEhAHVwlZ+y+rn2VZgeq5Y77h3Yp7sxOw66fXw84IpNmsUTP01f0oyJYVieLDF
vuyTzj/j7StEwmcMyUcOpJYVlLNKdf0IFQfxupckzA3jAtuurgaKqVcP19X7ptedg2zamRXGDE/z
kYXwqscyARrSyfrvyFmd9FfHJsSpz/U5GRqH2OiZPXkvog0H0cKE/Uz4l3Ak4o4KxTKZBetRchcG
OsCFmeoKbJVSG1B4tW0kxWPai7ApbOf9KUIsSjQKFT3CJi8D+WcDlf8Lsc6dEPoV/r0BF5xoMjdR
4ehxgb/nFOlTPz9YnDdL6l3WZWbwV+sG5/HOM/IYWA2ZsceCqiACKp4QFR3oc8GiV5F/dMrSTreh
MqR6LNfRC71H98hRTs3dYKdDrNRfJW141odqHweW3dBBUIhydYW6mHBWm1vJVJVdqBIPVs+XQuvQ
vjv0GBb7rARhLQlxb/leuysGYMjbirU1tvGS5aMG8jSOdOKHpzxh/DimWs2PR1a0LSUo9hyHX3lg
wwu9geWUB+t5xs7Q0yADNnrbNztNCLQlHF/YuOBosLSlMghzmuWAsxoBrX+xpT/N7DBZkXgBdAz5
60ntBC1+HQz29F5NdCt9fE0ksG4GkYBJYvnIXHQCPKTEEJcNTz4cBfqgGDDxJ7dEWhZrmU7CFA+5
Uvqbn//cu+CvDhNNm1v38asQU4rA7MaHRnnXCZBA02cCdagizcwqzbGLlqxqEV5jdisFcvIkMGt+
lWoLDw5clh+q4fQyKwGt0q7Yr3fetWSJi2J7gCKANf2iFFWRhdOUQ9p6aD/nWQGFtYQtFh2WchZz
XODt6kWUihefajuknlfAohQ6XNWB12x9Mdvxh8yholCiZh2EtmADgzC0w2/gi1QSx8NWeBcDID0n
q5fgMfI4NvUjA0wT4OaC5rybZwkwCVyMxke5OAnNpOgP/vvFRacwSKDiFgPrnSCAp/ekfPi3Qca9
yvMdK7fBk2nxVBAj8gjtXcZwcLGD68hunt4X5f5dLPbd76bjI9EGR2VgEHuUPdEith83OWgaEDiD
4soT8gGLy1HSAKsP1WlyXGiu9uXZ+qFzABJ1PaNDm3vkOiac7M9YziYJ5fIQ4wLL8heKiTmliW09
Mz8Rc/AgAMRlixaUbK0e1ksEREJcgghHiS+dQL2mnXhSv2heYpDDN9hhoZvUz8Nm5EINjpPPXpXy
wbP0i9bGDzRr4Q/YQixVgtOZW/V7b/cpjNJGiOhFnyT6K/uYmTPiKiP5xRLL+49lJqDev5h26NNk
ybFYoRnlIkyBGJJoSiU726eN3i/30ZEQy1uGmjFZv+qxTKgCHct9nbtwruP8N40SN922ffGqxj2Q
f/haXnahg6e76fRnZdmQYxjoagap9UJ3kb8FAqqoyTSaHlFy40EPBwjNmqpVoqksEi6F9uL6El+9
nio3TCOj2hwZ3ykTUzHFrCK0uzC3YmITLlcJlXxpj6U2JgFlWkUvUgyRnVfKk9+7GMRQ9sa90+F+
tWK56iDmk0Lm3/okIePHnlVfFWDdlqIa6SLKXjdIxhJnuP2w4N9IHOC0q/AD1KigUSBQ69acH1Rh
iisMSZgqrkhSvckFIF1eoN/NmYsLWUDNPrHFWo5ImUoJ6JPTPV72jwtKpO1JTpOkV5UTn9umW4v3
iS6cSBCrz+3fHzoc3FduOO41egIf1EJqbLylol16W/74ohCfKZbhH5VWBubfE1xRRGaPOhUJilGY
PplssOMng4QScMK16EQOmV4XSDsCA9laIfvMRIaTuriwqa2FY4F4G1K75C+Ta/yB4aCZRz/Znpye
z4hhcN2T/xOf3SZRSYHL8B+K4QFeDkI2eHoCY+tURAsqdbqsWsVKEmTJUKuElKE9i9Ms0Jv/m2nf
/0uoU7jDqEA4ogc0LTgDMUsXo/dZsU5Cndy7k+Zc2zrrYQ/a6lMbMQWK7KPM+iAN/QSk2W09WSqO
V7LsrLJencb4UzdLwvBucm1Iv51eJE7CB1XftfBEjGwaHNJXVOA4iwbzNNinm40+H60ZKk5+64b8
bZxeZbyGFGno7cvuUMiDGvK6YcmMgamoUwS5ZsxhVqNObfl2pRvhXJLrT3RHH+TSGgtnxa1La21I
vj3utlAxjUA/KloQyzaAN3Vr7ddUorF6IJwz4Lbj0VC0EkLtWJCLSKZE+mXVvRv/KWCGsmTf7lxA
7NgB9JnAwlP888qHdgQK1KNytA/7JOBkVVppD8euerjYfjLvFbZuE9gjWBBW8j1DvoK1aQ8Oj0nz
YPFvio2GNqXrbYHEvWtXaGdtEJlYh+99cZUJByagiLmmtGTHjwRJf4pm2VVml9+MdQtX4OYbWfl/
sD8oMu6T3yX/xaVqHBVnJpurKl2crhztubvqDFsUf9PCDZ88xoRac+gMAmXxdF0pPzj9wyc0oN0N
Nvfee5xRzW2SbEQDfrbn4yoBPn4r5wCqMcMOgyTLIOWXKUYa27dKT018D+4rTOBZG8sBSZBDtwb6
g2NquzyQzuzR9YrEfv1NM9VU5HzH6fbpXRwTVIsEPeErQDu50Q+CSO8YxaQOVNsOzwnTcsVUhvsy
s6DcR54If7PfE8g929AkUyc0OJeC9OVkmDoSdhYyIVRKxXg97xum4XYQwXh+U1LenrMF+9VXswqh
2xBkGP/DNkIFYw8vs0gUdwj3z3Zx0h8EbIux6oWnjp2URcm5pF0ncUZWDFv22RZrpsxNzlgJNZ/G
1l2klvimITp9qvLyEEUTpsYav+eom/D+XHV782uiom4j5h4JtK4JFCFeboYMHVN94BM8cWL3DkGU
2XkNZtR+02mxsne2YVXRktgMHKI5n6XSJ+TO2sSRSgIYeC9sHzTjQHsGR2se8tkYo63ZRcQZ+DpM
eFWnA16wFOlmuRlNSWRV/Rv0NrkK1ukgSz5Txysz6yMIxeJ8vZYwLCsMBBpCTXXhSubnkMU1g3j0
Wf9jSVsoLRqFyrHpfBm/k4hshU1COl70CSM3IAedhFoMkrf/AkdVLo7UWId4RdtikwSAQuAsyNkH
QkRKXnh/hLjvXukNo+GVyjHt1dip0G3WCq+U336loKP5XfTMPKDjX7mCjpoRM/A2a09JlhhiP2Wl
A41JUXLqgYZ1+LwSz+NZZzBYL3X47w9xWBLvABYo0909WA/+fNCws9OsVhPltqYWhZgceChzbP6+
iJi2bc+hW7VVjuMBFOECoIhCmYUdztxC+9X5TxL9/wpGVQOjrIyaAAwW/PUmM4lL/B0Ik7ZH1ekv
Oxdu6ozZF3GIULVa1E+LpDoZRerABNis23EhsPg4g9sP7QiETybcpILplvbaFc+8jgvGtkYNlFxL
24hGCU/6rGMbR+1QytBqwsUO34wqIwklWzhsuVg/Z7tNpFoomiI08nUZ06NADqY9dZuTquG1qy76
H/dauek/ZOkTYwcggjSBJu3GxqQYeP4sWvD1+jTGHhnqZz351BGhJi3aUqgOMZXC1LQqpJhk/Ozb
JF9N/1ca9rjVBE7idXBForilMUmf+Py7K6U/G8C/+NVODzMaKQwUap9703Es09xZtlE+1hT88zgP
1wBH7IbzkTMburKAM9vsa6+aXhPAPTbyGkXC8AQlC6H4g9k/OheDxGf03esLRQMrzBC1qb0W0k72
qaWUWscmp/eccV3NUSl6R5ObuGg/8M5i9fabr9gR9zRWzWxQ4lXA95+OlmVEuYhUSC2Pz7o/5Cf/
azNekMZDjoAsIqcDi+vLnDsW28NApxeVPv2eduwZ61+VISYLdlSl1D+z7azYW1jk1DEyj/MkNVGZ
6YRwSqxlvrIW2J036NF2LiwLverpF4Modff52kxicbauPrion8g45Qm/VvmniQR68VHKA8WQ5Kr1
Pz+VGKiryIkuDKxnEyF6qPAokeusQ1yjEUoHnlNdv2SWmgwpsDOA0VkhrDZGF1rrdbacb652U0lD
ll46gbej/C8aQvn9oM4VgNjVy/gk+zBRhqJcSvYY+MrTSxacPqgUNg/ckGBCKk0rgNWiXeeaSJf5
TUBq0SiS8JzypHEqsp5SF70SZYYau0c/VjquMDM5Fm9Ii0dvwuBJoXolLdpHNCOXYqmDbKExW/Wf
vL2vjHsVFbWY4tZ/aP4LRBzw7EII77NCfHKJAM6vCkoJRK8rQmddl4PYJEifj0Ho4S7NNp8EsoME
9D7KxCbyiVVsey5q9CNA1J4yicZqIGvmYJbZuHPD4A/YoMHE8h6gZa7Lw+xf6PRefRsvQ+MBzEMT
I9OztHl4+CHHX/lY6eLsJ03/rYMoFFWCNgj+ZAlol/nDe31bhWDdGC2A+aNkIXuP6FgdU4DtFxDa
FfwPshXlSh9VaMIYz2eV58E+R+MfPgDkwMmct1tNQlVTIhw4j/sKV9gi4vQc6FtY8LBXApKRN3ng
bev8xTHZc6kGxywDXAUlr4U2hEkWG9lrBkaVsWOFs1awX+Bv7G81Gjad6OW/v/tJkMs6/CwQmDv6
M4eEsaYBkhG70qduXZLHg9YIqD50F63YxqIQjiBab8Qd9rqV5SeHpty9BgCPDYbUbdiaEpCyWc4V
FK6oJV79N53l6/WowxH9tfSJ5Rdg/zPYUuzTEXdnw97JqJwfdAP//ba4qS3cj4g+20B+QEte7o/I
x+xVM1+4DbiYxMlWwsztUE+yxrPb2uxX63M+Qa4Pa8nar+Sf7++ygTzZbkWbHsOA5WV1zBNP+XMs
G2SLidgSmkgqIJIiWtIO1Ku8mkkOIbN1Tl370XqY+vk3DFxDfvnJuuaVx6n2sfXM7S458uAHhziw
YRhd/ON45z+GgGv0pXnm3IViYnXv2G1bzcHPeTG3yABVWbL31W0jU0ouNL2S0T8iSEBk1cVxDoIl
6Ng1zHoPnMVtiKoRIQTP+/jp8UTHE1uqxzIGqdeJd7sh6hkHiT1KfPU5gB4noUU3Y8QIabtOUSgF
EtxtiTDQWGpZoiBHy6zJPj1uCsU4C5NWunZTGS71PVh9/8G02ey3d5PG4Iq5uAbk01OzUA7pFdGc
4GBBw8ImGNbmwtVMCB5h/pfpz/TuJ4tAxJYouITkwNWCRBP6QP/hOvEO9+zdJw27JGsc+B1ekjvB
iwZbUTgD+aJes6YHT2L6L9BS2UNeJRMcGc2SA/Fx6Lal4HZF2o24BaUKUGxQfyEj2I6Nw3MTTAT0
IUxlHBk9u1AMdgYwgGzbYHsiFxclRnY9urFdfjg4Q9btMnUtd6vBPTE0llKPM7DsoC4YKEFi7gOj
UmWOkoZnTyq0L/7AvNo5VGlIY1loYzOKzlce7AP7tTLJxwoE8NyDMaNhXQN2WFpjyP0gXHpB+oA7
c5Dtu/aI6FNex/c4GSiCoyB71IM7wpHEVenox39vlQBljCfbz/7mCchC9PpKtg9796qmefQPgd7c
7a19jIoJzgFHSnv091m0C1BeWZxI11t+zlPQDKFbVkB+mFfjTw7/1x7wQk23/xM872Ukqpk6eKvE
EAz51jjWRTT1D7T8K0lrluZHw9pVdcgy4nJVTyWSGgssEv0r7E+vY70OQDX4Vd4Is4N5oXPhZBJX
4vDJmCuUpnO5VPEw3rsGePQ3bUmxQUg8SM/D1P8ayDUskJVRQDeg7f1Zm/nlPzeX0dNksH5jWwqo
DgQI1ujhU+24C2JpIvdHPXANqw1Ubwgr1/XWUbEIsZQFKSGhYeXPXwExmyTdq7GPn7arBXncCtfe
XhSYA7BYLnjHynyWcID7Myc/PH54I8ecj8btJDH3Gqqr+LhdzJkMS6mxz4Ym4Z2/HeJXICScEK74
J+KnDneO7DIQoqim98v/OFq+HBdod1/UvakOgdPrcYtjPN9VSQLP5DeuufmL1TMihMY+2MCwdiCL
KiLXvGBWZvaoO3+iXnQoPKzJaivEkWjL3717/w9e1fah8m7Khdt7BtViV7sfNSgR1w89Vuifn+RC
iGAziDxMPL9sgdw1n08gFE1NuSnJ7ZdLakn6O4u6GsvURIXgCJ4m7OfaTXRKZ5D9BO/bNH6vCJko
v1HkDCVmlunoNMcbUn3M1ZQw+VZkZ8QpaJS9ZuPjH0HbEDRiFqXdFZtxjFF8NFoXkvsmwHQNtxJm
AxqHYSAoI8hfaTqGdEM8AnmeEQvRb7r3mh0W1nIvrFfCfIHDE1qawFZwrtjlNCoUYXwZvq9NvcO7
KQfMLlBTDrpsLlDr3qTeqvNYSrIwsad8XBqlkqx2BD5MFW13zBbwgR/htsMUWjpT87fNSRjHI/2b
XN8Qc+yBc9Npnu3b86uuIKdmAqzbnyOLwVkTCw8FDMVXoVvd1DI2mlnYqle8kPXO/fBMJy2YbQLW
aDNHrn4EmYsV7AJPBCkb/d4LWj1SFM2yWigdvCq0syiGgYUYSyY95hXF3hm7OzdEUstt4HatMlHD
4SQuBlgaA591WOJ8s32w5vX4W7gE9ZsTslnnfU/gKksT9cBB10GMqkd2oz1x7LQepDmaHZkoZdTx
G+9bcSy40jpP2Xb0Rc0eIgSE9RyJrtELHcsh/iKyNPc4YwXfgbaW/wFUVTy4mmBh+3N8yKhVZm0T
FDc3I8Lx9UcfzVzYcjZBUTV7SyIQm2+xFK/oGX4lyPagCb9+Il+ubsELWXwzcbz6XdZEA7oOFcVV
oJ2MlxVwj463CxI9ENpxY4X6vSA9wMNgULQSpwwS8nfXcasvZvoUlkbP++iSe2Sqjv5umrrAEJZP
nlE2IanCUYMG8P4083sggczevprHgCuPoI00Ojgkis6MSDBa1XP3SsH+CeTd4WxhsQ3tzzTJzvYY
wzfsjs5ihQSwiz8IMDv0/qz2xaVvjxiN6YujWONeVcN6L+ZrTFhqsNpOBbNd/orfA0n+mPej+JWS
sRvzUxTND1QZ7yMXqfS3dLMEFDde1dx4mnOMxRPeq6Di5BGZC8GoQmQMDWADCcZI9ud9/P2i38vV
kssvhPF8kcK5umgpDJG02lfjmtW94vesjltdB+DrybtuKSUeJTm8W9WotqcKQ4HtGyr+XK5oAHyl
NT2o8yIoz18Kjl0niPOWWxdjfSkAQbOFDVtRLwwFUaFfxiLk+0OCYb0fP1wELoTDrvIK26kuMfyN
7PM7s3vuWhT7zUwLq3I5j1wsqSG/cDIdpmxTwJB6ETLFPq9CczcFConwjX3OtzLWvdN2eN4oPPo6
Q/9xVz+RzWt4xe/M6ioODxuEoCnZxtF/F0DDHuwSvabfaC7N//NIpGJVNrzA2mCtw53vtwTfeah8
52CYc4DfDUHU3S0ZaXQXmmWE7k+9aPkKwJlNoNRmYjkZI0+9n9pH2wb/WlExdVBxEF+oS5GCVjGq
qZ8gaRXG/EqbbitFR2pxwim3OCfCGZme2Bh7r5TWPhm9y6QaOIo+lX4cU5lh4GDlpMojNlQevklt
GAoqm6q5KVCDg0jCnb/WKLuoNLMlVI8Orcii4Boi7NN0+mVrn+zywIXLFlQOMAPQrMcPrW8C6Viw
VOK8tuRvB6cMmEg2NZtwsggwNp8quK35WH3i6OFRIH8zNgG2DA0KJDgfFDuO9pewAbnckfIwaYgV
CR8+64PTe2trCt7UQ8I4e7599a9wvpFv0AiYezzOjl/vTogoZMkO5kdUujjWttu/9JJXkarPrc33
UVY2ghtRW9L+Q3ewFIiZHQImsNFoqFIvP2tZgnDprDRJpyZAGlk9/mKx05uJ8c8U0KUgL4YdIANB
AfxET5DqxUwTAAwx4lqo9NBtdxMbJ958UD+ZP6rm/Zku7FQY6CfI7z/csNkhOBVTWcipemenEwrK
kj4t9vewpEfoBUVHHt6go4ptCf7TCGmLbFtVqewrpgl2g4o5NiG0C4gNijdBuUJnWK4EV/vc4ZYJ
iw8743Zp4X1riDY7oUKoY0YbihKYSM9NxmRQdXUFP58vB2ykM5ClprZQuIZR/WEqjB7nvobFa53+
QytcESvbzyo7rSBg+/fiz8+sItSUx9nUsUaVlhhjp3o7fzv1jhcPc2cV16ggFyoQdFNu8zIyB7PJ
7nnzDhF4Z9Z/qY7k/gu336QfOS1XA8W4853ozoW6lTwCRCPlF1Y6K2eGmIFAsgGT1XveGAtJNAkr
iilzd/2RLg/UyygnKFNlwtEfFBNaopFZ0aytcPU+60AnbYNdvj0oFkGVqlk2a3FWu5xXXvpwCwhR
TqTyFIFvgQ3V8CbAc3gtFrQ8O5b/HIDPdEXK89ChVf57OVtxATVxE6W+9ZTWyy1xeE92O8a1aZge
kh4Gg/exXSvb+UhnzNCcao2MHsFEpgsC55tU+EusR4nINukRivp0Aj6sSqftVMhTEUjSnziObYQC
sGFhsKcPdbopT0Ap7WKvbuE4b0DYLmVKxGfCMQeTi5G+kRk69BbOqr5+QwQw2AIo1oaDI2kAZUtg
3qbrYj3o22PbjIKJpPwPNY4h8rOuVO43QqqrctFmUNOOPVoSA02S/fpARebA1HHDZyKshHM2aVlU
Jzd1CBYfcRSM3OpqgE0p3JyZMONOJmSwjT5eF4eAJtP8o9+Gr5iITs399ov+IKj3jZ1ZdBb8CGXb
h4vg/yl28u9IOpXYPxO4sPcz6FwSLTZH/hsdBsqcSR9I1CnWHfdFoJRspDouCjHs6CwWI/fHf4uK
fM85lzQPLZpHHrfstyNsI/VqtO8Ood16SQfDTVvKbUiiDINiSzw9PgAL9CziVwFDrgdVQjKm7CxA
DFeNBx54pfYZ4f+6K789E1WTdFvNoRaVmuGf4/+iSoRBf1CAknkzLEAVG6GXkbNZeaCj57wsYhKe
QYuLF9HBaC9KUb2/U36W/qAtnNIibRz0z7gMefo31I15D0UNKmphN9bCVksd7gm2vcMsf/nuFJn/
p4p250TAqHP+PCp3kAKZr8IaKL55MD6WroxzkzhCJFYgKTealkF6tVaOECxw029bXcncEHV+R6fq
b3c+5TxaXdBBomiuCvdW+gt2is8QS6u26X9gIV21Zcu4Ngqlq9nzx6L3orx4dHFEFxBscP+ty26G
+lOglBjC4M8OludYS/4ryM4UvteH2uKv20FQcupWcgAJTS5ZMUs71rK8XLL8S2DetB1tQPtlmSMr
KwqM7D4D4yJE2WNoWLz7rOkE7arGUeXtE7ShtLPVX2CIjGDIIKXhSjJbt1t8/8YhUrEgT3PN7e+h
m/hXrmXxnf7nyOM+HxsaL9sxHKslNzb7Rbx1g7LUkODRVH6GRhk7/odQoNtd6YLBr1EvFAyF0Uqs
lGPiYj5Xq/M6T7LJx4dJUcOarhENrVuuyOqcgkH+0WbBFkBCAF3CndS16NcMRqd7Bep8XWMtQupD
8Qn7sASHGLZWCnSPcAr+6OGU6mMpMZReZd5jAgoXZQvE3ZWsUp3Y3MRoFbHvIToCMKn0Xo4nn/1Q
lt/6dWo/ux09IhYG8NagiCr2RlVKw8E6hfNvv/f3UBAwk9xZbv0gALPFmFxNypXe1+4k6UyzrHfN
bjspML+Y6ZF6Kq08BkCM+cYcGKjo7WIAaqEX3cHN1JZsUL4OixwK6x/Prfw5kiSwypkFUsZMkhL+
pEcD90WP5NFuFJOOLUYvZYz8NHS2k7qGtZgeQeRFy/Qg4F45w60uZNJjQUBqEBzTIv5n4/kEXKzY
8+Qd0kU9hEYnR8D7iYpNT0Mi8fpBvBNkJpAPUftd9PihF7VA2fEPcDNuT+CfpXH76qMf+XeRiHZS
f0DQg0AvGDhJvlpOhjiYulX7bg74VtfaVJjQwW2HNGjlJ3aAWR/sra/xlNUE4PpKGrmGpLtbI3r4
32TpHvb2YzRtFf1sjBxs5FuPJiYNprM9OI8ygVu8HJhw9vh/p++aKBjt8jDaA0ZuAJ2Mk3u3nFmF
p/I1ULZ+BTxAc6LpYTUr1C+ErvIp+j6Ju1kE7UrTp98Z5OaEUopSkmO5QaqBhcB1c3BaHwLaXfhB
0jZMvxaJHDowTy4IkhH08659U2vLIsvGshgo2Xf4dzQ8SAmhQ49IrXJbsSBkBv4UXBHeCOfUcpmJ
PgBAPih18C5aUaBhmE2AY3W0j6i/yGuYDA9g5ZemRUVJGXbRtMwTd5snfI8hStmUxDenkR86Up0v
rcKlcQ3omGylgDHW71POFR5rxrsbystXNkOiRsgbOJfSEd1+Vp/ALcTfecjMn/jtXKTogawsr+tH
B+lavRTtouoBtewBV5jB75zVGhngmdNaQYLQyRLWLjsykCR4a48DuFwhbx30T8aaO5Wlf5otPSBR
mxsEFlFfV8bmtMR7GUJqx5Y+g6kNoKPUfS8bbqvXng1lwc6LiaKSkJpohUT7ITVgdam7zKu3TafJ
mFjjWEbj1PNevm2ch0xlcmulDIxfZ/y0xMTvAkBlvWupvjpAXwRva70sNcy1BgULywIE/aeoaZvQ
DSEVK0SE7PTEqYcnxMcn1F31nfB+GmVWkNcIBjCftsbrzyeIwyhD7GZZtsx7gUvevWt/71QO1SAs
sisi7nfrDvvaf1Xn3f6cpffiYMFjUk+WIBXlnmmeCJdl+dWBBIEBevUUB9/cSnxfB2i9SLRfqtiT
EluzRBwt/79GEl6VlBZoQjTPZdbZcD8XAFdjD7CjlNM2KQORozALP+XV5DWxf96TbgyycRgIvWz9
RNoBEOn1g1jM/4XWp4dRN5wfS4KV8Kuv+h9eDFVfDjqHGxz44zGGtqEYSaaiF5D66xPwByzV8+XI
0yBWqzR/iYUQehbPcN8AaOFCb/8hQEFLEyOoAq9HQyss/mvAJ6KUL6a3NiQYCBnDqvNUY6A1cc9k
hEHjfsxrkNyub9fjW9PyD/DrWv/e3c0BenC/4I8jyEDKpF6esY/a3nI0pH9zJ30nLO+L2DHnQrov
SweP6JKcnv88eMlc0FZyW32UycB/c2qniaFWjuQ6V+PfEnMbGumSEDhfo0ZXsgtcVw898Rfyekvn
mgjY0hDT3m3Iph+xedly++EBlJr09V+TdEpYZDYwsLGZBzJzOrC7A+uOPIjJlicgroHXG30NiPpk
l6FiTLG4ulDBNkpEckZu4mUMDaExCpl1tq+PAXmXxXAk+fsuR/dU1LdY6hny5y+pXB2GeJ48U31j
5xHVSSp4vKjQYdTox9c8p7W7TPkdKfW+2OQAZJKgFJbXF6B28Ai4OkVZoQKxi5XV0rt+nIU8tos+
R1x/SRFqG/bf4oqanEKe79FtMBpjSaTOW8eKJMomnJRCdpmGWaJmSK2CjaYReoaU9YBDd1E2hKoF
WYyMlMydOrt+cAlmsHTAURBi23kcgBvaMnp6VKm3NGsd0g2GudAoDJKNipge5XlUlF6AyMuzpJCU
M2kq0hnO4oVkOdH1dAK4vKzn/KP+OuU0jCv1KyUBQfmxM9taxuUQo28v4ZoykOcTobEjyzRwhZBh
l9C6P/UNW3sABXH+RAP4Wp+ISeO0naLNWv9l7huVh2Ef7HjDD8LO/XsCV+IgLY5g58GICfxBTDDI
d1F+05IM7KYvbiuySYUS3eQc3fXrFVtD5ObM07ODrvOV6jxthHTirfi9d42FyUflttS/fiVYdkdy
Xl182WXnyuQ79jDifc5ONHs1T5PYZD2ZDUaUQEjJeBYH8iuFPPFN43NE1SGD6wIOW9I8yakwXJTB
XRWsXZ8W2lolQ2XfjSqStys6ky4Xo62K6tM60RPi4ybu8ChOI7Rx425wbtPVIY1dIN9s6k+QUwRz
grDYrpxTqBvx1feaYW1hISLUTdX3gxJSAtxVy2cyfNQxO47nqLxk97VCNSlfIBPIDH73gOyb/+2M
yyQcAeFxT4SYu9uM9gdzQJZWZ+dVKs8KYBGB3WXiSbJyc2M2hQ0mCPNZcUgvTvSzFziOGIo/LOxg
q24SZUdr8KyITTyZ+w4SQa09E2q9MmhQ9QLHDW0cqVZ/toJrdWyCDKMuA2f984vB8ohR1499Xzsq
ed7tSxj9c2Is9A6CED12IjB8/CbzcXrR4qYuAjwS3mt1HfX3kp3bbFLm4BBzb0SfQBW7W9yWy4Vh
PVzNyCZk9JFBHJgt/MCImd3ezjeivVxPrZd4QxUp8SkSseG5y+MWWJxylWMSh+rIAyb9PmtmfbzE
DK4Bfd/ctkluotC49nnbOiMGMljBqcKnO0clYq2qkABFYnQryMSlQW2BbjCaOepdAcbzdEfkAioT
gtMGLj6g5Qj5i3GLgXFahzAmzh8U0mfGtEawtObecxl+MrCchPiGORRvAJDr/cQAwM1hDOgdK4sF
JiEnCR/jswzhC9HsJK5xL10Ym4SohwyoHv1fqw8LzlOtfomCoPiqb5BhJcDh2pcMmzSFAQk1oL0Z
5JiSeBygiWHcxUtd0zUhCeT2vASEdbG4yUXGEbnT7IZbnwTghPaKR+sEj6yorbGz30lNUoRUoQgF
Txi9tJE5OBCqsFmKt4iSo8Go9tt2FKmMlLLz77QBORICZeglq63YizYj0j7ns7Qx1iv6OAvXSDH2
yoBAT9FckdBjV6siDdEHMYFQQryJQzc9Hcd704AES98wbs3YrpnKOlQcqOTmU0jToRSzIbl6RKhP
gEMKAO4/Gxn4cEz1/MJHQ86YAiP4uspfz5QvHFAZWNBm0f3iQ0RoK7cChj0/iTMgLytalbasy9BI
BEQFvmGhHMt1KC+Lj50Rgqp7O5XSX0jQwVRP5LRlX4a6VGoFMZH1RHKHdo1LYd49nV9W9VJ6Qxqd
Ov2gLyGWeRsB2pSZ2+p6wWj5BmbL7f60F3opXacirSztjzr42FhUc5ek6M7krmM1o0MW1iuFvyiv
pg+Y0FcaWyBX7V5Ad7yxVTdBxFAFhPGW7mgYNXsAykyEbpfDGVurcrUcKNhQ4/1/6h5mHgmCE/Nl
Qq6KSqINHc+itjYgvGfTwMd9wAYWUXouXKTLIQ4t+ymagbFB3/0jiglE7bfZrjVquFd/zgaIw2XO
ZFQlVjist3i4ldEDiMAhjW6o0lNiwLOuqIOCCcyW5K+d4iqo6jQp4F8EP9DBBZ//+rHFCrN6yqGP
VUNvS+0uNAx7hX0ForBszSxFKIXQdoWI12AFfkCiZbDIm7LIgUXVislk9NtusDHMITInDiH8QDKD
B63Pm7NoSfoDafFPMsMm0TFAq7VARcxOqNVdZ/Jx/McIgtsc6nJsx0jCqVpUJdSINlUhi47uHRXN
oQagiGHsvHemsP1LmA3ps+K52mDzyrnT8EJd9VqAfdtww4EfR4UOn9q9pOhsfv+ngRUI03pCyAGO
KqXlI3pLnQyF5HLTdTgUjoGh31ikIXzeGmzooEgqhI/ouSrCbVcngg0+F9c7XgM+pLxKA/dloF2v
4G8fqqH1Alm+/pvT/mOI5X5HTT2TkafQyVFxGIpFe/uR3fmJ6uSPDs3DevT98Xm6xomGhcsaLFdU
3j+FkYKxEUD5xXy2AADUu0Yfdg0dq9RJIdjEzxJua2AXHqmu3SUhLbwhr1RCkE7wbJrKC7uulhqz
5sN6CZDpzUafhvM2v1IGLhrGiEYsLPV9iqyfZQlXVllv7X7E/sVu9ZmljhSkH3Quqo45B2bCjd6q
j+ir1aICNRTjakvmqtmPw9Zs5wnhRAh9Kz4uIvJccldCqNUxEosZIdbduluykEYwF21TCcBWND8F
83wVvJfgQduscxI1RbM6p0MbnmRNvdCgvQjVNwQEZ0sugEnOvJpJqCxx9CoZuw43t1xTxJ7yhm6q
OC9Km0kN0TJPen6PfGWeKzCO0mqI2IKJjtCL8HH78Z0UbvN4fGO6l1gG4Z+2RjX46/PbSATSNE3x
2qlfOSQ3fFBPyNMNY0vKXv0RaxhXSC55ETwd5RuiLVHcXcChtTmsEQwhls64JJPpF0H/TLM3I9aP
5Ta2F30XoMR9+YwFOdo4fFTDdawxmS3mLLM+q1Ct/nLbAJkkUv3Xf3VkZzw3eF3L5Iu26C73oElc
AtfL+t5eHa5950SWxlwD7EBJrZdrqW7WLxx6djwL7DGGGBRHL1Qa79ifjq3RJot7oB6NTUzoy0Ns
uUm9+4PS6Tvl9rY12ssdieIEkA+74AEvgBB23Zdh+8SuiH0TX9d20UMayETg0xTemqEmX6GxHA/F
LC+88THkRLNZuCLWVT8+tiYKMX0KuVb/xKPUIHDvVshLTQM1BzksGBNG5N3KYBdw4vKBDbJeiwC5
+H789uooe504gHssy5DutcLaZc3IhSmziXUm08wE4BN2h5jCtMQ/Stk6mwWq76zlsoLcl+pwE5Gt
1GINBxQUh8BfIH/MuEbLbZwcF1sAStCQ6k9lsPgnOwgxtDkR+ivX+vZbUj4mom1NkXLSpFHzvARU
PZhSD9h/UpmF2b+PLUqT9ceOJX11Gar1y15LUifd+74m8I2DEVKfiB9QqZSPYPdlql+6GJW/o3H4
MA7glel9jlWedsMaBYyVvBzsGWb9mjCVwoUinGi5taKORV6mCZ2PZZMvEjk7A1hT9MPZyvhU/t/n
5fMCm8AX1McpltesLOHkM5VrZu7NwTODLnsmalfoXj5UR1WW4UOf2Z6m9u6KTchioAcoFRBovFU1
T+k7BWyeiPrhwbJWFOcQBWsshpSFxy5CvFjHzC1mSAyrIReaS7FhurUV9ffee06L1boeWEpb0akM
CSviqs/Vr/Rm801QjxcGLW0D+8Gi/WM6Ie0fZ9rMypyg90jRMG3q5L/8RAty2y3EWyQK9D2SCQ7h
eEu7gCvtDuXNQSk5sBodFCk+vy6/Szv15TH3ferhd4u7JExVF8h3lLxvzYQBI6nN0JpMYqHHgvLn
ugic5rDrDkWiT63lVvd5vowMXVfJRbDyhf2x/VEllrfJTly7aaVhHXIsrTccAuecqrBpqlU3bvaB
n08U9GEsRnjQh5eumn8Kg+5Nbv3fW3qgFSLA78GZdRm+RkpFSkaDvDNn2Sn56oTE10TBv7kUuK98
x1drM0WtWqnHEafZN0rbTbiKFqXU1m0TOJYdMqGu6PXA74s8+mkZWNkZOeiYkHEDE8tDhqdcqS+/
67lwYCl6Vf3AB2MpeXBxvWzuA9xqMVFpuP2lQf81nNAhhIMhasnbB0M8PWcXmUs9oUW0DKuqbBo3
pgtYLxLliB66PRG6p27vaQbGBqZojRdtCJCXtW7fZumge75jOhzwE6pJJ9cC7tamuCR2T2il9BI7
fPfX/W1v6bUURHka5fw+VqRQSOsQy5Cxoku0Ug6iBHnn7fmZSasBVc5q44z7KsI8bzhSmXgs/v2y
dstPav+nfgq0WqMjRa6PTJIfm42GKRS6XyYPW0zGAWFtQZXSaZYsFEeaUuo4ERcReAilFbeyQh0r
T1wO/qTgg14+EkAkxRFfw5O1czE3a3XMxMU0SlfCWJOHz4INWqD6K3C5h85r84Q0nSQTWOIyyaOB
fU+MGppyRy9K0nAoIAuWzG7YV3IKEdggiGqpJuoLox8ti/fpxT5Ws116pnmL4/h/T5iqBSid7Wva
7HXC8fzSsCaKlZds0ls9JkENjjlS7YuOyeJH0Sb38NN4qhNptjr0Iqaix6h0OXInCWbb9FhEg1bB
AGrnT2Jr5eBWnnBJFm2TZW1BzWpSj9xMKerWGn/YHaoXG0198n3c9WPlxcyzZpgiBRz2DInNBsC+
sQSEZeLb6aFgzcF91nSZW37n8qOioUP8cIPxhX2C4j8ZDgRpUhHTykcJj7CKrgre+Zx6zwPRGNHM
eydxjj6/m8Vh5hVt5lz+CdfzMAaqMQaw+pvdr2rBXfYoJyRtN0l7tqQ/sjgEUH66wnJ3JbffRhDs
jdAu/YKiJvrydqZPygHaO3oYWwyVTzjug70U4Vufnu5Sp0RMhsksPBfoKcOytjmZKC3zsasS/hMe
CHCvC2ucbACqIHfx0xN2WuPpIsEA+EZpKLzJTzIIjNGNGLZrsCLhMvyYsdcnWTa61peJ2UwFHTB2
bsj+gZ0TaeDdV0q2bYsyuZsBx3cqXKz+9LFpiqR0tZIBWfLvWKwFiLdrLkHuyXCW8siX/V1DqPpX
wio3l+ne5PfED1OPTBwQT7AMUMV+8JFIqOdgV9eJelmWsWHt9R+Ug/skwtbW30YjXfsYbhCuKywd
IOFsW2T+ye+8fNVIFa0AMc8Uq7s8Kd0Sx5isnRdnzPtZv0pWjUbdGhrY6UaBZqjAJiR3gSbL68s7
fEdUAqZkVXUBShvzGMyN90L3UcuacFBi83P7tk1zv4lJCNkzOhp5PuHsuAaXKo84h/QKColJLX/R
PMpeeSZ1eyvdsyPxlh4oGoHYuhAkg8kUWZ2Kxd9PNRTapeXwdAuawHFd9PhgqjlTcb1hjPGcBAqU
EOLscBN8FxDrWXO9HxnLWc71pL+iEMXDSI639A94xZKznmlby9R1HIkUcvgDurjv/BB/WwWNLHm/
s5d19ZeO46di7CjJEXyaGUq+c0t0dvowSTRWEkjK9hzZf3JuVj/QW8uacoYwUeybJVuLmrWq5bPY
BassyxKOk0Rrw9VEuFO6M4hHp9ybYyo/Dw8DXWWTHbgp91zrhpfmIqZhM4lklPScOOLlS68QGLjo
U6UaR3PCRV2bHtO/pKdJfNlW3IxmxrWD4VJmOMnW9m7HlIDBRMnZsyV4/5vtWOx+9qlwmJ/FXODb
Pla/HUAYIoj72ZWKYaUw6FnpBCl7QwLVLE89eiWzQ4WblzCFN2NqUNRPdooCAGsWouUgT1XaScxf
WiL3ukpTiy7kntwQmL5lNs+nzijcUj+bjh3q4kwLJTB1+i4Xsvk8qSUtVJB9ICRgBfm4AGKW98PS
Vg2UmRzeJ2ac0TSm9fVxBDyt+MGtPVUs7RYjUo6w/RmN34mvFMNlHG1f7jPPQY1XjEb7ZM9H8yCp
zz+o2fV9F6AI5oLduAX5S2awBzXb1kRkqTn0MwakBcevqDs1mubOpX82PV9wibRpdgnKfk2Nzcw5
WgU7PZsW8CQzz9QQ3RFInv1uVPOZUW9IiSMVTb+8umKes5MnPqNvdEVfQ42moZN1mS2P3eO9LGO/
Y4BBs1Y5W/cqeIaFzfBha2EvM4VNZjrLa+1q/fZzTz8o3W+0BDJzWj8GrNUcdr2wxJ66h7OQlcLA
cTGPznujEzAQNHnoTotZRdfRtucSREAOiHfrWam4MnuZcOiDlszVgiWOKZAJAWXeBtq8FUmeJe4a
q+9piuvvcwij08VwDQWh6DAAq9mUN+P0ZLJhPqZNTNE01lNf1fYi4Noxvkq6rhZEO6/Rsmk9dkv+
PrVIvZ7E9eZ4st6rGDPA7qY/02Vrh2BRrMaCWS+wIuK4Ay0wYWJGkiixv4IPr7Oz/S4nCSMYK2v7
WxFFGO8E1rpbtOY28JI+9dsJTiqUIcwOn+sQsaDIYAUkPD0jBMJeusN9fhIO/NoA1H14iDIvr3mW
5YsOkd5XOL4DOoV3orOwJ8RkpA0nhRMgJIMaI56317UMin5/3b4j5uuuXlzMEsDJhQlcouGEMGXm
98jXOna6w3KDtjAIWD+z+AZ5eK8tP5QobQA1q5Jd2MZRfVrxXtXNg8mlKWVTKGOxAQmzt65NK2B8
kyz6wmOxB8fTgmLycw5WEnwV7pZk8NTjqFjbbTtCfp/vzGu0pFzj0hKQgVSMmcRgOD7EC7wJPbvP
5XXWQXfbksWyvZeiGxzj3sOL3ghY54AejeLUZstg1zFF1zsZ2AvUMuzQWmAr/LjwrQXU23u/WkfO
Ac8k9t2dwH/HkmvUfPrcyQh/vU08St/Gb5adaF/pnwQvoxmcjmHoMjJzdXUqX/quJ7q1g9fZ1uYk
4fZ7+voXFT0OrlVA0ju33+E/CfH2sbqIf6P098dWcGba8nhRFkUqri9LqLuE0q2BkqHMKpQy4tMX
Ta+nmBvGZO7/JathV5qf57tmLJ86odgO0cnUoVVHpt876ZE2zS0yU6ugY4v5rgp1KDoY8UUOB8uj
19rF5eCfAoLuxCbIDldhXY4gBKmu9a5M7siH2/0J1OJ7ztxGYd9y/AgEBGtOuCZrr9njw4L81913
Pqp+TuOJKkvDRFVQN38XMozgA7t2PM6bjlJU6DGtekw9gLdqsnWnLqOeGMEDFglCAE5jrMtE0p62
zPZ4R7zhPe/cbi1S8zC73TCitWmUXvC4TbUvocOfkfiXtfESPfzxE6iAZlGCJx960wszZ5EMfIuu
A2QeNmIUYFK3cKtSTcdEG7h7GisDRTbmv4U/08GWTwUBVgNj3+uwXReS+XclgKociqkMOFS39C3d
5yDvpCX8YjcDXumq0zPEodItyo/S4+MeWIIyCtOBKHbOCFJZcpFHmZKu8B6kUuzutdoZynRkk7P/
8JhbIpsHJSV2SWjBGLzMBBsoB9EZenIXm1O2v9KVQM013tUv/F5l2rmSMzJaBH/WMlWDdlo8n310
Tl3krILHLiGnKlffEdORVZAOe82RbqwKsvAHv2l9frwE949vGdzfNcqxvxujSbbjn8H6GrO5VxrX
c258KDDp2txdp9nTcMi9K3eeomlR4gIrIiegTVhLGy1blAYBuWJ7X+RUsrH4aKYygL6yuCJaUTgD
lJeGsIH+3kMN2/eHjfWfmLmTwYPCeYzgjjGuxtPnNcFRT0h09CuXpWKdj7vnN5cJv2d9X1aXNtDn
2O4H6jv3RnTs0Hc1SGBohyiJhrut5PkTZOihottP8i0bK+80OYNWpVxS+gLcLRnkvejoNx/fVGZ/
VYyrzED4ai4bkzbdZoSCMJ4VoZhvb8G5ZF1qO/pxL1TpCKZ/mf21U18HCmMlM8ZM0NdgZr24gOYY
j1w6Q8uhww9nv6+AgjaBskIBOFZ0HSxNqdXCcWoD2HPc7n4KVbC1ZLKr8jHL4iUXFRU7Fctn91I1
G/k1Nzu9US6AvnGwPA6qaGxryFslmPWprfQtEWz1JWe5qsrJvfzF5C9sudm+jMTSntrreCAyn3O0
bN4XdmYpUUUpWhVRRR6E4NimKYGbdy9fxBoSAKqloZhMK6h4yo6350tRGWSOR8WEvJzfOZ9Rxtou
1iU1GBj5MzbviN9OjK2fKQ+JVs4nQZ5zy2GcOfBZQC+mkS/0PBuNFyIumpjZdf2DJeLXQ66r8dD1
zBakTXi3Ar7hTJz45ZTvH8np50ExDPnIru1ooCtbRv8PRQ/W1G2n/fNECC+rffVvFEHgiVliXZjt
G7Ght6XqOT+lxHYcBMK18xM+blncd5Uk0W+rmYSRL+kgbekMyk9KMcg66JvsWNJoalbEq0TCfT/7
t980CEE729YoQKa5Gq6ONag3zcO2TBa18UNS37XfbVIThkfZ9zQ4JdJSMlKsP8pY1ZoYlYbWlTXQ
cFj6SQLMwdbCzVo0kHfJTufUSdIvDtpqKY/j0XA2r9VDdi0FVL7rZw1FetXrkAmnC0UE3uw7gvE6
jNhQe/zxIO6YNF7Zi0OwUqukEgjVNvAKHgPX2c8AbtW/Y1/PCIPJuW0adAdslbU2aRlZx0NDnljq
ee+XvbixYgtwdJqJ3+XwKg8dE8T8IoPRl095plSexlGVdSUsULLwMeCdnAjY8lTktclGvtdCt+oU
Zow/N2TpPVIWcZ9qScjDgPU27pVaUJrXRUJqYFFpj7C/5we41s9UD18RrRWnzs58AfztVS0UEU0X
ie95/5paJTuVzHvFjNkx6AaJaNTev1miBLjFySIgIue/g5j9sOflaaiRYcIbh8dwV0P3T+9qVO8v
UuJ1FXFQQ7AuiCTbBTwSQ4+pUNwXEsScI42mJmNzkqO/s4iOvKm0GU3hjJibYaHFqeNfewRT37FV
pytiUcIJ5i9baDY7pTWcjqKnvp8OqqdaXjyaNv/YXvzcMtRkLw5WQ5zprQOauXlzYWugShWJuVMB
McHSFOoXHTiyvAhY9xjAbHhPdNhxHsnJQ5iNgKTcHnD1nz469Dlv1DIRxUMzcOmGJNk4WqUfbmhu
Io0uCCqjXB1ijhsW2BX25M0cVtw+hO9DTpCMSIGlI5pF4PtxAdZWnf2AA53L90U1cQ14/O7rpp35
e4QFzdjx/b77s0bxhHvpkAGUyePCq9i3N02mDu06Kzk0RFDjnTHew9rd6i+4h8MDSBHUiwegTabw
Xj+yfhXCh2h2IPBqbycvmCZg7MJ05ipkZdqPhlTI10SLIAVjdOmqBXyGTehap859VoBIyGJ8BJIp
qr+4/KVdSp29Y1B7Og2t0doMLObOSBA+EDoRIT014oQgcfiGhkWv1uD8R3EIxMXdk7DWBPIu67Gs
6Zh5gQ2WBr6cp82K+khnMku9jAHwVpIodIb9gJe7+jZyPfUMTdp3CzihcW7NeRzeXWST2BTkv9iV
79iYiach/Y54VllLjsmhBnIeSPyTaLiiS6jPxLFOJr4nHUZlp132lv16wS9HFiugafPaTq5ZhYeh
sXKZcMNiXcl728BxvGgPUwYWj9FpjMg5Qn4y6K+bpz43/9/eu+SjYC9x7AJVgQpLkFfktyVKLm6V
j73kIi0wmQwqO6VFDonHVVtTwP3Pir9OS41lkBmV1z9Yt2sEGuNGS+dsgdsjRzCRIKh3ChyBxFDe
2pgCJ13pjOt+AkhayUpdiafKcTq/ysGdZyLxfBrGsdMGeMA97gnJTOID++IqgjJH3luHijAVS2Fc
GUCcMvayHO22TnFbEi/qmdj8g+FVkOtCXMdL9H28fRwWW7REO4mIrFkdFhetDBK4MXaf6hAGm1i4
H0diQWS5xrAnWnd6/JaWhBNP4MZf1f6QNjsZa8PPLoLl203jU7sxBLjT1ekg/msCqmZalbo+Q0Ev
GD5ltWeptzXetju2qLCG3nUPn7vudh07195vMh0jvJOns3wNlNmhxZngh+lgxQr+jzyD0j04w+U8
VQyEafhmGQaoquR0OJrpe+kfoxH0F35BsKzbEAy/NCGP/vYpJXx5YV3wmGa7CLLMh+6nj/VD79XD
2QjFHyJYqti9BwXEhMT7wp5y+6EYw+5Iqli+ih8kux2OaypuNyibpr1trVKfwJCQ5wpAwlhzgrYe
dm2E8XjyMAG13HvEDVHpfGxuCkNaawya54I+jIqHmksiVfXPZkLBa2vM+WYqZx6DbU4JV+kb8ptf
dcUu24VwM0J/yyRO8cUzfl7psjf7BPYUr1P6Ad2P7kxa4lkyGkoPHlzMG6UzENshjoQrgYRLs63J
22eUvOi9jaTk3PzQcrgxH2VjDeSbxDLbjQVjjg+3lFPahednH8zRgeIyFPKfZ+z9k0v8R9kTNieT
e3cTLruSq05NXg3CvvvWKe/VUI7nnl3D0nsjuh9YVF2fbMuCGqMw/Zd8UxweDgbymZzf0UgAvusW
os3yeW9BTAUTF0TgWCPNBOnrzRSvx63j4wifqn5WSfBKflCOSQUfdr56kvuSjNjUsn8mYQ04yx3H
JNeoYXPK9bAygLy/gv2/AT+7MpfoD+7tLN8xX1Psm1iUV8R3ULVtXSKyb+kCnuI++R8zKiWmnWsz
MmwcDghHioyPBPLeSZve9FJ2IR/2fRv6Wy6ViHx1zG6pGx5afOVhm/5y6xRkhRxjLNsLi8TUe53j
euCrSVOU/WnYBqJ8yQwIdCy0BlB+O7JwNSn1UMCOzO7+pI5xZlmEaIgLBN+HtZbINHCVozZlZnvS
UZ5oEpMRYPev7NsPNzxjs+wvSOsyXTPFOdr1prHufeLPG5SYzWr0ajl8/lfGvzW7Wa3xyBw4dgEs
gekrMSjqmUhFV3YVCOQXr5gaMDA5oxfAlQkfBYjnBH1K65HrK+1dHY6ZhpSaT7YiTiwyuceU8/CB
o+7WcNC5QhyWKb5TcugeWxRMzaY+L8M5P2X3nT6oMVpLKDJ/y/AczUgmdjy7euHfG67pJffgrFaI
Wqhu4L950bXjf4uyFY205TYCPlr2byrKDLlf4DZxQsOZ2x37Lt9BAUnUgFEqTJN1pH/8eyNpju5G
AuuOoZ+wr7ePLAx/NGzrqixaqR1aJlj7r1x3iCFAhWlI5nrpEOxKTx2S9cq8k0MrPMMYW2OWCHfg
OzlmtHFG2pGJ6cghy1Qi3mhzDEI5G0PpieIcGAQzcaA5i7T+beCkKpny+Fk3zTY5mRGbMsCjlDqa
l2oM3h7up1E2KdUNb2aoATLhsGVc8KfhLV0oWrZiYH/QRzPWJKPAxVksILqBfpPpJEAEZvvEUcHT
ol0fOKGFJFuwuhXd4J9Rk5gb9zqMH5wtw83+EfFyia4GlaImcyARquBdjOCO14GVHi62GsDCSwWw
rHEmU03ToYLSW7flPgG4JpMavSrneb/4MwhdwD97PuLiGOND9m0TE+sq1NfGE9LU1Wld95aK6YfH
uqP8rWfxD5MTiXHjW/cZmXrHLXni7SGaPpzPJXinPAvCrJ5Z5DfTUvwGiNNrNtOb8Qonyv6ZYwfR
aDKaDY3js5vZa4QYb5CHy7p5Z7xDg0OAPH6eFooabkdHhenIPw1+R+HgMHxCL3xu/+KcevEJDZ+Q
Mn2ZpGjCTNQB7npSMJg6HlOhbquhl6wZqCpYLJ3F5tXggQ0rQM18V4nbjaoLM6bBBKalEJskmdIj
I8kbI74Rm1rr+6dEHKdhSxLZduXfGTrbYk0KbrYtKmCRzx+yuGmrgEz2rF2igCWMqNzKheZnwI4K
LR25JHWS/jxfDMK+CodkzKLeWFIodE+rRUlImads1Pcp/pDrdG6/3dlXk4G1sq9wpSVHj5EEFil5
MF2t4v/qKxs2Roy1Qu3rxdmWDeb728jrgtyU74+c5EAe7ezAOfxbjefs2sNndX2dqkyMdObnCDRv
IAxphv0oBO3YS6b+RUDf92xW63qoHq4naN+05NpZUL/kLHO9eXrcRuMIzEvahwVApic6dP/kDyA0
7h/NKtulxNMwODuOmlR7ze2L2sbbcOXurSYym1aDmZ7kfdthXagwtkNkDtnpeS0z+DnCmSf/aa09
jESbyIAHLgh5CjDuMc9AnzIXvv4EiYtvO2yeh2XNPOxuy6pIjwRB5dUQk9fKy3lKdElLUKR1hWh6
ZIpL+nhUa91RAWkwrbR6COu7iEFF9m6gjHOfAn7TcE9tBye0YzZR52esRg03crNt3mmA7y086uPX
nU2Nb8b7tfCuJ2P7vOn7YAZBbqScePxfxvBWg5eVUzGNmgkNPj/CORvmWAZveW5ubXp4fNAERT1n
6regB2iOTNnK7IA9NZl5KtXCfUq3QVfoILrFbGSEs722mT9T9UPT/FyF1+y4hsAbCz4PlGdUyAD3
H7deTnZ78wTbJdWIk8ztqQZ9IzojRtNZxsNE8JEJWUsrkGHv9Obo3ptiNb9zEBMoz/JRlHBgsqdl
ctKRHbY3y1nTEm4K85WQXOunuhguFgSVbyQkNoJg9/fW/HeIHCSeAKG3sruujefFf1l+5pZ9v/S8
apcmyJof2y2cKYUP3PW3WYYGwuZCWkrob14WFQRsV9n5pE/BlwOJQW7MkPU+InzIirfXKf4wlRmL
wMH+rpMcT1tBCvvuNRwzd91nt77c+2WW3MttLbcm72I4kMUKLxTFen/QO6cHvhuXbZ/gsvZMlpQb
ST25C2iUyz+u2DW4vdu4HW/SPXYle1NCIqHzHYWM0TZ2ceiCSKjVzFjRjNUTJqtt7kIcaQLwx1gf
BOjldMFUFNf5sF+aT9pZ/sxugB23DG5M53Nm9uNJsjNh79fODgtu6Bixgp3nt9iV8Zgcj5VFZojz
/15bNcz86JlpbaKcY6O95FIzj/YiZCf+IednWIjQFScz2aRFeDW9gfFnhdr7wTWJtTe8QwAMyd+l
WEN6/LEaDZprsVY6J/LWVgrOu9IBvkbRKOutpLsIKXhTGqm5bdabVwRZPrlMugRTHQuCMIv+7MIq
hwVVPy+26PajVfZ200Ze7vtybkEFAFIZY26iMpZ5AzFvg3lE11N3m7QTLZPwR47RBDAAnP9wazDk
ImPYuybtbG9WUVeHe8or1PnxhcbBR5eAAvsLsGT8c1YTA5g4krRVPWAQvtiaJHAZL34u458o9upY
CdeKHFIPUiWjW09etlRWGoK6P/grlmeKm8B80xl34hX/ZWHo0b63QiWCw4mevLLawujX8rwzZ5Wc
5HE8/Td/r1GK25MXMCZiUuxSquDlBnCwZt5LdFi1g37hQRY8K0RMDaLEa960u94J7QwbvDE9gclh
+iLCrtG9aK8jkipwJeJOrycuzn01fNb0FEffVupYgGzUZ3jKj/LTOq9ajGOFtIRSJukwtOMUTFsZ
awO/iA2ZJeN/iyER84MAC7TDqYce9oy9mXY5MJCC5G5NprlMptta8AqWPFjwqKvfSu80/kxbBPNn
iZ+0qrPs3xBkOXGJut3QmHRd0DpGcTKBNxWZR4PxSsEILjh7ip1/fd7wYq+dWrcjAiOsPHWl0wzA
Z4iZ4Wn74edfTAGNe+xoIJ9jFRBFkjZSm0ELYKBhYAUxXaMgrd81pauhiKlE5KsBB79VFK2xPeNJ
sBk14JslUm8s4c0RHitzTNAj6QWeGbrpRGWq4DcLcO3Lkdwl+12uzqMMYAPNDPnpxqgeFhNB1Wkc
4qOZIEbO+1lkzSaAinDOtLWawrXicyemJF9OWsP44hGEuwRLNPlrf5nFQ0l/bJTjqP56b1H3eZjX
PCuFK7eKDXEv6n/gyg9xbjEGrQ4ecYLA5w/kTkhyOkeOjrNfTvbuY8FhUcBym1bab3dw6jlcb/ob
r9b8QNAvT/sslla+778IQkPo/Vww/n1JcflO0N2gUTHYLBTMHTr5aQ+XvdcIVXpGeZYRldb2UtFp
TWx9pvOJW8Mz3A8WUFJt8/hrXEziN9dJmzFo9BUg4AWWqZ68OuQ1kaxsKPjGu8aQY8Ps4mg9cm7z
97A1/C96GQDSDlwkt0NI4PIwG9AE/VuId4Stfcr7G0Wijr88nSfN1DMffX7J/tSVfxKI9T3PSenk
R8Y2c3yGQIbcGjD8gON4pEaZzmvKjEANw4RyIYOGdFpAIfRjDLuShmXAtRU366EfObH2xsPQrOGk
Ed7TgSfvZp0KcdJSrg3RRhJ28LGbmNvb5fB2dZglH3sC6jxdY412gMt9imj4EkNFXYMjVYJ3Grtk
c+P3cIbbtWMtwptPqu+rZpgLKJK1npHMkrkFN85BGXFRerywGo+ukt9UEgAnZm0IewGLfOTPsNyt
0Lq1qhNUNOcvtcVcB9QeJJo61xgPROp3uYFiSdfSS8FlDokhQVoSCQj/HZyuMsYUaWokLE/TvweB
G2pvbalccwoSEuEI+XdL4elYEg8goUK9rpTEKTSm2SkSlTJVmxJXpgDgA9VX5baNd8CV057ZBVSe
weq0MC17GtIqapBE274CmBig7qbCGGHnz8yZNXi+ustfuZdczRGibPll6iqwWQ9mqIzuEuac8hYB
o5FSXMMpOQKUjJR43ZBsHk5EBHLtksKuIT/cfJbcnMXlHx/csEZ5rQbDK8maJ2BMLdt78Xm9wxid
aSn2myFXqg+Xho/Eg2f9fgd9bjv3tLbTMrc+56T7dzj6dVaepZw76Nt2xB0lLh9SfsJCFrbnSjAt
kJyEQa3k768QPSvJ4IBlt6is7IPRTS70tV4KNiysfShpzVXM7W9vFuFUjkrPvmk621DxT1Dr0mq6
GdGjxl4lDZNudIqSMNGd7p2K1MwKS5uzaEt2QVBCyvjb0x6Qv2eojMSTh+P0RZbKYsXsICx5LVI+
2DxjsPJ1vxSiexCC4Kqt/GB5Akv5K1Owy7po1dGab+1kZMUs66c5ejHmdPXPuqhGbgw6kodC/T1R
C/meexQVMHazITO2oyBcltP9gHJODxtdDsWTS1P9Iui8uzychjKgcfJgyJGf2HpQkcbtDo456fbM
5Z3zrxM4KEUBeMibv+eVKg1tDg6ClWI0E4aSaerZltK59mpkKe87D++/QbbBWDNzK1RqMqzwYmUy
b6M0qUfO1/7EUhd5CePfFWIEkN4pL/pwfDf9TuMiaCklutkvIwLj/ZK9A1bPRfaJUFB+ctigHE12
11tiZll1ntdHfi6Scu6Ldj2qmU4/73/N3maGWxu/6ulRt7tpX4hsxyDXWV6bNfq/VX9iSYFex0Qu
JpkZk+YQ4bY5lP73ZZS9U7mzV/7ZmbQycQEHzNys99ceAyGYG2drQftQnIcYmK2G1Jg75gTl7PLN
93Ba3oqF4SnEgMtG38sb+Rg5Bh72mBZx1J2At7dIvNNw4NKXG50LpIO4DTLa+GLuOXobybKCt4FH
x9nGe7zcvP1shmw+FifBBUySIgWbO5H/D6wKQEkT3VtT4m+v5Va01zqrEPgYKCWJpJLjZnAwXF0A
VyA8NuMZtjflyDzyjPN+6bhN0wUYVPvEj90MicGt7XXTcLw6aDt3TNrGSuYw4V2Uesfm+HSmtopC
PWgiWD1tcfQZfEg2577xtv2kxieZo7h1aWYRhC1uOStjcm3ftv5wEBhjnGijbPE9RDAsSt41F9+3
6D3eJLs5E6q2UW/g8CzL8kDJ8x3Dv6ft6vM69SX4/P63ngKBi55r6szJQBMNTI92BOx3NfAlOfYB
zdrdiT3U5c/BfDijbOSjr1n2kKbS23BmmVF9sYLU/q0vpbISKMBcXTLxEnRs1upuxxyTHX9Sw3qB
xKXrNLL1GHMyGGgfvEMbg/+sAX3Vtcjsxa+TY0pv2nczYpAJo1ajZ0WYC2p8wrkdxq6eq740q6DC
X1gPlclZHyz3MNJXWAqkMVs8qMXS/p/bEeVo3LjwL6SrQJloSy8kt0Km5ulSLZRuDCy8c+m4h44o
xrekkBWC8CuEd8U8ZY7BaWziEWQyQnNgBaGb7NSyr2XFMU5PBcWKFazy9XpXzNmoeq6Gtc9D1vKA
yLQjKII95FkJMEPQ7iJO50NC+Iz8ZXmfa497VESmIb1auH4bdaR8mtpeLPJr8A3JiTmuXIFTu4ep
Jft0lP02D8i+thRKW6TUVLFXDm98GK7Z3IQxBFjpEHOkeJU9WTIC44BZcOlvNCSnr0ok5lH7aVMd
NEMP/jIDc/cvcBauieoPrLZckL7B2YNKTkVjYEgzjmpdr5zvD090acdrOSDiora30yJDVyck39bi
evX4FeaU8uzVyxvxDB8EY4al68JTuqGg5E2aiy5OPWCf7+exw4n7DPToVArf19RsqcEBykJIgAXD
dWeR5Xbb/CjCSNpnOeNbTK3Ut3QEBWn/f+duYIBiR+sql7KZfW/ZwdabQMeE+Y6fJ2Mj0kzKv4nn
baafIrFZR3EX3T+NXGQ8zSdAf5IDd2Tayd9qlcHAdmTLfQP1teng2Ehy7JVWdDeoDQpM5+t1yqde
WJ3NyIWSmvT179tPyszJ3T6g67hSB0jZdfn12j2yyb8/RyIjoiiqeFGrC38ktHKfjwhcprxq67y6
Y/R2QLLQvU0PnPf5+WIw6JGQkHi7nUDjAC1wvd1cPYWcnrqGQ8Nmma3IjDvC14FH211SGlgXbFXy
mMMlW+dCuWLzE8jdRHHKVG11CPqg6B7apaMlf7M7hb2MoZTJGLhoQe3C4ULzsq5SC9qjVcCEe6Ka
8UdPowiZ+XnodkfzCPpP1PR7pj7hgmGdwSywTc84C/yzo4SAolUL9hc/5FLLV7ubKdqZPFEKzurO
QtpG0i81KmaWrA7bRVR9Ph7dOpdhaOeObZ/NGBuh+r2wM6yqdqpCs6Kd50nlIxaDUaYJbZ8Mig7g
jgDeLP5glVaOfZqnDx//ADA+HSRlHUpmLgcVD+cAQyRlz3io1AYTM0wqdGKSs7BCpLqOH1X85jJN
19f9h8+LQmAp3V3UGvQpuMkt+1PR2SGqG4fj2QwALXnr8K81dCi8EB6Ld3wpWHCl0XzW8yw4mkzD
3LQ9Rdp/Ywm+S8zSsND4AAIRHhzqtZ6kvOLuo0SO6/N2d8vYCcG3QsCgASbmVwVuDBBzHNFrdY80
zDPGwFKOdBnFEa7kqNgJvq76F19LC224gncngiR0K3Yq1uxLezdS7jbJFMwWzwFdI7mVoP85sWNE
vvLYUy8iu+86qY9h1k86tMiA/tMQacVbxBAl3gB4ErzGIJDkRKHP0QIADlBhBCSSCrhiUoYtmx5v
p3s0VCEa927cQlcMNX5qBm8CC+46g6oBSND0JWutXRJfVxZ9Ll5Dtj9yAwBK45DO2l4oQdkf/mES
hLbO+/kBhbG/xKXfdKOCsoM1GG+2HM4f+vuVDFTIUU+3YN66oia6tuoWWoJUqilv7Gub9mTaznv2
n5CRhixoVzqgDbOVa0IleDkX7wdkmWumAlMZS2B3rNGTmXe8g2mZkTc/lHnOtnNhr4g9pMKvXsW2
fGVSs8xagXWlArK27R1cK9Esu5UJg8g/ZHG08E6hlYfwURnbrYhQTF2j0/M0wpe+smyhM3NexCMl
kPrNwBdqa1Ndm6uLR9kVNkGMzsBLL/odfNd933PcyrUzvJ+1JP4YAjXrcH4QOEubbcZC03xyGhpA
TPi4AHKiRSX332YWtq/izJgptfSdLjK/isXEXl7KzWIF2hhl9bAd9aNIZRemhxO8F9KxI18c45Aa
SGPVPOHFHt3/kMGHLxBdXtFXHHHeDSq0n5fmspy2T6srQZmfAtDbSE4gyQkf/Rqll57NH+dBO669
OXQOZ2cXuh4Brt5RF5L7ITCSUFTCzwo2zqqIbOAqtEQ2r9PI8nYfQAOjo5cMPPZxyi9ypWh9IIFl
YrnDO0DaimENCtG3kRWuI0ulkR+fYCoaC5EEHG/mkJlyvCO8lr9iqWjiiLbMsYK4khR8fKB+7HO4
N1O4uBisAyUWrWzlg7dVhBSJmyR3T3BvO8fDv0wRH9CYKZvjLPW4mDI8DGsLNpFt4uzJULi69qTg
OH834PnfpR3WkizYuNYOePE7wanE2VMZv+upzQmqbETwDc+V5XgHZEiYG4usMaiudlaRdikZ3iV9
ydPMmPma/kH0HSrh3dIkN+hRBTYFJa3GbT21hc474ks+ZUY0bnJs9x4RYiLuNv0Y7pThrblDFU6R
zFnj9ZfdSuV0eRV6+cjieSa9iRuosAD4n1vhGEVhdlWkp2Mi+R9TWeQr7Fr9JXq5B2Mv1Obu7+WK
W9mLgJi7Q/dsWCadgjVp4LjCxX1rNdh7vmXPEOWVC+oj9uJJu8ISOmcybP0UY6PsoptkamvFW8JJ
1BGjNA6QIPOwmQc+Wlr3n1/f9MFXg3SkFCkBRRXpz/yQWr+gnSaXmeLDiUbEsH0jGbEkER5OieNA
D3hLlo5lQ83pIQlrGoSOgIPKDAubhupoVutbpVjJs5hBrXoD0mM/Sguaib9vLCFMR1iSCyCDhVN4
nkr3VGtuhqfsCUbWi1W7vhw1crsb2LwPxFJYT75aiW2bDiayK5p3jLxQCZcd2G6dsijjW1eWxJLo
zPxDEOaJtKHQzoDAQrUYllgoF6NF8uZ2e703fa3ZXvYf4wLizjB7lTqZJPy5psBhueGjhGZQlr8e
Ltsgw5nxyiO1D5ysnSQ7YhDFtFagFpbSXPYKNklZev19WWWWf/UqxS4wCz7IvKg6j2q9uUkztYTz
UQ+m4TSpuk8xDecGlCvvxwzL37zJkaDkixGOwVJzlEqIa2avs50yBPnmG6JfZzONNDlJSMyU6UuL
qbPXb9kgprQP/dZa1sVCDkNfxEgm4AnM1T1/gCDtmCzQYG+pEezLN0LS3AX+QvN6rNm8o/Y0D940
lzJbHYa46qf+LvW7zjQRp95a84YU4Nxxqo1o62+p4Gc4iA9Shkd9hMp5l8H1/8YQ+H9BgVYK8uJ8
HCWmXlkHtt6DQLsq9AoNqHqrtZH8h8enXzynb4HoLCKXXCULAsm7lr79+34Vc+s/EvtjF/I5Qssh
8QlyH4Rdo9Xv+LCa4MxSs7j306ka3AwDs9cFCYbExIXi2z7dJI4x/+eW6GM9zehMQxerVxCvUEea
AfEyKvC/VqR/F9wlJ2b4mXsM3n2UYwYX6F+clNiNScNtfLfaNq8qiNKNV+rN9XO4fae9274vOmG0
90b9U/iAAaQXXInNb5KPVaHoGe0XO+sOMNNEqCiH4pDU/dp5T91xx5MACXEUxQoA70kboGUIcGGd
Wc2ul7ndK8lowZFFlB01XV+jv8mL4V3DKs4dGywFCbsNaXHHHp/NFcdgy09MYbi89kUNo3Znkrgd
uelJuG/7KeB0fCc5PSB27JxRW41DUibmIuFXeW+1six+j+EtNeZ6pcJFjFWs3CPPnN4MWzroeKIr
29kpYfBrnOQBvRBoq0fmK6qBUwcj9m0mlPsxZMLVrqNeSRauQ/2jxfZFVBmXRu7PCuULdYAOFBjJ
E8WGJccMVuBo20+kGVDyDFguLZPw9yCy62C0HgWTj2psDv25XjZWaKr5hhkvkCS2np3GLM1gC/Hg
xpLqo93QsIuV5YJtnrMVeMd/XjpE13o0zRYvMM67Rc0+KVsdSZHXnZqp3FkKLlBUadzyBLKsCEKG
tGRGd7ona6fqcPz7Hp5G57GKs4AfhXAsy035ZO1M3Zf9Gep2ynUUDJYEaBUYRjaHNxZHCBBcfytS
De+Qc90dNCek5my7mVzmFW5hWDO/fil06TkUQM51ZBK00dTMYXTeIopl55T+n5q6bHJAmUsiKC58
FXyNwOX4SnecE+JJ+M0F7ofB7RP+Dl+sNDsyJkI2FNIGaPR7d2fglvfg5l1Lj3hpQJVew8lvbTNw
GtQWPC7tFP7sVBGAZ+5BTbxXOkLA0qrMRPVU/92KPBSxnYfwL1fhyxrLDzQPdPcBYg9OzrjVAgeL
zG7LpatirYb07jrmUbwSpy1rhKTqAtURX0M7UuMyQaCd4eX0GiDJJWwvgpMgFUed8Kd+nEYM7MLj
1TifAoNFiEGHt9xXrvZvpzhUrXi7yirevJntzTIgS7Zmq2ljQc8lqpqYYEo7v/qGZcLCzHmdLZdb
ItsMHiuLgmYg5O1ZT4JPWCiUeBVNClHsYcJodFa3vU9cx5hP/Rr8sdUExxMZUl7UR6Za4w7BqWgu
a+LkZOBclLZ9W8mVgQNGH/HCMGZv09+umFAIqhO6QA64GWrvQ9yGAxwU1DmVQ0SsZ2cZYY9j3Jum
D4HKmoW2xbI+9Fj2xBh9lwXu066UKRSR2H5SttLl6J/jWa2kDxImgS+A3QGqhTqRhR4sVnVloTWW
qXA85oJgvnXrtJUCHLXhwEA5rHm7z8K35Fvi394cSpjLbnnmU4qyaOydsWk1bwnUa5DZXdCaTjg0
jY14AeHtyLGPLZv2vFqRuGnpVcjpzIkeHem2M3BUTWvLv2oq2otYHJ22C/PzgQLt7xRxcTqiEj5n
1R0usWHY+9UVpIcMT/s6Kn2lnZ5z21Rp6wzvIvs3Ys8f9ZvV+8yP0TNAse9zHG0paNC01iN9YMhi
mvBApk895U/QgdhtPlGP/FT69s0nKB7kaMqeaRSf/6LtiJgWAuBjJjyNVVcBNnVyAUEyQlyEHmHp
WFFPIc465yf0EyjqUyV3nmEjirBZxsyuxDWhCNib3vyr5w0v+NObcyGmElhlwhdeXTywCfBWK1+j
JrxLkdrHky8CiALKP07JXrl/cUnOdk3MgCOZtmm+YsBcgWlcg6ogzeCYBAYivbMXbCQ88oqkcbW9
3z1b+kD9Z2NJCqCDVIR3HblwC0JioGZVvnyrXz/k+sUiV8GK9YaUpGMPYdn6vVdSOi3ML3JaR/Yw
/MCY9vE7EoLQG66jBKJ4DZwPUQ+IZVmcRQZmQJGDuyqZze0vJQoXj4kCif9J3ZXN6WsoRcXyB1a9
/aBvZLsR513nxdKpp4VRLLaGjXTOXRJk15Chb1ORxRcR9A7WS2z2Rh2N4zgdDi2fhzBLkZrl+JaA
0eflVzmW3rd/5ihNFMurOR11piDKvK32Rd91jkYrost5L9aGt0QKLJysHcTx8WWlvPEtGz7RhpHu
DyjEHoa74pDv6Hp6jBI+ZDRvVpzkGbshnph8CPjBHMW2b4dAGJUH0vzzf7prLNq5p9U0+FplIpAZ
FEYKuPa+EU7v5E3PG5t3oQHdoVBIE5CnyfhC1dngJ4PXHPto1Kw4A/u++vpjWHIwK+uGNDEekF/b
+BhkIDKNV75Ar/A0fG5KxFnco+3B6Q02tMx3nCMfqQ7KIDSH0Db2/urX9+D/i+iWM8neUzYcV9Up
z8FO4c+XpS43L+lOUR0dvfXZ5F6wcFZ9K9t6D25HId5oce97X/OGXYoMfk/YMP/vXioZkoVkGptz
FfdtIWBFxBSdzwk2UvACneedOAU+aF3wynWpV81zVZxbotPUjbUgmw5R0xsZFSUXMT+lHI1deHMF
1QkA48XsT5Wf0jexiPK7CgH3at0OWQ2MWzEfDz8UpAJHKTYiTmtVDVAflYJQ4ZH6x2d6f3tb84a0
/hJ2m/0YkgFO4sdC/zwHTBXUH2jx/CDcQBc4XfBrgvNQj3lM8FIQxtnRQBFeg+THcvOPi0kPwtC/
M2pku1xBjWu61udv+QmYF+0N5SV9tGU35gidflCUuSJf9YT6LuCLyad9JqLxF//38dzV9QrnaT7O
yv4i7DhgmVIwoYDRQgBy9co4ViRfbRKX44QBu+zgOKSzNNlYfarTlM0YtOdl9B0IKoo+l/RSBoJc
RBPBW5XSUXh6h8/2R6gl9/bFohBDBf1jdZimVa2hN/3RPq/L374beIWiRRRNbffhkDLXOt+XGTBA
gP4PK0jY3wdkrdtncrEXjSIvz65PsWSqWKPObq6AhPMfnGVTPqswZagmowGZpBxujJU9c6B4+3+R
9d144DE6T+OZomPeGe/eYAirpGiiOh93gpAqeyB9UG73c447hfQLTnlaXK5eXcpCvt7qyyjfgoIZ
wwYzWmooMMNORBhzvbJXhzIByISp8GvfS1Mh98OPLTohdoppRGFhO/wQfWES3zHceAuGSRqPt60y
XbGjAOtJiu5IHfZ+dSKqcWjfv+CRy3jkRsHaKXpWSIfoo9kTmCMgtydpnoCmeLBUNRzkQQaL32Xp
Yn5uCke+k7zlBRiWkdYFeHdsSdnCg8XJ8wfggwIvCw08VPUMP/Hft/ZgWAuhnKXEj0Q5pjq+3h7W
Gh61g0o1m8jueH0OdFBvCTGWgqiiY63LNZCrdMAlMJj6tnwg8/YUAhkiRlEW0APj3qfJUNE0EDaX
tGg1UXhpOIrHv5Bt8tJVYNFYq4PEMkKzmg/wRZMPpEB7LRdq2PxXeb4E40JSd3Th1YR8kSMoc/xO
wiDOY58AeLk/HtK0DVXsyCaqXDSj5YrZ6hWNZ53bh/r3FNayACCMxeZgaBjkPi9San2PhvZw1Tp2
LjZJSr+J2t/DYQWd/YwjNzdGyVkTDB/X5z9dPNXRDfziSDJqEWa5PhuYbTMfDzkHqZO5atD8lzbI
DWo3E31x0pUhAsXbgUTYqs3+8/rTvQfen0H03gkqqBBcpLpcOZJHHPBi7udD381B/nlfKQeu8QQT
R96UyoEbJP2sn8nDhcr9jUzACmO8MEuv7tz2+kyFcw03NBSwVu6j3yoPaNuyclt71+D35L21X1AY
vmLAS92bySx4V61NrRx6lY5oJWU89js186pa0HryObng6/aceQonrkQa3Sbaq4lPBCk2hOo1+02J
LNFFm8aQq4tAEBokVj0bQJxighlAqH/v8U3Tz7AxMy+skW90UqT6Yk1iV/Bf7PaIHK+3FXmMrd1M
Fy+BXfvq7jfpsJdFhZjbtkRwpUPO731pL2PUYsv2qATX9WSRVGo+9WyhcHavSLUjKs4tfeuv1Mif
4EuLEHZcEP4EXj87D4UMvZ4JwiglDAqcNHRIM5N4KHII5FAG85Fhele5xLDtObU8khnzyHsCC/em
43WbWMck6exU24xSQpzlETFi41aVuZ+sU244g5DgcVgh+fWI8337P/1ffOWQA4puFZPfDqSZJmNZ
yQ93OXNXgnb3zs1g9yd2i31W2DPHAX+chFmsza9YIuOmGcY3J5mJNwjIUViQfY1onDn43RU3Dy6q
0E+4JKmstb3njnGnSjRCF3PU7P+vMdAhMB14KO8KbManMfnHAJa6kNIxX5mvyucQ9IrgFh4UwJoG
ElYCv4xPnN8vnTIreQck4SpG7TFcEFXOxe3jKh28/rL5TcHyY1CXD7M6RZwQZiWZTA00PidMxj4N
/iOhI0+1YtkhrLlzrGP3h/TbOFnIoQ8vTrRqCH4W+dPG24PiPhf39+/YWduIoKmVEIMzeodqgqSG
DiDgT9KQjb+G6eaVdP+GqSlqZriNhACmz/ZRiJffei1WBPkkr1vIGAbkbZwaKon92Wby8vmZECTb
zXo22wKqJtq720bzB3LhIaX/wNRGLMJPNrq0Ga0WIkxO1kJUEMG0xf6HliOsrHBhx4+s3v+toUn/
5TGwW+/jAPqbT4t6DxwBodfCktt6dB3E7xtoX7diQIR9QMiQYix5zCcd4hIT0KfNIowWSRrsdT1C
qW2u9ui04FEgtG6pw1TOQyPZIs6UfhhYMPlin7D2bJEzL1U0YrerfE4Urpe3DqVtOeFAo0nY2ghA
rGViCV4diQkQzggHsM33bHPGZ7bdS+fc9QTMVjxKXCNqanhjKYQOQ3J2gxwUKY/MfzpLKo0EaKlf
B9hz5RLrBqrCET/bAML4eiu0ReoV5CXDQ4cnl16BgQSC0PX6cOK9AshQFxcW5GP2QwJKPcYFoOvi
wZRQZ3RhZgwWIZdgc7n+KJxyJnQYCqvijTso3bxznR540ZYFX1n6LTDeFwZ1CCMe7gbU9D8tdJQ1
O+mXbGO4VMJV7WVB/PNHRKanA/UaCVkBIcAYW+s9vWRfOygq12LmzmtSna61jen9jsnkyDmFlsMk
1EbI1WYtb6GgJ7jGXcpBQut9UipJy55qXU2U/8jfbDu3HpQH1by/C5RLgzAr2SRr1G1VRDkztMuz
Wq9uOav/J6tcTL23imDHWMxR3L8jCYIcFWr9hmDKl3+lmTKQizu6jpS21JS5MtrT4aEfQ2IN6afa
r753LgB5wm0GKHLYX0+uDNk+2Oioty6MYOnx9o/tlxTCZMMK9NBn5hmpx4csPwiPf9ye2o4yaen8
TtxlvEGx9ZzzSfImjUnAmhLMGqskDhDqN98LUSGj+tEHztHDabo3tG8IkdsE6woDQqA0T51sySkq
pRlL/ejTci6WJJt/wYyE1RW4tuEETuBjEgEUNU6DwyolhBHlg4c3ySyS1tnUogTcgQV9w/ffpVA9
6eo92NqbH1ep8pHfXqVIwUZwYoV/xpKGeUl4+v1L/Az0FeK3jE0vgJXDFkfZS+aSkexYwKCZO1qg
z+1Pma1YI6EzvvllKv+JUZ148C3L1fsFFgC0lcSFOOL+0kfCHIZ8AG+ZgdEe6Xa9o7zfbCNb6fJE
xrtrn9Jb1MAjf7wUsQvN7NdQN2dbk2N8EklpXAHVydZrkKYbC+/1Ii4QnATeevvyszNolDXs4t6v
zBwotFyzHJDM7Ze/ubxNNEV5zIKDGM1OsnSj8+5cUFAsZdYqxLaDEoLxHz0O8GfghNdBEZZjjfut
f/bDJ46Fue7XUg9egvxnH4zBOF7myqmM4d7x8tBQ0Gt+/M9YQpc3yNBJttJtuXshRMeKOQPirfPp
h8mBoNAXU2hdWOTl8dmrm8fJeNlUzyoUJcKpc24ubfIid14fePJz5M5rHmukhXZS0L/Ab5zMS/A+
dx8Tr+VbUTZF60+PJEzGdcklZMeX66ZQgbUI6vmYuj5vi3doBafjxvJTzgWnN5hDaFzxy4V4cyLR
hs3jtHFsP2Wivuf6PVgKSkIx6E/XRMclKLiGiuG83xG7szfgfz9McPQNK5+G9627JYTrQpv4uisu
medCDmhr6Hzeipc3yLt4yCCfjIsUTQBfxTczitClkSGNNRBujkqWSVXN5YUmplvh8KrNq589ZB4e
cgjcNR6RLGIUDB/x22JB3Lz5pvz4jq25GvDEve37XoLjF8yQm+9uAZtR3VDfReXK/IcnJma8bXq7
Oc8nk4TZ3fS+K+yyGxjHm5Mjc+On1UFIeYBiMXLOFABzkt7rN8FYVObV6bcDpR6Ny3B6hIZ/LZsg
Gu6EdhXXG8a1I0ymAWkI/Wo4uv1iADRlW2e+vLQuVroj+ji+8zCRL1mdDdVp3sUe0GPyz0v6/S0k
zOgJ+MZpV0+Di+k8BNokbU8WhTFQx6kMMbn8GMtdckNz7zJ1CujNFWduwoh2nnhNDI9oWuaLU1Px
wLdUV3eJ5DFgZgXMj573WlWzLbLFewtmNCtjDPPtxI1AJ20tOmCDoLo1CasYG06E5HVgHbGyZGm/
7pSwCccwttmCMDpgr+TEMcYAujNGhoQgwNGOayXpB37I/kwjM67Ut8TcRKSxru8KScmomN9dj3Hd
Q0JUjw4YazQ6knM/u7QjVa/7/N5QMMVgQcZSl1yLmzaLElAU8D9C4crkmp9xhpk4OqLk/k62DsxY
pMXqq4SDXm3pz9TEcSQBpECoUvisPuCMsT3srLBzem4Ln8OAD5t7bzHj/ZtxijDPJawACCDm5MZO
xq6h2DIUIYUhXMsEaQdaB/2rx+WGRUv3+PHOYUTryIL+LlP1VGCbxgR63dypxYic4f8S9/W+HmZN
t0r19xKC6QQHnUAWPEucAh1Jfs1b65xewaAB0d9ttLrK5OuuOiWlvNflyUisiqOt6xvt7aWBEMfd
Jombv1k7BuBvfzcNw/G81jXt0/DkILt7x4YE7G7NsQP0KYejhwTXgOj+23n7Opplq3FLsCdtvBX8
+8KlrOQzdY2Ha3OLycKgGTKAMFUvBQA61jBYQsELGgZqj2Um5rYFo75KHQTBZ/xEzZBHVmTRWx45
5Jj0UUJMEgLkK6wxYNOKg0Lz95RI1D4xBt7Gv9KuMQPvhvGOtujSgjdO6lX4k9iUGIHp+RfGWRWp
HwT3rMHUCVG1jCvPAR19Swjq7W+Eljdl6ymbgMvAIFmiCcULZquehbbdRHJen0JG7kQo06m1YviC
b+B3P8mQLMMNja8uY6w3sF1JWvJzg21Bf3EmtCf4hA8zOdqqg+c85Oihgr41IHrCl7qPvr5odb1A
zdbEG8BzLBiD4NHUqu6dY1iIu8341EHNGaqW6waQEXvoANU8mp5iDhXUWzprXPYeKvOCDlpTGV8T
uoN4MBlzl8gvqTn1ARVshLP5R8jKrh9U5c0zRrJ5C2W/gspz1+Gzc0srrP8vwlQmJVK9ggB4Ik0n
DlQBzcFgVwkkO4FFvJJasopoqTWegM91TypIb/Yv9HvomiZrYUFPbNy6J4wFu2dXxuGmqYvb4a8c
OJOULQ9/6WiC0b0KWSakPp67es7uI4IMLwQ7AjQJW42Dx3mt/nfJ+pG1ibnFyJY6biarjV+U/vhU
NZYeUyW0l4bLrBX4ZEvIncXCG45LIp8+HNHvnTkww5ThV56zzbR43Alq1QGQ+ihQL1JiaSh2/Go2
WEBHC9XKov6KPhjbReK2UeMcj1Pn4ATq3S+yCpwOg+ntEnQa0Le9L0SC5UdMoswgGjZdjD12fgsZ
ERRwTJNjloDB6hZT3JL+RnCCQpoZnrCWHXbyhFcbEVto/HYdJZneyt6zUlXSXho8QHBdnOIOK7UB
Pa6x76A8WLZNh+sAeH6nyvlD8xvuulaHmA8g8Ul1hkS+mH0YCbfXJzqG9aUNEXQiV6hMgSICktHF
q+L7G5hCTSmeCwppy0Lr6GCWu9UxCOmi2o9ldd/C0qQbPI0XV5V89O7SEzdM3PfWtRlZz+Unumei
+ntl6vM53iQj0dZPBdbwKT59Ppe7WPflgvlUouGxumdsZFjvacOwcbRgb9+euRE4PaSlDOIaUk8C
ZmKhi6XSu0NH6Jgw5J78U0wk4i9kWbW0WUoYiTqcXr6tVm5vNwNgZFReWAqhVnNWlDpv2g52GZJ6
9+j62FiI+hGmMRZSimgEBz02Atl4jRCvIXNm33/o1uOzPeCYu25IYQlSpvoBTI/sKCD3TddW6p+r
TxJocR/O1BU9H404y6YPNLM7tmBmeJUP4DSOtIwZcDsLGdVZxbkMYfLHleAo9382a8JeeByEn5Gi
ewD68LMWatpWHNJtOZkYRtpZUU+Q74UtfMD61Y7jSwLV2XhoJvRF5kMp3dBvxhBsQhqrPeujHetC
jmUz/1WgyLLFQvysebNl2+codgQ6Z97xZRBOoG7kjQdB9nsIV23RIiiikLvjSv9rmic8ksHmPLdC
7CoBZlvru1B7ZixGCsqysV8bHz6w3Fd82Pr6OWwTIrnQkSbtIq7g7owhE8Hj033LdoUN0rL19oWl
BBFKhcLqj37rwgo57fSWLLDpvtnlTVZDFpRQ9VWS9QxjsiKzdkPs4edW9URKkogdl3KH0PF53n7G
z7cp7DpqvpRcY4hELCzI3BGYZwyZFTM7l8eA9fjFyq8JuI0aztVwr75gFFJxSVmWyksILpyjBDIs
Q0Gy5tEpUhP5eqw9HCT/K5YkLqA6h+ZAkZtLo4MaJZcqwOd1Oxdn5cVek91co8XQo3uQiTczodA6
zmk7dufVlq357IDeBs+AYZOT3GGaa2ACep3gFuN9yZTAVki1rI/Y3Sq1toa93zEG7OBl5EWfSzKC
HXgzr35AjW8kSEIWFMkUnurFb7sY395dNZNSdNDKy6jdSKcp+GpzZnpyNY+U7Ydi53YZQWK/hmw5
6Ban134MtKkKtE32BqWHSixcak7A8KjBnZlyQQwRy2Fj7sYQNi9DGUlRJGQ3GOgox9K9tmcO9SQB
jElXxQ03wtAzLNm3/SuR4vQjKrumpXAMH4rjouSUYTsDLK5kBLv3YzLfcQ0SNUNP+deIOpxBLYJT
PCDWa3zxvivt6qVW+eY/OaVvfghDbBciA3RbkvXR5ks+lvYJod8xBDgfWP4AdlVLKZOnimyXSrfS
A4JLkD4jKFZOvXOkXP6Res1txbvx0vacQOxSYbFW3O0IU6aspcXHO4e9ButXRCK7kZLValbhj5bJ
rsRD4SIGJRdUMu6/+F4P9XMfj0HhuI2FkD5d1XcnT7BlqpxYDOsRvejKnIOnq3obc/q8WkHsTNed
OilUjsCab9KrtrowagxA6+l12WGlLnX69yUfNNoXAGxFxnuHZtyq/vWB/GjVnMJBTfsxtRZaRahh
y8GShaAGVTwgvtG6Sk8EQEocTospUbCnGi9alttp8rQlKaLIn9U/FgopSLPJvt78noTmTjlbh9A9
wfpjnDxoC8fW3Jo4gRfPLbk0/GF88Vbg/WX8G6/m0SIA1+GnLBcoSIWrkfP2g/6TngmKmi2qAbZC
vbOK475ShBo3q+gqbuwg1iPlj6BhPWcaDEDzngIJdJTWczgSZI1LFQtgjQIiUExu4n/uy4O5tYYi
aU5QIWBFwTVykZFjAsgzTqZI3b5slQvz4q/a+4d9k/7VW5ZOF+P+tnKCiDrQY76cJGVFbM2bR/Bf
aTX0JFWW10ydBF9Xg2Z4qb4TN0oXEaTuBEfU0J7KqKGxnFcKcsCZZcLOPuOahfnh9LB0Q3trMeIQ
0wb1e7vS2mXHaZr7H7nGAVeNY4saDeSFCoY4ChA6UlGwUGB//0IMVVu7fpRSb62mTuq/WPYXTptw
M8cRIzWq27lY98QvXjS1jRIlDMjl11rbuDPIxyJXtA/9F3hLj7Cz4Wpi/s8FNooWCOcnM72FcT0U
OjCTsSuW5Fbl1PGZuxS9HXPRQqvbKR1zGQKQ2A5x23Okqh7jagswn0laNS/VdEKGD4B9h2H7TBBw
M2290eWBj8MOppDfcrPbidTvVV5sAo2X1aAlHrlGE1iMP2qQBrHE3XeHR5jeQgIi8KINJdE9hMhr
HSIEWknneghQveXvcJRYk9RnSaZ/wXTyG8fx2SUsaiaU5dwmzUlE4IfMbvm1sglrqEDpw6F2N7m5
mpC6bymc96SK8t4B+acufWinyQkVmo6f9kf4wRzvOXPUhHh1TtWRekevoO5JBY17Oz2x00n6uLtI
MI3IPq3T6A9fpTFd190SGFe2zJNYDE9GZlhBHkRSKj7BYt3fi9MwCQmbTHeyuiNKN6s+MjvQi2HC
yiCGG1q5/mEd6E9Kt+vlRT3it3ENMPUCWRLXvsMXfQVE+F1C19lHGd+KpUH6pz0OFoUD2EjUjbXQ
wla/bcbO+S2TzmaRWbq2SQxtqldM8Zx8i9rP42sB/T6g+qxJhymCawfjKZYaxGACNcKqOzgstQQT
J+1Iymgq2xEA4Ip7lgaAxkEkzbmrMBZRCuQdi8Zb/ZwHc//3fOI3VdkzyA8inDQ3OXmt7Ko8S4lC
rhzC093DZsMraBDnPAbtlpfMX4UZ1hnzHWEpibejPFKwJwf0bWs0QwOGffv8qePn1CIk+pTcUedp
kUni5vV4gkoAn6FDpqjFYY3xSRV77/lNXdtfixVphh4gvr0yuBsVJgCV3ztgOY9WNQ6LQOwf1mnt
70EDCeE3XBTimNNDtE8vVs1qkpvSmAo0scUyNlETdaZcVL/6Sk28VxLaj+btAfliWTUTGRiEJTwF
I87eaD9ngSsPEIz682udAmAGfhJl0M3bUokOH0wd3PCvtQFDUtHI9DAhRpGNu7Iky6V/NeiAdnFf
YIXaF83RwdFhazeEvLYq7EJ/3pB3HpDCFQ9UhnLRyZRDCVxZzovOTZzlxYW6B6qHh01gkSdimc3c
5xaaNT0ZRQcRMSLXTiY89xNUvJobATTiVO3JumECCoeg5ie+v7QMlCNxAyy6t4vMBYJt+bIvEABM
GWkSdkkqMF0Zoh0o/DrMzRFd+yYXb2NWyUQVHDpI/MXR112Cqq9t1xfQ6P3hIHtN6pl2DqwnUTkJ
1gF9HlTiyFsPk1y+fgmRVJ40ZWH7KaMuhigp/wmcQRE0PEbGtwe8ieSmvaJrL895OdG5gxMlh0cR
Q1au8+iClNubHNEudDFjIPqmR9CkyV+eJYkVcI17S83PT8PrA6CGPelLP3MObz2lZ5hPfgubaTdW
fR70+fKSVLv6DIEh+QtFqzR7wxSSP4VtosNP90xYULZXm0sYIepSWNNga5a0Yo11XbbzGhQ5D2jG
P+IpDbdCqUfNGqsXySffOdQfhp4I6QHcJ/qmksFvXStwpJJreYSUSAZX5EOe3f6OWqnKVYCQmJDw
nyYy4DpAkplRmBHDPpBT14MTyrQcnZo/qAbiLRKUs3m9yMt2ZkxvP2imATiZPQrC+PJoyrsUPAdM
+Xv2SMr12xBEbfjtk6AlEPSPBjKjC97NyJacLmFt/lonYTWZBudiBF5co2JVfU8YLQl29NWnIsHR
e//9AIcXOPm5UR41RCYW3Bj2otx7BlX5rK/NtwKUb0jx6ExjGspNaKTQXjG7VQndRSLD9WWkor/W
KD5Di/Y1zDRD30ahXU3wi/zPv1Gfo7AbxcsBMioEkVhi20Yu+2F8mjm2V/ZTpoBmR6WC2BytmhHG
CzFl+14Kx6lr5qCrvRZqYiIHKDqAmbvzc4SZA8e5J9GrWmA96LMGly+2Bu6vyRxFydUY0s3WxqTf
Dc/RZ4a8ZO7eHMHJRJrWAaNNvAxWaHusu0sDdJlX/VnPE6/cNAIsNZE+SpR6nzMUeoCrLUy1H4a5
XM3zTRPIcwdh4qYXOIlCd5JIrvnZQJN1JeDMKhwL3WTpT1WffjTIvOGVLebHyPkezxv7bqbYew+L
oaUj35NY/8Q2V3M3l1AVaG5yzFS4GzAG28uJW43VLShfTYFpNBwws5qWPKxydvNxAWNnvvyyNxGO
PxOEeZI/T0NTwMqd4YK8SQ0N6lxYGHlY81tTmnD4zw8eseytegwZnb7keILw3ESSkUEFGmdq1oDa
XwWmPF2khXsmL7Tgw+6C+Lkipw3OvRxgaAOm9kSR5TNu99hnFTCSc6y6uVwe2Ofn+3wA1CkPLtLh
bWoGC+mFqbwZHTlbWVgN1PJFqzLIl1QVtNooqReDuQRpkQgSpYXxYqbNr2GYT/5wy8LkqggbQJKT
TKWU0/XbudbhYBfywdUr9bMGlUGGsrTVNZ2KesJ0YgYs9BHbUNnIzNUNrRTUp/ciIg6qoxecbc3p
vhLxjScrZfYP0++ir4SJ7DoMJfdJAMf6DAOz16IooVtXA+LeLQgj7gIjU+BkSEoFxAwf6HLw6GTL
/c42wM9GKJ10GgDQ9VcrBYaH+a58k2zszPCocP46PNxZpgD/T0K2ysXYtfFB1kSzHWFrbTtPoMnN
gCbPXKYeO2DVPppxKj+tci3i0NQ+IKk78Zx1mrwUcT2NMUv6krFQJX9C3nEpbhqO+222y9n/8hZs
VR0XJUUDOD44WKCnHRQlHIZizCLAcd2nPYknsJ4nACRaWvA2X0SZW8/lEbkVC4BKZ/JTVBSMrJLd
r21NsQrtKX4ONir9q/QMJaRye1aYtnqfgJBw/GDtm298k//FWvAHwAGU8WVkMM2IMx0FUnBKbohh
suuh7B5beRGBirlO9TyggsA9eaedn+3joBXw0VMuw/3ap2GE867z8zkLAG3Ia6IPVjteog9cpqMh
HOGGidHhr9mKV5aKDK+t/+7xPwdBdNANPHsdLHIN4XWe7U4v33dDfpoqJkGK1fu+A+PjxRtxqc/Q
7z8f/BlQ8Cf2NxbRr5kWAds5V1qs5X/8IH9L0iuge8EadRzq8zXx922hKq+Th8lp+VGqUgTQt+Vo
xk9UrLJm9Tfb9TLERspPo/ASbBWGzajr6JnREFJNy1vNW3tvmrbMYMGS4MuW1vGL4UnmNHD631vA
7KvVCI0kTp33JWofrptx91EsWQhuflDHs3kA1rso05BIy9qbWsNradWStpk5GKhTpua5WrgP8ISR
zblyRAlf9eqHH/WqVX0ksOKyShH0rcWS5dtF2sytE8Ng3Tm2vruQS77Tdmcn5spkWKgKis8F3N+0
RnK6cvDOCSdMWy6xtrCeN4jZwd99SVEnUGLS77Qe3LOkH/b7/Tju3BYeJr/TPUbqb/iz/uP75LL4
oRSg0PV+Aear94Fodl0GnhtTA70o0hokdzzmApQA1kpMuLidz+EW4RvZgnIHXDL+SHeh4AZO2N/A
trgeJaJUOjNxj4Ticz3V6h6Ma73bc57kA60Jl+eipNtfS18yqufh3t+AXA43ft7kdn7FedbDoEir
l9h9ydGFVZUipHLP3rtAaZt3NWqOxIs89nREYqyDoNCyU1Mj5z/XkNWvBR25KnAwVwgXOMt0S4ax
HTyfUjGFqhzyFcvIs5iMf6U7xxNya36E+ycEPUgfePh50aU5cNZTqhMZxX0VFzPLgSq0JVtH3K0T
OvvBB42CB9G59h3TXd3o4xaOSPFpkD6Qmz7SKT37kkOevlK9OF7jQ2AHd1TDqY7/xc9rwcE7S9yM
zbjvNYeSyQcRH20Mlg74JvfD8BnggkRWU6G5SpB73CnQoyq/MgHCOKEczH+1igmkT68QNq1KIP2M
GU2gnrUJ0HbgsCg/Zl3fyzabxe15aEz5ZqRu50YlAwRn4e17l0yt8GBsPwveDhkMCvqg/Sn3rPD7
2jnieAhoNP0O2rbRju4xKUxtoHyEYKGwdxBL6CHBPxG+cW75hjwalEmM3YWbIpxBiKHvkLlmqaI+
VB7WYbHpRdC6yQavcj7H8GCq7CWSYhpP687BBVhxMQsUQw9huNvRWxNl3YCGTLNp+UeLEnpgrOzx
MzPlvo/JE2bFxbXCqr6XlWEHYoAQH1q3gqTXeocGBBqWUkmWrCkC8W23pAtbcmqTcGCcGnqEx51t
4apQnSZsTvliXLs0LO8TcJIXydLRTb5VVW0sxloKXUHxglzsnPjulcqBZ53ep09gm4goXWe3gSFZ
MBN4z0fmzgWp90Ilke0lIfwFWCM6y+9wLXANPqjPacf3vcCDa8AMCDvWKR6bfYta/fvu8vGW/uaV
htWjWGijwYcRm64JmghBCz8WOksLfKhW75GBUsVBYHaTuPe56p1T5/RCChjxBZoknP3FxQoBAHGj
kdkYa8ddyuDpWTcqcMLHccdf2wSAFg3FhJD0JoVQBOObwLfrUrVhA1NvSxw1thnutK8e9XeDao7J
HNh2HJrdub22rwHQrge0u2pAZFcp9GDZ3h4Ta3QiZKQkZMJSHIrWovjSL2vi9aT3BJdSeJhXP3pB
c6CorwMYiY4bhdVSlwZ8xDSvli98fASJtjxZIaDrHj8Cn60esSg3KK9bMf4FeHdWiXYZTGpyAf5y
Nj0rT8SkB3jPr9K81PB2OkS9WeyBdYe4M1CgG12jycYlp7oqcsRUIF/weIulGF5m0yP9mWBxMyCi
6KS9ax6UrfMcbK5oDh+bck6ot0uWMR9xesZwblKcDI2WrGUOXCj2Jcg5glVrm9/c2qY5G74lrf97
bEZQ1DzNEC+5KTa6WbxT1y+v+1FOrjLNOwDaQtPHHT0xi+1Px1ww5DPJZcGowHmgza4W6sLIFdvC
+gfnQy3fTBS46ixkr+vjE8bbixN0iMJED51NwFbiRN6eaWw5CfLWWiH/uDephbD5Qo2Nq/mWzDRN
O0729lhyWItfTXvL+ZetbQ2OlSPQ3ZUY4c4b3vhOYY8FqDlxBysbkjV5PsfKzgxZeHgyqr132rR0
u1MLya3IKmfNedJC7n/xgjbOPKdanq1GPfHUv508c2yufoU+oKI3nR58oYrCxee+o8pFSiIUZ8Ja
3E/429HPM9971U4O6VohjmGaJTeVDGn2XSV3wKS1OLc8ufZ8I2fbpXtm0lXvCqbwDKZNDbf2PBN3
ocvo+XQ+lfKVjkE7rfz8pgftjfg6C3hyToQ2/RgRa82l0OgoHv+bVKx8y5s2A/5HOXsWfvQDIGIS
dYI4Yt86KmW0qipvKSRQfEU+uAcbEZeFovsoIQ/a52qaW7qksshSs8ecvMQgETEFeod83gPTjaVI
lZrPkryCuh3BY/2T+AT2VxmfHcoGycCNHZlykriW9EBzFarg1cE5XJuLFA0wedDiRiFZzcvqgDa+
SaB2t2KU5ktr6A3imBTO1L2UYFyAnhOpivIOK9vxIfbB9TRTSnUcS9BF7BM2MOebcIbwdYsj1Clt
H1bUagIvXDjjwKgQ3Ip1XhZJ+exfxIc241QDEuVBduw3AMGPlXmcrn5aR3gKkeTgFBtsoA+XZO23
EX2BODENhInc2rejd4KMjKQmC/OYJKGY3TxtXKeJcLhryOj1AdqMDvYxH+aI3aTrC9bKqBuBSIGt
5yjCpQiwoN5ReZyKYXAOzd4TAQKBd22IvCmUE3Pkvw7YlMBIHZHf8y4oPgUr3EwLMo0lXHuYO8Ak
Eynpp6AudvggLVYowThVNeejhfsKVNTSYEvf7TkdLkrgykbt1I4joV5jRHbqjlHBHJyj/B/0G+KP
RHb7R6YHloOgNcLRwoKNAIchj2fNX2Bh1HfxG/ozviztKDgMZ+T9cDo1dqSNnoc8UvMT2uHdz0qu
xZ+IUrgPNHYaOXe/bmDc/0Smgmpl+iFBD3EOR3rK9oWNRj/pHWOZfuxOPbMu41i0VrtLVPg49dXM
AmWvpYrzK3X1tB1NKluLuJEaOQ+W/6U3PHlQfVQJXe8EIl+EWPQoTaE+wm7GlBO+LlVd84loEu9G
9UA15YdqiziS29nadmLRo++5IFXxjyJ2iIt1xL0Ba3kJLfotbjBO42T5OwXolMhLFGFJA3BgzGD5
lAPP9L0P84dMiB/5WAoAMtlbMc7LlwHlm4F+HcxEu2NYrt7oOgLOoAB/CwnIgYH4/bHCBQZMIXqZ
WELNCYAgf4DVbq6WRiCkWOvRIJ3F5Ot8sVjdIiuHvZW8rm5ex3Sdw0u0NlUZ10P0eevQtba8kMVL
gO3vy7lBrHBXIFnm9XPYNAoBtSsf3Wb8A7KLxoFbPclWPDMxbMP7MogPH0Pw00JXGwwsLgOzrLiX
Wa9i2CPCKGAe2EpARJPoURrUi8dHx8lxs+JLXvNfnonY5nKUZPBm2ywK5FMRcBju6p562MUlvonT
KPWXL3ZSfxPiKi/4uwTsHqrDXJivP41+/YAxNWesxfjnJGQtZwe+hVg6xLHtB4lmpPnH7xNRYSUh
puRLtRSGl+yq3hk3nnU2TMynJNDH+ul/BEZDZG2HYmfUzz17C6zUThVFDnXZEXtRPbKipaFDKoOG
ohXhPJvvGXLC9wP6LTX63kK8m3z0oitRsZjaZnWdLj3mk9JUOeiHJtSsKjLzsgXD+2+cTfa1EL+W
U8aKawX3jwu/0f5aKep2VXr0e+ylbSVsrsQs4xg1luBZK6ba9K+e8cmHse7fQNK1n7AjwGAoRNC5
DfloPKP3vbxAWa0CLLwGgZ8Ls4YFHT6HbpGS6giMK70u5igeJ8MGuySPGubEyC/funCr/5sqLgCR
w5cYS349K4iNZDtii+xJH2BryE0+xI+hUWvIbKtuakgAQjhnJ5uLizu3x8mTw7DRZRsHansZ7kVY
o7XWmIIhh+XJYSUee574l+8KMfs9459+fctWCOamo+wFMj9vcZAaVv6uMzq8VmWWuDhFqBqFxtHM
S9v7Mn6X4RRvNjdbfBkOuwqhQOJf5syrHB6V3aW6R51zClDw/PvsS6Hc+QEyY8Zg7T6HIMi9bi54
pzy3X+mcVM6kYJzT2KHuBVUW/mVKIz6VoHERMhHvbAhuRCuHCcCcRRPAfb35Nai8Ysiou9r/VrL9
pN9XNEipvq8WOx/Di7ULNOqTjdUBTJlBoRgqluklnFI+dzoT8AScG5PVNFuBXjzRvcj1LE32KVtN
sSZ7r4UCYItrUHKzHCV8bu6qyNULazsPJLGPj+aWt/iDNY4LpWA9zB9hgcXIOzWMRHfbjkCMLy3G
rW2zQqeTpSSrPBRh9I6PFgAlPG9J1XDEChSIHY2CKYinvmWQ/ZydtKY9L42hWI9ZJg8rSBAvWK7h
c9RJd8yKDsciis2v9lDbsWuAsgznGE1I6NDBLIZ4Rxcs1+w84SkG8AgDZqbQRZuYJyJ2TIsau1en
m1v4JcOecg/RzMn8b+rKWGP0zH6rOdiEz5+H9z5soHBGWhg6SeyFXuD10W5vWmKp/yTb+Bbbsx0C
iD2bW7izQknE3NsdBYNar0BWxjpbqBsxLSBvhYDi56+UWg7tJKuLnhjLMbwEInGIywVex9uGVR1q
qBPZtMm1siDy9HpAt5vEdowY2r/DNEN8I4ko0HZe1nQYOKjRbhKNkuSrn7pnMycjy6KCo6/UQXDE
oQdGh4CjugoSlZaYMlMDiCscqhDuumfiaVA9gNo7WKosZ5Wy9q5VApPEmAO+EycPUipLyjjMp+CA
1r4IH65QH4PkGGkbcy2pax+KQpvYdnPrK2pfveipg7sItvgBe1tnS3Cdx7y4yrab5h/NfZGpxNlu
RaJ18lcMeaALv2rZRpv/21GOAIx35+so9sxTnWaZHICQ3JggdskrSD978EqZk5XPrzHrlsxL/CzI
DQ+OJ6Zz3K4emz6Qqha1Gg/7/z7/Q2hwHMqe+VYcDhzcDMY+uDarlHXDxKExJEAVIKPyup0/amTP
i6g9uqXg/sS1jgKb1JklH/0wwPbURNLbhUHIb9AUZkFjxrLUrUQWD4KA7En2cleg2cuW1q3tSlcT
oKn7wh27/TyQGouYarvjnvipLd6bIiKrs5UyCIBD9JnYV2FJinSqhxnVgg9sbluF5RsBhDqTpkMi
2gpovqv/XJsBIj2ow+4N7hL9rZ47q2Uk51YXi15ZEbSazOKNJ+W3ecKuWUnlzUIfVdpOKkPyyQTd
4bM7AkrNJcQB1jy6lOpbEH2oq1zDUGzzeaXLHZ4Maxxy4yiN2Oo8HkC53AE0glV0gGCPrL/w1w4e
ykCKFk8hjQmMu3ruIMNLk9UbkPHjkzhXk4iRKVBiwdXQ+8NYGOWLZjO8MPeu4qkyiyZ1XSae86VO
HLeRckfqwIhjt3oBtZtLUdCA40AU3gWFWD/4IkWHY+nZyJzd1UI1e7n8DK6ZlCq3oK2MTSGkyuFR
PEJRYWFvi4uttgxLHx+W3e/Sv4I6kXocPjoZthnw40Q4LIwb5B0erBbkC/Bejaw2gdxMAkcuRK1p
E6j0xX46zUB//GzbOZghIordM49aYrvh+A9scXsq4xDsHICX3D2VZO8Xfru5/MU4ZEuSl6qUxJvh
uZ7JUthUZPlVBlaWRzD1L0Vplc4J1PTF9xyinR7H1adO3N00LgjmC7Pk0w23WM7qAX7JxYHTSKm5
ZxcotbSCh5JrA1lP/IYlIa4R2qHl2mUjq67+kSp2UWK3C3/uO9KnJeiZWnD0agKF97skFYb62cNX
Z2BL8anL4bAdSillxezhqx+Q7ALGaeLvK7+23pEyCnJmyU3A2f5U5oSDqwnc2ivHCEOnLczXallo
lr2p+W5+fspG8fcjVU5BbJcafriUomXDwTQxzaX7B3F1hXcUs3Xfwf/yLBXHg3pmC+3IcrQtzRnd
p7vNClkRJvjEITeqntguU2/uG+AERk8EaAH4E3puAqGz1f5Hx57DDXzE6v9YZ+kG8xxTAu2B5Y8I
gCymzCK9ARz3CORqteQH8x8O8UL9dAzrG1M8WqOyphBAu2BVxQngFI4GLVolKI3sE0UMgifBTcbU
quuKhS34lk4GKmbsiNLoex0qZ3HzLKO7ryc5PNlQLzD/u2euANoj1BnJJA9wIeLVJ76QCYjkZ2JH
q4ao6xg2YpLOYvjd/PhjZijEIiO2lCSfEU7j9eJl79luk8ZPPfL4+C8v0a9lfyAblVQ4wDz6jXHA
oB/cZi4wrdp8QVJbeKHTjj+OzK2F2AhWPve3Tw20tsl4WhVkJ0AMtIhHoM4Jr/dXissNhpjGDkry
+Magk9y2bCihJWrawD2BBAaMlb/SHLBgiGSBJYfQKiC0xMaFvWw3Hp4KwAQPpWuqprv/DzY1VllE
405gajHU6D+W81KOtWuIW7LTNfmJ6L0OuIlAMgYsNu8widB8sBg7o3LrFU57Rwv+vJdIrGp68sLf
Xo2HR1EC/iQWfcMbzvV4Ujuwp4ZHlqKQNj/r4q2VKjyZObhRJ469hgK8UG8n5/LIUDaM7qQYxFRD
l86d9nXd6e74yBx4letONTS4V+yBCdsL6W0ZfS7QpS+fUWBEuiMHkBY/Q4Eb101Onae/A2r4vvww
TCCqaNYPIudfoJrZWKSEFg3Fh1lQUOJUaVxDMINQ5LY9MTE68msqsis1vqe3mkCw6WTw3imJzliS
RA2dat+DxcGdaNyI1MN8PlgpffKbBCOnobc0Uf6AVPtzgbJnZIrCzKgQUHU9WSCgFkx2fuOqBZp6
43QlNgdqh/egnEbSoDH5lYvMTyccd4/spem8YCnb1CEHIwXWr6ixmrSUd3PJE83HJRh9yWl8ZRlI
1pJpsvTFp2IRpS8q/t5JFN62N3FoPXc2LgYUYXaZmHTCoXOe8y5xorPXI/63KyIfBixmjY3GaBah
qMpfPvpSKpOEG/s8r4daNj6ReWVnD4io77njegxVkZfNtYJDTH4NR5mf5AR6IA+d/Wi1fgXJSWKV
0ruCQyeArxhtQKqxAwuG11jzyqiLsfmNy5tKP+tpeDXIA0wBHOQeVhRVthXFo3AdYUL5u7V9Ozte
4G1apk22VTMCRgqQ27GrsGW8o3wX14oic8Axoxn7QrAw4aYt3AwlSPtU4Tfj1lGoHmxbJJvNmSRf
1WGdzwFl9Mm1v3xjP7CKCeRQxoNBQu5TaNjEXCRrkL8GKV8wgBLNJKLgy71tlpcRcGz2OR4MExIG
3N/uhJN+zwAnv4S/BthjAk6cwj/OPBYEIBgHZavjvGdfF9/oF4yeuM5xXbVkyByTDwyhvs7IvyIP
evtNTWWtW1Tv38Du4sXFwWGxssCkMblVoQs8HfEBYq02RYSArdymGuKFTwdkvMZLv/LO784JBlKn
5+IvbcyQ4cICAeqKpXCsx9kP7+k5ER/zAzlkUISHOPgDkn1H2cfi4gFUc1UK88DsMQgRexkI2myz
+IjDmNL/fjtz06XAx3rCqzjbV9R4FBeONm5zckxkE1N5RTt3gSzv5I0/afkl2ste7BWtevL6SJcP
57oSVj5WxsiXwJbUPgQO2X6VMQnjs/l1+fWGoFR9GUqeJhP7AVKxrQpXUnqo/DapWVBUP+sKfIWN
BHNepRHTPDn4RttLhuNqYoTRRNwH7K9NMoEM0BZggfSTwnCJKmjR6oK8671FHWZjXAgn15CrNz4T
AO3+uBCUNSkHfQqbsmsrYzb+D2yj2LwNXZjFv7Nd+VGuwrVPRBy0tJdgq8ckcXsgJ9G3QFCE2Xq/
V+yYC28lIubWVLIhH5lNvr8vzYfAD0zSZR39A4P0rpE9riTmg+5JjZ0P9aaY1++PllF++g63FzfL
Pc90w43gGDtz0XGDZqY39kb+S5C3tMq3iaSZ+p7A95ikwL5OqyBFt2UHb91NHMxYcVqBfR2yk8+S
8lRYzb8eLNbQIRPHuqOObYAmri4tAFTF+rUVdX3wttbXorQtKCJ1uNVjKVj72fP/Vdbq2YuzXS6+
/oZy/8gVv9WgO3Y16kffZ1oxTrsQGG73bhSX2oo80frkVRwQaGZwzdH3KIuMGcfsNuWeeMMVNvpM
hqDczYaRy7ZM4m3+wa2R8C+e2kOJFU3altoLLW3gbOQC6ohrXPpqA6xgfuu/6bs2qPPs56SFzKFE
zCJPZHo6cjqe0HDV5u4EUcvZEOhUo5sVlQVBbiVUqWWlXud/JxcerFh4Hx1qJjbFa4E3woOc0BkN
LoV6dPmhfAN95hQSV2KnefZvshCVlXHG8+04DEoE3xPWYQei+Kr+Brlj4f8/tJjL+pobItyd/mgC
wGNb0cN1tlH30inSzaWbzH8IluBm+cCl7paMIObEzWWTo2SMNJnA2IwnFH7vn5vPoGEDuDgNAqND
M++3vF/uoLsAlw0kOOBJYeBGnl2Y/ZZiPtM6NljaaNzNCtzocdjtux0CYQrTqYCvzUTjJi7qRsOc
oFiaXLOj0j82IrfWjrNczn+F0MsuFf6lmX+T31NrfkTfp3yDiBoaiJQL83iwW5jy6bi7qYAWcsb2
ZKv4RhDMDBr8ppZqMEwNg3U/YPuwIw4eDsm6HjPKxtxR5GKBXzyBH1yhZ13a7UoxKM0ygnmhLgy4
4f6REbcoi2dyL1Ji8RHo0KOMH20UMMmn9/7p/S6zm498zGpn7LnVShuzsuYJB9CwKtJSqPwq5dKT
lGxElSxyKd4xl3YnO5/dniHgs+uj2fwcWbtwVXLj0wBKH2dHv59TBWgvsZ7bnl0aQzs04/FWnBHT
UScmTheInGOXEPicbbxh6Lh8j3qXjXpMCw650GjWyUBL99710sdhnazOsuvEWGF0RpNlaFpWon0q
Fdpz8kiI+3nqt/Q8KHx8Im45h7Bg9KmTflWAneWy4YbkeXqmuX8NzlCuqwMYAP7ZlfKca+L7kamC
Fcjz1JkUduw+ibasFn1IyivO/RioADl3ZgfWrpNxR5PQ5JrwaYicwP8QGAJBtVDaZjniJnPvThSy
jyDyUeWbobJ9w0K4SdbPLp0JaDig+KkS5SPZEzvCRk4xRen/+6T7ZabmgY6c6QkGhxAWRkEeyorQ
R9bn3eviCbyFo8DRR4TZNutofdagarTGVnIk6fWlz9WKDUZR80PMFlosAGW7Z0aJXuapjPufXgJD
18C94JJtdvMkaK1S75ggKcjg57gm0V+jU0zggE6gePXMuQ0FThKYxm17JS7hPbX+K+hKteJwD0TJ
iT4XIHpolmW5jebQfmHkMq8JTZUSZo924R/p5OwahbhBXN/P60ZBAOSWKim7jbeGnpPUnvK7MPHW
PcObOfg4Iv76YYpglsS4cKo6zhUYN2DBFSBT//iZECwNmel0QUBnkIcgZX0cX3o04QkXSmLCTaqf
/5Od2E+OP+sPenZgdtnMs0e3zYRYC+65LSfUBrVXHxrq0YV5ev+wx5FhPTvoU/Xh8ULCyZdC9HuJ
f1x86yOdWkEbAIEXNdANrmfNydWSsoXvYrrqGyIfmxLjVsnrFfY/qmeSFwdorXvlJYp0TSc+Mb8B
7p2LQDeL8hDDwHdIXbc5h0A8A0gd9qWUdGV4V+yRgC67dQcfFTc91KN/2Waa/wPS9HoVIF3PFrTE
pj1+mRytZI+EJ8PEuaIMnRbop9iboifjWbreKnTS71hMunLvsGFAc3j7onj90EsHd0noOWBeshpP
4YQ4KzNcnbfZmI8SEHLa2ZVABKXrpXmjQzMbTNyPQMMtlevUZL4VhmVdpkbCai+fpPpvm0TGdX6d
DNEnTP2+z5H5u39Az1Z3h3UZxKbvSPGos18N5Vta3JcstUTfbzPegEJ8gSN7RXiOLRlvkNRXrvGD
cMar95qKZufV+dfknSrnbLzgD3V3p5jaz5NTNIV41IkvMGu6vMm1mmomQJpTwhsoBXmbfn6yp/7G
v30xkgPsFDhCs2vWKJY94c6gehSIrgo37diUYF76dnG/9vGj7rWCp21ueOwEO0u/w7f6+3czz26E
1/FTasieY9sXEr+42KOb99PuDQ0dr03OEUc8l4iW5Ba9JViZWkSdI+qSQ345wQo5YAhOh2Fr0CYJ
oT+Dc3INjP2w0Y1sB2BxpahFnustsH3aQvSv8gXYcdfVFnHO6/yWex+wkZPXRwmVUv+cD+5Hc4rU
QTzemeP18PPLFLljGZTi4ESmHcae4eQAyFDDFyXP2m6GBVDZBJE7m8sQIDPTfDMxWoiCxjLHLRQU
vr3lBRRwJCDEzXFB6yUy4yvS45IDWfemocPl/btMvEwDlH+tf79+tZmjmIsD2jW+U27r5rJDL7BG
FF+e4eH5jz+Uj3JtEvYZgm09TuLq9pzjaqJ/2Psgt470O5y5XGeU76VJdJeMoTcZW5QTcPkbKHOd
uekmd9vY8GiXWZdObXuFgboL7gCbAeXA5yJ6BEqDL8Vwj+QXYi06hQDaboxJ64SU/+lOP2jyhgdf
I961L0PjUty1VE9nXm6XRTt2ZU4WodevK3OnyY/OsgJY8Pib6Q41XrRR0zCDcHFz5wrRsfmKGJoC
qBpzNbnnOMxj/iQLk9tD2WGUWHpZx6xK/Aosyed/dsNolfctTIGS6lfpicAtUmYsgwpXhWQn2veV
tRPrXwc0Tta4N/Qu4hHyLDnUwhj9oxSZ1rkdY8nQkWzpboWot0BvvhR/EAvNUwEbTUdLjSXIfaCi
eF2UIrwMSegN1q4eehbwrZPS14M3Y8laUNsByb1a3CdwztZ3UJDFiGjW7TDD39yWObHciXBKw0yJ
h9h30l65o8n1kQoHP6PlfUb1sHyrOkDRtPPZJEfzgru8wQe8YNu047nqcYuzzL2U4pf8c68Q9dB5
g/IrAcW/3Rr4IX/OXBpwEnnrAwayBbAoC93zeeueJxLz+7zv5n/AbTblRAgeA2OsP2kpv28d+9wW
B+es3RCdHQU5KTMLRwUT8Xt7QsOlv9swAJ1ISCtQaJZUpRST0iEpd6NDFfm94r57wj0IfQkTS1mI
6flE46Ni8FRbrXHHXze8qdO0/RcgJEKKhL6XcMNeLHFAB+9/2IPSEyuNz7AEcN034kWGsHS0x+pu
GmxeX4/aWvOKQ8XHwsAGNUuVRWsjLvELc5xGYFWFJZYiYScYwP2K+LUIyMwYNNZ+wfP4AvVABAzT
BRTvE4M/sMiWPe9KrCATFNVl+wD1W5eXisLEPmbGNBc7Yr7S/OG0FOdbYKObkX/qJWw3EfwcRTlm
ZsAzRjFUE48pnFcTg0OynE9VpHR/2NPYXO/dUhL7g46FO4NLnD6w7DY5S8jHsm7t7oBNAM1p56Uo
9avupIjORJwRDIWSNT3ijhpXu0pf6Y+YQauEmHeRD2tF9JMQBln9tiIwin28VJZ0VoBr+6S9sS/t
g0j+pOOOoefCu0LL9jGp+lCK3FgSQB1NsS4iYMKsOVAvvzLn+4jGsF4wLrgpm3tXnbI7BQCIHH6O
c196SvVsAFlLvaN8TL2W1eKW6zGR2b9kjM8YY+ZigAbDJG8/tkV3H2LUaoP0r6yehS3+r2EugEhr
8S/gbvBiz5W/vQjXbOMaCnmulsrG1d+QmM53GsfS6o3HBFw0s7o2DCXZIMEhIifNdE3PBtH6rK4B
0t0/GXgZy3i8f7IGLgJ/IBRyzkYfejEn5cThue7OJDAjcBwbu2TqMaCJMJOjmQAS4s0sadYFYpUq
0ga+8RxZcll/RSPef5z6STGbyEdcL/DB+VvkD7X3E0Qco20i/dB0wDDWxf1Yu3wGYzbVghCTuwNm
5Pcv9rZ00zBCXTqQiYcFEGpSsetXn/8SeS9v/avuImRs34nJnd8Yh7yrWYgcm42gJlTvj/bc97eK
VMaP2IDwlNaFWT0CXFoZPO8xqhBrYrwFoga/h2ETbyRr4zpn9JLupo/Kh4K/u75i3ZJoGX3nOh4I
LTCAuJ9I5l2qrpnn9Brj3Pjb0C2SMCf/6LWnNTSMCNq0Ah+ao+7Md3x4I47Kv6N4spLbBDYw5yir
Gr9fBSmIkVApAK6mK68Q01Vuza30V34xJpnfcuq0Fa5hJzidC1iTQ7NAuzm3AAZaa7P895qIBJVc
ci4EajikYzmpyXUg7lZUc6DSWhYAR6r1KXgx2yt/IWBh843waL6RL4ZMrQVyw3IAu1Hro9C8bCj+
sHHncxsrHLFPv/RlzCAPohco9idPi4L/vpE+FSOHsit5x6yBJYH34dskCuLhdtIIvFoOX0R6NfY5
Okoe3wRcLLdeoZVizL2c/sZw52TFXmswZaxXMuyvp1t+0+RghZkO5dCdPmFcdjaCkOXMtlk3dsTT
pUqGwPDRt5Rw98EMHE0EyTK1WF6UC0+ELuW5tgF4kvdoKLMfoYC4k2r+LkSczLT8BGMVMpzGER3Q
d4VTfrMLlO/cjDnAP7bMyxiRvO/t6x+7CIU8Ix6STv7ljRskNGot7lccnIwLrGr5yyFBu5qRi/1T
wZ+pRKGO7Rc30m+NYw5LKvRC048480b4wjnRXLpNbqd020fM051xj0/+brgI7E7mpxkoAaHijv6X
WYDXzHSCqaYNg5+LaCtKXpukX1wqs2zB0BWYJWOIJ32M3sPXF5OEbtQxgfaWMl/BMH3+vYghPnzk
uxxvl8Jof0+s3VznQy9RmWv0ipJNwXQX2W8wTjKUFfyv7eTB7SCUpOXLWiV9YnuRsSMxTxwUbbgX
5tYqqyeL8mic43av1DKGd/gR1vSc3jyW38f1hjy34wWMdufeKHx8S3aNwp1S8aMQMn0uDCXlgXuI
nCvGt6GWI338Uspct5aBgQ6qQIqcSdbqHXqA8NDJh2NFi4p4mQvyLoCkLJ+oBWbCNOv5ZsVz7mXp
B/Jphq0HbN37jXmVAsampPalSy5n6OQfNRQy3VNfYnS8TrYGIWz474ZNz0dft5m4J+MrrM23U3J2
E+dgEPc4WqoSBCQjiiKBaC0L2T7QEiLazL4e/Ry1/qePVNUNjQjZFZQzFYmem/ipayiUj2WjpwHT
O44dszSGTWYnBiZ1Yhrq7osG6Y82Z2gY50G6rS+IskYedxN9b54vwYbQTXDFexZufsLiUz17i3l6
YjRQtmDucm4GATs0EV+uSDQhp8GiZfv4N2nA3EP9PpANSfZC2rTUW82H3DrqXN+TGoqn8uDi9QlA
FMyjzRN625EogVqAqI44+pFjGlwGvyQ2PqeafQihzPirzbXUrKiofPumpy+Qa6Xi8fOlbFLdjzFI
ku2lbydPkAF29k28yg97F+1ZC3lB//mixoGRXTFY5GZqkGhMilXlTwPWaGy33L3o7IBHDQTSmnsl
r3q9nH6MXMyWkRjAm7e8/TA8QmCNKg2xGVgnYQ5UKr66DJVh6gGz7Cw2/GDrT2GXiB6KuqdtWmBS
fLfDvvsZ2QDBboEtXjEWhxn687WiTcBoxck3EPHiiGEgiU2Cw+FqRGuImqickg9bxVtRxLiQ3UUO
p0YDY2nGGNV7eKZolZsbhoqenKqxC2yN8K5hyvBOSu/uwLzr3qiTXZaBTRssbanFa1xc1HGc+P1v
dckjhdxXg+ujTz62JGu2nuQMm+cbsEwQQmiwvnxg1OlFiqfPLMSYFmNJLUSb7kEs+IQ0iUkh0hNA
nswng74+MicZR4ULRMn1O1b5LW2ws+gPG67ORjXU7i6lsJgIN/wquNapPLcom7UMCBtvO3xuQ3gy
ldMrhfMQNHXHjRG/qdzCMnzvSF+N1D35EUfUfyZphHhBEZtS8rtT3gNgmh2SNXfLiZbQ5764Dk89
csnhlLRaYIyWah+eKJFjCrVMUb4KbLnvf4rXEN4+B7ljMlEEgyLgEVbnyixjPV/bZYv7DgBo5Rya
N8MCVmOkQM5Mb+GHG7h2osS75R6rCsMtmfG/672mJ9uxJ7sDOzVj7HRTKX9/UCVBNSSSts76LtED
3qI2y1k/9M6zdAzFBFsA+lfexETpJrrneupEL/TozcTwWa63H/1yyTtCV1oKc0fQE0ctwe+OSHOJ
AV69YO0k+p9QsYQjXzgiqmNqZLX2PtTFVh2TRMX1TYFFrgrzTmoV6Vp985QpS5JrgDoBPgGsnS3g
S8zQFkMRIIarqo4sKSk+74vhsBmh+w0SzJmRp/XjfS4+1P/NCdA//t9MWY75tJHpoy8wcrkc5FD0
e6Fvk6S+6gol7geqk3yFt1PnL0bnU3TG3mp4bLC2re/3V6KYFH7zhG9PnfYalmCzD5ySOujCn9mQ
vhhkbKrqyxMIV7As0qO2089LFTd+alMuxbbr/2zeLNaRWwtdUJHlljDcv1tQv0TE5QjctRYlRSx2
jJTG7uSw3r8POS2YaRa1kjYwRMUBTSoqklSPcWZjgrUgsMFH9I7U8VRLS+tqritol+eaD/LQTzEs
lRn5FVsOpyvKnXEX+EVSyN/b3Y6xXeZr43IB7ZJlLXia5hbXWVLkhRDQEFRwVBJQgiU6DQmMF5GV
YDHKyLWY5uf/fZASZS28LHKVEl2jNDXeDtSOeI968GVshebF/sKMi1FpWgiW3ZqUqGWB8g2fFljX
jvbe2H3SxGoCQbNzJWDDE4/F7952tsIul+TEg8pL7kLxhtcp9dWGHuqWYQ1M/f/lgpBI/MtUcW0N
omsk5j1kul4antFBqTpl4z++0kARbPJ780HHTc/vT0YQBDKA/TUZoYdfYA8ygoL0ApKI/+dhgmoK
Uzr9doTd8qmb9HN4IxM81Lh6T1GlikRLUh5RtJlgY9cHO+UuB0EHLztYZ/JFSG8+CM7/dKN08mzc
FN4R/Go1LtBAeC/SZxv1Jl/SSO84iqisqLHA7mOKa48G1dBt75hMcbcxfiLqvgTGcCiBTRytHxKa
wwtHLIx9tFarp8KFhtii6o4d2DLgXj7ltTvNfPl08xpslimjGntHfycGDjglYPWFsAmY6fToaA48
Ru8FuK3CrvFvufxYPbLJHDEwX09imrmDJ58ziPKlOX3hqeCG2rTEq9nKaPE8jOTOBb8IM1JfPevK
+EX3gYZtMWOOU0wqHiypglB5SjLD+a6gJbSF7P7a5MHH2m6LMWWkWLyYhdjMZCjzS4Irc29SEgew
8yzMxnl2SzQXxgPUZQEyIPeGCw0ufi2xH7slu0cWaTpF2UpjboOxrQj8Jf/ouPktBBX1DEPnuvCo
UQsHMdrYCZFGguSqzI/NIrxCsqR7usFwyMSDageOasLtbJRjVEerZlzqXq5CKoZnQzRbBA8jh4k0
UyY9sbWHLhT4k/xtUEm+B1qFbUBQufLqMBY3TOuBJlWmJyAUa7kwz/8lXdw15Tc9b3o7PLDRiqcZ
SIbtLc5/HqEpILqtEd4O5uIFeP63qcJhfaUgJ8bEtbEeSvruqLt7DSI38S0LjBeTeDuKnCdS7IGE
2slo4fFtRneYAf5ydfwimfBt8OiiCBXe2POpE7sg3u5a9uGuD7X1HQc6bfLueNf6NIniqgEDN6dt
hsk9nFSKqBLyO0xuV0U4Rnax70akRjWoxGy3yxpZjQ1IrzoLc8lMt+UmbGuYvVNMm+/toItJaUER
Whm6CaTRwTOiB4hwBf52A31xcszA9QN5i3Zycilro3q/FXjaRuVaX9E+R69XnsWfoQrnLGUVpOl2
JO6XHgsPBW55jBM2M1quuAPGlJrk/t4CaL3XXuypOLmnIKpj3dJ0RcU+yVqEPBGnHdh+Gjn66aDM
Ru9SwogTJ50e4qU2qyOdv2G/cS1RDx8/SmiIdivYvx4HEZxvNAv3TyebGCkgCQlfqPHE9bdf3LKl
lPcHW04RredDf4eW0cOur10b8gDzpt8PYFlnudX09wzrJ2xGvP2R0XXOGEHBjcxksMN0m5zO+thA
nKe10DglNKop3sCFxWsi76vzRqDvPPbvBkDJUjR7qwfIW4IttpPhZTFFrpl9F7XGHc5rYDCRrBbg
NG/Jc3TqFHzweJtUIKSV6gpk7tRQ6PLsxwYkfs4znKk8xXZGo4Ulb1oq1B9/a403ZOe7BiTjrKlP
7e1sRd3K3D6KFV5KwCsBajzyG6BZmCO2k+ksSdjAnqTCUnwa2v9MVekMEaYQuNs7mWhDohAUZ9OU
ITjFTWeTuDKnJ+tN+RO/+Lo1T+yXfc1SUsu8V+sG8LO4epivAzEq/zlVUSnJh3LbaRheRiBsdHRY
cixGLbWp0zLyH/8NtGj+OYmuo7Z1UFCsZZVcUfu0mciI96wwrCV1YMvKVYEdpNE6jxBP9BDWqthj
LzLTcsJM2w7QTC6PfipscU2xHxCINCL9oqBJKP4xW+nMoOl1jNHJbld0QDBvlCqWnG3Th65Gr7nV
IfJfcDvPwAikAtNVWgUPYahpP89VDNMtTEbTp0OoBD4snBrJu/18YlchdIxQsMTg01kVF0w0qwOx
MrGGwnuAou0oBuW/81VWiflTm4wdeH6JgHoNea1+pHWp1h6jPzNRgRmgwazwPtgq7zxU707rCsiV
BjAzv11JpzoelnKPJji8srZW5COz+qYJ4Iv+YaPadSmAQOGhkcbmnMO68R+stzmbHkIJ1Khbu1dp
EZVv+GxO4s5j5szm0AScrH9mbrPy4SXqEHxU9XtyjUJWLSGkNIQ5StZShTEpsvbOTnjJUw3Hny8K
LIR2Y1PhZ9Glx1DmfbBrjlIuiw6I7CyCV9Mcd6GZQTwSSd++oLHjMYQlNzdQHZNPK0oU+dDev5Be
x3SDkv2wEPTIebYU2HF46GvkzZwxIyjdz0KUyoM+XqQq07wxbQ+kg0JqsrKarkotD5lyHw+8FSR4
gOJldjznbKp8e/kg8ST53HyH5B/VHfLANPDRO9rwXy/R63sIRdWvTzi7FHJGlIX4wY0V77Fo2BiK
ywUJhBFLPFGlLYfs/sM9djN7NVutN9ji3LXb0P3V4w1XPhgBDs26n+zqd4X4EowO31CkYIXDFicx
UolXWbF01nMJ4xHWNqXCiMCfT9wtec7OSsBfmDLVg7Uyayq7+SC0Ld4CwwdAM+UEOvfXzWlCjL2S
qXeypboqvxUVQg5d5C4787EPaYaOWQebpJi4fCQxDzzEE1ShFEzWC0q+Sl2u9kDreSK77yYwlXph
t52BUH4tw1NJwmK5Yk7pODxQfV01jduGCL2uX8gJeKio2dvFhvRzRXLoE0Ewv85YGxkLLZ007/Cm
/6u7OnptKPwzU0BZWagYYoXoaBoI9us7Sa/6ds8wcH3iNMeZ5QDvHJvhI3ZERFFfb6UCqodCiJmE
x8fN3PVUZ7ZxmcZS6/RX9qrrZgA/HdDwxKeZVHJpzq0mtN43HXrsG1Ke7N7FL7i6ju5YCMaWyZwf
0nnRA2KXDeqULqC2XjXmQbN6SEYskPtMKuV9MnVhxSadBV2N/QjPXXiw7FxlTEJVQumgofEpUM5W
1gHYX1AumiRVWAtR2wDe1KYCaGOedcqxZ2ghteDyzXtfvt7uPEvp/f/vXvptA3daGnbDuMeUVlvG
Qoul2j4ODS0tVz1pycApYvAQ1Gvz77bMW82ZhJuqDCh1jzzn6utyluorxHCO3b6DzvfldxMyfRpP
F/VJNvNjTBTBDpJGywqkCiJ476TzffS8W1+RkXhKekBHg9Og1yaXekW1Cb+HPFEpRt975RLuKys7
50w9NKf5wUU29IWx5VycX18rxecDjyr2aGnKpd432EoJH3cVwb4laFjJRKwhQPjgn1hnejix0RB0
PORgdsWXuR3BlArMFA1hyoFKdYHhhwmXy00nMonVPLzwYipqxHyeJC3iwNhB/4rSKCaTYkNc3zRc
v3nGbJLjWYetjW6U2xeg9i/upzZioZUIXdMawylEmjv/KzD5OgYklW8iHRyFZhjKil7HMLn26bNm
6Io4MshOK/jCCuOgAVsgiJ7XLiO3z/DJKoHNyIaZT+rC6R7yOos4foyBkNW5YWP8RbzsrNzd0c3P
uRc91Xd4VB7tHhjR3r9Pb2AfRJuvhR2/DHJDjYEf0mz4nR36Sba+Tfhbv3REd5K89l05XZaEk4zs
xB2xA3O6NVOAPPh0byTEzTELKuAj5BhNepiS5woqEeGT/duzvjT00IUdj2pN9rtfWCjjXf2pa/F7
aJNDXTnnqmOXVf8MPlDoAm0NADBBMAKOshwrmgZObtP9ObRRBW9vxxLlz2QpwVaxIcdK2sh86afw
3xPuUyYUxa0DemeeM7gueCZ/ISWTu6E51mB/hN4ZxbDIm9rmq+Mb6tVCfbLtd0PbOX9DCi4etK/v
MEOL3KE57Gq0OT5n55UMB1xsBvkUoP3t/7qT5Ub2kZ0eyuC2EadFyxRmnCTmwoi2jhZ5Fjs4xbI9
H2cuP51B4AP8tFKL1fEs14Efc1YDz/L71//DVwa41EtdIVkUTJFZmCz7JzYdrkr/1F7if56dS2JJ
sgMrwNyRFA2dlKPtcyWg6LO9slN2XYQwSV2MOxRBc1e5tnMm6Hu3QcAvOCRXzEVzS89d8Q4TMC1I
kr9OfE1rY5n4Aj+jGLgbWMdiMnPQ3w/PgfL1mo0iaWD5inj5DiaMoccS7YoJP7zp7KUUlJA7QFZC
cQxPd5ljkZbaaV6aJ6E0Qx2EGeh34VO115WkUBUxFLLltW6MVSzZry5tALCKiVZpsdB38lEDjlwb
DjNa/MXf8dfeb381p4zar/Fox+eiCHCoiaTzDiVt8scwSRBzlSugYymqNJyP2aclDv3iC5vPRLe4
fJ9yFOWaSDW9FiS/ixzm+FbMTacVzcZ8yZ0O+qxAHPzZL2SF5sl9Bf6pjzBC5hiSgRXwiMDv8Blr
rEW8e+6KbYLMaDNx77kGHq78PRZyKVNW3O4WcQLhy4BiDyyPrG5yXAr/ojLutCc6YpeXpdo6Y0t1
tpYdfawD29eEVxf78ZQykDYrls8VYuvXiT9vBID8qkUT9CDIRAVpHq8RKbfhY7Lmqd2QcNo8QTkM
TxAOX3NJTG+d7ABKnO2nl9XVkyaKO+6XVmuX81PZcRoKnV1Cw4Zy6v2Uxm2lE3vH3JOBLsWFfzsY
F2oeSqZxfTMlCVrFL2K5f76uoXGJAI40d+qo+uhXB1+Z0HedCT4jAKo23aruiG84dQ/EdRXbbwKU
uI9IImk+BgRibqwaDCLatQvjLEucipfePezwMWDwpY3cnhmGwY2fVyFAUe+C6QcctuWrI8szBqEI
bwhV4AOVaE5exP1/mI+B2Tp0gmtyScew6Z6R6BRIl+msrApZlhHESNXiyJ4l4PQ81DRZr0K+tfn2
Oky5/NFGKdEm9/8oft9mN8Bnc2eBJtaZ7biH+8Bk93fJVgn5UoKfzBx0fQfkE6Bpz7sruFTwMUAv
8daRGcGuSYzamrSIED8se9a4HhCMKkIkpav70uIP5eXVHlp94lk5jxZ5NbqmL/0PP5FPPQ7ROH5D
hlBq5iQHwGGSaH3q83vDcUKkSyZtxebAS7WU9BK+/FcaN2GgBEHYLguSOsiPOBSBLThdlW/HuIDA
Rfst5lSdHK7lopUG7ZmR9LGIYtltl0GtOh6MhFlaUA2KwqrUDF4RjkoKP/mskVfZeIcBru6lMULW
LekftFcs4Eis6XPoA4pBfsA0FxrkIFZ1Ot1/3NiQk0or4MOyzAJe5NaQ//+oIteEZuTz8XU8KXWe
6zxp8gObqTRIVk263Mue56HPSNKSsC0bvLdKY3zr+t2baN3fnaM8zeoyUkDd+gTciEavPeMC3uuo
vALWQJLvEE2s4LIZwoKpzh/zHaib59EqU67fZPFrN3+0vXirp0BwRb2BR10vj/KtQXcjyyoHEac+
k/FGu6HRRwAudT/rwOHIuZFU6ZA+/GUWkiDCANDXgGw+Gxg+Pg6Ditka5cu7Pu8WjxbHePV/Sy6B
knkwIxA9zQahWiGUV+9wQQ0xl1/qw7zrfDVlzTQqiKTwBtJP3SGlYPfuMB4rMJbLBDk/YnAK8Fft
TrFOHichqn/T4LgO3+Tnxok3xxZacrrfyHr/w3SCVaCQBvOcdE8RUjdiXz0Bj8RkA1j6hiK2vEoK
ow7gqbpSsrAoO5rjU7lTbSzgNQh/UpqeBV2XmcdGeN3iowhBUKXTUvmvxh+kbF8AB5Ty0KsVudYw
+1YXPJlrtwjRxqfAqAlHraz7EAb47KK+FNvJqPol0nTHgTjyaNrXxP18Jbli7nV8p3Q+Guxf3hp/
yRKaeKOdz5NCWZTusMWGgutX8EGTvKd+QAQ4FTp3odzSvap5DS11WyBu8mz6dy+xHI7y776yNbqe
LAJ3vGlp4n7gMXTzIrMYel1U6fZ5G9IdOkkhVWNZs0L4P162yVJ3N1zjWXTdjf/ROtjbtk8YPBco
rSh+sWct1Ua6Lj/smNYEE3G0FCFgBMA4O1YdVMEfgVWRCbQjyRMpX8K8HKsVzdUBWotCglneor3W
oYIgpKQyYi2r0zGOAsZBfthO2Fk/i6ZOEcs6TU3andb8ICoAIeBcrLzVPBPLNn6qw5CjUjeLZFPH
abMZEzFNr1FJYUU7+2vlzQJoUbcR3y7b9JRmzlzPqkD57PP1ho+214j01eYp9FHQnwrSTDflw+UP
/vCyrEslygZDsy25P5INpGnQOTKobXfKjxgT320mgXhfbhgLxgGyHsOcUN9s8SdZ75EBmZO0yMWN
/xUITfuUQjqsosnbz7U6nR1m4xrtCk4KVK6tqzj2FUaz5pAHx4xLl+/ShwVph8SzizYAsFHfHjDS
9iEC6rObh/XIu7j4azpEZDGn1lXOjCWVW5fXY9WCVm3w49dyCyayFMf8kAxzESWlHscO8+elSm2I
wPv5BiNVLv1QnYK8Mk1xgQi56IfajwVGsCrgOY3tr7AIXYyf0EWmbwrUeSZh+knAMbiJMZ0lCPiV
2aFW3PzRZFdBr9MxSkl472d2Bh9SBCsYgDZ1zfP6L3LkRrHaKhwXMXfqjka6TxmVWXwj6NRANv6n
75MaO5QzvuJCoPaasBNfRw4ydvf+4xHwqz6a0HbTF2e24Wd06qs2etmLi5wwWHIHoNmmMV0tGYnp
kay/T7ybJX8vgLIPUnMaJy/XTZbW6toSKQPQ4N0cJO8x8MqY/bUzqU9hbKsAANEVLc2GTpHveVEC
pEVTDEtt3oefjN/F0g3fMOL/uj5+omhtdxFJoSiSjc0LofmzzGiv+OiLxSkRabk9sqMvD1Wl3OiN
WKTVPDfGTgon61dTCMjgCVu2VO6RLm/Y5EtReO5aAxtlD+vhebLRsgu5Hr0ZA61uXK67ZGpG/9v2
YzoJst5CA6xosYm8Y6nWRmgsDZlBYvXtJnb5w+LKG2Niuuq1axtPssSY4ctIV5zF1hqHMHv3UbcS
Jr/Qd3fHbA3vIy2icWY+2RKMVnQukzFI3OVj+i3+i8iPBMD7aK9la/GF/j2wqoXCwiEGdNOFapny
N4cyLzkIZ/cniJ6kQTkPDBhDvAMt3ICD5u35VBMQ5WP9tULND8EVS2Q90lOnrcj4iyjWWloYO52F
/pVpjx9kY1eVTDVVQ2+qP/0unnlt5whspKslOemShJW1xK7iq/WrDTh1QqSiFWkUrirw6BHDoBHc
O4iBEqpCgQ7AvffoKxR45BEXxJRXBd5hGzDscIDHXmpQxZ2gOxQJ+WZ4u7XJqgcMRcp0CG7Mq0cd
CzZb0akEnyFcwfWr+u4gqES6avcjXWHCSd04DkHFePMgigv0sE6xr4kydOz85AXmQBNoRL+IwyFT
Z20SdoQYglEaA5c9tOs1lSJWLtdQPFRVhz1BoQrkgZe63X0ifuNV7z7Z2IBsvRlfhTQHnOiHbw3n
6DKnuofEGyLU4NKBsWfSWbt9LsUG27nDEQjEk+RO+pbaJUEUnPak6yX6q1vHR9xVDIUSEmJ1R35r
JJfm1oZZgXMG86O80M4hhtGL6lXcPC4uEc32jPf1q3Q4KfCLzRcWgxmI27STFmf/UWgYreATL78G
fvLaPcKhzFDzanqCDstH054tEuqxe5qbVkD0QYEpC47F3nLXXgaa8JM0biy8BNLyj/4miqWYb0O3
n3KE+yTcruKgpzmeEibWkpI6dEJqmFPAVI3nl2kzZAv0tKmhnpDKil83xq9o9uUBZzEW6awhsMuq
cg/m6XBDouVCGKfTznk5bgjiKo3p7fIeZNDgLij4e2vI4bmlMPVXwEqQEibCt19Xgx/ZMiGndcH+
IUdLntJTy489AMgjTOTg/N7NScss9YxucTFXN4fwBIyBa7N+6m9EEFaR/X6msy00Z4WOVSECH9ZF
1erAPWF6gOLQGqfRYAwxOgMhimSvTZhjc/ICSXcAkdZqSMStw04Enxz1A5t+eRgE9ONFc2JZR89N
cI4vj7ZuHbGORvTTq8iGQFtSPqqPOGUObBNwDL6HfE6XBhDEYcMe73auiYY7PhaB/DKGT5m8FlBK
IjoA+C9JLo/NGp+gpNqtpe9M89IYLWRC9bbUsXb42UPNkiZ+64dtGWLXSpJBXsFZWhhW2+ujffDs
n6uokuVCa8K+oNZRAePS3jn+Znb35cYbPR4gCk66bhXk9XOsOsv3y0a4y0UJ7f58rJosEXvbHB60
2SycGAME/39K6fcb3q9NYJjecK9cm33UoqnGOD7IFgmDkcWSBSOmcIACtGaZdLOoZZjg7bbhXohP
QD+HL0kfuJ+7uny+6sx+YpHCXpTynrHWS9oadjTo14jo7pxDmThlhMUFuSEmlF30wOc/FVHEMyqk
6b1CuluhhUs6OnsN+Uqd+J2K2KOnWtZqNX1bc4/as8PGMpim9EYfsaWq2P/9ZXQ4CPdAfAqtOWsK
wlzqwUBR8NojCXWRnBIuosgVDlVe+yPBHlbaCJ6nMHyMWVotOXfKuSerMKouIY0nTLoDCC5QGygo
nHAt/Lo4Gzavc/rPl234GheQIL+S4kTto1OIPy4LpBWYdyx+pP34/3DVZbippAsoxyGeTpwcG78F
AuUtnDSeDHOPmw2bYco0MbJV8SH6SFnXIfTXRuDg9yJt6G9ZliKHsPeFNXMWScnPUXvUH8aNlKwY
5C86MZr82SVNicyUZOcOs3RKT19ZiPj1+ZxryCaoBsBYdmSBpQEq64Q8osP+Y5CCZ4g30tQ6aYWY
7ZTXe21PhGBbU7xpesbEiQw9WepMsjBeP8F/gsEMvRY4KQwEikX6DS/FGeX/ij2y1QNIEzTCPpoV
2vw9cxKhb1XD3cq4SYeWnp8jGr2kBuX3Zvu8IIirbNESLk2WqKt+NNAHOlkUB770I6jWfi7zqwyk
KeYLUrhyrTz/NHM4+8KaD2RuK3S5CH8lauSyAK3lH76KeJwRu/LysWQW+G4bBA7j6j8PQw1SfASC
+7etwCyefFs3rcHEA2pgbhnSx6InLjj4oi1L/B0X/3XpfLAHQiReWBXfTGhWX0Iuy2y043AIM3Ep
pemCPrLxqrvdhfjqDT/bspH19MDkwwiyujCnZsewIXiOGSgBOiiRevoxTQBiwkdsmORgu8CZgrsp
uvcGW/c6+OxJ9I9hxiSdA1DBS8ApdRctSp3rrm2YA0Sf3nxGOW8JUUxQKrkKID4GBgh2b/fwAiYl
DFzYlulgExv2xsYiuO9yF/iP97tdQllkwFxVnXMcc8AH/KqCvDCZrycJ9Y8MD/nKkF9SEXm5WprF
vCcGSjY1twTip9xy3TcNzx+j7/oYMdnx7LU8QhQvPwP0pngLegZssVKBCsNO5UTTk2eCkx89+QKT
h3vAaSLi+1DLs9PUC/JJp30Jl1sJjiIwk1jhdr5BCAZv3XBqT4n8dQehF9/Y2BJX7jznyCdvCsN4
dgpwnOmcM/VxiSwGoUKvkSPKO03vR1pTW2ON+D5B8d/CyUX9TdsqJBpejXjFIUytMnTrGyADEIvI
cdSEvOdi1muvk9GikNy2ZnKrtc+sdG7ba4oiz8Wjj8uJaGiAPEmCnW5n+aUUXOn0FA5C9AddFff1
z6xtpRBm1CRdxK1fvxX2K6keotusHYnUjyCdpk2Q6HjUjcHFGlTPU6fsVAvKP0IL/zehLYW9zohN
CxkYen3Zq3wRyc1SlBJxO1YZyty6EC7h3rUh0Rn1paE4lUmldWWEuVP9r4+BAJVC/0JcmtzGufFj
zFqS43RmOAJCLaKNz4SZPB+qHYsbF+sBB4M4Ua1bMrBesWA86Bz9Vou+/axuL8iGACTut7dpqOpp
ASHgmG23HK/+CgTsgAWfPnlpb9XSNxG8Jo0gkwqh+LqrRMgqEICGUSW4qyzpeLwUJraHl3H+4BxA
gH/gQ0/mLfDYmlP8jPBjA5flwHTQazCabcfW+2IgYuUS/bLJhpix8vqL/7ggNbECSlwZ3lULRwlb
puJe6flirFxEYeF6Y+YLzu9onlQYI2f/UPuX8c+jG2i9Eoae3D35SlLX0XvPQENMnjk0LLY41g1v
rdNsYH2cTZekEltOW4sKizDg3D+6tqd1XrJPL81SrRJv+YQP0q1+3T07vGMxs2AkHte9Asju+WnU
g4qL+hPGH7dou9GxdFdusxQX/3jxrhkvj1eCVlt4rM0Eiv3y4mrHLG0cory0uRnnVwwPfW2CWkZ3
NEgalnFALmd93OJIkusRJ/iABi1FUTsaiANlxHUFqDmbSNxJM3nrJe2yN3VqZUhPgxd35zYlmpZZ
T613PcFDPRWWLICISOz8Q6GhzQIlS/TYsysRh1iePPE9P6icgAdr+Pc2Lzbsg5DXUNs+4OB5RDwn
UFZDjdlUxExzam3XJvwt48ia2dUrCwJCR5RPkTchB7lVp++5xsJMNR1avc0p0eWwKlI0tNALxNyD
FbGyeqfJm73+/wrtRdGb4DLX33+MprNUTerITf2RdlrOWIiM7birPj5/Y4OG2MZxyEhli0OD762r
fxvdsba5vnptfjnKdIrNGY9b7RGCkkj8N2ZUGhoK7T8HPVetlTFsoty90+pwDiyyWktqHPdO4Gfq
dSZ0vUcTX9BsORP3A5mYx/9jdJvzQot0UaV3g6tR8SUCks0FW7jZvkzthpkSTrxSvzfV70x4R0WW
dOjweDIRh8ZTFzmEQ2brgE2hUUGqdcnCBQmHy+bw7Np6Jk6qGXPqQIqQsdwmopIORCmdO1qhvBV5
MxK9E9/KniSHXU+Izc/oRLJu1yLDJ8N4WH0bVQZeXNAJc0f414zqp+tsqi8wGuCHzb6NW4+zUFA5
VNbEbOPsz3G2eEqBOa3knNAI70umY3FSF1I4Vqg+8teO/AItzAkflLlCiaO08IGjw4q8Ct1N7voK
Hks52MUdmbALWuCheVrI0zjL0HVcSdFjCvSzDLOABvjos3k5NLse5SQJq+D+IgrCTW1HARU8x6hq
PebjXIGaKBz4O0OUi/31XsCEPOZeR+pcrHZ6VY9EHUpQd95hoWj/6nwG2rz6QYmTtbIs3XnxgJEM
BdpGrTJsfVRbPS8W1Ze5IAEZkVoDrKV4RGKFC9jIjYcYB9jwLNynK7Fs2B3dAucqcK42RvtsEU5O
x7qG3JBR2JHunAEhm6ncAstQHSe8NY8dNcJ7bElt2AJbBY7Mqs2i/KQZ51CI/f2pUMFGs+4wQ0H2
ZO6zk23ukIl3qrC8lKX1HYnOilrJ5AGDDil2/9pVGP5plNF39UPSY4hJ8IZHKspUzqYWGZhu0/lJ
2L6mqtWDaDb4gxayeavPycFEyYmqXQ9pcOpxGY7/Zyxk168L0dIyO7PTBSjNOk7FONDzjJ6yLX4z
auNojLyv4jF1A33FfgZ2EBnaEmdsJeVqERsBuPhzRcLjSr5ScAms6VteB6jkUWRf/UGUNgSRbGib
c4L/ruqOSTHTL4usu5z682/qc6dPV4w0SiQnfAykExjF+Y70CYRaVL48p4IyL5E+MQcE5rB1R/5U
wSiASDLqqtvoVZkhvA+J+ZKFhifsYNihOL0UjfMBw7W4eAPuti331hcYS5n/jmbqMNzrJU2m6z6I
09B3DH0YN2p8mepsvAGejo3u1Zn357uAlIyDs9k1H9RCXaBll/OY3bwNHtFctKWp2XFL9/fBkdrA
lc6Xew3eVa/PyKDNhp7KOnFtHcOHg422P/p0HS8J5qKF6RcS0t9nWG5gyjHA6am1rAILvVnq/Sq5
zBJg9abyxkb5eSPEcO20qfVgTc5IkEsCxhWlA/PMyJTWM217Ete7nwpDSmd2NN0bc+gwwSm4fsxE
iTC6P0OEOZKHsWIS8AJ0HrhrlJ7yxfTNzv6rYN8g5tuDmObnCSjCeal/Rvy4n9zWGKpVanf/Ss4s
Rrpd8DoVb3gvSY7ItFoWKYPmaxH+F+c6JDQhDTwo/wZV/BvOV9o9iX9mOEcNJ6P8cdp6APGaSipf
+O8Ywnx7rrUS1XnB6D7BscRvjc/fkXmrw6dEE2TOr53N202jDSD2SFY2KDUAP68nRgnU1pc6oG0u
D0tcOGpTH145G5CPZ5aBXK0hWhZNpCuo9GYYvgAbwBpR3kkW3x9Tsr0vYYFsqj/jVug0CBiTsTLE
tz9WGaPXFZTFFPVCJeQwLDNFq4GNodGl6NWXbODvCrlXygBhDcMUKmMcJ5vKpu/RJuuHlHdeExeD
Hu4AetjsWOpg/de+uqn1A/E2dgiMWAYJiyloilJpkOAN5LNrQdgSqJeiJHy4cMN4dOYa6VN9463O
plPwI2cwvMSLfxlk9xHHnWGMcXkWpz5TNPeeco1mpt6SLG4X1EAOUn0GqhNUUQEdi0QVQX8+r4yC
7emdLMVz4a30W6DAGPyH99eq/CkOALdsCRBa5OMC4REiRISX30MDgCTtR4HZIuF0d7oMR7UAYdHD
wLxgL+ogpeV3bezLTinS3DTCggJBxWJGQEpHr91gVBcTDrdVjj/uyt0BFYiJQDvrjwP0kzGLAMyZ
dHNcdhxwXBuk6uTuANQiMZMjpupq117Y0g4MtQpimymEHHrc1jpKmKhSvLEDj/r3oIZOH7j+9aQv
LB9YR/0K+GOBf5UDMt00lRZy1UxExQGAFWgOchcwhXXmHQQ8OvMJz+ZjZDuBezRsyv60MGUIJCn+
q6HhobOvPwkK2FrAtHisiOYk0p/Cx0c86oQ01tPXt1vSbpLJPdVDSCYiSLQA0HpbazhgT3hx6Si1
9weaGymh0rIcYKDcN3LdgoUo0hZ81W/R3AjRdzDVe5xSGTzSuDAWaZI/si0UvuX94Kl2Akg+z64n
OP1b6juPvFhY99/UhacHndep39KAwisG+uK3HYr6ahqmNFPpatZKM68FrlYonDCrzvssBcjO7BYf
oSh4OSmRuzyizIgMjn1ODT1W4TV3pXJb5tDp20RWfgIdggm0SeZ2cefS0tzJPMpD7RynFnXTMBqG
w+rskveHUe4igmNVSep410beRIjfmIdxJ0N+7bvHEz4HnfSX8KuHu5GP0DiOc9rXqCnMpmF7E+Ah
4avM2pvC+UypY7asNcLD3Fmmib6fOFvkYyj94tGAy0OaZheu/O/QAVWMN13vwfM3I37TC4fjTB5g
i5BNA2e9cbQqyQ+qlU5H2Lr/luvItsM5FUs2NYX6D3nbfzvl9IaB9eIYkUL+TdgHme3+vYhHlme3
lk6gmIFn4Jgx4spvW1jzW3Af6dOdjuNydbeGvLI3oyl2R6p03m4HkI3krPtdlufrW+Eq3Yt9/bwB
7UIMVAoOzXGkujGCzvPP6Kz+44e7Fc7FgFjVZeU7zTQ9KoP6QMwhjmVQuFrkRKRgwR8L0eTLgWnB
t6Wz3SoiAMkwSI+K4sZ9JSQt0K7xWxJjVdba0foBHntV8X2UGbt94F6h6M+om6OpaKdcDgEWOdyv
9JmWeTraeFJODzd7c/EXwcExmUL6hzZSWRIJ8nfu//5QSkh8OY+iUC7Rqv9X+rin2jZYRjheesbd
Wbo8nouVffgfP3juq28DjsdACwzgpG7qZakVshVhhJfyiEPKtsVm1ziiG4JQ0tW5MvMCEz2tfaGT
vcrYSikvGHOxU5xsEXnWpxloqp+lcXFmDcP0Jx2TIYOHH4/GDTTMfkzkTuBHng0o/BCZWBJYJrWJ
07ToIiH42fEnlhUAzYv+RIrm7M8A+WJ3DWMGexQIHD0pqXEOrwk4/5mxV5H0JM3Uwnfhv46sK/6G
2U009YrUnoV4W9e8EJ2KJ62CxhteCtplo5/j+XEZ0FWscgxIvHt+Ja5Vx/nN7+lFON2s5NjfBRKm
J8mag8hRqv12B52PHgZUdthxtBYIztIKXQ6c8pfDpw+leS+Lj5TAfWFZI8Rj+QuxNrW4p21K0ETH
QptbuCos9SGdUb1BBfMYsJwg3/KgMWZoKGftjRl+BE4sLtczYgtAShTGK979+uObPV4adx81L26d
S4RElWsAZOW4COUCzABjqRxD6ZtJkiAFQJfwTVRnrmWxLhSNIjJmJRaTSuvcupyQWO7xbem4qjBk
zjSH5bkDx8c2P0Z8ciTepn8Iclh0mX9KZV/Xr9BY6skD73MbYnhoECVqWfcMLek4xQyN/BH8JtNU
jFUX6YVgluURQnZFBLc5UvQy7+qwv9OFQ1qfKGprcz3wmf9WnRA1bzVLaZ5X6TR9RZB4xKgxGw2I
HT9i1ZDpXPIxxrUe11GK3zuIBEsL3rEjYm2PdMx/LfaGtnHDS6N4hbQRRY0NNe6D1leu2giMPO/m
BugjcSmywz07zir3hqwNVqMdVDTBijsZCcxI+fdbae6bcu5WUNwLGgY62BtoSmdWdYh74pFfdd8j
c6c1DvhBBdwIpCigXIucONAdx7Aw0MK8y4mwHYDD8wYQbimhakK2VNny/86z1aCJS1t3ssZEtCSI
AbfuvBf0/R9wNAra8Eb7+FUfT6DWRe3kuN75VRTWgbJRhhfIwyMxwg3FaOoSmUuiGP6NloRrLYK2
q6GsO1QjZzAb/YWEKx00MrAkYZUxeIm/Rynoi2jKaluZaI5AHEsHe7D2hMpb9j3zntBcT40dGEWE
aWGaaxnfMNCL0v3bE83Q3M+xeZGDO/2rCXNMKFBqvMlUFAe9ZNWZlvERL2BFOYQWhHZeDjEbCXaW
tK41L9JHgjxFqNots1Lnq5UmabzvyRgsDSbz4h16FlwnjIATsvL/C4i4+l6aiHLrufTEnlJZNbFE
15wmcLPLZ0KN622Lkf9xWI2ktFCJkvwXbgl/3dDKmQffmI1GTs7yfUXuK5EyqPjOOP3D5SqTu2oF
Sk99wu0UljtRcdtefyOd2g7NNt8QxiRvHzpmCHlPagd/uB+sPDxtK+ngbLyvJasiRKyKA9sGMI2t
fR/JIPySGKeZgiznfUYf9FFcOwoXZCF+TC+o/P72I0a00jIbOPx3i1JbY3MLgWI6hrQKEBDSW1zF
Q/cQbPWhgEW8WM++6lxoB500DDLPfl7J5CJnNOY88/3PQCBpC6Tw0wzxBfqizrQcUFHMo4GMV27s
aP+0qUOf1uRJ8F7Rj1iYjk7Eo/5w6la4MKsxCNtRFwuZcz5lckwMRQS3Nh9WAsyqkkUYjhRaHZPR
sQ5I+lfVyP6YiLWqe8+x6K4z72l5x6ZET7QJM6jO/Y4eFntQf5chmknuaAU+tRv7k0vmSA4qFRPm
WOgUoiQ1BTMk5Xs1h+2mAHikAILmyxLE9XoxoNFXO06ad/lbt8S0X5phiIhKAXEo6vi15rtSViel
QugyN/7+mgLk0DdOFR7MWSvWCdI6kjJ00Wb/lSuz8ItJZP7TRidWpJM6KgpTpbRcUkuG/6hUafTd
dZA21qnupuR++Ovr8vRwhCazVz5HcKMo63X4yl9uJ/0+hBlc6J7lAIsZDBjXV7hnhTbUbOna4Vp6
82zif6H05y5/lsO0RGJQgNcEHsHgX0weooknIkVy0S6YSqVNHhUcL/XY50WwhtosoRNjebm+YLA7
gQ4B49oykeQMOzffvBa0ZGcPHxl/noRhFnfgPe/4+IQE7iKThsDUd6TfwPDOB22CRfEjWgviXdgT
64B7ORIEWCAoNiNIWS2jV98frTIz0l+V2l5IK67g/2Y5VKTl9ZzVhlDXRLKEsuSVOmgHq6jdknSl
rc3CK7hk7wOy6jZ6furgUH1nFZ3kPOJYm67PULMfjMRJMAf0pK95fBtP5bZF2pW0lkwaPIiv2ad+
Fg3lILR426BUre4tR3fHEgS4iKfO969z+uI9g1VJhEavKkzwl1HR8XRL3K2CBZCrc0IH7cyP4cc8
b0cs53Yr3y0zleQ8M8AKDvE+9hTymAcgndwkaFqv4eDZR+o8WzND9OfzDEQ6NtbeFTwIt9e5e2q/
cbbsvaW81+aEo8VMpACBr6bVUTqdAFs+7KMmDT82vo2iQr2Ag5wQsDLdNSN32lfjbb0k87kxNVsW
qf5gRJ5GIBYWf6qKQg099c9RsdXOMowZqdHW5mZhY8jyTnjZBYdf0VTtu79ma15GdNvpJrrgex4+
S48vlwn+JaugJ4/7tOlxvrOOob3VXXqyJH/Md5XuxkZa7c3LPGMTu75Uj6EjslDTIHX3+pB3aCJQ
eTYN639O1HdE3cbGg4rtcd7MOC3eUfvhwcgZqUJh6S/ldNYbXAdGRM2ExJc40OZHwDHkhiznmnIM
kfdTzIr6vrXGomVvDB0HQuR6zWWfoI7aWo9BOcD2SrZeTh7cme4DHPG8hJ89kOXlXtb03vaCuaiU
fJvi6GWnddI8lqpAvg2YR21lxkN+CEDSSvWiYvbhGTU9zFZF93OPQJBPMVIr8/3Bm0ANqs7v8MnL
lUjV14MDNJIPN3h6sHhD+Da5ryuz7StskamHiPEIsyXDaKbRLCb+BVmLlrKMSjyZuLye5Vi9p+PX
jfTN0s+Nx2nM7vVb26bPxIsZ9By8PsEbBWW/sEVoP/PvB8einmLzYXZXq6Le5Oz0VJDyMEbk1eN6
P2k/tLkaTV7cv2Ze2ei4VZYNdyx7iGabvLd6yDIe+nDFyzqSzWvr85zq+K5z5jmJpJCA9SdL1pJo
3iU66XK9p/cAehTSsu+YoGkyO0zRtZflSWpLtI9ETu+75IP6lAiWf5GkJt+WkF3iAkNtWIAOspFu
qOHa83qvRmQK1khQV4IH/vAIv6pOFk25gJduqLo/rdVU+PMWhwOsFJdJgVfposs7WDRs66JY+JxS
ILaaYZeny/pXIXwZtZzyBlHVKj00gsPvp5580F64C5owMLH6QRqCTbE3QYGU8MpxkB9vumuVS+gP
64BI9x377vdnq2JL7f09BNKdn+M0TRmrp/JfapkGuEbJBl+QV0FIWCuMOPuId0y8gnTjbJPNx6i4
aANrRD8VE1V5vAmh4IZSezuA6zQd7+I+Yy9B/Z8saAvTuVCe96kYBOdWa0jhq2QaMT9RnQyd6jsO
wqPua+NVgssvId7Cu+W6QMBAHUhRibVRWThmW7yftfRAHcZEcb4jC/rkINnv7xV6L6X2dlxG5ya8
b+BuuOuHQB0m8rhZa1WXd/6DSysHFonpjVLmPLM1ojrlzRZ2/3NDfhFpIQUFMfjY5iETvPLgKJeu
nsTzhjZHYnPJx3652EJcaje5wBvMN6erkBLOJgLP1eviCxnxC7kGCxpOs3ehV+yppwSymw4jplLs
IAF/w4dpAXnVm2u+sspZPk9HJbClaFoLxZdlJEAvIfrul5Gby35tmmiNaFeOHtVHWCnaHkC7O6rn
XgIaRStuOcGRQA6OufeAmNttP5FTrM4MhHdrwvZHm90t/jRSlo0E1nCOumMJILUBF/fafvhC3Upk
mKRZydLiDADDHjgovPtZPvBmbIPZcNYw7VLzc2OAAdWlTmLT2iptpHjIY7QLLAdLv7cxqyJN4JLZ
iE2SaxUlwU+YrpkMdXsNfGMomAamFiKtvLf6wVfv/9dtHIyRiAz7N0Jd/VcBmwKYH50HmaqFkdLP
TKuLhiMo2iI8muB8+Xcbhf3zZJD9hR3EAq7zP/cRMWZoF12XvcKZO+hWlge8Y0Wv7osXGuBxTCFk
AoyP4pIHHZjVBrixVKNCE0o/eIxG+Nyj070aJoTImx5XhO8Q8zSOmU2KjgE8IkkU0AvYvfHY1bxO
frudYHAB/680fcusStzQUYQetxwwvEfaa2NflJ8TrNmndGLJh9ou4w6dSuajPCLXDXYI2e037ryA
iQ6puWUdAzUF9diEVJ9vxdfTM2DxSraHjUjzQP+HExla90xxRYMcZ15cvCGMjIC+rs2TYKD+eA8M
CzP4qVHjf8orShR679FTlLGxL+TrZPl/dhbJJBtfDm2/pd0zMQAHgGP0JUY8cbmvfCTO3k7FZH6J
ZJoFy58SYUKDh7buSJmT/N1QY+959+vttE8maEUK2548AG/i0Pb4oxIu4xmT1LZf8vYW5orkMqUe
BsY5CDDsG69MJ/sSJ7tmIlW/Hv4tFW3XQutivs1I5qnKJOxB+Eoc3jfiyrCZ9pxb2qFtJdaTjl+A
PLylxqZWLehxIAMvTN8uzeYqoMv4sxJsVydpGJaJ1FteM7I26NrvIHvnuH5YS3L42SOpK74AnIBh
W7vlwKx3uiJeG3MTyvJos26Ba/SSsM3cZusqGqBHRDMs28LQGLVdGMaZcKRbtALz4Nkby0HrHRJ1
A4RSSC1bV2Xth8cGvZCa2r223+MBi8KVpJ1lu7tKjKqkB1tIMGvM458WdT2iK8IKZXiGLEj8NAXl
5QbK5JwYJCJGU5GSQ6/WUTqlvbmYEtKbNEjzfUfA94SpSp8SYBQpeJd+a6cRDrr/5Eafnb9lukng
78MbqQgEqOSlSJ1FhNx3oTo4aF5QT7yJBO+g9uFvAwuhxLY/x3iQ1ojlJrF6HnmaErXEtXv2pvjA
pDcz/VwdCC0d7XMl1Y7LPAGybPhVjb7WdZ5hgjILBhG3ddZvTQJsPtSWxnQ3lQ0Z7TNDeG90KrDo
6QdwjzLwAnWVaJqIY0WjcvlaiNxTfMKFhq39+A9Jm3ipfN5UB7e5Iy8dpxVDlvwWRlWjT5QHVlfu
zxKFjcOAe6zxjVDTIi+xKLvLXg8pzuSa+yVRocf2nAloxHxwtiAqsdWKKTz+sX5dRyYquPaiVqpU
7VpaM0/hRyvxivCvIoNYD2BglegHkDbPCcFD6qntLRJsJKJllxScCPVM3ChcGBIivEYoj1EVdcZi
nImnHULfVKt2J+ixbUcMVEzdDaoupDH/LvW3Dsli4BQySCaNNpOYlGj2l3f1fAL2oLmOLybOClVa
+1VUcUph02FQTuAmIFZKAQVLYZPhQNeMN8lGmcg3o5WhiLT+4SVhVl2uZmsKp+irsEJEEGXc3Wsx
GcziCy5CFR3nKdv709tkJGzLZlgHssjNYo+LJJb1x00JBMrBYjr4kQ/+4m4vhtt/R3mKaJzNy2oL
BZaBDzm0vKaQiLZ0/Oy85lYxC/s2LM5e9tkada555sCfFeSN4ajllWpEeF/qov532qaEyBe0FRb9
ZolDrcArWVunU4jb3xHmPzNXwD1PpEMLeO1Etsg0UDEnFty6DymelTJ1xv/J0sfUmL5Qk6+mxSIM
ib5FJZ7+ewdNv0pK5lonkzAolQIUPXRXPMxVhzCAR6eN1YLzPSjuUdEjvnUP+vGpZpxvw+VgOd05
abf9rlRrE65V8BYK4IRQjGz96ABb0FW0OrwjjCiSIDz1ehWDKIX08hZUamGUFRCaWKma2orPRM6L
wL7fPzREirrQAtFU+zlgVDWyPQFMMqezkw+AlM2Dl76fIRIHqjAmtQnTTh/oo5dJw3+eJbiwKtj0
O6cxJ6LP/dDErW0c+Ada4HAFzRPjRAMNjxAuINnHn64vMaxigjVabT6FK/wgSgJpRKbbFSrFWhPl
iZTDb+7+mDdlR+qVucs66QkYTE5/4D3kHoJqtsHwtyv3no/gG4852q65j73Ijn9AbGa2FBBLOq0d
Jef2e1fXs8SAr5N0Ol1Er2apXN0fqk2zzx6tKPH85L7d2pj5AkpgK2o8Rj1YYMPjw4zJOShVWR3L
cBfF2AIW4eKDomCHQ4Jijx6/YkM8nAjsDhA+BU+n2Pr48zJyY2yCAEl99ir7Ct08K5XACnUHcq7b
/kbhnJvU7i02QmCXObcdAOPubMqlhIpVmIZd9pZv692nRRQOCZAaZ0duZPbSAy4l2K5hSl3RrItH
Wt9V2hUQADtWNkULkWtCzHQITREJ9MHZYeP8WOacWJh3koAyfLOjlnZLd7phJhyDL4CPwnu544/H
xOy7WRPRMoo8150RM77csIp9Jf+Wa0afmZF+pL1n43Q0OMe8SvENeJpIcUYoK9naxYFWQif6FmLp
drwHrAh1yc6jfCNK4YPBsr8YuNAI6V7KjeMNCeP/H+wgGpVm9B+NZtGPe0rziAVqq3vk9N6NhzYA
jRWQB3JAHI9rKdhFoOhGWwBCyNjLaU0lIMAwdNlukbxCoCDF4kWy1wO9m2RgJdnRD+KFLxk7NKf0
LxphnEwO+0ZAZAJUFq9XdTMijWH7uKbsxZaSSNf44wDkzCqUPIyDSUx78B+ATE+NFsYh21fWhpuK
DqR9WY1Ja3cmU8PhWeOJgSo8KWnwJwstEhzeRKw/f+fd6SnQxyqQnS9zBnEQm4eICA/pd7Q/QKHY
hTPD0OARj7bWW3HNng0GRIEHmeEEXCr6cCGguxnZTOgv0sAnIi7mmX4Y5vU9RY1mPG4y7xEul1e2
MmzrixXREtEcTW5YjMArGaRyj51OpdUJEhmN7ya5B+x/Qvsx77+Ys91mSGV6Vu1fErOKwtNFGPQV
nwgcpeNKsqNRIkTvNXgltNYwC8UJqSOo6kLWvptEOR+wY5Rarooas5CrzX3ZKzgOX1owW/g25pVR
JV9dI2ugI3OKNwRNrhmm/Z6oKS3jGc1MHCgdqJNlsQr0XdZ5IhI5VvpAwnQNrgbSDKJeNrnblW9w
Tr5Am7+Pwk4syEZ6fi7D9+xxW+jHuxYEDxEo3CfRvps6lUxOD4GpZ/fbNzS51k+ZOgleFu1wWT/z
KAQvvK9/Zo0NqAt2b3pBXZCNu5OT36s2FrjL26YZrFlNeGk+zKj+L70lDqrFhH75+mcpv4HkKDUW
KgKgE/Z8FpBMsd8vcAqDTc5M91G0rK4M44/z85CbqtdVPPlJoymML/jbz7Oq6jQIfH73q/00XKaO
oeIh5X8XmrBc7wCYlMeuuaOQbeh8sX7DInaJcBQQOMDhFddyfZMS+y+jkGt5xuoWBnaA/R1LL2Yb
nbE4KsZbdtApff4DLrKJRJC8Lk2Rh6hSR0YB0WrVi3nXZNEvhqq5+g9OKCp+V6SPNfO6GzqTFvXo
CqggNtNf2Go9GPoFWnam7ZwBChTV+ZnkasRtucrUI5BPO6drDYYfGtg68po5clDayZu5f5Rlf1pu
IZxNWWeM2kok6Pezc5/IUEz5SgfrsFNcF39yLsRf8ah6pZVkHIQ1Wlh1hAyuI7NgU1MDJ9DD5GUP
JbhIlJYfMaWPMQxFZWjjVp9wb8zbn/Zfjn2IZz8+tvDQrDo6wuZ8sYbTdAuA3lCyIy8vonQPhXIs
iSj1nT1wmi0oE0Pjw4DQ6hKl/6p/bWfrMIyBur7tGV7rCxb3gool+icd0qwSY9XQIfA7tva4ifC8
Qf21OgXBmbx9sgJJNPC1pZCxSgP/PmqgvzFGjTLj7qDLSvSXR7CsbgOQnH9LyyKeXwsdixGrcR3x
/Uypgqo5AnkatdT8Gpv8+ly5NgngXwcAxj5AM7myXejAClmdoBfJptw2HCvzgbSNtdRgGSkN9+Gg
UmRNlsO/0SI5qrdAl4NxeCA32i8cEC485OAqlOShA2zjQL52pKc13Vi31oplsNINz38VSzSTZDv8
J6bysqOO3zl79YUuW6P5p2c7sR+EkovQjviHIwv/pV/UgJJm2xfv6TWbfmzpOYGDSIoZe7cqeOyQ
8KM5m8Q//F05qKzIf8eYKcxxiavWsNNW/t1IeKAA+Rz5+siUWUosDvz7N+9QLXbTXlYpEVqU9Gzq
4Iplhg8yv6zhPed5mpynF1ps/t21p9AE6HwBGS1TUEjSAENCIbHott+sB3UmOPgK0AEdAm3AFfei
XPohu85ws5VnLQr6I7dLKXqDDhZI/mjirzUvNbkzkcb1BfxtW6iH6WCfxoYZn/GN+eK6iDkbYXM5
jJy/RG/JMTQapf3Wi8Tlqc28cIiGPJIzzvXrnTxgSJcZUmiG/FqlwUFti01927FEaf/b72vyshHo
B0j2tS1wbptw6DY/6rg9TuTT/21u7aNIvU1BuaU4h8Qcz+wBBAiUQh5Y6iWv6WcvYB20l2hHE3Hc
rUsOM/hz+ca6OlZsLwmrwcq+7XlwkmCtdohnQUoY0VYiBUxLkKAACosYO7+lTQmKzYb7NRuMVvK+
XP4rGnM5xSLB/0FMcOV/81Hs8EFvO7w1QNZHelt4zFCq4zzHP98VHPTGX/f5N4XTKK8ZmIOM3hiH
zRbxfZywCojQI9lPwMJ/ly5nMA9CZ5O0iAes4su1sep7qd0Sm8CWVJwrhNh7YK9XPh/4whXs+BY/
KO5PqZt5zkJU9bPv7KpGwxXSrvLxIy4S6zE/WNvdVmT3F8p+shZpCPR56XbzsubCuTL0UvezpEXZ
3JJQ3MV8jGgVJAcaheMEShNQ8OQpyCzjUU+FAmDBrmm14MIXusHU0yWLOVHU3quc+wW7lsEsDl2G
GlYxoscGeetJuS7L3XjjHMHJlQ6gibttmWyWHgGdyVLwgzIblfVxSXAFflLVpu1IdQLsMtuZZBI9
03VqD4LKQnqo3K/WNzZ0rps9StHeCQZyxRZnQ2EXNOKpy6YRXQYIY8DHsoeTa1v2ys0oaEEYqhja
LEKBZyI4hFmVqz4onv9KF7bO0BVuxqy8q5e9++LKFCuH7p/0v1Z0Jzlkft9FyqMgVaYZf2LeTwea
GsGePmUfbiv+TPEWKgiLW6U3EFlrY5OChuV8VGs+Ewd1l6zHvnuJ/r8nPZlhzbt6QNnr6waj/XKT
/vme/m8/BPpwaSH544YlaPNzTXNlkJ3gejitfkg8bUZ2fdbzBd62qfiExyWIhTurcR4+BToVU66O
xG+CyGV5S93UwyEBAJLepo46Z33MbIsDE8hhk1j0JdVfwF+UYtHXUXn+NYGUvyGerQ7oxizvhxc6
M0g8TTQXPH35UrAD/lkjPIDQyoco7pJiyG73Z/lUb8kw6alC8YAWPSUQCTdN5hcbVXaU16NughFm
n4wkEu62Bo5yfOFqS5469S+cX+QvU0Ptk2yH+dSoff+1aLh5qC4XjD2J7KFoebZCRqdQ6uMCGJC1
HqhSq1WhGzEzRFUCA0rdqYWCoRuCfzrUR+77ppSCbuo0BuVQEV9NwMQvGnX0BC5Ja2IdKcFqwS69
X0hGF58vEGrr01fofHoRhfU+UrZ849OVJGB7+Zhw/nWgzAQ/psaDHVuQienWisZD0Xs4+f9V7Cvu
JmT9AJdiEPRFQDCoxpKdFKE/0z3roQo5twGqGE4GGRjS8zEM7v8NPLfG6SKa4gtTkJ1GWNeykcmM
dWz4v2H8vlNUHMBGOmAQLKFIk3ctnn6z0ofD8DzzA3Wo7gwDDq9o3oGbMQ7jWLm2xmvETWXXXa66
XBsMTZDefddDjME5FnOJ5vFuokYhmQWbkN6NXj1JlDP17VPeRNrbJHJYg4wGCmJXyTg/SZZMU143
d9cxZH0HoJJs24aj2cyX20t8VnoHLUewBaxaOLM5OufoEOsqiCJsgIfJLuP+Bpz8y1/nDIXs31b9
V3leSnSSRhYCStIAXCOsVWtzQb9jNVr05Qx3we/h1ZWa/bsY8vc1GpJBv+zSSTDTiyw6GoqLpvZp
lSwFMldz6IX1KyokJ1rTo/77LfSkwATdXnHDqxDvtGtiqrbdO+LsV0RzyLfpUyqSOvhBdqOt92Hv
CiH4O/cooUn+e2gxh2y2CDZXmEY35rpDgB74eqAdUtvjUtXJy0EuK6D186rs80S6DFWB0RFuUVAN
pEm3HZpkOyi2KuhuXknir2emUczSgol/+7f+Dpsb2Rnr0yIwgmd5h9N8bKCkB2G4J6/XrzVW/6aW
RFWvZA/Nb4G6PatsMXNi5UExqqAlQQxWcDL4Z1a53fL/gnV5fUluQLecB2D7DKy8WnUiRq6SUzi/
PMDQQB+Ac2v7L6lgvWaYP1kAO9rBn+RCgityKHE9teMjq/bK2tt3snZcpXri/VXf0v7B5knb9kER
jFSPQGTHvLb9i44dihrh5iZ8bCZSr6uQVJ8KIN5CvbDoJPm4sdm8jOprz5N00V7vzZFEBfXNuxPm
iHfqq30nC9TeSiBI5XBFnnupRk2JCrcNeQL+fR/UMu505XOUHmPcpQ6kJ5fDMJaTJypbsIEuPlSY
tOt+q4lj4vSk7zrbsueEpM0K9FCDgsMJznXHEdKGYJvmNH43+ID35SvycVOk4LQqS6lFd9/venI6
mNznQaIpEVE+aTOaoOOAhYxiEoI8as3QVr7VgKfkpoSiHfFn4xKUvWABMuD3a76YRMCSIGgwHYn6
dOCjU7HDBNHbmf+F0hkbQ+u3hW/CHt/NGl4Q3BOW1g894ursWJq+iBAf6o4soUvYIALzqVfOQPLq
Bg69NO4dwTIarcz4mxprfO7YBjvWb2T3rPFIUSgv9aHURDeA3/knBAVcw9FkTtO5n0mnHCvpFF9a
7W3Zpwf417PzsUH/difkXhkzWvsDHQG4lnlxI14aEDvY8qMA0yU8kZqeGWdZHj+KTWnCmmRm514Y
eQTvG0GvRafSlFJzWXA6Mkv7znai3B4ydoA6FqBsS+LznLIzVpCNNQfHjCezfBuNnRpRuMd0Sr5V
5BA0CVLjPzsb+/6h4QoT/gM1MMLqS7aL0FUWgtZDnH2J644RiPjPGV1BzgOpLJv2TpNEGz0XMLdZ
Rz/BDOMwZQqeFMSbazcm4iOazFyPUBUL7I886dtFCdJVGm8HNo4hWr1d0NU5G+nxcdzQDzCYEuLl
gPwfgHmUeZIO1B1cxaIhLAWAkMJ6U3enz38/zznCYA4YsoxEwXebWitBZA9+zsTyRDJdYC43FTsJ
clyvGNn8HYaHoCrMrYJl6Td21/y1tHHhZQjNem5s30G9uQNfGZtPlg3tNCOGR13U27jZPbYN6U3h
d07TtCglmnz8THAHzEU7hgf61+HjKm928pE+QB/HHTwbL/rF45M+ujEElmjvlFnF0HM+mSYheWDO
tF/vcq7kMrFmS3pRaqgnBAdfXpVtgx+LvifDddbmkEVcBndd+koScEI+DtsqlBxC+dfmqzPdIB3I
nCHQKCia70voOD3YIy6i3SnrLOmL9sl5pMnilQ7cwZlSVgNa8gd0cneGvHq1GOxvMMNBeAKDt2+C
JwO4LMLriS1xIwytlalk9jhbDXU1mBRICypGEpttx0fnA6lTyK0Bwdjltl/iAsjAFw6IU+7eWstp
UKSlfxdlBzHkcyaxN+N+G+K1yhtJkBdhV4zf6TYwEd9uIiA7+k4Mbbz/O598qZwK37XZIIKqzqnw
v6nO6n474Cio4VuegFCAoK9oBcUE7GFlqcoXlsoR7UmopULt51BUwDPoYEvZ2hM4oIEG/EpurX69
pre5YZICgYF8FLeyYHC9YBYxnSRRe41mqjR94TstpYrtnbhvYCjoRhWdK4oNMug19SKArTXkhNAV
azzHBhFYDvqxAHaHrFryR8ZtbWB5tJ2BBy7ERFsgfjs1wK/mhZ3PrCLlrYi7JmGTDjnfixwkaV0G
321LoMgDm/6l9uomd+4mXIj2NATlcJMLu/9GEdsrpJBh0xJo5xTAa9txruedw7K/n6Iec/3AppvK
VQ7MWjj2Q71OTEY8rs/aNWYUVCkhtc7wZJ4Zop+oFz1lZ5auPyDqnpF7FEH605+UibsY+URMLOpm
t4zuTsd03C9IW2okWbqE7WcTCNJE2ukaFDo2lkE4ApqadT0WS6SHGY1uQlhAZ9Xkf7haKpf6OXaf
5YGW+GIELPWx/VpbZLabmERsDCXV2+g6KRGVLs9TzM0DYRFtQZidK8Yu+6LswBZOAqrg5pSnFoSI
bFM8cO6SncanfwKndNUupazBF4/rpdWXLnpKpSxt/iJHYwoSKCVq+NvuPgzlw7Fm5rLin7buFLQo
1wFN4HPlxjpNTvFU2fKScRDLJV3NZXWihzLxVAn97tQ4Nb0aci0dMkc0DgBmHB6DDiPTQuWUobjc
J86L2H3abiPUtnGCDeICIqrESU6lT2Fc4y/NCb4grH3Up8FqL0fCOps9uzutBR64X323OrypI/hj
Xva41sBTGyul9Tn8TjrWJroBOVbShc6lC3Yw3Ni57k6wRm6U6cySr1c3HefH4Xc/ZY7H55X8aPf2
6PYeoFmbCjaN9b9BjiiHjxt4PvB3T2Z+cZW/8Xg6WGM5AAqGYQwjUzHXOhwcZHYkT4gNNdK46SUP
elNl0zlxuLF1VWPxN6AOHdLD0XbUubFt1jPPRc2kCjFWuA4v4hLvtjxIhugpkNF6Tci1EaPN+gKu
gWfsNoxQFn/NOhPuEVYysRHNyRvXWcAaKJr4KygjofUTLb3Mb/HQGbXcOGOnRTsoUrNP61MSO9Un
iiOMrazXCGNmzm1SWW48ePAZDOxklUY/zF2zmtHBlszFZr/O/OtaCGaXppMZQa8qDPL1ccQaeQB/
ineuO84FctnEO0SkG9O7GV+vJv5d73CRhAwEMyzz2moj6yb0WR6apGRp+NhFhA6oaxhBVpNtGWCY
mZfVTtD7A2V7S/0WuBGepji2SgMdwMBUGeeMYukAJ9lg5vFkzMdFQTgMoLUpR4tElru/NF1F02dz
mlnYwV6+VrZBFQ7kjdo2LC4FA8poqzj019rG1K21AR8CZOAuX8UW0UceTcUoZSSF8EeW11q03yM5
A2NUinuQbpCBhqOSAetYhRrpcC+kTQUQSsgnp/A8H0m8tts0teIujm4wQA6TA9C216EVjt+sB194
7m2h7XwJdOseYMzFAgmZlQJH7nxH0hZiKxCYwWABvj7ZgvNIcq07VVzrob6MlpdsTfnX1uUvqgdB
Rw8HrJOUsJY/BeIHG28TOuJX5p5IeLIEhqhd0v0D7Rg5NFaatgUvgOTicYLfm97Mh+IoLUG1qk1A
t/1N0RZpGgMu0CTBneBb9+LIVw1t6vvaZ63wcwnHUHgGbQ+ACsWCxidcm+y0RwIUbGs/xPUg6aoG
7d1qHfdNYt984Sz+PAQzVDL9FF8sHuW6d/Zt1Q9MO9jxm7eLPxEdcH2DYkY4zx6azZokCWevksBF
2eO8eDfWpt3GM8TIUZuIrErlzsZJFzwv2zhbiRQK3cVtmpx4n6a1GYK2tDbwkyd96McShajuzQWs
UeKvUc4xH2VjLHdHsFgzJJFi7bqZqGuJb3wmD440xhiDguf08ZLA7u7yneviuaZv3pvRNkeNBs6P
5AFdR83BXvhhzGxNDlaMXYhPCqtlTlie5ECvpm4PvDWcwPyc5q0JsYIj9uO9/KCP8BBDEWIkISHA
46mJeRD+Jfvh26GUDEPD8/D/DwGByz8nqzigl1i9YwgHXgG5CC+bVVO3ImauccGABzVBuJqN0Sjs
agrmvMbsJxzokrSAl/k4842USrs3uHCZQ6mKcMb0RhvZynPzWbOPFn1j5dBB5OCAHqvm+Pbzx978
ypr1VXhUZnzZ7HvxvRRdYeI2zBEADogCXhOgQ3jz+U3TsI1QZgssaDTSs9S4EFEIlNYW+2Vb6EBn
5iUkG93SvrBkPszOL6i1DS0qRSXP6TrIEHYs3IZQyaAl1SFVot+HTcTPW1wd0AaBoIfJ7R5zWrzB
Vq09tO6OZBcGCQzIGyWu6BZcI7c3xcvH5u355ux9YPLWF/plPpZJNIOVuWKZ5dVg7Thtc19xUXcx
bPXv2Yf0aihqx3BayBWs8EALua4wOndbWjPNg52tDQ17JsxsrQ9D6r9mgceBqEdxwgMhpE9AFBNB
LgsNkShy8FIk8CjQ4jUJCZCxXRDBkWoDChe1ka7NLUe2pPKdah0xCQHRuSINJhFwDSdOPo3c5i5n
ezMiI7kpG1DBtnF8HP6k5nixDKuJpTc3I64jSocySfgC4u752dK5AG/Yn/6iA2OBGMCGpq/c47DU
7imQUTkiFdVC7Rb6ARlPXaFBNyPo85t9pDZcS2re0m8s4rQHrS9F6jPJxaH4xw0eGxWCjk9AmWS9
5AvIryWhaReb/kdP7C0cm4qFERcs6C9tpbTvWzMgqkLTeOsrI9HhrNp8QLPLZRvHDXp0/2LWmpC2
cvsDZGj8Sgq89TjqElbdheNAPjuOiwglvt+pQR57yAiAmqczncFW9oTm0UN2fC6MhcQ6dYk+maa9
2hrXz+w0b2UQchA4iX2QPs25hbhPm59oO5oKBlw0xEAHKOtiauHb7WkRoNzxDpwtJnGYFfGgQzuo
Ad2+obgy/rSjszKSEg9R/9B3r6IcNW40wEUHrtw6IBZoQAcf9U3cz1iNStvqam8e52czRhkqvLDY
ijWR6gSL3YeisdFbwdR3xZ0VCNoRkoAnu3qk5DrLuRhq7w6UfW5fzMaEdNyVYZrb+Ae62qU/Fwlz
eS/9eJ1MF4E/Sr4c7gPiKzAry6pQDLPC48xH680d5xPWUPyrRrBbgB1eCoSOWVro0n3OQhwIKJXv
XUjh9pi2AorfWvmpRNIUqX1xJZobPNHLaeBbjEV+38KTjYxliMcUhTYZzQQPxTsx+AxoJTDxT5Yc
4N4G/vRXqXSalhUcRX9IBXeSuY9iDQuS3L50OWG2z8m+SeR5a13TauuJp859o0g1x7FN+x8aZVg6
r/O16/8jxqWjZuNCf64UFtMCwEiqnWg9YEENkVxVUsnMdKP1WwpXJsG2Wu16z8PwE959QAJcYC1Z
IPWLwvFGPPPLblBgPtS+dWECEYMBP83PBsr0HJKxwgzNQW2/rKjbe2+Zxg2hZR0sxSyadyGR5GDB
v+Dj0wp27jDGgyTww8lTo7EUf6pcfeoaRgEkrQL2YAjvmvCmNKDBM+R5/jCzwYNexaDuJdp1DOFX
19K15nvtc8lrZcErxd9V3pz+Mp/NIu/ziiWsrqJ65ppNweCdbKqR8JV0Na/ADEf3WvDdzbRKQnzl
d7Wr7wky6Xa/nzGov/gAuhB8+SFvLenfn80K5sR3OTQAtvhOhAaT9ED60fwApktTlo1EFCI7yhUY
9kmDbIPiuTHHxusX8Xir05Mtb1CbiDat01bDqk0/K+jHZnPiUMHHhCCl54n76Ty6UWOH1DiyRGBA
IbtG6kiwrwSql83dDAeDFJ6VocgpBXE/qOyWuw3M2zmOwKXT0CCJJt3IemRAxlp1wzsPZMGBQ/bh
4PLQS0tKVPefyrVjSdLta683EHQOus6JKhNIbDYNJ9F/22+qB9GRA+J28102SQHyFBwy2XzpOzaQ
0j6oHoe5OiyRhBemtIRBDlR6m9Rd/ZsOvPrjeNKSCpNp0s8xG82/Xcg3kdBeBQ2VDtYTRDMMWz2M
Wcsd+iLRU+pOHsMAFf3VDIPgAoELocSjqSZAvIVtr4PvhKCGJmnGLAuYvQc/BpeDR1dtLRlfAZhJ
MzPF4RFDOLOolejuFNGcV+2oKREfQwoXCwFtO1duBYaaaXLIZQSu8PFFnePxntdNiKBLxRujKVOm
el6coEBMwOAqkmTd1QtVTkLJ7W5FOh083vBS/uz1/1Tsj2tpuvqqG8cN+6DFu3M/f3eRN7pjZ4kN
XhHj6ZLG8lUSNmg30l8J3FlIUOu2W5pNw6Wih5hQ0hhGyfiJ25x1APlM81kwrDrd0COmXZHgDGsn
vBKBbLJQ9SmR/6JsqBfRuRxyGJcWmkV7uZ98y1yY5gKgZr0T5j6yUeugz11dFJMsmHU2JHCqUebA
SNqO8Em+Srd9ju/DQ9S/4Eo5Fol9D6LJmpeSRPez124ApUgbTGhOuA4WCyf/Yq92zf7n3n7GPjPZ
VQ7LZX7N/Bg22DUxQLxn8PpREP1fx5pRZggTYJVTI9jmbpkaNKP6n/Ixax+IF6TK/DB7rMA/XyAp
cdd3tRyNkYZhZDrXNwUJg0fTTWfeT1LkS4oH658qXgBXdEht1IFD5YR4pXt8rM14LAXTa6b1o3q6
6B7xXemrYXfMcgvKGY4/M/18BDbDN8wgRi3atqtWfz02cgf9QIaV5ZhfxGQIZEkuT2A0qq7e73Dl
Y7gd2b1BO+F+hXO70WyviycPSOs7b2YIGY5AhXgD7A1GEyJOdsB2WLKl+nCPFAEiWp060iXMVl61
kF9GSyoAajSV+IXMEYo5EZOQ1JWyQ26uICS6c2JhCiLi+FUwU9/Y16vO4izNv3sz5hvX32ZNFKVT
UfHde059pnprHsx4YIEXCfHcw5f450oDFc17sBtKmzRNNyeO1DFFaNB0p0BChHNz8ywYjgpC8pbp
gGgmjbUlTHybBLYgB/BObkaK3ZdpCoBYaf1wQhosWcdA14vyuI0q9iFpIrvBKF173oOJfnzUIQGZ
LtsyGXj95mnBFO4/QB+HV9MAiDNghHd+XqPD9MybdanwG1hFEBMi6Zyxv5A2WUVIS/zjhhWBrS2P
2jdJr0m96y9x7Qo/qIvLiZitehf61ge3LW9sEh9g5LAKkLCfchhwEtymboL6nuNgY5ljhnc8eKtS
GseYsolZso9LoypYISNJifl6g6QaSKlTBKFQ/I2MxK3ThkWQjdRUVBiJcYsuk20nbJWcZdvIrxlt
FZS2aBO8G9r+eVXnbgOyhPvEVjxHGd8Y8CBrZ59awqFeioLYqv+HsuUKdgus2R9NQgtC4UbOySqB
xbHsM31CEPx1VWbfJGRZIF9+gD9mldloTHPVD4ueRoJumGbxm3FO3+LPt4/TUOhHhIIintk6xWy0
SX9L4Tp311ShIZtbuGQPgMyqX/QgGUoeEtXYvDU/4Jnjpg+jWEP7iFgE1PpxxCKjSkm7RSk2601t
tpltq4OobxKAXeOpzj/sHbI0bwLpj9KdQ+oi8SjSfIfG9TINYN8bPCgupk9Inco5H6giKiJkv0TY
6o2W+ZjycrooFhqjInTVDEV5p38Xj82x8N9EPmczu90Dq+QAR9eu/6QYQDqNWoSjjdDmVU9gvq3t
9tGdfgl/0t0lRTfgernanSKjhdBYuRIVrl+D1DkakEnfMziUrDhhQs3IJRajSlbrtcCaGxMmEB1r
OD0L6Sep76fXbVPTxFfYcfOSs/lLbxIIq0McvLZHXRVFX4qsvZcv3Ia1GI5iVlnMG3pwoWGX4QOB
zjDDscvrBi2dLVB1h8uEL0lhtGv1z2itOA/fCdWXf3XtV5Bl0WMIy6ulKrnOC1z1cWUm/fQF2NBp
UFPYKXQrgNLN44lzoDWJiariYXgfA0Y+IEWsRQUpHdLKSrUyAEfaiE6BBaSbw947neo8XBstylS1
Z/gsqmKttaOpJjhUJtlipd1+pmUUBah7SufmHOjy4I9aAzrtikW78Z7s3dYbUvc8pLltvv8jV20X
0k88lm42BtMjSP6teoTucsDQ7iX1mCHA5/CrK9V5Sr2k65E2EvRJUvmjhLhkNDacHoTwmcohMh0z
KEk7Fk8ob0zt6FoHNq3TrfN8hjj4b+oD/zwG0J/1Orr1Ki9jGX513O66ZX0i9x3zzKypCsPnPuqC
YCAHyWLsEd0jhBcf/xCb7zZjUjkwMC8cmUrtQOrZSbvEeo7ec8Bg4qm/Z3Lt4/m69UDXJJOuqffz
FLiWXc97LKcmrSRbvtRDf/LVIh34wXeFF2YY2ryQCxQYeF4aSGMbf3yb4W7rZ8AYLDjr4MYZlYxB
f5v/ovL+kE8mnBWhHO5qHpLaqbBT+1wL/0jvuh1D8v/FOp3C1kGD+X0Wo+Je0aEnrzIJ1VfDDO0t
ohG82D+tLAnWUSOsXr4zSwMWf3ujpnpXNgzR+zkF3sFu+Gnw7nrCjMneQSfKPeh8pQsozT6MFNH4
5ikrGEr35ylytRkQXMDnMUygahzjo+84pWhZHeBhR/Wd6oh1aVabb/2NcMj4xKMZ965skB2Y9FM9
0e7V4wD41ToxowgYRp0GAcQNXtkuwfQWFXVljQwv6o1DhI892yPPVoF3JjW8q+7PU/NsTkEMaF/j
N+mV0WOUv13gWsMZeIBkS8HxxVfBSF2o6gvc6uT+YfbsU5ZRZYeui9WuU3R8tK3ZNoulSD3LUGZu
PyfzkSOTuOiyhFoeygTFKEIYr0Z0v4UvHcokUsprJ/b3ycuH9GoCLMRR1whtyCgeYHK1jh+J83Vr
xCH4FH3LiY7GFOyzsBNPXxnTG9+sFPHQ7lUycr2JcJ1slW5XHHbxwGkrWRPw1yPSuoDgZ5HS2WgB
QjaL5djXdRS/gSi0i3t2O1S/bAnPz0kLXWVVXoQeFnxdVeHDc4AAl9+jUjDEa9NmSJMz9hCB3Wqq
yufsH1EuAlsrkS2JT8pHRUO7NTRC52cu7oxRRrHDs70dfkApyEHP/52Al/n4iDkLDYwsoB0o+7E3
BISU3JFNarhSH0sWs4RkRz5MrFCF6Fxh0sIlAcXuaDi5RuP03ipONrSLarh7uftwFHZC5BeEPV18
UE/D9ZmWOaVlFjtNbkwJVLGQFLxgyIaP4FQTH7IcTr1ZVjKmEY0Z/6Wyh1jHlq6ppin0ftjwadef
QWZlUIKIfJ8eZHxdeyiQG1IOp07tzZM7X1MDcV8+jCTzUACi3Ezj4LqsWBPuCrbPIlsu3eyHqJJZ
FzENcYpqymZbg36Q7HPC1PaOZxHQavYt++aAcN6nFCcnRdfHcn41syeRJImKVfD/AuYFvVbaUx9O
cutmw65t3oZgEHqgHxmdvIORVRLfjt4vGG/GWRQIKVIALvgSHHHTcN63bNhAXuFhK82El31kmOjH
+90upmIyQDqCbuvutBsYIIozDJXuD1BeTP6YRc7jmjq+nqyEQ3jPVyf8Ni5NAuXtmo6WrXeFLmMb
Q0D1nY33J0KD9SKyRdKx+/dCq3tCmcgvCrxK7FaIDVTvbLTA1hD2dYNV7YYkqKUJiQB4GcrmgGPD
u6M/EWepyre8Vq3BVPp3JPbMBcdOSTQD3FLc3a/kBkXsKMWBxrrJNmFXiMWGWklpNUPH97+8K8eL
gfOuUbfOP4+BFP6POwbb5wlqge5r82gasLCvqJqNdlPUKCrj/qY4lJhvF37lv7NHybOrwyFTdmzn
YD2Lu9e4oc2BlwszYkU4OPn/t/I377n2AcUZ7DgWLV39NHn+LZ8OmV8FuyyATYo0beq/8VsT2rNE
TYSaJb8wF/rdGxARBlRET0cQMiWolEgAjn6ypm38w/7jWbAc6wogflxIQ4TBqupQ7Ja1hXRKrDnl
iEa1SG+yVMy6q45R22Sa+FQmxLJRumlQaJrfqdQum0cY+QonGeIa0jbdjPVvG/iLLVWBm7+Tyw0F
d+6cLxGH0sQXXn6Ly7JkrwvwUaWMajgklfb/2bCeq7n1StEOS8sqnHVSRQfYgKNpLtkNPrO50WpG
8KVPaW+ebX3uxZL2G9+Z+frz3tEcXVF/IJIzbSelnj5cGzTJ9556k1n3B+1fy0skqh0KevE0RypU
WJH4Obuv07SHwLtUH3jUNRuutLC73jW9WL0KnhjFYOB2eEcklsZbLhkbyGJV7ku9bCzbE63f27hj
yQPh6WRFDpUsH0I/0zAnjtLb4aiJ/Fk80gl1LGQTg/VydyOAaCc6nwca8LdKTj7J39P9s2e44XS9
Il81qgySJMDkwr+FbsnN1cAuIWdlfHvMLt9gBTXFk8RVv9DrrEqIvUU4RXJd4mym4mnZlWpvAjkL
/KhCjfwWincDhRHYQNewThbzMmkWKe46bkN038zC/IR50O7vhmwlQ4B2vaBQUlT134GHMjP0ugnS
OMzYNpWKAsuK8onAnRSwr5eiwprH/Om/StlGMtJ/YYFXSjxqgTzLSSr1zQzhRckWr3/rLKkG+SyY
v2HX33blQ4TyK2k/3cTK5ShqP6mZtb9G4gIj85vH6+NzqiBwaB+lJh81IJLFZ61tYAi1hyxofMWS
6xQDMqGbu79WtAr6nY++0gtMo0+Unfc3Q7woMuCu0wq3H9TyA9OnPIP50rBD+N5tkgSaltAUDXdY
DhS6dcHlT8LNfXUccyDGWCxTRujc7lxlcCjqdjBwRP9bnP0CUr8jEqdK8QYZKsmpArGmPjxNI+Ca
orA+8QkcWddy6ht+NRriIiwxRbux7ftySyLnnhjK0buZehONuOaIciBpKCXAeqyKjNbdbxRukkBz
h7EPp3dG1Bk+a+3nCgSU4zx7Kev/D8TWTUjDnjLev1i7D8vHOwWQ9D0W+VJAaeraT499YFwwvaRI
iRyGiPrru3RFFXd0hHGsJqeTZhCaQ1EZqrIfkcgpZOpdaODkgDzaPFhRJX+pngRnaQ2oIvNZ3t1T
azaW8E3qOYqTg1A0yVpgipEhO5Yb3NXlQnRdhWa8zhF9WOihKywZvf6ISfVZTDJx4dzZJWaCdD17
WD1M9FSHGhqs/GiPV0dzFMFgBHrObNMGoa/6glQ/ho0bmkXuGd/6UG7Bi9kyVWA0T49XSwJt1IoN
m7AukuRCN+OUzltZvkPp/3xOUO+2GEKe6bmSc8xu9R7bpmpylxZF8pF4LO5q/NXZK/wpvLi2k3yp
MOCSx4e8xNO3me/x1wa8ooR/VC1g9xQ7EPJu0p/LmWzwDXAfM1lydNDRxssQBQNYQUIniLhWfjhr
BRj5uVmNnelKYsQYQ4Z9jJXFvLIb3/36XdC4LUr/762rIECCQAJruSEfedjUNFeVNrFqOlCzWKv5
SI016CXy2Ah9a+dDNsKsmfzBMz6q8kVdocdWWcOx4PD+r51H7oGlytspPi3VrcdsilC3txCHPiMP
DrT5VTgdVrYxUKdLDpRDiXssiIhBzK83b6I+8b7aAjca3+bH0gTuLFQq5DPmZFnuNY6akCCi/0WX
VNM7daT+W1eywZ/8rH5ltRadxjZs0dSaHzOAKtwct+RsJO3fXVqQogsIPUpx0r6qKfTDetylEGHb
SKUjhesEk1+lz6dMqvUIUvO8+9HrOjjZwvQjx8Y6qyKtGe2rMdhLNBWoKjC4ncSqCue1KJoRxrLX
3Wz5ucWHPO5tFJ7NZl16WXVrjCwpOHdgXAIkFMU9pYNyCOkkSU293Edkg7jVstzHdedakjswg/U7
yulw81rFLH0dFIIC9CNWQPKAxd32vOgHfxAQgr2UFad1k/JZ0XuUns7f+k7Zbn1u0MDj3pk5Q7vm
+0zA97U0YG7pVK6c2DARkq5fGu0vdnpGN87h3yTTdbGViA3Y7faJM0W/D7UvbbD1+mqCn70Wi+OO
jibNc382kEBMo4KKQpcuyO3DOCxTH7tvwig6D616oB184ZdOQym25v0lxT8u1VVr53wLN+gNb3HZ
gsqbrwo8ncsBLRRNjaB+wIsbVylFd9jehEyWCvNTi03D6PN8tGrZgmqVbvop2TWh5SjP0I1xjhBw
HxQ2JRxisoo3XfT4yEzeAj+IoUMxYwTUS6YDr5FX3zqoaaYXff5zII3whypYTuosgXkj5JqhFROW
n0fJhkM/shom2Py5E8WbUocUabm+C8g84FXnjx4dWT5X6ng4y1UlI3Xw7OxaPBK331BVw4oJa8ob
oZs55bhbSD9QFodg1Waa1k+e7VXgT05n3liz4F5HmGCAR/TMqfwy2J9i+oB+TqmEm/LdbK5jEHxa
N6wxqIMM6y55o8yjbm4bup8OLJXgC/PS5AsFmg1zLnm7B/134i8ZfdcMR1JoLKsk8+9shuy4BnHc
+g+qwbfYEDdBn/UnCx7oKvDJbr7yJikV+OPdclAD3ac+M/djJesbzQrpHejlc6TIJoBrAYX1Vqm8
/n6tYI9EA52IEpDeUMSltWI+2bS4ff24vC+wOON/pZOHSecZbs/gQuBH6mtgAikpL0nm3egOiSwI
WPFD6iNcuTZJ7A8Q0+YZPDFxHJ0m9yCjyOkLevEel/BRK1ljMFBPQLxd9p56OIPVhimru420rF6P
cp2ZG7cAHguxugcTQFY+a8p1FD4RW0YAELleY9eE+6CL3vlvMwnGUGWzqsf6FwJBx7TXcF3z3NXy
+NQHM7VV1zsrG0Dxv1hQF85g05ncK8w7taiHiVvm23kU5vnnNGS9BC/3dMNRXQgAyupHr6Yb6Myo
KYi+rVPI+euN1nmplFi1jyWQVl/Ji1h3Aa9Xo8W21zSx5vi2vpuxyGObK6amv7cJmJ9+PLRKXqfR
JyqKZjWkDTdUL1aEtrThrYwocLoqLdbrvSw7eKbgGaDDesNR+hdTCZHMSu1TSxgSbyNvG24ehTh5
VKKTRi6bIprCbxkE7Xp9JxisTrEW7BrvoFlAZqX4N0SjqF7qcCVTWMzsqE+1jlaadH492PndvGrg
Rnp6KhUzANxjAivsBJGT6HlVPVp1FyzdQps/uTZH/j8M5KCmcccCLyhFWazSPaxj7n8e12vuqxFr
Qlz+6rTPGQCF1VkeQRBpwziRH9f5W2LpVqRHaBThI3S/bQIEugI/rq0mwu0uzMlUqGbWc+HKfT2K
5WRdw8lTd/GHqcH/VGA8JJ2QvZZX1Fn4ht2H4Ja0LJFB8vQUQcN62Dld4NeTBZB9jKY8Izc/tvih
rXicvpxV0EWu45c0kNM97qYHAMA9gbypBsA8AIMzVgBD1VsNcZ9y3X7du5XKbo8WDFAfe7A8N+FY
faHl2GN3BjRN7fvajLw/J3sj5nVpd9cIv3rbW7JjQLtf5ylz1zl3D44YN79p+kXFSf9Vquebl8k2
C7BkTwiQd+VqUFQzQ7er7X4Fy6tKBFWIaS66C5YPWMdNhepED7EQkWQ5bM291Dg4tZMZr1/yyV4i
sgLGZaUlxZ/XALFxUsNeXDOMCiLQSyttDOu5Kp8jRIFy/4nykdupnlVdf8p59JKtt9a9meCvtq/L
VdSjM8eAc3FMeD8+0AMy7VD0GsCL2BJeX5glxfHmDHFT1mtb9daj1j9xIiNTgoMgZypElRdRCsw9
R3OTdVTKb2QTe+kJT16xZK0A1Ypox8motfqELHvLptMZ5ZtY9cLEQODdNYW5mqx5H5oo+3tr2r0x
IkcngVoc9lEX9upPQ+x8f+4DcnXDl54w8XSY2Cg8wwRkDaFBl7OpZ0lKtWU3a/EeNu2FlQq6E2dv
gnJ8b/uOcIUwGhDZIHUxMhDP4RICCuZ0N5WWFxnJpr77IxBd4w29lBtSDQVbqogTLrBJGk19v+4V
3NSpAl3unTBpwYcyE/4Ou18T3mXsmRx6N8GVM8HiiX7h6ySv4/lVM4CsWenT1sZBjm86o/WepvIV
pP8lsPehQWk9AhhkYAUxeF56EdYinbwBqVnCmWhGvSwkXqg4RFRVcyEEoxn8fxynXdHk6ZWdpjab
/sUG4djQBq0b/H09MDNYgwaJb78U2DR7LGhb16x1wpgrzaiBKiXNMZjATfUTezuPtn0zahg6Afal
Al2c3pOk5Yk54F46wfOyK7rJmuk7KsbKWjax4yxLZkk5qXbnu+qCYNORJyyqhxuiEaw7KsDfLuCH
7nMzJG8t0wu91kchxmoTA0EB8Yi10kGCtPFs10BuvKQpEc01jyTIENmYvmTEElBwGgt5r0v3y2Wk
4hSwtdgj5JL2vvQKJawZIQZBmJJAy0xaG5Q+AaVfjK6A5bkYtkd01hzW7nQMFpdRdfgWtbtrZIe2
zCXg6j4SZItPwlhBFbx63Hbww3j/pNFXLDXY59RU0r9sIY7bLfb5NLbPHYr0EfK7qofxxLd3OC4I
/9k9pST0PyQgJy+ELmF5TsSpzot68FXDYe6fzsVRumuowNYurRNJA2Hgp3jw/ohdaKzMIZ9pSgbB
kyjvEN/JhOq8jdUkJgDXKANTt7YirnjpBl26bIswJn07/LSl5VakGATREe63RC2wc8Ua8prhIbyt
UHo1/73WoaII9/gzEuQdCdMk2g4z0Juz2hK/Pp62JQU1RWBu7DJsPfwmTLdHSrUtwH8M8ZpiUVKT
aWspjcMHjsQZ25VjGqSdRkWo3q/okvu/TOiYiPGWoFuRmSScEG9m/EjWGm9ERGD3i+yJQuyAF69/
0VQ3R+7e2ecA6YmOihWQBA22SqW47/gzo/t1p90tJrhG08ZTg0zs4SyK7g/NUily1007+GqVNlUo
JVvBb89k82agSSQkgyPDj4yb0K6CDUZ0+1fA3tdotE2WLpk+zRD5DI7Vq+qPJMCztPPDJkS8dO1C
1Txe1IFeguSJ6PfwqX9DgBaIgrCE46Ab0CDHdVJMRPCpx3kUIz8uUbsCSZUKm3apLcLDanJP2GBj
TMB+C/XDTYbxpQu5G/Tpv98hYA0bjr8LJPYUwaYg1WReTxhX4lDUxW71AC8X2mVfzyMFX6OSZTjp
n58flgRm0izAbBfhiMxqj+vkY8Ol10VhgUtUzHCsjFb+RLUF1vlJggrO3tYXODOfcJWf2Wnbk/fR
yqPydKvDzO2ZFNrDwiPNaXEDcvmetPwrsv+Y+pmrdylIcvzx0XpIGKG7nOJI/NpLuVHdbqyJcyWW
f+ihyf4ddr47aOm1PObwVjotGdAGNZ8w+1MropfkS4+FROGCvj+73/Ft9LEHj0VeAwr9bsC27jW6
Ux2FE292sxYg163v0Srb4gb8a0mTcYqpH5OfndnTF6Pydi83nXy4/v48catN4P+8P7Vcj9++qtnc
DjUYsuGF7L3JNqXiBpG1MifSC8P/WnDt+HDgG7xP+TPGcBcG/ouf6HzJ4TV1j2WrNH4+PiLgct92
tMRR7XvMInjtYHeCHqe/zqEt+vhw9q1KJBYetoAaQjVLIBaFV8brHP89kTr79G3I5GmVVUIxY2TI
LAeMv3pMY28pFeXTl5PapsXiDGbMB1+o8ry0eXl8mKLQEaEYLHsQxWmB58QdqRz9Qf3SniEex63n
/Z4SVGbV9t8BlZ2lAdENEfGQ+A197Pvpz/FgLXWNB2U557aixPPSXimyIBgPGYRQjng6MtEma+Xj
dtu2oinQ3M+BZdYCN8gv6+jbh6f/Nl7dY+953gP3mjyQHSeIyKDkIGtscaaLwPsv1BQqnXHsb24d
W54QKcg2ivVoevAayrSP+Bm0Y6ydzx6PaGLfxBzjNvHRGhvlcshE1rXIusghLLfcXtUAeuP1X/UF
w88ROJgo9V/Yj992RO/DcGIQqS+HqwqO/qj1EOHZ7RH9RT84hxqHZl1wTROM9zP+r7tDYStMzG8w
zGDplVlJenIEw/7vPeluN48uYXMZqYOb1/6LlhyTAS5D+cdz1SYxsLGknSgKyRl2OKatFs19U4se
bHVj7oeu4nPfRDDU6O+AZxos0kCoWksp71Ce7FJWhzTBtnnLgr1F8VrwUYaTTeXlz9c3q6+eYrw4
BgAXomEGKy0PbX0krV4dpXushp7NfItVMmWYyxMZaONOjbLtcXM0/iA4LA5GuAFtwO1SyYi6/wR2
Rdtri2/0On/9JvsNUeuWGw52vAoZUROqHdS4JOsgS4N3dqKgQr8ruJzyA3iwaRyzm6ftEoZcSdNs
1DUm8OrzAaoOD9TQnvu2MOFgbQg6MniGodzju1yazsUpcrinCkqWBpSJCXySyZ5aN9eIPM3CvEPO
v9fef8PgbvKwRJZgTPGx1ntdBJEueJi4REQg5euiur6IA/vhMgTOlhFmKLUlH/ULWHqN1cCwGTor
0lCsYKyV83ldkyA9QDc1+dCRJrFGrQnx+M+VGOfNfupJFoHefr7whguVTEL0hGY7GbxtAHKc8yup
n3TQWM0PyPr41z6doM2Xm1FlXmUmwTV53XC9hsoVCl9znzAGaY3QvsyIJ0Oprk5/g6oSiE6B51a/
rJ8SvvwX6AASHYs4EH5jFoqr2rXg8Qnmiv6CsIUg7VcPOKfg9cKkYeHFxtaiREIQDnsRjfKkFUuW
lhNalW4kGxzc1LR6EGIs2PxPZ5Nu1fLh9MImd7PWn62ePNYEs3NB6X92NjvjTChJksNjHZudha3h
sZmvpPtJyGvoC8iHaD8ulfBXRlYrCDkwi3FWwk7jo+4XnRRcqLm41nk9e5BEKEW7W0cMMPMtKdOC
BFKwzIKcFOXRWrutqkDSpBhzEAgmlwDf/pC81krz1X7kUh8+gIdsT/PO5fHttDgVH3VW9NufuA15
vpPThZQ6GelsQ0vXLy1zAKk+RSqyVU8rU8BypGCAkfKFZkcfzo0PckJ/Vulp4BSO2e7P+6tjhzuM
fpFGVm71toOphNeoBrccfKN9qGn5oyruLnuZ79zE0aAN0g0m0MLPoGt6X3KEwVFQCV7yXUXn9DDM
yVl5gizjPVzwhWB/ObfX1LwhQ6J44m1HESIAFYXREvY0/P0j/T7yKG1wmflO3/yrivogxMnPJkAC
iZHKvkoWZlVsgmSdRV03F7DXRaM3G/wl20XFbQOsD5I93dJ/flBh8Umx9A0gWRIdzbcyNZaYyvNl
ctH92pG1jn/jCdXUV8gduHGXc1P+Yq/kj73ktcttoQZ99sqL4k/qtT4KAXa373FcAv9NgayrsfjV
WDudgNt8/SuQkkkD/BWrj1VptMMbK7kd2YIPHX5Ld2Ctgw+0xWzcddJmEi2Y4FAPuDQiPG3Zj23K
XT4Z/PBaHSWWuE2BZotN5da6X9kqP8zttVoqYn12I5ono8XRgdy/3iSyVZrlqQLs3QGwJapJBsL4
A8PC47WHGdMyCntXAnvpntPC2qeeO3fFUuMOOCaJcjaTcM2MYB78wixl9Pxo6h91/oLXKxZxyNwF
bRHO9m7uDJ6+ilfSKLrlDWY/U/b6qjqH7mcxYrv6pEpLA4Ejhk/rAcZDSl/UQ+yh0hV+3UAIeKGj
Dwdli67jxR9j41b2NAxskDer4onOoG78o5UALfYvu/CHwdoZ895I0jp3Yo0feDNBACUv6nyLFtX8
00scZJiVFYA5ectMS3N9KJoMUat53tiR3tE0Zf8K/OpTTFAop5ldI9EvmoTMOL9v0IreZmS3QoyE
9/StWA/H9Ep16tMjHn8v8iDhL7Ox+mMmXMKIcQ8B0RTEw3ccPrqfPg2HFcnOXAJMPdu5lAkBevfN
gTDfmlv9NwuOGtGGeKyeu2ZcTNXgPbmATjtuphQLIZZe/qQx/7RAnmy7j5S1gCBjTp5l/xfxKOQO
tV2YuCHOyaEFkh49vvOc3Z36LiZf4cYhxx3Ca4K0YAAOf+X+ptJEx+7/K/fZS3Eujoj696+FmnoL
GobAr46YuCPWECHcPfEbotZwCTZOWauzxbRyIMt7vTrHkLRYQb2VLJPcEQQ+07TTDDNYaP7D37Lo
v91fiiFAxK6AKDT7ssI4IQk7xM80CnYirljDaPLpwr6XlYssm9+1r7iQ1/DUN+tcKHdqM5uWX0XF
t7jeYdFXBLEMhs8PW8yvTLRxSetCMS1dCEOO/9gYAnHUP0wyRzPN15ZxakIeYh8G/Rzyjtk4KFbh
yvFJOubuG5zOjGcmcKrAJxp9gNmSo5/3I5Wg7aAwdIpxupI4VHOm7OJ/r7TPTtr/Y9dykhso6bEh
KWaV3VBwwWCCAOc9dtpe640o0JeYozkzkfapgsnLGFLdL2z8OFfOENh7NrzwGfpyM0Fmz+xpsjOG
akWiuGd/jJLk0f79QNztSRI7SjNdXnqJg0x2Aw0vS5yxWNjIJnJft/GLkAKyKsWmK5/l207M4VjJ
sdjAmVampgjac69jONaBQJdmy8fOnpqZGOQ+9DtZuDuaGpiMXwxiV6Sj85T6geP8Q+eEIPAaHRRf
wamb6u5f4WOytU7ngasi5iyHdCMg+foy/TmBef5N5hQa7ocm8/l+QUcCgtF0DN83rV4AyOTTdShG
ev/il9mXfdCZ2zIQqwxqFsNGEeYXAEFPYM5KEDBX2ZQ8Mmzxo2zyyHiCFoagu1EFK+zeGaKNmQvs
rMHobnimJCAFs1RCJkqiZl+dCseI1LRfd+9XNNpneLWussk5h/nU/gO6I89DT6YeMYNfFZ4CiSDV
MCg9LcMdQBSMrHgs9utmjgTEKn35hr/2JaJV5BgBr9iVs1aKIoTxkf/vfhdnD++4aN3Btnokv8Ei
oCHI+vbJj3U7HUb8L5iiTode6NTbgtmXFfT3dT6AiczaygR6HGGvaeXmo7oLATmnCrFGhrTKZJse
5Vfl78KUgkJFx1NgicB5PnbIHaFxB6zaA9XsopKsd5jHBMJgQT2rbGgvEG3hN1EMpZi5IXMEKXS3
T90gfUaIpjJLQLBcGbbbH1hNWE8owXKFcXiFz3PYTEsVubMcXWMUaO+4h0H4pWEBgJ/G6X7sivZK
mRTdTMa8kNp+qo8rN3rsEeRPATPtXs4hLxEOq0lOvO5+yHZ5HPN2bI1DHzbXV9qUz/4j3Kb+uqbU
1fhdCBXdm4+dAwcz5t9/1gpykmKZPAnI5qYBpKaRAY6Yi9DfGB4zsVYc7HEUecEMb9FYTPa4MZLk
VXPlfwMA7U6/Z7rozuoCUAiNUSVN/ort2CYmkgp7wFEG7dMnMPvT78t3sOqsLcswo8auV+qc7Xqh
IftipPk+UYxYgVj4Rs9f6Yl2T39VyqtccvsjKtkcURmt3xnkjHTMI2kHV618RzJPYIpw9HDCHyXa
YL4KjmJLZGG/XztZF+VdJNeaV8kRWnvVbdtlbQSWiUtEqPL51CjKLYqbFCskyOURhTz6lP/me9Xv
w1ncM17J/QKBLNSTXaXM2vIIjUCY6rDkhH4p+QYK7QuDdwDs/XU8PGaU0CBruKUXQSZzlKYv9eEm
tn7Zaofc+eu7PCr+i3Jw80lllDgotf1nUDrajPfuj3xEJ+G++VD1aVFZQUfhDWaMwvuCugvl6sdp
PAAZy+fXgNE55RxZbvlsULOeTpjUwcwSPCa8MmwUFMwbUzF1wFNxRGHqOnlY/51mni+EowZCgg+q
+lEwECQQh7MIqmRsH8kmdZJPNTi8Pn1I91OmP6AUPfrjG0dIuPPkJB3Xat3f8eB450lo2zFOPI2F
3OYisSJIhOZ9Q/ixCen8p23rwNxiER14G89abgIGW6ljtwdZDZm2KZcluRpRprucECfc/2TDnj0y
my/H+LGqIsfB0jwFmTuduItY4QiJLI6d0Kj/QHMheJop0XdUGgamj+Cl8qRjGzIHnaYoGtYMJXu3
WtyRMpVGXNoWen93l+RctvmTllqoPpjm7CTuCUxM9jJ1Kvfr3eeuDtKKu8Rs47pi+dMe/klYUZuA
dgz54oj1+xsHlV74k0xhOH+YuFnrClN9PxWAEGWMMORLmEJiZid6L228M6VhR8eroTJFGHJqlgjm
8wnqOtvSj62GjPgDZhecciordlVIxCGEsKNaJpi0Sghei2H0OYCy4hw+IKupBI9pfPiR1CjFmIRJ
1WdXbj+ypKjv3+DmlOP+aBkVxOG4g8nCntJqnb1l/I5313Ye3F9FpADlHx+TvYbq1aUyA6k6vcTl
kvhr0RQv+J7Ry0BiEXl1UGM++XnUyvc+VCbDhNb+iSjAYxMutuDay3oxpgx6VY5D6kkhndTkYs4c
ZJNFdA7lVAwpKgRYu/6DaXam2nGjvTYZPzZ528xmlNq1aGEzK4hgFK3pL8WlSgDcDHkswAq9lzot
XBYiM+e6ROIZpnDhEiJIRkasYRNq8ud9EZH2bxODQgRrtbKBoQcm3SEHs3S6q4g92Pb8ubAcEWq0
YOe/JyEgrbrxudzAAqsKdrQMwvjg8ezghM/BYcD6PoWJpg2hSQX09sQI5FpxSsWjBVXh80HPMEP2
FieXIYOagDbNck/ZuD115wz8Eq3lsMOzNhOuOttdLB9WJdBJxiILPM6pGSdas9d0neZn+Odz82Af
jLvYYMQlyfjDMwv31btIU/TDOWIkbNtav3sbN8kROTchd/TVYweUkUwHDWrHR1DTCOALdoSpkhI2
MHpZPf7L1ZWtWRpMCrcac8fWxQsQzZ3Lh/bIq1iCO/8OmJnJV8cAQEkVyIQeP2BcE54Pm8SJr+eI
CH4c3IfMtrHlL7fcW2sVlV/j7xegL+qHb2k07j/1e9lyIYKd3xRstpT01uOd09DSIlcdJC0cWkqF
PzTGbflhAYSn6I5oSV8MmuhRRlc4Vvvw8fSQ1TbWniFyyKeR2aTAzbw8q5N954VQpr2StdATPSIK
yP7UQEuk3EGlwBKy12ml1IMS2+q8XD2tbWPFCk1cJGQSgL739vrgAmUbF91dyqLFQ4gsDf8Xu0Qw
6fCbLD/Xr67T5iEVnu8zS8QmUzAgojsVmGd0+rtq8GdqbZdAP9L2vzCNRYqxc00ttH4g2GKZFa6e
2aTka/gSiYO3d/rhxV4T2eYTaD01uT+RYkEhY/6BGpSC8Q6515XOWQrdpqscgju4iJWti7LknO1g
4nhBsNaLpDSoLwI9nv/VLkuK6N5q5P3Jwg//w+QMd5Se7bJvOgvqMvZ2ajcp9ah3KIzoQlSinCyt
TIBOpz1cI9lW9/Grndh2tNcimtx3wuKWYpB4sUBRenv53dqL3ev6UTMcvNR1jj4YS9un4WBKLcy+
pm6ZDtbprip8bajuHm33FavM58T08IxS3Y14g9AcwMwqfaiWJ10i3eeVpiPTQB4ss5qRx8MKoV5q
mIBpHjte9L28b2RYi7sFaQrHg64ohcZCLsnLmZho071qxwZj5ksm405+YKdWotx1RIPWWtxWeyxl
4oz22MOxhf8stXEWOB/7gM7+CimepZP6DBBayd0695Yfid9PZts+DhVgh7+nIIVgHx+q4r+GctRW
kaJcAYror5vpXySqqVGo4ccRSxEY6EniuZcAtQAkYE04aSv+X3h04dHzogdph7fauzQr6Hvst9WX
sA6kq9Mv6m+gN3/+lJqVt2k/IIjWHLt/xpHtSxRWsCHbazsfJ0T4a5FVjZ5Ua4d076wti4UALFv8
oUd9w01OTISyUX0bgqFcCcys9dwFXa8MtNzPASXCIeaqPR2xKFtFqqCPIBekf6VmFrXwjVfvDJ6z
1Gr9qCqhI8pmoNEP5+Vpb7sj6LaM8G6nGlMgK/Yjh1d3VONSic417rFyWazpCMpOJHWzRHbevblU
HyiYyXFmZ3UgYO2v0qsWI6H91XkuP+v3pd7wBuSPub9PZAtTDc4Ihpv8nAAEh8YsGCGIV8q6ekGk
KiWgJWTUpzNJJzhOV8T17OX0s0Fyw5wBrt6ethZD/ClCzqlheyVrDLFz8qVAwdWdkAXfrJe8D1fR
BfnO/ofynx7K+Iqk8LtEOCOvtYVJ3Qzy8vhan/fu7oT37IeehJ/3UQU492hdM1ABLfwdaZcPPub0
hW89fH+omLcngv3wDwwc1S4tdThEQJuSI+vNuZ+kJ1Ga0ubTrpbVApLgCywhmr11Th0Yer+IsHz+
DVFdaENWkuSzS7dB+NftL6ZfgVsILfDed7vcKKdJ2ux3QgZcwVu1zRLgHWIMCQk27eaABAmA9QR6
lX+wxemMfFd78vXn/K31930Ui685F+f8TITWBjBsS9LEwIaH+Fw/4dhLvtRgmchintNDs8yrvhEd
ejjHuQebxe+QVjGWUcTHER9DSJroav9t5Zr4R8sjguVjsD+1/CUUXc7wYojzgKSJH+YqjdzJFTuP
LAgmhohxTDbczGgoZng9E/yUUDCYDQ+ywW7DyDw6SMrIcN8X5HDUJtzbMKnOzN5U50C8hatUzK2x
Svr2gkpiUQod7Ydc7TlekTnpmX5m4iW9ox0IgRnEHkZzesuKfdHcSoPEk5H02Drv5gNcKyQ3B7X3
sL+VLQPaLXFfH4B/8qY5FWkFdpclAX7kK5vC3NVh6N/72XUmdj/6FS/yMzul1U71f4cKyrk0yd+j
JQsqQARMfDhWgjY3kAT0bYb6V30Ntsz6h+Yo3VTxJhOx6IStsokPjtqfRppSqDAmAOthAOxISwtz
L8SqxFmbehxmANt1QrmcdZVUYt83ES9WvPX/fub7fvZnoQcWnAkLlIlPuLO4z3U8L2lalPJ+ZXeT
TAWh2fc3HcUSXc7/hnYd+OmN62FzkorXyKQJheX3jqOrUUIOLVDvBe6bGf5Jm1X52842r0iYsQhB
sKz5ICDmjOdwxhK8NrukLb6b6YLYWJMrujOp3QCxmedV7VMV8uEllqHhh5DZqdoV0+JzaARjcma1
HemDDOzrbkKSC6bnLGRcsb+PBYigKt6zCBbcY9IwFKUH77s4tdQBZ7z/2tRJNShD54o5Iyr1ZvVm
U1neloBmEqtz/NtX8wIit3N8cF6lspPEMoKTJG+NOSIRmbAFQOmT7NFA+i5PdTcDeo+uHhicGf8D
dh1WKjeSSE1qVe0jGc3rL1MWlJWFziOfedp18C0IjOL0Aj7fWJY9/x6H2nTHzFy0Wbjy/ZAk2MS7
bLvnMX7TwNN3fCCeWIn5Htaw84phhJusmIW23vCucxfCBYzn+WFGmflyN8yvIL8+Wn8ujazQFnWO
48pJMycRABw8mTtrEeP40yMYoww80oZLvX2kkG8RNhCty81VlrN0Wkep30880I0V9vo1U3fCpfzn
JBCcOy30AQNsz98w62eT07kmziih3b9xgQb7cVc9O1/Av+9J7Fe1/vOf4Z4iairBB7u972vH37oo
qQvM3o9gVuRwmo2UD60M+mDo7EqKJwwGZ5e+bLVvqCqy13WjAVxujLoxqVNEhY/DlhpxgCONvjci
MgiQ1vdqBAshNq/l9CS3C2OT8SE5zR9BKMf2tOHglBLiKtRLRwWosMZ4/bQ8CMYS1JR2pixGIOgQ
RTgtI6urVjC8KCjvNIUBztn617a79FKAFB+2v4sg/wJpF9/c9ryvelvgDBxDlz9CPoVT3wQzYv/w
p/eW1l4Ejh7PpefrMP3LDSQWPav7feM+VdEHo4JMO++5KjMR6UPAV2XEuWYeqmcC6XFUrZJoEE6p
A4RK8DZNeyNmnKk9n87zqAZ5ce5qjgaPFGDplsO6h724YqnJuiNI7wPbO7dn107N+VhE4GLbLNkI
rLjqmOC6hf79DJB1w3Ucschc6J7j/WgYQ75qwt6c8MzKnzBA317GTMJDpYqQd/lY9gZDbxACnFAA
na/FdIEjUX5KpCwCqqQS8ixzT0zBcuFL7QYWWSYm32gGXri1A1qXE8IHfR+SESE91v7Ql+SbvIbd
eS+7SWCGadGg7q/l0nbnsHMkpGC+qoxniM8iroa4yHf7GWRBVt89ZqVR+tqhUJ9YHizq10uM7ApB
bxJgmr8lNQ6kSZzNg9dLgTvIt/AySSXzUVS2NYc6ZKdUv3z3XhwjaMQn8tSWiijLl44pTlDdpwxS
bsm4PQawBZwPlAim/LrNho+dm8hQLO5Yv+tFrGmZe0XjgO865hMxVto/txFxidbQnBAbzh2gHdOR
jkt7ybxnxgVH8g8yOAdEJ7OhaKQDaLeXsJ9ulYTIoHoWMgORZiZ3dWlNhyJb+Pbo8onmOFyWSwCY
xQepjW8yUmrBsMwQeeEGLtq99JquMV2yxU5hEAl1EmsoLXdXsSCSztYRy4LqWyOz8VHmUMlWTwpb
yDnaeSnvE2Q1yhzkNqB0uTgrmQodf73tRAYGF3q6OYOXaeAdFS/2PaLiPwup5c07vdCzaEgZ8fLm
tl19Wt8Y+wZMEqT2mPc8lvRQSkbblaaxavLYea4yUm4f0ZeShfnGfbrVB05O+ymDegGge7YxjfqT
zgRMmLhNAyKWcNzbHufjMH49O3AmEb96G97r3Vr170FgL97sHXVWnmaOgxIqTKTiEj+tcj8aL9Ej
8wQ/fbV3r7a9xRquy59gPJ3StMBXetjGp7r13ZYZSwZIIVdCVcZNLuDALdT2oyU5o+G+RX9FYmTi
oHOtIg0QdOO425bgHrt71lZCf6jHz3O96vf3hn54hPxwvBPuxJ8vipm0xGxxFk2DVdOxZb21QTMy
SiuIw9c1e9tZ9e8+S9mo17my89pqPSuZ+GtdR5S9ARXWwHrc4mL5RSEtsO5KCGFLx7K6Noox/VG1
ujU/3nev5Q35nLEzllpfTsFJMq7PSG8DGDEXPJL3pnUIj6qWNYnnbP4ceNpboyIHq1M7XutJkqhV
jqZB1WmfnTDQnxtPxj2nVJtX2OP10jiPCPdFJeuJdNEKY0IbiV5yKL1X3SpBrvkrzo/kz1SpInwI
Ggf5AiJEhxCpC0PsPRdo+rnEHMTIF8ym4ihZzyGJhSW7YbnOdP7bAWy3EGKS65xL/PiYbBLqaGpM
jjLtxIISebXW+yc9qWWIX+6YNoA/clD7nGMs6ZdtIJdmomFwNK/Ym8tso0XABKP0YJ7Rk1VTOJpU
PObtg8xN09vCcNXuLKc9qqKcP1KTikX4aZQGtFF9BIrknPkQ9Pl+IJNf4xZRRRmuylgDs20wYuoF
Bqam/XdVdMhzu9rtbv8HCupRQ4ChmZXg1vLBqK25CITSxBmAYWKBaN3mtwjfff8NZrfEUa2/KJXS
hl10mGoc8azRhJQ+O38qy2+WOEq3dHCPH6CPoCkiepohW+JH/kV44TsXt0Yu+Wuiht5+MC3D5HLq
d6fPWJORVP00u1BgYcwdq3932juAn3qU26YtNXl3Df3s5dHSvbSejSHi5fxqZN3MMBpU19JUMLnX
LXi1lSjwfOPukh7NFa8nc0SV4R/SxcQmgQ6ea7hpMp+nRkTD9/eGFPktS4V5JuSxvehBA91Wn1J6
m0ujkOh0t97ecCacnKhTJtprw6Hb5n3UWiTF24ryV7Su4WS0aPYO5Yxo3yPBp+rup1dIjdt590AM
lR2TF3YkKrm/hPnFhGqXokWOTz7QP7qL/Pm4MtrrgCJpYBomHqCgKE9+Rj9Ch97llf2uu2B9j4qj
VMay09xXVnlY79/YV5WFN9iftNGnlMmAlJZ0JvZxWDgqwv9l1Mltmw6aE2o+h5hKLSy4wpXDGcGM
6Hv3heapAZ86BMEs/W8L3R/76KWBKOgJjFtCnvcZJME+I8W5RBgI/36T+xP1Z7X+AWD8R8Vmh3pP
Vgda9Ox3/SNrVwHZuvIP8kdyt7sDlbkA8tyiXyfTzY0EU74brQe9+DSB4fWGe0jBtuP2kTxTQhfk
3R2uYz1nFintswZ6lfZ/mQrbMSi2CLYjbCWbMrOdFZiUAuSsZ3Or0W4Mp2haZREJiyJbpmgYL8E6
I7BxtRMeTI79VLioxvVDGQe5VVvk0wIAi+iXqYVLYtQP4STtKWYR6FZB6Vlo6H09ejsrz5Qk9aVy
0tmUZDSBtP/hEM2mBUQEsS2u6Z6gXqMaq6e1IDyzgNMcO/4Vbu/EM9JxN8Zj6Or2+XzLnBiH6zF4
SPm7r4empfd1lh+N9mlFjL+4KLmhwncckIIxb14QXlRslkyXQmHCJtBNRttLvgToNd1z5ldzGVNW
cw5BtDI1hqp8WV6zR5MuVNegnK5JawWp3ol1by45amGleDxomKGlZhHe2QEh+0VMb/tZVRIbEsvM
mCOqGmXxYO+YFxaE9lVS7CPRRYaRTGHpn9xAdUBZKUt1xX5jU+MY/ZifIqb/TqYfS0oCPVLoV6nh
964LwYn97rthOZ2G9s/TwXaBPXn0cYuOEw9KgeqNa1YoZozINctimK9aeXKaeZY1eSdj5h2vtkSB
IFPDxxqQbD+LsskzA3tRe6e1GNDKVvOBYWq/2iTHA+HQXorQxb0WEh1ieW6ReKVvSEeb6/0rXhn2
+3HW+TzirjJj10JV9Puvr20ORWDsXQq4PXfCOVHa4h4DpHXsbpgryGoPzysMsaj7IS0kSiMzpvef
Si/6aXb3y3rhcMWRNF7Pd7M1Oe+v1u4giibaG0OVTmqGbRb283S70GTlc31zLrVxy6MgeEjvOKia
a6ER4BoxPJnFuhqf/q/jQJgs29cPxc2NhcCEhOKzYII+Kdj+PHLtPzSklX5YmdOld1MuKYFu/RHZ
z2IckHAtcv4q1wyuKwE+2flDJIyuCdVxtRV1Jn/S9bKuobD3wLKTWBXAb6dq0xJAIUhOoZY+UKdQ
/UrZZSqOcaGacPa2QPdhET8DSyeqAnhJX9UKl0YKSVTHxcdfwsQCsNPDFMwFWyyj8DbrNGYM12dX
iqwHLZARDrjigrzgE5UPnqDXyVYuuMxjWtgzuiG9j3kdIOIk/GB4AAXo0FQjBeD/oQSW5rbnR3H1
sEqmhU0Z3ojNRffewVEagL4p6TJkL2f1JcqQK85vBvnniY/Jz2BK4JKCESbPfzC+1sJo2b6dR4QY
aZVBO7ChfjALnuoIFzIzq1Gnh9NUnCl6RVSCN9QzLz7H2pwQjIoUHLDQYRS9j5FScwh1c/unZLea
On9vLSBPmUCiQEjA/mJXSTwzxwqHTkilTZDY/EsyjNj1FXSOVjnuPpuugGL+nmysF+ZYbYUtVCr9
lPqBEqUjGfSzigHR4VfJ642WCNMXItO+gdJHh6xv1E7q1vCgBjZdrsWWEGnmG/W4VBg+LWP8rp78
whFoX+MyZdVRUI5xoknSZWv5KL2td84zUEtB33uj469FCXP/aEMQPspVQrdFLHol2EU9TwrmjrM8
1fcpHKvnzAX4EkeY8wb00Fmpvt4BwMpmy8fVh3XRYeXhJ5L/ja10prFDMQqQjWpFKGTAabVAqYwj
nlV8cURja9Re5D5gGzVtHyy8t4HFm1V9Td3HvVbX1Xl22GsyO8nXZKl/KfwRC4N+k18fP+QckTY+
wyrnMLYB91Cawkf6oDEY8ODUC4vLitDi9YTh+dDgIpaTwbX5R7porpYSJVmLm/LgLO5cE0Jf8Z4W
fxCWvA0IUz1X5SKMNP1PyaCq9q1s1gvLgRgCvn7xvuxxYYn4+cUXfHDKS7JF6pXaekU1C2YjlAlu
Kwew8Q2JKe007Oh6BKjXN1ggR6grIUVTGAFU7cJW/hHoWJ6/G4LIzDPth05vGwbaDsciX4v3g2rH
mtIaLV6SI1GSwt/cX2qSRyRxNWQ+dL00g3rRq8dPhWBhUmUX5I8weu+WZGRRDxXSyWrAt9ov4K/5
F31aKGdTF6R8A2jemdIylTq1G8nenTIxkPj8LfUUOABtm+5HcHHrjQKWdtRPL9z+FXMINPQXqQIJ
bjVzqqa5UpIORDawIN4A/8gURHlKBklEMyfjSJTP1e9hmHna+6/D3COwlz3rkXgd087uksB5whAq
boV+YtF3s3OWe7lOonqDMbx2V7i/WYHBg5J+Rp+iE+am8QB9rHbwIhlTQPSGxx56Dxe4Ucz7JtFf
3COBH4etMQoj0LCfGidmYSJyuu/A892hrvI/SAsoCooxV+jjDTQNz+pBV2xQ+XW/h9v6ml+8ilCT
sT9KrEXN4u9gSAKQ9n4O3WLnXZEOrwaRSAzk6BGKjr7131KZmpPYaGV/tyC7YI+9xKSN5/PHxtSa
rbwJ6fONHTC+ZU0ztgBSQ0gHuidcyJttWGEMA47kqytoY7nHdrxmeHz4pIRZaHJWygpi5VCV28kp
YslpXzj6o/6f2YFAnYaRe5RRsN8qFa03pILn3iOdthAPBzwTT89QDgqMmGFqfKSaAV11CNCJ9aNJ
c2jOzLRML5GGU1cLza0m5ZeSAsNO9QvQdXY1WXc3LT4dkD0h2w6KSZ20OPBx7UP9xg96HkYONKJZ
gwB8aLQWqCSunB3k3ku3PQK15aRbcPlEXlYy2KTrVP/vVOTZs5WR8rMqClkME2mvLm6nYD0jYY5U
V+/7XHDb0jBm3vFfnrRt5nvtEFK9ShSAYf8MUknrLy1db2c318qp6WB6ikTBZgTn6DIBiwGkEdTf
FrGiAAzOTefI4Me7DiKia0vEI9IRXqT9+saZNCFb8AlDY3FOY2BXm+aRJlry/PxVrpLZPI/9aOcZ
86YXf8oSU/9AQoR+6kq4HJXe7iXy/q1W/nneaJDt2IIfxyDTJV924ff/TmHLfAvw4N4DlrlsQaNP
mxxHIa7C7K8rmWRXe8FswMvWVy4dfmdrrGFgwMVxEXP+9RiEcJbsOVRrPB3cqs8nnkYj/mgKpn5r
gajFNlNLwqx7AuoZ4rllBUmxTs+t1HKzp2Yf1YTY9x/dBF/nBgB0bzLflhkOrsBGgvbRSEt33P0h
Jy1fzO9mfxTTd37RbC/xmWJPFj6KiCBtKjBJK6jy6LRiAkEt5pkUTaq6ji79QTKVvio7F8MQcZ3+
41jHy95RQfLZ5gzz3/siKWJk6ldgv/smmql7dhj496zek2rrUpZucrcH6Ui2rSfVczlGamVDkI9X
+valKc4EyilIJOkFWcc0Lv6z2ZHviA/vDzhf5bOdOEwIvyC/v7PvmQ54/TC2CkWCJAfN46XnWDFG
IiDLn/IdEZ5egy3+zJedjf4fbVZTNKgfFWJeUW+Qmljc8vdincRz7NTnvEkaSyEOCBxGyH67Hhx1
u4+YM6f6nLvr73yXn2tecWNFSMzBah7+e+bh3WMavViwCkrCNmfpIHyL4b8skd84oAzP/G5vlBMn
Dx+uoz/ojynpYXMF1sm/h/r8/QVtPJbW4dspVzD6sUG8NI8V7vCxRP3b1o2tLasojhr7AX5ChASg
P+7F10p10B41Y1ULDH2893fyvMpYc9+TQo/0Br585wNQKnbXuSEW4bDhdI8CJ+PWLqsfhpDgsD5W
mZ5Nuz23nFqFHbkCoL3hMOAwvu0c4bvR+K0BITUOWxJyxKSPPUO2lpFGT5rPQLTHauBDpOWNhzwe
b1/9GbBVQ6CTU8x1rQ10ZnXfc/dA0qqj2rXDcpDBFZwWli4XFWbhfYgg/EHkm923aMTHKKZI1jv2
1wrOhk0SApMg1iQ+CzKbtUYG1Q8mxV6XB+n854lQtR59DqKhLP/iaZc4HcNy6kPpfuIGQ148ecrl
VM5zcaMgn+r52ejxoSXcawVlB5IzHFJaWa/R4x71+6yDAFeFkxlZnXYijOT6xMUHzpM4MI6dxKx/
0/0a7TtEsPBxAwDDA1M52CnfZ52/3HRJe5ZwNG/aj/qeGq5zNp5ppTls80j8uOjdiQBXuWgyaTCz
P+zrjmjwBvyhp+4Tp7v6p+X5/Gl5rr2swdWRKszl/F/Lu684GPGTscV+ZCibZRDmaWB0+zxe2dMU
BExgoOjfTyAfhWz+EBHqebbylWoT2c/tT3cBWxbnGodIYwKAE+tb+0uhJwusBZlyWU0o5PF8VjyZ
tPesrTp/FFE7QM/g+mG1LiB/co36bubpM8XbbJGW0ikfuuhMwovk+E+LI5uvPdOzTseZdaVEs3qg
8MkxcCm3g/k5Xn+hWqaLCILAYtFGnDtw6sDucu/DFbM3K46UPH1xIq1Ha00qm32Bhb2cgQP9TER2
J4Vrnc8kbIMAfyW1hBG0HDjsyMJ92NPh2gIB035ZbUSrG6LTkCXZPgTtKQwjGNX9559NXHVFPPI7
6GNqkQK9Y0hHvs0XslXBq60e2E8IunwWwKei//241AN5aA4p6Ie0SUnYdeFXMmRjci5sSOr+M9cG
n2+i4U+bIF1cX5ud86tyzTvVqop8UD1ZDOyGYE5zgEAG3eZrlNyasvy6Xn54OiXFB6MGh8STFava
fOYwiLVxIPfnbmQhVNOALBWzAfCAsVjZXkPt2DPeX7fYS/aSqZAZt0Tk6wDSFYZGj/wNu6lDZYt+
TLQIZYkS7UIQBuAPde7+cqQDjSJC6vDqvtby2w8ey8St2RPx+1A4YsM8NgWwp9G2U5Wd2zzI5Qqm
QYkOyX2evNiJbtYGuIom8OOgmgrzo5KnVlnQDYYb5R8pAwuboAGuBeQe+Fn0p3CRH+s9uSx4et3+
N14jKJMHgC+Z71EHMQfDHd27wGKlZw8opn+NB88i4jz4lT/FMzLRlX9AMkffHh9EFsur+V8Mvebx
RMTPD1L727SC+y8gsYtNTzLtZb2ZKM7XpBFNadpQUc51CR/JGj/HvofB0P/DuKBLKOF748y4OkGh
yqEq9lIppexAmXzDw4ozCmRVfeYnYAV80dZEYZ5YwZvOxrSnrfRzufi5xpJmrz8iH40JOokylORH
SufowCw2+6lniyCHYRDv6m+5zp+Lx/oaO3l3Zz9vLuWO+q5p2q7gAwbwb6xyhbfpK0mBTXMiJq8F
89cMIY1vZoUC4QAIzFVhY6uU9Srpqhshez8t+/8RlBJb2uwhfomwHDFEkBCxJ/mMnCZZ5TxbqNmD
ynvXBCO4rhfDC2CvN/xw7sBEnm85iWFGTIapb6RYFUs6dOEZRSTpIoLKLDvWCRUYcUzNxkEh8dOI
skxkBCrDoSf+2qgIhLEr434Cv02o8OzC+JvpttDWHx6ck5sf3Bs49Ej7hRRekBiQHYudoopHwA2i
ErJvMqCmi2sfigmAWvGcuufKg0fkkuhbylVOCHRcvEpa8q394OKe46pSkYshZ5Coi6CXDOhmGxkr
BtLS+GDJqPoDGGLAcoAmtC9AwarVKfB9mSFBXC7KPs1ii27UNKw5/d8/z/SAC1ftsBPCXqDGfNUF
/DvB2mrCtlyGe8wjpRzJfJvbA4LChNqHVjhJPkI+1DvU8d2UFMjlDHsNhbc8K2WSSjsYN2rEsD0g
aLhoBXHYmW8SnZ5MBIVi7nLt3hu945iqiC3+1KqJ8cy0Y7x4hWUoSPSBiumfF12HlM8ydKyQFEfZ
q4mYSZuuMxADK4FiUbB+Bpt+UP0iba+3APXMA9n5WPbgtnsbBqYZYi98w5d+LQAp62W3Y9JgsuWn
+NF3u4VenNbQqSWY9Trcr81CkdRNFzX00HA472mUk6Zpg8395Sd7RWPShKGyoqasqNYRJuibKd0i
WeFFmlrydRbshd3tBXRRXloNgA2Hgkg1aLVDAtKx+rF5Z12WGVcMr4AZJhQFN1B+VbztswkKQDM9
ZdjGcsI9KgMprH2Z7iG8O3RS7zdfuroVs/woL1jVIcQ9G1cMwQxa5wWa5GLODcefmItgLtM2sr8l
dqgSaATPpHYdpuZh0Vgp0BjsGTantEOUUxvME70moM+MUvuZ9juxSVxKEjW22SlRE9bRzwxTH4LV
R7/UAjwHQnm1isNRL9aEqLTZl+l2/bo6e2VZlgTaLNi5t0N4K0MfezTe1hlRAEcBOQ6CZdQv/dRn
FM4xpFWn76a0YBAzxqdIyZGdxhzoWCDPwv0eGl3YqC3UKWgpxQZIhvo40YxRYtLigIRX+96RBzyD
pAw3czVpCakIOk0m04ukKoFJSxEuo5q4jyb/uRPLm/uLQcl8HENtF4pv2U2AjIVxtLDgYpVnlCB2
mGjADPb4zIiygR/iIUJ3XmQGDLXnNaGxRhY8FDJG8xC676ga2KbUKQJJ4Z8N/aCETnsyyeMwz1uV
X2ITga45KhxeMz0bKewtelNyjHsePKyjKdPl7ZZqkqoWPh4Mug7yP3mkR6walFgj1aX2YjaMXHR0
eU3xcRdakH0Uqa1dA/bF3f5xhp9fO0Kt1OCCAYaF2/Y3C8gSBRqfvmHMnVSz62/0NKrZ98/E2SFc
2Af/g4Jh/4sP7LXzmBnjd+GueghjfC2E5+g7Mq8zOSqdZDpwbRWRm7126xkI9lw28ELmm84k61s/
kwHXPu/vmTeimcXgCT6H3Njdw4eaeSlh+6XkS4kSP/f2/EeUIePmiCBYqSmQfMoLlRjyjHgWMGX5
cqIlu2IU4bzf7P9s90J2VqITf+hMzeEmpHSjRHkRDRFBhiQNk5TZEVNTCCqkT8QBVAV/uM/+vqE9
xUOXOcuCh10Igk1lKkTmu3vTiAoPLEYr+aUynpY4vY5HdEZns/pbinEcMoE/elwNlQigyieBi3Aa
+YD/Pgm1lILVaHgXg2Juv5DoOm/1m3HGY1qfh8Vs/1W5Y+bN/Ay2J5wr18KK/72R3+PhiOO7CRSU
3ehvLauZxrq/4zJCfxcOgq8LZ7EIddn8UuM8wnCmf66XmsWY6NwjpDMGrNtWMeo6sEvd7UmRLI5i
HvhqSwDzvKc1+uH+LNlxWb+GE8FR/LyOzI+2tsh2uvxNkRCdZuoTGORU79dqtOKu8RS7BbpG9WXs
ORTlQEEyHe+4al6LCOhc6noEvH2/PY/CqO1kGyuWBRvmST6xDPq7/m3SDq7qAQSBkqoUFbD6UxQT
dkYxA00/CZv+nIarSdvBJcjxEmg55LWSacRXanlkWr2pT6Ai2/5NzdwAvUmN5SmqACRyh2VQstc6
2hfxv2GCq0MtyfvZzkVEPFUTitSBgDeyfhG0dWoOgHUYq9GLrVxUTNUq4/ptjVthFflvAJ8cLg1F
sjQlm6fDejuitUo5ahINRdLJwqEb2XYROouX4MDNAoxgrpFGf0qc75mDm8F/Dz1EBHa36LX44bp/
jFN6umYW7rdE73i9ualYcdu5uL/4vt7nU8f1Lm0JTB02semtRSCMcvg51bdWPdMiumcaR07LT2zL
T6Xc30SyNQMBDlVFAX9XJai2oji1QufIS/GXIP/23x6T4eSms3+fEko0h0aa7KjXCg62uGPH9InA
imEp6hfk20y9mVe6RPCbln9JUKAtmEwE9oBXCz6O/lfLYz+bExiXs6IAqHnFUOpXNCzExLMvGSG+
ln9hRqtRRIAw53tjaO6eEtMsTv/zj0S0a7yNU4kyWkXZPZLt6H9rH8OfGdrL6Or2DScGKelMEWLg
jm0aMfEhr/fVw1/xw/SX492fjelAc3yBMF4mta6GxXj7toiZOtTjCWIHTyG6flsbIwNAa7LcWgA2
XB0lPSyDgA/3oXdw6kEsEapn3VPHY9Uf/oQZyB8ImbHjfAEi2tcikcwFCmXauDPZYW3aehq2oQQK
Hm8qCjldw2ree6etUlnT4/zgdhUi1Xf6k+MDgP0A/PlVEojTcgNOEemoWC98z3NMduolFKbaHHPg
o+kIbRJF7x+hSeM/XqcgDY/3rS5ZnGck1rk4uss39/8clXHO/RQ9P5w6lLsT9Aa34c5+ecaZTacu
i5HYYHKgCGHXoY43+VgdDikZDxLQyLxs/H/t398Tg0LSwOrCyh7ExmCs9IrpYUIhY/Qdm7y/BTGK
Khk9QAONgz3xA8ynGjZ+FTowrZkttDR54BGeC0tM4nW+K4eJXF7nOhFVSuEvRNu69ZsgjklEiZQl
aRhWvX/AMT3XiP1umF4Awt64fK4TNWPmbc6iCTYup+jf1mW+DAYmx8eL1/yvrE2BeTRJF+YxEa3A
DKjwiAuH6Q8tVbs6OooG9ol4AmusCw0HuhFfJX4zEjaS84UOziJzadZuQ1s3gHzotgadketWrYDU
NY8wsEyzUjLotlg9TX3jBl1EIStNICQIL1WVtFhZApnv+KimfW2SUSvbtnm21JK6xzv+AYLU5+vE
Na7G6Y4D5G895v6B+FJ2ZPUrzd9tJe5NmKqfdrCsJqXqti35RBUQZpbc/w4iiRlfpS9+JKMOmo6H
KXSk1dnrEAkepJrNqrYQbFg5GBXGOTWylqBEDiVm2eB8xDnpNUVbla1q88ANks6wIARt8JhbrkCj
jH3as70Ej3lKLhm6g2M0o0dPCET8GoW7l+oltCzNFABg31bdzxV5C0FQqw7/wWLuDEFi76fK68PW
PcBXqyk70tZe8mrLoi/44z1q7zIYG1T/A0hXBsMAqQNYt1kuIZfMCIMmDkhQhsO0OvACx5gIjqhK
i+JKjWGgKAyPlX0oK9/vkcDqrJewmxqPVdohSIOq0eBc5HZoDeYmS6DgXeDlx2AnRN6xUxSnE8Ox
Qn5oza/6XPBp39i4yoGCHR/m7CeZaeK73eYrVVJMV6wu4VTwVz27OzDnwByOLOjZa20PXkFLegf+
svGgpQhoCzwPlRXFK/o6iMdxCbrqPAtYti8d0Mbxq7FSwy4SAca7/kzcUhCFP/nW8VAkyczOdc42
6kIyyZO+PFtIPYMLqUToHZvkOWY3Zb6PVjaM1Xb30xkJmmFZTNCAwQmBFonONjgF+31kQunsbdJ5
5oEFSeAm28HipDCCUTu9LvKWQ9lRjUxJ6gyj3Rp18DT6vwV1KPYyvWMW6/2nqqhU/DOQUpIMUSIT
VKdhuOvr5MYppgquCQYw622fUA5kGMP8eZMk8IPbUKhlLs0ZyTpmOWrivkLePepEubFcgx3r6Zuu
09g8l7RE33d8MxU2eEtnHKnm/NTtlqryduvwvwuOq/J1u/rImq04fzRe9PIVw3wmUZbaObWKQou9
Q/xZcqP8D/0j14feshw5MeVq1bnIbaH0ncroDruR5w2WmjZpn9C/SnUqSFP70eSx78WHyfBa1D7s
mcqOlSW72qZ9ZjfKDtiNm7LMufeNDdXfPa8sq99QRl6hyeD7H3Ni7S7EwOM1oM/9kS4ElKQVxM1y
b3VfbmpDwbiOsll15Wpf9u3rqIvF2KxcF7jMkvKbyMQHT1UGWlSPi2f8Xa8WURe0frw4RxJrxxlA
7YlbWr3HvDQ+DfbwhsVZC9Eu1vAeE3JZcGZTGHuTOdal1Ytq47Lkx1pFiXQJiaG1X7oYGd75MlhP
JPXRN3kVRjCApNIg+fGHq8q6n1zjblAXml/JbWNK0S2EBtoKE/ktrvv5wqsf40+qAVBEluHZYHoy
jQ/9HeVIVtHY0bHPSB4guEUpztmaZamA4o230n3HZc2Jp9QwLSv2iRSZKXCFzLsHkeYfmkwAMUCm
xqpyrbRnuwSD+hTllyPzXt1fP3+D6yGr/LgHEWqcZi89Wj1UrjJjup3YlGXsPTnipzJKU/LFdrJ1
RZyjwRQk2g4pWIDjfUHKYe6VhG+9pAY4++jtuGpkac4IP0dZ9d/zxnoot/5Xus8QChLAo0RAqtmI
/aDig/Ervlf8o4nakySLml/7BtQ0S0U3JBbTo/rrSLolV7HBKTqKOvpS7oDahDfnvb2j3f8VS5Re
DPA5IRcanmQiPMnChncL5eTisfJ1qswoJYhTjWNkTOodSGcYF9kquP6bM5+8Ln8PHEbdxdAtm4Ky
bZQNT+zM3mdCqaSAz5SxxEnR/QXpLSak8L0WS6/1ztm/JJOK20ihM1SpqnY+7oFIN12uUVd1lLb5
zDtFGqn5s1SVe/4727ruTFr1kZng4izKqrFYEETSWZQWhuT02gIaefwZNhlbr42pUMemFwD6WMbZ
HZ76iEOFp9mnkn01USTjWHElGFAMYojVSMvs7xKuZbXeQelpGlx3+ghfKpgQJwIYkau+2eK+BCfx
kQF4DVF7zo8XuclbDkGUqN59GOe594x3VwU6FwIfLpEcf5zlzn8T+hB4RwMl36J6w2Ax4g9y4+Ua
TEmK4QofP6MLh0K7VvxyUHCS9PuIaNiLRP/IXAzUOVDUz4Dvq25PqwjL7Ip6ihMneao2GGiNmKw6
TUsbNFR2M2AFDOQ/uaKIvvnPJj1ZPQKKoGSMqOl+xjlC9dI7htsdX7sGL8V4MIEWv6RwFOqLzpMj
lkM/eC8DjS8lCA1fEJPvODJNQ2+SuDbHNNEpBiaMZ0MTJnQM9CwVNTgq1RC4eNaH4Z5d6YsrL4Ei
kao6RdNlUiK47SY/EhiXVntUy/zbS4/lMPYTQ8m/KnWEbSiwm/uDUOWE6SaaQcn2d+yl70h065/T
sttissqynjTHPgZCBmAuuDDfx3PavmKqmJaTlZK63WUMhZZAnLlCmAJ9U4RnQFO2MRGwOuk8prTD
g8d1uhEBX7S/IKT9MUNOHCAQe5eSt80kipGu9DmI6Is9XhDVUga9WirYfuth45lO0a8+Unoe/54N
jNzKoEEHAsKWMUAfRdIljN5Asu92t1dOFwXw6GnXl6S2D/pQzhTlOcgnFtvBbOAFAxFLDzI0+Ecl
lXbiAFGkIzNJoCixFwoMDMIsFLHjQMNsj1BADA9ogejpwqBR9cY0wo0drNJL2VbbYSsESzvAbefv
Pe+RVDZ94G6aD0tDc9P8UAY7YZcFWFqj/N3OwHnJog/gEmErhkKei7e+5Dn2vn8FqrepShMgF3ZR
QLKpQ1K/OYjQ5V0+HLaD5HQHU0L1ZTqmcuoYC+sDLrCVjSFo5sOqdU1uvE1noxO0e9ITR+ESRI0e
4DQVYBzJDSVeIiWxzoLDxUUg5dZTZMN2O79lZvbFpLdBlzVT2YkC37pIikzqTOWz86FqrX5MTJI1
NyHO/cK4/B2vUk0/yXGGqN3Y3WzRHBECR+lw9YSyyGwwTKD1SuAMHAVi/GGHiPpUaj4QgqSRCgoy
LNi/Nycns+KsKmU5PkHtvdnL14cDDjyU9wSTj73nMzzyTbv7IaQBe92PqiRLxWoLIhoy7kf/b+K7
pbQobTv79xPEI0A5WG9w/a1HiROBBFXN6LwU1sRJLOyFnxCH2kE9D+g2hLuh+EHumIGgu+ZQw/pa
lsqStXQL8OMNVi4Nmv66VyXlmpDgN3hFCvfKg3xg2CqpUAibhoJMYd9wAFYsQTFRZfSjKIlB/jcS
LebgxdkxT8/owdnf5ZwyjNEJqd/UyGeAM1yPecRcapGsyJJXkvZPBH/4Pb9m8e2jheKEWQi6mZg4
aSsM9GswMdpTTMfofF+mPTKTKoPxkpYLrV4vkuGDTizBhhMjyxH2EQqpb60IXofd1/l0uVrBVTNn
kHkjRhMMfgR2YgDsRxstJf19GyXvfYxghJ5aEF8BkxQgiTI9p6VvLfxM861ACGxke6BzcHIvIQIV
VOI6lwltH+tOIwm9xPhyibRHcv7OVQxWRhJ9fq9JkcKGDs6fmHWsd3JIn3+AdqAklZLEGU6a2frR
kRQMDVHYOv3DphLF/IXg51UhBnuatf0XF4zeJg4HsJiaemcgTrr0RFTRpX73TeRk3U5WzAOIPrNB
/wKwGcWh6BS832IjlmjOKShpRsg7I3l+ymu4XK9de8Fes+KLXfLDVpvHggY2DG+CUrBcDd4dwzWB
GencBlkVpQZeN8Tt/Dtm/MN8wUd+E5FAdO+OFtUJBBfMGQE44hh7OkJYLEPM9mISFNVQAloLmaU1
jO4NpDlMKR07pyMY3DQMTZN4P9OHRVIFn6JQiyLQBYvEmzFOy9r7dW3CtFEchVk0i7D5bjzjwk4R
wVzIqcWMmChjZ77XeQ6AwZs3E0I4D10E9xaP1oA2bWNXnwemv+K8xVmfPWW+b/L5pzzJpqkZgrsF
4hhCtjOpMm2QykqLUX2kPf1E87Q9IG2CtXJ+ER6sSPBLA1UQoLfPTEdUko5L941X1ZU/0KSeBYWZ
UbkIklBqPwrm23+6PSnfjVm834q/EMgXHt7I5PH8xZSamtPRf5BpRvO9GEBBBELphyC/8SDQu71i
7ygZPzakOn+OWfy7pYv7wke8LdVNzTCCWMVRAvK5cYOx9I060NRwtT4kxN1hO97LGqr7rB7RqKUt
pgjCCkRJGT5apFDusZDjrqAa50jZUkAwauSrHl1ncjCrDzxouU8gyvX7IHTc3DT68FZ9n64iixjL
Y6eNMlAk/jMzoWdHyPQAlfuIkTItzcKqssglU8cJJ7xHtrXr8hiMX2RUn4zc84JX5YXkyxPpedSu
Qrt098FeoMRNOeYiVQ4xckDJ/igKz3Tv9/cxf4a4EMVoCXc5weBUPwgPxtsX3azBzjenc6OZUqG6
JoIBGs+iC1eRi5pUDkOgsj6jCC7ATpG5Z6mS7K8M3oWMFnusfZKfLuxChTsNPnpHt2E0/vnuVLVN
V2tL1PX8Ev+0q5jy8aEQsHNqIturejb/2F6E0s2V94DV5BjigSXfiDbHif2AR0G/47u++GF7uQdJ
y9TX9GRnB910KDkfd88miwh0jFQ/bgpWFgMRuxZceDbRCUdCi0/I7Z31jqXQAqUHetCqZKGKOCb0
A5fZFElFDVPFsC9jyVicW2O2wpfcY713Mk9z3UdtsHbKPeWHv7OtSQ1ATjvYy7OlRRfaMdxiLZ64
5ZiBEmQAerTOhfkwy4p8uYT1m8rja0q9ViKyHA+CXCDXs1rhM1YauCm23JtKF+AUOvpb6YR22bDB
QxgY9QInOvjNtYgLDpLm1Zq7iHK5bRZPZqzp++EkihkhfO3qvlbDNDlIC6fQ1zy4K+LZToypucZr
OKOqRtmHbVXwZoZ6sT9z0dJGMzOmiGMxHkcouxYLr190Uf3d3SMIQBFsHA64q9s8mDh4EKlyNOnW
WkCfhO4N52UcFmIcQBMKEhPnVwE4n/e2apEr7fFOQQ1M8CMmj13BChrhNOjF1VD8IYIKt4RRunNv
YDzOoU3fqr2OaxcBSJR41aqnlZy4Ek8IJy2VaGl/CYrLLuzcUj4wBZ67edB1tVpNprmKjo0gU+vC
GbOVefPSkzr1TtkOvU2AnRdTlDl3QdvsK9+yqTedELCgllaBc7tt1Hxja7v+bxiItUgl6d65xziL
Q1u25ceurj7jVFSL5HunUK0saqlUfgeLPje3t9vM8KShFWU4RzCvfr+nc1sS39vq4smlqNT0r78W
gGn2TCScjtpotpoo2JE/kI+kbabMajNJIbssQivhtHgqs+jEBBwtxBQPyEDZMFX8cfOgsVEBq603
wSwM57Ps6calhd/2cmsFcDnB9TPD+nNjZqppSwy/C4fHAKvbgiCXx9ECdaxDTa/0kyU4Oip3TuOH
lt2OljXahI7JFYGO7+FldLVcp7lMab3WuFLWlaVmmTXZN1eXmBNmO5Ju5h1w50vGX8nSwz4NGxqt
MQkdD1bKXnSvbVH0tzi3/c7kbRa0xHnWG6Ae3pkc5zu6pMkZtF+kIg1fjSZj6MzdkzurQlt2AjTd
WopwFTXopJ1Rtl10SMZojJO1xFw9x+YVLF/wi7chf0tp1jB0UfIgL6JCwIMHtLlc0/KFF7xvB6XK
o3P9RPkpSzQV+9mZBVhoM/KlYUrevTsQzM4BCFta/pnF/1FTCu9RxsZYzq4PBtLrYIiYKuB5msJq
1g1RJnhj6QHbdizTxC/JZQJGj1btGWbCnOtjEFBTGNYinngAIBOFJSvFn5iSyLdClrCJ4X4aEmwj
+IHZcYn1JEgj9uIc5IiDlzqaXbdAEHozhH4wLVrB/Bb5GQQj56T3whLlCp9WuvAVlPHGhh52rZI8
aH+VZMe1qYmJezo2QS4s23QwmxuD6edVIGCk0uGEOi1hgO/73n/SybIJOzLRh1BE5KFd7oOG/fMi
5fJE0veojGUWcSI5UQrR4fKZJuSTi5NmDye0L5R5UzrSme3nTRjLjMOond7730iAFlGRvyia7Nyw
Kwq+6g4/7TMBH++WfkddSck4Ee7wNtBb+RfpI58wxlvJTxj6D++B911uMhUXwil33b80EOmzJBOd
z2XxqzPrrWr2RxZ8hkIUwxlpiHBqpgU9M8Hne7OiegxeZtcVTAJWEm/MDBWOMKCnL1OcstD0IEXD
U7TeRMm+0I6vvUauP80vu/YBP27Lt4Srd/H1wiaYq3ASocoxILzIhdFIZIRNBTNKkaWNMhKZZMBA
AqIPNP9AjhYV0RYfl8nbXNXh/4bhxJZvg3k4dPaWdb7sMTLCbMuselro8xw9fJY3DxTeedWL8lmz
X8LNHQOGYHrr/bRyKR58qW3ughVsuRFZg6v8pxoBuJQQDh250lnpeQfcJZkUQ76Ba3g1kL4i9JGk
fJp7CqxPLsw/hxwqHOy0YQ4F8IiPEOV6fXilbsAimTjes4ECIDwlcj90JA//A3jEvRkpm0HEDK2L
lrQSKTJQW/LqdGYC73sTTKFH6tJPyT73ahpieYmADPoBEyaMc1G7Rno7ZG+v4pYsXcQlS/CPozKw
j302rG0wogA1m/N9X/JhXe3rfQEkodOWs/l4xEwsC62lLIvBBew50XKwb+BnYSdzKV5e+w0vwlc0
Ubttj0beylgT4wXKubQhyRYHybwQGAE5rJlmYGTDFv1X8HxKqtky9tDuq5TfrgWxr2TANK9AN2WX
pvT4iknt1HrbAtguBIH6AB+z0bxSEbFiD5iFsQR46NlKTF2sSRoMS2/azyld0zy2Rz1P/2jU2ZLD
6dYEbPJVyqT4NWtfJl3Fi+u7JYzzy3Db5mM5fgDTX9D0Gw80EQuRwU6ClxWAxaMzqTUdY8XCLcPI
wTUMh6fX0cFiEQ9EAfoYSfbstZViXrjnwG6yo/HRmH1STBf8QUVoljV2O3vQ0lB2N/Gx528gTLkw
oxxW1ZViVzLGQsXeuhS0calajB/czZRnZIAvk1NIPhL1iNmYadgoLQPdrE2Au1dqizfMZ9HJbnhD
W6P0C8B41xrUerf3OLuj+wcBA1FupV696LTxU5rFNyVhNXZPaxLiarN1pczkm4KHu0eL6nsh5BtR
YvG7WuNF7X33gC+tr0dZgRdDFXCz1I9liiDR112Etu85hSbNkZ+7RU+W+XC7rzzmEDom+Kjnk5bS
oTns9kIlS430CVGy7aVVMSil8wSVj3teKQzrb+tQvQZcnarv/atyP+JsoFp1Wj01C7d8/irS4Koe
BMVz36rZEWGVgpJpXRpeqIpOm+kdS3IoEYQGwsa+Op4N1BbSrqAJ7Gi4kL2qasH+flXvDp1F9ZO7
W3Dk++P+p9ocNatiRP+NfuPrLx03yl+0RohwwrN5WOY5grC7t0XlcnSoAmV6gLOaWKqToaQTh5WW
ahrDMRkgnhQMsSLfR5ia5U3O8TLUUvcuuNRXp6XDQJBTqEnUwEDUPslORxuuhBlGGRBS2n1qJw79
KtvqxY+J4hbmnmpLFmJumtOCRz6QSE9drqxzbf2y67pCkmqF/wC/KFUAaWqeKPNkSUefi6M+T9nB
Z2pI/WQ58iyJP2NG4W02kUzmDaFtMp8HubY95NQr+4HuE/aFa4zjnLxPL62kTK52B1KwMZpe+KO0
hsNng64wdFuEju4sSVQojxV3/xtP5q4mA5Y0UP7sFtHzk+FoAQKZY5ZK8eAzffaPILxf09jOLt9s
0KeP6ZExv3e6ef8Smw4zcETNSxcKjVIKdlEPOqcrUdg9sv23f9aEmwCMPhnNy31FnvvOk+8k8YRv
J2LcNUYFhm5kyxzDdlxB2HGvbegqithJ2klK14SV2V8HDi8RjGoe3oFsFF2Q8082hpQyCLbeLcER
s8i4NylA7h42E/BLqAzW2+T4/pDkBO7rH5MdwXnLmQmuD0CsK/1UcjXUFprC+EyVuf5a3e8DjmC3
uJJRpfubcL6qfM74ahEZOhpfurZz1zYZJCZ2NXJ64rWkSBajuFthJdrlozN/sGhMjiju/Wb7dkGm
+a0sNtbE9htftjnPQZ+NLYX08W9clKKTWrbB5wOO6yo3wYLHZYAF8En7alfTvTibrirws3AcCR9/
3ZAMyKTDZCo2LO5EJlavTz5Ff8X0heZh4a4z7gvAdJCsxH/yNGkH+WqKVokhbYOWwMX324B1hcll
S7pXt2iz/D1Ru81ao89aHV6LBDaAya5Jvy39iVL/BfBCqvnbMy4FCy9M/7I6iZUbJFoiKrvIpeFq
j0sUhwmrFj4UwOnM6eB+KWQWVZbNfSm+AKMO4fmOQzPLnvox+uyKEtRsV+Rcl9uKAE/V12vWZEZj
iuW/FYWaa39aqca17ioZjYakwz5Om4po3duT0lUEsWebxk1jFAGrI/Km0EN7Us3h/Y5wAsD9oatB
Pl2WkvHcQoHuwRyhvz+mPtw9qGS/Yv86mnc1eZ7WivZsmcvBv6qVgZsKkgCrV/Bxz0Usd5mRxuoD
4HP4u3pUt0BgxeZTzIxMWTAajPeAamGZhaqI420+XTlPKMWy0JwNrbBZOUn8GILW1RRcWHWxKY/m
ygHV9m7vBLl1Bk/HF0hQiGrtmXzPlDDVG3rY0fE3f1pdqQciU8whJTG29JPkSdtBN93tPgEyJWpV
76jtyOVRRNNtQPnqyW9uDAjS8QoiczXQv8It6LtT1mVOIvmWsDLqYLLnrbPM93KD046vztIr/KiS
c6hGFvb56FEC4E+7cTwRlkQo24B3N6zxvfAWxQa/Xq96jfUBdHjlnmnJw9PdHJ9qmVyP3DFTVhA6
XwrJdiaj9lxIogUL0avXjRQGiNdzpfllx5KuuzSOpJMXJ0fZPtbfuLQW258DDLAutkdyCcuPNeog
3+0N4dp7JlPq33TzeNrjxssLwIVVDIqniPZ/1GOzgk93Vt30+OkBCJB1QReZrrpUYYBHTqXEm6CN
fGRhzMidfW/U5+NXoLI7/87S1SxRIaCkFuQHoVL0kome6jV5t8dxj4MfZWlIWlmpCC4Lww4ErZ4R
tR3sP474+IOaIm+9sL4WFBd4Re/oo4VGeCStMJyXxsxqc/emZj3iQvH7xmdYX/m7/YWOrNc+Zqbk
03sCZz3DT9lMsOikKPX5fpFYh5UxOI8TclmQH05dxFicLKl57ejZVdwvnvocXfjHCKWy48j4OLP/
dMF+BoA69QYrJ9hEQIL5gtJRmvlLKCB/Vad9xHhc3zOrJupBsOYt+e/7EplebxpyDEF5QNnmQHDf
CA5CF+ErCOaMt0+/nyCMIZ7AK+2bYrAvHY2q2YyHq30cC9e2OSN/xdz7pjtEgtsjUeFGFoYHrac1
vFgUF64frPsfdvzyozfGHjh0hovmqd/PVKVTBpvRpjm9otR3JwO9pu0KI8lhwFUEEXjGsCC4Jtng
mzYqTs7ifZunrO+2s79exqvegn0wb+FMVePHtnfxSWjD3Ea1JzN9hVTA1p5gdDKUDNULSMuewvvr
M5SL5hKhzJo/LCeYbFeIbDSf3VBTKiBmsHJf0OJIU4ntd4vyU14NobH2+u4QIcKQ07TmLjHW7Aj5
ZgvrKJvimxYzGclt0SkFybzytix22laZTyRTJnWPNy0XiVTYB+bgH7NBeDCFVnOurdciYqMIdRmr
Vr0pVtsKIlRKx2RUQmFmY752FAUMK5XVdyN+9A4Zr+uEvotiVj57vMwozr0PyU7+ehcvy0abCYOR
aOjb7lWgegB0ccfcRRIaHluMJ/KgD4nFfevlVsHElnVWDBt+0oYq+3ljGk5zlYwMUet3er+cLbSo
NIWcIFcA8bv4oIaWH2HgJHUKiNipgPoYVsjZIuQ6jzo2VcJnAWVC3LarplnNE6J7TqP6oyhpJYwx
JBmcT2zsMDUiiMf1VrdnnkR0e5XyYBd4QSBEm13NvTMiaFQmou/DTBRWVQMcQ9XouKDc2hm1EQI7
x9YQfNv3uaQrFcjCN4c+q3uOYeCTBAqLAWA3AmECS6J/nMMWxDJ59E5AWVx7fqaF4GVu5rvj1fRA
EyddsgKifXbw6EE6YGwilQJDRcZbfM6pLFQiQ857wf6/t0Hqmew6qlXfcddnrFPfnsMVO4YSDqjU
/7VgvrA/+HeEgRnD+mQk8drPcQoemq9NTsDAkWKGKuiwCQOFAIRH+qQnhF9i2wdo3slTP+F+9hDC
zR3lnkEpshDEC77qetuHSF57tCtztMhPg74cOQjK+2n6xOXcfxBpyAquhN5MONDvOUB9+2lUQfwI
NqUK5ySrGNCMLEaN6ecLE509W9ISPjb7BzLkSETjpDs+NMRt78ewRevekjCpeBGEmB8jIU4J2mp5
OXd0/KTo+BYvwa3zF+RU1eP4tMjyYZkScbqovcasJzxsD1suBUQnH3rpV1LiZBIcqdImCjyrOYoV
8zXa392SK6H7MMoC5vDn2J6/ZgoXT1tUkD2n44rc7gCetJ2ddaaB/w2L/8PdR6gvCdCEtQTT3T4h
rsdV6y80KcwnbzDWiY9z7seO5CuM4pOD68XciIH57RDzWCwtqyrFNYienkYngvGGMzVLW7utwK5l
aUXdVqAlCstgrFLuevc333uGF/v0cH25pLgGwdTb48p5TIHTjFPmXuB2RYu6f/+bsmt+XtTKvu5+
shbF73Mw2DprQZAG/Q2IjLgpFeK8iLliAqbEWRbcpk6L55vPEfhl/8i+4KrjgvpmrZXGbVQxQrWP
KEQX6Wzsni39duKXdrUMrHsHPJ+JZ8OXr1VHT+mdoM4r3TK3tXf3TSS2w+cMrJsGkBP1cWX+UvfE
+3Je0g+6KYWY8s7/pnXo35VTGmWbojn+NwWw03fUqdptddK+U2UgfgFpfVMUlFMxtT6WgVNj1IRt
tXq/ZVJKAuHnvP1fJ+r83gbaMvMSg56R2i3mXG4KS9jW5QjQpOZQx1eKabWfpYJMcVFMlD+dDw0z
thALgwajhyNANcO4gLVRKB/iGNtDfJJngHI3/hSxEgfGQFwa4cynPvnx+RRb8Bz2MoRddSGuyJ1F
6GS92sPdR52bMJx9q9zJuu3Unb27ucdA4ViWUdpLemcDWKgf7wFLWyS7qehZW3KG5/U762vOAdzz
sT+fAQN2D6WHXWfguuPp0+/t6ob+BI+oq57yeSIT9/Qc/4X0a+kreWxqAhWqbRsHLQSba5MgNQQ3
Us72HHK1SEQ3TIeSew6qcT18VWJkZ2io26fAhPqwHMZ9SRFMq0zmm1q5uHYMcJS28rVzV7PsS1MX
EsoW6L559BzgcySgDDjEVZMRweIdWtdRVDR8Hl1HzyXQg4J3MWqyI1kU9oRT8Wd7hTBkCykdwvVK
3pO9gehsQPQYvZoguyDRUjYWWUMEpfjGYThZcBShpE/ugidTv9ajyeR/XdRmGuaKPxdJhyTQrlQt
n4TFgnRewqFGNfydxnJr1w6v/fwK6N21kkhyF29srKDAxWT6WRa4Ng5dEBCv6jAtjInEYxbzI3kH
JYF+v2OGfIODLseuHwqOidoRFbyHUDW4naHJ3IrCqCbq4wMtQTQn3Bu2zJ2X3a6UBQna7WDfKJw9
m+GoA5yNIJmaySZNNH1eCBevcfszUumbqwMKd2WJLYtn2FkA0Ww6YcCThCVWhw2AgNYrjfx4GqMf
Ykd2k39wyp7KItPSzje9Hhlz5cWmLDkc+ACB7ut4iYlqWRybvleLrpufu8PQUL4fR0NgTuXFtL5f
s7qR5wjt9xYCdtP1IQCoieoO/VvciiBy8W4cm9Vimz2IB/jiI1iKWScNKwjqGQabzBZrtoyK8Pzc
Y8yS5qmsqz1UDREuH65IbyxwMWDfDJeJHft/ReS2gtCwiQ85PbMVX9J3pikbIycFoi/tzy+yFACU
HG+ClBnoGMwZEH9CsDwheZYS1jH0OBWpFu5GGeIYcGoZ7KthJNS2ErpXahocodcJgldsTs6G7ekU
AHNRQTrpGraHyEOzlx28wu5g8trgh0O5PraJZyPmBULmK9EddtABxEmmQanu1q50Ml2BeazV5vST
dVcnIWwpqRP6fJ+LZkw4dwyyi/ffmJlP7p5gBYkwRUEXsYUYRzb4Y/ANn8UmV98usmb6wt7hd71I
hybXuIzKna4Cl6ZJ2x8UanWFAfKTwcxYQ+ql4DVO67tQ6BFeAkrHTCByTwF3xOEegQG9OPkIWQ3F
hHBFJ4tQfG3DcO+p5Bp12HvQIR+OEosioSd1O2re3Blyz9ACcguEj5ZiVOXrEYwXJe1RRpFTJvEu
FcZvk8Gz7uczPjG4no32PNkMqrVNW7D0iFolttL9JdRqM+jqdnxevj17QvBKDYAKJliIN+/X1kQ4
KZqXV8S7IkSWn2vqWkVX3yq0zwkLXFuYFdJAn2+o71r2LKcSVJ/epowQ5z+nAtCzJ2ePBeuML9no
ASGCEjngcik8SwH/lCNZZiGfhtrMaVnsJfsmJ8DgMcxObSHV8wo/9DFsZiukwVgwB4hLtFTUBati
63G5p2Z3MMpgYmcqm/0KEu/EYuZOtT6pc+ulHvmdQOKvYnOuqsg5WI6WOmfI/C6BWNCKNsNSE3By
O7gKjFbBqYeSI1yq1vn7LOrOPJWAJvLIP4lTeuEY/AW62++rrxHHLH9N3uZixIaVVf/CSpBxgY6r
Zq32ZBJ5fupTV6Lc/4Oycj5WVLPyAjgpm42JpdbpN0GeFBm2ah+2CzOO34f6k5WKgQiWQ3U3q6Gh
LHO4TdvYPUVgspECDWJj/pN+8FzX/LdK0mPcwdMxl4tq+4IXIg8ULbV+1v+yGef+dhzhOpu6Eekk
WQA2Zi5VKlbf2DE3iPJA41GA2FBZwFecAGTN8goDSzb/zp3LFbnL2qc+65DAJ6aiMcFGtJpqW4hE
OB3QoUtEhLVkHgWnqmSzj5sK2fnmZ6sIaH71JvfrmPFuwZmBE+hvEDp+G071Ow5TDl6WV+bRNMIK
NqbL9zXIe1jqSgRGv+k4ZRwL4LlJD9+RsFAwqN4KN+JcBcSJ8BrIzhaTAYu3EkBaMHt4/441Kwer
XSu2k1AEl2RrrUYzL/6Oqg+2IGZ6M7Y6+YNdb+getPZKTpEE+sOqu4SjgWsyCSe8OYbE1FI/0VjI
/ZJLYWS1wGlB2xQCH9f5gSGOGnER5hKgoA9jQdpVbjeU2htowlWOCrGRVGCS+4ilJuP7u5/XW0/g
GocJnVjUWMwCU3VaOgIZ3yHToH86GtaHfDRGark+5zQ4fVdIE8xRN7cAsws/7POMCh20e2sciBAn
JbBw/d15KnbpBHHVmTXpTfSI9dlYD8Bg9zW3aPykjku9jvok2ouUv0TxArr+dFOFa7+AcM9WyHZ1
hvCIKcuYhpKOfLrz1i25mlK9tZ1nm5ArV3+ggpoVzwIV9E0mIGXtbdr5FjcMTm27Y4zvw1e0ODje
KGn8umkmiAP3JCWXB188r4vy//gxLew2xdrIMCUiTfXg7caV7L+bVhJN1lYYBPrTuKoH9ru+IwYt
poMpnEm3DwqJCRHPZ18HAfTFdSb3GFx4UShJ0UF+i/tV1kbRsgC0GLcdeI6uAPggqe8OWMZb8FON
sQQSN8OCitagy6J4VxPNMj8dyTp4T97S6GOdWHbdfl1iptqUPZdfmasgmhv+nyOzDHoqJG1jElbh
oCSOLDS3slr4xQWqGGR3oA5J+Oc5fasSsCb1KsizC1Yh3gcOmy186sjhXIxiOeUBew6WtG+U6aXX
i/0H0CeSicpXLntJ3E0nmKeUET2ushJBdqko2LebNJWxUQ3Ar6Hm2BhEcu8ZRoSI1or+PW1KB/4t
uJmZ1O6tUuFdwPo1k6Sh0jFsyb81tOaxHClkbGmItpBT6zxR1HwSMMqpG3o1bZuw+kEOGS7KeCoM
wbWy4tZmPJ8pNSGLdulZXTWaNpIAgtqSQi4CtROLN1+aeiBToypclISTL1TL/uqTojcX2XrTRYyp
x0ffmYb1nPbOQnfQMI4BVtjO1t9hOSBOugtGUJA4bSa4JVFZV0NUx+l7VlI0jmhCkikfXDbP9Bn8
DWxJuEsla1lHgfUTE4DBiIlnEQeHs8Bw47EIEF7vjgB6g0J09VUKPlEup6Y0EMgd38XJrnp0BJlm
EI20jvNzYV98lkBef+TMO640VMGAIGdRH/47Q44DZjQnxzIszPa0FTnkDZ/LjiA4fTRW0qFugndt
vNPqoumdYB09xtodxlrsJbLy2eB3m5h4uc5C68WWDt9IQC0EBl6sWOESxMEU0ci4hp4G79Z3SIUe
In9uyAv7TmksKwG+e0KKSjw/dp95dr3iLnbgqmctIdCTozV2VmC6MINF0KlrmLMUaATXxhA2KsGL
D66eJdKvIlsO8pLmXcPJEzfWNmDHyBsax4eXUAo6b4/yCUhEEMgSmhQHl6CQp5un2k2R3J2KxrwU
5PsGKU0HiDykoSJ4Uf5e/FjxQ8jwzbizjotzDaqifSqaUcJ1C/m7EseDxImamLMXy1Xv+5AVbeVb
ppn4k5fpV4lmYw78DL/1lPiptbh1fKPX3Kr06DZdRk1GFFIExp1LKAb5Sq9XaIW/AOqABOihnxiF
cCAJ+wPp+9kC8qyx7RebJRpA/XVh0G++DL+Q/wusfF05GzgiTDJntnN4+ehNVH5qUzT8e+qevhHP
hXFVoPD3AqnI2dUv4Lva3fj9q92//SqKf8oXlCytO+jLD49oPsKYV6JllDn+DhhH5U8BWq5KjaQV
PRiXu/vpI/uWaTfd0BKXLDXXfVP3hcXziigoqMb8dSCY04sj7AoQhDb0C8J+2KeFeabcu2ujr1WT
KBIlLMngBtHXhqe+StRAVa6PRjTB9LkwCOCnCEdHFh2bnNWktmdxxrwu4P8+aVnXlb6Pk3U9TmeD
Xr0axkOoBk5Ix7lytjny42i3BGHUlHCCOXwzp4Hd1fj0ZysVV2z/TnSfBiA9dLsDw//tbcTNNjHZ
2lfuL/A2pL8VQnvx4De3MIF2cwBD0/Iv5RzrgK3iGjHdwjLsSL9rUZcQwMmTAFw0a6R07TYY/Q2f
e0aeTzoiYqVfGbr5HQ9OVPJs6xtIVkUy6wWNhKh19YI85yByhgj2uNRTF6+YDQF+78JDUV5oytGU
jQRcmLwngwsNvWj6uuBhOjjxQUO8SksJyhNxCr41zUKfbkGuhU2g5Qxf33lYFTJE9IWvUtxW63AG
VyZ9+bk/fAI9u/dpWIg+FOUQKXbMWFTnF9XtgghCzO3Rb0MFxIHzkKvaBROL/radh6bD3/SeUVqP
1tlhdapwWDsRzRzVmvP3CtqPR7TffXVWqvaWlqb/4Rm6om9L3vjcE6Jinu23YWuKlkGFSgIeCZL8
BC7tS9gFXXSjAhuVXTtt19wAJpVJj4R1WzlMjAKK+jFrfZOhlS1oRhAJRWyXFWeH3qPGEgpGjxzB
cGnHulzTNXQzwyiOhobB6djpT7Ldgz8TmowzXA7KjreMnFqzKNWeGIQTm71b9x9OKaxtyFSrm5uy
7MuqXIueMsszezpl/0kgAb8aQrJH9hEzul2JvcfNoMPIZn9N72SLUVrAK/EaDQrmQh9Y5bP+NgAn
SLHLwdF7j6QybMZ3OWnqg8xiR+2tnJwzabfYCE1rDpXv/W3cE1HEc+UUGxbmCJPy96c22TjS3jS8
dbtk4kFtjGVZfckCt346NmdbaixqQR9n38R4/mHppMS2zvRnpAf2Gceb2YT0I25pVoLJkisHopbH
X+wihaUhqLCrAbyImj57JMxgK3HyW/8otYQMcCSRztDl9mrflovOjPDNflRjQjRJSIdNffFN0b31
SW99GNbCq2VlXdwEAvphMg/dRLpE3v0YOOZJVHpiJBU/+vHSqBrtuwUkgX70JvSP4/G4Befn6Mh4
xQcsYyfxIFm5WaDNRCzsMX++MciCzgx/7EyHwcO/RONSChlkx7BbIoJB0jZTOX/1z5LYchE7WPJV
l15ajvCYUPdJL3olfxxbQaAv2gGVNZNTlrKkdf+Ns47ynCwVaVlXjqWGBsZyIzqwGM2SQyXRy2ef
uMpsiaIqY3aNWLbKCamQYd68HPHUNS5vJNZuaJhMnRSDGJLfb1drC+WEckuJa6n9bWCMMMYk59mv
qNIHzPT4ZJV75vJ8RtKiQ478lzkFZpFGcqCKt4AEmkWogaG1ze9AUTWgh/0MhFKOns0XqPo/9tIB
wzilVeM3D9fyDsX59Pez5rdMRGEQbwZ2BxDj6Pm+zJelMPK5DSRgLYJP+/+EIFDdQ+OBCsQZckFR
pqVgjzdxdLyvnPlezrIQFrfRw769+jzICx1yHEJSVSJiEIah4bjmIUxtQ0i8V4XSLZqXIwUKslcQ
p0/AA0a+mQYXxJDxyQTNCVitmwy8mTsHqGHvwmqUVrzdI/JDV73kvY3dW2rHTpfewv1qzwXAmU3n
bpG2qK33ctJzA7SL9nh46EHLCAphK/gCpPwI9Ul+pOqkfl7eYwGNRrdMgOp6A4gqriwzbiLPmncF
OVPUiGwIKrak80oBpb3gDkeVDP1F7TGN2K7TB/sxQoPdAgHzcKZHEadWWt+mZxCO845CoZcCuesb
iAkXZRDM5mAvQjx+bQqbXEVkpAXVNsHPNxRKm6mrEpgERqEor77DcNKGPbtR/wgnUx7dVCJQelMz
wqrziGemZlS6hQWSlh/AHJFDAVHc16+INkhX+AqrZutUQtVvVllAeH6S3BQ5U6oEa00dbT1LSxfu
16BI7BnJi10/YFePoUEYBwiEdutwJJQwR7oJK8yIdblYFrSuuKDNlSb8bP7HM2Y9im9zk4IThHuv
Y15V1RjIS4wQlPFwYHKRVsBMD+rg9bvpIA/G5k///EfAcpOQOktk8k8KlpxFefKkz8pGnixNLtDz
1XituzDiiNbIPc2t7wZtilhEPYMmZbfR4kCHFxou5o/uZgpCj41zf42JvU9F0tOff5n/ozgd+FHz
XqFr6q3xyfVfjdRTCfOsjiGbgV3h03zv3HdlgO1uV3QfViJImbkzIw/g2GTO8Ll0pOb2GsDUFpZV
dO83iEB0ueFBJS9TY3YuqIVWfNHvjgrKIaRHEx2MdyvtRV66NmP78+0K2C27rvMgMSyHtdwGOY5v
DGCckmNDJGSSv4ZAaiCH6/OC415MoMk2uVGaLBeK8yZOE02/qOegoj1o+ctBD9WmQYKnpnmFcB28
SKeeAvEAIyvWHD0bdIhGUW2ze3JjvfUMlValWXUcVf3hg86SbkqW9YKk5b8zZh1+vt9QShU480kb
2/ozVGDEDJ0oYtNiL6WhREPDl6RcRgd9gwAp1CGLE5L/22bJrYhOCh+NnaufdRwfIR0RceS0LF2n
qNILO6jZBXvjmAIvAvJzGY8RASVjq8xwrGMOdGoStMufaecglZbyL77KgxVVV0dKzFuNe6z2qVhb
gRnSVYrqVIpjVpT5yxIIJuGjWakR7LyLXt5OWldwcNRYKYmD9/XCAnBlRzQomPz7kW3aSx1jg0tf
fPdyOeOFGuUQ2QvCWIC+83AR5pOVWeYJ0P9RpgSiEx5g+YWhpe3C6APfQtEJTiEfDE8ITp7lREuI
KV4opDIA7g1JIvzAshPoD82gjRdyBpLdVI6YlpNMsAxozMT3DnYIhm3k7DxH/Huad/Nwo4R+emha
TwzT5TrmSFC++zVhmcz/GUKcDH1/+QdcdwRtJIUyXuUUT/JDiCFUcdWqsfW8n5QO5ey9XDGrqWZU
uDAv2GxiGjFhkY2qiJ+tLhomD4l27EqP3aTsRhD6WCQEZdYVyQD9HL2GFBE5VqZwPg/8A6aHv+jl
qYqHXfmTuPTGpyxtXR2lXuPSAajcwtF/3CrXY1LazoBZ8/jbe4fDutFDJpUnkJnrteIWj+RcJDwY
sVy4fnL/RV8/BIljnWNcw6honTqsrUVZO0cwj6JxJjaVFJD5AKoM+AUc+ZfMb0hc4l8VfAtsma9J
a0iysacM4Bm6Vb5y2CKUZv+eDM5u3TSrt2c8cYnfda/RvWIWAkezqEq5X+tzhGj0fJrLXRTyHXTU
PfwealxYBLUaTx8yrjD1SgHYaLjWYHxXXBvce7ZyS/NRjOue/fDMnoHVoFn/u+hBjOJbh05Gs9as
mBHt32vmM82R7evw2qIhpIdC7064ZpOFYLrvx8vd1A7XINGRWCQavinHHck1ULIw+RWXw7rFeYG3
y45/eTFu4GlP+hzi+IiCpJrB7CiwtXcaU9Osd/XMJyRuKIZwpQSxGQDNlDD4mvpWkzjoe1mwN/jA
pDmPv7nc7xbW36pMZbd2yRbbE5qu3+0FnVuX9iwSh3zmShm8PtFU1nkAIdxXf0SC9xgbh1bd30jE
FcxDLKc0wGH32k49S7n2xwrN3m8F83+todIEsvFXqglQf/huFOG6p8MuNh2Ia2Y2cZrDLkM416OT
ZnpqCWVQ29pprxOm/R0nDxTy4j4e4AvfgtO2Br279jIpSzXnNQvSQfnZ8N/ICPI3LrJUHJWuCU56
4DrAnHMwB9yZazYAQiQ/XCqeUZx+PjXIxaXqkVi1TQkfeHamAqhOHIcjoDqkUP/ms5EEcoOJCXE/
vhXXcHgd4UtutqdjfiJCtYREUN+XrRvVgCmW6joiRbYxuoY2Yp4WeWcGaAywSnKgCwazAnvOX+yn
V+LecH0DNhzlglY/gjOSYiYw1iXDwGAP0AVnuuuwwH7tgO5aq7vWFllMnwjt/9mbNcZMepBZ8e19
h/T9rLh+sFlJrNMVNJZgwttPxnQoZ8mqGe2wVi5IXcV2GqvplI0I4wjrB6LC95uEgxabN3oGuh/f
2LJziBILkN+YcbxyU0JFED+Q6iPm58g4xyB7nkTET+79EY7tj4zX07F504CHHkH5q2Ksop/YuEX8
IxuzK52W9ZQ0jUfsmaU5Ak1axqmvcrKG60c3cEmcUQQsO3aFx5HGU0523lfwnc9/nOuxg2hmWBIe
aJJyHW2+y0uWUV7ZbmyBIi4KPT0o2BIFVXpO9Ffl+sbziJWe4np7PxrurT3kDw2KLGWQyW1fH+It
Zrstm8OTa3hMOsBiXwo0saEnRQ3oRI0+CAyS6rVE8lW3ZFTM5ZFAsxm5MGG+g3jh9Ykls9bqDMNI
XPA4D+kYVs8dWx3J6ijtbiNY9yjIdRNOCdEvBeHa6GK4pgvxmuZeSqzDigjEZl5nQQqf8S3GBnLE
0PNZnkUUcgzl5kQeXTq84d7XinmfZtcZBca9FGiots0nlvT1nY/VTBIuuxDICtPV7oZkVHzA1/kn
uSAfQq9csUUetacmjTQGMwuY0Z1F4F1v3u+niWSDD5mG2zBEKf2fAkI7/7DkjI0goqz2yMb0Q8Po
04XkUzsxd5vz2eLXPSkkWfuJFDumlSbOKqaU1LGkFU85CDS57RrJucF5xEAXPbTtgyZh8BMk/uP1
1Z0HttC2PY7btuGx6GbDClnDyMh+hkhmGbWIpafjx9TFJdaDKAQgkNSg1Phaw+EG+y6JnQjHRjVH
VOqqQ08K1vpMmA5hpQBItDlZ38y4TwW2amJrGXIf61sGhxZXqv5cHyXDzCOEATxq3Up6zOfA4PUz
XdS3ZDLfpd1M8blrn8jMH4Qw9i1MSIf5JfzE2FFhOJVFsIC1nrl5MQSfR/ZMwHiKckS7QLPJ4gIK
XyQw52zukMUiF24mbf32lNhIpagYurW95XiCd8EJChA3d/pK+EGYk7oQpxAIsOR2TEfyDdGbipEC
L6Z7M0g9zOGgWd6+dW07rBcPcT/7Mt1DVcVNTIM0fG7up+m2jIORJ2dpX+1E5bbf0r7Z2FVqr3Qh
zZPy/jKd+zjMOJpRoPpVi9F5kjylvofSjhKcdyZUjiWaV0idRYueKfiQO1Fvxf3M0Cewqu/S3V1I
L70b31oEixvsL8gBFkFgjHbToqtowQFqj9ro5ZyGBIuKWHIupHnmlYTUkfDPY3f0Xub+Y5i77754
1JujDR0eeBk9DbIyxuMhRz1KgKl+cqzP7ZsBV6ShxKNtWEi/Rl49/9mAMZBIgBSz1VQs/gBu2HEi
Iw8C6r3PSzJkwsINFXcdcOPh8QbB6D3mBf6PuGsJS6avvo37lcuZqXyU+3LpDuHobyNz9RIXp03b
zL2lnb+r34eBNQ9XkS19Uxo22n4d7l1tc1HOsoIB8FSh9osmRQVVAsdH2QCzpG23CyUDfltYQOyk
dOW5ayXZnnEOlWFnmPtiVne9U5ij3V06JJr26X1DVbC5nAZ/h/7TQuL5Qv2tNe+B0kuQtjyaf/iC
bcf73tooZDuTn2DEASkyckGzBRE3hy+eBSdg2eeZr2unvhQC9dylO5YUIydZ5XVEQkwvD9TlveB5
KKlmEQ/4cvJ5olVIv4EdmCoLPSxcHWgsI9BHxhAgt0oCv1lc3su9tOBm+er6D+pkCx3vMpcAum4f
Yh+CsBAUCCYOUTJNSEvu4UU/REPjQ5GL/kQDKt1fyCNbm/8O8BT/qOYFp7S0D1u8DRNZIQMwvfN9
KPEXMd8foVp+hTefc2R6VEJdjbtxQJgNn4Xs7ek+oPoysH0ij+K7PHNM73a1IssvekiPrDC/rWEE
nDh0vUYa8cJMatD6xGJjlvSsCnhyuHeSh0n1Tg79ShTRtCBYHgMyeDeTLY2Zyi5SRkx5UIn/aPua
dtPR4J6n6v7OfmVHK3EkLt5CVT+2aZwUyyf/F50n7DxEgB4GEwf1SPjdFqfG90UX5bzBfaLXqAGS
t4LXxF6Tqk/0aDppKx9Vsfzx/Mr0fnNFRipsyS94/rHIHylqqj74bfxsN7Hm4Gx90U1mG82poK48
k0FfHML/QhCnRC3K6lZXBeKrou8Su8CIQoiJfFuqpG9LEGG0ZH3e2TNfHoAKNfY3rLI+Vt1qeUwz
7ZdqwBKXhiWjbRl/qKpeVLLstOZnTrnsuptLPV4f57TZaUP0/LCwidSeNkipLKgdkzekuzGfb7Tm
1KwOlZ5vmVsfSdTFjT5PGKslQClsjAEmF5yqWGgtskRDTk5f+gTMy36SoCypY7bNE8Pk5byXsEUl
hobGABFzvstM0/wl7otVBCofT9Hne7i6SFqvQxrPA0fAcVD1aahli4sf1+qOnz3MlCKY8ixixNB+
UynQwvCNYHkk/gU8EAyyoxRWH0usLKq3bgG2ZD85QRaPN1QTcM2scc7D7zvZtLCOPoJGodKrorRV
rAsOiAqp84IwJtXeTjZefEYw+Jey1+bLDRABwTwlavG0RY43Ojg++CNsrt0nOvKQ+OCFDMGGhrWP
HaNNvXskm1aUGwf0OuU87wztDRG1ZdJcrLPxtTZHwqEg8gwJQzbkcWGJsuwc6ebyOA38NKVUPNYf
2wmU+BlUDg0uWC9BOSU8E4LO5LbQ/LsyIMIw9UWVTB0KsqCC+Ya8PfMoKYpyRo6D5Wx5GZiJMbMq
4sb0tpBib9Zne94hya0ajy80JSNg22dSxBm1NLITpw6AYojNqRmBj3PAqCYmCs2NkGRtYl9GptU3
NyRjTVEKn1CUfXdudDHz8m1E13nuCYdt7qodGVFA0JD/csR2TTsGVcmip87uOD/PeBr4SbPVqWKd
wTJ4TppXs+G8F7IjKrwU/i0xBX3ZQL/Onyr5gAe6DmcpxRuEdD7lnnlvNXx0ZY/b9pL4RKvWJIsw
kaXXYoStJR+IdqI8D9MGPnK2Rekv2JxGtRh5aONYqu3tcoDpCbFID6hgFKq0fo1FvcWe1Ju3Pb1E
2Db/AuCwTxY7Jqw2nGUOFssXonVlBeHgkC4xTF1ezG3lCGv15HUK/4IIVfb1E4I2H6izrXFUGGOK
60AtSR0ABc6wdG/QH/IjCWnakjGvezhZ2RZ6PY0jkrlmQWRx+98OvH8Wxlx1KPh5Kv9aq/Uzh2kA
Ljl0+wVO0+9QL24nZLWmcBt97wdhAvzpMmbxLg6KcgXE9zrDELH7Hyj6Uxr4mX92Fm6SO8aN4+2Q
Iagk7yMqn/u/Go4I+213q8Ihj3GVqAp9Za9nrAYrzmuX/EWvbMQPv7ktcq5zr1TeCGqfCh3Ef3n6
kjXOz9DESZk7oM2zbh0PAdbb5mpUlNlTymmgGDBuokAD206oUTP9nQj5ZLgBf960sTYV3BX2HzRo
FagtHrNBjPug97e/L5lhhciK2WTA/oxS6ZTuY0gZUH/3YJx+r50M1gSTRwt5SPhhGtKCJvy0fRk2
pjvKxP8uSPlNVtp4Tg7aI9nzDLak+4SKpwX573y7JMFs5OuyJwLoVSv1NOLGHLdaP/JDvTRBp2fI
1mxgDmvzGMu1UH1dRB+1sstHQUiBiygejzDP0AHyqwCbWhfuRDc8zDr8wHboYVQYWoZpQsCqqGWR
fc6/jcfPnvEWliC957iguZhtuAN6+TXlYT4ru4azKzrBMQoYN2SjIjVWUk58HESuRYS5F/rumS+M
dbhk8lNwZea/V10jArvFfwLNzy/OjmygeyWK0IwbuaE3yGaubU1Ns6nhjmbH/kc+zcFVJ0P9AlNA
seNqN0N8HLFWztzCHw830kQM5wK4lZQOZCde/Z0K1E0Oy7ofLsonTn8DpCXtUFW5lSv6yCFw4QoU
4fVhAN8yGQKi047zh60HjojWQNW1K7oitQ9SW6XW5M1ATQMtTQuBro/TXndtqr5EMe2iRRpVQNPu
O/HHctqt611PouF+a0c2zSjsRLxsfpvX45BB/j21OHU53NTnCGaZvWyiTzSP9fTdMLNyluxe9bPA
4El3cslH0U7skkzoqQkO2TkA682JAzz29BIvz2vPjaTZBI9sqFNPpQlCo3hlGeaa3Ibomo7PUheA
ya07RLTbZRrhtrTZ83N8TiCNW+QpfTDK8DqOCaLpGWGZ9P8pj1ns0viGezgTeAON1PR5UkLznjs9
lxPEnikIwzp+5uMGm0wcB65j/+l7EXNzYwhNdVwPVbminho8X0qhIQNEsPF+fUB3cehdAZYxiq3X
ggmAzGhT6uxeL/+MEa9Hl/V8VNOyz3/ohqVUHKBRYcBSO6vQsIszP86pefBjD2AV8VH9xQeYU2jt
TocZjOktqUePiApiCNnw7dSNh/7lmnvhYxsKhvowhclmelIfq4YColJU0qh0pZEZbz7x23cK8tXU
ulla9Rd+LPdJCnGAxrZL4ku0YefYfgYzWXk3iBS9OKjdUKvmCa3RPFFbtkQ46RaDB8xPJG+rU4VC
TeeX551DJ7Ltqp7AgLfGQd1QYYZxetPZssUMvNAF2BInoou0LF8Pam3erCetfFsyeJsmE+2Qx7AV
hw+ReHCFWfOw3VfHzUa/Ou4WJC3/aVsYlWCbi8jJbUz4P920Bf9zSVnhnJogQpDVSlB0Z6qhjBA2
jX9N5yLF8bpStefZbZP8Xt06zuJx4BRqomXe6ijsC/HU6vCOOgCZjeNOQR0tu9R8n/Y1+Vixe8Lb
oHXwS1vnY5SES+GquWkmi3vTEmRpu7v6sillkB9FI1buvTp+6Rq/c552TG/0ov5xWvIrIv+wOkSX
hvypts+d2MLbS8BZLWUiVG6fvBWdTmbsvcC1MNz2BLAuXkKlvQ4eedimm+oPSHEjB9p0avlfFByg
KO69oSqbjQhzfYyh2LTJCML67jeL1jNiBRGbAQsbZ6xdJbEXqe9OLvVAJBOTYlD2YxObBFAHJunf
VxmD4fmBnhrZta/QJ+t2x+j1eJeqimEUqYbzNGdPfRPypjykkA9MV69s/cL0Kx7jM0gLKLw+AqHI
XfDw6jIoYjq1qPr+ME9jJer46mkmKt8KbKNQA2EthmNTSxyXds6fsFNKg+4eKOV15xL/Mn8P13lR
PgfY+X45eNX5/juxtZGSThuwSw6ifLMYJ+GpxpDFLKfuedgGaDnepcHiQJjcBeRU1K5AZHyVNvOp
+Mq75NAuUa/X07zvwCoPakgX0FycM9uksoZhBLkaQF46tGKPV/+Lr4Z+yowm4bm54Amiqp9ofsdX
/Sj0PJbXwMQi3div9HWa/NKksHG4LO95uExe10CsDVSb5c7uTjpBciwTNRHlTXnUhLUADNj+w6fK
wacscJftqn4tXjhGjz2Szs8AqGDpyfoeCo1emPoizhopVLCj81HEsTmY7mRzEUySzY6zsgUwMaui
DUysIVvMrtwLsoURNfgtnwktYdVjr+JTcIkGmna66bi3kkBriK2WIs3KaBgaAPR79b993p8nttWb
AvbZtqB0b+cdYuX1fNyv4tRBX+rgnkxfZd1TaAV4H87bEdgpCPwb0rdjyOnJy1JxV14ggZlVevw0
/8yNfOww1LqkMi5G22rbQ5ZuSUEOzrZjaBLuJm3XIcGfiAmkPNHJHa7g2ra+m6VVibb3yonD+9UQ
eZVwMqk+sftka0Tni7VGKHEP9w4WYZuJpGTyIyx6f8Xn0+jv4uxWMnZONTx5e+OkyXkGZI8ynSdl
qC8j27H9VkKzQjue7JAV10BI8sdmA3dKDZBPnUVoqm84KUfiLqXOGfLK6sVHxJpp7OhqBR3J1PAT
loutnsyiXer/Xy0k9rj3uKlYDUFuY/UQ+Lt/3rp96xdwXajIU26pmSZ23tM44xvNsQBWw2CSmEro
J1gmTsPzy/mVrnYMysTmQAFvfNz6YEmpMjyQ2uAQpsmJhHPr+gPYNP/9/8rKaOhtAWZj/BInZeuI
BKE5Rac1cWFPccvfHVPQtmmfWcojj34xfQhzvJ3KUePNDodqP5rKxZeGXKQVz9vaTOdUbG1jMGPd
1F2gv3VXjJpULGAJFjVmkicR9sH7UliaF16xHqb3/qt+eW5PH38W0T1h0c+fIVtYVEBgahwVl/LR
/bKTs+wUR4vzOacANSnE4o6op/JmUjB5lcQbrhjJvzk8k+U9VHWpbf0lROAXP85kjs1/9u6Wyezo
alvI9IpfoZVDPc9kqM3VlSc4zXYBAWZ/mqX7DH16EygvOBvzN5wIuF8GHmG0WKKjq3Hww/Zxd6RJ
4/I7JHEDRmOXinQuIDlW5v/4pygZwwZoCZyRk3u8W1nO/FwQPL84T4K6LvxM//kkEBtBhXppbNVz
toKmNKhn7kYwZ7qDikugMJbBhW2LmR48AgC5q/Lk3SHvwh6izDutJ1d974X9gOjqmeNNccwBshXh
XC4VkJyKhFO8FD956fR0xyPLleB2kdI6dVt6oicLh+jAsjl6T//nvfYyyHhXQ6+ISv1wIPt9Gl6d
Q8RS7cKLia5IeV4nWN6hiHGIW7BIRP38WBrIRQH/bEWbz4EeWr3f5LzCChys7B1q3JoWOmNqxJeR
meKVUBhabKvGLZlGQ8U3lkpFt4Z0oc3cWZVBj85AVM9UxfBCmZ0viu7VL/WrvCoZo+MhcweG7jnS
+tuctSQpiy2i/xu+DYSZnTU3RYYEXLrSRiALodjwR5RTCa93Rxtsf37e4wTXyaB7lyVn9WzAY2UH
H99PPMIUyoIf2fSzc6k6xj4qZIU8iGYX6BosQIhrqUWnFVSHXPSj2FbaISiZYaJlRfUibL+FZd2j
9FPQjTtu8kZOEWVsuWZHLvX5kU29RDW9odzvlq7moLkKeu0FK3uA63RGvrzAWwOvdAA9kr0HSfA6
4LarCw5Zx2giete5iepSoq50RDtAQqfY6EjJfay/rWwyVi/ey38y4woKxA5PXAZHe2U2dNdGLEOa
9wht2suXjfREhvrTsitiWI87ucGhCh7l6sVJkuWhXOPITvvb1kk9GLKj5eC5EbB3j7k+39/1dCn8
F78uj9EZAI/LO49BCrYFwFug4y1nlWgIMl0Mq1FV9J2ZeylY5u1konNsQ24b37Bg7DIwR8qm7GGz
24MfRZXgBNvC3Ev43mKyhbCl3PTJVGHLJ2F/1CYrmN9WC+1v+vPEoZjxP/k2bdHjhiuS4TKWKEPE
kWFJU309fGK4IcUTo4AwMPmAr+rvB8jVEo6KapAzqLGWCockRwJPGkwp0unPXc2LU8jN6iLYfdpn
WYw1jQ/2gSzGPGSrfALQlF11i+OYPp9/XvAv/UsKwpGizIiJiUFGeywLmX+B0APvOdp69CjAxLcd
JgefYmFpEhCjcRNfAO/7ovBAo3c9zESCrXIRIVbUgcuQiXkpAeEPw7wCzbiANg8QU+emukhCQo+N
iSPdBbm4no3DHP08bdRF/1A5A0vmVJHgUbWTPKVfGMGkMPMVOvGkS4Muzz95Z+ciiMNBGjyGH/ld
QDxTiiNyrW3JNspvtWAHEms6gVFrEYgk5/ZvU15uvRliy0EyvU4ilsk+Q6X0zvWBkmXbN0CVGXaa
P9xs42zJmFaznaaceCQ6CQsfctH7I5NXq70Y2XwxD+moso+/ookIMlMbG/zTO8PBFJ8HkWsznKDL
f1pG9MuQG7HNp3hIruLDhCdA9Nv7a/zVTtD/Lmera9zUcyFwncyQc8zc/OgMOUorTM6bgDmiS/DF
ss/atHZW5mywJ/QLcZ5bEFGPGY4fxdA+pIPWMBnHBYLngyUeAKe7R3hKMqE/xasHB7SGkYN6wVe2
w0MO6swSqGOg+uO6pG5/Va63HyPhVCNGLdUzHn4Pcl1b8dHEqeX3+nacVDsJHWXv+wt79OJeC2oB
HRrmLe7VUxyzdtZkA5eoPMxrgD9E4bfRaFDlT8UZGwsLcDQJXVwLlMcPJlnYGa2KaYBbq2sz/eCs
OktOz9JWsj+VtrJvvJVW9o7aRxv9ghCW9l4BUCnzTYqvjrpGLx6eeI2EN3zHqTvPoiGctP6+Gva+
/6G8JGoO8vpSrZV8cocf4RPeVKsJ0y/gdhZEb+3pvj9lqyQzjErqlWuhZDkIPLd25Rhmiff3hFCM
GljA6HylCAZj72N6KBqvZ/6nm10CjemwbINI4YDcWQuMUdpkwW5Dzz7V3WIYpgFu+165AXW335Dh
CBNyHoctvXSRA+rJzilNFt9h2ocA+XrXnQx3zE3ed45md8wfwI83oraEo098BDuP2774mejhXsAO
T1F1s0nSf6l/zyth9xUIz0ZZG0JWhAmmgcAXd7gMGZeF1++KI9z5317IkMBC/tsYrDHVjCglbjjz
8qZyK6BAwbt50k44mrgqWH9pUTvn/SwSymYcqI9dEpzhLJsUWT+dLc+/7cZwWw+fnJIvgh5RMDrM
PlsxTEHEeJ58MXtueLc0fRnR4U4vAMb6IlAjaM1pjww3vMm0wstexF9JxPBryFTy3qBPGt8CZQtp
mV6UVmYq3SIbiElaXaUqPyWeuFYMGwYib7ZCsNORDrB9xK2ZChRYMwbvtFgxqE0demGFcIQXN+r+
A8OD07Dk+12HR3JUgfa/3SPuY1aVR6u5UYzDcj3nDIXvVela04cxItoebTO3ytKVe/QFIpYev18+
B+tfF3WCk0Kq8yL5x5vjEb7/zuMZTR4IAMWqmhMmVRVi2QuNBb+huonw2WQkEOAytOYP92Y+n5k7
YhGe90TCd1plNKKwTQ2dqyb96XdbQKOlUCfMHqS1y+Wwjr29D9x4YtXgMfe8OCLiIwTW8cTp60QT
GcEx94CCtRjrC2lhlbD+8SuQzwBRcni1k4SAscP42KS6tD/5JxUr88IByiiMoZrHKG99W2jiLvc7
FRyxOzRSJ2ztQybsqavWzJbveNq8PwMZmOh8eLsRt9gETw6CpAOWshJIHFts3Bkg72ZML6ZJaBd0
RI4hKTPDezX2hBuY3UutdUVMPt9ZdmKYS1j9L/rFWcfrPGAfT6yTL3dugz6KQyCjEFyiRdjcElH5
Scgu55tVbkDq+cuoozRwbeTKkfyV3dKRled3UCidN5fdQZ48LTY0ywZy43PXJsDFpvaagheybqCV
g8PXMBnHMiG0AJJ8lRUVplxPfX95GZouBpqHHmr/hUBdknJm3M46+hZKJah87buvR2KVYEbVTaOn
y2mgVdXmYUoGHFqxJXR3mtbNonEGdEQCOCrc1cbrmgJst4M0lIx5t6FTFstI7r5Kq98fy4OJrnA0
ioWO5EQ4rw4xQDB49TuCFhz1DUq4ugVaY9EWiY4kOZehY+O0N5m6r0UkWIsLm0JEbCuB4ww430+R
GIQRg37AyxynbIbIXS6zSwczAyctG2rHibDH3HbBhbKip1bIAcKmJ3eJRJTu1M/a/lie3e3ulkwa
4JCF+NtVe2gy9cgpCgHwzFKYRG4Hq9g33IQEcDF/fK/o8EDOcLMqEPzhWwKe178xbyVfOod5k2YQ
BBE+sjfNcOUntxT4D7WeyEUnRiVEjT2yCPzUMjLA5YG91ZuU7kW0GSspavkyYx9RTwwJ8ZJVQ9XD
RrxyP3IOyXVV1UCvPy3T/lrMXzDzHN36Yb0fcAn/2v5oPalixBHEsF9AkxPI6fiP5CTXvtv1FQKf
RJ95bq2o7ZyphLSRnTr1Qk/W851KiioZDtBMf3Vn6chTExx6KG5cVhkLOi06Ym5eyE5LSVb434Xz
P8lpEmAP7Usf9DpwiqcLp+vL+0V4vB09qH2+w2Yx7nPvfrUo2LrSniX8+JZPSEotTQ9qwKqHtBD/
vryzObuwTXzKihGTeuOaSxSaq5dYQniKOdYNzlqdvwAexZsJHlUpr7+doYJzoAsWeTl9WoWPKL1G
Uo5tnVDD0NKI0x09Aa9EQBOaZvUlx8t9b9mGk2xRDNcBXG29bXKbmqBJ1wtYCIey6e5iybH2rsI5
XvqLoJ1N5YP3+PZBfttt/G90qb8HSot0vwOC4zXyVYrAugQSGnWhs+GMbyQq8VX9MMkwYXsPGsdR
hOXG6IOwG6spdsKJ8NfT15WGMrWKhOpM7rYeOa6tbxEsfXSdgcCW7stCQfN9FCb0AObfn/Hla7ou
Q+uSPLqnLuDZCxWDJzBnRmIjbqeD2g1FNEpdmxDdHnlEsSSpuQuKq91wZupPNThU/Cz6SRiP2lUX
EgZRoal1Mgl7/3qWTlpd1j/sSc6++yuBWqJuC0ooeZJ1Mh9f7xJ0wuZ3dvxYZ1cSUxWKum04tXB1
CDNyBblFJG/vP4ieOuS7HQ/NuYos0yOC2Sh4HfC9xWMRqkWALUlT2U237t5KE4ePe4fHq1ckYJVo
MYPq1G1XFomGvqBIVfS8vULxW467/WOw9hoerZmYSAQ8H5LiTRDfO58qHGBs/GHuCQmhtTjAvd3b
9sruEFfnAlfyEjPXzg8fQT4ZVIgkOZa4vrH9x7E5LmymtlpgSTHGUwKgxB+5s9Qhe/pQ7DJbL85J
2k6f/60+PoV8e/0kSS+s5f6GLsDEqDWX5gkEVoDpS+Ya36+aMzPpjj27qqaTcyuxNvewax2OmhXK
1L+XLweRwT28gM9qvLjYVM4UXkEHH36XW0RCFbElW6puWXxayWhYTQQkfqkMFNyyOBaFvq72GP+r
gxcw79+9EcM3t04jYA79MAQOUfcL3pdyUk1iVSk8d2hETHAjiC+gzdDB569v4cRodLfsonrDo3lp
eAjH8XbjKSFMqvxYjanuEzYpozn182Nk4k7Q2tHg+PXqCkj9CpWiSwrHEVpuUUrN1ka4Lfj7XifJ
u4vgpu7HbzRF7XE3jCIaoaMrvygT0WuS7Z+j2XKNcHxgplaebOkm/A4HZv+3gjTXBsegC0Rc7Au+
if+yra8ISJlZBuBVpvQ4hpYSKVKEVEMtDtm3mH3TGvV4m64XhKtXgrR6tk3bDbYYPX1rZhetPhOQ
fRpEfiFESI4r2Ea+NBtTd19DLzMjqamIFtROgnwZyi+KLOygsj57HmeVK2D+D93LtTA8CsnlxP2J
nj5aBvMPRNMXRznCvKTlforazVyWncv13BvkwrcRJlsWmDtACfWhEGMfpUf6ubhHSzi/1+0rqz5e
MSM7IX4fyEb5RpdB4G/uW6xsM46HN1RtSygmIFPC70GC52y/kSH4gCZxDuW4rkPsRrSq/RFILI0f
zgLIjiXG6Y8V3cGN0M4PZgZI82yFx+MwKz6l5sXnuGXrOo9XDB4k7LqR7nOqu3XZHFxpfQEs/hOu
V0iy5w3wBaYctKhoN3NAvMS2DbISVOXPAUlr02TRiw1Jjc5ibKyE8aVa+wtEfgxFHo/D7BZ9qq0T
SvTFRGIteky4+hEj9dUnYQ4KWxajnyypFASVVdyfYSfLlniym+yuPHi0eb5/ung1e2pO6M//+6z2
yIouMrKgVtLCc7ZnyrvlGRpCoXFG2lMGq+osG3JBS2S4rrupeXNmHO6U4h9rgNnhhX1BX3V863XW
kNfD+dpwRqHCiONEuMFeoOUbdWN+PXXFC17l2h7HWs1Coq5z/FOm481oEE6Y1hkcGe/P0jA0G/Ya
5rvMuGbzRD4qQgnmcUMbJsC5wn+Jk5V4Q9v+PuUTsT98HAOMGtm+MqscVLIGtgo6V8s60Pgjz51A
j42KO4equaIq89SF9poili9HouVp7ShhvgZEsGhoS3rhPja5AtiLXSQKX89KPRgN/HuUHkB6qtx7
JSWjQ5QRSMRS9ACpP73ioir9DDTBMz7AoDnUphk+8vPOgCQKRzru8ab+ZRWUyFkby89iZtr+3ZJC
Whz8xggVInuKLIPEGz2EJMQ8aVXNJAGULl9oKJ8tpQ8uOd+XJ5EHZm8oQsmLIp6DIU12eUuYCJBo
F/dkimwyUsiVZb/In5wnOX9C/RFnDaa/nbJBbFWTIWDYCkSQ6KYFtRnwZOjK5C2zKH20XJOe2zu9
3YMJN93POcCEjtCrUP4J3HV8k38216qH+UxwKc3loP6zzwvx6EgU4eJlJMmHnJ0LvoPL86vsAAbP
wGQOUS0iVaD7bbMmFOtVELOSAgrM6XGWVJpDhZfqVA+WFRgA0t/XedVu5TEydEi611X6//WUfpWd
e4OqIO4a0jbCq88BhIisnMNOmKX3NWJmhFLdvuy75700ywRzlKauP1/NiDn63x73TqXZ2P5FxQVO
Fq4YOFytqPOMitJ1kQ9hhY01AF5qijhK1J+e9SjGAc7o8GizCkmK6jacp8ttKmrTxqUzD5S5dkI7
h4BvJsVjdOX0Pv/p956qGee9ZhKZliDLNHb0BNdf3podIppyb2QZ20ecqK+ZtfTz3DaxslasgnVo
qAwqL7sGM+fCNYPLDJX3394Orq7E0knR2BDYg18xxTavEuQ21+4a7a78pFz9/ScwCc9uzTi52IT4
xAcYPpM2G9iBFgVXc37w47pCoIeox2yR8ffNnAea5BZ73ZfklIyPrk67+18TGREqdeLAn+P2NI0X
LTea0i5TUhKgeDpBFHSOQ//z55kjZCp4yq2Vk6eS0YDrTaOE3jRRVkK7m/+GUtLnu2GDxvrYizza
Z7dY6+6YqgGMyL4/g0yfM15bWJJgWTt+f7GW8mHi+ujZ3Nd30ZqzfNh/Uy8SvmFkmKbU1MR1e1Va
+dBYyxHbzgVF5nonMEIWxxMR2pv5+WZykIv3CEB7xJKxLmdZF4SZ9+qOoCeXIixT3RX2c7F9Otca
Fmkwtp0A8CLTrG9O1Q3xVpZ0/dw/yJnymS6zRhG4rTwVt/CheKqA5ZT8fd9EuTZuwi0v8zgD6B1s
ryFMftA10kzLu+OkMLSSDZNKrwFoNNLNBw7LbPs93zfSeNFaKfwC6bI63hs5yecMGa9qJGdfRQuP
VONo2QpiczyZDMuoT3JyiEhswDNRJMW6XMx01ao2d/EpZo5IHx4yClcqvy3q+qx5SHJ/aMHR1Hv5
gL4IjMCiYqrybzKQHrtj79S70K6bOZAabTtWKcJkKFMiC+Lfkbqkij2pFqIVSDy5wZcCpyowQMK+
jEiFzCFuQuPogaHw3QPuqJ9agvChoPT8MIZdZWFPOQq8OREJGW2sn9UN2zq9fvPFaLjEHqk9F40K
SpG5KwJBJsWr7BJSBTdqufDDBgnXhENAdNcZC0IpdGBCajCb1FbCrwfBeREylZU6ItzlyzfWYUFG
OdOc8mTWXmUDeOGuFcyqq4qaNUuTxjUIvN0vStNPddeu0w/GVUe0dpgsgBgAKsVIbimJWrVxDQ00
gwudP3YzqnhFALQpWbdaxA3P4K2DBZWC5e6YPSyvzd8QI/2le5EqyEzreC3smDPN9zZIsA96NVHN
TKKVvmd3q/toAI+7/kqUb+jiqamj8409j+fK73XVJFjjc88EYdycvh3hrs0ff4DdArfm6r5fODSZ
4+Aitx0MkOyalB/h3AhHumrDC84aLJWJeV5euNoKuYB+oZbQBgqr0iQqygKe9Hwis3mxLN4C7sxL
ot5P0zH45N8xhGQoaBua6IH/ex1923oe9cjkcbOG+RIMogrMy8gMWDWlmP2PkLifk2aFTTBba4FJ
1SKxw46+UhRkUyAP75lpk95suKkj/cBYxbVcwL6PKM1bVQ1HONEpK5k+10qPiv03OaGeUlfyurnn
kKecBCpu17zLwyqpesO3gsV4cfpXkB4b5E8HwIWHImBQwnEr5f3kKPBXffDQ9kjJeu5OCyETIVXm
d8l0IOLPeMY2baAGLPHxRPxAMdYyb2LBWQOqhEjmWTS57k7QD80dq2yS1Cj60VpZKeNtCxvKfrvx
FKKjAUSEgHrSNla+4qYQdbD2ueCpk1xd36DDZHfSf0WsqPFgDN/u85lii1nRPCLMTG9YpoDRisik
xVFfJmSrna7mx54gKG7HjrGgLYwKeJynZUPjMmWwvx/uhN5fEXdET+N6lE70ypb8HC06ae8DSOwz
DA4ADTbHUao1AS+tRH02pvaws3HT63wdfk6QzSMjjz7Gzkav4MXLS6vkk1Dwu77uUDK90nYmyH7f
QaR8JtVGqNFdRSM8/QLLmMgp86zYxTdvhMujUXsEq/1EGC3hP+FV9XIZcsEgCM5oAhwS3NLOyZEx
AjvBDK2ZE1TpVeMbV+iOBkT7hwfOUbHn2fln3Vr3qBBHWfPWZKmpG1FrgysgA3DlcM+egVVpb+E3
u5Q6PkmDp2ZRSTrvkF4qkKVjGLxNjp1pj7mT4qyE0sT11FFg20EqRh3rg0E1JkdsxagoiyCddOU9
wRZKqytYZ30qR6iFX9eGyDfQgzQi6Nf9A/NdF32a6pXEMNRG1AJNBfGarx8u3WG0Ik6ACsAuJxUJ
qn86dC9TLx5L0xrpz/EQpeSs6PiMhXqJjIDzgCZYnyurmefiztigoZKN6Eesb//7QJQEKtLJFj96
1D/ubmXKCGxYeSUClvLLkQ1BOXAMGPz+MYNtG3Vs5wRvZ1BlUk0Ntqd5e2GQHyQbDn3hyUKciSEz
DIRn4+sjTh/N4OXi+WI9H8EAF8T5p/7SOy1amfOYcAo1hD9QoYxbToqePTHSOtVSJg7lOjcQsAPp
aGaJiQqxRUrv1CcuaYbhYmlXXPOo2HtAaLkSTIKbYJbqb9wYkMJ9//pgn6D4Ny9DnholL7lD+XpY
Xp6nGhwZ16evx3aSNnoU4RJXu5BaUUD1mofR/WLCyRVRsvfiax5J//8vyatL0fKPh2dOQNuTxY2T
b7l+xx83sqKnC2IyVQ2vbdKPPFZqpCAm2mC5Em4x5tUXOyYOo+vj5uyZa0YjsxT6Yg4JeD0iKmHX
unHs4MC9+AsWgayWXwCqsjXZlxtRCquBuqhpKYA8LZqqsAEQL+kf8ZSLkzINbxbhKuIIqox/Mkbh
jOZqAMofcJO9dHsTyWij05lrmErOj+iHOGAcVVrKiZgXt3QX9I919wUWjZGj4kD8oLnirYhjk178
OLOMN4HU1+4e57V1GsSqwaAHQXjU3yMjL5a5Xlcy4uDZCNDs4aEEQMJuWS0RBXtD+EU2RmGHiO7S
X4fN+MLmaYIQuVXIoxwQ/4iHNqDM7TvDICDOVb9FlMLCMmAeTtxDm0SY8+hFdBaPH2aQpntre3Te
Lo0xgmDW5a0kTvZ7yi6I3bdRj/ogJgzqnZ4egYWUWzwbqTYw6s0AyjQ/ifbMP5zwk3lxNdVHxiL2
7AD4goKj6CM57EmdUX6oOTIh0VCEzuA5IMH05cRdtnG8thPoc4C7U9RCDj9ewRgCZ/ePZLEHVOJI
+4bIsaEUWjJY0gOkNK89bqsQ1vN5dxDU0EzoRSU3HR4dwuzuzpgkpDun6wbLsBQTf0Dj5jc5VAOt
borE4ZAezZf8/ewFcGtU47AVvisGL1VwJDhoModU9NONthpvh4c1aNnIBEC+cU0EHk3VX7MMVICu
uOOao1kqqD+j+A0EeDy+QvC5rtcWyMYadkWooLb+tVGUMN9eH0AEjhyBquqYRKzhMA59T1e20h2A
Y5XVT/ISmySh+nWCRQOSF/kAPJFKhusuD8psec5HKMGjoqEjjErpKpdBvFBMMyEsq/5g58PfsQrn
jwXU1bTr/UdEAPFbmrt/XQ6ppaz792sEYOjyy9LlvNmaW/jecEwJIqdB7RNqNXJplnFwq433ZoBh
bCC+g0Apl6NoTfCesLyuWfSMnghwfwE6q9PI3ZZAaAOnmm2x+ZCApq7UKggeLmQ8+v8Q9h8h/5/A
tflhlDneddXDrm0TeOmdy24+QzNRrmq7D86wxzD1h9H4O/zUy+/eT1Rpbxgo0/V+1pxU5spwuS2Y
FzDkwXlnqXsgePPvY/ylryJbYqUcpp9gdMTjkn78FCKlUN+aW9P5Wh9G0Bzz0QhDOlqmp4TSP77x
QODzPIMFEXjvGffU9W9eE2RbOynmfd401DOIY1KppjbcBC/D7uLvHGITvw+K38fRnHWR1RFdlisP
khYfQMp0Q7+xF3wHH+w/JvlN6IR7Tkvj6bGcTIdhmx1H7/1nU4KVts/gHyp4D4UBWk/ecjAFgYK2
rJC1aQnaKItJSZf+XpgOLHSuHe9w7wUMRmAP8qOGCUp29Sd+03i/Lf4q5W0/ARZSkGCNdYKy8Pb+
a28Cy1r8vcK2xsEJRz2paQ2m4DyWzsiZcPK3KSUrF6m5uF3OonNm5enAVTHVZd49ZstWF/zIKnGA
3yN1ONEaUcE3YP67nPlk2opE7kwUTq5S+7aSPQbvKpIQGljDhvhXF5+5DWgWBhmNGGQ9JpoVzC8/
gzGA9sqibBD0q5W6S1CKpvweBC4kW5kB5VsRsVw13lPhS4n2vChrcIlycFuaaclnUJaCbLKCmEDb
lvpTTiXtwIKOf7JWNP8KPd2Lvbxy4dZh9fbj9ClQ9zHcGzzdTsPTL2LyTyN0Ts2eUKwO/Rw0tVFT
QV1M02ZaKxrKtfEjvlAcO9GBTA/LSYVr3FFU3+BBtltvyK434BFHFMSVFYZZH5n63C7rOxrzhlUv
++8vtUzJ0Q82lIg6sTgzaI7/FYtWW3KWcL5E3YTrtB5HkkRk9Ip3EmWqRR/ka2omZAyKHxh0iFjV
WYL29eav2fVwkkErPPjqFa4Tg5bh6Rs/IkBUEz6cIvvavw0ByTPjEm20Das/goYRmrnX8lhMjBvT
WSjqtCBdfhSgTdviVLJUv/pTvIDbxFYtajSWYsf6Hyo28oF8ad/xWDX3iewtlFr7cY2JJng/Mqg+
sbXSEyrQMAGwOJhdFV3g9wzMMy6lQCF+dK6w7ZSOQlBgHzygWjYfvFBieF4+iUC9ExPpLAQzqHP+
MlMxg8KlH0P66/caM7fQ3O5PwhtMOMPjlPmDuyeMvx/dJazZ6LSPU9ZwVtqcXpQDqfUSTr+Y2g1s
3CGXNnhQAeD4w3mWEQVx2n2ELCCMJYkb7cxWBFAqCp+MZVv15tZhiN5qW5Z3QygY6Tnxx4DS+NtW
lJhiGpiwxQ09yG9Yl+2iJCSa4+g9V9wHhKWUP3dnLAktFAeatxZlCheZuTTdDcLnN77+oranIy7+
xurrmpO1FlyndWy2lxFODIcZ+nhu/qLYiz06tbYd53ePeSY9wTU11++SkeOdL64qDf75+8cF3JVl
evhhF8CmlkJRoyOcMM6hi4okyhbcvH1I4+xfd39ogxDfsfaoZyifuxNi581kZGrRbcgZ+Twx1dOG
YNP/rXLTsA3exfnteDR9AcD+M4f8llEcXg1etU9Jqu0qTnc02ubp7hlNBsLofi6L2YlaZoiCoYFb
tmerq4kK2LHHZ9AtgbLy7yd6hAMYpfdhp+/ysjkQWv0t5JQlwp60UOP6Nn4AGQ3d0IOA+3DmEwPJ
S/wsHocKy9VSt8mAchx90wUXPiS+2ibZewa9bDFUnfVRucJyuF8vHfpV031mwgtJtQQS+0tROQC/
jRwjgm5s8ITzKck3KaaVVkVopXcEmGQU9E5kjV9Eo1gNqWCxj8yO9jYMVoKsCRAFurjZobwvThgQ
HKJVzYJgh6/R8niABf2cysNpADeXEiG4+FIN4ckVjEM5IbD/QptLhYkMPvWkcZ0hAMZrAcL5wCRD
5gyV1hY55ss9CX0jRcQAqxUI8QMhcQI26wy32375pqOCSHGDJuPPeA0ubriBnfUH0TxyoYNESNVQ
tN/wkePqxfSUfFdLmfW4xRWd/BDrmeFHmR1ndJ5nLXWR8qMcs13cAe1T8jRwR3/ZWi0syRRS//hY
rh4W/nrZGiCrY+FY9sRlpQL3nvV/MRGEkMBqv4aTnpRwZMiKTtJTSKRIzeH3ANrfW4kxj6WWcc8t
jJjYBlWFEqVQubujTTDIB0k1kxV4MK6OXtTlYDZqwtsKnrCrBdzs2Rn1RbWe034POjahg0zcH5rt
d/ZqwDnFCb8V09GOvhko3GGb7qrJ0JvlqjMxZua07XivSgvhk21u15jfiCFUvBeQ49v/sR2P9c1w
htxknQIypbInkNonXDfV6u/QD0BwEcsi/cfPq/MYfpDL9PnWCwQNtPc0QcWTDDjPwyNNporFlirI
Clhyct8YYKskXn0zQsQsv759uCifX3QXTbZBQuKaug4zjcrnzwHKNVkqs7LEmvN+zbRjn3B+k37a
3NlMvwDsaz3r+g91M91xQgSWCD/ACET6vThB7cvT3HKZD8dx7YVO5pjkM8zZRagp6QniwmZxSkjA
l3jDQXRbuFZY8/0vU5iDHR3EsoXxHHKVozElK1i7Mfdn03511cCoTZdeAzYbWIo2/t1VAOg2vTWH
+VjqPwlYa2NUCL1bQMamRI96H2JO03RqpItTTNfs46tQHYMJoe4iYQwIbx7Xl3CKlGtXW8n4og5B
NSVQVjiJjvST5kP39DFQ+LxEOBKjw51j9BWz2dsNhaKmqm5F12SenauN4dPbor5npZ0T20ty1Q4e
/P32TVeOsYLpal6mvlXhZiQHfV/KroGutnm3gO7Jqa69KhzhCWQ252jEJo87QNh+akOwfUmqGWzA
Aq6+A2r+elHuzsVzgJ/YSLSnri2pEhQfbYYMjUUOmW8T+5plUzta4EEhoQIDaS0gdPnGjnr2TGqM
doPBw5sCoW62HW6bgHNTKGFcVe5anyldmjGrJmybv0izmwdDhsRLDSytuW/1SQI5lO8szXGrlxux
+FqEi8oRNBLoYYyZ4gVDaM5SLItyou99H+cOnZJ0loA58KK2JLotkcrSPH17ub9DA4OQriZfg9ut
/grjaHB23HQ53Qi/zsnpHeI8o17Fq1uUlT0htlBdAkG0i8Ne8btRIYzL7SOXFzdMyMzAKPfCybHV
R/t25ZYAnkq7sQ1+Og5MAK4+f7+1PRocCZomzRV+cyd/ENVj2piP2ml5nnW1Hhzly+1C6qS7KGAT
AA7er5gVEV/1dvqVur2y4RonRN9nU9nlqiRqoemeYvEbhPPXXM+g9Fq1vXxWXP5s4RQxjm0oVdrn
iBmgTsSonTRk9xYSQ9P3xMIt5lwf9IphwPRORkcqvtwtM4j78zXC3rQ30tP/HZL/+tFeJGu6lhHB
RYvF0hrwUbD+K5RJppS2sP12wf/j8PxcyQHsX4Uxu95nhi52y666EszZ5bSv8npX+EBhEWCeQcNd
wdvhmArTFudFMeLrAFWp1ueFsdRoJp6RYWj5J/JHJiVoiJNRVmOYSUNTNM8zmmfT8aaLrlwEa7l4
LRnyr9wUdK5f1jvMkt6MKPXuSpmruBwTGTczSGRiZqwenXlcEBLxje1Igj3BTDhq4t+Z7OeXY/Zx
vE9MwkMGT4R0So6e0nxH0PtLhNuuS5/mNwyZwaMo1j8Y3Jxltn5f2mYu0v3ABMXIEXesuIzxWooN
DDau7uRSX3PX14YNXcA2KXP96di0n2pUwkVarH8WTiUXlHJ2k76K3KX9rE5degdAGZdBH4e9XUkZ
MKqy39SDvuuh2tvcPkM8Vb1uMc+AflD6pt/DL4MsTURz/SL/0Pp43RmQBJvVfefFPvx26HIiS6jI
cy9hdD20joy6TNRG7ub6OOfeRWt/gIRk34SqNWe2Ob/xu3B+jYa1xIQwJZyUEuFdYNBaTQM3/RIH
/7380C1R8ZviTvMkX3oeeZ/2Mw/BLDdWDg7W4sxncEfTXIUIJDKpfLXIKK7Nx5m3PapM9uxgZ9I4
VZs3V+OQ9wy3/p8YjYFQvEZ33JBECKmqnx4j3VG5mv7QjkicQ9mcJkIx2mr/28z68yl6CzWbKGat
e5zvjMOClINFLHJuxoo2OgdVX563dMPH5AJbmjpUsxgZg5AHSmQC3aWtqGnDMmvyaKL1Ee5MYVeV
4RJZsy4VmgN6spT6jEapJcqd0YxM251IoMnL12y8x9ahqpCpoFx0xARTSIqyWlq6gPjxluUV4PW8
yuRgvqP63h3WLfCjWysGed6CP1sBl2qJlmrZgE+5WVWbhC/dRX6Wwohni3WOAB3ATCtEnkJ5qZ1+
G0nDaWvJOCrqR/ZHsIJvPeORK+FQBnqDHDOp1b+vtrpVCWQZ+Mim7+ONBNFREovBjA85Rjsd1S5r
36RRrxY5L119GVLx/J1rQwfwUPHUNFicTkgj1p1icmdpkL6vbJbMyw7bPEadlrZifv4k3tyRt5oQ
UgLGy1zGa9O2W6uURwILi4H3DC+ssKhaomyjqBfiP6JIW9H1nHch+uH2uwzFNUbgYJJxfN3cl1M8
sa+2XTCeaCdRMHAWgp2/itoRV+9H6ugJeHAdJj6s1qlKCetVQweVyp6aOPjuQ72PLPZqAnMd6D0V
rcQYO82SY9hg0x27tIVAlSUOespv2QeajI9+0lNGNZWXErfZNZGGXHPiAq7+VSFK5/KkCG8agm6B
bGH3q6Z8JH/x9+6NsSXhe3Br6p6D3AGev5QOAm7czvX0yoXsP/+hMpMf5UmJ/IZ0MeWx6FGNJc98
FuHieKPJXUZ+aup4fxzrVPNmhe9NPCzFKdei/Jtc5BEsvx6EuIEYGCID0yk4IrAffXpKYx1X3nxF
AnRV7wP1cv5C7By2lYu5C9cDlJBw/AW7yY/5xAROQ5py03dpV9PPPWrBpwHds5dih3AnnJqCvWLO
UO5V+tR9SyejUfFR09azEnEux+mgZosWdi8rlOd+NUr6D4yghDkizSWtzE6+1fEye1YryIECE0vC
q3fUAs8EaIgig1KntX6o17w0OMiGe4x3+PXkiXaJO2J6cy1o/HEkKhu4krPIIEoDxzSVqS27H23R
FX1m9v1eM9+sQMDFf0vWb4MLq9z7pW6H4xvT7lPML2V7ZIp9oTH1uKOY0F9xUBE04/GMAr8hGvfu
cSckadCXJXVL5KbmmupsaMwYYCKVaeDSNVsAfKdr3VEpAoNdWczoUPHLuVO/47ggkpOLoyGtYYQz
EoixvXqDvvJMpYm61ny96r5tlEsbgFbZZ7oFqNxC8k86XuS/0U7G9Y9s0G8tceDaK9EavKcLjWh2
fkkkweeW7yr+FIIABUJaGFbCDD/fUmaGXMnh1QrgNgR4biNiDMLVmJZBf1pte7q6WFsJvO4q4JkL
csgzUMvbK3sTN9URlLGvB/GikYwsKdICBL14kqbPhDIX3hTBsbaaHciPtCLVoumbnZamvkwgpNre
q5ImlXL60Ze4BnLZRj/S1JXp8Y6OF4OwHCsUEwJeEs2l/+PvDpEqlyTuEGe1foo0lme0YSxOno0V
uxRKRa5qTBBHUk4g81nxKoaPK8cLoYi3s2/rzEgbRGk07u5HuKqbA54T9YmnbNq3IaRXBPF9PJsk
BRMO4Al0+Uj88INniQUTq0pM5s28IXEYJ19Zs9A9ZEeFPnZvMMLaSvElE4L71iRcTH3Bk/Y9KVwM
ErH0xCHD8/gRDbgbpqiYNknk5KUjac8p/qL7pSGTowMsogcu84eMp2D/eaG67un/p4wVewMlsitE
WrU9G/mvfPV9EIqAXmxoJKN7O38ybR1Jm8cihYd5QdI5FoYXXJbv0mYm397RCzZA7WIVOpUqw2QN
Y1mwdS7OUXulTtGxi6KvXWt/o03ybtmRgOMcgEAU93Nu3pWfvVZ6LwdgMtb1sxtxsuql8NnjoEet
0DiGf0Qv+TZXKFd59A0O14MYWIffyjjRdMy7cZoBOx4fRYwiKceFgWriN3wEZSG/bvyv5pcx/24Q
VyAP8fRtK1jIETEgJk9X8eqotl0easOQ1bnmBL9r/HWuAYq/fn5wITwXObuiEsJJ0KR8FOb2fUzl
PKmFJdgAFjTwbE7npcv/tmatI14+u3M3QpKRJUb8GY5l2qWT/zwH82A+xjZ+bApCO8Ou+4v00T4G
1h+9iuFb3VVhIg7GKJ2ZM109IZFh9WFhQX1lgb2s7seoCwAGBhNCaLUbvBI1hTGi/6EJNxafr8Bs
FO9hz1nCJFrk7Yc8rPdMnhlS1rldTC3N2TzuJOkp8MIv/m1oRy+S7Cavu41EoULBN5vJCGBdB52m
/966+O3eS3EFjvk0PGGMRmtC0He5Gh2sZf8LI2wPxz9k1m6ONtKmnrqVgQJPAtc4o8fwN+0Q2yKm
LhAfhT+drvyfFmIQmYPKrYanZCIG1B1TXlTP0Ter5ucLSP2IgUmbhzRt//V2mdw5TggqbWnyURnr
WpaMFX9bOLSo/xs7bFlFnJ8qjJoZB9iZSKUQehISYQH4jEA0rRS6DA5HSA31lufV0UiF9T7gPa67
RLR5Mi4i58lsuUAvjTaw/RKkyBuk18IwfsEpqXRi0buJwlgsLD4RhyAzkc/ZiYnZZ8/A6TlV83qI
1JLjoA12nqVprzjIQnMS1hlap2Ft0LwF+9+w77wy8tgy0CXx5T6FuNe+6ho1zIChF1RvSnsRZfne
xPQRGJqskf+NWLqPIx5Fo+iZ8PkHz3EdcVEuG5KRJ242rRBp54HnySp+3xHjdGUilHxz3x/ynw6a
P1vokVgy2r8OcJMp3NNpupI2yoECRFcFlxwFuglc9yzZrBAAYUA3CiAuRCAnWDXbreZGDUmJ4qQQ
ik+eoy/HHFffGPssBh9I9zccE5XrfAkU4SIzs3w1bywzl0PZsyfN+mD9je6mGSTv7BR1M1PGQXgU
4FFFlUjEIcS8dH+MDNRNn4E7o4BIAjEP0q3GzJFPtXhYb5pRtyFZIqaAEz9in0yPZ3CnamJ89LwK
VxzqhAu8MrzmUZlhE9efFXQH/0KZLwgByeKGBxpWNqX4jCxmEfkYdzm2lfnSo56sTXKfUWPNsSoS
W8wtDkOq//X51hdUvmnGSNS7lnKfELlwtPsaVdJqStQU6rh2DrJsSDD1ZiloecxY6vfXNB690onb
PSDsQQ//4XC1bznVDpedVmDgK6g09AHQ+LC57kK9DtLlHsG1Liq/mtiXGBLkHTP19hslxSpNBpuW
Jb62QwmQyqLjWmMDlef0HiNJMxm8962adh9vItWysV3QsksvB7ynwFBXbA2O7s/4LxWEJtc+uGqV
CSQNxr46CgskH4IRG12yFI25liITmD+9E7jaQPOBD+qyvxDCW/9Lg/svBG0zf+VIfUP3W38BIzTP
rsWtzYANkL/KbaNfww0rYt9FNGyU+M3xJIXoG+/ph1hUeqNoGoAxncHE5FcdagaEEBNd5Wk5xZN7
I+CXFugpaKRzt74vdZomfXr8NhLjWBaxaOTF1bhlJ4lBvfyFu/tIMlKLGGRdlK9pHHzlp3fo0AjY
z0o8DJuzBXOqiyvdQJihPg93oqcBDcjHu74XsEinFf/OjcJ3jeQuR57AxuJHnWudXv8UueGepYkY
L4q1gXWlFxMS+kzLvk4026dUZxxTVEgyDTlKK+OaxIX+ijVwGFiStuBQV6dR/xnUjKPdKW3IDJLQ
t6xK4VGD1WPqmLc7SsGlsAz27CfStjY0DXr/7PFbDaFQ/NPQv6aC7ecwtSoXV9v+P8jQDl2Zce/2
ZKnZLPPfdviQjM5LzKmFl8t/kdV97kl+mbEB3UKX6GhljUVaZ8WUrfoK90krjcLZyfJ6eFydrxyx
TysBWB8kX/vkRsRyg7lzijFKwBjxV3JVMs1OAJNgKg8ac65m/Nq4/DATbuF1orslwiNVbUfV1UoO
DRV9f8oEI8CUpdr6co4BhCo7GQN71z2tnG7aP3SbBBZ1IWDMjoDy/YoTHOQgIfH6ul9120ZGJWMt
HzBIM/GTNl6//ihDynQToHgHtvfg8FlV9t1X0OB6I92u+ut2GQZNMcbD7VhyG9FY4sggPEniMrhP
Z9E4O8VM+TbQMl2BdGQNwLV1WO1UZnPY0OONolHOB1ghaaAdxuDvxIjFM6oiw/4UWV0h6PhF3qkL
inUoIYpGtkhKFawC2fp/LxQeKqc9++fUWAza+mvApaei53b2sIia+A0EH2TphpInqBmRPvRQxoQG
p+OFnP+hNvtZ3w73XiFlIWVHyPzpdnxz4SNAV+eA7F3uluJhC/paVu2Mea6jrMvpN+2QrKLeJxvm
YqU7inQdFF0NUj2WORLUmraCdJIh4Y19/Pu5clXtb4OiTcSP/6s+ybj23FLmZWNEBr4ZSmhAtEQ5
Ayw2WX9gVmRUpSkRF/quRnP0cyWNKy9d2etkKeb5bW/0PE9yt2JXF08rgedvwxKGVRgsfi0j5BKq
UmC6c5D4pnqZGf7raLOudtE832a+pFxBLRVHe6SbXohydOkHASoi3sRSZThjiMnFr5EWye+px9qo
cCyFDNI3zzGpHsR06cRh6FbtA2Rx/MslMG7PTGUrnm5s7+AfNfaYu2s8mL05qKIOs4c7gkXfXxsB
jO4h9LMkp5znnZDAJQH4ZAq4GdRLeBKQjLLbkJEkGZtvLdPn5Pioyvb5Oozp8LvSlGaOjvSsXYkY
atDKoHnvq/pJdO3b1hDldU4VIHI3kNVTArt4Zf7yfH5gjoKxI79zFIye1UZpWYsith60s/OVMFfn
ndh/MY3WoviGmMXFmA4xljYwu4B8m3Qoa/CtFvQLntbo5j5hwC1NdVgqVqIzzxCrc5JOwicF5inI
2kXkmNHN5H3H/2mYyHDYK7MSeT+qMnzS7Z6Nohh3LtU+GD97195r5ckEgalTf/XujZWWbJoEXgpd
mibEboVXxm25RLvDKT37OLgHjJdifC7W1mg5Dyj/Q0ryBb4Sqb6TULTFhz1SRzqf6cjdXz8blcsW
Cs2SqdruFY7rZUfKeEQlrcKCAWbVK5I/+Fp20zvPrg4hSyhOM92gwQb0+ogdscihB2svFVVhjrVE
T7/5GTnXxNRMz8EltjT6vV/dexU5pp+EOd5G6x8oH4XEuONFnFbFWR4WfVOjby6K7nlQS1y+WwS1
B+CkWcGeC1/mbTOwA5uGPOTvCTXriCxIBMXkxqKVv/y6dmg2Z/Z2LxJ4SPQVFQQY8fBFjqgkAv7u
Zd5/L0YVMmSfck7J3SQpNI5SIBhz9P173EVZVF3dcuzn2/q2HfkTLPnJjKbxYqFYSvi2+ens8rGu
+nawqKtMQBIXt1C41XCLZNlUVk42XxtDnGcMQUkFx53sZnDJopUo8w2hYcXFPIXv2k6VUvqNxlOU
6QARoTI95KFu1I6zC3U8INzHMvFe0DqB1/DjqY0WRnmB/NQbNATjGz7yL0QNYCRhPQbV0vfJOqtg
3X6T5DiTsWscmQgTmmRd/4ir/3SQB2cIV6qnEwMkjPcX+KIfqlpm4hJtXqyODlld8iR8MYGD9DCJ
06bZlQLY9m+IY/8kiGYxHLEVGP+ndDkXHLgoFQjQF9DXEDv6bNX5+XzKB+1AQG9OPRiV7GejKxmj
UCqslmqpbMSLRkpni2erP3yDqIK/wFB/xj/g/CpfUHd2quLxrg5QTxns6o/K3e7k/Iwk2n0vz8p6
mCnP+ygFm4ulJCtU974B+C8pztZ6eFpQjW4ILR+H7vfbg1KKdigGY/NlAPt4eJdfanpERQ0tiXnZ
T2pvpIMmKny/+lSa6SMkQilRi7YFZ7Bv73ShQwAgCDszpaijBBB+L8rJkUkn1yW6jpGX78lyyBJj
uGw86izAqH6XNZgKqr69pS9BRsMbYQ3YzjaiIV/TUqDmRz1Oaw69rglSEqgtGwhD+UW7Ka58ORJb
1JtcsRRaTWEOWoqxPelgt5xg6WOOOAmKcWS3lXWS0lvpoBrO+nrL+ugNxOepBNLspPYDGCtk3z75
uDxG07HMv8V/hUvRS5hLY2VOq9tqAi530ZGKQVz8flKTphAws//eNNoW1cjbz68/lQBWyIBm9DqR
Lsr0WDGDEyByEc9v+kpdtRBYFnrymp0+92Bi7Yg28NrM9TWHH1QoUwkQbCu6WzpHhQkSyQc5XYF6
KFh3rPTOptqS8YveYHpsO3wCejHX5p19ZmE0+sLz0vFuI8E7Kz6Fm7sxIIMnOsFQHusXkBj2SoMO
VcFGWQlXRvGBYQeJSec3ghSlAr51dCYHam9zzCvOx3pR+S2ryvrxZHXoCUt69NgYu7pgKAJhVMAO
VYODTA1CZj2i8b/07Ui36smk4XAxpvsTcdVS9aySPuY1yaWkTybNN94g0TX61IrW2yjbAEmZNHkh
Z0nOMNAwwxqp7uvXFtDwUf/p2xbVqcWIZ2bfZ/FrXtk+YDBjZRAvwJgy30dVDS3i+aOCBhyy7jb+
vZ/5XUTgAvzaM/9KZBN+ed2WlS9JvhZGqpr3/WrhhObMOs8nIJSB8c3kgy0H0YSH33eXUKe4zufV
pT60MaiGTFEWJRzCwY30Hukf1L3SCVRQ1nwRhF4w5Wuaho1fH21/g5pbli4yKNceS8bcWpGWBQQx
2UjWJ7kSpK6BnGuIBIG873ks4S0uUbJSCjo21WqEYMyKpZ1++ctGK0sjh9R2ROHngRQi28jt1bWZ
Y2MpstBAot+QDu2+raBedAvbVXG3lOKAlLlWKuLTyRnjZO+ZqGb2NTVLdanyljHc/7z/4cJiaiNF
gDZlEqLF3dtl/gU0qLTRZAre/6w9ZkHF8gcEsKFGdjRLA20mSzEgIHQo35yOJb7lcsmKbcrH5UvO
H6uLl7VJcLQgnSfg0AdquOqeGXWqxWU20K08TNfSOTCXwYoN51IdePXbdJQ6vG7E8jw868wfkXOX
v4Fw0/0Bo9jjUy8wLeF+q3yHfBr/5Jc0qhUpkk1Un/AYgWwvKcGNoOaQ8gCq+6Qa0gqNrJksWqJF
uSlecC3hry1TfW2rnrTM+tunZPjV9Hx+IkyN2FYv+q1yAIG2ZGAzN5q76tLdp14POb34MKek13My
uuvlk9rL/W3dRU3474VgY9U8OiB0JP5DFtv0ueOwUl8bG1356DrnmRppzoLm7W7miiOqzZ08ZLZ3
RU0a8NgYRPRj13KiSnwlFNSvXcJD9KRpNmXqeUyfG5Bz5dmaF75zuVV9mZG/xa06X3GvQnSS08sg
p8Oph5wF73iFi4SQLhyGwbHJwnuPAznKhHwjnwOHsmmwCDuKUBK+3jAMfdl43VPWbtkCPKn3CBEI
6CyZZeNfQ9SBNncFrj++SVoXwJhceGoYCpvpOx6kBRgNJx24mF6CPW3P9BvhSqXW+RBQfltRIC1l
2EPTxfQJ/RNf8gb51eFWQ3j9Z/qDKLl9Rq9A+1Y6uMIgGC7CckpiC97sMNyvbwG2WETpZGT/U07/
ufzV7E7mqjFLVJGTLC3kesugn+ul73c20JNwF0ZdF2rv7w444BILLKdTVuH23zLBfbR9NIrJ6W7f
u5ZPmUueVYTWOprb+byQvXmqvmzoLoJJQJjLLUegUylBFH45y1H+jZRSFPG369a1vxMzwIcNnKbs
uKSPHzOFmkUDdsPOEMQwPETZfSdEA2zx+d3lY/ZD1kmm6DAwRRDy4yYktYwWY/EflqJVk/sGEsZK
eZNPji9dBG7ciKGU43hXyJYMM31AoehUnX1vG8KIQZwhNnKnXij1C5/WR+WZFyTJX7WbfPthjiew
n/ImS+tyMGHJWkc/UKYEIUHXJ48hTq6oHAWFp8NCb+ZH38vkIG1i2rOSywO/FGKdSQRgzmuSwvmu
zf7i4C/BcD2G+mR9uxcBBO3VQQNmwMh0b8Z91G8abQ1U4EKyKI6ACdcQmE4+IAoRixcUHel6zRbP
Yi/COAqEcYjFl/+LiQRkDwl8Fj+bBJNNFldurl3MtUV4AMvIToVrJiF60AwGf02vxOEfXUwYD86t
raZ0rihNRlz8NKrEv3uvdWwt+xWVFDxnBB37CJN5+DkZ1COL+wCYHFu95WgMuoARZ5uAKOTvVxT4
50veicOB9D85bLiUvhXBGu0NY2zOj4l2G1koYVBjEVnNWIRGbiifBnI7tjc+NrJpEwZrwgNh/JLh
+TyaibahcePZNwjlKAP/r+2xYDwjPsUuNHppiK5GyzSjzy8fcwau9K7b2Y790bfl5f5ZqoVxCbDz
UOgUTf4U3tE/SE/9gPppTBfqETFqz+Os5td8dgsZPQRzlN/c7XWVXC5BwWrh3g/R/Yd60kyH+4Me
WNxNcIVnkVba/os+Z47LZk+OV5MwajNM50ioqtTKh74iU9DfLXMbnbtTi21g7uoTnlA5ePTm7oT4
9eY+iWVpJGeIuHyujnAhSGVBPZzKRM+LvFEmcLSPPe6URztIgq9RwsEwUKFouyKwgGXMgLcSa7Pa
q4m4M9+kV5SddCaBVpG04CROl4kmKFktAE12XRVhh7Yr95mp/HqUa+gVzo16YBRAR8+hHpEQQxcy
8EM74XVF7GdYboy2x8aY6Vo7qtReqzUWHl8xk4RmmbJHmHPwLYQlX0/m5CiC4bKDXO9kVwXH0zuo
mg963YVZ8meIENnQFSk5mn0bVE63/2XL6svj4SOMXIyZs1LNXll4q2cUc6ReSYqk59mZ9C9zVqGw
Tz+G1LLjHfOT+lF7hBO7ZtnaptneeMO3EmfFjgCGkQDJqAOetniaFlnsUmOIaPBWkwXqnH2cJRfJ
TELgXQKN94Dsld10jiGTBht5andcjm3JE2X0gkthMjX2hbnWuXPl4yhcF6O41A8qjMadguSPKTsm
7RnuknAW2qpDzIrKNQy7tK9XTUHl9AMwU7E/X/F8i6+fmrnybk+yOf21XVSuRaSoEvCFO/pNchJy
WTnT8pfOKJeY9DFo5AvWWUfPqbVJED94+6KhXJH6/3xJ6BJDEdfpOeInxu2KpQcqqBJyV7nFnSt+
i4jm2db3siN4ztJu+Ccf1687xfZPtenGg8r3hbAkCil/kqEA1OcPViWlmMSrWh/u5qXGfcs2Nb51
MEqa0gxJXxpQ5idndygc9RJgfIeW0rL3j8vkSh5Kxe1xvGRpLXSHZn8BX56cuhwaPsyaoxjZVaxQ
bYY+Nb2DEkTqNkDw1/jIOxB0WSvL4X2O5lL4PtxZcE1ajYH1o/Oa1iTqi5PysFgN+KYKaHJZpLQM
lQgGTKtgGVBpXWhBATNEq9fa1Styk9TjLoNApO448MUeaYOv45WB0sLI+qj+T+1ZoFMg24MGN1VI
Le47Scba35UcKank9KvvvUIWJTXV0CJSD5fxUGfz9l7evSegkJjrj1wEMTcdNvnCleriWlBQvM9T
42Yx1d1opA2fN7wuncsBfcoyWmCERuJTJh1nKUP4hjpeTSwlM77PGldYy9E2SY8Xj34FIU1C16ux
JaU4Cz3wmwvmkxMImAuPtli7n55R+4Xa8RTYFXejhIaIVJ1iwUl8oiFDikYtwJigD+Ndy7/GAMAN
HgYmtkWPngRK6yLrGni8iB1JALmL65H+toI+N3PdazCc1M4iW89UGrGWdG0h5fsckiRQ3nLOLE/g
aYOLgaGcaCr19o2Cv2odJ2b4k2XDZ8zjzhpksZVoGya7X9OZjS+0dipvHbI2H0U4rUfFqb6uQyHN
S/lGRrzYiaawAqVaGZozKSuvOeP+SCWw7w2lvmpmZ/AYa1Z9iYg4sOX89EerJuMztFCehcmfNX/s
o0X7unCy5ofrft/lMsRZrN1XLSeg1nMawNZqCDhIV5HDGrz0ARf3Ip1Ui3W9NeVUmOOOqXEzO2Xt
dHCsuUD2s/WLrcxptimxH1GFNYRqoqt3nydrZ/hwGZKLUdhT4OOXBI+JbO6Yo0Jfoy8CMl7PK+l1
LNRIq9YKcHCwffPbGrWksi44rT6GjOL7bLenXihRM3qujkayV+o6tYeJmNoV4wV73l8Pqzoh2SEA
X57n8NW9aqCwvhsQhOCz+haAOaxKYvEZijHdPwMqmLqccrtgdJ3j3UaV6pLaYEcqG8pBnFNlUW60
l8KYVLjBwRLpaJeNw2VJAYLrQOvV4dNMiEEC5yB2brRK/105uECLw461uw1AHDNTVCiiFMzi3ioe
4/vZ7hZpHy765ej1zVgreJdzQR9mSySEVfWqn5/YvjC/AIrRdADVkxRsTcpDCWaGFqU1gAig++iv
qAZr/m2VI8RQoUT0CCJV+/lVDW9E7+uVTQ3n8TyY0AquG2+J87Wyt1s7OyNzmQtsG9kV4riFiHc9
r7GcgOhcOVPWTKtxz06BBiw6AdMkfhWe3+0ml5SO9eiYjYMRnpyfHKHSqyTmV/Db7q7+7zLSy5d9
GpAO14vGxKhXt1FiGi2adaOz34A9KdSVbJk3GhrL2joILc1QTh6qsX1Fx2bOOurmufdpYLxEYbC4
ZyKP1urqmaBSAPN/LuvCuX2kxmTU9R7X7vC3zPiy6w9IGyv/wwj3At2aIleMo9a8I2S+f/V1da+e
tAHrAusr7RCXMBIgXpdw4JFE/UEQgR7xNXBTr+/wTZzj5L8EHDf52boFcckhPLbl4BD9cHP6rz9F
xRYHwyIiNR8gh9HF0PCMoCxyeh8YlkDCaQu5dDwIpw0nUmIB++qwP94G3fe7cyd0RlujxbLBQTgO
OUBHOHds2z4rzg3w84GxdkAcUvjeecCsmf806bkPD3E71/GNmMsh2+Fc3SLPiAniT/4LJ/dzpss2
veMrGnXZ9hnBstlW8m3aCalpZeLQHWV7icBpO6qdngl1o9LjCgYIMi/DrTVxgOsT9a5xYsyJKeDN
F1y5IB3oGHDkAKZO1owNFbpB6R1TY0BmJ4+uAB6OzQlCOswJCMFUVG68f4AfAMdS3s9blSOC/mAB
gDRKwyLgoTtJHkEx/FVDxtL9A/gQ8bJdg21c1oSaIu8fnWBmvdlonITqD89phltTOlaMJ4pdh0Dk
4IcsJPKHMrHjdirnMVOljimajJYdbyT/ioKIlQOiv1vONvR9JyARM+sgpMAmVKX5UBorkO6bahhB
8tRj6fNpsvLqIAaIstaKQYAWIYRhliGveLe7pt6sm4uSWm2Rp8vi1vzJNB4yeRpHYTp0PcFQ1VJV
DP7O1gmgN07RqmSATab23ZZuTGskCEQ8DaXBBGKQ2WkGHztz8hRJjQFn8DQix2yKogk+2oqcfK6L
0Wjx7Gwj2+IJGu32OWvvKAVa/HVdNordeoDgZysxy/tIhG0SwKs1iMgEAHDNmgUFyIgak+nDB4Rx
FLWYA2KoLLPM055MyWJ7dtmYpVZQ37NYiG+Nm+A0jv1zIP4Qk6ke+HrWBjYgU62fC2469bl4vMtd
jAiCAXjvATf41lAGi4qv2aij57BC6pD9I8snuu1uirgHIe618RlSYLorsJ9cLpAVdRYlfETkZ/5k
q1+VHOLUK2f2cU+GkhAuXt88Lc1vvWiAvga2YznEAMeECKDWyVtQiXWtU+DH5C7wZH2KVBspN1Rv
NoRv3yL0FfU2WSfzTGu2yxavwOYB0s4HFNhJd76Qb52e8ugg9DuD+TN6oJrfL7DA2pb7bqkLuXtY
f33ZJxoWob96GBRk7r1W1oAeW9xB50dVPrQohv3VlvOG1nZYtXww4OSX0k7iN/oT6wx8XeEQD82s
4L7MuHc+j3omjPsrmJ/aLDBojA7ncmHoaSM1nav0yYWFqC5gtQQSfiYjQ21rD8sUaZ0gLAETWKAp
gC1Ze7Qs0nqFKS2L2xH5N7HWYxoqZN+zd8R3pf6G5AxPSysIDzhXo3vvqqD2PiAF0wzmQR73sEnx
7/ZiW0rD+D+j0ErpDTfLpDAf/6SQ9VaxSHyX3Q6RhDQ4hsqFXLTHePWxFMlARj0Cdj5Nv10zZzZJ
gyxaaXrqDxee8NvaI3dHbvtwqu7kl4+8TtaqeIG0OwoUJfxE9Fahi0NuBPA/7aQJ2DwVWgIJTR+c
3ASnfsSxYodx9BZmoiPx7yI6pZ6hun4zOUYnDU4t3Ux6h2pSyVsarNr00czg+gevdvOzmBrLZ+lx
QiyzzbNnr4w8L7Z+GtLVbVXlf9kEm6kvaGDmGYrJ3Q80ZnC5vm39MhqFbiGlLGSDCL6EgPzTJ2/I
J+a9RGnHKMwNDkgN2xOWXqJMfl4H6FDGApPJce9zwtF+XAqpKXiSmPBbR+ZmaUUi6JWSBLQDq1L4
fI1lbKrUXtiC208ItHuuv3jASSWpLRKlS9yD5j6RGkmZn9U29Q9AXaP+CV1csFDcNR3ZgJ+V2iH4
QDKz579g6Q9sQvqFDRW3QubAACX73/WyvR3xfNBpQ9D1x+64pSsmrLGnjkPT74ejEDtjVRsfiz8T
OAdT0mFfd7vzoEFv8G259lSzRymYHXn0QtJL5CUUBHa72OgTP4N/jmmQtDs97KoBY/VDanzpbtB9
C8cItoVH1eHmnIbANMNddqhBYlPp25wRRTx1Tzpexp6z0JTmpz/tO02e15wrtuYcMtvms76BN+D4
twXWn9wxJWfzCdzF5iZQKJ7+Pvtn8ve76bMqQkiDYRLVJBvZ1ScUFW+TlZMAj7TuBzwuM8siVtW2
zN49iAvRZTX0ItcdcZyJfY2m0M/qKd9pG/ZZCkK/RIYiMaXILd/79PrHrDMajgBOhvy+064T6jxB
fLRJ9oI9XwG6wJb9q9/o/L7mEDm9vPaap/YWmH1ohrRQ7qZq1OR0R6r4ne4P9zBdSsctket5IyYX
r1s5wlQBX9mMYJathB+QKgqcOGWvmJ7k0cyugoFWeARXAHW/fHRwd3j2hCqAEYFZxocKlSUyEa49
P8VP46u39GdhfCFNhdf47l5i+rdRXHlGtIHykN5cqN9f0V49I3dMsHzbDWmCwKrL+3ORCX3JUzOQ
rk+7arb6mV6f8pKIf31yl+L5yU/E4jhgsNbCJy0WZPlOuYuZvPxsrjHWjPxKGHLI0IbeFLZjOGE5
rTqde83vBN32wOjorY/NYLpUyVxJkmJJsusoJ2ri4ULK/N+qRa9r7b8z/YwNyS81ubIBIty6QPMS
ZO1kwMUOxWnrAjI7w9s62pzHwtGwZy+nUkcMkW1LNfSTNQ+DZ7eEA+KKIM+CC1X/R4CWxEKP4hZn
xRJ4a2VF8BrVIicduU5qP98B04WU6Kgh12R3qnZA4cWC7PnJg7TzXtswAazvUxDnqqrkp3Kn91Sc
s4mvM30O2W1ATqoNDkJS2QWMKubd9jUT7ZWIWsrPDmpH56xsEhdql6TkwWij2BfRK2G8fS53QXen
VObEd03/JRldga6ftYuJX5T4eFMoDM4vuRy1cT64bC45dp9g76Qr1Bot5S2/mKoT/o8I8+/W0IBM
GWi6pnTBSMDAMqdl2AKQEaWNCzMgR5woEFF8x7RsocCsPZBDJ8C14tPa/682Okb+ty2W6WegngdE
dHGxJwIeg1RuJDO2ltj6tU/8lrrIz8Ezm0npgOrNtSfqVbqZ1C1yu8rwrjqbMVP9srhkJEtRDrDN
JJDr4RHrnWw1cDIUk9ETYKGaFHGoWv1ntz97IITOXsuyOZF8/OFjhiM05oGMzTRMKip1Hnuk4672
nscORGQsECYhSaTu+2L/mNvpB+E3myEK84d5oLs2CgME+tk0Nlwdr0FHotsJIUHl7MpgwbBGC3UY
1QBm9hJlzM9mkwPYMilCQ3DBOQ52+zSBj9gJ53V15Pm+8NCdSiAO/noIcokTLIbkkpkf8t4ZBBpI
Yf+yEZTlV3vTLSGI2G0daeG4oD3drI8wCJPBFeDnE7/P/9uKuyL8CaUiy3Aylj+KfIZpEPXCMhn4
fu6YGeOAGBJOt1FrYMmXSybD9uD7Z7ik+cncPFQPuGeR0dKYJN3ZmfzyPtlKtQ2NAjL3SdhRrAGW
0gGX1Pr1uksao3232mw2Cgu+TTszVFnhTYdqhN4SAHqC8RcorNIo34E54pw6xMSl6zl0LS81y+RV
chQp/k6TIjAqoSfDMLJD01nmQ50WX9exdJcivjxB9L/SkVQuO9152rARFqSiPRs77M2D51fiWa0y
Q//jXJqbjzoiszhXYfFQagyplChUzzqCBbJdlUe4s+9ArwuyvfnCB1qr8oHePdCne1enVp3E0/pT
FhUEdC1ehl5p3/rodPgdcrcAsKZXGyt2Y6iZ1EW5Clul51KFFbQXzSU3Jj2oMKKuAs2oDuOJxJbv
BuB93vl1+Rrb0p76lIp8XYtiuyazKcMDPAtozXuW0qr7knLpAYXjTq9/AAaWrPgjSPmZfFJFZCgJ
aHjy1GIuntVx+AZgmyxjG0sEJ+zVRI+5XDu/OLdT8jW5DzA2APbgC07iwCLmcaw6j3VNz/4Yknbu
72sU9aGDF/UPb9PXHuGcQc0TYAIpOOFlX+R5Rnz3nTWwoB+lxWaXLIJ2waGDPdSgSpR272K6zPvv
5g/7jIo17PrzVNl660DgV0GaY2GlSw8273qc9uJAG0dCQALasJN/5DRZwcPq1nOj1zGI5fg8PglU
OrK5yj2aLGHIjsYIomlLRm+SCFqq1L2O5KQl0Oxbahy4vMlJr5dAPV2czdW1zoLKxsdcF+PHYv35
llu5jfMF0QwLG0O06pfmFpbbSRqr+ncufnJdux2LISjna1lxwuO74PCPXajseoA7TinPrPIGYQpE
xJ8rtkZkBJeqCNzZR35qBRU0rWhkJucT6HZaat2dYhvhtr116AD17g9UuB6yX20HlVL1luen8qKf
eCcxJurrAJCVo/32tWpFLwpZcwX9f2Mb5S6U2b+slJ8lYK27O4LfgsIOGco7HxUFaxQI+pKiXKOR
EsKfYulJ1TpdOJvtqQk7XvUp0sgbsq8xzXf8TudxCHLr825FXwXDAg6c1Fgd/b2idsAB1xJyAGX0
Jw8TPQ1dE2ATDBFt2LszmAY/j7L+Fj8/il4BAhosd2iyWniKiS3jniWE7yxMpS/hIVeZ1ic2TK9t
Td2P9JE+3lzfE9paULPiQdt5zm0SYgs0lUE8NXN2HEyAWilrWAVYlJ4/9V+WctcHhBEHFXaMgCBp
icSjaYS+0Io+/c4lav9NN2FTwXsKDpTs9t2+umcZuhomv6GN7bCcXSisxCt8W6Qq2Xcv8fFTSnPy
yNmLCIucr/JNMAKNfzYzuQpAeY61S5jmc85THnxuQJWJSTiTL0MaEo2iwyZaP2pzukp1TEqP8EGU
sX4gLRvZXuK+I/ciIM9TNMlVd9JIANPLEyDBrNGwvHuHjQHkiavN4qpPyFLGfLrKIc9X9/Wm7seI
1kdwYkmulnfUeTrWwpQ2yDnpL8tKufve7aYUFurgo9PnrBwiV2ZF4SJ8OPNuhewlKF7s1H4of0ad
ViVEDtxJmuL/557+Y+07AUTZ1rlmsx39eTJyXYCm3uFPuRrkUmc2i41d4uQCxZ/5nzvj6drvpFjr
f2fw3Yz0esBUY1m5kEHJvopaG97IA13r8p/+7mlAXhB8aYV6kLQOg//6SqXhEDbl1+3RtXZBd+Do
cm73HUdyk/9E01jQfD2sLRqsdEj77ZLRCEWxLLM34bBThZnktObniJwDB5oiYQjy49wNATnVO6XP
HwFEgUH15RBSbYO+MgONWkumFeTdElrzhVbYjcP2/gG0iIuwqxgeK06iLOSW2bhd7SgLOc1C6EyQ
ajl73m3acch5K54k8o4FTbmRpWYlWfL3YzFW842+iSUw5kSoSxl+i2o/y6IqME4Kw3dlu3zZWY4v
K12/7AWSJrBR75pUlL1GEpQK7w/1vduogmJAUAb/p3p8om8MvFxdi0s1O3gdB2IDIy8UNQCqVva+
p8wnL51hU5llsVnTPDL/iD0ZDQVKA6SdZwbs32pj9VSSAZpSyo7KXLHCfFL8b2BsTtsz2KLj5kkU
C8JSjS2wI6RzU+pj7iMe5s31mEgjEySirKteUI5VGzLiC2KeHZDSXXnNMWYd0DMp52FyqeRllxIG
WLGEXzsyZ5Gv4AzrRk7KoGIJU5Kr3a77pmefx+CXV1r03Gxgf5G0kMgVlzYfcGLRf9QianfOW1vh
X/DQjrkYSgYO8Q1LEoUo5HaaL+DLoYSFAZCfTzM/48xMur+1oPAREFWjE7Rvs2OdP5+JPtgPYyj1
q4S9rGQ2IBhRsBzi4vQktLFlRRpXnUSLJepbM+Pq47LTAL/g9aY/dowyuEm1RH9mEyiNaXPS8jSM
3Oy+5db1SSVESnxoYkpB0DirBY18Ymp1GIZDxoxiDNe574D9OhFprBOkB1rlkT3EMEEsHzmuMIVW
3i8Zmeq8ztbdVCR+YspIiIc010Fyg+9KrF4jqfLpruW+QIvoEOrWUczHmq9UHMpbIWDn9sBHmB4w
Lj86iHrzkjLu1u+kGBetlJ7Ce7+eqZVAcftHXve3wsj7LmRPzZsXwHhxXn7NCCjbU/LYoWKQM97a
xGj+YH3rgQtnSVbj+nQEtQh5UhztQUnIDxGy8+tBr0p3Z41y4WwYOX0ibFiA9XVtr245f2oizeuA
kvgEeSm0TFpmFOcr9/aPj9eW+MRnyfjONRbZusQIse1MKS7NKNdW2hGNYvEQ0x8fuWOocdVy/aRj
JP12gvQ6e89yOewtEUVJFM8O5L2CwBi8tOJ4n2jQockvWUzvpMd7VI1B56yREFXDdcSmOicuQMU3
33rvMcpLldC2/NMkd4rIHSQbjsHjA3JEBimVfAfytuTa0GSmRYEcOqExiHCboLB0o0YcIh68dq5C
G1PJNxyy4EUaW41GsEDbnXExzUXfmZkGRhe5mkC+lQ1jrZUEQrLE/0JO9HfU+Xde5J4tjmtcFoEP
FlGcAt84hzZxW1d0tZz33H89gSgtJeMEB6/akxZIBwujx2+3nycESX4ViVT+KJnQ2qSZ55SBk9ot
ZbtZ+PwSK9g6Bc5K0nfybjheDuYkH4HDXhRhfGktGn7ZSm1DKQzhRh24RFp7WBuvqX5iNOfy9hym
kvSVsg81/00SQGssCCG66ETU1hrtuDZtOBxTQEUX69PHwKDSVoI3SS3utXv8GsbpE07mIl0TAiTf
XTDmcgQulDhlcHIxDxv+VOIdo9nT6XyqLq5wwdfYLYVgyuoRpZqUoBXCuexrn1Yba2JDwFiICbHV
l3zTN3id+TQheSiLTyOQHphup9rd5sRIWLUMHK0wr85hN9zY8Cu5CrWg+vodo+Rs/Wc5E/WM1H2s
co18u8v42mNy2we4CXGdnGldwdyKt6hfmJiHOEfpCUl5IqYRibFVpKtYwY6paGfSuLTCcxxVuASO
ytntB2t/1XenjZ3Lwv3Uc1776aL+uyPqjxey9/qDJf/QRmp2/DckV2UJSE04VKGU3uUnYI7L8wVK
msKPFrmiRSYwbuNH8MRxGzc3eYvVbbqOfnJvqYN822mxEjCNgXFby0odbygT027YzWXJitLobTxk
SaK4K46k/+4my0hgadCXTnmkV4ywd/wVKZxcn711SYjfNP2cpDQELQuC+W7Xlm9ITGH0HuPLoOOw
ybB1mwakN8He3Hii2qztEjkW7tbwA3X/wUKcEGVFE7cRkAuquqtgA/xgCXm+Yn593xZetYwCF4j5
hdUwkJYaf0lQyIR+XkZRT5G66k9SV/CQ2VMnurEvvDd4Gl2sM1JEWsYptWJNGKz5gUP9fEGJQkW6
uI6rtnTennTIXcK44poVJK6dcZHAUlaq5Gjtr6tcEPb6EWVPia89ieTQorv9dtDVOV+/aQqvKVYp
i0d4GLfanf4A0xkE8UHlmsHXNO0H22GqvrCF0WRoMMeEJNACXiV5GG/b4tCq3+gFPaOYjoeyvvsQ
BPnSruz9c7Uxu3mQVTWjAS4rQIw3UiCrohB32U3kCKmpnVqz30aCJAJWbwPcOdAAeGszSXrVgUF5
FrCxzyxTYBWNwguM9n2aDZ+8Ze/hyMdulgLWmi7W8YzyoQJgjpSqHslIO9TBH0Su3aN2ARxzKEDx
C/Pael54f5AEgeQJuWj9VkM2DQpk85ifThs/aYk54arYWznE+UDNdJN6+0iVi3oeJB24HSNZPoCv
pPzwpUFyaK5ezzGJaz6RbEpMNVfduumz8hA4bOX+2wJo5kwSHb43FO/zNP84PISiWSErqXBBE1yd
v5iihkZw2El/xm0rQ3J3tg4C+roC4z3awVNPH7CfQJ3XxbqBw51MnMnEik5jCGNuKLYfuh+SyU5y
DTa0yWlONG6abf2PSeij8Opgyaf1OinZ9u1mL18sljrWNp4FVDlOEDfeWuvQfmpv5wdnxIASbq8V
oC/orPNxNcV+D+esir2HszuZg0VaOPmenatVhoJE481gioqfpAhH7z5bqrKpjkqIk6joUmGEk1tr
YyxbKV+Ne/cr3MDCbAtiIAEGuHWupixLfk4pU19kKRVXLLkrqrRQzOLIxoxLGfY5beh+eoAkznp6
pmG5mPtt1V1/AzvQlEmqiVtm7w8SARkOwB0D6GgJZj8QM/TYHZGooyk6Ush5ibiKT9X+ThjJGYGN
2OyenR4NYLLG+ne3qkvk6W2Y6IFdbKIkV4kmGW6MjxOmLH3BsSiVDsv8ktJPGy70alh0UvhuXFW5
FXK6i08HTFS2XGPvSrDfNWg4Yqz+DFCeuignDVBWnQKS1fFz0pK35CaKeFZf/ZHdqaDxcCl1OL8C
gXjnDSFqQCkDHC/IjsWkTRcc0G4Q1NndBom5KvL32YTnjtR+LiwKMov/5WHIZnJb5gPchveQfy12
e3BCzPpyVNxeG09EI4ypdAwl75FauPVI1xP0FIWh7S+Y59zfpNz/tAZoH64U4G3PggsmXWBcsHjZ
2ZzgFEE3bL95Ywfgm1h5f9FX3lGgETZNgdw/ikaX2urO+wQVBOY3yUHgXIbmQEe1qmEoDl5ENBgz
W4QmZYz/79WRqO5Npml/hTwRJGKBoC701SQf2285eM73EaROgbHls/Ia/PZb2w0rTmSdbHNa/IJ+
dEYbzeqTtK/ShF8OtutAIat0RkX4nQHRhUPaY6njNJiVPZA+j4s++cWRWsE+Qszm4YBJg+9UtL4S
KPnQvkHl0RWJFjn1nMDGO6aNSweCAxplYzd5UgmoeviY8MmHkDgqx5AzDZR5wOK9lvWLjenh747T
NrgrNlgjIMeJjscDq5FZwRtuNI9fWegSsRo6s8+5PrPbZ9GzSjQ36/OnQk9V/j4Jlyiob2z/r7pW
xKAC1iQM+YKSjHstGemQ2dWHEiYWKVx38RmGi+xKijueLrKG9FdELpWtqF6fLEbBAgBYR1XmQhQ2
D1QcPF7RGJMuqzN1wY2JOy17d9tyGMyYevHeg7rrOa+pHaa5f9wkHcu6lHgoUhVl7zozqSt0J9gC
WyGJ8/FgyZ0aZiDNbvZTmAITMLNqhiaPFnHK1y3Y8+XU5od8EN3DNcEMDRAOjN31AYkTCPQOk8wn
46njGjq09+Bf4PENcLTPHQe21fgIRGd75di9t3e+K/jgmlagkzaHRUDm0djbeeILyw9GhElqMTnN
t88HahmWckhfAB8PAKNdJS5qg1oqsf418mRSLnG7nKh1YWDGWU+crDgcID2/a20ewBubAUEvbeSY
BeYM2msC7g+po3q+goymWCMz2/itMF0OTOj2j8oKya2HhSMWAV1tNilfRhHNKXryEcg99hoCJAr6
TlDzrfqPxd/jmc6s9cMlni/7Ese1zLD8oFNYiEzFqQ7X2LvfTgK+AgFP93Eo5+65xfZJSbLQw0Ag
ym6g2N5msapp2HukmQxB8JMAnTe/18WOy0Xi3/o5dtAIb+7U+Ud7ymhYqmONUYKcxGOW8D+7JhAB
fbf3Ztfl3YizGdPDNc2oDgzNWcr9eKxK7jqeQGHofxp9rip2BrF3BGs77ot4QmgVY+eUXt4JOSd+
JerhJV3EDIYJVo5WkTKKP+kHGhTNexM5/mtuLc6htbhhB5icfsC1Ap7Z9IxEvB+6/C2JSn1XDJAR
slRvKdrmsKWqyyLgHusJ7JoqbqDAAKoM2E6kNGYDkC/umer2Ey+10CDKE7xjB9JEAvjeukjyffZr
9M3OHoelai+2QLp3pjDBZhOpRVGMWEsS+BB887lfaJdit74AK7L/++gPWG+q2qxEj2qSEdCPQ4mL
WHYzYZXYPRqJs3RYE4OSYWRoWAs7F4L38ngsDufuUOUmd4/QifYtSQAorTqM8ezgWYlF/HubkclU
cjVVJ0A1XKOa7HXMzTXS9WU8w6lGGv59aHls3eDx87sFqPfHNunpswYkg7wanvyPLd9gHLU50hhB
oIFJdNkQjyAM6AaxMq5zBaJsiRNhuRf19OAEr0RjuCwrks/2oQ9U6a3tnQvwkercXJM8q/kHMJmC
FozQXHVkMKckN5g3IG7Iub4FBS4AGTylUhfoTz80C0eG9+J9or65bCHwMpDoyBvCE80O6msUUVg4
41uq7w+lT6gsYwRN7/iCabpfmxjbsMHoqncHL1dKphqRN2lWcfdP9vUX32pcgerrKmNdOfHPOX4O
/GrZ+o7CsJ5xsu2zvPwBRsfY9zNK8gqtykVQumxR/JHdoTaJTzRVUBK/yrQzohWVrNy/18mQKjv+
8t9Ow+Uh6F6+EGhn+2MPTJ5Y9ST0+yND0hXMg6ftd2pf8SlO1Ehr958GmRkCtK+3HPO+gsJDV/eG
L1eIiCJnEzPbUbnyZ91UEYfi6VrwNnugj6vqFMNKNgc42MBOC0bSZXebNfgX6gQUYS2ZeDRaVwrs
a6HD/05Dnzs6wCduDVAvySPizGrX6oaUb1yFgGn3epxtGFdoUEwbOxL79tE1hWMqN2jsRbJ1/0os
8v9gQP3/WZPItF6GWlCi8Bgs23lDvvguhpjfebYQiy7wF305DzWtGi5p9/ItqU5KApMrZsi+d/J7
mRQsRXyVw+2NxQYzcwDWk9dYmpKUZMIj9DNslH12F8RW0LlDrz+uKvJxYBtxDOXe6q1uPnb/mzIZ
R91Er/Np/qSRum3f/+6nTQh+AZI/0k6Tpgwolt+pmCVNOaGoVtVNBFibsvK0B9k/yDWzVH3Tpvuy
1nDO1QzE0JI4U/tta3bFBcaVOQIGgszhpFoTxgHwvs74ez5K7IH1SMbKmi/aKqNweul01eFfzUfX
P4WzsrKge2Cwu6xXm+20FV6rogaEmgncN0qd2FrdQPnK1nrERSf5GwlnnEHNVqjzcE5oV24fZpSa
SsLvvWFEGjyXV88FkHCHUxMX5DViLBAJuMRfLiWeVhS0AT0iC2qpL7X/w62Ir1lz1Rug6vDT7gzh
qTDyzvofbKt2UkpftSETgj6QSnHCIatw37qpUuT4GwhOxgabgXasX/sHOHZsc9JV1WOb5QII6Azu
Imh9A6NGZkD9gEoBE0CjsTmJfXlxeY/FhI+M93hZQF8E4lTX86uBQ9nU8HpkAXNIrlDdQsOpOqzR
6psFfv65A4JvSzxz1cbXKkeadGCIVss1DC0nNJCd9PbBcY7wROiZapAgxKUFLuMhRKU6woNYOrvQ
Qu6AK4nAeYrJSOadbaundIGOpd8P8iVMof0ujo8yWU1AKkMbsyIODH5LlU/OOUJw5yK8U9xRCGIE
HAHXhQ4hy9WqnFm3PEJ9KNkaFojAkMg4LKjWWKnjxM6sCIWjWkhxUtSIYxItD0/hJN0DI3NJsKaz
fmo4R9URcYxKQWkpkH6PM3Vo9JQvzh6auf1XayTeMu/vuX5IDFcD1pnmjtC//ha55Yf8DORHyy+p
XwAhxlnO5zcd0NmLvbFyBUvLZe4+eZKQQD1wiV9XrDIhjLhOb7mtpvvq3ovQAVy8D0/44SKMkoyz
geZUQH3CKZ1MMdp90gWnkhbl4HNexD/9k6VaT0PsvSo8jMhkH8YyWJ8vwD1s8AqQt7A1ap+eoQ5J
AG+jgUmGWFqD4wD1NVZz11hWC9bztE6hzZE0lWfFw99mJvhsD6dopoVjcazuC41RPyxh+iPJ0tR/
tJ5j5xnBMkni04XJ8jIdvO7ChwCBDiAx2OYL8/OILiL9LFfzCsVL9xMAnsVUFAC06HpMlsgVEqCE
MD0BwhbJfGdHNPkTq6LeLpeWARR40eb4W+Tqdqri16OfIpT2BmLpIE4SjdV+p3FbcZ7thFkhLJ2Q
P3eMSrogbqI2hBRktuVzdeZqVW/d8r3jPniGYhxAtPqtFraTdA0B7uoXzsqqNi7iDrjT1jf+gBM2
vSeJcOCF5u6s2/XSPP2KIRhaGo9AVRu2TiZYiWySagLm1HoW1HpKjBKm2Ybaq8OMAEg4t+QzY52z
NRyFoZECiXd5q/HTZXZ4AoF7ZnFAoSW/9cu+t+0UVAbn+mcyC+NdOWJpM8Vfi7xwWBI9CWb+Eb5H
+O4dmVCtIU5lMSc1Bb/256qhkXq+EcxHHotZhuKWmQkymPRu4hQT62WFT1g/yBOYAkMI/i20yMVt
2EFCqUbb/Fvfho7qwhFYCBO9t7zOBx/56p3A9KjDmSmjfWZIpAS5wGaDQw38T08hx7Lf+cOOfygi
t/ZeTfifBPrG3tOa8LRgO49Sk72nhrciHpB+pzcl+W6WINOop0gYr2p3opElCQ7JJYPcuHHLCgnf
w4yFJ8ywa5rlIRiiveBv/96NhjwOExE00nczR2r3cbSnYFPy7Cp4x/MMEzPJw1hIIwZj75x2arJ6
JwqsKfsnR/NLcL5JrEbt8Z5j5m4JkroVCErwmBeu2EGmKGPWHouvd/WeQL0R+iwHME4vILu/y2yw
ZFi0MSC8yTJsRbH3YBW+SEd/n70aybbT+3QCGjsFkvUWzPuHWX7hIhTkrMtbsInO7xq+j8Vh3sI0
4PtVR+i+spBaS29KFgiALPDsz7zqI3aDW8SvDsIF0x/zPIfEv0yvT6Rg2m42cZ88UiDr0vLPYfqJ
IrE4ftsl6Ti+rm+OXZXmW95+BuR0o1583mq91VwpIP3/1FjUAaNCfMaczJB8xDzeWu+FWLCJ06Xq
HvnVohpEk7zDahy5cVAm1QT1IPrNiXX8NBQXCBx7AUz7fyvb45zSRZuEsfDOw8IR/tlhJks5k+Fl
zMkPgVFmLO1EeSBt/iNIOh0W86f/wfZkTU7DPUUPsPg12SBzlKdQWrFip8pYUnpwqIZ2/Xss4Eiy
fkdyKQCF7N1pmm+h2tyNo5UYpd/2a8rWypwoe12OAoW3aRwV0DBhT34bDjBneKMm0pI86LL/5pWT
GvEjPgHJa0fAdw8e7o7vxfrAQN4gRU2Z6O5GBORhWTsbjUkXq4wtFr1HHxf5geJDhqoeDOZAg3fX
ZaHNG/dkw9+LTJ0gcs/5/IIqijHx2w+6CUx+fhfaaduaWYoW7tv3lv/lT3Cf7Qs0puy9qmDdqdbL
JkF+kcSJr2y7/2Cgc0ymHUuUd9jjNmeLXKCMc9GQhWpcI0CFLN+nGrgkDSW7MvaKt8xrk8gI2oXV
xPHzi3Pns4SNKM9tWkAbaJfNJwxUMYTBhDkY7rlZyjHQEyN5uvDcirkRaS0usDYcYyRLcuNbPnEO
syePTg17dX5lL8r8TuGWoZxb3GTOxMtFEHenARcbHSx0j8eg4Ts0hzkPfzADwQYuTpHmodHpNCov
YmWzTbSi7hSrAJFJDfJ63G8i6rUJ/nPrGN0EXowKRdltA/wz8Klk9IOXThS75NEl80cfwxqO4Q5E
esJrpWlE7yJyzZ5JaLX5miMv2pKx51ifZY5PVRmbYOIfl1yQY1NA3ucWEA3oAKZh1Dm9IEIAA8Uh
l3ZRc/hr1HxfH0JmuIEuS+HWcOscSgv9yd0hfprjxt3CPc5ffgsYWx9WQLHbPw336mVuknNB/cRx
Yh/A4X4kL3edpzbGvaOOev2nPVlOVleu1O0OlNTmU7S82V/4IHsHUUZQGXdyC5egYqYhLynT3HFW
Vw48CTRzQNwMQrJ0S7l9q061T8lVY5WCtT7qzDykKuZW9KMg+tPn+mCkme5BsvLdY59WuakAhuCB
GoYUJzr+5+KBEYKg/auoYJGFY0bbUfw66JddeHDwODDCZ8/FWBWNSVcPk6I6k88YbcZ/x++P/BUX
WovxdQ9nbtwkskOywVwpAmo8uuAig2z6bCwE/HBl8tWAXj0/L0Kk52kOUooil542EiafLMBNUZVs
8dik+9e4SAtrfHDxNzyEtPi+xNd2IosF6wtl5Sa/anSmNFY2mNC6MNBClX3kUdCx846nlGqdHugM
d3gGe8hknWqOa+Fne2h6YVqBuVZgUuP9I0jGKc4rwPGT8B4eqF3ng088cHqouDIceHZVR9ykmTM5
CpLs1xTZxXpwvMXqWuFi1vbn3u9d574zhKFr9H51O6/gP63S/pdPocYoNh5+AexfrUuxbr2+Njge
KESXlx8f5lMwsA+ZgoCLmL+D/HQGFEZvmzFKBwinxdBDEq6mNpuLHm1q3DGiNgGZf6t3RwGxTf5U
37JHiMmJRTZcs7qnXSzRfd1STdedFpmQXXCgVsWAlvPcMJMyZbZSQsUY4QzbNHuk384GZ1yP5Mku
/REKSlAbdg6qWInmnxi+uivJHm3mXirsXER06fPG4raFfW+QK3vo91GBF/b01SgSvs4/8YuM3vyI
SPeEiUBr084Lqb2OBco7EelZfpZZCJsUjzHSaR9iBaltgs8EaHPIlOs55QcRqHG4ZmCdElTwoPc6
Bk/W+7+TdU4hVX56us1HOajt3E1JfetFoJIJDsJz5sjWYZ8E6yd2jdZvnbKJe66uarxsUvyvY4dY
Q8kCMuX7h3eG40UcnAuQWa6UQbQmU8skcdD9VfvOgXpRq//fErVy8JHVUPSPNTQF1F1ZlXKUph1X
NTN/9H32mZrPh+jGRInrfx+omXWlBQ4VZIDsuQV+790/72Ea8WZi3nuxYm3w+EZyEw2WumTMsmK5
S251QD3iz+FojeTH2NM6biYvaShe1P8/nMS40b25PIUKRI4fD3glP4CvCiZA8leMljnv8e3/vU1m
3hms7ryyEAKbiBG5vfHQBQwTpZDXEcNI/g7sX0CrXWpHbSiUObB3iuk3dxpAsZs/+1Tyo3N33K4Y
jkknYoKzwUbkqgsXcV6+f90vcr9XFEBvXBAEnD3WnU6mjU9BRzMC7bgJQ7DwLi8IMgElsytnOHv/
Rx0ocXR19a0KA5XsJ82fr2xxCPmgMSX9t23RJB88686taCWyULD1oHu4QNKSMzAFp5pTdkzbb2lF
l6YERS3gbplP2XtonPPCBW5RngPZ/ngcBJNKry84Z4nKWyWUtUmGXMGHbEUNJWV/rCeR+QEdAmQb
jkh3D6ax4e1RyUIp5M2CjE8idXRWYlP+TlsiT31x1l6FAhYzvAp0oHrWXhu/NHMNyngFSfeO4eMA
DsdEo02jN9+xHpvYteQpV37+Vs5dLwJo6objGrOTftqyf+uMiNeDeFGlaTqpyrCyYxJ9G44+0IVP
tFQbaAkw1K/evigIaObt16VfVC2f8u0tawNx3kdiT7CDSkVeEhTMYLORyKUFvgNx9hAuvD1zEegu
HagG4v2KwmerXZF4hSx/3fB7sPaFrwcAyPkLGkbFnvY2mLkwUW7O81AoqrK617VUtbywBMv32kYJ
IV+sMzTpdREzejTwYktHFuMcT/Jma8Og9uoCLlUMmFtDIQ7p7rX3s1QwrAyF/lolLozRt5cyrqA4
EJ6ILmtd+5O/BLjXUbTuktYfNH4SwM5xgSkVKy0lzl5mH+PdAyHo4LdrjNl0DTqotjHX8CfnYLO9
CvsrV9jOAmV1IunQa954LCBaUNfgwHCFRvhHtdDBc9L+gNGDb2brLZmkFbdhnYyMwoP1CLy8SgTy
SCwfDDBw2VNKbKUeypHHTjMeq10XU0IcQ3cH8Xf9UUKlsWxpkhpj5hh0gG2tIjSkfQfuRq+GDUH6
uhDvnw2T6+8w5UfNzwkD6bIplJgAnRrC7vBooJ5Pw68JMTMuEdBiYZz35ixZBpTKfeoL84dO4THq
5NSKl34AcOonLgz3rjBDgS/F7jw95H2gX6eyjXvbicNemuSAHxyPenyuRN4sp1dm9hsB0uSnU0Og
F0SAl3J8CKWKJECXcgMqO1/EW2s6nDxknwIT4B0HJHQGM8vyfjwlQpaPtAiHsxozF+4fspqiglTK
/RMkgQlJPpeZzgXeta9qQ+AwVTJXc4/ArWSQGEvNh4N2Z9eSBydgund3XeQaBGZfuTbedgiuEiGa
wu2rDcjG+GcPaGGzz87W0Gzhe5/HD/gYXuEJgnUwZ9tNSIV4lobYvf/IvfFa2YcdfYIDxvS6pORB
EzgL7nGPvyFeHyJ0HwMVKHkZ2Hs/ia9kuVurKpIczb4c6NOWkBtWhkUWsqkyiEbzoAq3KnqyWfO5
sQMNZMK4JpvvBtck7bhqQS17NN64LDV3Yr9KSKU8BlEiD/4UH+0UdL1C6AmbJlsHQjjcxTwWz53L
XCzN6wDYXT75gCDdoSMztCgcIStguRicaOIqx4XUCzpbFqvD5k2wYgO0V9XdW2+06PAtAJJVxm3c
r02dZoDTyetSqexaCs6DTKuvCUSHMHbGbMTXBqe8OQ1ZEhZHR5wyodtH0I81nqyPM9YMx9khR9Wu
ul0BdThEROHPk7ZwLOpfItvu9VmhAY5LZVgQw3+KGKs1fHk59KsOcc+A5leseoirpTd7e9BAL29Q
YCmi43TU13iMDnz29FvMy4Kv/sAUlqsWpE2iuhgq4uiHZ1iQO7t/kTE0TAts4n4y5H0sEjpjbIzZ
35AnPpOL6ixEsqw/x/wC0zbTiHDlK/dVKbxwnYk0nbWb7wPD0YeuG20bjoXdpp+Phh6/W67YTAU+
fPYP4alOE73I4CNs22ALt2jBeq7IiWCtBlplXw0hI0VSq/ZW8L/nWJjzADuR6AmXt+P0PskCOLhI
e6AoTyASqvz7ieLH0gbzZlsX22JERoX+moR+gzXGSARL+Abp4vHWcQFC76C6IolF6WPxfVjm06R4
NSpoEQVmE3aYRliRIDkpXwIJY6fw1/tgOZ3f8qxCg39SMo0nqu97suFL0qcXp2l5mkmFZTw7irkL
W8TZ8wD4onEPuhbpQApmKjntIB8bHEvbfEnT1kg5FmVUN8BWvWatDXJ8igshvZuyKAPTO3rY4yEs
13tmC82nvidbTg+tqpwlqCfG7VE4Yv/Kn4P5uDD7zOQP0xd/lk9Jt7qBcGdh1uGg9HefOaopuX55
c6JESQ5vCG6W8x/oJWZnSIJaUcrZtDYxkpP3zqc70gutqD1sy73EGt+rv17B9oFZM+LNvMOdiU1q
KDa8+tIedqoFmGKXaf38rmBkzty6LH2YCuZZxiKoC+fMKqGk0cgn0JOGwDZy63TKGrEMr0P7idDl
uWA33PeKnVnp6cGemOI0I2HE5R5PZtvXgcuW2z36KEXxV4PhghPtQ6P+tbWbozn5ru2AQY45CZ5s
vWqHaByKH4zVmp6xdkFthzGWFXTKOH3EO6lLU4kGBijJL0GzmaUNj98uvLv/LFVDkwO5JKG1bEj1
UMCLNF+huGB3Q7jnMsTviKH4QEm14IvAg7S//SuboNNazegmvDlFRdIDLX1YcOJTWaqhdIbe8Kba
3AORFj9/dbATXlcNTGX+S97IxU/gd2H/sLVyG/4Jkdk1ASQcpuS9RQUTUGm3+fKZIogH1UJdoEs4
XAilYm6IB6eem/BDEEEUP3KzLXMtUKy/MSZRE9Y5Vso3xX3jTAjlNmKh+FwSqoex7WDdv7Dw1YRN
0XZPW3K3DUq+yFYsYUoYHZAo+aeZfOUirG43ZIEmDYdjnuDCuFsX8ApcAfSfF29jod4q/x2mgYfl
kI3hZtB/3wFN40sRXtEsUYcWAwBZ0zJ3afMFsDmnHzpAVjYXRn2RvXbolu3WzOtTqbYUOf/3Xbvm
CywIqbaBr7Zo7nwc2zTFtbAKfsqGZRWatAIsqOhEIImdq1ZUa61gKkZ7YUa2or2ZoRbaJGWq+uU4
TvlCvWff1xEPQvU4BOE+nd0QF7XzXxGNFsa4mV/jK+FDxAY6XwQFD64MMKwiWqt7jswUoe1wBf/y
euYdHxIC+snUNKabx7Ebze6rH7pqRzqJooTiPuyKttOB8s9yeqVTwZUV+ds+p+JHyoKc288ZVwU6
BBH+wPvf/qXTWPcwT1v8rwZ2doUYkccjpTCGPYiKy61Hy3crAfLZsb5kLQDYC77q1oHqom19lBhv
INWe2uSvbKQYbjnLPe0DmRx/6rVoXfLqBo9d3EWrMRTN7jggf0ecMa1kSq92CAecPfBfVEvYruU4
q9Q+Di+RNvRm0IKHOd7Iet2R921Wgxic/+iN32JHvqcF7/5O2R+mFoUXSAMQWXuE0kn9g9gLo3fO
3DVf/oZ6jQul15/ts3QwSbd+yVINt6K43+s+8CBD0Yi1gcZG4xb7fcHAL30gF9GcJXzrtA8Hey2S
h8cWfA7g2wR+txxcxEor/4UzuqKfGBEPq40aq/dimsUCVpm2BLFR4OBnjiBtZ3AA9AllEq0GtP7c
hExXxRLVoe7THFT2zxGCx9kUZuh2LW5G8jVI8/eIsuiTN1yPXevxoFVAGKi4KbFj0LcXL6pk23Bf
cboaSif2q6VOOSddolWKoYgqI2ZWO74gSPv4q1f1uSp+XwURGx9BeHvG+sY/rpv5iZIX+tKTvYG1
yPhUoITBMdT1O4Gd0QgNTrZukosQvwWtySBQjECgr2DnF/GTdvPig24Y9JI3rf6F9zDBXIC+Nj7L
TMWrEsZN0GabwuLkoyOTEwlDUWZGw21YO4GskT6KEHOC6xiD+dwMGTh7e2KhGnZp3LHjRRe1jkam
JLzf7AMyBw7z098rRK20gFGP1C7BLpm2O5scUIhwYYMAbAYFhymzmsmBtautYROAdRdF/ibMUhY7
amsObNYWHpV/uYb9Na8kU7SMeHU+vT1j2Uhd+kp1C836pw946YPhdOpuPJVLOzO8kJhPDQBuyChJ
ogvaVy5+RyiwfNdp4ZXfgkPIwdJfJx9v4dcnubtuS5yRnypVYPwgi969L7t62LddAAswJmxpnKhE
tFZOz+9qrShxgIx0ntzCGaGFKVj8szpp7SRxm4mDYqPMZpKPF+Fw9LQawQhaTAKzJkLXSW5blDOG
sN2TttEKW0z7gy1lBsYmD8bpwB41V+IFzHUCssI0vjOlkvctOZ54yl7r8cj+Z2Gj5Fe2e75P6U2K
AgnVfEDXKlKv5i48UNriIrgIcn2HDHtlJwVxftJ/JyFlHySSgTpCged75rDtonRvsXyXfTKtVUa4
083zhR0iPNsD06ANLF8S8gSGPObf6ZH9bkVYXJVF4fZ9XXI7EaEbzFcjq8ur/UC5NOZh97FFt+Pa
AdJSccX35y51RP2bp8Z2aLE/b0QJAiHlAOy8Eb6/fLYuaFvHhSTLGRyg+x2LDxd4AOUKYXxxC6qc
MXyUj+porTbfCoV/f0Gp3MdjS+Z0BfJS6Sypg35zJMUBlF8Jlw37oQ8VH0/cj43k+rkQhjgwv9mJ
JPXY3cWMQ6xYqr1+tm8HoOguyJFxZjGsbbFShzh4Tw5s25k/4KhrirMDmH6nWReKPKquqEj8TU7n
6QGPJOsF/3Dd7uxk8PtbG4t+l3lRRR030xPdUrex2TmK7V+k/LV0kM8nCZcKHqXRP/qU7l3mi+KG
hIxewAdUvh4I8vy6iDAJ8Ybu/Zrur8DGRb41cXSEGe3uTQIeRcxZf5IceqggoAsl3wxcPY2ZKUKN
XVfYwgqa706v4vCV9XTlc6ccBngKLfMhKACIcjtsen9nynMptIQhmyXtzdjSLODnZIx6eF2R3hgC
tV8N6BZzSZFzR1q3QR1Xk6/eFD0E7sZkru0Kdek/b4naVwos8OBIO6dTcDgImhKoyKleDM2mzbjw
CNKK0bM+IQjIpu4MfwmVoQeH3mcy5ghPGoAbrFYTTOh9noQYVQxMbZHOsisELZ+WKbzIxUaWxlcq
TmnikEe5FVhfAzI8KH0rTJ48JXjWJrB/Sv6A8D9aRhvo2QxblluZLE3skI/TzwU1czDzPggHFySj
ribSHdSa7RzZvRLCdfvsny/4yDnRQa8sNMtyVgR85WyNKYSvf3oj2Z2EAMaRDrq79x5oh/q7Sjfc
4c9gwsCYsxtcwumSZ3d6Z1sfzAkjobbBFiONCSNq0zvrHy9YS17XPrl+rnKwUxa1D/gmFfPJumm/
jKgDLYOCaIIvLah3qQAYWtcA+bNnMsJ1u9sBrmivBT/IVa9yDgSyH/X/OaN08ba4p9aUv9oLGqz9
Q5rD4Te8/YER0ZHfNZT4uXQNxiNVP9+yraqmiHMBQb4SHR0G8gkuwP+Po6FGwBdaX9EdOLCTi4fT
VKlIBmo+ohVGkRvzjTqaoyIUvtYloCFLrGBTJ4NOKYEfrmfmReSbC53wtqkkOhWJnrbLp3RfRYwA
Y9T6opsJpvPT6GtNkYEgGSChGG9ptfnM5YvkthlBTtS1aF/zb1aw83ch9D7GCbASOgzkeWmOKKyB
iwYRLLiznkhkRouf+EQ7s2bxkAmwNOIXF+iyT5MwK+9b3DaxQHjIF6sAMreO7JX8i2YHse+5PKyC
5lNvAVmz2kLwatq5uNAx6beessyv0OKnHqv3cR67W3+1v6YXO1/133XTYylqHZqtN3+WUXqSmteH
NebB/kRIipF6lXOfj/tGfNsPJBw7cz5tMV9TM47DdMD7MrncfYzyhpMuhukpFZnhWiR/XyW116r9
zoAczPnQ2O3qEdmNV0t4t1UIeDrsgOJw51hWYGjB+BzbnZ8/c0OPUZMNZUHwBzGpQpP8XjmvxcY1
oTJeVcc1edlUe5czJFBBpUU7rh3TmVynil/qVEfONxgrWb+X4FK/pxs1geKp3jexqt+iY8Am5kc1
NhdoYIr2p5CucqeDLGXx0P8P4ni3cBJPZ18Pwo+iz26pIETioXee0rBx6U9P
`protect end_protected
