`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NKHUeXf9YgRiGh0nQgB1rjjGVfs8BQf0rId/uv0Juy2BNZdKwvVnfNrR8GROgukhKhJqe2z4lJjR
XeCdO8TyXQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QxSUeGNke012Q2lZQi5b35goYujUAic4tqpvKpKPcMTl5mk3KZUjjvo1yQPsjV/3SfW85bK6S1Or
cJOvNvUkb1u3yRcU6dKBIPFzuZa14AMfgU+AjJrZ3rQQxEE/D8BwAD6k1jxhCtMR5O8bzV05TQWd
LLfDZqSSMUoteD72Ylk=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ge07Dr8Rd7zw5guwmVnN/cal0gr44oCWWP1MSQCDgjk2L5tYnnyZCrGNnXrGniy6Px82EmbuDJ9e
6rqjpKluDfZ/Z3iYtsapjfSpWTP/wGMC13mDsPwog/S1d5ih58rqRPh2/gihWrIIDh/g++S/TXXD
xRlOFTWTPt6BIAMK0sg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YE7mz+9BtYD46oLTNe7TtgnXzx6xcCpylrBjE1xvXwBfXZVCuMXRWDhOvAkqYEbEqGqVLJFJp/Nb
etwQ0CSl+tcTEnG5O1loqAWn8YcCY8tEVoceMA69YFFKS2wgFFSmXzMbLujDlO7QelJqX2zrD5kI
/HAR+LslIr4hGOLXgRh8DMeY85SI6Y/JSuyR8RW5SA0kvxRdM04L9YnWR2CIW+uzZVDq0GDXTeeX
fWz5kERqHrYHgmSMxASdaVy5KyCqTrXZJPwiRwCnJJBVZXLCgF97OwCcxfT7f4s9sJgYvOyIyacn
FsL3KJMSRallHnabrAuNPZFULOl0IRfuvsy2AA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ankcp/PC3GFDtNywKf2jaqYEvrrE5tQncu+EWtcG4dVwQiRnKsgtPKWF+IUC69fEJ0F+flkzWM47
v6Ti+nj7IS9qwz4BT5LZSOIn0yT6+3BEHgctubNbQX+a7l8XvGVLC0LPxXeuE1idGOUijZBaad1K
8iahOA81epRxAEG1GiXqn0knat5DcymHaWayiE3T34sR7YDc2eaaz33/xpMr5+BaoFu7UQZTCOws
2Q8PWhSXJr49WuC2sBkmWYLo+H2M/SCFcifYmuZqKIvwxNuYBhWLnZNa/jMqNSguLFveTrxIwPEJ
j5svZHC0YTzrVqcBpmtnqElkLd5CR84PrZx0SA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bFKbVJAZVxTmdIQfa18/qOEE6JHVLbD7ggpPpnW0fKfkbpuIApM48Pg1d3swr4mwa6732q6kKujf
Y3lsSnteVjEfLqm6dHPgox7td+pkqJagpgtJ8HKxuwaaYupaapElRQYdJddShH4ZBF3DudS6mluH
8EiRs0ofqHB2BGv2Npt5COSQ348DMkw/y7lK/ynhfKwoDwUPI+5rS03WfD6DMFz3+Uphs5I9CcAA
i4oXOvtLSsjW1oTYNrfGtcYuvWEvQSOLIK992HJmEPXGWDVmVDIKQUUWWhgAiSotGxi3fK+4nCtr
hl59vGDUzm1DeeHm++bIgsIjtK6F5u1H0YgfJg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 765264)
`protect data_block
rvdu8xbroHwXS/F9CgBpSWvvI2kDY7sv/wiu2C+Flst8F37E5pFP9qanTWoAvn7UACVEld0AOwL7
30nt1VZMrnqXZ+OQ24jPsjJljbp+BUkxI5DATr6RlmgIzv426USQBf1du5u8FVvob3wOralrx70V
ZQIdNwqAzY1SVO+4b3WKejh/P4QxqfpVFyUdZrt7mOzlJjam2YVO0cwWbCQbcVUjjOLpm2G0GKI9
bnLFAMH8bznacfo82mFVZdkalUNIoAT7VlT2argvI6j4ow1Q7r7wIFxjDnJuQ58Zp5mbjqhVu1DI
rRU4U/RrDfIFywOZGPrvqx2TXccwFqD1vMr9GhcirtNh3rfgDtQ7Bx4AzhTLTNX1zc7tfzUfMAAG
NuzmJU3viaE4+KXTZRl+kUkbP2lD1zx7/Mmx0pJX5/rlIdN6duk43Cpny6Lv+Mb09AqaAOincy4p
yOcW2YsTXkggCrxOnnUWrh2Eli2KHuBOB7Osv4R6Tuu9zvyiKm1iU93BteO4D7AwZs4eMJ/qnRSc
E1RSrsaFJfHNVhQY4I2jUUBcnBNgRiRYbr7k3+KvB0M9oXUDewx9Q/0jgonZ2iidyCrasDjem01h
B8aDT2xS+reuFEmPpNwMxkFYJSv9sXvpCznZmzUHmtMilTtx/LgtbKGgynWPAM5uEcEDqgo3K/kX
5NtSPDKBmevu4NABqMZDsCfRlw9I5oUNk55XkjYsp+JTuY7yVUAnjIlPH0R8k6j9viNC1VskNJYH
2cP1RWhV/VnyQ6AgrSVDLv/vG3A08Ku0w58cELuyOTAfXtP+awmcwYDjpUkplXnkrzcluxlAfUYQ
yVTMM5xyS3OhpJhc2ugr1GyMpiqsRxTPsdiiIDUc9xUOLn2WFwHE3diIAo4M8dZWFmO+/WNIQmrh
fvoWCpNdrRqolzyCOqrhQkl9GoAC7IqcmYpZMZYItJhnw2aTmVNEyVLlnr3NqdnNaWlbwPWUt5r6
c0I5yaOWu3i0OwXQDtzjGPkgVKY4HyGWNxACMEgUFJPfsf0TTt6sAUp8F4oPavupeAMa47Mpk9g3
X5Yqz4BcQyly/6q0mrg8bboiRcx5efYx7s/1YAUxyfPOlnAj9lIt+KOt61RMEG2JjFkl0apkgo6J
pB6Z7o4P8Vq0tva+bxYc70Kjps1VXyRN8seAAFhUNkaStwS7LS+yVY01djxqqQWJBAYcRcau3DKL
8GRm1FGXNiMtAHqee04jaa7Z/L3QA1lGWs5D7PD7wdHe1f9xN8MRL7kAs5yZ7XsH88A0QY6/xAPk
lqBt/r5nN2IjUwhKueRbogVsENTALM07RzoYPrha0ZhrQRarymUnxJjdtLKbzubvR8GsXFFIjK4r
NUbxGFeTlrvaFSznlLrQCUV79QCMiTucBlDLMiUAI/6JUH9FaFzJ8vpXnpCpKXkRYB6zk6BkBq6c
0kxRgDXqWFjr0d3QyGp9p4f9t/X9OmmNFOK079EN2CJ2JsfPud6Osa5Di6gIhaROp3w4lojKVs/Q
PBf6FxwbcNlGs4qVe23tTjtvREjQWbiapF2r0wcDIxivFo+GkZwwSDKegWEgeh4CAS29top5ri4z
+p34HKK18ZM64rt+q+hQJvsgNj7tqE+AAjt88v/vItVVTc8mHeyFD1B3JAJzQUtbXYT5ymLL5ViY
RELR0aYm9gIUPjX2EFiqNkH3KMa4HJwVLnY+mh/Y6yK2MQSPztQ4g9GL3CetA1THE99l3JkxvrhM
iirjv4VQLY0LOHxUNRISlgXYmedUAghn6FPw3SYmOk+R5cTyXB8wea4fv1E5HiOnFsS+ZZWQk656
Ke1mFi4+tgXwz0wmhn/rDRXtirOS8U1pHKKdQFQgKusg8iy+q1IbNyYfe5LUS2gjfn9rndBz2IwD
Fv06iq2oosBg35mz3XwW6kR+ZeobazJ8AxAHw/DFSz+HXdYliD7EqIdxgDJfql3yOEJLCE3t0vzb
52coJrhqJmn+RfXVNpaZpmoT/wkH+oqNI+Kxx8BdFcI3t0q4RlbBiDXIfpyB73ZtR/M09R5JLMon
YBx13e6Vj3YBklxI5aKMkQezhQ6cMesMH1lKN9kcMGZHBK6cr6fa7PrX16z+lyuPRWQ2RqGuzkZn
bmCVy0Uya0GyX9y0ZpbdP1CDAememYw15mXdhvaoVKTMI5rbc/AQu6KQg80gQyhGIqif55/IJ0OH
n97plqZmvM352Bs0bD3UIJaofR7+I+rwBI5PquDQyUartqCnHNHl6bjECYC3ljfbg36ZDjD0RRV7
DEW8Q9GYdDs1+YOB5Q9PmCcHYcpcwj+Bse/kf0gSSQyw5jaRCV6rqdp7xeYOgIwuEHUi9+DhJX9K
WHwVw+dEaYaklLKPMwWgkwdCNWP6vw5LPGV36x5Ez5v+AgjcOs9RFt3F/uPfdw9gBEUgpmVUNoMr
7ANbtFIqNSD3YxwG3+qkdOk6eGtaoWfz/6Yb0bIOI0iu7N8UwXfOMZKXhobvdYS4v+5u6NkIVaBO
IYndNL5nsJjDHEzq59Z1PHQGToOw1R22i4O9nJ9wJsBulkUsIWi8sWUgmICjemJZSl6rVbHVVzUj
CCYCHRhNgVR3xCuTKBjOGTMNGo4pp051srvKEJCr86ZuRo8hAfo+z4YRygL5IFKzpdzXB83PKWeD
b6PrLGxoNkLWbk2sS+NFemzyidLwQuo6DNBiQIvHq/4Ltr1HEOvLz1FmP0RH8iUZbEd27hL44o6/
p4cC4B1H54syIyfRuezAfJ5T9QcXz6moA1cu1kC7vtFGAMDc9dsYLHDDLYUOSyUYGlsibDom0TSs
XHvu78GGmdxLa6JE8SUCaPZ12O99+GAW4JWF/0Z984AsXZXtlb3o57XwTcUifF4cFTWwrqoBgEHR
GcJlnnsv899FsWEPblXrxS7L0Kuq4/7OKtG3RP/UDOIOGeGjbnMKlaT7lc5MDqTrM9/BIkQmQwrP
2tVlajdTe1ZSism7k92W/+EtmqcZD/i0robqXnVpLJH8O8gH9D2EorB0H89fr8xwVDd6uKz3yy6Y
H0EWGnKO6fTc9yp5Qt/3dPfuyjmqxEjXeVeJ+qecc8KscbA5iYAlGBMV6rvAZkA8OXVq56SKsX2+
98P2pqVa5o8yal5+dB2fB7PVUwWdrwns25g09lOTOAr2dOr2NbgU2atR4BRNv+ExEgniQ6nIc1b9
fMFOn7A075W5kTE0m/kvERgAvTlKih2aTxMYSEkGJtvw/FMJUr02bJxP/jgBaQ6mY/qOu6GefQGt
X6PCCcslkEb8iRDJKEdu3uKqyswFSOjUAbPR2sCZc9DQDneI5F/mGEf3+7mzJeGTPDo7OZyWMAWD
/zUaet9+9leTubA8YWBHCkYNN4vx143tZ6BpxyG3eB38jYz/kBi9lDsTsk/InZMYsjYBq+sxj2bV
GzSfCmuUiYgOg+kEOVZTj5yNomPHiwZw4bnulIRH6sH5opfWQ6ifhhnNm3DPv0ky+cGkfjxL7StQ
qH3lbZtS6V+P/FZ/3YRbU0O6h5EdaEETHJXv4FYQ1mKX1sFxtdoPs+6EUG8n70ChgwqU1m/oazwP
LgTpjYDaSA0k0K7nMOb/RU0OTMvAO5yVZGmwGr9hRcJ0ZJMiMYDXPqukgwKAyTz9F4KwtUJuSE0i
ZvxCntT+r9hcB/r9Ao2z3G8bwOwYw1FAMOECA5aLQPEmNYqngULRcG3nIeYeyTAdmZOSvGeOXPpu
Oii5V3AkHFCLWI75HYZjNprweKfNftoFUx+7MIg7QBjc05qttOofoDxNQjlJegCGRgarW3nvPJfN
3johE81uZNoaUTUtnvrB5aEQIyxTyNGDXF0Xyc0bAupkawLRLI0qXxjO8xMKDIQNMieBtLSSJoNj
ma70tWdjKigjPKLS8e35b2nnTNCEBlBZ5ZGh19McTsJ55RxTCCwAvsTAprO4p2dY+OI2MSU+K5QK
Zl9TcsQhmSE5kiWz2IO7+D4CGwj0XSDQ53cE/yDpCmfbbJ/rKjBbZZJFKdolU38k+7bEyCEwQWSK
nrd1AyQi5gz91gLYgUG+5AUFdOfaZfxb3w0oXYl2AmvFvmIcOUFyxzPYa/y1X588wlGEel1OpanF
WpkvfI8V5/HMqMCzgdSJH9s5yKDLo+PCoxwfdxbvnxFJxkZzj1YUAlo5AHe6BAoW01F8n0fqqnbl
n9yUFKZvvSbOY/ui5z2YjYtbYqjhDfEBNfmSz0bKe5kymI2YieLZ8rBT+WgPSgD5K2Vh5+c02EQp
efwvncNnWx1muuAEYXb2pS3C+YJ7MkuA8pOzgIFWEo8sCUPuTu09BuzGQeDaiLykQYXOF72rMnnx
VjWkU1ZJQVu7DEfQJuWtcNzR+OzoSwD3d5u+qNH9Krz0O+r4IErgr18euCg+Wsw7fzqWwvTWdc1I
qLWCeEd2nO1GuXIZ58whaMVtRjBv8Ea+xOiDOr7v4PgeRC2JbH0dM6mBm+hMTeeokZY+jsIxhHPE
wm7gS++M3Rsds+Is1ze2JKCA9xomb1npaFCMM6u2g277Exgj8VMMKSChlVG8QDqmpRMChyuuADoY
0OJGC0vsi5rfX+1UwxebWGMHwo+NRj4eafkHTyABZechB+lnMlQLQiFUNXMwxDcEm4NniK5efBdM
HUstRYk/ipTJhiJ+pcEHStswd/ZQb6ag1r61W2YiWbz4VV11YofLrHycSKDV1CK3b1QsaTw3s5In
I1zDr6Eea0OqAz1jr4Hp9A5ClKQC3NVEfRvKO9jrBiwKYEimIC4hr8r3yRGwocXq9Vr9EsLaLLvL
JxfX9pTM9wolyc2Bl3mZIRtKpQODSgsadmBLuf+rfdCBkbC/Kq2DbYrsT6NQy8MXUY6psYYAT6/R
1WJ53of7GQZ6KsJYgAB/y7yfq/mTzDZk3AIBVNFnR7DTi69anlmYmYQsKMvqDed62pDxcCp9VvXS
jc5xA2TBw80Dwm5vRDE7qmt3F7+UcEthqbaLnlg6snyMl6LbTjgVp6inVnm7IkpzBndCZm3dlWY5
jcL7i73aUxVDWm+QqbN7WU9csbHr9ksf/9wOjzYMzQHCKXV+TIalWoRrOV7IHoswwDqKJoHLbWnC
ICcKpdNE+vDxHEmheOoPtABFjynJxi7Vxe2jtd1O8kLseIar3Z8SmfJkkkp7JIkRMHrprFkXf+T8
mVHf7hjRtufq766DInwxFHLWg+Fj37tcJ+AXl7aSAKKGCyvGrUjwy9P1vWvri1SRP1ps4PeXqmR4
cLOEV0tjC1+HGq/8NYWI3CBWcFbNEfNLzwSUapbj3m7qdCY0wsCBeDnZwMmEAeJqb50yeEiv4hK6
ZOIfFU6x/aXtsLfPqM9YkdQvGXxPA+HE8FHk0cweCLvKI5sO6eUbnLv0RSK4dxoXjpim89eZL8Ju
cbwTNvmnf0kOSZ80w4cack0EYqEbEUhGnep5zeydaDQnDK8KltbMj8fkt36aA5ehxIkTaZT7gcka
IcSNO+i9ySoUb7JXKaUf4yC8QDGuGRU4Uf4HEMYDDllM1V+d5e6JHXLxH3Xu+M82iotgoVcmhxmP
f6cagstHDFqRvVIEqVr/fqvzv0QmedR67j22OP6fn9YTzjEOcnCAP5BFm/qKKzQcb0w/tsP26dxl
hY57cLkGgPPP6w02JPToRhoBGgIw5VwNpKttkVwOQM6DxVYerUyr1MhzwiJt9PmXUIBq5+vdinCv
0TB2GCxe7eWOPaK1Vol7A/xAjTNibfu9kqjm+WUWgDSrwFK2UkUtZPuUU9ZhnRZR4QWIygqYfyPm
kLWcYYdqL7d2XFoIlWH4XGpx25IYFurpjRhGt8N4Eq8wkupr4LYOeE2dxcZvT+MTb+lFoHN7BKdp
ix1bIsw63ryndl69snXJuelKIxgrECb7i/wlDOfJ5WSIXv1pywtMGG5wpH0Pvvcqen9OWrTq2pdC
CaKdpjscQQxvatmRPWdfEoWMH7iZs0bJYeE1ysjV97cwWTsQkdqGLdtaurCK1Zpntr/4r0aKm5CO
ab1DhZhnHRmk1nKiQJIf51PavfYUf1c4f6TsqTClAmzhu9hw0h/zBixeyLG1tNl/IEz0mlQ4lLFD
D6INGcdFre/ApbvR3h545l223+kIr6nFV5q00JKmT+tJMCDCIOOyWn0vUP0s9Cwa6JtTB7sokFAX
EOtzPuGKMg8x5MBpMBx70XioQtl8yu9C2FF6R4DBPMjRh1SkDHgRphmwlWuJNkp+RKHkW9rPrgK+
ycnTtoxIfKsxlJ8YqOhSNTkgK27tWzKgFsTOjnlJMyXVUlVuFVchmElH8pgEaExvT2GnJ4iqrTDA
0tYXNULM614G0MXTFbQEBLlpjN2l981UCud3DiVogSPbHbPRPRiwsVlYwtNNRDdpdV2SbMAJpeDY
834sCnpWdTU372wjo5WP7abe960EHXe+asMp0/CiPW25erNtvSmuApEWfDswTM8ZpS1mbAMQKihD
xi2vcdBKPvNBAqYzH/18uxZb9KfrEx2owNOnEKRZBWhgfPtlPASBkjbEw+nB7xRWLh1K2wrinV96
lYOecy1U5V1vHcitCUSWromyBI/3MaArLhh6NJ0HWSC3qZOUi6pMtE/LstdPHS9h1FqKW5t0e2YC
QlgA6ODKt3IuHgGfgexQkQpwranDG9jvAQ7p87I00OJQquG9gJdZ4+QljCoXLZo1blC8hF9ySdzD
T3gjFhtVLjGs74ksBRWquLiUrAJiel+lir3UrpeBhUXAFKGDndKgCbMki32g4p36jav++9D+27Ho
8nthYR2SS9ZVirHmFVopzvAuOWoIdBY0z8B+TXLP4Oj7nx4P9Thhl884DppCFcslDIZyPsh2sOH4
Df57acgNRntD1fe8n4wvqAlrZgtu29jGIauu/mIakfFlTAT/LjTMCzJgtbd9BAJb71M0QFxVP84O
2ndQfRfM7d5gtTn49XLhwnO9FbmR0BnXI8G9MWokQC81nwzl9ckBesuxpNq//aJK2ezHYHMQ2jN1
qAk/fdbcz3gHrEsGMEW5Ic9zSd3aGSKW3NUW8vh4thu5BlpV5BD8G7AwVUbfYUuwVrr62h7RVFuq
vtwazofPdWa5CL7IHCrDd6ERhRIQrlJ2zfvhpO/cBJ+iZuoZTIFM1cur5SND107MwV66BG7FkVGT
pDKUTMJzYGjzS1EZSrRy/Y+W+MlTE1LXV8aE4jGTJ91x5eanvBfLzx4hhCvDlJaX8OGZXWjLfW5L
LDAJqtTT99G5M/HbFxGzbGkyzcPGEKzPzUZIYU4+7WZQxX1pmZZTGeoBmiHE1YrpMPMb1uKh6nHT
QIqYyl+z761IlOLBNzhLhQVyIOhJoHdZrVxjnFmMTTKajE4HcWyyXaoi8kWAAZdMFPonH8mjj8O5
uDnC9pQW0//Kx01Su3j/2zZ4g7LkxNfE+xj0VE74PR8fwyv8jnm/5IBazxGMn788kt9/bUnbgTYY
qs8DkPa/kj+D6kxPTI5XSOSZB7CLYwt+Y/XEbd6s1r+oVyMFBsDEBA5IlRu83FA5HSTW074hz97J
w6Ro3Ey27uZfb4M2Dpm3ap27CC9jqLqECrK4FtbwolsdyCd1P3Y07SkxsJfpR6VRupnpa3g3d0a/
/V5wxN22ptQDTQVR0/ZTktGAs/tkB15GItmhlN/RcISWnyWhR9cynloh6ff9r0Mli8T5XsCw1MzO
QQYyMbHFeGwEdoJKKAcU2y/YO+cGBhrKPkcgQxuql8TALgC33/IOYxOCfSOxdLDSAYYa+yVPTE5R
ei5EffeydnUzX7OWIsKoPXUQMKj1PXPWeg+NgWFYEuJaenPpgMy4D3mpjQTtrg34cVeDJClogNy9
4PUFIsFiTzuvEzMP/RilFy22IdlV0Z5PY8iCPX4yA4jydx1zb3MGMJQEWDECy6vmhFMMehp9F1JC
qzPJ1W+wGr3D7C1UE1gX5+dRA6c0ogeoxGIedNJBSt703HHNUHA7TBrwCt1OFJgvB7KizIpp8Tn5
Y1Khw/cagrvPp/pRXUmU2UQVa1kFRRL1KeHGDE95ZlmImDLncxKstbalQc0ObAkA/ilgsxBAQGmq
MSTi1dOxkXizn/RplQRbuakDTQ5bMtvDEJ0++cRb3h91qUDYPOBGTwBuuYCvBp5jr9gRPIiXsJnc
liJ9/CPGkwIsLp19cbLxbBzOPKNj+GR9Gkvf2oy9W7JUlWvu5ZuW7UKPQXsaLjnjxmLZfqt6hXXM
tTfOpHFQfTY6GleTZk0sqia0Wwg7ofhcAUlnYdFCZddTvd5vvlZ5re1SfxKXVJKGenVGLvdLMEoq
4+H5XtopIZhlc4JF7/SCSlu/iL6gQ9jzOGx7h0JTIOaGINhX37/9jRtFe+CYMWtN3OyNt7YLS+z8
2VicpITtWqYeGsoIXa5yMjy29e6zk1/GeWICV3FRIL1O44r/pgqS4e31J4vgfBcyhPMAY8nvBILK
WBNwk3ni7sHr+8SiZiy13olr45SvrDXMX9Sj9wD7cnVywphosiKiw4GXeZsZ6eFo/o7vL6dXBBaa
EzSaUDR9RovbWGgywKKPBiLHldb6QKWJaP1/zneKTjRMOTsJ1K77pXJUAEc36D0S5VJmErZM564i
rbfP+6vaiCYM0aPeMQhDvyxm1B4efDdPYYwgBMuLyFug08dkulaIf5sBAl0+9yq+708DWcZF4PE+
erCSnV1VqeK3teFbjpt1G7+1P6qL0b511MF47HcGtB58VoqrntUHkRA0It14G6qPtGIq89s/L1tc
8n5vZM3mgZO8SO152sTudiCrjYwqnytYqo6tHrf7e70RToQx5RbQ9ZY3Hy12TzovlYEAF+uFZpuO
+iFXZI68MBL7JrKciP5ApxSuTJiIi+U8t6YcNZcyD/z0JbKa+ibWrw32HUDEq2iCAfOb+YuRH680
IYU1n3fWEtpRHf74zznAcwws1Yn7oDVfDrQHQBHhVNxQ4WuGVhHrnJ1bw0Ye8CSRAPEIyZuAAcR5
dsysdHo+t/vJ3x7vAyh0wNErT/D//oSomOVNGFgby8IS2k2L7ibbNwxq/lFx50Y7qR1+mQw4EoWL
O9+y2QSZNoL5s1nWjdKQys7dT/IRIog76rhG5skTpmFAIjR/HUoXO5AQzb05dXyG6Vqe9CNzh73p
VhHE/+353SeB6oxfEnufmpC2ekkxTRZPJFW5hO0ngfnlSdFOwG95EmEKf7NjBeISvio7uqXXBqO2
SQd76ugYwdj+mvdqFHYi3l7WHe91oEQHXIZ//XRIfrc2cVPhgXwFvInce1XETmpMknPk60ocJN4E
MRfiioas4q4M9FwbLEGMXcoQREQpPvhnpABMBvuKn+7tYDQRW6iHNChIBDm+qWJ8mR17ipboyh0z
ZbJMQw7T+rAy3lKPgkYoXEIZ9KPH84ULxrRkb/XG21ykreOLzS6XYbibPQQ6fonYUqBU38P93Akb
7wxWMPtSBTJd37u/mU6jGf4EMQu7rgvA2s6LWrBhBtnm4T/xiBTKUgA7rO6t71aOjKJ6l0ufAonu
9wYke4oyXO0Zrk3XaiCRBejAzaJSjZlXPh1LXm6DndYoEwNUVJY6lUZNp2PK33iIpf+SpCb1UOuY
wdKZCehrq8/pLC4OecmDnf0Ut+spDVf/qpzITDBZ64Kk3nu4XEjVu6R0KF1upLwNF8mUolzcoIfv
RPd9GOoaZehTl6Tz1/u1r5Em24xeap/uduq+buFGoHqTZXLzs2BRsoucuHNJxjVw7Uto9DVwhqFB
G8rnIrCPlfF24TfT3/6LkWGpuIRKMvzZb3zdYfXafKQ7w6d5zDdRtmeTIe+0nfGoiCODu+k28Wqq
JmoZdURWb0XbFCnBPpYO9sWRj+zorQm/EnNTfMnTBg1gtvg7GbIiy1Sg1ZJWHNaszJgTb/BJDgzM
ZENGAZAk9RgVr6yBaoSWxUi6KLjMPByNRqedR/fUwdXjUSLH3kv2dLt7C74HYvkXnmc29eedHPuf
mmfyJ/NjyKWwUbfsHxlJ4mNN3GYhznjLvScNzt8bLOsJnh1nSxDkGqb5gZgKVeMxYdUUzM5oT9er
ngRuWAXZBoMyu1gOpavCVes8YD6g591nEE/u20gWpuWMMhCkJik24kK1n15gGr3d/B7zGHskEypK
b8VkbIQ2xQNUj+4zB8WkNTAzqJccdrZQ93FQU1SFE4pTJAZsCmjGQMlCcgHfmMXtuT5aIENZ8KSb
0TReQoMhCHF/8nVFsvuR9d/eiDmFX6/EJB5z7nRnGJUKw7xacRJW8VvDzr9RkJpFRjm/VKdfBy6O
DrpCD9wAH+RkDwawk2UxKHUS0HJiR4uI1cqeS9zOgo5++v/AuBUBlOJQ5z/EDZK31DbqKTCuw05k
0J2TG5tEJu5C6AEtZlMopN9La+z7cF1P++E9hHm6ZmTl2vqeRH69qZ5T+P5hVMvkRN7UhFUnWJd6
hlY1kKPL7Kw3gnvHDTuuxRxEFQrNsrDwyHscjo0sy74JaKw5MKeJZykO7b3U61cKCyAaZGbxaRuw
1yruzQb8hz7JoAUqHY5vXxuKIyPRUdREFWqWIXaZ+ImrEFLDNtzGrilPj9FE79RZNXMEHOxdCRXj
3IjpuKTUYL0kZVu+eMGJweBceoEKJaZtLAsogeXFBLLe3dAD0dddu3LRv6g1xa082YMtl9SnZcFL
AVLQ1rp3swJW5Ycdnn3BzTRFFqtSN0fQMV+E2Hi0PRmlctUhezfmYtOoz8zBNZdFN5/Mu9S0hbtD
T2rTPC4DNZwnP+cTw5dqB74QgVBps8Cf/OUitoGd0RCyjP6iXDjxzUTOIxeKQ0/p/gwym8rbOyUV
Nia9BpvOZdfrMImfv1eVM8kHhJlbkvdgl0hbajE23O0EVuGlPhjwTLihBF3tHsuJeq51rwVyB9Bs
GRmyDqYBUJSz4E2kZMYugiyc0z43E4cr/t3cCPqej2b0Hq3ve3nfQ4n+JQ2AR7iFAQMr4Hr2YqyW
BprVSkXXpDpt0YYqhNpO3ikImFMUe2FvxVUQRbTosN1YSPjqX7syRpdtoZ/hyJuoT0cikMVe+Iu4
KA1E5LU2MpRkoMOkP7lONLsZMGMTaOjDrvJf/1jG4domUqXNBIc3cDUHYVY+sbYKr9hrbovkkIA2
d1EsOn0g7ceyzFzkhRklwCYQcIEagC8ZJUubKGdapqf3ow2ow0qBY0QgodpulV+/TajkNs7wd4Rd
Fsh8emnhn58ro8V98Dku09vGlMMgZIaaRqF4uyfDpdZZYXwrGhUioXHnhWRcpauPjLLkhF0+THgU
xGW0jt9GnkZLqIRpuzVobRs0XIOz1WYnc3sUkHJP+QJy/WRBplAotsqu84tKT0RvP3GDEZkEzXb0
lPp7I183eVWMpYnBbamSKJhDn1Lv0d0fqYVCUv0gogv4nCSYFYzPmO8m6Db7e+kPAU0ToMvlxNms
eGifcOOIP7sGXXrzA1ZdRHt1QNqsZSoa5OL8eRvlRaB8M5Fyq4J29/KMEZ9mRFXj6y0i3wUJtd2V
cLl1V+Xc4SOov3MFQrtZQNCv/BPOptCE63BFoiVUPLSI/6iPtam6jJkmLW/ZIiVnbk7Oe+xr0OAV
YU6JmZ5T+BxFlxy5XWhonJrFPbWIQ+qT7sHM62gdJpmmy66K3h73s/7yU/gs3kJmEUzR4x9pf2XL
7NR5rVXLtbIYKMHZ7yNJbmt15vZqZyEx5gDBhhsWmTCtzd+oR8EOqO1j0v++gDT6+DhlVb2irqlr
ohwZZaodI8Jxw3lMh5YyUaOSQa3JsalhDTcAQPL6LdN+xbxF9qxEuPrwANt8u9STeKZKTirFw4Wm
fR+xW6QxpSTm0V+RYWNJX9vtpcqqOb5emKeUZOfCWbTKQnwq+z6HQZTASQ8A+Wz5hrKZmJkVT3yY
Rp7odJNXhTnv/1JMVmb57ksQpG2WskSuNdFirSYGxX+B3RVFbfPcZr1V+r5XNgWVnCtSxf5bOfJ0
bwHuxrLCMRo9jLm6gBeYjL1/I3jov9kzSrucwOnnFkUf9tS8a9Tkf4kzb79fTUtJ2p7E/ZUEkHaL
XK98a/P9qzeU+bH6s9Izz+KNnOcvowg5tfMsH+UuWSiU5JqJUKEE0bgxX8yJimdJvkmAVVSsjMQy
0qVnl403PCGPVPHRWOvOzbtjGuM214p9IXdCY5I95Xufr7TdZlDeaTnMcvFCId8TmO3qiRc380il
K7lXYeNkBvZTjyeTRrtcim7DYmJY6wTUgGB0RU/PCdvTdAxL/IB+Wi4VwPy1EMoigm5de9ZfnyAB
V+yAuSW8stxjI1wl5cvD8HfMyV8jdbhZPsZywwkLlGVMPzVJNlw8JCecQj5DDiSflgLxQz3yiQT4
u4l+5wJ4arDpqGuM1JKWrVnMtgDF5v9lUyoY0QtO1Fz/SzR7GdVZ24V2LQL+Xa9zYnGhLPvU4Zv8
avbPdA7e/HeBO+WFch8jkwS2tTQxdgN7MGhRYLHcBRKAIMHvk7HfeKwQlmOnYFTxYTLdGNyrc6jN
qisCHFe1XGpjZcn/MuiedadxJaCw+WfXnaRaovhssyjJKNUq8fUQI/Fu5oN25/o5z40RYsmqgBla
feQCjfTMcSVprhhO05zytex80Cqv3bmTVeR/UR9RMxmmoVphyagcDp5xVF4kuDljcQ6brMPySLpr
LNbcZQp/oNHerRjk/Q4tOpWE41UV5OMCQcr1hp5ksvbnwLYULDL8T6/yG3HRY4smeC4puJeBtPPN
k4DPhEuHLaOjgA9ooWmGbrzdIHjXWqJbrmOguGlZiOHeiV9kqJifr8sujCy0JyYmgMh+9CAUrreh
jjay2mzN/VI2enYmjlE3DBKoNtNXIFDTTd1+hei4qjMQ7iGcpJbuuysKAIJ/kEGwrvWKvawN0Htr
7EJJv2uvA4nCNgncB9i3Q/bOIgFiCqkIDNL0omEAgFY4HvKO6iryy8yuvy+JYxTk/acSu0YI6pWR
CHBS4cnkmlb9XIYwC4lE3ZmJeWYV3RdTcVLUagwtmlKO0Bc7ReXkcxqXJRjPVJVH6Pm/UdLk2KFU
QDk2ysoq9NvZ57dVi2VBFxpapkJEUbTl+E1k62Slk7i4L2bJhk8OHMDelM8nBVENoeCW3tUNnKbD
IskYAW2L1hQwqCqLqaNJ0oPvZmCMYiTlELdeIsf7EddISNT0vjvvgGbdzDUf6aLQ2F7zIo/2F9xx
uLqoiF+5Fi8j+e2cLrblAKMVXQKLYTfZM7xwNK18N5FtOFnEXZMnhJU18o8fgW4y84aDBCqSKYU+
/nsTwoemEVgyB4ZfhRvNj+PVsb0dLIJXwQUoivkNuhcGRllxqtlemgpUUIRqztYfa8LgtaEkbAac
42GcQVfyo4OFsd9/MeSp6iFjQfhV1wzfj5icWBhI7mNAaT1CwxPlfU+xahC9SDwUxzXzEF4jewHO
eTzkZz9/eUgewfSqOm+wZMwVOYUtB++9fZi/QVi0A8S6C0a+4U3e+OPNz1p+kJSqpMKEoYcwLhuv
ov4SqlAQW2X+kvMvL6Kc0W8ZufVIIncJd8r9PAA0kyUmvjWqmCqfoHw8FJjI8Brs/a1eaWBNOQKr
A8W5hG0sRXRn21h/MKpW2Yz9fZxId/WutioGat5khocQCnfsqCIGuiykFEX1hmm3OVZZYYqzWvgJ
7zA/bZtoGAA8KUGbd1FhZF+ekZ0BP1tUWRrkX+DxefHqIst/v3V3HFgD6nNkJxbZwparjMgHR4YS
i5z4MM/oGDbxfHtTvspU5DAWQjtoSnYs5FpBl7wtmrTQHNUw3x1aMclLDey8gbrIqZOiPDQ+Xkb9
6B846Dy4iI6nDIx+Qs8eYL83LWX3PVNIISDx6YnXdUgj3eK6aeY6Nbb84a5wZ2nFfmT9Zd3y7/39
dxA8kaqYYGe7O0rdMy0Kc+VqpSwWHnNA7wv0AeQL/bH+SlZ1BaOsjsCqVi8OEYQrOn/LRP8fiUEj
uGrFOuSvkOvDIOprKNO+1Nz50uDATBHlHK8XzUlfRKbJlokRHzQ54sD58HoMCLJ83JaMI6vjikQa
sG2Ol8CdCyEkZLIpXOmoGsnAxENW8fKhBediV0fFFPS1TBIC3ZfG8R0sSqCSTwRs1fI3NZmfSr9Q
7NEduqGouWitas00sorwK7jxA48i/oIMMrJy8iFs3fP/AFjK051SBHyQ5BHT1Q4ECnaifU7xMiXi
fjp3Q/UMjhs1ImkqbDcJAMETHBfXElyHKr1qnqcXGIp4z3zxSxfvpcYfNFFRYH6wt/MBM0VmJbGR
cVOx0E29hv02h/o+Z8iKUYaDBve2q6Bj1iO579hZxRiu24auv9Nwv/mGilk0ZE5hE+GzWhxIeGwm
038WZ3KFp7kticTqg139rhh9RGitjSaJGuoFEQ5zWEfsKamwGTx1w872GYcJWRANWnmUGCF0QEqA
JUyBsa6JGkx9soxYwfuyLIy+LJKokhDyADic4I6VqbLaXoWoOhze8lc4dZt8bpxlkE+/Hm9Mx+un
ketBNe6k90wiHEmL1P72+CbEUrrrs5uPhVSB6W5ulTM38dXtmTEA3mlp19dKY8V72DovG/tLpDd4
xt2Q8e/XG/rni4ZghT6KPO9W2kbSH7g1hCP5ycFxygLMCmoKoeXVMkkq9PCx2+CLjocm8mY4sFTl
DkljGTT3GaqaODdQ7+XMiV6F3uDxJJHsmWnzouV3fV7KjlUrXR9uwxLXDLz4eZNQB6bWQwF3P8jN
gtyE3THdiRIUps8OINCGl7BVJuceDm3+9+4K/tawrKFDYe/nRaKyiwIb2KTGj2JYsvePrSX8o3Tb
MV6X5YUBnnVCbtk2UX64uDok4QTwCCKZO7oByn8yN06Unc4oLmH06na/9myLs7Whi9JeBeIsMxzA
99ww7k8PPPVr0xIG7/YJjD1t+qhl+AZqnk2f/psSS8/9YnfIZjU+3vRoiwtwFvrDKigs+xKhffeB
oCgiQs8M8JzIo42eJXORn5joSNr4fsXETPL1aRnevlpE9vjVFaCMko4nwcnpgskk09GRiPJI3DwV
ZldwAPIMaD+2oJMDN08HK0YgzgiMbx8TxqHZaDCvjUHee1UVu0lD8yJCNZkMDANxXfRy5yjFtOUy
RQVTB3r5kFZmbR6aYERA0Sbx0vJ1HnB8eaUCiky0zC5EgmZEGZw+yYvXSy1PPt848nj7zkkHI7ai
OL6P6dXymUs3xt9BqJ+NRHlmMwVgdRmZdGyndjl/Ncfv8LuThoZTttvsTf92MdKyFY4s95HWiJDX
MRytpIQgGd4p8ata167qATkMspnzaPv2cSBkf2km9J2o39V+hCn8vSBz7EXt2d0brovqHCwuyM8N
u4Z0Q1XtYhy7/ggBXzdTHWyASOv6ytVKENSMI1UCEXxN78A6jLmd27tg0Tvn31xRd9CDYQcMWauy
29CY2aXWPoUuzCH2A4Q/t3TWycq3aYNjevmHu75JVdSKkoEiLzGc3N8NUlqweNDoKKrouv0dLBBA
KTJHjxhSLMRg9Y+RdjMzoTi4OLKt6k4KyPvmrOtqPdclx7gDdIA+ZbIY/GAt6VBFCoj197Iguw4f
SXdeZ/Aa0DMnZlOqR/DUvH5krMuu6WYV1JUcorlYri0RfVxnKf8kLVgTNUX8mBs74Enve0R/hHzg
mYmn1lmC3M4VZSEJ19V0m2UfavDBgkhZSbkfJXVReKsA0mPZYa2RhqOZxUtAKOvcscKRJ5c0c41e
T2ikIyA5PhB/TRgw7KKvAMfKr/addAOk2JlDDsf7FveBryVDJL+gWPSTV/z2gOYn0nB06dSLDMGa
whm6LwFx4mRh1M4FG5oxQCsLCkKY/Iw+oM7AywOFpTGcusZCNoFOzoYCQW+l+gXvTYRjKcC1aYhh
P/UAXrIh0JPK5KXSsft2G4j4pyKrqgrwLb1LcKOmZlOP/vP3GFgfJHLmlC4zqXRJQACST6PwqACx
OJHh8t5Q/j3WFULz11NCkWE+2coFw9T9RigX5msEVaSdVP9GQTxxOJ9gr2hnU5IU7mq495YSfnwj
9tA8o+vTV8gBNR1e8g5ZZOkf6HgG13x6tX1dOHSc0mi3SU1nym/Ruko0PU9V9zPk7HYYA1bYOVLb
KrBX9rR6XcWziV3yKWLE/4VmmF5quc5bjpvr52hp0j8/bJ2idKqI4iMJqocA+x8RzsLv7jGJeSmG
uAX1zsKEP2Y7Frd1SV8+zo/8S3xTdDY8r+DX2/bx+oAFyffyHIEMr7xgBNPKeOqmmoFhcvmIUmDk
6eoQqCXXLRcfWPGvD8teRyYzrDCwEqENbzs8MzuJnilU624N0sJ6pCoUGdMerUfIsPqsRbat5ehg
Hp8s9g26rz2xs8smBohYb6Pz2rrT0LC7ZK0DlcWWgdygNSIsM1OfyV8BQZbyfUuiB6kGt0sj/+1Q
olmwjF56ndzPArF3OAsmslHTxeqhc4hi1uNexyqYRcEoVx9/65cVfrg3T+KstmD8k8YbeqVMdpqI
ndBwr0LuLbi7HJdoHIe5/gy3vUKf2OMLt2+eZVo9GRXWiFFVDnHAwFKgmLnQLnEJJqlBskiyEv0N
BbooS15Ovu4M7E+MXSdf63Xws116QQGQRMOTez9duRoiO2kN+kPfojy74QyH4m5RMhkyWEP+Ltz7
/6JL2FEiysQl/1ndn03ZeTjsZ4xrC66IKkWsAQ/v6Wu8jAOgpEFP68WVykSDV5LOa4ACdEHS/uAr
+FS00JQNpQtckbhMz+gdDgLHmAofjQAyFPmE0OUUQJvRAtbGzMnAEH3ZK4me7Hi3agdjt+88hRz0
wpV8LfWmPeRn0ZS5dN/UK737Z9zdusvH51Yu7xAgLDmE+NUWkmoxEE4dt2EdTVzgEms4QemUoRMi
Gyg/+BinxscW4UgPYZFINbDC5TeaJ4HdE/6Z62WlQ81uvG2D15viiqJCtmjKLL32ZywM24yimsKa
g59tJB+n/Q1Gxv/F9F/XUcrn3obKM7uxz4Pn/pnk4j2zUh1XGC+ysHCOKTaLgyT2Yrg1fIUQo9aO
UDawK7n2HAIepFO4gxkd/fakaUo34i/sPBcs0ikSdGRexwGmgELnzurCv/nM4u8rUigscR4ihf7C
vOMrZUAUpe5b8RMGSQH/GkAFW2kXO+tRa5AjDzQmhRJeNdWF9PVQI4C0duEaTOcaqrAOSQZYGTpX
fHzWHlHrVsEhm2HKa/ZAJeJmvpKQKLYyZW0QIilbJoUcRKx430hts5kIaG0m5zdpeEa4d3/7I2E+
5WdLX7u9DSRXZUpwpug4aKLP5ccOn6QkR5mICZuqRTpJuEYGiPkcZlLYOHab3g6u4Iw05Tqkyyl5
vOJswsMiPro/bSZVNuErO2LMyprUxsupcLQ1uDJA6uO3fHPQCLxvefZgmLwAIT9vOB5MvbtnHN/2
isXDFk9GXGouBAklZnHeUQL32YAq1zH5AiP4uoPH+xVsa8pM0XUG1i4GRouPWN5hSFR4tXjXTtqf
AlLzWKWzGn9GRDH1+fhJ/prJS2+uMsiVKoOEdSOcHqae+oXfdSE0aIoZlzEpqTa6BStE63vG0zXS
OJHJo+6+89w7hGPGolIwaPDqfm8x07WEhymx14gJ9Ap6uOrM6KaaAyup6iErEPnDicxqP/w16AAx
C6Ht4dLoAVA0gCRXTuRRiixx36XVdKijX5Xiffz1tplzuQcvNrggCIbX8txqGpNOUxY58HZvCeNr
IEqPapWKKPv2THwNPvoP6VRkx9CfHHE9if4LwE5zB79+KjO20nsOaqnYSNGx4ZGJ7AVbcVk13p6m
7TwN7OW4P2I2gi6XQIUIHvmQbHV7Y4Nzutw7t2rFoOc1kJuIz2LAglE/DuZLvnr7nuxKZ0SJ1Wg8
VsRzbWPYZJqiaCtABTBuYCZhfe2kLE+ijOL8OGwc2WhcbGQebWOG7C/1wW206ncN3Yoo+8SxO85u
PpKVwZeKQzAxRiEOWLixbFDg968yDeKMhNJjpfQxiMxgA16yxcszTtekZQZVz2+l31hdXYNWttVm
O6JmykTdWJOO5GH5jVOeJnEa1Jys3PLxYcLricLxRlHcar54X+LxcP7kWu6aPedXfr03FqKM7tnm
pkheAqnU7w/9GJ6FOb1WSeLBY0KXE3FL1RZ4rBaXUg8rEGBxVeg8HNc1zggPOhcaEFyFkwvpj3Xo
9eqkOL4/Ql9Hyk9cV4wD7VUE0LCFWkGBuGQgyW28MkXUXjPzvwRdu5uldeTyWvSBtkqzjH+2TRcX
DCB2Fd31SBgEawjkSIp+axyojfSso1NZalkuldjnqxRzBe/FU8GFhFI7IC7SANTDunBlikeBd9nA
Vfzn06TcMuEBxNneRxny1ci5Xl5vR4fEtHcM7yJqAT5TAopfNn3GUlx7/eQJT6NiJ/rRKTPWBSnj
lhEcln3/G+o4WmwKCN+QYAT8u7CG5ScKrTW7gwge28nn85ZIZ1Mt01NLcS6T2XLQsOrLyaWqnfiB
cOO61HdBvF7YZufNTh5xZjcQLdGvN/KUy4acPAAacVyDC9TAQB2U+zJ277O96gmhDxvpywdtIatV
AEkHr061NKpYfi6Evx+QuqT0GZaHHAHitP/uS7XvB5zphC+jceUOF2pwzBPzrXDkolggDOwdF9U/
6NbdVvBOsdLBSseJsCzTTN9TCJtw0Fu102Vj/Bc5DxsVIpDDWTe7+GVhypyCypOHLPpcMKrvsTzY
Et0bUVWzlGyyTOGTS4BeFAuC4D8w2vCAbLsoLeQkuIIy0K01rLrofu0+x4pRZqqvxGomFlspgIzV
VukH6GH+ausqpEgxO3qebVj4vUnDbQgB6GQ1sKWjMd9bIHZgnCVFUGgL8Di16HSNHfDjaIualxbY
t6qGVnFzFwzKJtj1hqqfGhI9bpWbHNqCdR+SwPo4gVk1HUflHVI8VKjGjC1M+OMC5OTJM/XOIht3
KC3b1BJqNeftau6B2Ugzr1fVo+ntjqatffq0DQsmB5LOkj2PSVAEKHu/zSHtV86ZScKuikTK02tM
57j25RyEFixLkc+dIjgHr0VOMKrmRUEHF8gRfC/ykb14BsspjB2aPnjnRYgUDZTyblN4JGdxic4q
3fAtD8AWWHTU+ke3JQCibX2s5mD3Q1iAmVr7J/F+lVjrcBi1OlZ6BpuCjk32jWt6vf9KbuqmtP8o
nGeYi5Mz/6dc2vBM9WNlNqnI4WqSR+I9DHGSjBLEq9OXqYyM6Tx+ndD9A0Jp1xADwRXh0L92L9JA
HfRciIGhpwAserL/Q2Sc2KY6NXv7hB4jSwsxXMf02i1ldBbGgcBQKAzMCsuwAhaVlp3gIfb7wbfF
f5Can0ZC/HddveES/P5FoLxq16+NH6br5b/encqljT+BGmJVnHo2cPy3b/HfbuU31FPnoqnffS34
03d64OAIH/k2SqB9imTjILAzKB6yQigemzuP+4Ii75ZgCLA7tbCc7HkHZ74XLE20hLdJx1+QdfDn
FJi5xdmqoAVPHFDwzg/uLlXcI9wPyaQFhHTC5aBvU2OiYEBOFACTRQjO8vlje4Ee4E3sXzu8vgz5
YQSepUjWKJYhXrQj7ZPNX/ELGPIiuSu6fv8Qu12HlyfZfdsh9QVV1LqPPAHmamQ01sYzHW1r03y3
9z5CauzNTBT6q4H8Sctn883G08841tZmUOK+3n1CAi1aJ3bTybp+3kXIN9TEo8IPOkhfXyP9601v
rllHxXiX+B/PshqewjR22hMVsBe6JPJwqBeP7u4BiBB0OZzWf+TycIcWzK4vI8a1IZ8HTXgEyIU0
/ZCvT0wtuC+qKZ0nhHTjbX70TjZ+I9FpmhZEXWDhfW2cqs5ofBV5ivngwE7vxIn1azu1rtZCi+KM
+3/4V7HehKdcvUUvbStfpzSPJG4zaOhsq/UNlmy7vP4ptNsqSfP/WurODyVPZzwsuA+XyDgae6UG
aH8atlKvQBqiCo+TW8042y9lzdtmBwcxGRkzIBCrOzB0WJn8J6dODDhQoJdlQV7KlvBokuSpWo8h
Qzm8byvtVALj0ZDOckhXXaBY6b+RIPGy30pVhipYdsHJiYQc14iEPeiMOQLP2jDkeWyRmh6CaIhM
U5UhPZWOG5C+3JUQWnhDlxpHr7VAnF9IpgyvYKVzk0ullwhuMFMKmHGcpN4aErEPjbSGttd8J7aP
gUWvXM/siRoPsOQM6qtS0kcFpB4axLd5iQKb5G0Vdu1LMHUKtnG8y54SN8Ab/z0JZtjZmjuqU2Pf
EHjVb4QOS9qaSVMe+/rmg4dJs6qJG8VxGP/LvnV2lpE9emr0YZk5VjKrUDTQ2f2t0FEedXH1AtC1
ar5CkC7uozJCNmq7V2YVLsVXHYlUGfTjMn3rgk6FRgSYOgFfWnh2t8AVpDNt9/0N4J0Pekp3mjoV
vba4ZI3CJ+nWFfnKBDIRDf8nstnggqPX4tWP4Qrhc/987qk37mMC3phfw4qsg+P6kNav83qSu+RB
Hox4bjjNDXepZahAnNAx1DhEL3yZMHWzMZDe3PnE7Nzp9n3yXUkXWu+5JdaPXHIiMTi6mDxtDXU7
2xbve6mLEhw75WkpuzyZ3HAq17BBDDi9bY8u+Ruy1Lei1C+16iIo2Zw4uV98B+p7u0It65EcQK4/
B819rE+i4jB37jsCm2kjTu7XFxBxa4w0qqEVeQI5TBX9CaJI4dzMZNNSv9p8Km+nybks2K5dZP7B
+KgKE5xXBdNvZzmb38yKCw930yepTU7jXGm6qTxwt+BW9M56Bvz7zIYjCH7UC+K40a3NMWzhbi12
ft0boKIWP+I3jRoeaRKggJt8NcxwtvGX5GBsZJSH8Kv6j9l7otVa4sfP2kN4BvvqnLrFV7BIaJJa
d3A+8LsoXq73fRNAPlmlZKMD3L85khqOt08iIsvOCwRLDCWq/A7IfZLsPdeTz4/HMOOjC/KI1jDl
fXejql2sl6l44lwbZfO6oBVVX5lxjODYUIxDS11ZgCUfu7Hv1V7fmQ0axMdX5hhv+hFlPLGyUy5D
iGdcgoEl0GB7/AT2N71VDc+rphV3UHf5NjLiNlaiYbazy0hLTgbrLTfdguxvGU72wChHwx4llft2
xhbDK57yeWgMLTN+tmegjquhdUtIDRkbQhMhYd1KK4czM8snWbdsormQdUinBq3fSqVX8xiiqC0h
3YYnkJxc7yTTTA+8rQB0sXWOHhPVx/JcTup3pmH1x1R8JXrcGYanTW+hGhga0fatqzZaCzATsLyb
FS7gmfLsSe+hZrVhNdFeF+8Z8Mu5D0q+KaV+HaxP7HzxS6h2YRICHW16nIHuMFrmubGfWzPrIYqL
LKZorzHgzDYzxIbSOHPCIIO7c/hyHT24gk6KfmNvhBvLM6BdDu4GTAcPOfVE2ySx3bl7EeKPnlj/
UhmTg+80POVW7AYWZQX9xPAaZt5Y68yKMfqoKKgeaqpUg3OTb1Ooj0Q+fBeojMh/y18ERWGe+D4B
0wEASemAMnDUbScUBvYzYSQj9L1EWiwVp3ODe6W6hMzuqhhLdXEDWnyJyReRb5WnV452n7lEF54C
xcSDORJbjGxyAsRZ1IsxRRTYBrbDZ7MlUmbM8g7kE0Oy4f0yBqVoUUnGw719I1MIVCqwUXgMEeUL
zaoF+v4Zb1SXLYVG6VHK6iWH0mL7DX6IHWZAAIDsL+419p+ndswNLgYSiEwlNQQhjUnDuabN/zUO
50V6CeluHScp2wflbiXvzNjJFo+2M7Z+klyf0rOP4hucHtfBLlpI9X1R2EycYXwzLh3+ehW0CX14
OxHR9Hs73H0gtblRRP+hcX5YByJhY76zwu011Ttb6/tV0uPec1auFyLXZwyJXeOgz0Zla+BWjGEB
YpYLT/kLuS6ISOwN4FMVdMwbtalhFglNcdAbGGEgOP4t8xem8Z2B63qWBmY53mFCUEtLbIGPZjmm
Bd5oK9UaLOjYUbHlOTYSs6o7NEZTUbf3WT3IScNAgfOO/C0Xurng5Oru8HNb4c0G9H/Dy2A6OKNp
/rOdeY4NjMBg7ZY9Kq3Jz/YMdRyYTeUfcSlw4f/PEz7/V6VR8lpKjSLjUuPxbAhAgMUrP7GWwzA5
9QR4uEI2xIg5sFEIGFDhsYOBOk563czNWhMbUG+F97NF6rhKWiSxpEhJs9jA4HjNDDHjbS33h7Jn
hng6T5MdQiP812C/c/yszCTzwD87zmPCo4v2jTNbXJs8sE+VSQlAmljD3yB8rOi00+IOZ7pPmiHz
q37NT8oPjyWfHtkQ4EhUK9ySDkJkLtDxGsRdfk/E94Z5VWTwakxJiRkGDw4ii7rb8WSInu1l7YG+
4/NGzmZw0viTRsvYKy3kcCtnOM5BL6miRUQXp5OgPDYEvmjCRvIN7pSz/E4E3XtJvNtKV73rIwcP
ORVyku09Rx030sqr9p1AlV0O2eZaAL+YDr0QnuZEbonZjMuRbIODDBJap/4VWVMiGh5tMqKLVPym
kM5le2B8Ao7sap9jEdQYy37gGNLYkA6xPO8ZqIXFlBA6bDTyj6Vw2b36mzUK5/ArKuiBpgjf+A+I
oM+KTr8UAmgz0ALCeK7MIY3uELsHm/nEZ9qCpD0GkK33dwQHN+zA0yJfh4VTwdQvU0scgUa8nWrC
oTafMfIJhFO2G5ua/gZ0TvJp23kGFw5mvdUw9SnpAL5DsSjgwduPc+c8a/XdF8FClP7lF5e94cqJ
PTfVCaBe9uLmqOPm/+cN1AkYmDpc0gLA5QIFJb5jG23w8kLuuSsGDQizrIO5R6KiMqrRzYpLJd+H
ila+aqDej0JSYk+G2GPPGjhrLafO/VfmsvWPaFyP5QlxenxAvg9DmhPEfrc0TxdA/XFucm/4Mp5r
4HL4+Jgqrj2pwzz7DEwLQaOXPAo8bQ4v9hcpNleTe7YJkcHGq3ucIHwEJz7VzaAAiZdPNqsu5rGI
ayEPNL4j2zHYO74h0rCv8HqFm1tm5RhHbEnXyD7FDLpfnMrVP1ueWS8cyVZitvHC5aj/UEwn+nYi
dhP4C5zV/gPfEZv/64t6VYCUJd4cHk6uJBJUtEUOWwSdy+XBSUiCJIQRQpLIf1ayJY12SEhbjMGg
Le6E27SgUXwJRNxaSsuwuXFhzbLN2mXUaxqE+Ezsf3tsVZ6u01MvPJXxCH/+4jPh+1sGMpr9j1DG
WnPvpWkBOKRXusZbnuj1U38KseMHAkPX0Ocs3dVqxOB4ivXnIyupUPn7Jmn9y7W0g8HYIARjNt4u
kRQHxCbjMyqgrLASWdgmpXFswufifYEgjZHxTYJNJYIV71wAXkktRdgMUJwbTCHXycFmiXIe1W2i
9XodmNVDxA1ZgMJa8IlhkRxSLIlL1917u6K1k5uW5lLsPEzgqWcNNqERa/W4MVZvGDAk5Gpi0U68
P7ye64j4wLJBM2RiC1kAQZBRc2cEluWkgnDqGO1BgP85YcARhfxoaAuhCoakNqm+sI2KzvqaWmTn
Q+nNZRAJcT9U/JqnUU8qrNjH1zW9vN68cb7zCCVV2aGuvvJBfvqrRueF3Fh3EirmtdPaBVbGrkVB
6e2zJQnh3UY5Nm0skAv1RNw6Pa4JftDfiVM8IG24RotQ2U2s0c1GgGthddPC2OA1Ow2ZXDI+gFOJ
7n9NEiduvKuPYVvw9sdBkSHQ9V6j18a7xZbPisBxgNgRImxSUyrXBnRIBsfg8Wmq8++Dx1yvYVr6
qbmuHL4ERUSz8R3xSJovXzDg/PomUUPllGRMBjCPJlMtjc3m7frKN+WNoSX7wUz/ageH3wCOWxhm
EaHLGz7heFhpr9ieydetolv2njZOWchgCFn1g6MGtP7kZ6cq3TkuSyC24V6spXawhcpXMB7+oD3i
KWhaePLhKjGYlwOXj3Av1d8K/TqDNnadb9rl7t7y/27EofMPqLudZ5Dgw4yOI1WuaY5ZFGuVnM/Z
U9cqo+NYANRvM2srhBhLjEOqQPvAZb1sOFQ9XOh6gt8soTU7IrH2VDfFrWTtm7VVYiUVZcXnZr2G
JBp5cWVDmMmfx8OJ3GeZ/cHHbMw7nz4hXIRtCBOlAu0QKGN+ryIEQV8zBF9SAUazpLDoRAI84S9J
5xclnWzMwvAtr/bAESjWGp+YdaJB6YeGyKhxN1TXv7LY6pzZ4NL4jolv28QTQRFBn27e1YpLD7vR
8ArmBl24QYa9zi4O8YpX9rnEoToKqV6O+e4yJvI3NlxHSpHe5k4TPugh5ExJ2Gsp5+4TQ5htR8gR
oBfgNpwaonglKYmAp6khJvBWvC2TM5kpqPsP9dSgfyhMSRGl4XQUDAVtTxX5/dWdUDyQwnysr2y6
F+vvbKliUE1YoipYS7Vhf65jwlpVs3SI3GDBQU7LlamwLFOjGKPRGPKO4VKt9XrdmPtbCRq4sfVD
bPISY7iQ+uYA0l7grUCCAErbhDkv39Lx4z2jB7YSTSEaCrOzTRtEE8JZPXTEomOL+MkxcuTv10H8
1t6RslGvYkjbm2M+5AaIQyYO1YxxYskttX5ui5Q7rknpEzUDga5yyU7i+4wpsSdPWlhSMdex9Tm6
ZasGG5keLE3KyuOberY2j/7oyOp3N/mJtFlYOxgpoLB8WxyfEtnxuiAc9INS3Tuqf5619SlMg0+x
Hid9eYfR2ONVgO3x/Lf6X98jE1En5oRtcCjZdBYMqOwG3yilbenXh6VulpAnBlY19m8Z15h7oxm+
UR68PQQGC2kmSelY214VYpoYRQWgNtMXe5TImxytGBIPPYXYSyoVZg/B28ljL7L3SPn6Qf9lZBpd
wSB0IiTxiXSY6RIoyvbMwS2IYQa7vYmhCeBheoQP+7nv2+96XCfo85mdj7Mbu2u3zVcq7h8247eB
4UE6E+UF+Xc3GCAvkuQqbgJDDwVWPfF14kMHC/HKHoM9cPEkTiPhULylzQYrZoD+d9lpUscEab/v
hKL1/w0sxNjMcMSY9FeGBZg9VcMekZmFJyVXkNUoqBaDdCIcoUXOKB75jL9wBU/3QahOnVUWLIp6
lypubzzLft8B+f13u1Th3MmeUg9Qc4/mg/pCAdVzgNZoiV9u0ZZrD4oQ1QSQ1DYt/8LZmvy3pbIF
cwsTVCUTIfcX+Dj7q6O6LnqajkzjneB6O9VYYqdnI+azJ6yb6xmDa8L/v7gtsmlzwOFU+MoaxWDd
mBMmIekMYYxSeDHKncF/VAx6dFsfwjTR80pY503C0xmYoiF81BllO7uNgYCTBKTe8/5Hv9ZEgnE7
31qGOYO80J5h9XuKpDPAnYJamszglqf2276I0W6/ArdOuMyNVnuqifjo7klJ8nqFt8KB2oPvsdgq
vM3YX1ye2VSLsoR3m2J+Qku/FNv2gCBB4wB6Zlb3JSdMRfPlss1CKi4bjE7sQdT0D2GHwC96wk0a
16HATglSqj/ILSKlUzHE7LgiZDFqBS0FRLZUUtch5VbsEOMqgRHNYpPDX30C9U0sy989m8rfJuiq
aBiogV13sggYXADuZ0ZESCMlvWBlAQ1xcLiPzBq5wewOv0BiO8Qas5yBRA/CSXSVLPObxADYn0RZ
tqquSc1kEkZbU4n5uG5mqwdFO+Lkg0jXD5oQKBE6wTsFoQXGoAetfHw1Nb06cMAHKdOvVILATIFi
YqeS7HDXlbfd+cGv5gpQ6qOyzbKg5+VgdqzQ33dGbpDgtY9/iqR8/dRALGgGlWxKaVgiFnKzdZkn
fZ+N3nnEh/GncwbaxthFwM4Mjpf2X/fastYbP3B46GO07aWOB+Xul8Gw6mVGcaP6FxOAI/5zQPak
EZGMY4/Ch/ftayHLpL9UuJeDjRQI1pFjL2qAhf0+qw+zTXbZqQRpPgVZ25mhQ4+ZnFy8YDgj89T4
Cbf5ebiQNUFOKOwIjPctk66Rjdla8gMwjBPsj4QcKy16y9SWUp8J8MCzo3wg0fRzjsZYlHmAI5pr
CdnWjwAl6kEenKYhU/N0tosDw+nPKRJs2c23oOTlfybEA7WKcnbDucLW7YDWbpoNkpncxXoxLRtw
yN7+iYqHfu/yHN/SEVsNJrH9zVLXNSex7RK9l76RPdH/p20MHBxhfptsqSAdcXSPmcEY970vduQC
lB+pPz9L4jbJ5nW5JbrGs/9YSMHBQ5t0igEaG3TuDrYaOn54xK/RKmNRQCfSWND3wVVkQqOUn07t
eWNMgY0siYzgxo/SNDGTOJR4aT4iV02W05PcP4g8RI/dQxzQGK3uceYx5lyXk3ioIiYzxcprrmkN
kf3bths1ioO7/MXosjg7SQDLZiymV6+JewChm9peJwNV7+LSMq/ug42kfdxdbHNm1Ayr/XIwZBqS
l7jSXaFF5K8ovEx6Dh8AY0G2s5NujsavRUIhp9+JeUTPFc4oAIdRV2IeXZIU3R6hJosNgBrH8CYU
ZX3SMp9RxV9k/RyrRwg+/XKP+UISfVSNlaGiMST5Ib722UVqUUAFAQYRmU1aJK4pUDmmK6673Yyy
6iXNVud96y/ap3wZuTt01SODzm9hM+KuEoxU385LZVtQX7P9k+vrVyd3X5oKaeZpMphvJiE0EnRB
fPxyhyxDeJfXum5ioou8Yx5LxAaUIMd7qCqpPZ2ZxIUJ/Bv2HLPbfMjLxNHPcntHXjizIPWAByzL
rcQUFL+e4yNsWOSFtNvNrjqdXvuXwg2lp7SNYkn8DjRvMcCEUP6uMm7Xuh55SFRdtO72RMY4Jmqq
fWPqQOrS627gmElJ3ekJvc0n6B3N5CM4q6DTZDLV6dOaAyTy1mD375aziLXWQW48rd7xmtJt4ME8
IWFWMlMwUFk26BkqFsJwMVa6D+TFTzrlcUIlsP6ncLe0MUV/baMEP5Tm4bdIaDXPAQsCGxAQgAHC
bQxj02dBIupQqfrvSFM9e4XUYRUGOsG1BRiXS5de6LHIjxFxSkgQ82ER6+xG0/fODGQoBL8S2jvS
ZFF3+M0WYwt8wZOQvpgDTGBK9OteDvAzB5PU49PgV9eowwwUnTgxm4jByfT3N1nmAunUqoh9UmkA
5rC+uyaQAugDKCL7Hf9TYKZR+kQZe8pUHUwaKVQW+bVQ6h1NsrAZcyfSpwPk6BN0i90sBXWZ+IeF
umRE5CrP49bTxesjzqEJiOdwFW2ta/y86RR5YtZKlyVv2JWQ4l36JFmU6KhGmYFnYK/Q1oWkNarf
sxjEqSQBBMX6ciywIyUdhSctyFGygWTXKCMrj9M/YIfqCu7xzZ8ZwkrQsNX3B3i0Soh25+YPdPS1
BVQMrQhoYjuWK7t9unXb9Ul/0JLMEU2w6qUZdEIdkvGZ8EHFUmh+LH0GOgEWx18PeDyrwvBJY1cm
HO9CE7jG/zTjSXGPYus6LmtIo7/6ZInLkVCVrZ6wFrFIWUT79BApfyktfUWPBwRcjJ50JkD0gxGz
2bIbN3pJgfNDZRpY91zbG01tYzT4sybrWfrs+wpFjV3R4eogEeu24B2ZSabRfI0VnilHavTUE39f
H5wQ01zp9ZY2fkxeKZd1jJs7R+A8rHCCb5LAZrinRuhsqhnq7SGspmStqT2aSuUME7fhj8HoeUK8
XKJX6V3a5FXcsH0zX7xCGjWYio8C8vBfyo7bnwye3T15/j3gcKKRDpzXjrPQRLgsDTNFkjoVcABW
9uzpLL/arwE2CU7B2dC0udpF4eM7algo8drWoexVPKftXMnR9cpqegxkCtBfTrArd0/4vAsK4FG4
fL0oNyV8NJ0dc/sudqDqa6ag5utfSW668rHAfa6R9vPtDNoh4VD7tSgNXuMjnVmZYYoAFdSRNHTv
5EfeZ8PjdebblNBaQqUhglpcqeju8NWHBYO2GtLtlpNSHKNpecxK1msl8Q5LiAS5lJJ+Oyq6p0bZ
DdnpsAEu0+Olok/YPdrkvZZ2flp2v+YJ0xccH1liE8rrkMYVUPv0g4EpAl+Ub9L0MOpzz+Sxxp5j
wM4OmrZi9t8V+JObwr3YRk+81dRqYGYu2Rvg/LwKe7r/oGW8heOndDCHT9WxGrsHyBcCYZCXgjwE
Qjf9+2MjrP5fQx5iG0HV9+up/ukqjxK9ysW/npSONrLFMZUKwwDn0tacdojI4DYwBYbVO9XxJXIx
owXPaKMDMDYqPv4Emo7tIc4R6RM5VObaMAORPccK1m/PS3Li0HOKeE3tMRldT/sQ+xP9JOrWo7ir
NXCp8px5otlVm0HV3121vLH3AjDEIStP8PE5JjRCfsks+/lsD5pMrObJRX+py2weCaC6eyUkK4Bo
0G/vAQsZZoosu0KYkdAHaM/NWBZGHFOKSBk3W37IFOH8rVU4TShh21ZgOgzgWYucN8SgcSR+C05M
u9GjaDHCo30fT85bdntvNGSKpRq7Fei7PvEKRHdFgrlEcVcvgDu0/tO+xsRNOKI6E1bxlTy25hMR
qlAieU09UQLT38jlAhqHwDibTaPqMkVY4qQT6RAzFNlov/94+xgvfmr0Zd45nvACAYXjeLu43Gx5
/Vqt1mh2+VRYbayMASXBSMQVKcdq7E2uHGqcDVrRUF9smy2pvEtINgXEd7HMf8ncnw5qQVVluidJ
R3aYCZaxaXf6ww8ypqr+21/E+7353gEh1Wyj+98xI/AebgqET+kkFzk+ic+6Yusrq1qNqRNZNhGT
6zONNmpqgIxPlf3LYF58fY52itsSNSfdQdFGL1Uu0j3KwWRSTWQ84SuwWZHht9e47OvlPNJJFpXv
LsX5tusy/2k5Zygr9+pOF8xaRd3epOOPHym8HKGRNOKjwP5HtBQg5KDhgzMCqWQV1pNf2YFTD284
K3TnPUcHanSFXLTUq1azcHzY9OIvnnTf/soIxhxWrhaCKmBYHQjpNLE0VRRVZZ0RaF6E5DVBA0c1
tTU911/jCdHeLOSSBblcQBUZBzhq5z4vM2dXl/ILsY7au6pTRARnG3uFbnoC6gd3Yt48N4Znn8fs
xzoMX0zmTW9jW7A51qijM2gvadrbDQMeUr5loTWDmbB0CImub/7VdwqU7LWYUm3SIZrbfpycPzS4
ubHlkkqSg/hvR8o5R5xj9A1TW0zVZBzSD6fjyBDqol2vv1HFnwy0bfZ+DYV3BEKVFADiafw+73aZ
i/BeLpXGLIwnrC/HYlzglkLjmMdE9Bm6KmDh0AhJ0EIdHebDg0oudeHMXAHs3L8nf48225TBGA0/
19vmtJ/tef3uIZ75VGMVRZFaZs48kF/bQSXN3oEAZzj5HUCNkCgtzilvNMJ83HBm3dN931uxlFE/
eYPnc2nG2zpVTKWkF1e8nLzmTH1mIpXtsx9cu6UNJ9eDploxBmVQThP2qqY1HwYgnKyzFpfznkUf
SAWZraeNV2d1OBJJwarWe9tSy0oBlBvvYSvfY0GlOy177yZFiTd8scUWDi+R+q5e4SUjZe8NT3Gf
Ys6lLJ4lzRjl6VPLR9rX1bY0lCRynevIbIdgI9DzE8f30lkXssYO3shJTmNUpOooF0KfxFbSiqDA
0uzmJ2yX6vOPQoRiF4b5ndb4pLcl+vn48K2aUBYvGbKqHfanEmFhP9mmR3llDXKBoKjvtkLXmDCU
nbwu7cPxO2gLsgiRakOwf3ljs00yqho2rS/2GmLWJ7NryD6KUp7mHV+EcqTAe4JKG67Oz/WLP3Gb
ZRmuTQbfmkoeM5lQ79RzpN+c4q1dbYOgFsf+GKMEv/5AKm+s4hZjEjlHlS3Rb6wZagl1hTg7cEV7
BK/q+FdcEBMuIkM/tfUxMIz9ZxTUx51SoutKlxMQJsb4S/bppHpVoBkdSGiF+w5dAd+IhbV/Zil8
VTpShqYC/MlL6CHPV3Rem30QgmMMFRnYEqAspuLaSgQKFFihYRkR6iixO9Z1Ct4R2OV/n82EOS/v
INe9Aj5VDajC88+FM0mfLwAfBKCFVgtZnZpvLu2D+MyD1k1M/rkxTqEWFgD1WuSGRmhgviHT/KTt
k/8CVb8Jq37M0wHEwEfzjSLwT/cQEteaU/PRHUCF0gX/3m5XqLoJZBrrSOdcrNsl8MYsrw/ynz1X
H6ZdHQHfk3r5QjA36Fm/VbwQU7P82+YF9kvUFxponISiQfo+M4nyTNbN9vWCLuOs96/zrNHD40mO
DZbxfJj8u5RwghIDWOEotBE2xikciU+MxCS7B15nhepEsYnz+HRMWW8Nr3kXsasl3+vfsXQEGDXo
9fIL/iNVVzJDk9Zq3NU2IKjtbLGMOa1F1w6/AHeSNy/Tzk7zFZXp+MMgZChsStYF1KoAJsal8FBA
7wnkhwcGbKMNg7UQQmvPZqpqNd+6AX1h02+m5EKuM25hpu7C8OcPSZbyD9SgPwByjtldMiwSB4wN
pgXQkVcBcAW/NTb2a7m1GN4quP71PRMtr18ByWqIuECML0GxHDgwQi/koMb9H5IO61lvzBe/4eoH
fnZE7K7Jd6V0gHmNVU0SKxMCwKpOtmo+14eLEFQMz1RodHBx2bs/6zVcn2ScWkbk2YJnCeHQLqQk
e35ZlR8TwLjpWdi6wluvy/PHNroTL3GtLoFA+LLYdVnyyXbxF9bPCmK3HSX/54LjQYnP5evcdDze
k/mRPHT26qHzrrda0r+NLE+PNgbz5DXSIZwCivW6+Ei0XZWlcCTKHeMBCwX6Y+VhNLASKsyXQd5U
kxfbDd4CxVHU9kqlVHb7BVp7hkrH0lk6+2kZtGYr1LP3BDbGpYbnPtN8Zd2N0rXN3+dBNwkB9Ojr
8pTOREh42vgvJwyT6fanSYBdpp74ptePamRqDps6GwamP1726CiSH9XAJEmSMIwE1lAXLVwjglpi
p/+U6NEGK8CC+hVvgC3hag1/0Owc2YSWOw32iAsxLen7HI0EVf7DkF5tf9bl/AS1+dAqo0DGF4dW
/vAGeosY8raaZWOsgdtI98wimJXHhfy/6jLWnCZ5p4hsyfwHEFM/czuUiHV5II984XZDfQk28+lV
CJIVO2eMqWlkHTe8gJQfFuEvloInev0GAjEWGl3xi9xFBJlTuEbP6YvZLA249x0JT+/BzQnXHChD
QTPUnBa9HynVBSy1XM9Sit3tS5rEabTQ6YGgTdV+C1kl1sGB+1BiRaRPQAJkoMa4yHjMKfKApPva
0Ly3gec1Z+YTQvTAkAPK/6uR2K2SsdG/WDIaTS6PHVUUNt1Cc8ioGDYUHB6VW7QVa+4Ez8QbqdVU
efKGcIr3GWlcQ1q/GrMT3GOggkqvGzjp2WjGDLqO2DApd0Uk2Umk48p9vGUw/rmwBSc6QHDLnMer
lPr3zbk8TBfilUbvpEXjAFzvlrZYBpyFQcEcfXLvtZ11VbtQM7C6isKr7jlRmE7nqKFzd4EY4Ig1
JjVcanDSmY/sT2ErdI5np/+Ennm6RL5/A8bwDOHCZFKpEfpUxCfLXz1xCw96z/mFpSUmZVTsQ90S
/P8TpAZuScTXzDcK4R2GJLXaIJjpWShePt7nxosbWbxbJJelafuLS+62lGe0RDI+35TrE664bmLG
lryV7sO/srp5u4nNZYh7Pe/0eAFikGPn/Uk3Db4J7Vsm0J2aCbv6ZemwaLrces6qGCLRd+7NnHwU
oLRQENTnphSZfRyJqGi/B11jENSkrgfFiFiTwk3zG313HEfKaCCYBeb/ro0bgRffUf74jgHr52PS
j7Tz+nAh2xhYNFaDLXSKEp1Umt10GnjVY3xB+vkiTi8D/bH78/F3bGCLuU81CcL3NC4w02VWdDL3
Z+ftzw085JoWmMKe/jU4ugAAEuqjjsspENYiJlg2m/38GrgRE3qOiVeG4on/xbQzoFWa2Grbijb7
/nYGinJ2RWDWcugU7At15jmXfl+j6F9e/NxQPtmaOEHW4emb40prWi5HEIjqBO9cg9lk6fBPUZ/O
GRXiC6LFy8Aa76T2P0Zm7vqGUvhuLrFhJT0KoTOSQS+Yxxnr6DHN9M4jCtoQu1m3fTtIiOzli3/U
8eACyU79PS4l15QRQ3iWsHGEx3EUW78+A6rTch3IJaEDu35/GpLP2qxjXi2UPLGXzLi8RGMi19Lv
mI6VfWuY3i4TOS+AXV5t+FxAyl6hrbX3bwAe4DUK0GmSBXycT9vl4GCvYQqajUpmNAV2Ab6UeApW
LPnE7YnOZJpdVlUpguZSGlHpt7SlA1XePuVusfW8AuOB+uk+PWF/0lfaxWy/hcTObUZ65tW/sTvm
95kY9R/qmsbm/zNevP0YCNrU6PK52eYH0hzCpLUGJgWlaFrrcDnQLeAnLIaDTlJBXMYZvedM41EL
yGZ7pOj623qY+jwZ8tMtADsIhFFA4yC/+u/xIhn+Ad0x27gQ0McWKQo4P84Ka8/C/x/pBk3w6Gdb
Mp3ly0Vcnz5LOyXvo3opWWni84YQKqMvSAIfTChoGjF+C2+brS33qL0qdCt2JVxXHSQgdggPVZ4o
cWI9LKMqslijo3y0JBmmPxzfz3NGqYoEI4EVijGd8wo8OzxTuL3Qgc7KZUhBJgi/N019pq3DBdbl
K0L1H5WR/vg7R655a/l/Cc1EWZhb47mzKjNNB0KsyDeTTEJ+nfd3BfoW8pWIyMrF4J5iRvmjPMNC
+cU1vN0FL3l24+GuIFl2U5un7iMQ20m4Xj5DCNlBxD9l9z9+5uy4ky9PyX48DS0SyXTT+C3WBIxe
uqRDoaYtQ3gaYGTzD6XWGCO68mb//vWcDpEv2p4A5fk3oAdTUlfh2YU/M+yxeLgjEdDV+kpHkzxV
N6dgHXtrVPg3mu74lmx8CwJYGCrPsqryRVkvrzOyGud85/KRqZNF943+e63CuqjllyTVWIYmDo9J
3mzulbJZ5JyYNbJ0RawAwx+ZbjvwCeO4AuvuIsSKRJYwgl9ym4wRtS+9leZBdfkcLVFbC2RMuDVk
nro5TNOLl4veeyYDkDpmja3QrkMUQQGkzcTwObaACzRsOGu0VGObpMIydXyKOaq8rXAVACcJJxDa
edpewZUGq3VvbP9o1aQkOXE925IC+EcoJiRtq1sUlk3nMfcOhyUAiZne2Vbrg54wOZuFwkpZq+9G
oyIkJ8ly73auiGWcjxl6h6I7GjBEd0Vm0MW8+fqdQesPIWov7hwSXhEWWit8qWxY2waU9VksLJMA
0nWWXibOJfCuqTIg3eluZN4sukfNxvu32+qQM/l8+RfneTx0YqX0fzHjQ4p0QN4tGB+CPqMzXqQm
Q+SYx0dDbI61bmiv1pm8durYFXTRMyffnHOftJIFH5ig59VphfColdHuHZJoIdROgbWgbCzCdGLC
V+FOTV010GwUNt0DweTE7BKlxfjK4V4BaQhtDY+zdVsAZWnQAEnm52U4dBX98N9aAf2DtXP4A/0Q
jIuO+e1BML615fXvVPl/oROgUuXot/rOOohOJ5rkx9LIadU9H7xmQbx9WEanjWhoa75U75BI+Vg7
MitAM/L/8GCIDJIkpdH4/2eICMw0YpFNvNS2Z42Aj+4PdgiVDzaf/0NXQXPcIB12PPqVfNEJgwBi
MkggJt8v3iefo3GCwYcrLKjqprg2TtzYgihxIo6I5lxZ1akuJci1zLiYN0ZDNit/8UEuTfINg7eE
ko4xQxWjq1uFYM8Bp/ko6A5TH9NHELTPm3Z4xDuMTXraQBKp4M5Y5l7DTRM1jfzM4cMISbzEAfLB
Wwv8QyZ9DscSB+7lBqT0/aLat8TkcSC6u/MFUwKlDdRN1PaIFsRpxb9sIoECCd2Hv6v34Dh4em/h
vW2SaqnUALiOr+hDjtVhz7kIvuEZ4lN9pqKZwWar1QgiJt4sbwIGxejJQKxW8w5TC+bjzqu0Qo66
kefX4c9eiHpgx70KA3OTotrrpPLJnceeOZZeij3T6M8PT3UQ3IHw5NhgcSeVQ9NZ5TN+PRoHaTBp
uWBWynXAerYTjRq30sV8yUct6IHnQSJmr5VvqtG0ydD3mXmOWqaqmAZi36MQyDBpf1tp/8X447u3
0cof0hjukXAaZrF0QR2Q5lytDUyPi58B8aa9JzqYYiV17ZLdcr4C2qpkgcm00Jj3Ijr8kbgxTWEw
caB7LShxK052aNtzrZ/iBaKuihdPjflIcCDfgChPiB2+SF8B1GApQtL9w7fAxRXQRBBHyDf/DlkG
s0HaNfgCQiT4ILVvg6pNiDiQohJHPqtO84G9is7Vhu1PptKtjAe1z5h3oyGPRXwmusFyMBWTIgBI
b1Myvc9sWStgZ7Xr8+ihw93jq1vVO1dyhJGa8r7m+IxmNK11q2Ovz7IbzUplH1t17IwaUgB/YNYG
iKjrqxXw698Fb+dX+Thyuht6j2jGkhD5pIiIXX+DSWZ041yuYw8ItTpUsj1Ry++1Px/UjYoEB/Xd
hA27DWFz7gbmrrlXlrzURab+OiZAwr0wW5uzL/mh4TVjdNiroTmKTVE4Ilq2eFy7Gl1T72270gUb
s63/WLYkSuAQttC1Q9UrIaeYA32U6OzPUSrk8Esa0Z0/OSCcQDlRa1QIMje4BW9ZUIl4ndnkovbq
sRfb4YcRw9FWFRko0tMWp1uWytVmEzIp5JV1BBoHEB/5iee5YG4e2vz26bn3FZGAPjra5bcWIEy2
Xh/vAHWh7ccsv08wlIp2234Q2boUEGECfwiIp9sXnVgNE1gQg0cokc43BnBHOf3BsmVcApb7+j0V
gPn7opC6AMdclEIuEFpBsAQe6I0wiJ6X7Z3xfnUIMjLdSi6HEsEs8Ph1ppW1T7ultek/RhJQ/k00
fyJ3mPtUhTwxwenQz6cfbEfoWn8Z/OdcG+jKb9zY0nmh/zxPX2C22C9huLemhUni+I5pcEa6OO5m
I2P+cVefzU3lNWyUmyLKPhlm0uGbqMrlIPkBbjA6QVMd/lUMC7apOcgdrusaLWtxZVe4wmvjqdlp
CSRh3SWbTz1XrUB5oZPq3Zj0B83DpP584tpV2eruoN3CaOZHDBzHJ3375Oxopa3VooEZfci+V/sd
+V9XpnFxxdg+Frl9dqPKwRsUex3EuPreDVAjfMQzO5jeuphOmlOl4LlFZIeuCp3HrM5xloZ7s+rd
Bs2taSwFBGa8zpaDT0DIILofVZTgmtU/qnSFN2sKkezATroM9X2ykkymz+vkfpQW/3V6jz9osyPh
GjXExs7Bj6hOkgsnmqo4W7JTCSCMu3cD59Vq7KvvZtLaz4MYO7MnNBmUHuQkGivUOWjHjoPdBesK
Re06iChlega+i4gy6fMGOEghrhM3BV63iFHQvI1D85O/BXot+ZPrBkMW02s0tWRfqcZyR7pyiPX2
yCNAIz5BqvBKZfgzgjTBrFLajQ4FSMYJpEjtowx8HpFtpj4YNAs8aJahiKhm4HAz+gyk04/iDWWk
CqP0eKE0j868u6XyYKMMjWBZv87aIwqWArQ99MQ8sVVzkRCb9216308W2neIPzPmct/qbBF/race
l1+I2ZA1B5tymJTTjlHUBdkVeofpNUn84hFlBX8hkegg5Mstew9zQR5RZ+ANRgCQTscef/WkUSK0
1nFqiVN/UeJANyn1W/kQxoC7T0tFTMlsut6oMCK4UafZu/ER6bjiM2PnbPV7IBn+1HBmnUwCRRi0
wn5AKbmFY/CmED9qkcU/1lfQ/eyvKAjoo/x4KeByjgaV0GAxg4zsN0FvO4yHVjcdqSwBLhBPtYRh
YVoLh0oLcgY3Ee/dalwjIyX7V+GNcRLkZ82h0DB1aXCAzS0yG4Pxdl6YvpzIy6HYaLEIbY7MAUkq
3lapXpZQ+XGE1xDdBovm99t4JvGkoPh4xwbrmPuvt8AIFR+nwG5sWM8yhrLcBAJK+w9D1QaPEgW1
z7njUhH4sYj2NYaC3KXy0WDwUuXK+U4cpWdOJPHaD0oUgbVBSK8tXKiNewKQ+LDka7vk8NWW71AC
D6nUO7nPNFYTqAK3iwfEk2wNVZSQXb1lc6L9ZLgYaU1RW/liD8Ac+Fm681Yz/S5cafZ06bgTg20v
TeN2gjR/vcTtSJ6BMk+4wCg2/KcQuWLa8R41D9J7ok2dq0emKdfbtEvnXwkL4/nMpO+7kyuQa+xn
yJhBp0LcpNK012v3yKaNwDT9bLEPtCDJjObWVUucZ2FK7OacKkKNrs5ykDkSqUUQYRcZYLc7fwSk
GUGa944qyG0QGX3BLg0cEQVrFN0J/NMtjop6SojHbc6zIA3I1Xoq5w3OTJ2OPXWeVcMwb5qeACmn
D5Vh4rsx/bvppmLeefRFGCXCtdFM9GBnuOjA+Ob+2dGc1+zNo+MrQEwbs6OW5wERvGEyQa+CUvoG
AhNhNItUH2Lm7xVJDzBEVXzpiSOqbJne7m8JvomzFtCxM3f2OWC5blfc3dIfcaD/D6LCnorq4ZWm
WBQhwOkN1NHIYGEQOUw/9yxY49GmEzCFToJj9zvAtOZCV2xqX87t0WUYGfViTZSStT25dAfEb0R5
9I8Ix0zOyidTSBPD2CQOOIYueLutoGLzDBYnP4VvNMCjUbktIGDz+8+12QHrt8yGGThcSDIOBmzr
aXN026R/pCEQJvbq33sqM8yQftUi48G/mH4H0Xe+AvAbbHx5XzM+2AQZOUwLoloWDNgwsj2xFd0C
0GVUFVxGqDufPC1oycc+Sk63NXb/ardh4GR4z/I63foYj0ts2otJgNFWu8mDaMzixlz0h5bFOs2c
5zWJSIuQZi5bpo+pe12FwS7/0PHBArhLrSqyndf8KrgqnnUBoubY2VO+cZcqB8iYtm1gqxnNa2w7
kMdt5Esy/Xaj57IhJCRbrmqWI7eqBL8otEHXQTpGjXhLtIhVeGQLW+0MzgZHo8b8xPZL1EuSBF45
EvvcQ1wHMwYQ+YNY21Q9vjo5Of0uvlI9476we92/LFAB8gUyyh0hNjDwEyas9xQHmMGKIk03IJCj
Pgfjzem5C7z7hosLEcAIaA4miHKIoauuTMpvqclTBKU9wGL5jouFPmmKWHjgbdLqToz3l0ikGBu/
azPKv3q8UkUpqIPM7WainATNV63vhEm2T4eudL9b2/zLpK5/QgQinsDkQ67XRagcbL/fcCqZTInC
7QCO9NNRsaRldPAsH7llhI9MsQEF2rEof9XeOJrQ9uIHTIjvN798oxKrqhIjMl8sBTSRbQmMKHET
pK+DSYVxHtLSaYt9s9flPK2ucCO8sz5coK4iSkMgY+MGNTe6JFn/T8xyuwG0jKEYfBYPZlupirEx
sT2IAWRBQglM//Qu8eTbijrk91AC7mo/Fmf3F4NjEmnlY5GRmm6Ep9Ivyx0ACdQJ0dFKdKE8GCHg
RVh6dAs5cvAhuClKo9Da+tA1TK6vCu/n6Db4Eg7u/QG3/04iYhtY+VZI6umguARBHaCU6OO7x0Ab
GUKe+mpZx5+kuyve8p6u4GWLymz+nT1vucWNsOoVP8VnVZXnP8TreDZgRsRP3SL8ZNWfp6HXmooh
J3qW0Vg4UbSIRMtYYrRqhob7sA8mtv/HE5TJ1j9AeAXm0AxQi9q7obSI9YZIiajNaN1CrYGO8v1Z
MvpQdZgdc+H9oJ3hE+h914sPubs88lHMJv7qYf5K52mCirfudhHIMRXyB1xusOZsv7FWSAFi0j5u
0TswWM9chlKxXq83aweXXmzCe6OKQdPLzt0gm+AWfRxe1NGywTnWPvS03ArWUOaksaiDSeXFFvrW
g0U21aazVl5PNtP2KEsA7HA6kxPar2GI95kNEw15Di23B4xWrzW+ND5zUaoHuJlOO1xI4wrGJQ0K
AjQXrXp8OOPWKXC8mhR4AZYz8TlqocvIbKqMS183m9qRNqDaVRtO2jFo+IwV1evP3hP+ZDOLvwOQ
OQLVrw+Ei/Mqaq3R3vD7aJRp/1FvRlA2RFGWZRnHS0TmlmySW0BoZOS3MZuUe7SWwqQxdXslCO2X
aYK26lwDVOkS4V3MtzM72kAhFc4XIREbhTuaE4Te0vcL1YgXLg1taAG4FkZ36og5MzJqHPhx5+/j
jP3CWnV2JoQ+3MdlpauGT70r77uqCFYEls78d7KqCeVYrjsKGVsYl7d6ahyqGburo4KUxe2xhmdI
hru68mVKXif4lqjlN8PxPCcx+VPdvc7+lUjyDyDwNYTo9oKvjzEv2Ow5i2BNLBmV18Wif8O4OZGX
cPUb4573seVLsSEevU/lImbmZxtiMx0TbnOBOGbfKsv4KfyizzMJmlMcju/VmypXlgMmY2iKW/AA
T0DyCuO+F3ri0HvbVqRVbKyqCcw/mTRA782V2fUl5s7siP81N2gLjf8rxyzHVhIowbfs6+yCpNnU
NlBV4oO9E1/AKzZDCsDwsAhUj5HcNilJqcAEFvYkPPHf4BG4Jp/2xR7/woRPhutC9+6Go/5oXqyN
C8gZCKm4Y6w6crdVOM3pqAqVAqaak6OSdrJAycXtm9z8w1rkhXR15n5s9zN/w7PTJslABU7uJWPC
NZhQc5zDG6xAIgD75ti4N6of/CLCV9w5YzuRcUya9aYmCvatnJQkSvZjZFI0bNh0Ye69DMepTjVw
ILMD3K+hOYVIwKBt0IXb63T8q4QV01uvEbZfBRtnOgs4XX1vrbHVr+MXpSrU9Qz059IafsV29WBX
M3/jidtjgV0EHrV4I48FDFFIMNULMtBkFeA6Yue3w4ZJ4lFob7+evZBO07oHFmzJJJU/kKVWHfzv
yzBq90LwZEMXR7I/BdmGrsGSxgf63q4R1JSD3kcD3lfZrk1fU8U0k6wpXGPrwHPOp70VFcM6dlGq
yOKPhyqD2YSSLuugCu+5tXm6mEA2zpQw8DfY3NUPZIknZ/JOtTl8n+jwhJmIk58A3iGFpV7AmOpm
54dbR6eqBg/BJ1IhhjO071BeET1aS2IFP0BBYvX1awniBhAxtOR9zOKS7SJSkQh9dJ6jmgJjj6bX
4Z8Mv2YRtk/huKYMZERB/G2n51dcZPEcGvNdC36glD8m28Afu4M88rGp1fpyP+LxRCBm8f/pQFqT
fpPu+EQ5PVKiEVuVvUm1YM6irAeEyERe/SLIiu3GiBmPn67tVDTAY5uo/bQqjHgJZ4VsJUudof6b
lR09o0FU6G0SUtDs6cGs893M6QVuODrvfiQ7TjmRzh+G78aS0uMJpdKwf1Dh41MLYP3iljBJ/WEF
eZzOc/vyvrMwgfQeo2+C0EaVMQmX2g4aAXtTa0ufG17M0gZ6CAyDyY2pmd20PdpPHiKteRh/fEVu
LRf3p0fiQ6UjivNQlEskUim+Jc2+aE5NMnZdYuOl1Zw4F7toXE9uOvrPnONYJ0+AwDBwyqMiec7I
eUm0VJN0+GYMgE6DD17c2tPItyfh4PqqyNS+AU9UIG1TZhiE3J4tzSLvS7OCg53i/v2iF65DiB4h
GCeBHCIQbT9If9DgkQCKpvf0N32ztgK7oRcAQ0R5Habz312c+8uUMQo01J0OoTxER+FtwB4wrd9m
/7TL+Ovu6zOIT+jiFjSvdKb4znCuXbfWrOeMY0tn0JdWW7exK7Gp/UFxig19VDubPYqnYzxorI/l
jxk/wFP26KeifLzq4PXQBEYC1A9YhnLatv3JjxExw3urG6SBDq3/b6qy50lBsfRZXMkKi3Rt4YWU
aAEMmHekJnVTQEYwkMQxeMuM/pcgslvXy8Ej9yO1vnyK6DWz9hNWF6ZVDiBr72IyRc3qxJYFB10z
udyVwahhio+FWj2/P6PlVDtD5NsFJMMR6ppXhnKt67PVLxAi8YYSJBvnNDNSQoYi1p9b1yfcYLWF
dmfrFxI74Zr+YvOH1ZlKZ/Pv2+bAoNIfM5senViXnzIrdH/Y1P8Y3ptrLHqAEwgl4IGdthdq7SgT
C8UEHSwt/MTSdW5DoMK54yLWZ9EgcjM/AeToZAs/udUx9QT/ZFqLupCYjJ2dpn2TZ/AocAx+Wqy6
KYqXumjifk6L0aJhSHaNxe3IOB8YnyfMUovWXOCgRLHqBIcFec4O46+2bd2jSkjDRTp4tcPc21/U
keDxWrHViNZ3t62orXYgmRYpNT5vzW5HIhPz4Zw2+RTIrGgCTA4rmtL2cd0XhiQgEbt80tLQ/Af4
ftB87fGavB8LmGXQZuNUOAVkP69FoR3sSzzX0nNmZq3uNUUZm4lnSNbaoP2O3inZAnR8XtpFJwxd
pT70rMMXBAvEcmp7X4ZJn2NyHk9HiVzd2RjAjTnpupuClazniyUXn7P25p2L7+OW65mcWKW5TC/4
IPKJedPskV86jk1F+nEJAuENXkL+h7QMrndFMwizGlaWi/5I102HrkwE78B32UQqGp1xCbD9grnX
9V+c6e+NJpSV4gCIp8/KpO4RaJbM/Kxoi8mHl9aJ5dToDKoHjomygICBtc6Q9KwQ+s5nBU5TsZfC
FxrhKiC0plB5girMNPfxcN7ZjmIoPuWQnQCkrz6d65yhgHrZvRczZYNqov+NemX1UnCEus09egWd
kh70AbrzXiSIfXwIDPvpFdr84krYhFeghwuSJ1n+ReUKGe9/Opy6hUkLq4XnaNnbYuwluhkaiVZt
iokVGzm9OKzqTUIuQ73XVhz5rIaAUuK/prI+W7xXa9k2bbU8CuQtA1sKj5sGUFpfLfwWfd9PTik1
x+kSDAYNVCqaWePtc4zEsi9tVaAOPN1+xMQQj5ukq8Mh4CNz/I7wU2rrZyktddBqxa8OgEq+XnT8
0jKGOzUIsBQxCCN8YoNynoNwuMtMYWDPohuK5PC/vkcWU5u/6q812keVYsVgRaANrOrLK4KvX0Un
cB1KcmYeyCgb5fpm7D1b4DXG3bmb7p93NuXNf4KSucXcPc89w6wjpD5RAUCxX8H0NLv7xolikXiK
35QGVEaU17h0lR6ujUKT9IF8wg/uYVPDKYYCK71XP8pFV4qUaK40FMnZ8qxQLpy4uOq3RtMXX/xm
f4dfc2W7O8wLVXTyiqzlb0/Z6DSoQKGcbaaG23sOPbaxVNZCOHd9rEbrmZgk+hZp9gYM9eP6GuIh
YWBvDe16DdHKlD7z+SU+IjEQgXoPa46HZ26Rg68Ct62k/QBtlSqz4Z5wEEDlnDQI7ABSdHmaQYHU
5yWvjloKYxpr/cUFqTAzVutupXFG0AIBBVPO+3zkKphrp53TNMYeHsSSK/0EdFScRRg52oGvWskH
UseDyVM6Knr7VYJxtIrfXMxfByWtmKuBPVg8wxbJjPHoxSyHbxycBxlr5Ss3JGiiCO8TedOzY7vR
gVvknh0MhuVFOgxMZfuBKnwoAs6MOwmJBJA3lhLJREBy10fXBy3FaGRSQpIFxTcbZ3OXJ4AT+1Xf
qFkx7C6IFyE744Wy1bE+lAOpZMFyJUg0Ses9cl4Zdxou2KnguzjdAL2aPJaI7w9x0G8FR6Az7JlJ
GZ9u+efwpIrWLVnMz4Oa4Mdpt+2q2Hks3cR9NkP2nMo6eEzCDgK4PBCRghgjANJkGk6Tt3CWho2c
fXYypDiiTG5KLuMcceBS7v4xEy6sdDLsLcU/McC4dFZl736K+JaryhAStkDWDoIMqQ0iZsOarn1V
Yu/ONXdgCC0LGN9sKEotKSMyRfX6ORUFS8No2TJ8V6bTNkJuvxWcYN0hER8Iu8YroiRC0QzJVTVq
1KyHGbnxsjkf5fr85YnBV2TTs3kduM53AvIAP3zNqA86VaFAtz8XLyoFaiKm+bcM6HGvEqWb0kbL
09B2M1jIZ2oz0gVdt2YzW229eaEx0SUdGGnPgk4JnHBmqjeeJGeXeYhLuEAbaGJDQ1ETMFRLxrd1
rXXCVmsZOoZfz6td4vPBUGSyRMPJKxnhHH5a6XN7el5lMtWI4945JDMdCxJQQb5R9ji5CmKZ963n
3vQ/H5atosqjEkOGWWLECtDIWvjMymqwReBJiNBTOJxyMYKT1UCgnG4tX+uFqBm0EF7Qa4dIz+KX
cwwSaSdKPnG+8nC2mH3j6vC1LVt3UyYqUYyN8iuJ7agi+DfTDSYT8NfOpgcJrnmiDME8cQh1+aXF
6cwXDUtfhOE0OFoWbUU9YAyxQlpuEb6DwQO9aNuQQrrqFqWNw6p0LDMhQm3lJ3lIKMWnvWeDYCWi
xD5eYxQ8zYbGlLf1CxCGBbUpSaoqO1nP8pBZPuwcGzsNFwej6L53hqV+iHydm2jO3CoMo7jLU5R3
YiHvIG+wQp4xg6pjKunDhNOJWIy/yoqZYls2DmRjrHWBU67w+htilsLorDw6CSKUM8HYtZjJs5eD
NIo08wTx3M1w0LFfeJfkTOasC9UfNSO2yfOk5l0oIGHvO3j26lSHraghDLehuLsLc9CAEB34xCng
sLtWoAObY3DfsYSnc2y1kJppeEcEMUonn5VhYG9ay7jQ0SuS1gOsGsIbNXD0VpMRMNYNQ8HuxYSF
4Wlt4oUK58v81cUqV+u0p6+VCBwmDFjy6BcvS8OJ9gAHjCqkk8lUEpdl7QL31gC89ONmIxRjoWN1
JUFVz73xPFXMx5bhOyjnY1puytYDztVRs8Q/Fic/nSfS8XLlgdI5azX/x9XI8ivoUSinWWAdOk8t
ZgpnEUY5MNfyPrUzmQfFCDyqPa/E+5TjSDcH0W8xwFkDLxUvPYnrQz8yRenTkzIgTqfTrv4TAviJ
JmNh9cow52e/PdtBbtQnEP0yXLsIybmqXvGl7XgtT3foa9mIBhW/N1HEbmA/ENsBej5V7tViUdCI
OXREyJJCJepaSYSif4XaBNUVFmEfJE5wMDlZBme8RCeIv4J/EoZPlpgw8S11d0WskFMYr5TmuxT2
bZbk5FBvfcuxBPkQcQfpl5Y22lg1RGUl+uthxz55cWRMx5NtlTpdrbO2ViDQRUazb4chAD0naKVb
42rGCFmoG3GVMnpkjTUUJRUVBsIWU4TUHDTm0xqk2QMMZgi2APDMXoOvLWfZ+hEE6YO+EVaUvpFq
tI+ZQh4YAjFR8alvjlXbq69nCYSGQSoa54e9/a+b6Chh9ZZHnAodeBtKnqDOlTa/w+1P/gq1UA/H
SDAZOUV/xvY/K5CFRH1nEBsOcl1dG55MFS2Efg0glDIUBjk7kj3ufNE/d6eh40GR7lFLQaM1+NP9
7yJuc9Im24+sQS6qUV+yGB6uvSD9Lm33Bp/1hfjWDIYPAjbeHLpPNdylena8+r95RcxNYTx0WrVW
232cNQMc+Lk5qXagw+HTAHIYFHB5c/GFWtGP4Y/cjL87mtn0rt6zNiwmD0KpHuTqEjpKfYV9228z
JiLdQvv7DYapl1ywG0/G5cHaFa3KE55KjDU04taVfNfArzgi0zOgakCqaNi1tEayQujXVzNqB4nW
ClhA41FOH/NFALd8yfCMXfxbuDrFVI7zeqzDfyJpsu1ku5gTQ39YpYk6ZbxsWuT99RT2A3eoRFSk
VSvKSOVLUqqUAN9jykTf/9WrHQeAZbH7zGzBO+gTLDzSp282FyPwJM9NEMPOaS+sfJzxbtZbzE7D
U91DbP9yIFaIxjHUKgDi8MdtxleES2hyuNAzfonGd27V9il4rrbAjYIsj+zDMdLWdf8v4LyQB0Xo
nQo3KnSfMwAChabbcc8e8PuECN92EmLTuYWatoByljJeCI9AJ7zM2r7lQF0bcI433tZ7B7LBVXCV
x6+yGRR8chTRGEioh/mBJdT9u+ky7zJNxPMZLFa6eNHTSyq7LPc7qOodET5aIyHacAc9DgLa0tGt
XpWOFp8K2XzC5IWr4VhYwL6UIQI6tcuIFN0IBJighDkC7TOtmbYQsheN61UfdHPJ84WrsvGyzRqz
anhBGU2hIx+4d2AZHM+6zqaPrgZkVm7B2DYyoxdfHumz4f1xwDUyD5SBfHH0bXLOk9JSKOJoq+ka
zrRmJ3I7ZOXdmOvi5PU8cEViLmzh5sRuCcF6vq0i+8FX8pScRhleczBxMSOccROK3o+rZO4vCYhe
iD3kcxs80oBeobAM+TyepYyVY2FGnm44gSQ+YeV9ZZpIyypXa5lGzFq/o1/mIxfB9jWEo9dS5DD4
rWrWABQb3oXsMBprMXJ8iV/ylsevmrDIQE9DHInVTQrCKeXEUMc8lAA5xYcBLZQFsjeHELczVlk5
fEH7/WQzRSSpet+HipiGAxfCGd6pG7YXVUEWZiGdBMMrOTmJKhrVqNs+8i3NjyCqoKRNcXd1w/oA
w8zJ52APUhFOAFeTv4mhcmZ1AZqWNh9d2NYaoRK5/csvo8tQr4tOQqQ38/Wj9EpIjDIoukZlyBpM
XS752anxkDYEE9bTP7DjzqYQiXTT03qhn5CYJ6iCLBLZe0VuMxOIxvrBdm+LDs/Wa5+qEAeITeZR
9aRY/HDsv1nNdzmyBoLuMgInhi979rwcEqTFMOH1ZEdpuhBeETzjQ7RreZAld6hB0n0eZvqLkE+S
Dv5MW4RpUxtt2nxpladb7517ilvd6fNbI1NTnelkRuJhgoA4acbn+xVvmpSwU9GR5GGRjLFqrf+I
Apldt5JZCzuYIJfnIBdxAivq/sIEXXxDjxSJTiEQUrSgUjkV4nFKG5aU9RkJMFKOxT9pqz35qd3t
yBDI7vxD9j165X7HeVN0PXyU16cfcfMs911HqUSOBjVFeqEgv9vzaYhEimCbb9OZvNv1xIapAyMu
AfnQ152/wF7n8S/5u4RwKFM56J5hov3nCzCi8Dxyp0Tmf+HNPzvV9IBO8/dofMS0sKhN8ix1BNBH
A0Vk+JvksOnMaAimKl2PROcuwRD87imDZyTDtDH8I8Z0OMHDPlOz0ci401cnlf2zFR0yiAVH/MuB
snqXF6f5Djs1iLqyy0WVX3ffZGCk4MgFSxxn0ULjnG2CYrSpcTyLr9BuWDGqyzBoT28wWrUZUMYQ
9mkY/5bZcC1D2DrmRtqirmSKqte9qz3Wl/OF3VJkdbm4SWnKrKl4xNqjKLMSv3t4nZLOvxRsej5V
j4tBsVh8vuz0tYZq+HSq0YA1J+ObKD8N6kp3E9O5I6uMWTfDmC8KeXwNbIFOSCiG0Mvl7r7lE/UY
KHsNwxKMjbpgzA7dbw0XRMDWOd6zFLps3ivXQbLSR5pv2FeZDqgB4GN9I+HgoS4zO2hWaM7ldyBj
AzBYzL5jUps41IW2dewjGVDwnJxombvt4/eNLr2ufYNt+/cQb8HyZb7ucZTauRLVSTG5uW2x7wJP
jWhoE82WJwelPRPs3Ohn36cnwWCzwdG1woKI30sf9smUV0oX1u/3AlAxV7cZH7CqaMCj15IOLZJX
/nuVfYNgm7VBFbSGPw/kT/I4xv6buEJxOv9OAj6mXxYkUO9VcMswf0U6cuuuMCPVl0+XQTGkNTZc
UEO/02QJCoEwzJA4W3ZmHIV+HqKC5OqgyPo75r7C/lS4u+3jXRQSnL285JQ2dkQgOG2lzCahJj05
gcz6lfgfacJvN1zitn+nwntCHc0RFYugU9u9nF3FdbI/4+iOh+z02t+9rAlo8FUFai8WFYApy/qW
QS665mcudWCKCVJbKxusvb2+Dw6eMIYmuZEQr+OGqzSUzv0ZwMV2kBjZCuXxD48ee6g744TCwe8m
IQpl5JYIzk2SXYZxl0GKYaiZf/tbnH28IHAQErRIB/++IXT53EsMv2qsBMJONUh/uvBwjoV0LDGO
XwaoOAHffwqUc1fjyaSYrdJ2r25V0o/vBDpilyXiXZ1JSxgb79azTQv4GwqsCofq+QZ9DMzdEF8G
myg9CKOboJVoseErehMhyEMPa8EeKRWwCmgyn2WTYi/rWGXmNXNr5tHjtBA3wELOg1+UaIsgeos5
sikbXxODGNA7z+F1IbG4PJeYsBNvHphTtOF1Ix0UC1l4eV8e3pNnt8eA2BzEVTmNyGK2LvZJ1BU5
PUxyCdn1Ui3jkfYF67sjYTqevkasyjzEZGHjt8uw4+FHQtN2nMAbZRjY3QOMZq0mf7UPxa0f6zbH
xzroLSGGRNqZuDhcJQOJ1iwd68x6GnxlmgFGZAuluDVDtdj2h0DjvO7fNEGUfGi84D9Tf9tXVLAC
GIsHhy5YItUUXE1uJBBTimxhoJzyqVoOFyz9m8bS46RHSWtr2zCcJFCmSUmWvkCGJUALSazJYvbd
CnMNi0q7B9XZa08bWSh2U9b9N48qyRVDe2Uak+qXDjn23gKPbyJ461BEUnFXJZ+uSZFpjV99yAHZ
StQTeMZSkA3h3K5ZIM6qJs3kjVuD3vb3XfOlrOTp9likBpYq6+7BMk7YbgRsTx5OL+GHI+Vn2H6T
HPupXaehbv6Y9KgkzYAgCWPLfAYpSyBslk1xEjpI2RlfxpMr3XOK551Ltf/RQtV+SX3uhcYBL02P
FDFofIwPsAAyegTbI518Qe6lUO9CA90BTIYx8ffEkqVDg4Yia6WHkyEzTrlvAzFUhkaRWZ77TY2W
HQSKAFb/pIuIU5Chj7ivCxzN8jv+CXBNYXnaIkJEyEGy5rs2yyUnlW2T3JcnRTn5agGIHWKzd1zR
7p9wMajFtdo3WROXYlTZLGHKSTHNBAiI5Z2ynOAWs0rZQDNdoVL1gdwUztg9OHlzYaHsJ1X5o7fB
5LR7vipSi6X57IVzfzutLd++ApqVw7/FfNSeLMiiYw4rUdAy2BNUMMMPQ4UhesJifF3O+/I/YO4k
l8G6UX5wxAJQwJqJ/wMBPubcUjI3OE+87C1IBNO3eyWdw13QEl1DUAKejOiEGv87VRGzq+0XeQHv
ZafDxtbnqVqKztz3n/D0ItDqs1jX9pt/PyM0fYFvGjumQxfAwc+Ob/d2HN228gyKQGjHnNyLucqe
hxgA3etkGkTwSVbbskMw2igkLJ+Wan4leqQTHbVvNKDqWbyFtg4LZ7+6B5igvYyGOu/i4VkAU3MV
7BxqhZ7iDR8wmT3pNNQmd6LjtlS2l928c3AfKuKy1R3FHUJsBsdgkyzpJxyIMCjv37ZaQmIqFHZw
ZR4oco2kwexS/w/VEFye1rLP8VneMzvpgtlZCY2SgelnUlw9125HHPumbzskbi//ZbWAbpWr+dUZ
Z6YF4oDpREVu2PEvwgKR29EJN/pLV+Bsho9UDPE5cbaoYPyIyUI/syw/buN7COWZ4t6Dqy7eNMUp
5xEnmxPQZ36JrCLjhSQ2SmFZbasF7LyDvp1o2y4vxBfED6ykhELIKPZsM03LFQYBT/zS+F2ysCq9
JEf6/11/NomyT02CArBJWIA9fCQo0VK82NGKr1eZM1lR7QaIiUdTL+kudUF4bFPxTVzbE3LA28/k
Up4T5J1OqbMDSO0je8z5Lj8iClsSN9ZHSmdr2osSuThkE6CRWzmwvyAj0HmNqGtpGZGRlXRHXes8
Nz3BwePQDP3jDsBlPsd6yqUFn8l4CLP44M8YF2glIT0ix8tQ9x7FTH+L9Kx6jFM6pmt9c0oUymzu
cWTj7oPF0JuiXG5LQ3fGb54tPXul2pJDh/8z4meRMI12FwoN/J5kGckYQDOnCUfpZJ1b9/EBFIHz
DfNpmmzqvLbsBYT0pUmTy+ZuNCPB3BQsaHAvuTLlMkN6XLt9Q+Tza8RQoZ8a6W2OF9a8cUah6Y7A
r8tFYRacJ9f3hUzyBZClC9uCdeOVtZdt8yzn7IJMXvozP1WFxQ21hfpzosMUBiqkSGgQC0VEpIzb
FBHSfwy9KaNy5o8uqQBtiKlujZNmZQ8Br4amfemahNHVp7sT1p0iBQ9p8XbLoDPSQhnXgc4Cts6w
upmzClvXpA9UDm/vQ6GzQc+Fn5VBJw4k6G/DkWQw5GQKLkVnAX1BM7iT2mqNG8DM2TBVJ4JQX51a
IhB0v/VNERxjT3CT+vhfSC+/DDH/YtXjVFjqbtkVqtH0Eilg1gcqAz+jJl/52qK8ogz7rheOmXNE
uHdNH93dUlMLOk5iJsjGDZmzpMLDjI8S+wnBGb//jSztdQH9gCgxYbJCCu5LT052gc/xHnyMrmem
hjI5i8tU78n+oGPcF6rE/xCxn/0qf5HkLeaN/271NONNK1cZCDUV9hVbjdYS6Mdcqf8fRyRIeH/O
w6gX/ZKlQj5aiEIcxQt6z5v7O9mp6risAipCsHqZ00wHkdZzka6TtJgt6fF5+AQSGB/9s5BIsH7w
doxbRbVvNYIFv/y+Sv6KY3fvntNNIa/SHFdIpowKrQl4+eEtoA94x4wdyLnDVqkIdaO+SoMqQc4k
70nIRFDFG9jNWa5GoT8xFKVCsfLPzJvR232Wijbr6sDs1cix2eF4Cl9m0SAh7MNFF7W06kMtSSZK
9pFnudFRTba9w+3MANAhXF0q4ALdWsRx5NBjuYwK+IjRnKwqK8j2rfAxfrrMF+Ki3e70g1BFviAN
Lh1eI6d32200lho5Yvn0LqFSM+YO102l+0+aWI5f5P8yS8HXXd+rn8uog267Od5D9UmdezWgfAih
9sCh7/pK53z0sSCoykRn+GYAwEqlBqrhc/BdjspkQo2M1LOv2E6+WYgQTvH8IJWWqzS+O91u8xWt
qVCoEKVL/0Z23a8emlGyPxJyNVWbfMW7KJSBV/fsA3K30DEslE2YobJb1cW8cI7KDL51PvM5+8/c
+azrNWcgQExQsV++DScAAw4CfT5VcfS3GSSN/UN3zWVJU0S0luXeutMVFtlrk3FUdT45TU2DXTlE
Ap13qRjg+pWSlSmhyNtDFNiD2g4iRpNsULEw+zi2FZdSUJTnELb8f3xr3arYC5XRZZ6DeQ0yuEkE
sAcFwTr4GSdN/gDMImrqDd3YO7ZolxkmRPHjp7t38Mtk7fHVUWzJuuBUa/pfgswV0AqOQ6fOa7V+
rTLhPPAqAljdbuYAUwea4N3+MiU3B4Ml+nLuhi4L+EeAQ6nOGn0mJwKwSyJgZCOhUzffzKdddA7K
QFIZ1wFbnf/b0oRAP7Cv+NE5wwXgajsphRlyg329Rdg52ZyPw74+SDUDVaX2kE6TahDOIoLEt7aK
LxZL/qTueFMCj8PUTlWmefTQayJ3lWUZ2RVVy7m+itaMBdKnIX+ieSYbFTf3B6ZgG3+SxZEKPY6o
edKD8nK+vtaGbOhjvuqrm6vWq77OEmGFxecHHkn0DXMiFm4A3yp08MEtnGRFOnL3L2L+JgEOcw5T
i30jPxMTriwf5xvruxT6kele3P7/GUhio0wha+rCXD7n22NIu0qK/j/nfr9zM5t8zjwS84445f4U
18RsZZ9zWp3G357LwFGXr0JE38IOuXvcZ9MTBsNhONeK3EzenMqWR8/B9/0aeXwdQFOIQT2F44pn
/rVxZdpu6vYwqbRtoNkhgiUYdQgMZZ71SZjHYBv6NVw9Zsz/aRFhb+x6KYZs7H4KaAncg8DyaDPy
rySXujKI+cSvpZudwgj00DISug49S5f7STj1aFOPYMvebI6/TB7DgnYcdJsYu6U9f2y5krB6TttC
WqQ1SgBKWA3+fVmwJNrmlCgEqTVIh1OaVdEbdaYdQTFqv7frvLRsbqPsNczZk+7hU26wn7KXgn+z
TG9tjlYPi3jjzBxQzKjltOBIquaGVTjDHcGcQ9z7y6zmJaWb+uXzcrjgeSEv9n8ZcSdOIj5+X+a7
EsXIHNVmRZlfrIPO1bbURcAFw5molbCduqkH28K6e5xlwzTwgs+ZzXLXCslvLAyaYxWIT3UCRKtN
gH2wLz11b8VAoJ4zOMQAnV6Ft5E885FpoxFcMpDrTa66Yq4Hr5y4G9pFCXl4NKNY8bTlN+L+AJYg
pzZvb3kz90nYebH1knJrpN4jL6P12TJfxceS74FbutkA/scnfikHEiHRtb4TOjmnUNVgvbobMsnM
aVqnxpYl/SQOHvaafwxjsWSOeqU68XftisAmMGxEwRPLpW1q4uqYCNxWvJu/iJWSamF6Bpc4pOh+
MPn5BtqfCjUnoRxEAwL3YmdTdLUW2+66MF1v2rpu9tI2m+yerdu7Y1D5xl74hJRKfPjVYKVd+bc/
baApFB1AvXBSpLfY1ymGkmAy2rMlFUOs12GNlgRrQBiUX0a4elt4w3RfdJyuFFS/Rvs6cWEBwF5z
1dQUiwuEXZ5+oBKRm2+1SmdKFCcULiV1TqsMzi2FtQIhIsThgKeyBtWHetQvCamf9czNm79JQvk5
Dt52ppIMA0tLY7BRslAunTrAU0mmEIp/K7ASihxK5e1BUTmB5gLB3UNJGedQCye4rT8me7u2u+sE
NWizMTW6AyEW+9WUuCbv0ovJrgERWsA+0vb8gRhK6aZgAqYSHH/nz45gkREonpGbP5WvvfE7eYNH
5vhJErHy8up1YDb4EEKRe1c4mCdHkY1osZPCMvotpo52Q6S9WikD82fyRNBfj+JQxod1iUZIMHFQ
iQkHq5empBo+okCANIxFoVci/3drKuuEsLRtC1ruGcHxcIB3BQWsg+FWZWUyOKl8101dSbG90a9U
15I1rNlag3TApsm9F5JwvbbJQJNTPk8HP9xW2hql8pFhBMti9Wtm8EJNVasMba5yjiSLNbFcK9Sh
fULHzJEv8TIuahgZbFPWY7isPJZDxFQrz0S09TLinJTWRgXRffeguq7OmwW8xM84zppdmwpHM9KZ
QgtrdNN+GrcUgKEfYnJ7QlsGAA+rkG/uNIfbFSq7ZNU6HLiBAh6+Wed4RM9ZzPAbgPgQ4bhUtOXz
rPbMeH/VZpxYPzRzqII7ng4PDWVFUsxl0ob/L0KiWtbPjVhVM8tFPKjmPY8hFVBzUCHdyX1H00xr
ifHQLepMWTitM6ALAXbJR+K/K3PdGmj5Shv9/gvi1YFEiY7T2ZWCHiHaCjjUWiBp1/Cv5pPru+zY
mxOoK6Ya4t/hrpy1oG5mDxuI5puaX+8Aq7DIAIztMLjbIvE+2ltbtFLuHfvgHId5PleqS7NXgN/O
l10wk64qDFL2FzVruw89mPkvSR85vkRhdA6WVj0dYF9o1EK8k15J4lx7vF8ilW8w5Qd1W7aqegoH
CF/wlDVyNdQsQj4CSW1CjuqY2bMUYwh0kiF/atfpSFVK5yKkg+D5Y4e7RjTlCbZLh5IgglaP+TcF
YWZJ5IRNKslSEW+LpL/jz7NHzD+0FcdX0b2BhBhpk90o3QKEHlsqVzZXALFy5JnA+DUwix957UDB
3zNPilYyTsCxGb5mYt62Zf+4hEkD8NHSqDuEq+0SR7r5aGbUfc8Si51E91kMWnDGUaLnoktNR5ZN
291v1EfazDUMsEpiMsptEpX0KnRV5/hzxaFcy7oOojamwLJKxc8nUsyZ2/vy+bLjy1XQqY0bESHE
u6F13iJFSztJMCKRBtnvzqR0NffnJxrtoVA2neBEGjPsJuMJ8/py5xV1cHHz6m37JPRmxD0Itycu
rzo1xCYGm2BepjCV9TS5k36OLCc6jcVhXCzOZWMT8ME1DIT65qXzbfHfXsZFgIqjRr4gFhky+/zx
hxvTmdUBTOrrS7U5YUvCK8ZtcMS0mN14z7Dd3MmQ+hELlccl+8DC/61XUsv+tQ1gb4KJ967qm/eg
RbTOXZuiyEgZyBNdknSsI0S132cEBVq14qwLUp2btBH41E3lXaoYn92a+EjB8mBBApssSUmu19sL
VJzALh/DtYeOYUiQB6g7ecK6USL9DuGGIQRzY59OvskkPa7B11+MjDkF6ubwTBRab2JFavTfjSwH
HfU+qzwUO00HEmCFfEwlPvR9G2rV1vQ/rSCnlz786p7VQR3YdosMfyJUepKbIAOeC///tzIvlZ/X
oPDiSBSvsNNVV0S/upDMzCnEXYM0R82tlwZfSC7kZ7Tvv8EgOa0/UXwydY1djwUDPSk+wVv4K/Ry
eUhZcRUZS2mZnTbdLyHal6SNQdvWSwQWZdHMhwCrv00JoFX1AA+Qe6ZYYR5tad09jKLJyDU8CRSr
uamrLfxGTFJGExYYKwc6260hgODyAwvuH/cbGe4QRDfm05BwiTFlvixDqpPBQxOc2ZyFvpjQtPoW
Ei6pmCd2R+Ccq9xg7zFd5m+aFDnwWuYx3XEHlCCuHUuYR3EGKUeWyI8gaxvX7mGm+zL570VNDWFw
bvARkOOBtmIdjID4r9qY3Obosw/qQ/EfvoYYuvPOli8x9lh5w3z6Pxx2Si9vcC8ulAI6ssjyOp4Q
s4JUSyJ5Anb2nrDcpMLVEQpdUymwx+oyJwXl+IyHTAUvgo45JFO+J5VaWp0BMCXJRdY4h1kPAV0m
9pGo6NWXD0NnbY3P2Nuc42I65qv8lU6YkEs7XcgqggBYCFyx76R9UBaRfuI5Cnz8unAR8pHhLe6w
tlpMf8ktgHLXjGQNLmVItMzXZ33hdTznfWO0rMItr4CUOdtFFtMqOUHaGv4iAzUNCz4orK+qK/oE
T4zCoK0vd334Hv3PDeQt9BT3+sI33kysdEdg5okY700WJ9uTH5x8Dy1ZNbK3Lx3jjcolGJhGpTAL
9G9+RB1qf7EAApEpArdxii1HEqPK2tfykscwD3kzOmko4TEz4JDHhvM3wr7stUdptU7+JnvdNqqL
086Ki8LinE3YnVNU75cEbBqsi1MfLtOCqdw685H/kB1SgzC7prTlV+/wRX0Mp2gDcg+IhDLBC2PU
oKCuF26W8NUoIvGjwsQMy9jzyB7e5DNmf2Y/f76dUCLNitwP7JveTzu+Xg6h6nlcKx4j9aRYj2nR
TdV7gyQljK9hpPMfF4W9GUTdICQc3PE3vpD2Blct4dmYTAu50tPcf7hJHiZhLjM5hcwzrhL57CeT
X3f1So6JeVFEDHT9skskjESn92UEysEK9a16IgxOGhDu0SJTWu0EriZJAPRIzQtEs9MrPe4VwLyi
IUzYiQKKpZOUrpuswwp0OEeJME+axLMnRPsY1VtynMr9YeIUAOqwL+xmFyoMuTkc1dLQ7pRaJu+i
P3ikk2XTWEw8Un7xxWU0vw+XGME6cyv/MTjqcEkw7SYGpRVuRUfylY9QyN9AH7YmKni3TTzmoZ49
EMnUzbfMGqo+pZoVvvunHRQxJ2J5YzUF+Twvt8wl7Ilv5+2puFr7FXRa1OKpwj0DdEj0j1d5Pdy6
XNcFC/ZVEebNQ5vtomE7a+dYqD7pUaq27Jzau6Qjoe0GqQzeGzvdS7ovdJfLPi8+vwsZBFZ0rOkD
Qq6tGA9T7kS2cfCDZD0kkST1JH8JGRMt8iHdL232XwL11Di7znx6AfLzX2m3MZVlBQnuR2MXyOiF
hEu+iAukTP6iCbOPfzO/KtWLZWIc8OVuSX1lclfJh+umkz1FFemRHaU91lBtkfYvrxKynH9Hofe0
daiVLwPkNpvpxuPwUWay2qJFVOwSY/+oMt0a7UImVWlnN+J5gnEEWlHnkzSHX2+bJpBQuPhgTHSF
dmE0eBt7Ip/TBx9elMWsc9n8mtGuJ9JfvigJkkhAMLur3iNnFuX17I6cDUl3q5T2HcpeEph9kvqY
KfOAqXH+42RvPEOmBmLF9v0/6aB7JEJTlJWpfXdWyvnDXbBKODn/W7/U6GXphwFuERRz6mbEtG0b
C1MIVsTSMsTHvlWIZoIBIBaF4Aa3hCX3O4CVUOXlC7SQ5B5cAWRmp0ibOv2YXO/045YdcCVyUo/s
jyjWZsI4wcKd9KU7gwopaPg/KuXL9TZLA31qhVqyHmu+BS7Hfg0VOdeB1UkBr4kY9L52QqYG2IOm
vWgifU7jpSI28g0a7G62kImnd5LGtLpTrbovS7f3CFYM+nZWj/CV++YezQmrdkWnKQA4AtFb0lQ9
pziWRT90dEEqmU8LHLJ46Sr+3u7Qz6AHbhE6Dh+OKfUp1d674nwfUZjAJCR0gec7JsiiJSk5NgBJ
nFSlmnP8oW7Tcs7oQGGkeIQLYqRu5WSUNSqXCpNET+9P8sUA25cA0KRPorw+EpDH3KfKwF084+5a
VztSxH0RvdZxWfwQidBGkoRL/FGbIbjPxIdlDS7TahcmHv2WLiGmO1QsulHqj+Ezc/kiemFinizO
l00gSlUyOD79SI26kpAOmfrlmfZd0UBEn6npfs4FU7gtO37+HNXRU8VmDOlLYxwzJzqRZbhsHYvV
Ck2pJQ3yz0aJitH0p1cNvI4CDR22gXneG7eWH6F/EPBG5oyBZr2HHHjRyMid06vXJGUe1x8wHArX
epuIHkN7JI5fxro6qKix5OKyN4IytZYlQR9RPQdo9tmjeCZfNqKIMVJsxVgYHMIG4UueK18tOFby
jVU/MOTjAyTmiYA2FtMq95jEM9bLTekBs69iazGIcBoFrMOkNa7Bmt7yYbCkrm2NuJ72jctyfeNg
j0vVU/RRFNZyTNRWNRKLqrVvVV0JSRwuoY0qBFxxz/+1PE/mZYFcyfgUyPY5igmIV8YgpLerBOTY
do9yt0bRLMQ1fHOQ0mtJVuwOX/+kmLggWkyLSYGqutkHoIEUkoMc2k9iDsvNANED4W+F2pAYKMvD
F/UuD6aJJ8KIM6URPHRAXfYVhbmGIgvI8QPhjQjOc8atzq3N2lJRuUl5W71xVxX2i0mUqJC83upY
o2HzTt9/DcSQ20Q2TIX/OamPm/8QpR+BRYO5vjEJMIFIYYL+ilqZZtb/KPP4Hbrnrq03LUAeogz+
F+OLkkO48HHkTVvhE640ThqsVqlJTkyW0oLl/JRn277187BYYi7F2AUr4KDrszZu1vEo2Zb+Yg8R
HxZTXlnnjRgiS1eZ702GgXVRBJWoQx7Y87J4aQCPfOC6OVofreexBeaSOJFrZWX/0JcfmvdMRukW
FvFys5u+gktp+aboG+zTfCwBFMUTQA6kon3nWmWSysVLATFwL2HrrLVh0LWVN0Go9VFRJg5nDkGv
S3da2i2qkyyj0+MH0w88eldxAOn2hY7XuidJ0gHULLx+2jBNV3uCgyqy3AMA2nvft2H63hLN4HLa
1WdeFBFh1I57blss2RW/XDOI4wSREMoKjLVDW3mL2iqvD4gTQBcLizIoVWaVF1pDBG17HLscllKu
R6kMSRQb+W58dhpq5ActrhKWqVlxhAEJztZEj67dbTMjFcEP+6/QwXr+2zG9B5z8DsoR4OADrLH8
yxrHwquDs8xOO42T3SwUj8dOzQXzDWkr5fd7pDnsalcmmUrPpIjXWnyqPi7hn4jgeJ6eQHJ2oEuc
J0itjaTH+kgGqE1ZASGNlPN4o5Jn0sDuX8EGTH5xYP7aX8PgFprJBjIJFGwgmlWsqFpunM0Ju770
94Yqf5MR8NUDUCceCZ/7mggI6H2fo130nkXQxAFp7TAxcPu2S2GMPEptKrRQ3nPThoLWYu0E3D+W
3dezvwVTWptmOPEGQJUciTXvPfmgFvoRLpBiMwtc+/C+4WOumiz0BQ5adGeqRGO6tiYP0Vg4d6M/
G/VyW2jTvHEki686Kfo/5Hq+v/4wqWoyiDM9bKUU2o61zWdhbwpeDGNC7sjDo+lsbS/NXWz/m47t
QxAxHoo0B9tPiPfp4RTHTbwcVI6nMVpODGmDff0mTCm7Uj0e6fvpt4up0Otu2Rew2tncaQM9LFUP
2nbYEAs4BSli0ZCmPyAPM9e8kRT3jtOiVGpUjOTZ+KUY8vDZVbIw2HjhTdWfOd711fY/VpNGytVZ
UZKO1rmzRc7sSwNg8ayPWjYIeFE3QFNcx3gaqrYgPXg9MhW0GUqyr3n0F9fw1/svnXa1Jl4CpyAm
bSL4Qx77BTw4yBJ+t6+jQCMvc+4zV+SPJsYIHZZUXQsohIZKxOc2Q+1aW60kQvjzsuBe0v619y7Z
ZJk3kaies3LXaFjFh/c5Hy5NGpwRgr+jtoDSqsWdWZ8zARm/aw2JmB2fXdeYy23uCp1zG4G60jNu
K3ywjEnmvoI4qaM0fysR8+Oz12XIK6tzIREKSV/3RtGZl1lUU/NEZXQWzpLyL3WM2UC2XeC91uHp
lRNsr4qW4j4WfqQcJwOaQJ1jTm7o2OLDlKmW8Wv/CDwW3PiWUEW6HicoEJGBi1ljaVm31qo10Gi0
ZWYNk49qF8uVRqp3qzVD4B+smaLGkArrbWeSlHp/3JnxKno0fcIjch9Hu+YoTL/pSdk0qF+4ZgtA
JWqXF0cdhtn132khIC0mFLpO1BpfNKKE8fhX8XnS8FVP4YocPe+uSL1+oII/pfB93hLekOMX7C4p
+r5TTgpSTqvL40/E7gWRcf1F3P3kJ+t1kN4TDHVhE2tW3PUvyDKvUIKxs8Ypd4c00iM/RCxWnmLR
ad27ik2gdBevluaTptj9pjNLiamEwHXC4agC9SetVOO7UzQh+V8AZDC3NOes1Lv98k6crOXPCyLx
G1fR3BcoCFdgZ0qyGNvraAywECQ/6nm7Ob/1JKX5ZNaUr3KpYCa/14yyb6WBrWr42/C7jHdB9VlG
rjIqcQ2s+1zES7wFX6Jp8xif1nCAx90F4s2OnlkejBhLhaDyjVU8sDcX6gPG8tsMJK5Jl1qfcUJn
mBIJN3+7c8oepFqDI9by1eemdNglH0PXzTMKA6le5v0VCeRp4Vqn3A4ipNrunrvIfSY3velJiO7U
+bXAWr4u0TO/8jY8homsxKMvWFvM8bj5/BSmHWQ89BJeaW4elKuk8MjP+eoHSiQnavtwgjxExWkY
NG0sP4L9Dfv3Em7U6WyO9Ytq4OL3onD/12aQksi099wzzYEnJroKZEzvo4qC5oKUjlGTd8QaL1aF
1KOy/afJzdf2rx/ZGBXMqzjVL/PBfRVg493+XmXwDs1Ozeym+gG2uDalZm5pd3NbB2ztiE0kfVyr
NPSg2d5JBr9DsN3xY5f/mzCQxMrDyEIqVyOQw4TD2x2pKM8x25qcbIY7CypcyRMBeb3hbeupYcbN
8AdGuqRuIEiVYTL8jPbYxCRMMt47m80HD+bm0ltLiQGG9Kmifo4f057uvmHfrbGIITNtIuUkKna9
qC/LD6NROIqekIlLa02Waeudd0jiX+8ifKW4TrGzNu4dynJvxOB6RSaN/2+aqeAtJ6fWRlAGrGi9
UePePG31jJtuK1rzReqBM12tI5U39xnSEaCr5fA+uD4tHtvr9cNXFQJDcSS+YUuQcn6yOoUQaq8n
WBLCDo1/fLE4OscsQ4w6MBFHjo17k/9QfstkUiXzJraXT5fUHjxEddJ0zSKoiqJ+QjaLzmqAvEbv
aY7YNktiDDn1yrpCEz11i113+FDv28dGtUHcZExBsNs6wrPGWMN4Dmv8faJa4NcHzFChW5/eGx5U
rYwgoixTMGvc7hYQ0nrR3egtVjEdlr7SLLRq9/ocJngDMCKoFzfNzW49aMtYLk2TnhKcgeoLXYiG
LOKs8HfLBFLFeeRrdT7QqjDVD/hNsRdorbLR1apaWe3EyCtO5t6WUjnBHGBZ4A1SCbju2rHaC+YE
pWcgFwCkFAjJCl04rjpTboUy7wvYWctAPXlrG/64aM6qYPjnvT81JiTCG6ysT/rhi3EZ6WctwVIU
mCf4SgzE18s9gGLzPbhEXqCoYBQy5vowaSHyZt3I1Vc5lNGTsTA3Wq+QqLHPDLot/TM7rMng5FO4
nIlwilgzARrgiVqOvPIcxKA2DwpMWXcJrc3mGHzk03DvNfRS9ngn5Lbhmjl3xEh0E2Cp94eDSK4W
dX19Mc6KCe5jjHqg5MJW60zBqb3Hab+CgZvIOeGoXj/wnGSQB+9G+mYMxbJSI33NIqvcNqN1Aycn
aGzFN1Nn4MuOCt+2MuJs2tq0z4iV3VcdfRqeq+tvuWhOo8YJW3Nu5Htuhvi+DkhRPXcQH9DQqMhW
d7vXi+vSR1329SvG2orjiNsJynk3a3nAG/NEVgCha+rK3NW3ht1XuwU/HFZLgNt6aaiw8mu35dkr
Ff9CdYe6jr2cqSck0FmkQ4E6eDOe5bjjTDPZhFN+YRv0a8cwEcxJqnxf06XvRYgMwrhJ6prD7b/S
kVbvt8Y8SQXaOAOHqLs2LE1E3AjVhcq+V2sgQm9MWyiYm0DP7SyhmpAJVvPcumuI802ymGPlQ/kI
ZBOwmd94P12AxeIw8dBRxTLCcJ9ZcQnV8i9zhnaOPkvrKuRldN4WPCGrUmcRWly0aO4SwObhVnqa
89wcdAYjriMuLAuBAgNnjT5INS7R/EWXMre5JV3l81wG5G9lGd0TtACsBNRCYbCKc0iTADjssUsk
9HyAbzJz5teRTUNfUGEjIxPGoIKqXBpRGSn1vCPfGUS9u39UbLIGlhz5faYLQnfqcxr7F7r6KZum
nRYP/A+lCHvepY7odBrkYtIt11JgAKlmfSA+Gm7Lu5BYDPySKUy8pXcubJ4Q9ByRTYL2yxIlOJit
iYoV5hgNOokGFJcJkGvxKd9t3voLvQIuZTJgI3xwv4Hw4ugz8m4MUM/pbFuXRU5U+S7Z+3WFyhWh
pP8ioGjHLdPN5cnd0ohSniI8psqbcbOQYUbp92FidxRlD7zkWp1DRWK2nyzRvl6ji92SkbvJVqYB
epPJYa1emYzIISHNeFukKFqn+fb8naqixWJYlR1g03AIPh1C1CEw2xEydIxOsN/D3R5c749feAwU
Jx6r88Rc4FKnpmB+sKVpCDt7O1rLQwPTqLpR8/SW4y6PBNv82R7V4CJZTnkWofBbYBirIcoOpsJ6
TigZWXA4Djj9zM/wmYRlqjklFWAfwOkVLrwPDfwNWUzkTNhS9FFwYSQGFOBH33bd76d2T6UrZV/1
XKElq0aQPT6vR8pUI/I/ttGB2aYgTF2OYoRplxUVDvTOUOH5pQyiYZjVBywaAdI4Imr3kh2RxjIV
0j24NbYyX476M8M6dPGUqNchH/QRrEdR+ifCzb4PffxavctVJvOjtrUT2JX2MvJk/SmSi1nLBOA4
NY5sI5NlUYMA/atKocXJ1AjK+yPuRVNYsThfJQb6Qi8KP66AQcSxqMpBlKfjwWN2xS4L/ZDvNtwQ
BaLU4CD06VIZCkLlC03vZreucL6JGZm4pPJRkexFjaIAEHTfE3gI83lUvKgkfeyT846et4vtBYqB
yk8a3qtHGNGrVoknmDfBjEYJ/RAH+2E1w+G0f3+PgDQCfkkz8JEnAW6HbhkYhBCS9hbnB1jk/Ei1
1PfiamHkaHyccvvcxWZCKCNLMvJMZBjjbZlIlM8qJATfQbw7gTlt9NBYeN59Mo3d7Z8pgcgU/bax
PB1MDPUDYrT5FH8rSZwy5cHKTUb+ss6YVT/Vth/VsqD9WRQqgLD2/QOGjw/wz2ChAeX4eLNVLnPp
1xYKCOFAxLTp0HMUMEqKtFnQ6YJnBSXsuuDQ+TRcz9GwKibebkHvrM6jrCSOH76+pOCIPnQzL6EG
vRqDxoQwgbbPTMxTJ+ago9c3iKIgwAS235C6xLTHsXqXlEniaNa8l77qbygRglWbe6OhTL4WIkHD
50nY4LuwPSD+6BR6MHjiNtD4oECCvRUppDaR6DJc6TC3TVVum5/c4ycKe63eIsYNWgQPGMgc2zvy
WRPAvu2JalKNFTzy311JimulXyTlGIRMLNm0gKYJt/if4HFX/nZ27XumJazqgpAn4HtPHtKUhQrr
IThMZpswqxWZPcuqtD3T3uGfI20lTokkbmvdsJ7a+FMDYhiYonLKI1VqDfjKFUDZB1Kn4XEf1faN
p0smFrBScKhxIy9jtb3dv9iU9C9EZ44Fqr+MsGoZSPRi4dCkW544eIqd+q/XfOFZELa1YttiQspH
/3u0bTQXq8eUVEvQskw0E4jvoq3hi2FNtorC9yqk6OrgwZ7GyCVhDs32Z2DKL4xYropzb8/pv7y3
cYXWSF6AeHsn9QWMgW0T8ysCG4qFKAek2mLTcJFQ8Oqq7/YCqeSqFxPnO0JAZbEObQpzvHD+xeJW
ZmhH79t9EZOa4o1sIV8OwmX/Xoqzo0vvllfLTHjaDj/4oyk1hpQt3KrLVQM4EQN53bTbfobueI0D
N72QZfFOJvQ3S1ASbjB8bbuesFsbRGxPePZtPzGssMPJF5Qbh5PDSMePtn0vNA/CQf8eTuox6nB7
DevAMbtV7WLv8pRYCxAXev1ls1JWMoPrevzySjGkf62+zT6G/Rj+cLxUjHGEvuDxtS83JzMBoZrZ
fyhxWUybMf9aD0iz7hggvyrPLTW/jXoDboKk/tdp7Hde5sps/wUwkPJICPO7cLMs6wXSHA4jeCNi
RHZUuj0cGDJa2aOjvkAMOVlajml5k6vjmnd/frIb7hKCTBnRD8BrLLgJDOl+V7ZH3KbjhIqiSnvB
iUaDvGRHh7cQW7hani2K/IOkiYbY3VO//oDIUmQIvy3cqlf5kxJueEgyOD4Fy0SOVIRK58T+bFzl
4yPQlVtwf0Yfg8NH7rsI42VpeZyFx9mzIQDZ1OwGrwIY59x6CHplvAMq9WCaoVkMw4xtFWry569T
5xaqvK2ulillIKzJgYlvNolDcNCsFrQ45jctbjX+uH56N+B1qllKNQeIAbbpEKXQqVse83QsSMy/
nIxRvSZ0LBf+2QlgjUbBUqievrazxRa98sYr8WpVbTtWTQLkt0lUMC+TojfLZpNLfVkmb2qelJ4g
3GGDFhEcrCWtQzcGFS+BHYMRxtBvS52DZEXEqIbgWDwklA4gNJgDLf4xv7lbb7X20yuPY/nbK1zO
kASztyo5Z12sC8F+URDX3Ac6QONRNZ7svw0Kzuh/61LPiapFk5uEIBzXqIcDXaha8tYeGJgHNZOl
a66bj0dQf0chDaJ7dupOeBYhgPXuh3FyAe7mt7LKRfISJzqAWq0B/aKJox5zUVXlBGDvF1k4NwLa
z5962N3vHfZ4tlI5ssaiNrMP3DmsJd6dCyq4kulXYyfEkWeamCOLjfqaYNHMoNaxj3jgrJgEZi/S
ON18ug4xPotUMxWYFrPr+M6z3eZl4z8aLq9WoOZjweWuSVw/G0OzaQlIUDSDlXga4Xwi+fejhD6g
X7UhCYrkVhzIUx52by0cZHnqQKLksoedOBpXBOv8RFAjABcT5iPM9Tz+MxQzhjIB0iA74lBO8b2Y
jscxguApdxSZKGoQIfKz1PsGsjyIHOYGY2yumtA5E0ImmhIpdqsOumswFWEZdDdat7AYp8bGrCHS
nnqtXwjZjZf9J5iFSyD7LxbT6MNDn27JEI6u7jY/P5rytvsGK3Q/bqYgcRYqnMzoMi0qVOW5Dy5Q
TqYpCeyk3Ze2Crc/onW6nzbitoUqQBQ1c894z3J0REjY1lvD4rQeOkRoeoxA0eoQc7KqEBE645Fk
nOLPFifdEP3vE+pZHAY4BZeaAmFOlsRDOPY50qVptEuHZpbDSnjBRdYhRC0xFwzMGsywwQhx5Ipk
kHpiuPv8ctNf0WA657vXe82hfoeinWINF6ei5hc56w+QFvJiyUq/OxOucgSVpahkxJX+mvcLyPMY
bwPnMJSomMyfpGNa19SBsqLAjjolTWHraewGAe3ZX8LdjKjALFcwpgMWw3jn+FsBg9IKbej1hn1+
X1CdoVc4a1NYPEuWFcr/mGoRhA/Hbk/mt7sB9Q9h0spP2xHu9XT0Y/Nz9rmWBykSsQtCDJ9arXTb
UfCT3+As2kX7hPqgG8a5fDpluunuP4QvMnLlcHs8OcqYyIIqXBBz8yphl1NOmA1oeNg/+aj32e6y
MF8L4g7i1a0WgQKc0QBfl/LfA+tIE2HDLyhmtjpZXMPNzdtCVDoHd9G5B5rNrsCnt56i9wk0Ej0m
wIEnrCgTh8utkyCghRPwv3UpyYU/MgmwEymKRRo9pLPQOuGgB+UxBzhvRdgnX6KHE8f51hNDIia+
zgbkBcALvaUDAPfx89QEoQOaTEW8wVYOjinFMnZO16xQJnnwf3pDxQ4H74K+VLVTZfrYpPoZhAh6
PZeQ83zu9NgjHq6B08P4MBVHAMnEyIrEgeSrMjGWsXnljbkPfi6hYX8b+OTESILqajYvOKKQSnAn
z33pMDi+auxGdcDMVQd3bo7qMV4ol2nibFcWot5e/tQuM85IpfAbrzJXaKkwHXq9d7YRB0VKJG7/
1U66Z4wiFLW129WHDc16oNLemPFUScXEWp9niCK74zUkw9iaXpjC1vknd+8657poSuAmQYui05QF
5EMPEOzxg/N5o37VNr6ZtcWCHwedy4E04JCZYFkKOaykSpwiCuMWUPcVSHhlOcKu6jkOelDVD1nR
t7ZbWJHIwtK1EuqJWUBzCkqPkKmbrIPRLQJqAAnr8E+9T5LNhsAMWZVJNziODRqSzCq5qGvdYLjO
zk+08YMppvktA0p3oQQw8/lu0PA4JhZJe1qGIZuigi9zc7AZQqMBsH10h8/K6KuzGDllpo3uCiNH
Utus+JScP7v4Vj3gwOlENCJC79zAIVTpj4cmCrD19yOAdTJy2sJcPW1IzZMLS9pt9DPwPEOVsQiY
c23HxfYrtTuc+XekmFgnVDHXFt2qxUL3fEwU0/0pGcY3P0437CVJwlwcKHXPDodF4c8OLrOJn8uZ
XX7tporchqfEWNXnzNPbDcitbpLDn4a3q2Oae7OORapeY1P/qkXyGTDDvoqRYiwhQm4D56z73XtT
w13FKzuC9ScpfRXmyqfxipPGxuLhQZpGK0Z6iLNLuebXjFOK4n7kd7QAqBMQa1K8Ddr5/oebHVS/
uwKag3bK4xmNEFFsX24JTJLef8H5OrtuQD7WUj/zhgTn5HrOWtDhrKbaf2x8crmsI6iOO+DgmDQC
b6B6QnVrSH2l/fr+epLUhGnJFmXK8oWgZvIYBCblWZ0d0kUV64CV8/u/ptSvcua9/w9WXM/TpEj+
2F0EIUIAnRxv/3pR4XnxLh2a3d90BjRK1gdhZOIH2soSjK6bjohVfGYyHUvnZ1x/GyOycg/aBElH
yA3USK9mq7ljJQWKZTI8c3MepEgz5OeXBnjN/Q9+1mnTialwvMEc6imUfAIaBPro1Vl9JUs7RnI0
lbTTctirdg7QXdoxAjJLDhHLBwOxAfBqEITjXTaVRdOn4OZ4K8nrhlajSWCa+WW35xEFKOJZTUPQ
158xOzJxCfRjkcpZoYhU9lR0Lojt3rPe9p1o7NTgdxUlyasrtm9ew/B0YtnesgDKZw4bylSARu8w
y4Xpus6kGF+xAXrLcY6Ay0J5H0rhNTFkITovkn+L5X+xBAfMZ33iNt2t0F2TXZ7mlo8KQeS878j/
Dpupw7MLCbsZa3Jne0F5IGjQqwTQoSH1N4lTliE1Xjo3mnjDCO+AfXMMm0H+BleWxYDD66WNlnaC
mW8l0yxaGFvwUcEPMb7PM823x8PGzxy7LIPaGNhhMQUC3WnTDm1Yx+Wu7Tgjp5BOK9doxjvF8HLH
1Bllzwm9iE2og79yypcTH+TQ4yamntPv8OWrvw6E9Yz6Yi/jjvUUiAilGoojnqsBRAN8HcJ1Jf8/
F0oZZi65zXw4ct3AnCkSS1u7OnFHYN/DrAUBApzaGX0SyigqTYRhiE1ZhiPtusnHsM86cNgcVhh6
heOQoKvdzI2J3CR+Q5BFbT97/xZyEcMF9uPrIG3ayJb/I5SgGHUO28I5G0wcuil2mN/NomLVIyks
ArFUWdKm6vR2WrFH8mvKUWXjliQ3t9ZRhWWc/LffJj51AwXQ8zj7NY7eHBg2Kk9AwNNzKWkFLHUo
i/MJGDcgQTf9I50VcSyI/KxQmOAVzCcTpYEvBOBb4vYcOtdSD+urOGoXWSweSeMvzOYgd5pMxlXI
AE3UJxBsJHJOtElloBhyClKPHKh6bvVi54ML+ZKlrvy9+QVS4NRmZ0ICCx8kbyn4IHOhAJZ7KYn6
+I05HXu6uMITbnWBVnIhttuszR0rjh6WcwzY5OIMeW18TWBqvUj/tJvkCoc0iFNZ+vryMqp6klQy
MYn6wqCk+DjP0fIRMm9HXtBsyb/+6es0ig1D9Pe3+Wie497yPKsL3p2HxgY37YLGtNs0DkVJ+HOJ
9PpdYAkO/7QJ+NUOGqMsA1i6aqbi3YAL+ugLxiC03MnWi2hhT4nFBN576colvnh6id3NuXmvEteJ
n8gwiDAQV2xxi1itYgqWVFGwXb7U+Yifdd/k5MPg+Z1vmxFd47JIk8uXLLyjMlseIREp0e6A4ssK
Xv89rCX0+BdJH1nsIk0iRlNVMm4a3AzeEKLLGm15hZNAf0+TlLZ6YNBfkyHZVm8oNFFjXwp/GA56
YFHevXamPohFimJQd2tU7Sv4sygLjAnLK4GxO0Nrnac/R5Yr1sC1VqcaIQPC64ZMs4piGChglWkC
YkdBsDHZMCfoorC5Z7CTzgmrGOvFH+a6tjtblO5yQJKAo4GdmCKCjsh9Co07Yq6j/BQpLiO/vmhy
C9tLvp6EFhbDOwViAbt/PQv3oiIGuwEkHgeKbIUtvtazzIjoD2AoBwUMuIfWFgjk8joSbcUje5cs
a4xNn4uCQzjAiz5JUqaHcZNaJxYIkIiFebnTO0wolPh/sxuWqnzy3y5AeolqqYTTgDOh8q/uhDVj
LJmqF1kAOr/sUXHPyrZFgNMTzN3oh0NxEZx0qfeoqz6LcIBzT6ERyDAqnaSLpNYFH85dZvfKMUQz
XyIfe1xA2m+xmnfH8naaHSgR0hNEAvXmJo6y9kLLaZ0apheKtxgacirrCerppJTSI8oxrMY4AbiA
1qVfSrJwIjnC8SP3bDILC9Hy9CboB1gRPCzaKmao1LjKQjaBlpfACge4i06xwB+IDGry4jIiN+ma
xUPycxidnqEzCVEVQ+Z5xMQ5CRKXw09teg5WUgjNm/eLXnWLj9ExtmYHmTRyN6SRSmTl1YbhSSa9
1VFN2Z+CCasZ72F68SJ7UZd63aRbHNB5hl9n1a95M3qymRzjcppG/peyn9kP4FhwrM1P5ZnOMfm6
eTwtWlMagciaLX/MfzyOf4kkECLofZbs68jR1JwZEZ07BFvp+ElxCLygF7VLyLbZJkK4CtGzYZpY
VIpYkEiTIsabw38drwnNrUkoB6BhSvo3sVHgCdA422VASeLaxRHoFyd689/oFztpYd5rVKU2EGi5
vOzl+jT5YHF9xjrhTUrrtRnzryaV8Bcre6q8zuJvhXCeehfLkBGQEBq2SCgfnhrf3RjvGx81uFtn
VR7CQbCrsbXhTSSLV9D6Iw/TEIyBjxaEjzxzmlr6nJo19GxMXxGrst/wTB+gSqxbheJTBGT2Nv6y
P4oXnzfRQYqknpNUDXbMjSARIyETjToYlIulzrRuZ58JK9e7DK0o53mXMoUQqU2B9qbWxK2MiY3R
gJ5fNf2EGUohxoXHoBJ7zvj9N9lSbsUxyyQ0+SMDhXvZEI3fxJcJhnLIdATWY6qebq39NcvCTkWK
VzRhoB2+nPLGsNLvFkKGlN/rYEarcu/KW0OhrSvLZoKQ7Ho2TMWx/hIDKQJcPOAQiF9YRioPqw1P
MXTwW8V71vkQgMIMHR+oOlm1sVk1J/X/ltm+Cl9hKgqqc3iT2aJ+2yGR2LRIPLdh5mEoTkbf25dc
HGt4M/5mHhR493VZnuIXKB0QefacSTuK10iDgKfdBDPhhL6THGG7UGGUdBvuY9srMKlXSJf7aXCm
BrCkDhK+yTaPi7g+sZ6/zoLhXSvGgTjTx6i4Ug43P9CsBNY3hcuVAi6Mx8EYMwc4OlT0mNYxMusD
NktSTzS91sUm3gAocnnsbOba+u9hn9y8mSqzBhw10gX8A22GuM1rtxj2L6HLyBlV6IaV2haWQZFL
7zIrWsdeMg/PyZOdte9vqL/eDq+YyPK2Ir/XOqTqACeJ83qwRTM8UUmP130R9mgDnv8qMW6GZMtE
FtaDEZrUXILPJDP9mQXPknkrLArWI0kw0c4poYJFQuS4ysn7M1KaE4YjXomza71GO1FqK0n+V4/C
FHPBcHmiWc+h/Oag2MZt8cKXPhdTGXQOKKsLAdOl6t3c1GXfom0CnZD8CElzOgVAk7xZjEH+FBEe
LEVBvfEEViwPKpvicynMOWlPqj9jSb9PCvHF3D53AtbgWU3zSNIWR7Ba45PtqwrZXZO9Mp8SJrwU
NJwOJkEfVFPwdD+8vJXThzSLprHw7CBzipeuqx7vudZIuKdoDWATlt7oNsGKatpbwca7rKsdv4K2
pfM0gj1YJIyib9weiVPoUhJdp/qglwgE2oEPYolDTLh43QXTh4sFPtObM3Uuo/eUJUd+FoGFmVrP
kXz3G/ZuGTSRwLP0GomwSpC59zBxlPRidc+AXc7HRhrKI/81HhhoZpwl+4950w1eEMToOl3ofDO3
ZcDTA3CIo6kbj7t0FA8Bpr8la6HtaRREU/9AbmvPf/f5L/aOa8hU9dtNZZZvAb1FBCA9Ls3ilUYs
SrnhpkUOBeGYF2LtzRTc57wLNcOveK6M0HkjBRHgM0V78U4bOSP45/T9RjsvRKUCzI/cODHre8zl
DQx9gPXL2MVJAMBU6gdwEIzf1CYKZ8iFJIMIGK2n+hu7v5r8EihFjOtFofdmiQfMy4iORWFv+mS2
Agz4+EuA8BEfKIFVxrazkqxM3ixmX3yi8gMSDzAg08BXpKLq0FBQmwkmaGYJJLQsxZ9ZeSLzTzw8
Tjn70ru1Uhg6Zq7eBAYj3gA5hDft9OYcLZVp2l0jv2fm/lWyC2V549qnRVS/J2xwz2Z+flf+eleN
0UFFO9qQHm1rFvHQfTD/wIywZpI5YU6XBdLJgUptW4AdfJcbQ9XKLTQgoLFy4KB47ifHLukn8ro8
RwYvdfMJ3YRd4k+O0chUeGLTds5H5oGEllr8QvDQA3Ez0Roy9Qn7x9zOuGrtzbo2J/xtuJPi/HDe
UNKC58wPCGl8CsxBh3pfALEFIe/KyfiBrOiHyFQwjakYdv7CAimnzC/rNm/lBKnaMnTOEkkoldak
zYLW44mdzgVXZOhWUWZ251WtYIitVB4pe2z3Aq1pi6dmoNlkRDHDwuaE9/1eLpsb3pzSMpiZqAIt
v0ElKhswb6itAHm/skQZ61gxFBCvjMKttrgJY/WG/DZQ02CCVV9kHq46b6zpG3TvrkYXKPJ/4ntq
T+GQju/4vAW2cD9jNaES8cqaYg4GvRXu04oZaFNHR5xdmWVNm1/DPoIkFS1ySeom1oetRiNDp8Tw
mWOkaEoXedZeZ0NyGWK0iK3cN9ltmXjVQgdwSEu1FGM/mGKlRko+YDFLWRa8JJ3ma/D0Tu27AgZD
9/0v0gxcHjFwxpPzElDUThdF6T9D/rL/MFV+5VIqNSMKRiOUJd80mxaJIsVKNPFX+qwuMJiC2grV
qDAnLF33ktD4IjElKfhSa+CrkKxR70fZyjefMkr/jeciKYlOxlULCMUD18czgtD5kmOA5wfvqlFH
WwnuS8B2m2yzcw02MdsvFTnvq81t42M4z13X7M3zOVw81O0d8iqf8bbDFq0PuHhqiork2OeW4tKy
Lj8at+6SXRBOmkuh0DpFNfHXK++l2t2RyvzFtw4RVZjIPSsGLM3Yznz0Lc7LOXjM5CzqBSRtLW7w
n5l13T6Sd9JpYirIq6E4hcKZ0iLbbt+FkVxi0iGUr3ehSNSMpCSFsMm81wgGJ0yGqkjWOmINnvcR
rPhJykfLy+hn0FbXjgrYUfmNGUY0dEavBUzogO4tSLWpbjVVyQKumzoX4xu/26Jwph/dqnpfXxmR
Kg4GaSxF/M9Hd4LrH90UhM1WKDaB7XGPce6CU9aABLwrmzsDhUWIsLcr3K8vIYva8kR9A9xO0b4y
cdLPwB6qu4OeQrRpzTD3wVEBJ6uG69TyflLCyds4WPgTtrsHT6k5N6Or9aLjyBXmiIL7nuYPutPa
R5YKgICHacQ4NylpBR27583xFouoGrUlJ3lOJFZeNlyNWgOofhYCiX+qyERFtIXxqzhHgzaP51xF
xPBSqtSn4Nf/M3LxVxwoVlyqCWXYM45D4W9GMIf11h0J0B8ZYr5zTuNZ4YXsdwdeFSjbtN+JRahC
INudUh6sDxTva3MBsPTE8F9wwcb9AsMAhKiyK4fyqn352KFqpWl1PAQHwvH8xv3DfcbylyXykZne
5YlifZAbvoB2klLe2jYjxXirEY4XqUDc7IR7GgC8scFEmMgecfCA+Ssx1wb4HZYsnuN8EWXiykrq
cYpWQGq5LrMBA4v09sj0PqEmwgt+FosI9aAFV/C8wltqjP1RLNqE8yxKxzAS+tLKIBt+GO2ZXX3n
yylVMp+qK4y3BvDlHXz4CmKbS6PBjmbyuvywo09UYXuuQC5fg4mai48EBm9Olq6HMJIFrDvIudfQ
J0EwVjvGC9Q22xTB7DUJeXR062MEmTbgTVeUM3QZnAZWmXlg6UlYZI1rd8pYi4lenRKTnVdYGNj5
Uw6aGTKPjXH4jd+uYzuTmHdolvWiPjPRlObqCaHMnJZJLP/QkUSPtwnasCRgAX+cKX9Rn8jOCQa1
cBW/yz7v9mNie3gesdTBwUn/DA2w0MDxAdc9SfQ7VCe+DRXg+LvciBJDQWhFungoG4KjMb2mwCs9
npbzht7ILDQVn0OimiAmRIPGpHlbEFrCM99LVgzaush9411XXnGLuzJTcUJ2+8kMNRUZ+j99Djfz
xxGrPmUXWgAa4zEq1PrBvjSApNng/0f8XV/ELIiYK9n7NSne45t+6Af5DNkYrd/8bI5GTZYxxtKL
9VC4bBreikZ4Od0PfXTeRk7LtMiK5yclVzjsaQkwdlQsN8VD2X3/5tfgiPzngowt7WRA4ShiZ9dR
cmLVMB3f7+nZAYeojPIot/c4fF5+4OcCUZWD5HWVVY10M/HvoRzyBIrbfadDvCeN3NfHoh8HArVN
d38hZ6SscncjbIkayJHfdLd6kZoV8FSqN4xNlBhz4KoYhNbTj/c3+ejTCbwFpb94EsxLSP/0mBBg
cJ2BMog9YunsudXa3UymarnotaIQSeqa77NcKZ/PFywyCZFtvmnobydOG8zmZKy7mzhTBZ9XAeQR
x8NAgUxHjyXLxFrpalkgvuxsawPAvtgkS464frZFfMNcjVSxkXmu7QNdleaUOba4f3Q5mQ8YEcjB
ZwVGXQVp16f9NyhIi8uoRmYHPoLRA8Mm10PZFHUUuJAQ74rLh92+icCFt7zTHOC9N1wsl6bKJqUs
ahPV4P+cccAG7Mn2kDblYMZcBJkuQYLlISUapwLAe7DXc6RaEeKyyDuVNjqidxeO+M1a1xQEPRJ3
fb7+ZivCLqQYMio+7nYVEjJoZaLH+ZeyhrgdZKWbGleXaMk6GH0ui9NzkSiwhzvKhgP/ADkxL/86
KvimL+qdK2bC6iIxNKa4MASQFkan6asH+EB6P4eAsLL5NILnbYsjqt4MiRBzxDZLvYSPkvDT0Qbd
85YDkcRPdxE19bLxE9L5we9YElfgNaCjB46QXfjG2iY8X7V5+Zfy1lf+Ab5TCAWqpjDE8Zpbq4cF
Jvc2GFia1QzpxyAdLn9mr7zmgOJh5AeIu5Vhjk1PO7NWoDBtyMdRg5CqRyWMEqKxQwU7tZ7j0olW
4E792ntg5kkbA9mDu9LqaKk7zZYaKVb+/y8oP9tiP8HCBJihEfarW2Za3KVn7ssld6cGEtqVKVUh
3G3bMvopqA4TJrJV8FwTCqNQnI6J1PUEdmu46nw1vdHWOky+BIjF/jx29DHRDNP2j8D8Er0Y0GAD
QsrVHrz+QExVT3+kIm9vExn3jG6PSqDR9NpM1GozXGaGV8PCfEex/OzmfGGlDRjdVi38SF5DZWd7
AW6vTPdMAkbB+g4LfAujKjwZGK91CYSwk6ARiJUo6sYh30uQJEulBmp+n0u4eot5BXsQE3vn/KMJ
M02ROJsCeYxiMviGFIh8fLGGiQb2sHCuYn6+ZayfW7N83mvNBR54rgp/KYFCHddrklhWP0UdTC7p
UdqTtheyjkumnvqsW7fuDfhlTaz1tlbszdZrvcU/kI1ZvxphLfovNcNl5Q6Wt/b8GBvdrEpZutzs
XPFR0p5tHjqA94YY8fJay1vNu7+HPqW5Wgtot9jB5l2QgelmJnoOe2IyVuMm1HeB7435XTrrQT07
TLLvnxaHn6pqCLPefqDewdlphtmFtZoWzbwrFihC6ZMfEDlANxJmwu38P+gmA7F+M0ErkVprfmp3
zwqc191dOd9nIFEV3MX1ISN12AT2zI7UZwdsi7q5rpTzRf/GWRx3PRERdMFeKjIeKbf8RWd1mo/P
Ovf/4UAl4Xl08AQlQg65F+XyGMo2JAUhW64zDG/YEQR050iaooo4Ae0uRezhGm4pJetjL3FR+p/h
1mtpeduzJRGg7OTPM3530xdnnKGKFxDSo1O5pOWJDbufpQJ0W58o8Tk+fJ+0Z80SJKL78oJ+YUlp
MzQRUkERywf7t00GuENqwslD4Z3EYXg+EPX/AGRFnV+3gTZmfj/ZT7P8hDNPdlsuoobT1PgmoQO9
9A9RAhwn4/LFD/kuO8BR5o48mThxTDuCoh8voAY2lkLMQ/6PbUrB0kkVSc2fjl+72qDJ3E8cn6wt
V0OXOjY+H0GZvk550wbKNrf8R8lFMyC7O0MfskievUoPL4hvtKMFQAOBKeMZ+273NVpVuiL9KDDS
9KwO2gTjuUIb6woiXT01+mkYVRlwGqhOZtiEYz0iT7lL33/Bk+BwkumEnxQR4dsUVKS4pVdJT7+r
vqPrvl428LAeUNvaWjHPt5FsgTOmL6qm+h1Phmzo8NCCUMaJCfRSp03Cou24KG7tE7767WKhregY
EpIPNCK3JcLxrntDnRqyPC5hnAuiFGaoDDlMXiUkGs0HzD9RfWQtyowsSb7VU9tgTEIbmHLKzU5e
elbA6vdg8MJcEbBHeXslzDzkYpzdtWkXEuIQ5i40ty/S4lO7/NzGeVM1/lwoEbW70DqiqJdN1WMf
LIxDXQjfEw5eM6eo5AQmYEC+s8SYhY6FrznwdZFAFq9aWkn22TOmD+1esKebv/IoOA283Y1g3bed
HNkFiVRC+70XAy8WLUTBlobEIX6lRScWp+3nZdeTBzFDi5Q8OXJI2+yhipWKo4HwKVFrJl20zKdS
QX6TVKcvZ3jdI7AQb+UQeSBxBT6f3HvLXv/QJMQq8Gn6qfjVe1X2xtGGKYA8YFvO0BFBQp6pRBFs
KL84aSPtvHXGHyfnFxEWabdQcF4iVFGbxmjTcwW0FYf/nSriQmVUvLmKsNLZ+5CEhq/YSH0mnBe/
1KqGG/EXBGnFN3xgLqP3cWpfoM4qQj5pwTOOkd2fJWepUZZwNJSQ3AeeNQfymaWnyfj3Ybt585Yd
+EiufLDyhNv3ySelIH4+WlZkzu7B+h3GbfAZkw8JbITDkFem0BVls2zK85gUFLSK3UJv0IcQmaAA
01tjmyu5fFxxvppVTkX4og8vdQhPX0Y5f6r/Y9sPou2YDjt4vsG2LMWTr8Y4kltIUFHPWwX1He8f
AKH9ztgDZAMU9RQW7DrMxJZLgF/i6vy7gE0IyRZFUJl7Q2EYvK/gu7SffWSCNsfa6p86jla7JHN6
yanV8YeqCKjXO5OVxsyJAfi/bDXz1rzp2Ovi9hV5tfMko/BCVKxqOIZTyhJhGKWNOsWZFLe6EHlM
mPOubUPww5F3F2EFbJDrKMaH0ESduMK1HOovQuz8XO5pzqGQWKv3KLpu7Y1VZgCD8yHiueRFRX33
ddy3Xz2J6uc+U/2ct+oOqi6hH1NLyGZ2PldGVDmV9fwyvf0R7iVzMp6UjxGcyi3DREI0hrtm2+t6
6zamdfhPCYDsT7Fx6WFl9QzZUOXL/cfI8eJi/Sw8MDOwq8lznt+5tmSMTWEpvrm3shOhNpnOUw2s
Lh8fLJo/+cR1aa/N6ve1nNgXnunAanVZvcAvr21tzxwQ4amqj679uKG/BErd8SNj25jusMooKcRT
8Q+jlhQKGhfJtM7Dp+4rsZcE6YB4gat6UTFE7HQit2vBVc2OtpWAQPh/8DwoVB+BZtevKArUFbZc
H+lMGXWa5GshPoFRjExpgmfSc9KawX9cUK9slX4PbrItjkUZPHlhE1HKrc4FT1ksf25F75RJcf8/
ZuKXkc4SPsmh4EqebXYmd6awgm6zeQjRCXNLHZSfwMrJiSvMXEVDzHABaYeIbL5HfYxcbjJXvwLg
e3vvs7mFGnGSYZwpDhsdaIfcQjE6tU28TAHJGYLAivmzqalGMJLewZD/CIe4v9GL2ICs9GmbpMnz
BtCmDStTyLDHAelXgPr3xDoJFhj3uTbW7/xv2XIqMWnpbzMoroN+lb7MULGe0fXTtyNrvANmNyEq
sELvNIckgJDgvUPbk2ZzCeUbpgxEclkWTixZQ6R+jpoffpdVS/hLgy1s1cv0ypSRxyAv8Kh2wW27
5SfwtyZCJeV0yPeeKt60JIgA+F2E1DDiZhPfEpb4Z6Qubm5quyQNjX8vOJZ7FrofekynIrxD8M8k
tzIPVPjQJNcpWoruOAadS+M4iaY9ohW5HeK8STg/Wdt3WjYigPWkTW3UPZB4cuPUm4uYLHRz4brN
yX1Br6ofJZPy7xA2ZMRUNEdQX8fEbadQmnOxbqqKPDUuHgOlGK+OiN9bjf7mn5Tk7cyIsMcP9jA3
sk/fQTWwiM+6fJ66vWfjmeby8JRIq2MZHVW5bNdrk98htoUksPkBBg2jJNclv0i40KYkgT8p9sDQ
SYKKfy+4s6iF4TlIIVVg7RBWWonUgddK9ECIgml61P2yxirvVR1CMRVOAxIyuczhcmqoEgec00MZ
okQKULPfDPTVRU2trKgr0CjJ+zgFXdIPQcFWl+40wgNn8Dsq2EeTShephPNWcH/N4A3s5VURohhd
78CEzVwwBblT6XZO8IymSUgRTECSC6zWWzQZW0L8wUYIm0GuNVo4RyZo/zY5LgzLyVPAKoWbDtJn
Cjg15U8Icja1nO+ivUbzKVwqvt0YuX+PY8cPyfHMkYIuMuDY5zho3AOwS3Mg+2D//6Q1t7nHSVZw
Hri+rRJSZ3XtIixcbSGUr57tN49FBijt0EsgTb7acSn5zr/PZv3YtEitt8FAGZQtgS3VcMWuNlxL
HVOGEq8AnG4iYcIFjssYm/ZnzSS/WMovUBl4jKpB0d/mp2325KEyhQBfCmZMz8MQ7kVRVeIHBRZJ
rhLO/Mvj0R4j7Tuoif9X6jDHTmK2/xvHiZh6ra5jdJVimXmw/z+DOmZYKBWZNjzNoLk2Y409nqU4
VrjE9NHD/auavhBH/R4egjfNfNqsbddy95DvrXXD/TPF565ZqsW85XFNjzFdLMFf8vvJ/k0JZ2ax
MOV53XGZwSF8RDhKsmfJH95yLuDfgZPMqUqpL9GhEN5J1WzrOvFEasAiQdkeR3FpcSOMjKaKoxR8
xC04+kWd81vL4xYylWCcD4hoyuUoO5bbBdcY3c5YTI6P4rcwR25a4Az3tRRVb17EK7lv6DRWXEuj
2ngrKu37mWAMsDZwIahWfoG4LJZCVLotlb28AbJrdlqqhT0WFSA6j7h3mv+53GaPuMIeqiId9CSc
ho4XteFsy4Hjusydyl5z6/Tmdyo++1aTQRelyu9CWAUTgFlnykmRbnxaBPLRtgv42KMDLhFYsvFK
qsVq3j8GZOtLUC8gHIli58BJCYmkfPQUSK42DXx5p/VOI6flPzIPb2gsw3a3y+fnw5O73VkL9sab
+xiQRvG0pnRz8XWunTq4+UA0ABX5OVhfIQM6Cc/IbCDZlt2P3BEX3U5dl4K9305rGb/fg+Imu2V/
MqMJPRxXsqlrp+L+0QjqxUyLjbPxlq643CkCJlZeVuF4i8WudcEKGdKYhXSp34/Hvk2VNXwkrSUJ
6OrrDOCyGz4idDmQDcmEE1VGmVSL3yU9LFbqj2MM+dyjVCUKNRwgkAXc9sKWhXNy5yyVBz8YKmCx
vWgpLEnpqo3f34nC5v2SeywYbgY/gSVkYtC3xWyq5RhUgxKF6R2Ayd6fyzlhcZLLEGiIu6LsXnSb
EJYxl/KCz7peQE0PDSvqyZmhIGNcyvJSlIXVj54akS+RK+rdAud62BBAVYSpBSA80oRULGwm441K
W5DyjI9SZshojSrOmwWOJeG/07UZrefuHON75/Gbjl4P5v5hWac9E6SdJGt4A6x+CX3keStGgTt9
FxCp/sjq+4avSVHH5ARga7TcE1WvWXigYVRBgLEqwszGDcAfvORkLDtuuZ4KFDYYzQFGATsLKhCN
sBYxFZTd3HsnCT3weulc8sWQyJB/0u+CBcGSJTljUMoBuMgjnwvM8PyOD3P4QMyoBRyJ8vvsDect
MmFDd2VRpyCmhlKsCcbsMe0c11RJOlRL1+4Q4u/jizTSPHnvp2EqMv+Ash7J5mPzbFuz5QUFTvwo
3IeOtvka0cP7m/TPd4wFHY2rvkKw9N8QCN8kEmeyP7x5Ipn8avAPOkKzG88lvDYhdyL4boEwKnKS
oO7uokq9Yn8tJUYT+Uz4aW3gpyKCNFjNxilGic+x/LIdEBSMb8oKFymN54jbmke7fYG9OUxv83M+
JNoRq9a6cbupR6zwIzR8AxtxnCd+yer+bah5vQ0928vXNSWLOMjZRw/oraoAfqvwatSca6cQMFy+
q3VPsoDHEVLxqkBo82fXB7pXlQSYXIAp7HdKK9N3uwKLFSKQ2EX9ork01oVYdKiDmkzc+GB7i0ny
DJyYY69pkBQjxnMAnk/YvbCPdTMhaWW4OXqlWGtjRkygNnzE+UO1GhJYx6nDqcXVOhiSlnCTJM5e
yRJZMaP97AQdO9inFsVhBRR8fNP48eB4O4MvUWQ4DvrYqpOVxUdKoVQxuyG+AEWiOSTTjz+MtevA
LUTBnNBLQE/cH6t1B9Eu2lK6j2Q0LYA9fz6AlmoT4jBgfHonOaVlbIgtKxx5ZS7FxWhYj8ZvCG8b
4NsaJUV6WY8qsl7pdiJsetiJIv/QpwFcpXW/gmIdR1NfepNa+D7SDSxHMnBwHyH0DcfkRxRGoDlF
2pMDnM9e70+L/IkVLjvB8uDKrYU+ydf+YObr7yrZPXFFnU3Zuelg2XeUq47AD/UKLrL61arfrXZv
aP2jDS4vC5cy1hnEdOqlm7ywgnVkFoTj4d1AmucpPEoo8+nDDOngEuJUIqtTsny9a3sJ/40v4NDC
zjaWTCmXJkIUSc00aog7WOEyLuRaG4n+U0eDV22HTbYYlXLlLkRZXSOQ4YqRcavurMK+mdQumtcX
obPPUyfPHduRVv2tip6oQQC+UuyoC07fQEZTsF9MKheOnWXXZwWqO327gbP8A7tTerm3t9FzEiCj
Ym0dPMnkguuIZbaWi5qYzsXxwmqCnsYPx1pm+OBFak7Ukg3STx2crnKQ1VthEeJejfmnjEDWPbG+
N+Mi/tUzk6P7WpkM4La/H7Mnp93Bs2/ILVC8s2JTUXEdBM4cezXM7Ux2pktxBnV2j7JmOCpVNSwk
K3j9oanTsyVeO6OeKWasp08TBlhpnxCVxUflNmA5MO/VOHUcVN2mAaKFyrXKJL1BGhjVqn4+i6ZB
L3xPus4d2xnE7MlJC7QtjW+HZ9rqt954qwqdsHYQbNgU+YhTBZz5kEqUmuK0uQI51oIJgCqOSBha
+raPLYMJGZ/SF484DeXzxmJToBJEwIVZ6znGQXlZU1xU6gdmzJY2jrrOgtqPQqfB/akJKuN9w0PB
ADGbpQvsVYMQU09FG8JfE6Q9oOM6P0IiBcu5YKIlKrrSxKGNNS2bg/eNwz7D5+aPK7djnSyCNuOC
S3QYflO2p5vN3hcxlCTVH+o07XfdY2DfAJxDf8XgWRlcn7HXwf7Fn0d9hRr9cVL5CLLLHKERN26b
WP0GYAZZkIAEJyPEVt44vrhEtnc58m6uBiJJNpWnnH3gE01K+oT9jy/Un35/43qELHkq7jSmEsMp
dLKvmIexHQvUSyHI/qIGJiA2p0aE4Twh3cqlHOlehDUIxkX46/6UuxjdiwT8cLBNM3yMgLoU9zIl
BbBsD8UEltjIWWTKSM1ZJA9AEVyK69wWybsvj/NxWUgZkSDJctuWLFWlJT3YtazJHwoNMVgJk3tg
hhyrGG3DN+5MEgn0nx39pDOE/qrjMqRqHjJNEnJ91yrp+2/nkvCgIsEIyE5h54u7kuYFLHWMvqVP
ZGO53VDJ22QIY/G9DlIzh1Pu+QWZSUTzb+/E4IuYaLwwCG3rNa3/eB4XOmobS9Q2FO/5EnbXJX5a
rj1qq5TN2/h3U5Dys4EGzgBna2qIfV/BcIO2KvVQXGkQaJh4D1JFNvn7NZ1URk3T5SeIIS96hwj1
JcnQUAXdyJkuBL+WSH+jNwjdwKw/bP2+v4Mf6whVSDj9fBU0bikPUjNxRnh++Dyk7xpgsXk359gM
zJ8WYhnaKgFW2L5u16pgKrYRVQ4FsQd7ayBNGHEO9073UefCf4DEzdW1ldpIM/IrOmYoN5T2WXmy
mrsEjFOFFUEZnsbTdOc399udAJh5L6+wbhMcYzddBYGJ/rkM0OjXcIFSaVCcmKNipCNmLZz7DObl
giUzSlUUMZPx0gvxR6VCxzi47lD9LLwZ9x55ItmqAB8k9/RWTUUJIQcBIutHMu+XL0RUsWTpGkET
9uqLUIWisluJlNChyYCNEFCDzPbeNklSZBrDuN6+jDUS/QYTuUAL8X/o0u2Q0Nw4ltHU0GrvccaK
1zvKMRfdDe3ly4NwFZ2wdhDFb0FXu78//qZ4GU893pqvcf3em1bMtGckaoYKeu2MDk+vi9eNMuxC
aZOzyIx8PhtDTYeMyIZ+4CowcVAVhVoZDaJCET4UfchC0X48eFoGeLOiMZSLXDJY6keO+pvY/9zT
yJ8Uxfv9sBXtQlLncxeUTgOfuJL4InuE7lWnj8oZuDCriW0V0nV29wCJMT1ECQibbjNX0bMqHUM/
DzRegwxM2NKM4fqy1lgP/Mt+Ic3N3EInsPR5vYR4UF6N632MuHm3W5+SZSxOWx6jGxicgAkaM79N
5b59gp6LR1+3u170oyIY8+mnV/fKQ2DCWhkkp56st6PtZloJSU2HT95PvU8qb5L1nGFZx3FCIwyo
xMVO3VjORewHmZLWMePBfLBZ5b4xtjoYNw9NlSue9zt1CG69EWXw5r876j9o9vJVG1rbg0WvIa+N
OEKRs9fDiaC4GRUj/JUEZuojv92CywOxfEXyHbc4dyk9ky08S7FTWG+SYTPN1T/cuQ8KTypJWX8c
Iey59imWDEJJ1ZoCXMdXg7xf9Q7LeYKc1EDAy9esC/rGkdpZb+mQL//eo9l0vr35xN/+lf8QxRkV
EIHJp+xfkPrZChM2YoxWsInu0a95iVtSsyMqE4E1JDOhgoZzyJ+Khk9hsgMBDKVoNFVkh54dMV+k
EKgZnDMVlWFFVa8YIB8yKIfnJkh0pbu6tVlR3Jdy/CLJLoUsZ2NPnXBrK73kcAodTliR8E2CdUlT
jcNpZwiHZEvcgw6ZU6tZDWGYAtvz097XVQRQnWHV8dtlIdmlGZgDM/ugiADb9r0lePam3gt4cify
z/aNiqd3DaEQzahS7/8zb1Jt6GTaXDZm5RZOh4SrMaEb8r3Gbq7EKpOnIloURylUN0NVRJ5EXLvG
O2Md7QKkETd74LDu8ZuPdx8x6W+tY6cd7qyDh0cM9+JjHaGHMI488D1UV/XNNKQ9b1HOvBDr8RpE
L6cHxfpDjjThfVXuhjRO+qjuplSXltyg7cUVOVduy2Q2w8vp17x6Smmn/YI6gJCpPO8uWDvLntvY
TNYE8Mq3XzxsctmVYHXCrUfilDEIPoUq9WpXyraMidL7c6yttQxrD6+m2G1O3jS1W3a193J35wTm
PzIgFdByzYoiLTgP0m88XatiTw6sGX9fkR4Bth1ThmSzMy8c6aQyMY5QFdi+QSgaD6flPo4KOyBM
E7fdioJNLt4CFsWknyNt5EBv9YPtNqBBq+HbwA55+WAq5sGfTIc8UvBMAHOfKEXMFpt6mGrIIOn+
X6LElB9yZC2W42z4kh+Z/p/d0lEYZ0wR8Z7+XkZ3la7ENnlr6n3aU8fD14vpKOaXy+mJJx8eec76
adVJl98efalb44hpBUrUbxnGLpPQELKm9FXyx6dMOtros9h4GfReO4aCGln3ep+CtLzD8pTEsbHa
ggnWRNnhL+7XzBAYJnnZ0oYJfHknYz6yeWApgPe7U3KCxHUuO/kBZNaewMKm5lsy3m/KFMO4iYu4
vxIK0vSB/o+SFsOO6OJWdvKVEdPfjU07nDi55a4K9C+9oe+UeWJomeaaEr8Sq2GUw54gomKog+sB
JrWbot9q7/hUVwXhw7OdM74/BWRXLebCygqjz85xFS2Wn1nLQBD5rAzJJbWbeQ2JsjrS3y7qL1K1
LpTCcKcujypBYF5wu3Lo9ynkn1tMHsXOhI4U0APGwQtJXZWNu6qmQC9vBPyXM4al+sG+qSFl/nin
W3t+wrBF+nhS44DqcSqrRCLKXDU/BP1r4mSDzCEMUuAQ4peR+9ytz5lXrZuq0wmyME41bwZMgIQC
jp4IPNPKg1MdUOuZ0Gdz3tQRA/WNAVdsgTTe5DF1PAGRfXGeDndjMYd14BfqGYDnpJI109v1neLe
DpjNSuBHcWJ7ofVjsujlv3LOSqYt0N3CvwLD5VlfJt3+e4Z+vNDnkpNkbKRGxeMfSZHWSAWvHndN
Caw8F8yb2cdBVz7+Ev1O4g327mcF3ReMF/1SkeJPgn/9pBZrTX6mPKstEOsQ+Q7dh/6R2IrforLe
ruk7s46QlsA8QdBqf2q8MySE5Ib+VMloLdIDo36q+4kGiKvxlkJ7l1fWoOElLFh5VyEuh0cQ0LBt
zD1p/WD+ye7+MmHyPYOwa9+BhY0JrM42OuAEjx8Y3b66vXj1qSUQax3zxkLoQNbGAsv7m1gF4yII
w//Jro+fknKObLC7Xle3eiHK1es7vkXD83zSoLa5/9WUwhNi5UbXIHT/R03KeQfaGQewmOP15Hup
aoL1C+qiWI1DHpRZ8mw/9EeVT+59PRu3tkhLH1JApnRhOj5AOzbwefCksrniG6HmJNEHDcQMVgK6
Ip28mBGDlLSLZo8zpmGyS4f22+/Ow4WNe525bRSLfw0UQHcAx8+JyLdLlNO2yRyUn7Ybghp4mzjl
k1E/2vbnGg1IJF7RneZ+OXQbrG/b+B32PfOlat4pvLhqLT6uKCyOBKxdxCgw5f2VqdBXjt11KotW
DmUZgothrdXbI7f3oygjW6CYyiUcIbJ3tN+qFza8NXd/k8EbDl6FpcWjPeTGkAfVgg52HKqP9tDm
dCbhqqNYIQ6S2z6ExHzuoF9uWWt3r/7Ku2BBfFLBELGXcs2sdLelXc427uvN0MfveBXlVNZIe36e
ocM3rwiVTmdjO/RrUNs6RyduckRGcYLZqpmHYJYQ2eCZnU9KBUyoeSuMYcFEVgGa1BsbXaxBWZvP
73QsJiY9F73C0tYAGx0aOl4gTKmviEZ07CZhnWnhJ53jlY8J8oAf7J9n4rDbZET/tmoUu/63OIie
Rc8cYNHqgLgynD8WheIdJwbNxBbOxeoFC4eqMLRV7z1LiHB+yWdRGq+XPh1eUJzrLxFSn+wfuVVz
1d20AEqqRaB7FaL5b7pQu4OtSbP6MJlytYdnTj/gfqHAbSgAKl8faNN4MqYFEgyAFqqlghI67wK+
uhr6lVBeW3MH0ugez51WoO/WxXfZgfD52bp8tki1VBdJSzca4cr3TL5GdpxVTFMJIuj4Si17otpE
Fiz0Klqz+cXAIn5w0yjsaAYng7mvvL69CC6CeOU0R0zJ9l9Yk7u7JdeA7gkAMpkgg9/jTsr3HHH9
t9/ccj9FEEfB2E0vrYoQLdx8DW0whxLVUBQcXFTVuivA2YHGaTSCNVoRdavwjIMVknJNukMRi7vK
EnQBu5svmEAe6iMHFLKxLDGEcuYlB4G2FUE4RBelLXWgDLXT2vZiRqWOkj2Iva01JOCNatHEZJdJ
Qxz1Al1iyy0s3OCc+HoPfqSjOVeu1JnKkIEeiW9QYcPTVXYgDZOT6Sf+1Ap8E8tGr+3VbyCjIgtB
ZvPMoVayKsyPlVXVUFaMfoVaANSnY2ZDJP6/Ntf9F47j1sC0THZgPVKsbAqHYMqhZRCGpTZwkKr2
Fo2v3xIfQhmaXwWmeiBv0O55Nxq+8JBcLgYZC8aHsTejhvmyhEW/hhMrZ7ptTxxkJB+gDpd3DuGP
PQ+2SL2s1B78XaB4PU3mk8UmiMo/W257TdQ1lTmSn+i5vAJZ3ZN+6uwfUCGfEJCUg8iEIpKnnCLI
LPKJ/6ai14QuUCgJcYF0+YFRYKOybB47AM1F+eg24QyR0RH1bgOnqhyf7mb/k8f5eubtu1itIsaz
GopzvqbmijfLb3mnyQP1/t9bJNKnGyAVYuCE9mPcILuPLhP0Jpue7JvvNTtFzJ80pOtfXnKVhP0/
cP5ak7L52lf48fboznS111nTjEIAIJ/11T6kGoyBosClZXGmfpNUKHxKJE5wVqvEpO+0CRASnlJg
fm8XQnxFT2qjB1DT2KcqT0bD20bYgAIqwBLMOOM8eJDETDS0y5fcZtaugf/k2Wt6wsrsWaXG4Fm0
pyTRBOn1WQkQarh+/2tzjcotM5/ETjGwZCfARXXU8hvVkJE4glHrY7dMB+u7D3gxr912YE2U5Wh/
NKa81Ciw/FSLlISBTu3kphGZSgpwHFGfD+hCcop3t4ZTfrTLwTI9U1FbwN8FYcnuzU2jxLdNsxj5
zlSyNm8YZbP/Plvg2JGUXxCFsDbbTX2bak3BKYj6Us8nhW814oP2k3y+m2XdIhbuETVzjxdNp4/t
KDWf/5LfrrFNu7jf258AY4RXW26Jq2oP4eFtWnwVbYbd6BbkeQ9v1rxKg8kv5AiY/d5RhvNV6R1f
NgJwT+3/exzaJC8ufeGj5g7Npr4Bu9a+CnrYpS7vIEe156WLQXD/vaMGo10JapCeTHSuuqYnrGou
kWMDvvtyYY3Zqb+vK+1KvJ5BHENHOFQdAj8cIxoF/bf02nreMw912CKHVpCiPXRYkT/dMZmJn2/R
gWo1jZiDQl/ZpmaYHLrX2jfaNtrgKo/eFEh1BawV6Z3gOvB+nD6BLgXtA8zvXd79dQFn1gnAxdLg
F5G5uKMMp2ltaYisqgqoCzK3T7eYXAIRX3QV+4kE24dMfPRE+7LfXnCYiHiAqQpzJn9ifB0a59wg
rC1dNDAycq+Fjae3o+4+k6b01llNjRkiKt5FAn0Ek1n39UCskYPuBxbg4zJDrTGtipIQPG6ceUjK
T4ME0PKv62fISZuB7Jo2D4yiZGiTiIVZi1NjBMUd2nDgJnUomLP0zf9EpJaMWr7dQjI6w/vOpS3y
8/QLXXpZNlVxnrjLTZFwuU8iJ3yXHeZSUPGyii1COKkvU/fhtZokahtINSdq74lB7JlrmnaxQOSI
3lLKwWF1mfC9JdxZm4S4npgVxuS8GIqZO/wvFzu/zOEvJ/Zq9LgCg3TDvXkBsqVLkUPSi4bFHWkg
SO+JWPb0LBT3h+mrixfFDX3o3IbqduMqAfY2hgIuqkDs+1AyrlK3nu8GGp2XLbSHy3/71e+zN3Gi
Jho2vm/XQ+2NxZGukIT6e87mZZYBt6ysGJbibGqxm7e3Q4sb5SOpFKAz3vwlLsCn++PmbO3oPgVN
Ni0tnyD7RPFUqDQWNbK7jS6cunGcp9HXJowSQ1yl4JUjt1MvOOashgTpWDB+e8K3YhzRAedDt7s8
5DZRiHlQaYBxUv1u1Cxk9UO8z/Jzb8EqtVjb0L7bjmbYg7XIZl4VXZR9dHKkq3ERYUANQDYzuIcb
F+kJSs8FvU9reyi4KY0VMjGe82oFuqMWFBrjDu4oMI16MJoEInJGbRef3HmJ1b7Qbi8flIn4GI/+
GUfU+Ri5L107JwLPcRFtnERzLsqQ3Vum0gRyYINu5Qrh1CmDyzo1PnuiW/rTGnTpqUX/pMwnvhdL
D1tZp9WQsQBGVeo/KD4JIY/ZoVEBP6X9GjizZzvRpVe+Hk5OghWb+Up7G2DAMWnL0+iuwG71fbN0
AjHJ43KF09dSMRHRufsNKiaG/GjTXDqS3gzA0kG54sVz7KgJCrs7+Cr94e+ZE1uwznNHZ3ugj1cv
zLpHRpT8wFNV7HLqGLAlpyatU3xyj33YnJAAv5hi93FKwrldeaNhN1xqGFuh54YYdnH9o6TTy/8d
q2XqbtQtlMhIwffXL37UMoybzwAMJBeo51ltHsoP7/ZUu+nmV7xPTR8Z1xsuqdrSUx/2BYvlhI+0
O4ONLWos27S/n3HTRCuLPFigrpXtWzqWCbKVpWPppZWOpS/WQmrA01XNMSHqHZShcSEoak0Mb2LK
Rj7F3BD37Cy7stZsuL0wyrW6ltjC+Y4pQ6Tvq312b4kcvL4m96YDCWuyKM1L27VGpVVx0p10i9O5
MNjA+Npl3TkQIEmLOBzUpwdXW6NTeMJcKIgPRkHPwX268alhA0HPtF/MUfXWvpYFHTXwveFVyPl1
gW/hxXC3lKq645O5F7SM3YskV7KOA9giq+WsD54QK/S3+Mw9whcf+FXzMSN8pzTk6JAQR5xFLu0E
LeBMbki3OWOqvLnFVKaHiv9FwN58Tym5PiyTxi/1eA3FrTQGP/4nXLAxHTe0XQVMNbBguTCWZucf
SzO7x51BYpPJeNLCHG7zWSIfmTM2sMyJBszesdBFkJbs2VYC5wljsXL4U/cUMFH+0Ij1CWb2zVzy
nTp385d4fW/CIKlGB2yAez4Lrm/nKNV+BAICioE/eN9cE/HM7XuSS0QgH/ZjOaYuaJbWoFqYHTfR
1Bsx60QQYmShvZVYGsP90MYfB0mqpFH46YiUcY0BdGmHACSA5i8yPJgtjNEQzPrN2ffX224bMH5H
e9ynm6Lz6bUnX7dcB7R5ZzAb6oGkOYUf7g893utOTQOBekBnHA3EdPUPXtputJrfr7AOFtqvdyeK
xhh2FvZ/bfAHT4Sni6dsIPfhFKkCzZuudmfo8euDxfWGTEZS0GD7N6hPc2cD4JZn//G0AN+AWruM
WfJneZ7vpexztu+l8iKoax6NFMixzT8HPRzDfy8SSFlBxw/kj/ZuNiNhZvbtfJcM3qAzUrE+W9kG
P1GOOUMeFhhAWBcd9elp+6ogx08cDQcPhRVl60slzolv09TJrSvKzLsTW6/DG16AhpMLBaxgnu8l
HCYzhkQnWPhGPZbzIM7vNLzaBFWqFGYuBOmuAkZolxxjm1uwLTGNLtxhpeiACZrybo2k9sE7+5OA
6sQ7ydJz8eSiIQpDxM5C13a3dHgtvecT7pHAwJVw4uUIZ7ZnY2TkCnF5QiAFoNRKx4bPh07wScDs
Zt/RSU73KqGVfkcrbNCWhumi/LFeRzBZWuwcx7Pr1sxrj4wLl4DcpNWtAZ0VNSWP2+xdAXtAdg/G
HemGNufXnJe/6WcxLjWdTspahAnkC+d8mPEmvLyQOE+6fWahYh/Jt5FbSOcMPE8lj83fugmNby50
t1R/5LAuGlwxaJdbw3/RyYd1iIiTArvyWMuk57vXEzHrr018+ascEhuxDHYvcxGB/apCohZQ00jb
1L7D0ju/ePXiZLl+wJXiOIXOv1H4frziGa4mmRfB20Jfhl6vPgR5rv13PenskcO+d2DY2aiWcSWh
yQRkYkqMrfWvW7Oi++2kr8VMZXDzY3abAxqtYFuC3Vrfn6E9QrNwKdHmHHSmcZ8CTHd2Ah8/0f9i
s+uQZ6KR53naDlCZRgkfUQA6G9+FZ+D5shQ1G+wB0RgtT9Aptkm8o98wb+9kSwzFfryJyU0fWhxm
BqV4nflYsu/th1vvLojPAAMtRrYWj9yd7aQjs7UFEAM/JoSCRF5j/aGDtHXC17CCZ2p7ULYrjdCm
0Q6ZUsoFhdyLWvflEer5CEcmGiMgG4iveaAD9/rHGlTsfxxUrCeO/73tkXmyH5TTe4vcLIoq/SxW
nZtp73shsk0a7gvnq+y4GpegKjq1v5vyPbwdE/QfC3x09APv04Be6S7XlaSZzuFc6Gy8V5oBftQu
CTfqs6B4DSN+lLDtwHOmUns/BrbpIfIb37qQZ0mNHnEueQhmTMKWxRznsOLecEgGjsTtUTNuxvzC
GdfMDl1ZrqMoktoLQq/ZAjjqVz5RTLO5dVXVgRxlQD56N9eaiEOaa7fdKuyKg5TbgDJf7eaZsT5J
/yMTn3vkj9L2rXInA8VhzKMKIzAQApxIV6vROsiQgYviiKC+LPw6pyDRSYV84HTbc8TjzxUBsEbP
9SHOD480EHX8G38jwkUyVbDJ6BQDHKXVUZKES+5UDh/rPNeyBtX4BezO0smoiQUF9vnmMGTvcPws
yyZD9lskEWssuCX1JfhhLcNDTW5h5wui3deuHS29YCAzImtNafXkz3DcK8dWrtTKot67mSikL5Xv
jHrhDhMOG0sjLISOztgOpheSLyT3PnZ0lh1FYntMvB4856aSa1HKpx2mzeUSG8d3B5Iux2/G3WPA
MSGbC4ZqwdpXiVhy2wPfTO/+Lwu/7snrMrN1mg292AoefjsfRc/eooRox5ahTg7S5Eh5O0u8qiCC
KR8tWpvUs6Z1wdtK6INUB7qLqKYi6timDPyh+Tn0M3awy0zNflOLkpOH5dsHorqB1lt63eAVLLnp
GmoNTBqmBpnBLA/3m2b2hnSrRqCF11Vz/Vf0NBPAQ6DmwduZgvZnONjHCjli8srahGDEwJfIGPfQ
2ef29xNXPdNJSJ7SjHCm/5s/5qUYj6MENNPHRzhFOy3gY8VTRNdpfnI+UHp9Wm2HK6Eruyv0D8ZJ
TFEprK0SApmCxd7kTvDzbfz7FPSjr8u4BwX+LdFn+JUiDlPePfVZixC/ORH5Yyl2cho9rLVAErtm
LxjweQt1pLHIL13ZBDtRvrVvmY5Yhqks6UX82hnCcHnOEl82UzIv6zda9WfY2YvHWBJnj7UvQBHx
HIZfNIxZPhK31vSpEfve4lbAuDbb1Q6hO63HJJx0lccv+6MYGlbcG1wBw2gZ0p/aJRKn/riPVdFm
vbmZnnGNpLvSEbnpOTMjCCUF+c14kkv1LDBZCaFuk/BA81a0EuNB9ez66C9t9SyYBzSarMix3dlc
k9mlgD+mYEnYqKDd0TvMBJVNZfF4fgIaA4Fy90npeXDwJB3DbA7rvrT9+n9LeEr75L/MKnnXCbf/
x41Zoo1n4sb3SKB9ziJ9hi2Futi+shOGKZ9qpzi51U2gp41G0/MWnX2Kayfddd9mYL6qwmymdXtP
t7d4RtQnqOLbR6quLdL1AGoK3u2nt/cUHbXL+odecmoLRG52DI9pjnR5W9Oq5oBetrjLNfbdYUow
h7P1YR0cYf9z/LOMszuUoHAx4Ye2/Wqy7KMyWZvQlzjmguEBbytpfATOM1Bff8cUKlHkoGkW1P08
jo96Y1xRmHkUD+I9Z6KWDxuZ2reCWgL3JUFgw/sYW2z+97YuZOKLCTzrJvaDZLBwvRCamyh9F6uq
dWoYvD40mA5vym4jQqLQriY+XHxqe5UnmZswap+LHZTtIgonRAmpDT9+qgsaEWzvs8SxKf/RVFnF
MPu++owmDQSBIxPaq2HDSVt2uQhK9qyUYqfGgvQV1Ksmu11k1snCisH0/3eSuWbbb4+xJEdJLS59
wSy9Vok/prR88RUHiUuKwp39WP2sbMVdVtLIECAzea+9O5HKokJPCzkPZ0WYnd+wFwgXBgTL7aEy
YfiEhbVxkZXrESC5qArLh9BjULnMLtdiyMMnswGg6DdQDy3f+qpVXUr4Ol9QfY6iWHa48DQxH+Ca
FiacqwKiu8YJ2cPgf1cyWZCemvtxmoc10LqsHdOgVgj/DFFtPfJHXdlwFv7xEdKMA962lwPxzLQL
L+cj/dzzu9A9vGr002ZqCs7TMW+skBCGa4P/eReTeDxgh3SaEFa8b9dhKgvxQ9z7LS+9wWhyxGBA
EJZXOcYlY1idHj0RBqxAoxMMTxdMw0H9dU76ewhs1aWs7pNkeUMWWIRgbLZ8dIlyTxYt5WbOO2lr
OPBHphRorW7PlhiOWHu7TYmtoeaqjO/b9aI2xCh/YbSIA3lgHH+KjvXVgj+y7plizdfqAvnam2jO
BbH6ud/2SyUcVR+WDIMVxryV4CQVymVoghuI+ZupFgLCAtkkYIC5YpahFtYb1YFL6iwF7/RJRuKa
rDOMWKbz40KrgWJhgSQFlBAkVxE1kYhMf72weYBD1g+FcVBo1EABQRBD0K6tU5BxWl5TE2lKlZb2
u8Ku1qPipf6z79E2+qeUKAh9UpbSWHrHT0GopG9+ZgSh7vkOHVUuxd5xl83Y6ZvCvEPUvuuCzhAQ
hzO5yAXZmDYrQpANjl7ZPtmNYNMFH2vfWORCqzRVFyMPqbqo7aBzrA5u+nmeig8Wqov87pNcdiwC
VuU0xzEska9+4/YFUOzbpAWO0kt40wjvmIWTWUMdaDy9j0ocR+zGTxV+jIlOa6xWgorUhyTpsNP+
KI2p2YpgBz0khJ+reNOCTyTDC70YaWBov+3X71Nn3stW1TNhPIOlHIzgfGIHynf1H8f2nSckPS0c
7AL7eBNFHRDAUTlc5dkX0AafnkJ3r4P10CEmwZ/ChtckUrUEo2LCFmnBoh6iLgG7CsO6n3Nm51i7
hbr5uGhVsxJsZxPG0zjUOrXB8+HdvN9UFBAl6o4JQKLX3aQwkqDhdCkMmz3FKy5GvJm3EOWAxRg3
uQ1oA0o8s/dmRhkqsd0ttYl2Qyfjx5H+D4toGS3T6FFSWPSp/EdxTmg4GhJd/C+YMlcZmDtIg8sj
DpExS6XcZjRBmlcm7ry6gf8VpcoNIT7+BnnMSdITRu+fmhrfbml9sHs6CRv3kf1vKQVW1WNRwCH1
8wkZg1MmMfoLCHoL1Xwm9yU13S1upxkSzqScHg1AFY60cmpk8Hbpr5UHk9setKYH7e3PgQ4feqKb
g3W0KppC9UUhmu8fpuBQq+U9d0qrn1Jvv31NYHBNfVkhFvOAK/l6B24GF38zBtmdQdfLY0Ltyb4P
aD3fWmn87rusYhlgvjKQcpR9CpBs98Ey6qqVqFe8z0DZfCBur1yLOjJX2t0tTKT2M3vn8K6ANQcl
GL3JE21eRYcC/WEfoznWvF5wayPpWJs8Y/pNrtoaUe+pwDShA5L5QrkksuVdVM8s31GCfwPKWFds
NdOirXWlf0dJYUXaaKRGi1BaqOb6cVVdYhO05lcWSKKTVGGaF1lFczn6TwUE9OMps4abyPQRXx96
Oog3yNA3ksyNDBxLiGJbp9G0gfE6Z2II7JP5tINCYGr3xkQFQH0Sinx6Mr0lh5n8p/zo9FpJRkEu
I2T1tTi8BfILZmNfcZO1lPt7LBd9EzM7wWtliIkFeMYfsHDlAYqWalMRSLI4JWz1zGXOtCADyYCW
Qf78tORVBrbMCOz42c24AhNtq6sbE0vR0aO1KgnRRpk2LPiLtQueYw3x2YomMRUy+KfyEwC1kt5+
nH6Tn3+CEAdo4lOrZpui0HNA7tALzJv6AlJFAnt64Mx2GH7uNJJJIbKuTSjBrNjg6XIv3S4G1Qaq
2o1BokeoLPgA1XOjAHvQ//cd8ck6LWbC9zsoUv+b5SdWB/m5BNofS3dY8l5JpuX58Fhb4+skl01J
n273XAqT2NUbYTgXZ/ZhKdFxtapXwbDgZ3eobFfXO2TNtZ/nJIsZUJNH632Nu5HpEbmlWWtxfr6o
jEveaAf29g6CK3/GdJ6n+8C9eI6+3dLrLU5N7+aKEv4UXnM3Dx62ypLNmVxnO4w+yZWc2Q17w2VP
tEtqs3aN7e6JW+aQNWKScLaduvmkkQVtzsvztl4xh+fuLqVkAmaF6iXdq4oEod0/KD1O+mX00bY6
yZG3x7DkXTJQ2uOWMIPPANm6Rg2zM/gCfYYsT2V4e3MQPFLPqULZmxkyIsnPZUuVocDwKa0xoMN9
Xv0HTcaLKWxkOJonhST2cmkznrpsCbeQB5ovZQB05URGWchdOFJZa/uR5sv+rfcz06q6m8tNB/wD
IJIe9VtPaG5oVRgpFktQjSgMz+X7AdNkNQILLMTqh1ptkwLTSpB9e60LiVBE2oLc12xTzmftndKV
J/t1AqXuEJaZvSAWUhbwPbGj/xbG/Wfy410AQ+eJoyeVWP7V0qa3zh6AC6nUlKcbMhQWLbviSLBg
qE6TLyPqT0Ao3N+nq2UH/EXtoT8/pgcnKlZeYTE0gPXc/R2CjjpXL1cco35YhEeqfizrLGSKU1kJ
m7sKRJqkjvV1U52j6Kd5xT2cFSj3tcI1AE9RaOSadThOrQdx7wsNZ6G8w5E39OGD0S43LCD7cLMT
DppfnJHKU9x6BU2Uf4DK3W3GcFY59/BqdwuTG9UgoXzllTI5qsBXYET7GxW7AyW21kn4PzgNZrVY
3BuBS51iYad2j7f3WWWenPiVqqrhcWbINyKeIozssW/q/KyVKT4tT3KxLXDQC6ljQM4wCmq6or7O
1RFcdOdTzdMr4ZVVNv9YmYIwNBx3/FztRnVLJGuiyv2oxlmctGtVCeTqbx1M+ilwygseOIliWWfW
aUsVu1llqll0zLmZ4ElkNsRG4p272064pmybaok9H3iyF8nuzCNHsvHmL0iLs8SIZlxMNu40+ry1
9wnUosBg89cRYQeNjF23DdZ7y02GBYp+pStrpPSNVxgezgDcFBBv90IVAGtwYBgsg3g09KKCpjpq
PmSoCyZ0p79zcpNtQe9rFMfM+FlBLb9cOqmUzIRBm+EeFkN6hrj8VE/jmTkXB4poSphG51iKs7nE
75HUDcEQdOOA8LvOgc3RBQVzV1pBZU713KNdqAtfHjHVAvmAIhoQDF6/Q8dx5DuEgPO68VlYK7XT
DZTDqsIRUZz/CXGOnGJFLCAXu2fQ2pvCgpIro2rQAKYakqvOjmx4ro2V2w/t09AL2kqp6XgvWiZY
KqLRLYabFz13YtJxgoxQ+38PLUQ7fX+rkOnOsUsQql5+H1FKRAQ/V2S6XL1eO03FVpTFsXnEOEIU
DIt5b0GA4xcYzGIm9HvOYp/n5YTkJFvE0CHzygVlOcfPUzz0pj+CYLcjWz15ejMNQLcY804kOVwq
qZqqsLuV1FtI8gaG+ueByqn1FKEw3kIoI3eBmEO5r5Vn9eNdV/u4DTE5pQZbVCjIUscacfqdcijJ
oRyUmJlvmBDmB6oZfci8J7om94JW4sWUGI2bX+q3GL/1OZb+5778AYNsXW0CEiqJfU81kfd8q2yX
5aPP8fI5w1vHja67K/GxjTsywfko0yDFCumMCZ5EQ8WeMJjtBB+WDgI7sNQWVg9nr5nB/bU7n6ak
AajZAR9u2qE8TG2UgFvqIAULjnNX9EyGhJIcLLpezrj92mgNNRydVIXrFWnybHwDhBOQbX4I+Kns
FglR2mtbURZG0MIdrBfhc0VyzYpM8VfRr55KA3J90U+JV1XI9YxZ4wWClA/NHETrLAErvcjb1Y42
zzzSP+Aw4Nn4mRsVaThpQoEu4FqWR7cX1js4vtvEkgDM4cmipWFIctzMhPiiAUtVH6X326njl61o
DW5xA9johGs/r3Z1nj1vbyRiC/8e6ucFVQKyXi34NiRIY0BeLSVIezFcscPNeH+JjQaF3gPTpao7
xyN1SUaNPePS/lXBZKj4WmbE7nWBlwPCz6/B6P1fMBU9JYKZtcAkawmnS6p0J1D2mHYCMImvf5S6
80DB0tz8HUEkRC213qEqEV77wJhWx8o8sM27hvnSSiT9F0ponCSp6kjNJsqHmpyN9Pyczqyqnzwj
tiN54K82iOukrUW+wlcBXUvOfoOQbdVW2R9pR6EbkuhH38YBXsefkPxCRPRpSOKdoNxOAea/wphs
j/a2SvM8xLlAOxptCOY+bjspgNb7z8Csn1+0NU+gO3SXI2tdCLHmkQLuO42dotGssUWsFKkaSN3w
290XJkesokPpI3nUiKp/zieV0hG/5/E8vIrnQj19ONCcPviTFWoiRsPIn5l6qc+W9BmBpw96empx
CoqX/8IiALMVFrC0gp1h92krSy1v7l/hZgrOGkngG827j+/egzpt1MtGdxa6f73Jz5wk23oobsGX
twPZeCCBejS5NNKR5/uWVO7LqQta8ZHIPV+pYASVyRycs9a9KkPJDZQ7Kpvj5/Lmf7IxOJRy9bvf
dbDS69Lo6VwhX+Y53LWCisbhQ4X7v1BGheaC6mSeMs/7igmeGcJNS74dKJ00YzlI7HWd4bcSvY6O
gqpS1EEbFHlhi9jgcRso9ogA7tBQhyF4utNTTxyXn/p8bTLb8uCOmPpBHUDK0uD4/H1MGXwdKAkV
9M5MRAWTSAC2x5lk+Q4STEcu39t8/yfWTKLKs8KkjR7O1IXuwiZu/VOk2DYlolxox7OonZkSSf9+
g1BjxY4jiXPIrjPRCxmIBpvp4TV0mfYV6qPfklWTrwmUBqzD8INVmN/9uMm10UxeucRKnbrPkscr
cwWPS3YhBLUIvUu3dloap+60GMXhVR70MYQN0yr4pwOLmO/zcIgrh+Nmq5pb1LU+B9NSZPwBRhJD
oyN12iSvzDYDhNtXSO7KFUYhEKxyZEuzKSMJs5fRKb4v9XsR9aL2oo66ZKRKSHqRaCoJRuLi62Ae
wg8AXaZj6CWeFEJ0pHXOYipmZcIRxhipIqE82NXwgD/zpBXd3QYX2oEJqzOoshSvvJTrwEJd8QH7
+S5m67T9z+QD051WO0FMTdedz/OpmL1LnNumHWB5zMTG57XMNRrB+pcojJYyJr3Zr3Kvl2EzjeJu
o0aQKGatqpKbLGg65IEnLxPoz1yTA6ioiOXGmo6l/RntKERQ6w4FfVd+gMKdQnmhHK57H+PLaHgk
TjidleA6er83ORUr/T2/lhZ164jKPgPUTGEWIalVMlDEcqnz2gqXkP2zgbNoGe42QBOWyBZwhpzg
+FKNNRcLv9wpgyQ7fZq2zPTqVdUTFdBtiP47X6SgHRAg5nxeM0mPe3uOb8OFxqK1Y+7Iq0JL2gmt
uMpgPDADakd3CPy1M+Zslf6ycrhqLxJrRqLZRLmMaoXBk0JDOzgUDW7PqrVXe7amLd9Qq2llrU19
BquuctCNDaBC23wYFWZR/umInog14gqlCqrcfqT4noEQSVomvn6c1RluS1e40sfnSk9dTdWWYjQt
l/hGwF2LwPM3DqM4kUwDUr12TI84O7U+pLHQZ3DqivfU7+w3+Psf7SaEC77c5hR6Gf/LB93w+wnL
vw/kHmFAUaU5G6KX40akcIg6kM2FkbpB0thOFlRcmNdF5EuQXh58/njnMi4ORz5KiPUZOpjTYwom
snNbb12V3DiWVWhU/5pVzme+IWXrylfZRMG8ujrnKwqfN16RsvKyj0ezLo4KoAwNT2MoWIpPmqgi
Xl+tgTVrxikDrbUSOhHF3vpZX148C+n3k0wnaukFgHUkLf4qznFZSk50WxFq/gDE2drTjTXIbgMw
bNKYTfuZaXO+7oApEqbfHJzOhTpmynoNwkeIdFeLPSMdby8indED9NJpBXfdETjPwbtvTSgH32hq
NOs66Fh3YKB4pseZxtEXCuye8XEAfu+HaCwRcOkM8pKgHUuyLwJiLEP0dhAC++PEUML6CzM0AFOU
DRcpIm84ghQC4Zeq8ctcyPfNzGJqbY/fAAqJNwxIe5cvY6kjnpHhqzmuMW9yonFYiDZWZKCIiZTg
zutf4Xj5fHPdkGtAZFldt7DTb7pmAVJ7ThV9/yT5HzJKdzTCYGWvEVHcu9SZmYjU52ZSPGbJc2zs
DCLD//TMh+pHe503Rk0JuVUP1KjzdjFW0vrMC16FbKFAZdOKqSu6emRJsfGAtxYFS18RMw9jjGXW
iuJrwyKrrFBQ/glL0mgpf8nQ5v7FppBmHQOYeAcaIfEU84Cj0upH44n66NaolSpBThOKn9A1RlMo
R7ioa+P0kNf0ErGA5e1rOlLMowNqpKdGXXiBY+qCn22f8CJZ5PCVad/EGRgW1Yis/MZSWbOhJ6bh
NFBD8y1/lQB1bez8wb0YvIaHluzfJzIGcP1W3aMatWkdvmtqZzncWTSIbStVay2+3PWb/CgEquka
5W1Oea98C7Dl/vUl9yfJATygIvw4C+T+2iKFXnxBUckMnRv4faUhsQez80NFNkwLkQnbXJ6dJtz7
wj9n3Nd1KfBAHr1QBKjAMQpZuSMH3RgGIoxxqIppx3qZdK3Z3jwwSz24XQkQGmIm9D2i/8gj3NXV
qv9DcAig32wn07bW6pY59I05U18HQLIEcutleL9Za/nAM94j3+Jj84JUCKijlRPAYAwjadbWgmZj
DjQagd8CJ2JYpK2AxK7H1aayc5khXXrL9kA4F2jHqkJW0Q2KnuxMHDyyjmcEZjVCNa6QGOq4CkIH
pzowAtpSJZzWVh1MJW82lbzvwYfXXcKXxbt45miUKhaigbnUV9KCnw9C0C457HOWFpvVpbP2ylri
Adljcm0UbULkg2/34k+9DAoc94pkGzHrHp5UxGkn7wpi8y7PTuMyeLqjptnrDxkmg7rsCk5QMM6D
KgLXtwZp/gshrL2n2O0zRJRx7pMIDd8PxAcvAXs3PQupCaoZ5Jj+PpGc1FQGzIn9qaU3BEHM90nn
rwPuA9fj6UYVXZPKzah33g3ILnp0XJ4TuPbK40s33H/OIhGvC33zT42IHhsH48GDnUP1Fnb5i6EX
m5nuLXMVkdEZSLxwVQxJ+DOHtRhJEy52SYy7QOaRwcTt+pwafoy5z7VytJnLFsgjH072WWv/a8GR
bAF7CL314gTf+OHnC3QL8vuG+IdagUYDJsCB2puPvEc3qg8mRpb1QoMQL1iudjBoRSSuKGykR1Kl
KYpZgo5Ms859UTmAAtgckTeiwWWxV4SC6GWPcEHAcbwxD/w+rWoj1Ntye5P77etiYL/ld5WVe0rt
7AblAuO/ueYDDPe7cq+gciwfJ/YWY3t6Bq9/NwPQvRfQpspqG7AAWfX3z7bO+WKc2BDZtXl2ltJy
bE7GwgbhElYKbho7qvMYFfg2jXheApAgxlxNZ395cnMbDUaC9Sx0FoUEcjAt1DnT0Mv3Gyr0Xt7e
liiqPvbom2uX+3TACxqII6aZQvB6XzIDrb8HKi/xMbULaNmz5pLN/kKWX0pP9QKqHqgo0PYHx0R2
0XPkNMqIDoY5AYQFuQ7hAfkW/b1q4tG5ju3GYYnaybRiAaAhpvToZ6cpoZLtTjaaE2n6cylCpGPX
LHwnZV3hHGIUH6Pf5nF7pGXJ+s+gUe0EPXS4eYLSu6pJmns2VM7IHybTyo6YXI3bx9AP2pd5UNex
L9MEey7ZIXSljbwjtWrPYZWrd1hv36pXFspEn7MmQZ66AT/o48OiPU5k6GbUpK/CgyaZXJB4CnG0
aEvnK/uvURXES245H/g31wjxfmNsLQFxPI1mcJ+PO/h4JXvYBJhGJnGyhthUG1zOxjzEJ/iGI4oO
L+pgMXMwu+GzYfhTlFUTL/C397K3aUJdlrohUpqYJ9epyrS0HnmTHzd2w9xMw4Z4L1cdXhCMUgxl
DcULgXYVxlzxwXM3pu3CGbuVRC8a/cHZZvbe3Ts06Pq7P/Fb4g/xxbIpKrqwC1RarGZx6XGiGyUR
QUYfLvPQW3MkGXb+qhEXSH90zdJUFjM2hrYJJC3kV8aZzEWz+yZqUAKzgsYzMtk6j4xso1DzqCbF
rRXP2K8LC4CQDd4foAg+5sDx+JO2kHXr2b1f3SX05zE+J5szkeUBqeFssJrVNaVhLW5joaoCILHX
S2cYZYcCEL3Bc4PwAKwnABvhM2JgU2Ggdd5kC87qIhVnFMLnZtNddKSVyO7oMMrv1ONvXoXY10J9
WEGZxP0TZa6PKN1RdIcJGJ8TCw4ahbnqjqYK9W5W15GHmV5XhOZPR9OK5uovZjdupNVOoynTXKnQ
P/CH4A2hjlzQz+nU2nMoea9WmbNyk7gQ0nAI15cuxLIqhpzsSEeOwqyQX1eFCpnuVJCtADYnIRNf
gQq3kQTP3D8lxNu7SKEcaMmlplrcdi4O0Mqf0WMzmKwXizgU8pwvLuwiLah3eKT489fY12VYtt3f
rIa/M/VU0Jb5sYCX243PRqktmngvXWPv41ulj72dpTVXqAV0adr4MCbWWwDpFQJ5VsEkY5paxLuv
bM1zPXCOddE6VrWrqJuzLZvnaULJSnDszS+kLXjeUrTT+dtVjSr361oV+sJe2IBQzURJ1w77ZFeA
CU6iqhorktx2eUlv2KO2cI9uwyPz4sUheBXQesWSuTwC7O274ySLingfz8Xf0jr8i6J5o0fM/d4A
8jD++xF6q+YQLFBMONIfzkWm4dzUgCU0Sho1AFgBO6r4PrzwojHYS9ncGD389zbNITigF0YyLlwm
8TBks0CXIu6BoQ+EJcMjcyS7q/OP8kmk3RT50WtCSF5879MkiQbyCoXsOLNVkuxb7DJvOldnZY3v
cjk3QW8vv2KplrDWqzbhlNkzvjiPGwVqP9og0pw3vibDDWbWCaLF1eDLUShIK7MXcIhMwtDaEDrU
D47GOugE3Q1KWP7pwqyzfJcP/X3ykPVme/+BkTI8v9nJmIaEfhZ+TVu6xCdiJQmbuL3nxDaKcBuh
Wgwzb7abk6BKAjJoQjbxSzaeh4/ANpXyXyCGFDfSfM68i2ms/mZO7jB5ZFeKSLRwBvE3peEqdFKc
7rLkvHL1GPDOsyjZK5dUbPJBqRsNmaydhWAMxXR6fdbdWMfbJm+UjxlxbRkf+liIdS0hpxGd97xv
TeP9wnIVI5A5sAxPWC6HVGz9U9XJZD6NlzW2ckEhqK+/3tt3Zndl9fS+CkgJJ4NmZAkU02LPQKC3
dMEjWi25udMvX4Z46plNHojka+pgc8b4D8OlnAaRMmktOP77BC6jwE/J7SKtDXqFH20+ka5OBJNM
wuxHFxzC+Zp7HWFdQsJUgl1dx5Lv8fhDeTL0G6VnqKfhG+2p6EuIu3dOkMLqfk8mHkO5I3TDCpF8
wC740Ax+D4dGXauO/qdSy4Q1W4WpnoT9iPyii1qlE2dvgsOo/KvZb8km86fWQngJ1XZBwH/gtf2C
NNdIVgau7n0T7F0AXNBg8tWgc5152qKeevoI/Sb2oC+1hUCoYZIwNfvQjWWEcU5pU408eqiGpW50
8nPtot53sNdF7sByInWTZnNrDgi7wZzVcPvMMUPqzoqbYECSVEXLv3uF14an2CGNxFHjPbMyNwXk
InNeSGhFGR4iHN5zrhixIoKp5KIPx34ppnTA+rwC70MCZwswKnrP0kRMJivf7A14DyUkyruAGspV
eu1I76222LQb4fW4rP0UoyVOiqak/D0JN1Guo9zkJQaCnS7CsZy3LbW+/zVA3S0N9f5qSmD9HFXj
pc49hpYtclbYjtNPjLG83QknOQAWk2PdXyIKtLpvyuNpLDsJ9PimckS4MdcnmEVc89Eq1nNTJXkZ
+pkmQd4QlCVtNIbFMYvVgCO3VSN37iS/K3PqZjTvIpYBgGEHLVkyfaeUlVJT5jqeZQ6d7GH10zdG
NckH2fPLexgOUj6stCo66Ht1WurUnIBBDqhm7+QPi2GfdFJ2SpHBN80TMdLPLMiBuTkuMK0WulKB
j1AAsuxP/9NBPQuvVV+ePhev/bsPSTGVdgSyjKbCT91NQyOcPCeM27b7fneQt/vmt0Rw6Zx23X/1
vBU3+EdGZaNfPF6ewRKEz1yq3AJK0O6SEdSKU0OjLWm9/mRJA6dErt2li7fOr5jH3sjmtXApC31t
s8YAQAKwBHGVBBKq9htaMaQtOO8n606FdoisxCYn2szEswWAhn1NWgXgPQbULKiafn+VsUYovaeQ
fYMV7wgnIs0tkXXZJ8Jzn/+sRSc/bSGN8DXoBE0+F1joaMTDRomsFyJyRrjR80mHaISZ8x9PNxmI
yPwuNowpTCTap3X/do/MWuO9a1FDLa4F7hUwFYuj6fe9pOgdpr5RuLwe95Qdb7wXKaNgk9LCreYd
LuIZ3+IFMb6qwVerJb3rXnavtNeob8yag6cdVC12OPAE5X+IeQu47BbtXT7eYvZUNNbQEAC7xRus
wiw8gm0sRvA8iNm2vcoaNWT3i3IZN/YkDoYKmlE4u+xGGkiY4keMW7h0h1CyG2z1Dr3zqM00ybPT
/qaD3TNN+jwTzvxjri3mZ9bVRE2KJV+WWi1l0ttAfTvinUaO8XUs8ZInXkOdzng/hhMt+QSexsNa
28hR9Iix7PGWY61GLy4Om8p9aIOu0p/km4Utj7tk7Y6U+iPxrgFx114P78e3N8OwS7FpBtxYwdJQ
J8t5vIrQMOZiLww5CvCmX22kbPqAnAOnDZNsl4vaLCv5TTLrkcFiNVop9yfd9LrWOmfLfPKEE7Tm
ZYa7CGmtXjYVPGLXuXDdi49oQKv55q62sSljd+gMudQ7dTxCxW5aqWkEAyv1oL+D/Ourykuh09DD
rnb0zMsMyWw0hxqzpzp7Axd1zn7sEqQucHwcz5nZG29Vw6MgGGmZ9kmzFt7Ou+dcx4c1X8bYT4Ap
NVntUc2rpcE6bUot0fr7XYTUgQY6EpXxxYU5rVMLWJGxWNVqjGugYaNRYtoJSupaJ+xDAUtnsC5n
FvpUeGwL+xRd+2Isqf5axvdk4Tkw47DgziooOLRRR4aKjTpb49SXc6+S0KOzOeHHAJKNkAkfTLFi
mCEu0B1cAoNK+TCrA8ddtPWJ5mRc+Fg1uFBCXIgw2kqSZyFsIjaiCMLkWfIxoZYg7WAdud0Di0OJ
IINfI/FDu+8iksl4puhoXo27agmolZdZj4pCfC1ii2TY1qxOzm2Xmc4QOiGfbkEs4EdmmqaCQDMk
h6z7GfqJri5K1upYdSqCk32iB+gpkMCj2VOcdHow6xx79sMCueYSoOYvP4BxRFPSYKZjelf4GL3z
cmbylYbYrSuyDVwnZcUAH4ua1gxBPlpz8+lEdx3UxlTvf+LYE+rr9RD4iuYQ5NHbWBO68Z8ApBiz
WHaxX7h9QIhgkwelOJaOV7TkngN07ujdiy8x4VGFwNxCLjObMsxYZzqylDhKnAFuGGZRW9ncFNtd
Sd7uvLcSRwkTLx5TkAHyMAN1KP846sv73XbsLFZsednMLbZVXj9AuFEnm8nk0TMAKyTYhfZEHo/z
XihyriiU94xSC9Y18+c8tS/VyuBzuheYg3jMGDNctQKClLKgeIc6KrfSUmjDp5oGE1PP1IgMtNSJ
54CdU7t1GQe37DGQ8YzBE0HXMT9a53t1micvw3pphqsGeV0+qluAwViMHWWXEXrRk21krVzTIBND
79h2uHU0hhiQpawD/Vcb8i9AvUXvq2H/mcREvNpsPAj+3I4TU3WF+AD/FyxirVvc7H5KUmlYnd66
VUP3chtLjgdAEdYfas0po0USNw55mx6/Uwf+EpGa9ha4eLAAriZgYel139MzHrXSYLuzfiRk+3tm
TAgAxueotkfNdvX4H59/Hv7VtZXGWpags75vJThyZeHy6H/RdotgqS8bzW6dmZOjpt2wPHdrUDQQ
npCOJ/NOS9RK5wqcRoWKHB+VgsEZJaayToAc+b5S0Cqu6Xr601esFU8yJEnJa1KUkH+ZZwQWYMee
NszObHYpfWCjF29huUkCb2/EqdTMIEEJbGC3qVXHEH9Jt7gTsUVtsi25HzpkxmJzMRbZtnnMAXuR
7h1xfOm+F40zh+ISmv2o7cDxG6KnjgjTIvGvEZ27ZUa+axbCOkf/N2Kpkqw+wDJ7xvumjm2qM9sn
KSqWh+Gw2+mqOxTHix+Br9mcLg6JiLLqsK6DF+CZ4Bgyi+IBuhuTIq526I6A0oSLlOv2LKT8aH2r
vvTasehHGEDKnia5N58QkhalN02V+eCd7e85HWU2KQ/K8SxvqADFRvtyrMJXhiZlZ7h4FroZ82e8
K3Y362T2RZ4FYCpvzdSTjyOyjLvkSxhLUl4A/s1l7x7I3fpQDRpLO3jqnokodeeM95wyTKyJHyHc
61SNz1j/cjQGYPDxSXr8qvNKKlqw5X7ukpOLtjKvNtqpIPIibU3+e3qXyZQZ+5SpRiibteoGZ9Qs
kXYCcvIKdhITAl9Iy05ADTlB2tf3MyvWxBrO2UdDLhyE8IlPxXcjLYLsBlenS4wtD1aNpHGrjCx3
o+hEKa1leB2TaQS516gM6hv+z8nzh53dHrOVq7U433uEK8J9ht4aP9geJAN0oz6gkio+jw9Ek6ua
tHLOvHgsfXSHA8kFeOI8HoCMurYIFhY3B7AfdDq6TsZj/GUNMOKi/1fg131trd/Dr1xsB363ynB8
LGO+vR3iNobT9GF2qGVfR5HDQNfwvpwhYOeTpAqcCDfJX7lQ4HbNDMXGh8sNfM7kfKSTOypeTWBv
sTWK+z7WsmiH1w8ixofF+aLPWxVHxnr6JaEeL5sQ4zrLBLkRkDfe/VppzFI1NiZOVWYA9nW+2pRp
5OnoiUxGygPzqBbb4HPP48RCfqafnkAmjOUE0M3KeODu5loNjprjZ2vPoNFJP5yOru3TRx4ZzGI7
NerUF64fIIqcFF9qAGBNTpj0nKHgNvY2L+AMENm+g38PSlLAXCx5dtLxwq/XXjnIIB1bkcnc1Eho
rpRq45MXEzSIRA0LOxtAlfCT8AMlfhYV60rsE2WgQJPizcaaDNEKC7GQBcEGwnLqITlM9vK5SW8/
twHny9MBX+DE2KNrQot9w8G6xa6st//zo8sJPzBmKkGwiFGeRxkZsBr3wqntNu44uUme8vXf7FWc
amIFCKjMeD1F2fm4/3P3NJ4mtERU2RtRl/VUa5uIfYNNvtjp5ltjFq0+mfPQr4wIKVusDEnDW2eP
mn99WCr1hzNXxTiS05ursFzNO6RnWjfHKgNt0S16TcGx081K0KuM9D+KnbzczmPrpPPlPECk3rNt
NLsL/LxMUf6LE1/evKswwQGxhVisIkZ1ES0BI44+biCS3jdWLiSZ+qSLalMfrMlBsJM83wGEdzNd
u6Z2Zo++HPIzZwt9wrFP2ODMFaUuaqVMoraKkQnbwaG1dSjo9VytqYO+p7YjHmNUfpcrm5Ymia+s
eYX5Ump8OUNokXDoCFOAJLouXe2D0eCPq5+UW52lBTW4QlAcibH/tW31RxblAnBGxaLhprPX6LS6
fPCAmt04KwbPBOXzYD152zIQfNJt0Gn/7QebAqCZbUoEzuOCZrXRYfoVXq9Gvks7z2+/+GPOvG9U
5d1fk5KTvt4ZCgR80++lqDSF77XIspxQwxFvBe89ieRz47twzxYMUe95LQSfKRQVGYU/Z+lYw1Yp
xBOFlXv/7y2u0Tlrrhadpky6WupffiDrGgI+VD2LyK5hGBXQQwm6JNp9zwYoh5mwIWUuZaPgaHou
onIuS8dZngQCeq2Uxo7x+26aHzJMgzXgRBaxL/hbatdfPuMd0loIpP7gj7IbCfs5++HfEDEQDwfy
oqh2JoGrY116bZFINM/ojdJAqsJ5a6iUqHK+6axfq8b3T3DglmhEdFA2XN0AuLo71n9zGTLK95PT
5Z+zMRerBOYr44HFeHE1Ajb2fbyHdu9e4tUMfJ2eb84JHgvvpuei0yEoe3Vt3LGO8SaZprRWNSE4
Gxv6ds9SDA5WhMrVsYPnFIXUE7KahpxM1qc9WnARKg8PO8E/KyOD9W8nKet2xrLZ9K1em4q6aG98
kkK48GsTka9v+adcFx63Bv/UoUVwZlqmi4Xqhw890U6KajVj1o65Nt4SDmfqYp+BID9Y1RMjoQif
+I5munoYoj6ahOstojOHhvz+Ts+aR1kRnpu8sZSrbHPJtt03sUCNwl8ubjC0cALlWygwt0EVjhn+
ELZ0aJaD4yzisVse2HjKSufy/LxXcvIqrAsdnrz0bvjXxLeGqkSkV/8yq5V4PGSOArgD88m5kTKJ
Zv5p6igg8M/4TtsWz83D8Q8Ocpei+OiK5Da2diYIclD4UHDppgelWovKHbGV+1yo6zIjAMGu/f6B
9ylYIPQ0Wdmq2wScXYxO70DyO9lpuqr2SaEbu5oM9xlcoBLhA9T76VJVmHy67HQkt2c3gEb8WIeR
cVLx7zd3/kgfWoX4SMPFN3F7uoAmTPuwpDkzBqDFuf94qsC96MQ8PaeQfCaOwuN5NCdVvIZQ5c2E
vuUM9MHAaWJjDr+WCiuQNWMXDgw/g0mqAuttBZ5sFh6zUXFkh3cDjo5OdfuauyHHp4Brj1bzarrQ
BnzWXTq5Wse9Sr+UX/4/ZulK0c1u0undADxoJher3sZWzHDnk5XOJ33wsKuqRHOnad8W5FH76CGn
atPooCREoX+ydxtx5XSf/DpdNJZVNJauBUeJRYQagr5fyEQeTxHYrrS+y4AUtjni6Re2RGMfpevz
+okvzIrgEcnmLAjqI3e+ihGAUcSKk0YjbddcVu9QaXULSic3qIuga09OWmbIar0TrylXAUnxd14W
UfdjxDFTl/1lK2OeKthECyrbAChxlz59p2lKM7ctYzFfBhlqgYfIUk7Fl3EbZTfYgWE+x5GDBjnG
uhHzqqxLuQzaBmt73qlQejJHepGyHcceBVq35Y1w7sSuA/W8yrKetLagHFDhIoOfv4tWmfspCbyk
DUvdPx4UGiwfJuQIl4Coe5zZohV0ODyGFJ9hcJ2ZxVvvqSYBam0yc1tX2Uw5ccfj694b62wUqdRz
dY0uU1KX7k/kcIpZrhs8xqcN2br9V9RJ/suM2PdEO2NucPSxJAlSGbFPBmEtB2YrZDqwBvsvBdAs
1LzJrA4KzZFz5aiRzRkPrLkceeGh8BMzfjMe2I09Deugzl1Bszzj7mC9XuXOiqb5IWA1Hm/aSCbE
BOo6rb6SprDXOVO65GrpcmsoqRJWN99CvcQH7hJBnM3xXpoX1w0lESEVzJXMG/P/pLkSPHaX6qzH
sFAF8mSE/YTgCB2hQf20mcRC8E4SVjSfCcH5wqklCu3vHMR9TsoicSy0K1VXIbMloTUt6aNgjuUj
yTTcyJmcr9CrN5+2kj+kd3Ed78AM01Y51P5i0fX6QnGnlTVMY6d3mHvS0GpdLs2kVdeTApUO8zOx
zk2uNatX9EGUSHL6CHBBz7uhWkPxjAr3ZchFB1p2IMY8TYdsmohtQv0DzFjSOGMlrAFg8B5NbiAp
BKSFM5LtztEMlRTE+NqZymRjQbjwP/SybFFhPIrSMktRxY4eh5DgY7jaIK2SkSpg7Ev2Y1o3hYi4
Xaokb7RKvdfmKR1WECgkW7DD0S+XGRhUsNnrYyoYJ2lpyKWrLHUNg2OAglbqG2m1WBjdOhLtodQr
gobK2ZfZrziUEtjy24p1A/jimWTBOV1p+qOT7fHbVMRnY/fBlVthR8LmafFF5IufJDtJRFkqqJWX
3jXViP6Wxpr/hcrrVfoH8ij3f8cPEy+OaAkdfgJwRs9MYmoF7cczq5c243n4fmrL+3EtqH2l8cQN
a1NACzWbv31dwvxz1Smrabi1EH1EykesDF/dv32hlBjJaDqsNdJwDwARAxZS8UlHd3Y2TR1OjFsR
dTTjC7pq7E74n2gmMuurOQySct5k8msLjk/XpDpvg7Q+VY8j6B8BfbikfEKVJSQ9VjPW9JJyuVLD
QflD8t5pFL13Zul6i9zFcRE6lYEIUtL12daocg2xm6kDg/cM70CYT+HVoTDTx26ux/OaVaFIpzMh
doqIn4hF/gRDikxuUYmXAgtBn8Lpav7XHj0fI8NmqMSs14AxePL8yXQtiA9H2K5aoBeyFderogse
1lm8DGVkRRbMusEPfs9sMsar3T57s/gz8HqQxtqLBRGmrh1JQvP1n4P+C4d/yr4pQKFBkjc6PAJD
fXuznDxfy+ti8xX9JxQFPGkO7Og+ldwVONGMFv8bJ+S8XAw1XNCUDPxPoBMvtXxGig1qhy5k6pSg
7alwCJDdWqVD7rL1FKmdhDh1WElBVQSu+ltD3NzYd5VG1RFMsu/FhX5oXwx91ac3j5PD/kKyOXfc
zAx3YgR4tX7BHtHrctK/0Hk4DB90JS+cSbb4uyExNlpB5HVCnekLybSN/rVfOXHYWag2VayrjK/K
7GwREsBOaXFwxqIBc7HZyYqrI0ZAfbc97qJx7BBCFSJq4HgXXkb8hnUb4P/zpBXbDCKsKmhOC4qx
bdatpR/y/ZLTg7Zg1jqT5HeAYmrQlQLprQCCTp8ydc5o0H1H0ZMwa4FYel1kbKp6NT9TyRmdVXWH
G1vsK1JAmrXcbF+5X7Tty6r0+gaPexWAdYENRdbtoGCDcjzXq2CjIuTOwMw7URCtHn2HDnVtkdCZ
M9Phq6RWhaJ2it4utdWBxabc3FUHk464glYPtBd3QbL4erazwn7U8AeHIGUyzCPqAzdEhdblSskU
oiOecoe/4zZ2CcRQg7Gw2Of4J61lS336YflZ6UaRV9Jrf9856BHlELsf51eCa+hXoeCBtW/csqmP
fXn4ZH1tmGMJ85simeq5G60CWGsI9UKy448vJGo+5kAEGHNcQmBDI0biNyX1hp7vk7DkRazDJRrn
ls7iMthA0B3w7JB1gNZxkit21MNWPBfBD6TcVuO56dEqjBygxNTxp9zxUp4nlrwOHwNPBsn0yEOR
tR5I8CEIUaEXi5LPz4z/+l0TKmYBWILagpH8POfsguQ2dgdlCcyhT3HHTiIRIvAVoagIZzXS7WJ7
3MR6I2TIbfYL5vVw1PX54YSYop9s07YvCSfaB1xb91yPG6Xq/SXzW8R2l4+5Au7KoolwiMVbfKiC
5U9CGXCjyY14l1zenJHyANtpfxRVNEQRATg5A2kqWRhJrOAukYAvJiDZlAhzWD5dv9hxHpsgqbPC
Yb0HT2iy+0RfCLtWxmeAzLMlj4yssqytNaqJzV63mAej6wNgoSsoa/DguWNRdh/0DvEArOANI8Vn
KCLx4j9WMGT4f/s9hVq3VtxnQNhPPacjQ7dMOlQIPgDr2WtzRCjuvax99Qz5eIFn4noaxNewplCx
42lnXYgj5GygrJ5nGzla5/ppAge1ZbJ3W6LTVkQ2OJBO6oQzYSkm+RMxx4fK0sZ4tE5m1KAqjHfs
kKDw0+MK9VFiCUP/iwBIdd83PYUtO5tlFm1uDvJJK33qD3GdYVuuKmWvCM3Sfpmem7qeeuiNMdK0
gjELXYyr+RXi3cuybbEEqwb01cyarcoieUiNERFEF9u2DPvNRcZXzPKixQOElTw3uebx+PBkwSD+
DdezznbV7iFuq6g3GJhCJSG29FrMy+vhpj9cqBgQcQZCvC4QLKXdCV18nTsZd/hxsgL25NEI9nUc
BLaUMOdwO9ruKNH6h+XojeyT2LjGlmpxw40m60AJHaWJc7vQByDWXD0+PJNdoQMzrdKQTn11z6jG
bsD5TXWSuX018fleffuqaY58MCrAzxDBvy5l9iC2Gp0z2oyGLLnSsFVUZosDoVziO5CFyiY2bqQG
SDhIoqA7An1HdL8G8Zm3eM2hkjs55z0BUVq3maQ4PlL0pCIrtEH4zZIEZbtyn+PB2H2PELl2BO/P
Jorm9g+o/uzq3ckPVAOasUoPtmNE9WZn169J/lEF9cwDgkEIA5A8e//qt1qXbNC5r2tvpFIAgQGS
8ep1dRV0hOde/sXkztbx+56YJ+/HQTziAipjOtYijbdfrs1W79xyMEsB5FfqWVPD47M+nzhsmhIU
86RBcfsZoNizawI5NqiHmmaSn4AvGd4pzikvhSRSabSQadwBrgFgXsvruqy0St3ya+hYvkpSF/Y4
7xrG7ENQGWrjxo7GcEGOgjZ0Yl+ysRzB6M/uwu0oDbeYts9S31VrGwaKRy3M/j/8aoIae+og5+xo
lpOW6njwDUYF6oH0yYQ/e1a2fFuoaLG8+9w4JBUbL712K3aFobqB8MQz9GjnBBaI4jjqhmm0Iumw
dTjTFKORXOcGILPyqTqrc1elr5eH1V8k+HhnB924jHZulVW9k2H84GiyxuMi2aGLmcm92Xx8U1Jb
9TttoaDIXah6qbraz7C3fk8ScaiWPgb2i0HQOkSbcNWXylsI6ILg+bIBH99kq7ZK3VdizfII165e
jROaZqtydYhrmpuGIvz8TnCRILnWU5YsVBHfwxQ9jo3F1Wx2rCjz1QKjPjOmSnUU1cyRks0fn24Q
9wu/EkDRW6qACnqd4DwV5vC6P5bNm0PQyjgjfeLjdVBlx0ZLaCHHud+n/KDZ6mr9oH1nrX9o6khF
DgdKaAL+Z7RlUCD+c6VaaPuyVuiV5Qxfz/+blnzEEY1pSiqvz5c5I8UhMS2cIhQxPrXpZ3X+ua+j
SfdJCQR3cT57389Mmyht7xhuBOjVmYgvQSD12QDH9MO/Xd2DqlrS0wS360X4DlAbossBj0upyWOc
1nmsp1TbwFhqLSZ/3on7eXxnmI1BeBLzILzhFfjVprVXj/fGbMz/NvqREPX4qBPr4dLuYBC7YVxM
KTZL7CKIBszDsQPab/Liw2P6duFW3SJdfzKblS9tKp99fNQW9HoDdHy3wTTcUWi11325LyTcvFbA
1a3EsXHwuhBoSwTbvJxhwhiIBm7qWlPjPyAO/3wHvO7fSt5GxtYBOkYebXrZIqzCIdNfyxm2mmnx
aViOONl3YXw5WknAsDgHRDavU/QG4WwFbmETCjxBPImuHhsBqQReXeQWWHENJzCSdVJNc4B4SyDh
RL5kb1ub6itjrtaduV77V/PocPjbxA76m6oORue7kzIN5TvNzb6mk29cEHeRRky2zOdt3KHcELxf
WuVWV+ceSF2n92B9Yv7q7PZ7SoL6gvRZueKnNAQdQrS3RNnvtwCWFKRupwXmyhDhmGwVxUEWqgkI
GfCRpi4gyApAjSeDA6tohUPv47JWyocgdFlMcVWAH+M98jI/qzy1fBzknRmVs3UNIBQmd/gBp9Oo
j69LtC6TjcCpt0Oa5LhHJbZj03V7I5VoFnmKt/gTU86DrFEj6g20lmCO2do1WjRWTbTEU8oo2f+m
4rQ8ja6+VpKpf0BJTZfnzxw/X2GEN/44aXz7gWq/2CH0KAOA6U6qvwKrOzB7pO8RA+Ds0n/6UdgL
p3LmAA3GsaeHEbHi8Y5JqqgfkoVccqXHPnNB4Fc2FJygstjM/8DLED4n4dzZLsHKRerod9TP/WJf
RYDMZRU3ljTimprfIwiaYjkgvVPuKkAuczb1MnP3QPHTRdGm+6x+IlLYl3z8IfdE+ccvTu4y9Rc3
s9VLv5IBKtSQg1dhPz/HKXvvw9Me6fIKWsZvdloE4szfLx9pfS6y4TBntbOZq5B/tGkCwd+XuctN
jZjXgg63+MgY9M4sySfTR67Eoha9KboGT3WV0XEcqJvtRptpA2rgNDN0AY9OpbDvXNx1jg0AoABZ
IYHIKTIzr9sX8J8qhnTyXEqPNockNZTtqROKPUTLu6+5q1d0VshZ12gMhnNQXi/omUG0sGpum0S1
jinN9Eh0YPdm5fGw3AvgSuluX/+7fQ2u6vRCYhOXdXYJnrWl68zdJyg7WRlYR8q64ZPClV9kT+th
jp/SwW74fgXnzI7q7/ykWBvkv5BI+YhIBDXqnmToCfbhs/7TPYgTv+2LBw2u8oHSMi0wcIlhCq61
omvUvWPEvNMbJXCUyV54L+AkP9fmYMyaIrzzZiZ+cbEI4qD81cZpE+tIVXiECgIm+IpzK6E/fjdV
+xVN6fDZkJySRNjVBMDO86903X1vghE56oq2EDKozRuyc4zs2naKLFAuUj4wh2kjsvOvDxRnDnly
cWaVfxkiCjuQmMwlmG66itNeMpw9oZPBy4t2PP2bymvEwYdXPOH93sv+5gSFM40UAsoviva8ssc9
wqYNdRlur2QhfFYnlAp8GQ+W5g2fYuXDOTYAr1Q7JUn38FmmybCDxkVbJVwFtJxdQmUCMyfsA2LN
lRRvlIJmiy1CCkcdGZgbUBBCIYeuQg7qG0YJ6nDH2bi1qAziKzENB4Zv3j0DXn7RkAuw9wVJpMvi
sUdE3j9Q73m9gO1SqDUiKUYC2Y/GJFcltH0X2PhlKTo10z8KJOHcFYXyyYfXa4GCqUEHiYhpnzQx
y7sDKg1zTATResJQKG4DVWKroQ7DCAWQtgG1sUi90M4HESy7WT/VnaQIz77z3Y5unG3wwE0QPSHV
YKJETGgzVSaUDhhAVSW6mnPOdV1jMYjqEGLhJHEe6YlNr17JN3IlmfZC5Jg4A1QiRZCWSHQyoun5
D6tt/xMrziG01hhd8JuY2ERP9hDFDf5K6xbZ4w32dQK3vjCzsBbzdzg48cfCamqAdNes3grpTRGj
Z2RbjAyn3v4FIH1OOgKvUVWsq7sRTSjW7cMLP3awf5XBAxuTktyYQ6y7u1vQua14CUHvv4UyqR+o
5pYquQl1RsmNYlB2XpS/Fb6GpPBHV94wey1KWWa5Z42PS2h/JTAZO1XI7IVjlHNwd2/EiqNw0nfN
BrDc3exoBIhbeyNHCsetjcBWzR0ZAdNNlRfI5Ms9X/AuDQqGgq6XOFhM+RCfIibnY0XFdfB+GpeX
MqRVfXbA8WLE7O7nFcunzTUfiJ+38UPgYlsSLA2H0UV1FKD7s9Hlz7JkYwZ2EZFr3hH2fP8E19Vw
07r3mPiLyXxjvk+wGTIZQdXmzlV7ABXP8ZOda2LltbdmJ9Ym35tFpStcAr3TZWvU0eZCpkm1o5wN
wU7qT7k8i1QPnMnE2OyhSWz8lu03v4Ik5paLLPPpS6a1j7apfmaif90rGw2HtOqZq8lZwPLa+OhW
Rz1oD1TwfIos7QkBCvhpj5UqIiV/gpMbmodJvmWHtc9xyKw4GWlplW/Q2K5wAtqn8awPlg88c47U
Hjz9bBnXYhMeovj0MpbvEfG0Ba8kxigFs7gDJ+K3nBrBhPH3aUxv5PP9cooBl4grZ8JfkgLOs9VH
t6RGB4tBFeDcbI8M82HmvUoObk7kLvLXngEgtcgPAwUWt9geyHl0t6ZGbb6z/J51en+z20+I933f
Y5+Ej7YlKNc+Mo/42Tyic9m9+Urz+MpInTzMa9otROPrlwr90N58Me9Ea/xSwSdFgKRGHlx5EI9y
fedPw7xSAOMP+3s7dEkEJNO2kyhirGkPtYGkHHen6/180HauAYfHIR/wQxoA4YCwST62RvzQE7kM
HlifvELsz6bsBYG5kZWBsF2eoKkxwkaeBryaAg/+9kgDHW3sEudK25oUM7KXJ00JUYr5N6h22wSl
F4PjWzmBkUg7DRBDt2xTBIHvI0UYs+G9lWV1Hy+vo8CwNOKXJx1UQT+HFZnAcoFf06h6r051JQOg
DfdvaTMsR97bDc3vJmEvF9Q0AG8rY+f7Q+9HQ2a/4nYyzPtUGTeKZIAAW2j+0zmj6ph7yRoV56/e
S97iUhnVU/eYy54B/jefYcdAhiiGRjhQX6xFzvhltLHCQkGakURAf2Lg9Bi3I5lmMeRsEHHrHRcM
q4y87wd+uaDEmqB91gfaAxplYYpNvXJFBxbqfe/RC6wbpoAXwa8IkCScZPZhBrdNqPX9xN5yZsV3
yL30mKDC86D2VRbvv9v7fYevT20q94YEXKKGYPjDyBeqh5R/7/4PRpjX3oOYvsgXi03mLmTMbu3W
0nCB5TC4d1HmWTRLhgDcMYsuQFWMYscNikvpubdO1rpNC4pMiKu2L7t4gVbMAsxQJstTQXMQPJA5
PRl+85GxazZn+b5TCAUX8hJixvYD4iFAFb882isWv9PRr/4MiQXbks8otVmv2iL7DiRUxfxyrNt7
32jBUqzDeltxgEh23JtXmeAeMvCN2m0KLG1n3Ae53vppgDrWNwgJEZW+tj/8ph/kn7fuUKg53Ozz
zGBT4wPOTNGpHsQPknyBu1PVGpF3EYLqJyFRx9alkSfUOw1nAJ4ybcl0a76aQBSa1BFjPqDHTpUO
uj7ajhmZzDc40yveHDqcL3cwKaL3a5xJKQXA7kGbttK2SEI85SwkpIJu+FIRmbIj+lfxZGIXPtHD
u3sfysESD7T/YyKkXqiC198HGRhsl619SefthL/MJDbBSOSsGo81AxCpG6e9LJ0ms9/kGyMMJNx3
ykcFnfAnfF7dLUsGxd2Ebc7Ls47X3c4phlokPGSWKYUTK8RVYNw6OwaNofw8SNQtEqwHOG0XQ+yG
1Wlorrm8/BTx02Z8ZV9Rs740VnYflya38Do5wFg/0C0CR50y653EAJVSLePklryRXYEc0C+NRWD9
fMwYabEds33zrkwvlDMo5F8Fjsc52Z0vyU92A95FQWOCmoEcMW+dWZeRAzvGCb8FH+3M+F8MtrF1
7frZOjcFkuo8CpJ10VK/kwr+oaEm70ubrC1sF251Bhkax127puFR/D/c1MIWe2nAKT3fHVZ+G8hQ
JoBPXfCOKrBqKcvZzTwS7zFSYIvFQXbUhyk8EylgQR/OHZtqXnGtRFqNsvXJAmPsbGVz3quzgXxg
SV8b8GDLM6VjBIk7BW3eRNrET/FzzWEpbL4KZx+zppTrVMOEiA9KRpFQVIOxGOmT/EQXJc1P9P7E
MciQAdbE25ErFZ5kIYtMjtPoK0hZk4L1hnxk9QtOFEL0NJhQ9zVOFpGGbD44XmAQgu2G6MHfwrzd
GlcYW35EG/Xy30sYxuaDHlYTtBpNls1BxJYbe0PWuR0Zn2QpKgjQviz++FGZl5LlfG9suf5kV+kW
zzsdZ4lCoSkMhlHoE4Pmo0vXl2RcOW0eJaVMDO0yY/mfrnjp5FYErtQsxdI8v7rKXd9h6iBl5W7q
3X3XQY5znAUEfIyp/wZMSZFqdQ3db+Zn07TEgyVXA1eYyXYKYh3ZyhleKdvDKAVYjTkizX4hWwr5
LteGAAVIo+Fwt/uaFoEk4UwfeRh4idw9ekvQVG1VaAlDnDB5KI8HOmHq3syreUn3Zse3d5bU7qll
cKpQRPLv//sdNXgOkYGwb54Vyz77BMkbHJaHyQqXj1o0D1d0/3f+0sZuuYh66Pqrj0TnQe5EX6rZ
L19eotQTocVrITiqSXcPUnSmTsUcnQKubLtazDWI0hxKipns2LdLK9yqn8RPlfHE2UgU3cce6cUv
7zKGeinDn1jzlXoXca0KeQtRnQOsuDfOynx4EcLR+96YuUa4NTKLtolrCleq3R5APj+6htjRUFCY
92bPwmUrt4OWhDT9ukcqdo8R3gViF1GW7lSVdm37sImIavh4bzCORbkfkxfzPigqs+LZQ2Md4zC2
H5XeVl0itXD3khRDBwj3izUjsSFctcre+KhGpC2JKOXr4wXB/ElpFpDc67DbBO/O64vM8lu+/O1D
HvthN6ynsrgPKNbiMgnmUG69nYk9IiBHPOKkpJ/E7/xxM5QNG/mYeABIy0GHds7TxkCRC+0wfQEU
0ypO7zABpz6DZP5oKbLglLIRNb2D0JdA/QylJ07jowkGKqFHqNFQkI4oo9w3lRoPb+fJtUVpa1g1
S/kimTCmrqrMXx4dHGERHGtwhfXxcGiTKnDj1eBlxbh9+j2A1YYbfcHKI5pSxD42v2lzfmPcfsML
zNYwv937eFaFSOFYGRALygI47334dNIW4L9LJAlhElF81TiPIK00+N0hWWuXW+7TmOFwd1pgCUFv
iljd6ZS8VIa07R9ur/KsmVvzD3ZEawwMq2huya1awc5QdjjfgQoaAsFPfNM3NWao4rJTH6BhYmwf
veno5C0DMv87pk+Hl3qnZbBxYovzDJu6UTJAPna71SAypi4M+f5EPLTfpcno6OGwuRroWCyURMEH
KG52tYtWJpNmUSuhCgFw+Hi7Q2D773PMrgVfRTRgKy6amlE21q3zPj5USdWOGIlAATtPybl9SB8v
S9J0PueOacCGthMENc+hwKxuH3Z3FJRKc6wkye2eq9IcVySI3ZLm9LE6GAmnKqV1CrRPsSiyMpfF
6i14/1CDQdbCyYT/ZkumX31ILF5EhAz2kp+3itz+AH4LoeLqYMEOtnnrW4lfQymLXE2IaM6/Tsj6
h6ymU0BpMBFfIf4rY7iZ6zfMdw+/Lka7GsuOBBQvW10twTzBDD1M3BDC5oF+DDWcrTIoBJmGxvTU
1M7ZiQURICTNXJv5WpPaWBt6ZjQdXSY5xWssQ05jgsQr+RZ7tlKz7wy+WWxc5T2a6dToUaVQoBXB
gQzs3KxWuX4pgohe83g+e/X0ynbHiBand1GHdVDPR83icjIMiF/oqhodG9V05kL/s6Xn7uKbhsXO
bIzTGxkmfmJ2pvV5VATMt03YNP7ssQfVZWE73NEM+sOwD/VF7kHt0q1FAz7Gkc6ymc9wZ6x/GPqF
OdFDMKhr56+atuq/wAY3ZxwnduscspkJ2ANSmnUb4gr+Sd7c63PgD5Y33YuKxeCm0f3H9Gn1RRpk
RrVLGTctq8TnA6+parsaNAK+UaQsbjILuKSRNrq7dX4xIPRUoQPy17Uf33cohvjawJ8eI/zJo2Cm
BL0PXNVrzpehJ7QWmNFV41uyYz4UynGv7zpFoc/DA1EeUOxIvVNlnJUA8YXzYePItWdNHGO1gKeI
0MBYGqkteGNKeJ7MlXSTNPy2hkfVjfkw6hkXTxkidJwByD66Jp6IeQwSPQrs0CkRl8GdVZASYcrZ
UoGX4NBZNXhdk5uK9VW+q7R4HAIZpW7X/kKsHN9tIxYz3L8lVHdHc4gMjcl33d91Z2UHjEBnmSh6
bzGqBfR6le6NDomulW8H6gi99CxGqPWgA3nV9WZduq02Za6ox7YabcK2TU0l7s2Cs7bDchcHnop9
pgpK9+y/lpFmG+meqb3RvIZtRKJD9uvQXR3LbS8qCKmXFIHbY3B3dED3QpjuEEzmpnEPBMEmQx4I
fWO4lfjkGAIHHpk95pj62Wb0cOk+IfJ1qUDwtwenpHA2HnDxlPyoIidA6DXxeAXZNJB9LQbKPRle
VHr24pVNqNMF1/3CSEwd8UC0q6rjiwftqCGiNEeZxrcX5HD44+3rg5WFPgRQ8F5gVmOQ81UITTSy
eFx/o8BlFk3SQuBblmsDHh/09UwyDoitmQgD/pB7iCI9f08z7fCarUMRR+pYSAq4F2Vtwxt+uqS4
0jS2KAC0krpoK1K174N6XCQFgHuv3KzaUrr5h6zF5QKy/OctiIwsZ31vjJ8G20IRRR7TpH1miuNK
Pwnl3uCP3s7M0Sb+OvyOjiz8/jlxNIAtg3NRP0xCx+rP2XLfuESTe6dREpoLi6s+7qf9Zjuy7u+p
T+rRRZ5inYpL2a1tPxRW0/4CEdIbLWVyICuhkngUwFmptwzCfoRUfFbdCv9E3mveSSqGh3PF/SF+
JUoKRupjsHP2v3vnoB4QdqV14wD2Ll0N9WoLBeENCuapEdhTuMQauCkssKFqfipC7PDwt28YjHFJ
fKSvWajWpqVbECaZ4pQIWyVuFeqQK+xMSQJcKzAS7YmlmWCs5dtS167nJBNx1OypmbV2OxJin5pG
RMUN4BAUCW5RXIAK4rC94pvdZMsNQP5zsm8f4tzATOz5/l/cLVTDq10XmkNNl1u+8DmRB5WW1tiQ
eo+ac0pLwZ67AT/JlGVCsb+2GRODzOioIheE95w75U+5hIrz7kATH1mmLYFrDb5oa2TWqehOvk9x
BsX8mAPP5KjIZDAVvL50PILqjv+5qWlUyoKYPluJoDTxUVmJ4+8T7+kDTkD3j1DWhK4hZAvlDFUa
T6N8Slnucl0TvaiXByuIrNAyu+hP6XpCKGiShPrTbz2PjaokLtrrH7EYRUgZqMAUCVviwwAfC/bV
H/14T8kKByYuYnTCe1jfV7aQrcuC4E6p3VGpYF1rT//dN1630XUgI7hwooBl5l7fDVqIq9B3vU/P
t01PC1gu/X4V9cMxC5l6iCN5ZumAY92HpCbHEbZy96bSkRVMd5Wgmca1jV1eYmnpF6UJetERRKPN
Bz3rfxUPWwKLoLyqyVLLO8AGG2R6kVR6GEx6tS45ehrEfyewKIDtdWko5AqD199MILIcP/SwuGmS
eHDrPY67F5iP7MCfRrCZt5SRXaY5h8D8as5ePGMX1EekZCw0Ry4bYuw5rsbxM6puwgM1/aejnRqt
VDZE963E9k9/WUpGwFP4QMnjwXPVfSlxPWiJDI1k+ll5Ue7JZEbXVAxZleV4MV3vSx8kqZlfVzPX
jj9rqGfaBfvyQw7G8Aawcwate+Kbc6pP+oeao8HlpuTN7hC/EtN54qCzX6sCPF9n+a/qcDcRmkHt
OlcLKhiuLxjfjAtrChPwqqdEnTacPI2abw8t9QZtPwZJdO7qNY/6SZS6ej/017SHmhiMMwN4RAQC
TF51vd+6GQAy0OIuyArH2DL6rbf7CVxpaRzYeUvE0/MXiAiqr17hpsU9Cjo3TEjM22/ZHlD/pneT
6uT+YSqtHs168/dgSYa0czCmHfOUJkh8deDiw1UzIo3+3/KnpLwcD5Pb0M2Z9cbcSZpdOR9O6s5r
FggXYUTj539BxDYm1IOAVb0O5HQnQTVJhOJSzmq35FL6UPRcjf2xxYpJdKnE0e6fJhxsdxasmBUl
VzdXR+LnE5OrYgVFJzrsOqdTdLYrYIMcKpjeHhetpUHIGOBPo1D7Hu13Mvu3wcbTkvPvFMaKJe7o
2NWBu0mb6+U96QuRFNo04lHY9Eo7xOnRAMRv4HM9SPPtEimAqbNyqqx+kn8KPgKFiMRntS6O2eo3
ve2sr0vSFVjxcTrlT+mMI3W8xN1kWYyAFKXQRSChG1bmzTAcDRxOwoocp82WFyL70ambHQDVaoFf
UAonsJj4hEm/5JNyW+H4psbp+KH1+r1YYs1r18w+nVvhUPjrIa6kT7eEQkV+qR1xHs5WFm5Y13Hm
yQVJbM5F68A4/IUU2pK/9iYTG58Al28vVmq+MxyfV4UASsCC3OI/2iRLwRl6Q/ZxJhWAT6RB9gV9
Xen1TBEUD6bstq7Rs2LJ8lwPzi2eh6jxvdxSf/NweQGv3gdtMwm9mUmOU+dgOnw2MTAx0t2sqL85
HCRilRNP03YR4G/YBxUm3lPA8Ic0qK9beczvvkzUbrgDJdBsa5aFGQaDucJqek4bNbs8ILzjHzKu
ZT7kijKZwz5jN6JrlKO/FkLLacAxwvB1ibf6d4Ovkv9jXfieUwMELxzwXgaCPhMBhgSTT0Nf3sYF
/0H3CYeg9OjgFacwazYeZJwSb/+WvroZmeSmi1GAGJRuMLJBvezeSoWQS57q6Oz7wHW3nmkVezRi
wlZ33j25QVVV/O1loHi3yFSEJUe7gD/yuXkkkIFSjFp35tv5azIn6G//4KInrM79Ys6iC93qFcN0
XXZwfV5WYDmA8Ut11GFBsfXmspAtKOR2vZanPbDdKSKD3Twa5BECOdpEimuwqIaMO2kJvRWBos9U
asyj84ngOGKYnI3LRMNKgOEiOpLWpthw6Gp/dPIwgA7eFxnpyQ+WHWDv1NM/t8hmcZGHUF1m8gQA
VTaLg/hQWpdFWiLTVLucl3378qfStoVbvTv03apOU9HVBDMpw0KPughv894d/FEHl8ejYvQUrPU2
T/GanKH3ktS+AiCgwPTGsIUpLI1M7H1hlLI8r6qgoBJmJHzsmPtaYZWV9jx/arMI4tRbu2HLsfqb
kbsbdqT3vic/p0U1U0fIDfFt7RbBhSE3PZAV+h6cdXuIJcdY5vXjYINVw32M5R/QGiuaU6Bnt08T
lpqUQjg4GfjU0K11BIWPJp6dUQeFRU3p14FqAe9lnCiu0QsqA4wT+hwzv5TwXNaHHd96jRLgelES
T6p9aAl45hClSgEr3vHc9A72GywZ1ihhK8J17HnHsnnQFm2NdXPRBRea5voRC6kUaeNUE8MpZZdt
Ujxj9GMPUAZxQiN1ZWmkfUssmm7gY6+ZX0FVa3ue7HE75nSW6JyxQw2pP81OZSWs6gebeoP6ye3y
dIKS9IBIsRjNG/BUzUXOol89d8ezCvDRbY2mIRoZmkHoy5ekmsbGJhLOvVfvOVl+x2Nbin22a8Ip
6wffgIQ1lEHo1M+P7lSULQN1BJ8j6cuS/2MC09sX1ea6Jv7RgSdpRThP9/yH13FxvzdcsNt1fLOh
6SPpICJIW5fKbw/77x/4LxkMBh0ONyle56uePH0OOAZ9FjDxPGE6VmXTPMqwAo7xbX79JSGZWRi5
topldunkW6VOp8m8Exnga9IeQfy0ZdsJtQlzdZ4TGP906rSdk3CkDruhTdK5Ib99JeyGV8i++jRR
bz98KWwT8XA8EjfTCxLwKNDlxRsh0ThZMGjU4SoKAZGAsbwAK3eNeOEgwOA904Ujutnawd1YJsDZ
1uozym7Ly9xSGajKmcET2lVb9OrjM/v5OjZHT2+tD9GX9OD7p4e1ucw416K3YXy5qwL6KA6Q2G9V
jYuvkyHkMCeCSvE41MhhQO/0QuMt1O1KNkjLrLa4vJojDrUO/x+rQVWv09VFi5jzrnOH1nliKpgm
ELESFbJUr3kVNeLPk1do8/a/D/P2MM/6pEHFokbeY3gw8aZ1q8oQPKvfiIsDrL7EhXtgn1j7alP7
7dX883CaA+TYiGUXQwDLJyScXPqEXdbkhnNAlftYQOhHMP18glSjJ5oOpTjtUrBPDIk1nH2IJKiN
3DY74/6IYab9hUmTkpK5w15/dzpej4zKbiFOIrfwDQtdHB4ZPvrWr0TZT/Ll8OQ+o41BsA6fFdPE
dpxlYx4hsIjYkZPNsH1N72vc78zn+d82L4NiDhtcEw9Pf8L2gX6paaf1L5VKkYaHYOXH0ia+hdlW
iD0gGKRQFv27d0Mt0bYLB2MPehocsbVMslTmupOFKcvWoxvyN1JSkwipAeYQlTvdBlpAm1swedDT
jZfbjSgqVlto++QwIXh3n7LnGs9h27d+GP6VNfDQv6TvsLgN5PijNkq+raFTw4slXXxwTiOS2BIT
LOmLYyZp+NOS9kpQtZpxVpv4f92S3ljkGu/+NR8UcN7Pf2gMYI8UhclxMgVFkjZhUrfANvAYYb/u
QA8Wf5wSu7t5gpzWdPnmBeSr5J7Zd4OOPERZcC+BYz4sk46kb8r8XJVJQOikN2+zxRcRtoVefQMZ
UKGzpkCStM/Uz6CrOSISU2JWnl8CFB7YuSvajRYcWGsNppxcsQHbN5wB8icFL6hxbumm2a5+vuVu
iHvabceCSyklurEphwgvCqljmCMveb4cY09dlBk8mbUOjdnlHLh1zoyhGIF0tnE6Au9I9uG/mgzq
IiFjVfjr9joTdMsNMojOd/MvWb3mw6mo9cxuMEQHV91poW+j8SvDA9qex77F9l5OmA/zNfN3YS1y
R4GJF2K+CRncBR4Xp76bHhgTM3E4W4qmgsMSoVMxGZ4oYYzMMyjZ7jKbHj9u5VXKXPbyHVR18VlH
9D9GUcvcogeIEfkvJM4M3TS8/Py2qqdhgXheg+c/gIdPLqluUpmPvGU0JRl4AWXdyfUZctqVebLh
CSM2ru7Byl1DPtQ4zVA8fKaYlnuVFCVA05KNE+R/SoqCdDVbiDZdwxFDiYWN0v1xqzAamKlpx6U7
GgXwpcZX2Vc+vvv6eWMFiOnz3Rd9XWwgu2qT9ak8xxOa7/OQy3SX6fZT9x35Iwb9rIXEDGFRoAyU
shICFJB7I+4HP5bF6+Ve9pEtAHB4ldiOtBdwUfwn4afhWMT5AIXAI3KUllou2au60fx/ns2u9i+t
Cx1eCl318p2EV+uk5cEI48Yzw1L2SPb5HID5WTi9fYvjPLGaG248/2jp6rPe9ZjR0ji6m91YEmyc
Hzfexl2rvS7zoqDDvJVQC8AhGtPIjf16Zz1G35dIkr3thNuPIZ26SSU8W3r7M9WavbdGnksVYt1c
XHyjvBMFbJxr2FL2mEhvYs8Uq5PTIPuibUEhmadaKpn8urEbti9NN928CeHIXflh7OWJVH2Rfy3g
TjTP5Pzu5pmdejnbiimjd1SKz2/FJV9Td1Xyf+6e4MH7PFx3teEw8e2KZKeWbVBGIElXqrWqauNb
HBxEE3DGlB/6B6h3U94nf8ChKMWG5mu/RH81owTap2laXeFZB8MFtOqxudGh5FkP13iFpog/8jeP
i4sPnC6uDvcB7w2M9+pI8PVroNF6nz5iidFtgTIQiwokP9oEvTWLxAeJWi3RO9qmNj6PU+Xb4ab5
ybBvzs5+sYp5lrtqYCTvleNhv/BvoQMC/YkfhZj53cxDekXUgCB/2efi2IKnLWuesi/3uNpCkUFB
LeV1EUcz91cBF8eJ6I+W00ObxPulqvM/zYDgpSF/o57ypeCdml47fxbsF6A9Ew31dKq3HE1Y9LfJ
A1UpBVZb9as191lHnAzDU1LPqJr3FLBu6Wd3bnNMlQuYBbQO8RppZHbWZb+1mTnPSIws79RtqlMg
JPJK70bXW5JjADLWsb53yjxHilo2ujxsp1cp5okEiPjXDI5RLSUE9Dx1Q0OM88rg5z9JjW8K+jJ7
ird3lpUUWlkZJHSxje9r8/Aj1E+l5kU4Q0lYUWhkChaTZ8awEWAx65Kg6ZjXjlVdP3R+dN3eev9h
FClUooDDGYewDbABvC8yO+hhIs2GoElZOpbjhD7hQoBuR1GTqahIJ0esrtc2ClanMW85fXLm9YOG
FaPNRHb3bKT49XDqQ/2M9oYszAASqiZ8C9QptJtPdJWbpA0aZSsJO/wULElmL/jTH6lvUK1KF+1Y
vbLnQNrBIOQbOPX+kuhADFDAFpTH50zL9REUHknIxEvc3SXGu+X7vMhVyxwoIgpAQv+Ski8HRPDF
p1xpsu2Gdt+NwHIodaw9Ur91yIyFhKZOdZVs16v4T2ba3zt0ij/LfjU0JOjT6pmOkvvXXscSTMPD
//L9uCiUpeTYaf7YWv1y2jACwPJ9LZ6Y/Ks/og7xWkL8XaWtlUWRH334zCMKQelorbpPDmOHKifx
kIi/CCLHGpHlULj9Qmy/SbfN7fGsL2G4mA8mY8LOjdgN4Ae+ACkVRNS6fTSiP3nATfRUPGppfL8I
0OjqNUKsWdh7KjGCLe69gzGlmgvQ1fU7za2iSiHWLjpZvPyTukY5tLc30Zl10GomWIM8gQv99MI5
mYkZAx2c7f0HdA/gsrVcSvkQfy7DVo0nJ+kS4OSzKxzRIqd4ezAKqYuoQYNyqyXBfLnlq3yGJqf2
q/2ALCw+tZ63DtWPIZbJFuKuo+QIfAlhUpR+XXkYzOvhMHJcwnwBTe1IGIOyvjWAkKU75DZ78L96
8Hlem+iOPoiK+SxRsN2QkoIwqGb9PmW1Aeln12sNOU9/MC9JyYMTQEjLp19skdEtXqpH8wPLfFQR
hQ6f5pGY57BKUv736drTskhXfaCyBQ/UyEu3DoQfXdE8DoOR8XxLGToeUWu4VIMMtgcj4NVIMLmv
oci9Ywg4SauHsBo4GAaJW5c4yCAtxStm2pP3DlQbCNaEj17jubcYlv90k6fdVkZ4gMfAazhQ5snH
7TaiCLkbWltziEEkqtgYp92glBo/OlaA8mw+WXf3WEHpJQS4Ye1U/ukA75kEFJuPGIcu+uf5mxZC
iDkv/ljpWjIWoSOZxySbclOUMuEPVO554kopFbAf7mtS+LoWgwPDj+Vp36L0Yn4nX90gltN6eQAi
+4sQ6LS43vMIzVretV3urxUY3emlX9wsgPDhFHkEUY9lPfx7xPWkGSkM+Qxl3O22crBz8mLxFnyb
+1dwrWRTumdkDlInGrO2m+US9su0XpBil42y3wzGLLHJ4AD5U7gFje4oEW+6O71CUNvEPSm/zG3/
PCHu1MqViNigAHUtMt9bGMDzWNfDBOB7r/FVXqwB8KlniMpFo5A9M8LlbNq5oCRx+FTUaSikjcDb
hg5vnF/+IFG6QSKVtPqPn5H32h0V60w1PLPM1Q5vR1CF+C3jAPSVF0Y58DvrwFxdFQnHeYjw923j
CRmgxWev8DQt3tSu/+YCVJGztYVMjfATEWvn2jv4+o9iuWIWJMeQnx/RhgwBcf1Uj7qUiTfhxqmv
Zos3pqCaAWRs2jdj/oXU/RHVs2RMxxWMyhXNpb6wNNa/pcjSYqXp7TSZ7+EBEey+kjEil4aaycDI
WSHJOiq1Z4hIjHjrPxzazMMQaaTWmwW8DgCxqWxQIlQuFkcBDXcCZ6d/n064vPcxXM9ZX3xJGUEF
MwcKNnHB03487agKdKGvqaTx2n/utSzMi85sFrlS/SXmW/HtBU6Gk480LCjK4v6Tilh/R22aFwH/
B5XVkNdRveK+zNGkxEWHhhJs/f2s1C1eyo+yF8PTe+Cw9OytAPxy6ejvfa72mHn7oEV9RV7ZUPzv
ntax0A8TT4G7/6oSTnstMgKcndWuShTfFL6U2As7CGlpzW8DwIyWiXR5wxV2cu9rQ5RjsKzKIHCv
qTkyqbsoB/XtsB9pvPakwGfe6SZrWH3zgj9j7SfA4JmxD3KMKBMO4Zi/Ck9KK07mTDtEAa4kmnXB
ff/UZLfU7+b116LDkAdX+N1K3kwI68v1HUxD4KXh6kMlsjUTtV3jeJHKCOhtFLGmEAl074bi9937
+uTEB5tXP73FXM1dlS/4yDGGb1rvaV8VIDSysTrVGIQErnoBLpNZH1YQnpk0mjiOn1pmuPaB9QWd
whLQa2ygyVeX+DEU213XSMsnnmq3v/NVXlsHTr23yTh/F1fvOraCrn0zbtj1XcKOYmuVhAczXTWU
tWWPZd/10DxsurIc+d92IecR+s9MSB6nCVZm9CkkSP23zRhZg8fAvRew5odraUgN682pzaoE5vm0
AiAIhEvGZLcfYDUoSEfunAa5wRqcZkstdbZUjtUmYB+gFChzSADNgACRky9/u26cm8AjnTtIX9wM
FuPaB+bs8J8WGkj68O+ZXWVw4slJ1OP11h0oJNpg7R+v8hcSUADr68JojWuDjvZksHJeyv9FmgYL
3AQS139FJfYurzWx9ysbpd1OtlWfxqyi9AbXCGVkvebstwl4o9d8vSrBWpl35i2whAbrQWgcyoSy
GgVyUGzhJKfGkobUn4A/vDb4y06yEIRBX2F+STChAMPJIbykVVePeKkqvXlTL6CZQrocD2EYlnf+
tM0iOo2dxlxwhCvW9BfvcipphRoFN9URQBlgNmxABVes30yd0XHAxkvA6LG9PeOldp81t+iW9JEm
7m2VSV4tgSAUdAy0TNDKBZyb/AlmGEHTh/u3mou4dqpdztIL1S8l9nDKcEbm7PnXt5rCOyActMcD
ZcFtL96TAC1wTLUpMoFq51FDsazokbzl2Rw+KVqS79iJ4X8rUDplbJCeEs6LFVtPSloxNYe2RTj1
tbsvMKm0hrTckJMtdz7f6s82ZNg8MpcRxSNhlRnXZMG47f37OnJ5mju6E0wGRYuTHhd3f52DevP8
cvE7odX3jhH9e+MsAYycse1msF/YMrZMKDp02kepETDd79FERzrUuRQ6D6wDzoQskVioIOjhag3m
fiEehacuWNwlxlhANzzHli1Wu+5Mcas8yuamDN5ly3u0dVEMfNvAK0dQ0JZB+oZSrOmdXaX74On8
wm8RgYZrI95dlONpYO7aw7rtLUGfWC4KZOIqXCK2a/Gl8Q/DRDq9WFAlFFpnIVcg732DwaiJO/Qb
7vNhzPPlgPJ/UdEzHIQifrzXtHAup+x8qbnoN2LOPw8fD0dgxL8hDj5MKwBAIe80RNVgEhQUBPvD
WyRdymmxoAbyBB4yfs4KzRmou2ku0h7fUfv95O+SDL0aeLgJzTO4yrZC3bPVRFhhimE8Vz69VRcD
W6++W5LjWzEees+rMpUodaYhHeRuktFChBToFr17kY1SaIAHDNPA2GJDq1F0nFfF/3vPZrjevAru
ZqQdzow+Hv6HMOREuxo0mumpjptL/Hcn9aroN2fAKM9hxcD6KJ20KacDw+vmgSxZqJn8c0/e468e
Vmwi7nSbLlti/B9f0d2+HpcYwHVITl0dUl+EY94HRGLFf9U7fdCGGFAYXOHjogOBq97YWjgpHay+
rwqs/u5dzjrA5Q946FsrbW0dhtHix1PF6XEV92ayQFcg6hK2LVoReNYPwqAsDgHm/vf/FwweoAq3
F6wthLewVfhqifLRDlke5TsgpAVm9AW2nIHYR0sN6LdxQzz96s4MLdrCtibttsr5T7OV23HyG7Yp
iK1qDF6gh17DOQl2/iP2figlXwcH+xIKYfv/Juul/+IOUaXgrCir/olitSenR0augDR1B50cJ/zF
u/V8hK7kDkHo0X6ME41li81j4A2+beemb+0X5f6pxSdkfnEink033kSAUsSBYzXaseb+8P7SGEVW
lhU/oEPqznArfgZXp14uCGX3QR1GZqnIPgi5oQogFwXNzLcugnRtVjio/eNqDGkbMjJkrP1LLusm
dhlCh7oRCRuN5ai/zPyBNRLprcaDZz+jgPTCGDyV4bmP7ezeJMMKAD77IJ0XGcB8IgxawkE5mmxY
xFPmd+kXN7JvgJEmdMzUhp3wK9TVlphx6R4a2/vOCKz+ssM5rG68cKLtjfSYfX9keYa6MzH6NViX
qlHNHmTssvJ5I8Wch/iMjYAtTkmmEEfwI7n14pdwbCErnN2APh6r+pUjupkWabLprCMBfaiphZFe
MxsYXq0iNwdUl5qJB5dTij1gzy02sRkx9EUV1qQJIc6v8BHgE+Oo8W25MshrhjL1lcr8itLfv+RN
l7vLDmCXxlIqbTDdN4CHG+4xQk5g9t+WHllIzRa8rVB1nlF/laAL0Ttz/hz7ySb5moZO+Duifycs
i2itZtLiYT+bFqpmpdd1zV4BYzZUmypyoD/XMD2V2OZXA+qO+3Kx/cGwduLpx7eYmysVW8ImXumv
9hM0BfuzwczZam1tUUJIyyBurEbTOldLl9tt67sAGxxl1BGm7aFFZuQZm1zo7rPJEvr8MaWAK18d
iHPwERTlx+0SlHojL6GAI7KxmwQ7rBRB/HnC4EIktNObVbd/Y2B9OtW1BECHCgGQF8VDswQGY/Ul
l97n7ob9kDT3oY41wYWvPlVk5NEXS25QPXC1tMSZdFH7G4KnknrWs79LBAsUo4dHMUINzCUYx1VZ
QZ8uuBDnqwxxMFDJB7y3AzIDKdrrNrdzF5CqWEEvQQBQBD7SQlzIPCDHc+UMaVPu3UcbT06SP2nW
r+8l9ktV9O9meb9Ty/sx3rG4QqhesQaQRMUYYJSJa+CVmH/gIkcy6RAhuuTzZyv+dXBkLiwnRX0n
ZXmaJdoCuduxoAgtVWzswNA59s4i+sTdUTtr36klRdo92AFXSHGw7FQVsWfyJCjji++VMJLPVCdp
lyil7pcvBUaCtWu2meSJFY5jZDACx2L1Y7GXc3IYmZDJB3Rlbw7A1z5hg0cMM+oxo0bVDsNnKmC3
9lMFc5RLH32hUE9BmUKQrjwcOr/x9+qbCYyn76W2u+5++/7aTgiCMu/4fWLrZQXQV4Jd1BuK5jOc
Vjtq4rM6WQrT9k1hDKEiERMzFtEHH6BIpwpl/3ABjXZgdo8AvSAYPpzqyPNRUeT5XphkqPHKn6qy
vBMszE2powmN8n4pxppxT0/vvOI01prXoXXkbzg/EuSsHB1+WTaC6nevWyAZp34quo2MBArP+VCw
KfLdaK9EHKYcYz8aK8vdAGMkjGAzvJ/CTHZ1jIkV6uy+2X5AZ7/hQx2m81pcrs2dhRvZth18PXp8
/p5UIhibPaouDR4eIrlmOIo4OnBmQmHBYhKCnrnQ4AVT7qqn0Yr5ZEDJ1KVrO80fOq/m+NUW64nF
d9EBF6fqwmiVbRa21QP8CWeqNU0sto4RpGUoS4KS7GSWGNOLatnncL2k+BwyVMpHOVNmYDnTY2Tm
dlf6eBehtx7Tn1/CNune0xg5JQ/7dPwdabxDOXMtFJLkRVopdObc6Tz7WxgL5GdBYxuJBjMZjeml
iz8ttmVvCz/6z/WAk3nXe3OCrkUnY8mSRzgkcckVJte+hVgolx0amT+CVWaZf3gn3epis5NSbTQv
kLbe+/AcQVvwQ0rYv2VKc49eYNGH0HV57ZyHzDCDIjEXEWJLp08tFkgbxmx30kEX/h4kOUQPk0JY
7CyeB6niZdgeozlZYaABarLPNXAyvNPMZt58eppcmoJHKU2/k8vjYCpi7SE/NOzf4XEOmX9alNBe
2fjbn6K/d0HchTvb3Oo0xbrexipDfy7+6RSpLclJVnqeYT4jQEBUiy0qZWxjAGqunMvi8XFUJvCe
AbPU0QeqTlFt2iDH1MR29kdHwyMb34QmrY1CRH1mpbQrVjmSIn+RsHmucrNWcwedskAuYZoEEjdu
QeTXMSH76s8AsuJj+vQBe9sszAeqz4xnK/BBQTzD2/mzuvLkLYquCIju0N/1ySmjp+oaOFjJMOgC
tafdN/UtE5vhoyVkmSb/52+DyH9/3IQgc7W9vKd+5QhQZTR2FTxJl22oRLD9S9izMFLASAwY3d1l
+SLXxXDKzHWwjVKomABV6O4OreZ9zxd7/qOH3XWRauJBVNnx7SNdOwGVXD/yHV+Be2DYNRxmxNS8
gUyFE6nvc2BRV8THnkS/WiXiBOpBj8j+LSMH3+yDPgYkTnWSR4WJ/VgAlC24clD1Oi3IB3KpfjiW
VFsNc9mi8JCbFJFGisx0Kis/zMPXPo/+EsSfhn6IpAE8uuVLW3V5WOghaRajY7su1rH4JS9Yq6o3
M6iH0eF9lKa3JMMdvh2PaNusvq/9sJ+0304SMw+rDYAQngHtzWjNs1KBICmWnT1FTFAWEpEqTve8
wTTRZ/t6Bws90SIrkjWnmeURrwiHT9bT/MpS248BKWwAHl7OiwZxLtiW/1loASB3otYWHJsJm2Nv
a9Fcuogw0JEKudUoKWsMGS/N4hcmPa9qW65SSyCJIdA3w61rHe3cqzELkOJFlxcn5Cd9lWRM21gv
PfvvQLJlJLZMwNOXpVMKUc5u4YLKCe0E3GegJpcwPpzMGEziF2czYj8fV0pZ63Sw36b3k94Fjcl8
ldc5vZXjzqEhczSB6S04/mQVBugNrLkDdNUY1WnRT1yq6IA9J6gQTh1yyScBvAkFREpxW8wFqMPg
x8hX+zMVpkUvrrojCN9cEa73N2oCS98fZyAaHOuRQj2eQR5pMkWr8ll4rMID6I8VH9PAKAUSeFgK
VQ3kRRDwT6wsVQMFpA6SeJAQomWhYE+MY1QFBrwZ+1Fu8UdfjE9r8t3IoKgGpcAC/XqNy0TjYrmI
e+ZiLnfMPp3VLOEwvuWMUnp4WcXB4H6Wq0uWNL4ShCuYwSliK9FWxIrfD552AWvEOeYKOpgsUqtD
QaGGy8OcdzOunWaunMKCEqxIx2EVSsu6Y8CCuTdkantSwsxr4bB6C+eW4YChIDwsplhnYY1i8DSV
yaNpDPadXRHNgh4oiiY8Z77acKPxSiQDaqdn8ubqoE+00UmNw5zNm/xzFQ0OJXkr4+O0dLSWicSr
rJSe1+/oi/TNLnY48mWDAQ1JgpI2N07ytOHt2C0PgT6T9FWyGLotQH0a1JfzD52tjW33dSz1x+EV
QkObPuTG6JOjG89ZdZwuiZIUtwxjE93FKJ4DsuPsjtBTGyHz2epxfwN9t/b4kRlGraHOxunxemey
9vtJSd7reHBfuRowTzRk3u+0JWVcnqSoYXI9dSGihroIb5+bkHuISGIWwiIKUs4sEssGRXBunSfR
YYGsnSURrcu0j3xXo+R1+FTR/MHQOK71hPc+qV/VZF/HF/Ba2icD9NAyLUQKQ0gKctGMm//foil0
Bi+ghQrQ6hayjeLJ+/bFbC6W813OZs6Yuugww6zMU+FcbSLkc5nKzMwTMkxNqhRcHxNgASiVBtiK
Cp5y2h3wfVyNbEPGyGFR1nksJzO73uR/Ic52MY8/nUN/qji8G9tDGO6eGTPo61i7gOjsRpYlKYGI
1+8OadFRXaNBEHUTXPU1WmCGph49UjuKrsez8Nq6Qg8ZY0LrUlnT8vpe/+CfFiKPtAYw9Abi1Uyk
+C8r26aP58QtAWDFDHudObCd7p2tjf/MCGG4SIwPJTdecbLFU4aBjuigNdUrv0UsroOmKaMlxPB5
qAEDyW75i81QnivdJ+cIpaCnTirC3X9hjvn1fdmSF4GUqHydav7amGDQAK1mAc6k9MFDI9aKugYz
5dO9lBfrZV01Ryeo9YaQROGF6/Ry6fI68X2Tjm7sy3K9dQvqpU3Cw7ii0bTBHeAmtfXCN7QFp3zV
mxFfNhSe71tvIFUU31HCDsGt3cl5+bzNh/Y/ZGnHtBJQ1jMfx6FTH1R/jtiCxIMGIt8ruY8pyuUP
W5aHnM7qGB5fdy2cjHtUEwy8V1TbwH2wjdWE2DsAD5vNQP19iRSnggsf9IRdoApppYmobMlEPrmv
fV8za9vHMZmQ1VNohVhmy35/ln2bKUhBHWwN7oBdqB+UyZL49WfZJvmhP/Cdta1JlaTmTbBhQXz0
LcYXG0Nup2LrQBcQcWlK/ri46/EMZcdOhxehACiA8OS+EtoFziEAaR9SS9eZkTw34oEIQRvLM/Ek
fTPwVzV8/00i5Z9EzFZ/rFQtSIRw0iBy0QJ5jJHyZDqscdEDOB7quUDgNtdDHi6q42ARIDGfEN43
QLiU7V/T8t3dD/hkZ5UyhpAKzA9NDq9hkDhQz23ctFfPXgh4NMwN9B8a8je22ZW8CPj9MY3AGdK3
rVHK7B/aAlKe6DEoIXk0qM/iC4y0PtIina1QLT0o6kGeyErzPuWb2OVQSxYePhiufnHn5etki8ky
XBGYWSS9C2XE69Nw/IemoCgNamDDiJiEVspsMsHS3q4ipCzAWrthxUpp/qU4swWj4upXiFk04936
+9++pKNFYnX/U2wa/r5zDo4x4Xm2ZlYZ3iDknyp2wunUoEIFm8vwVXghX0Qn7s/cB7cCDheqkc0o
AlJXJYpnKX8tI/aI7xdU5LaTfS4JYnG+0DpKENcRfwIUo7nqJYrXYzmaF9riUpklA9sl8HnF7rA1
AUqeVk5WmCVcFWynZQ7+DPWtFYjbg4OpHZo8SJKmnHRA4uZWO3APmRoImKzsA/2zlPBEPb6qpinf
7trxuUbdbqrr4syQAgOPfBzggOiMbmrJl0avkW7tZYWKjjsXCFQ8694fXVU+xXLuoLNQ8FYtohcG
2D8OVc1UE/KGxV39IEjPxgliVN4jhaUydynwK4VL41gG0BjcQONrCy3uLvw4hl0orz4UcHkQUiPd
yFsa1u2pnifMq8BC7HZLfj43UMXNTA1yAdeVvZrAMGtL1oBr7Ar9manHybIR6ICn/h8lS87ZLHnZ
XaIqyt7I7yBUNx9j+wYikbtuVkYdILGaO9XffIH8J219Cs/9GJOldbsI9GQhozy0A9drCmJWwaUI
ncXdKoyDLdjoFULF0MlmjiBNa1ueC6Zxe2fdIxWOaM9wos7frFqYZ28HQ94CkdUbh6GdjTITDmIj
zwCcTDPyEccbWnq+BkAChBjKacD8B3PiiQ6kDL77tn+CpivmyDad4nS42ye/ZS0PY1KhlZV8KeoH
QAZMPSsGSbn5YYgx7PDMGKDqCJ8HugB4qAQ7pZGpv6h7Lz6q4WimT5cf8cRSNCPaRqnzEvAUpbUZ
8wR0agVAi/wrfXNp/creBzDg6kc1X5hHXFHCTq5nE6RNSxsD9R8HbJqhOLqyRNz5qraqMEW4dj35
mk1qGSOwMx5T1QrZNnmecXexnnJWqXWCO3Gvo3wrIOKoKVEuUG3Hrq3QipzqZAl/Q0/1vBumfQDp
d+qVLFXai0rA+/IvEc5inaCHO0EkFPzyoMEx0F9cuoOUYler3hzNgo2EVVZBpBGDOrHF7nc+vvsW
oCL61G0N74DQz7q+DyNVO2nQ4ZCtOICQLXlIshnrLsAt6pRYOEYJ5wGydSYc7Abb1oH+ih94zn/q
r74d4HrqIy1LXcfLWZqHYJd8X4FVEgdapJIlfUyQdmBWlCnYtyrhFZDpH1615H71sDAOW9cI9mdq
9Se1Gb5TsTellkUQKvvr1mJcBFCUyPC2e0+Cqwz9ZQN6DOM941JZUCnFEUmr1gWppInybPepxP7X
gVYumHQTcGMQbF7ySVIB4k3su5aeM9ogldU9exuimkGCHwALI4bHonvuEOnULmbkrXKQeJyCjha9
YGhX4YRBocbtpiUbleJfagDFRVecWGUiMHvh5CwjUOehFv3wUrgiVUD8sUm7d6Yx9Lv1fUvVfR4o
9WlGRiy8qqYP+H0UqrHzKdOAN0OIEPBodhL6Prd5DnbFrbrO3LL0oLki8AgsOsjKppZUtgi0mQfY
G9jCchtVAJtqXSOaaWdN1mOCm8mTSWzHFH/aWbZ+JI0l/vBc0Hijs48fItqehZ0yVM2Iewj8COc+
Kn9gTlCfqFb33jwTB0UXfSseV+q0RE5y3dC4wa142vNd/E9zF0+xJFkZQCrh/SnrcbywF5td4nCq
br4fYe/xK1Xh7cNPHNUrvPojd3ytgmH1CHyOqU/Q9KJHVTF+ENLVc/cZQQn4wFviY+R7XhH1y8es
iuWQ/dFz8ErrkWWQEaZRIFzeQPjq085R+D44HT63l1ZwJobvrTy99e6StwGxgy6Np9mitBupduRS
TP+cV479QdRFuGGDOADAjOulYIwqs0iigeIXU8X1w7bjMuco+j+B1XC2fEt2t2Lq4ugWjJk3Qzrs
O9VBLj5iNO7a1OSI8zFpB8anUpda32OrYjW5q3jD9yIjZ6ep0fhR6okRcwCmAGZjd3w08+BkEYH4
kbwps531F1fkHQVlB925An+kuJHU33xc6rmpBGXbChW+Yufb4nvSSXBtZFc2l44R+lim3P25Xlvu
ZeWORQ4MREtT22L6Uj1mG+ryS0VuPjavOAIYFbT3DpUsxksIuI+zeEK2sdoz/OdXSLIgKy88i6NR
3Dom5q45VaoM1xGrFd0ZHy+8FfIakNI+BXEKQKMBKq/9pS8Lgx3eA2/2Vxhvv/eicTvnaEPt6q+X
AT8vZqDUr5/eHlEwY9QQObOf7gxK5LhAEICBdEW+f8S3MWtHik9kHVc0wsnudwGPgQyYvgxyFUoP
/az1DRFa7csFZeWq/CPFNe0gEqdboLiU3mBLwXL4S2Cqrww1I3Y6k+zd7Rwme8bBAFirIhxfH8jR
ydmfaeK3SE330xnmFI+jf9m1WssAU5wVh0hzyJ9BLDvL9/4aUechGoP5nci+wVaTShZTVmvedKL9
1J9daykqN5Qc8jWjTaOKG7m3g/atyZHNEoX61t9ZItI9pRiGU0PX15v7ti3g6cZi08rjB9j0VlyP
VMj8EFUcOVQrt5q8BFVIqrtnkl4zTqEJrekLLpHzjKFqXw6ZbD7fK4D2MmDaSqEx6ib1C+HZcTde
gmlJWgARqQQN0QLOcZ46UFxvOML4MOZ0TQSooO4t9Wj5e5ZOvVW+MC0u9tu9PsLaOa23y72pdjiM
5IDSi6DOE/5BC5aiRViCsF0WWeBZz0udzQtVb1OORHtbiKMB2ERPPSAL+Q9FxLfCOmwA2SsR5sBd
JU4SVH59Hde+/JKyorH0DIgcqIyzh7L028OUXAR3czu3JeYncY0MdV540IkWYS7tdZgwNBWLD5aw
u98JjIvKsi4ou43sIBtG6Sr8Y1swM7AcHM40PxKw0lghYTLvvEDnMyQwxERpt4hHXnotaqZHeGkU
NLUOTbKat/UjVQf2pRdkJiSMquYNHGqctM5fzMsfBlzbDgxbLyJd+SXb7BPBj5AEOTmeQzfm/DGW
bRzRc7vz8aEko75+c9xlBgcRwSWLqTEJwNj6Mty17ogdbMrzteRafhvQeK3KS7+vhKleMYmGXjtr
GfZnDMllMBKexpqUtac3NWglJbk7JlwKpLQsRFRXBD9ew/zxHiFbWQ4fgJE178q+0i1f60HtKN+e
DwZdfGKR268PN4KodsNgrCsf5FLTS9wLCC2Pr9evrzJtGHluEnyOqW9HSVBDzffeMG/ELLmoO7oI
hJ/SSC7ySmo7RvPq+0cSYYGUkC0xKmBBfhqpC5lBPFhEKUQ4cUxjGaq1ibeyuaw9aytss9oRbugG
vUb1jZ3mXxYeOVEF2ZvzO84d9rw7uhWTXqh6g4SJ4JbJZlCSj/a1uErIsELYwxDRjSmfrH+TodAE
Uuke37YlqgQ6K6pylPecqpBSKWWhlE7aE/xN88Ruu6UfJmmi3cfRUkfy2VPgBGiGR1NJTO/DUym0
uM7u7/ATNF0i7l+vauvDBRbna4BLWO2dhPAZ000bEhyrPALU+U9k6oXRzh6RyGzuk03zTc4aHzAF
y6LR8zvmzmwUSHhymZUuvmrmxqudd3og1Gi/o6eKQvVw8rNQ+5JtNQ7uADEKHcVILVrgoy+1D3J8
7cx+75Ii1eiklPx7VkiaPI1E/tOUFSxpqdRpVrx+T619yasvSBWFp72JaTT5mouKLwEu3NSl8kQh
UZHP1T+zhBTTvlBKetmfMRVnNVRbx3A2sd640r8ex5XeI64gls+aAuaAYPO+/dmWX02U/QJwIQHV
zd/dy4STDg3/jm3O9t1XOPninO0PSFuacEYJ/EyP/Zi0vzaNLbqDViVbf6w5N8XEBY3CuJ4jVAyq
pviAcyTYHvJZ0XtNhSOdXE4wb8Iz+qafcFteGlRsiYJsCNRsSTf2l4nra7MdQmd0mYs8/RrZQy1g
ea5mmtanFKUGXCspgci7wIQ1RTKrOsFzwZ6f36jRp2LEIvhu6CUuq+pgvStXdnuY6O1FBROJc8p/
PFCSkOAhe/qQQLrM/Q2Ha5i/nlR6yTvv6QpXnzAvQQiC9Yby9LTymPB+74FE61W81S8myFedqZeT
+4nT7MoMi+x2OyByGJoYKT4/0CmEW2lau2kqdWshU372dY4udsoPgPK1zESjrnztgJ29l85QwglU
LlrDOlD3rX7gXQQeJTj3Vdq1zF0alqkPtpws0s/kUyZYl7j8H6hosZzy3hwDsLjU0lISYvh/MosM
S0gYXUwRcDfA/K0B8Yb38prahrHq3PkmDil5DWWYun7p849PyolH9nND7G8jCa4zUnh3N7e3Z4TV
laSB8dHtJAzdH/uCBDXZUonOuwbh0Oqw8Eb259ylF3w2UmaiIz/LLa4Xf7Lz1a5ExfKBY8LrWHfr
15ceLFRZjKG2KAKqnVSz8E+GfZ2MPvqeb+06UMXHleN44Nrl3iN9SM478sKLHDX3zd5fxEkK2O4a
sGRYKD6EdNvXZ+EonaEHsldyM+fSoGliuUh4KTMW6K+jp7NMnmZF59DZK1z2ZZdybwn1a/EktgH+
tRD0m6a2vsB+EG7vzperDCvXKAlWN244N3T9Ku0f9XJqiCmiI8wvu9OThqB0XLWjKPaGxvlQGt2g
fdylFQ/8xXPeCajRekTRLXA0EzvVuVhGNGdqjQ1DUnTXNrsViietcrJ92icwRJNm+bq5QnUAjvNE
kl0L0FSe0/dPIY/bjHsy2yLaFWKK6DMPGvdgKNyX3mqYmN3rWbHk79f9WbpXMI+CYfzYAmeSTKej
ToeMCNUz5qFtfQ3g6EC1w9RtxrDwOb6WZISq5qceU4BHynjG6rY8LLv6ykbJBdjGfSYLn1jpSYGv
wZ8Z4L/L9TtP2ToiDF3gsgrSrQk39YEhCvxe/ph2/qG8rECkdFEuoBtSyMLhQDnEp+/sRG+BJU7T
n5pLd55Vt4rLTg22EWPUdBM6kS7baatRhPX/ueZA/zkdCoPWHR/9j5M74L9im7IwwppeErQsnDlq
ojXtMHKNAnD6F6MVSdzwuPduaEgbjUjTM3QpCOyXc9OgC03XCcQ44b208lmf4wdsTdgdtUxWxcWQ
/M1B0dp/ZriQxnseWwLOr6WyduqDwcbujvheRI5jnbPBQR4wauLAlqTvLw6roqD7Q4XDzxtZ/M0E
F9mvD1nWU0IAzApzfMJUGhsYtaBP8fztl1IWJYU3oBQv8ECdRE6xA9Sli4Mt8CDxT5LwlHAB2Mja
17QYQcIo7na8mR9ag/NhkrwsSqum+FlSBrDysrH1FaOLjaOg5mRuKV4Lk3foMYRDcJ4M7wTL8Vdz
hLjBBk/trLpZpHy1OQX+158xOzMu9Nz/f16jZ0RmNTDiwB8c1t7T6aoAcjKWQcaBwOrefR2jAW4t
ZbX+irfkoVEf8RtkSjkZol1GSpYR4Ec2iSk5WcTsO4kggZjX7ptD00QOxbfjg/VopD+ji4wlTxuq
c2gZAXVNADt1M7Hymug9Qr350IKCahNYVM9lYGsZKUYWsd+fjnn+/mHGVP4Jg8nE3DVCMcWcgh6Q
Da3JIfu6dt437qAwI8T9jUKVcvKBSTVKbKx0Q0tNJOPHorGpmuuRsNnvdnG3n7BdCrxDLHedFNds
esXI26y0XeO4X/lDLmDQrVribWZZ1VuzCiKLqAVheqPFCkmXKOzhuBpLqlbL3msAMjId5bJJg1Vm
1DTa1P8Q6tYkuzxfO3kgBtLutv+yt0kUIe9LedD+DoBKpznoRDO6xC5U7+ZzJ6p6f263yZsqflyF
lUROiJ+41E9Iu0mD9RX2sTQrd0UFdTPHF/p4PuuRFbSsNrzr+jbHTzXPWn/SFKu4/dLtoCXONjTz
luFFI0hceTLPMs33msiU9YIPfSwAGTJzTu0y+0Pgi5NjJNO03lae7Ift0q1NW17pad0wOtfHwQfS
yTE/SdRh2cdvr0OMg+V1QFPgUCbm0H1V3671jEOZYj2LfAwsjSCYWOs3teGx51tyRENF8dUo/NVI
9pR9terxUD9pgS1mL45/StX8fWkViwJlypTRFRnM6tvR40iqc5eyY2NI6uiCms5M+1bo6bkgRPQe
yc8Zo2NSG1b0JE5lqMMYMRSpRu+q9rrXRBPVBWv2fzy3UA6W/kP7kuTlwaBeX6HY8hPsiGP5Lpyx
N0hBqA842mg9oyZ+OPfNLGSbax2QrrHjvnTgP6f+MbFzYc3veI+d05N9PgUkFY5pZqtjA8IMcqH+
aDdJeGHzlfkZzy4uL2W3/expcydZVktCSyyiHSeXSN+2EP3hcSGnhySM7n0vBTNqz6EdnCRk/fda
PFopcECpCnmNw0E3SXOTbjZJbRViy9yGveSrCk1sePePBUBL3TRVt/YAP8hiY/kC37yL6ljhGRVy
jHGCg6o5YGLOKr1sKL3087DFCuyyvZgQ0x2157KUxzQ9HZaUPT0FnW7ftXYKg+tdrifgXbGS1+hJ
/jPbHgkNhsyaq1q/5Df8lgNX0l2g9W5baYzzpZ4mrOXuOy7emLJuclV24kUKeo+hTvI58jULIvNv
cgBigJPOVKnUu9BUnliLGT9BsH5ZzLufGGfXvGFVnpZHWQKy/hbzJ3U9iaeWJ0cieKCyf3ylzif5
XakjMvj3HpsEfwZ9gqdV06QhRs7ZPVhhEl8sSB7I8AYqoyAThwL1YOz8iBXk3qzAp2v+/DKzTaRW
HQpfUkkqRsPgEZknxMBFNq7At3uV9nydeMP6KLwOxL3VS0VHFvf9QrgqBt3zSMz0DI8PMvK70i2M
ZdTLFozDjFHNOl5SL42o3cbk5aTaf0k1/q6hXVTJV+dA9MnCJgAT6SzDu/NveTBUEzjwg5gLpVex
hX5Z7+3d5CCfhZyZasshgXxTUEftVrp9fgkALBZ6rbCadu4GIe80/fOZHge9F52NQQmcfaRvYfYq
WksC5DEfg5BySxpBOPHnD8BLE3qIf7G/Va4Is93XSDUFJqp0eN+aKFpfQY/aluf+YchUxtIujgmi
Jwx+7GJiXvzAfrqlallm+x9/RMPonKbhglEPUqrzaIIRYmQQtGZpHlA1EV3vGj8Y+vBZrXRE7pNb
sX7Tg6FhqZ0gkXW4LNSN/qubLPKP12ncvCVTUtSZ8xrqm00YuYgYwFXAREhyOnXLWm6+G1QjAoOi
wCY2Sx6bdKd3PfmwaAaG88w0bL+aToU2mvUslExHIXJPeDiAsNhgI0HS4Wl2n25dWdUI2+iJ5F5t
p9A9XoDA2P9SgJp1Ya9b/x85RoOM6k1vrc0OygZWx6wiUkFXvnq8SSTI0cCDnGVZ8dgu4HtPlggV
Ss3likiH2TRZPofOs7ljzmw8odzSVXX4oxmRUhkDMvZbfEKLhN6kk2H2ZAnmOAAc5eMpQ/k9MUHS
xVwG/El8Htxo7qtcgjwKzVGAhl89pEJabSIxZ3VEA/Z5NyCCIyv7xmFLPWGh9jkK1+1lNuMGgJHP
9G3ORGU+AfzQlCQxzwl4gqxFWx3ctk83ghbxyQtaPCX+jgPVPyndSxng/Xf7NOsX5F+pUezW2k2v
/q2OOZlpjbRMVrCkE3zYDc0/Fs7lxK7MRV4dQtUCD7fYNYJbw7F280eCQpdpy/SHcF4RCJlyHHe4
vFlX3FZKj7Oa6jT4CrPEtvHir3Pkq9gJEFDM6PqNNpk/RFExErRibo+hkeFdZGoI83VJUiuYPeuP
EzYKSodQyVBbiRXE9X0zFoUrbTYNgbcAKXQPldtijPMbF8nyEpwskFDOjwaOUoApIy4DWzXwwXbT
JJP7lEYPhRgbabxNIMz6/7DUZAZXlBjpSj6jBdSqRwe2b4AdHzFg1QJxOl99yxnGQ1I9gfZAvCPd
baj11UigSD9Tz3N3ClIEfRwHcGa9M3NAvnu2ZKdJklwWXPc+2COTU22cUGii8+BJU36XQoIobcxH
6l7PwhznDVdOeusLqbBrgOj9FjvuZhYRhQ95ApF5DfckDy2gMJQ/K8HhK/S7bhqFYyGIJdXhH8Wr
C5N1VmqbbXtB1KK70LQqEhjqfvG9nMnztxzwKHoHNIhQlys2GtJt2tssZYh3dKyeo+R/ZdnUmz4g
ZUNisZ9ZrLsmOAh3FyegRdMkPyEIIzM/NnUa4sWNAIX+xXk52BkvfVC6coNTjPJfBrNuig9Nlcqc
3dJeDiyTEUpnZNxmk9sSsZGHBFvgCBtitwxYWXjc8srByYyqbrziJlysszrBEE1cg0j5uzdIr9Az
HHT7qGjWwhrWZ/UMYROld6XxLuGcoIDDrDol7RgduFWFUnLjpfP8hWsp3gyKacPWt4/W6fyf1XIu
dQVwrORYl8zxQQr3mhjlKPkMP9ULU/HKfqCQYJdut3RaTF3GVJKAGtJjUt8OMFPp/7uOGg80mRDc
klVd9NHaS3DzKYlU7wnkH6p1Icta1yrtXQd+t1AsBeiryHwOMgEX/g2+hirkxPU14szyHdioLqdp
5wJHQuh1+E08Mm4ajBBa47DojUfxo3X/pwjUVqDKzLBnesYS9aHLdEv+sMw4vtpK7V7MwFmGA7Pv
K29zDChhuqyIpivcIR/uCyWs0sxm5kmXonHq4A5gta59wDDiUK4BRxs/m9a3e8W656aLMnDIaT9l
s6Cb6szBxG9ILP9oAsCCAEwFIukOWSHVqmTPYAlTHdkdM41lTgmTCVPAN94zPI4ws5AabWd49MaR
7FRLu2wwpNJh+zSOoJJdT0a/02CsFVZrjF/bkyCW6XcJKYB8hu259KN2m9Dga3lw/RgxL2nde//p
dk4DOswnCYuYMyaA4MJYlRftyB3KVnZqNepmxnzMAqkVNPO6O9UgL3erKUmPfAKfeZ76+HG2H1o7
O8B9rFM0AM9jGVF4VZMDtl0j66BNo76clOqXeRX6C3SDcGsBlEw3wb6U4E1jSouWAPHLV9o4UeA8
tRseNjh7tFwqCBqQU1gOkh1nLcaq1Vqn3aglsX1HxwALiVb7VmHYApjahtadVzir0omZ/eo3rCzA
JeRUdMjqvT/eDC0+9+k+i8/0qnFSihEnem8Xwt/YMybPSVCoX2s2DotlF1pVONT5zHBbbW130uME
yo+0DeMkHn8EKbHzMYoCZ8CSgxkzyOuTXeUzO5EzQ/DzmpbDVSv1nlkOG2vnle3J6Qz1/LHEcheB
ULJR4MeVPFAWiwS+LOgfZPOWHC80Qdr/RrQdr4DeeS2/FbdoeNjn2aYqf+Z66QIY129BocwAOZf8
ipefcV1asd9w8DSRrSCDoNS2cP2tM+PMYtzFHuuDdJUQW/HN+eBNYowyfOdMjEs4RblBfHuLUrPs
Z5A/a4XHRn9qwOAADsYxH5NOYRKi3KBpbftBAGtuToAN+Oe+ikUALmsDiLNh94Y7KrefPOC1mSWm
UhJaDNJEXQYRcauB3eWM4AdJPVa5Q15XI5z63PfdWX1pLMYHBrCA0UswjbZHnLqp8TORSvpVNqSJ
6h0ztJ3AlCxvuGxSXwzuw+KzJVfANQTdNz3hNNZaNB+uyCYr7s2CZ00HUZgIcXvcfiMhskREomkr
YEi01zj96ZdmfUz8qcWR8pOLIolAT/pligQ1nOf8rSYzNHaIw0vJXD423PyIR6O3RyWlSEhjep9O
1BOSeP3n4AKxZtXeo8kJYhSoYfIQmM6Qyn+Q0UaZCi82U2h4OArCiLttRX6TzlmiSYPigcBaFZ6B
Ea/NOt1IOLEbyBJYjsa4Dok3054pKm4uRu+VnHYBotX4pJ29KRfNZGfpKJ3wrOOXZ+sfhFcr+DQ5
VeF4zZGKPI26wZCAAIYap4jgNxKwTQOlp5H8Nf8RDQX2jVbJwURiSmaK/e4BRpWWrDwNqHXLmaSp
zQ2u3PNmcnhNSdBXyNCWh+s8mWnJ9Tw2YRKy0N5QtztEj67dwnsqUeLGJS64zv5ttyecx4B3EjHn
E8zZhlXGELVcvLyTLcQ43mx4HbasRt9Wld7o/HR5ZcM+fF+rPOYZC2LjfWQBkT2bIqk0zzO9daaT
wnrHTWasa+zmWdmQTVkiNZ21SDK+Ow1mou/2sMzgWGPp40Wv6wA0cQFqlfuRWiZfMoZEza7gU1DK
LXOJpNzj7kDrbXmjh8O4MzNww4kmgdZAXu1ubj164FabOF9uKOg8mmktSqX4azX6Qrf3ts0zZgyu
Fi1AsmecazJ08Fsd+vciINzWGYmebtdyh2/C2/uqpehh5VZtT57fQZN1Ehoe7rXBP8Pw2BxatKeG
4FkurePzcAM+ldJ3e/pxRFw+T3QmlLHv58vZredj7BZZgzkyoevoGYhsVxj2vAAOv3k/D/oOD46G
dyB7Y0XwGa7IZjspa5VgmauQPQTAX5F9bRzyQKL/oSXixQdrFzUXzuVH2C5Pdf2N5497t56IWwe8
pkJtsePSK0WgS68a9yHmUPi/h4WxFhcwpOQGrUxCLcfNDJVQLMbRzuhrUTx1QagXv8EQBKobp8nX
P+1UiPYJtuWD8A7Fx7eDtC4CkS4yXoIclKFqwLu6cfR2wPqxF87g21bp2wuYWjY6bMFoca1R+MIo
NtN1Cwkrs9aO/XWKh/Bt1MDNfLqPp9jH3DVAj2vYinI2nXIaBlbXFLtENmOJKkHxQjVPkhf7Q8RU
Cusy5lo4fqlJ4AQkKkbWNSB3LEhgLR/p4Db/b1f+4YN5ouoj31YX3/plIeJA+gzGT6b+sU+Tae3y
CUDmyVqGPcI8jCkGVzBbsV2nl/s0GkDFOvJFQGsdNNgOlqgiDH/cMv2NmbYwWy32TsNPezJRNzz5
vnGBpHmXy6vSHiMEcF2bObmM2z4f0iemqApSjXMQE1A1GpuNsuXmtyYEtDV/G8FyU6SBbfeh2OFo
vIjSnXWYZ0WlhsvjgQYcnfS6WWeC+ThFCrluadS3oU936EGhuvM3HZWig1V6hB6lTD2JQDVp90YA
Libv2DZ7cVCKnSWiZVls8ZKOz8bqHSqn9RmNk/N6salM79EvlAGU7PUsuxeqfTOD+OClTr1W94Pe
sFxG6YcgyyzUviMm2JisbQFmZhvBWJhmwsVxQhmNN+fNeexAhJSXdfs2qiRxxaasAqe6Y8PyCEVv
wBqM6onzQif2bHQrrL1X6sk7P9OO8532pcURXs20HsaWFksQ+gS/8zANBnPnf4HuEwd3aFqJehqw
fEtxx9qgkcQlyevyWqGOTk7DjQdrI8zSWjP47Dve7YzBuxYKTMGxaCBuPnxXK7HPnRpxf3VFwBst
8Msbi3SshkWWL7ywF/OqytYBS/J1qnxoQCBCOcueizu3KpzE5BDj7SJVAaDJ9EOZ7s3ThJ9kYDc1
t/fqohVcd4KT5ZneJ2NiVIfZP65LA1a64ChBdX/1HMUpQ6q0V1AvfUocxhqwtSEAs5FNI00V1dtt
Zm5ygmyPzTtFSfjGtaLuQnOpw6McluLsKjtQ0hx6bOSjlb/iBJ1LuwQnsCcjIqRtJkR/oZWpavhE
eizy2K6pZF1qHj9lXLLNae0mAIDeg9yRwGIh3xHWrwR9dU/PxUYzWCTcLrY4Ty15+id7hgVemzI6
fpE7/FrVGMamyipKwfGQux97OyxFLQzEJK5Csg+bmp+gUUAx8Rj94OT/2JMou9E1VgbaNN/Znd9H
+yzAA4Nubjo5u1+58X3SJp0GHJfXWWcbyNAq+yeN6ELDa7qdZuGfeGAhJXjCT//ISmDBmyCkLGig
q38em0RohGiRvlSLfs+6nGZUWxrg+lsiGXMszFCFaoylsZgCfYJWRptyKO7SMmuIPGB2gn5NMh/w
zAo0IaqrMnt+JP4xZk2gCAlsH/OVQuPis1zPmphdrqdkAxj7hkNZurtaZo2mSK3jRw/jh2dcTH8C
nou/xYML3Id71+gaTPuHLbyXflil+tnCKiM2xAFl/l9rloVFNVyo2v3BqyaA1KUiBT2W26a9z0Qa
2XM51FHCHovKwT/EqbSDz+YhCI7C6QYqqXkG4TRLUVT8yrmfqY5E/GL5cKRZt6mfpkdnUTAnyZmT
uiBWWZ0raHM9mb2uI2LAJ9yxPiJT5bldxOX0mWMrYbmganQ8SqJ12jhz35OpF08yG1wvZpOUg07R
MeS9dqIQMKPlWhf2ont3nEwF+zmeFadzOfGimm/BfxNysR/7WD+OtCxljVyyr5HApUZJM9nTdZeN
ol1vWlVuUHv8FeMQTWTwvGWEUwoGsBrEUnGXBM+Hn/MwB2fOHB4MDwXt76kZSfcuVqp6wy0Hu4zQ
2hYgugsvz5X08IP1CiLh7Qs0HdVGfnCTH9Zx1AHTNrOJF9DUNOXKp3tLOhtW2UzMaxW44Dx5MT2v
Mhz/jIWmEXsnyd+jDy0U3gFN1OfmeKXwtZ4SnGOXrawCBNy8jT3PVqIyNzsnA08hn2VTxojxct/7
NoG855c+YWaWlVSMdrrflI+xcKldQ3DKueaXFP0TVZskDGOuFkC9oOaAXaSRq89/s0WnUWf/Wn1f
AGrm4cvmuimD//uUvKkz5D4EPahxpHcOjT8XaMov9HRZBzk9uljJ0eTV/U7IEzw4mmQFTGtKmHyn
l/iVBbsR+vinHZVxfZkIlXS+yHTj7XEBO2Zs8VbW4MqF/jgS64pNMfnZn+s13lNiQhHhXG/d29x0
A42PutlhyiuFx9JmsO4151Ggh2deiAUIV80bP+rPeoHXK6Wnh16koGx0hNoa1wbgn0dbzbJX1mFU
wDcVvD2hmf9B7PaLGUtZK5BP1IyFCjRmvNA1Ap9lkfheRI6JYuAhnN7QMcFHsCL6iGvxupi1MFOR
pDJrRfLb7SGebN3oKbWArv87ayAfx106KpHTF+BSD+La6mFPyLyKm0uZbXV0tkKSnJMKSOZf27Vl
2b4IDLJ3kPUEzSAGm5K6wcC/LhPUZm2MOu04YQCwLHSevZgD1QNjWfYBBXCJTxuQPt14WNfj1QeW
wlAY73vX9fhbPpWRHY0uEmIA3wGJwPIVE0Ua6NaDp53dDKO13FowbqVZz7sm3rvIgwCtdk/CXPRk
M9AYeBaHK7pN7xaSGjYvIVUGVJCH8SlxEHaaSknJPOcTgrNRcN8Y+m1qhmjktsdRLgqafLeekRlL
otzp1UKVJyYpBu7OX28Jh0DWolJByxrFtKpPxRlFTytdUBELOGTngm7+BfFTdwlE1EVj+F9paTCY
mtKAZwNRzJ1rJYwNrzQpWh+Au4pA/OBMV+61jWoQhLJY1TnOlc8J40VtjyVnvKcqBSVPYoHqeCy9
vf/T5NhNAXmcb6qCn3dAWen8YoUu1oRQIxAVyiFpOvZ1Tfjr0jJ0YkWFxgU69wu/4WwtBu0shotS
7syCEMBxek2mJPAivwViX3bXIzei48mBww2CKqK0Rk1qG+ydzwdq59NqaqnPjW9OinSz9dfprOkG
F9etQeVBTIZ0GbPrus0qVKwR6S8WJqKjUn+KIh8fg/aBn+FnXWZpLVgU8UqjgrEW2r1ryFW88zL0
7qOLuMSeNOGfJW0IRGrOHp78Q34V3gJMpMyb1XQz7J/qphKLErFSpcczVQ/Au485V72+mmM5z1zm
pEQtUQ06foWU4eNNIgKCz1d6Rx09jbz37OLeOkXVfAV2QuvWl0Nmmcxnm7Ppo4vMVXFO3tCOHaJF
35Wktizsnpe7axcudJYkQUOZlBsOqFBypYrKU6Hf8Ji9v+8J/LplJd5tcUykKMvHlCkuzgYQsdl3
qTF57hXbjceVMOAQjJD2+QgUe5laa9pMEoUwW2B9hDlGTtk9mojg1JvkxMqV1B3nGf/3uJjuuaVA
CLA9lTcGI6vWQvVQku1ooi+uja+OAK5zK6hlA1vi0AVELKrBVSKmva/ubPq2iRvT6d4bJ233Mim2
WRPi0sRBUTeXK8SqNax9jcxEM3W5uLm1RMf06qi67RkGqM23njLmqR1OPCKeNjz2LXl1/Nn5yWXP
3BaCnsuMBjPujmd4iNL81hVMgnEJp++2Qf5X91rQKCF5eL9fTwcioGk79Q499hbtaCbGwg8bW9NE
945yEmctwt3IW8xd1JEEzqx2ynNY6h/G37Y9euhIN3ZHzvqmkhNRdmdrATXZBQUBxFpAzjhl9EvV
jq8usNCZ+w9Mgu5XkdA0DQ7ycTXnKMD2UdfQDmXo09NReKHzdIkdXLwLloGxkwIDybVh6U7wRWlo
eifJN9fCX53FwAuVYBSs2/yYWZ0AyUUFaN7YRqInfgi/hRJBWYQY89v+KGgb2je8mCB5C4UA5eZB
E1B16pltd9/wWKpmHVsseqr0tznG2smMoNAR5GaFTM0wS18BAAC5bt+CtIQ2OEWUY1ghFmdaJvO4
Cliuf+N3lxKIc7hWOQrv2D1REvYrRreAQcCtSBRMpkcFv5EJyJ1ca6eKcf/QfQ0olPLJI8Ka+sMS
ykGyHon+bjgFEf830ybpFUt0uh63pLhi7ii5SHx9COHFeq6LWlIZlItknHPwyr3mOxK/DuXSx7iU
JfeYGzecklgV6DUnQ9D62XhYZyrkudsqi+hQ1byoRSswqq3wydgmhN1/8imlZkzAyJiZ68/7f4zo
ltZUS0IumHw8FdGbm+3D6IMMFk1CtrE4Sv42Ob8/IKx/0899iXkp6Mk+6W5pVzY+h5JZZZtwcPmS
KsxDCK7xD1KoxP//FRKHRA4NM/RzxjGyjMiKWUgx0krCL8SyLoVpsheMVPPuaU79v9gHnH57OYMk
tjOXH8zR1dkkrDkg3lUfKkvVDFjmuL6FRxZkWuK/fjYiyFTEIyp5jFNwPrq/vxvH0S29eXhq1Dxw
ZATISf4l8og7xY6KdQ7bw9KlF76uOgfWkyvtpM+6iUv26WwaEUN+nt/twb1bOa9ie5nwbEtioZ/X
/wHVxcJvW4UKt+x7UFi/z/36LUaBCbJhkEIz2SrwC5YY9LlPDT6E/nf7beQnGI8ZWDYO/nxHNYFq
/tm9QpjYux20sbk7j9W5IgTm2Fx9CdTju0DJYqUAN4q4EVcaiJQOfeq+nZ6zXrEQ7GHDtzYOyBjf
wgJMQ6OoZ76lpEE5xMq3hege6t+dxa6YSsTwpdrm+e81MibHQkV4FzKO9jCXHle9BKgizseYVto2
0GR6+1se68BR9fJRprmp++J37BfrmNQVoVH8FqN1bJwVtWm1afvYu9Pmi4G5EHF0nuUcRQe8u28P
L3eBO2FdxFTQcD8HNUvAqul1su7Q3B+1oYqEqR7Bo0P4fgXqUC15hoym6PXb0qvHT4RF4ouVrBc8
aCpLXBtOT12Tt20TgYQpcQSCp6n2CqqBJyupPt+DMDwmWIUM4I0VdLKxfTq7h+sQC9CvHSb4fkpi
T4YRjuXRxNF7GNm1YUG46KuOijYSlnOG7VZDLRjTfI82mykpm32Wm4QKu0dg6OSeEuTRv72q77z1
lENc2VX7fQmLDDTXnQBRRP0i0EToViAaPV1eSZFXaY+wfeG47JQXhUwbuyZ6rnPAgF0nL6bw/lqU
L9B83e1S4krlWtVb8Nnn2n2PiH9kXDSY6v8iIb2s4QsXmYAF0vR1DlQcYphRmgF7KjciN3rEAOeb
RgBt9uvmCnByGa7ffECF3224RZBLeRgd4ZYHGKqhG3sLc2J9YEA+u39oymmBc7GuGu/Lv+U1fXys
w57hF9JoR6yRUp3yXwGq3rSnt6te99MsTOnzB7LDK5gDq4gQpWkfaw6qUwMAw/FZwLYv5w85PC5R
RhSMLVpjWx2e6o/iX6WBguu8fAOCCQ7Z3ERnUkw5io8erMacvAwUKVKEleibRMznwy/UOihRsepv
7Ano0VafSz551gCHRKtUHgwNFhZjCVkzyct0/l5WXFxg/Q5EESQ4uz8YSDSssVrVF2gzADG9zXCT
ouFmcowIodUiWZ6lVkKyYGDNT3UKrmYyAQiq16J07QhOKygwNKuftzD6WTieZJG3pyna7KKXKItQ
L7Pnxq1FD6FOcybePrxFPoYJkE3tL74S/FyRepqtwwj3mKaKHpwjcxbrdqlFOuJ79seMhmAInSAi
YpmxLU33WCv7B6Jc0b4EJOyrYa9LarEvoRBpRtRmrZgtNTCiLFKV92f7LJFcpzo9734g8MFXK/2i
afrC42C0ES/3xhsuupe6WQQYnGShS3pc3SBbfbE7Q56RcQOwxcet6dLQUACICqbIpqeeVmurKAmP
rJ5yP+DU185nrAl37EUm8M6EFBGtqNNvS3VRAh5PWSmXP9HktfXM8iyzMvMh7g6/NkVWGDKJaWY5
LN5cueorTxLvrLqRY4vus1COKF2DYyQ1QEu6ClFxgx3UNaA0xGCWWOfR47KoJr7FRssOIAQMtE9m
KoSm3uTFcflzeYEEhpCChk2whd1sUDYjthvivhuPadrsczoh+Gg0NOIsPhDgwzlnbgRoJBucpn+y
TeTBIe71uVon5qCS+Opo7cRh5YZEVe0RsTAx5DH0izC00MqLUBndR80zw2Sbzv6N8mDzP5xdi3Yd
ylxznL2QRBuF8i3yQOAyvSmw21SJgMMNubW67gF/avuUu79HD5e469lL7rSLfI9OAbbzX3M6A8AL
uW7YliY71lxkEFs+AqaHgGS5tVc8Duf4YOVZnHYYYPvhZJDRT1ONG4z3FKbQnIq3Ls3WMhvZ/svk
G995P3vCsjjKnmZPhgeKUn2Sf7bXjOTxNSdBvKDRBpe/UjSk0eBLedkR5bf3xekjk1W07q+v/ZHk
HcnymwsEfeKDVWNcCMgjKLvhVFGb/qR8vc2vQCwvy7/sEeDyB2llbn/UA1L7QABku2k4I8vFiRH9
YHl3avD9W/SxASNzdZz3yj1+RxzqPUfWJqiLEc5GKoGap0L1yu+BzylbUpl8PH1Rr9vJBpRxA+x1
/i43JcvgapSo8s8xTb9VWRYRz2TJC7A3FP2zQSRWNGCa4Dg8H8B9zrndtpK6n6R2VTMi47wn3Xtx
DzC2o79reQjip6VvuC4+zI3zkeXo6A6IKISLWAE9e0TWznOjYAhidtYmCp3NAo1szyTfrMHqcAPt
ngXR/RbdqYEXxIJZ0ZOhBV0Y/vC0udusYi0RAd6yVDFOdD/01dXFyddN8Aa7nJGthjPw3OIUGw2x
s7hnTqkh0+WCYpuwNF4yXq2F5oo+LX8rG5aVIAu3AL+2+jncXzvNhYnIyc6nNIw4qoQBieqS5dpQ
mBay/B52Z6SNWYoUm1BrGoHYtR/vLCYADNjJvRZH6tMMMS3EidQCK16p135Jtp8yYeka6MMVhsYn
T7OsnSONJ/E5g8cfU9pylxMMV5131np9ZuNyMDamJ99L/Z2NaUFRVxm5QMXrT+Fpru+tJxnPEVOb
Ii0UIhQKLHWxw8iman/UKyWdc5uQWcnDPZDdjJ7r9zMCGWYRO4FzA5pqjivg4ImgPkBzrWbcH7cn
sq55Ee/e+xLw4UxLv/kEX5ntdP2na9o8hegBY8LE3yixeWKqlN8KZoBRSZL6ROolEARyQaKV2zz8
f5QCbVlJmkGSZ485Plf8XyQvVQDdk/o3B2xTj2pEi5I6gBoEx7Nagqen61BvgfCumUfg6rXX2SmN
cnTN+bptF6t1luKVoe2uYtw02vodOL9G6ocqxVZn+E5H/UwOQqJZgCfpt6bCY/tOk9jYu2ZwHEGp
ju/HnUW4rBFLsq5Pktkr88yCpCJdOCJCefXFw+b6BAGbZSlEAI8IpkMVv5eBssE/2FWgQ2dP3A3K
BtTR9nU4x6UlBrFL1wcU65zrD4RjwAxV3M0bRXLk7YHu8u4WYGed/QS8oYDQaAE+zFyVZ1JXIZLz
P2FHXV/gjmUi5LtD9+vS/MXpTzb3wWaBrcd97uFlNI52Bhhdc2Jw14GV4OF6t4wBoAIGYII505IS
u6iBCebXEK4Gt7N4+FmgVmeOpspVnswhfuxHVHUyhtJBeSXV2O0ccUck2oeXl7GGygp1NPu3Ca8e
qKWxmYXbYWyM/JRp/fhjLT3BO+Ak3qJxNngWlKXppGgCS5G5oRX2oJlTFtrkxmZTRZZHOVFJ/z1B
pSV25SE2tv/6BtQjfE/3GL3KTf3T1XMhbbpjGVNYnKC/9S6K6dbiM7dak+BlsTFpuOjrLAvcfJ52
GWoLj37hK9CSjYWpby/FcJVZXt30PaUq5M7YzZYcEnMX4wE3wsWii1d0LnORgz6RFqo0iH9U5AxG
XKO4KbNvHCdpSgB9PeodRLk++jzyvxtVxLm0wtxwirUrpk9JgTvPWkIIDrTc3dGGttqbqR17Ml8X
qKLFylFE9F/i2D2E80LtiEzar8X/7lBiX2En3sHTyNrBKB8BKAopy68eywRwxgok0iANVjn0xruU
Pl6K4t0UdQVpw+EAf+QpnaZ0pnDhHwI2jqt+PWlJQQduDtz0a+d2k/ybMBwoKc8vr9WpIch+Jxbk
pZdma+P6Ml6RvPh7zRouSKzMqQnSTJuUuVfUQfax5nQPe4P3dEQZVdUofiQT4F/rnTchXQ7ENToS
6uRF1hnaqujVnUoIu4iLRZGe2FT8gBdpXhouayAkgeGGX8ATNi9jNRkOvzfoto2RGb2h8LCU9kwU
YRPookkMKHD8USKGWfp/JaPW2QPhbU/vZ62m9nK1GcxQjpDIVho741Cur6M1vSIdZxrdrCbg6EZl
XADEcubNwn6JsfGFQXEiZGTXDlv/FofzBo4f2e8kwip9sZBKKPEnnZ8/TFhnZVFTM/ZKylco8lFD
TBCYWLv31MoOj465no2PNFiQ57M2yCX42MAQZ30EQnY4e+H073rTqxMPPcfc5PQ/JWAK9kuMvLC2
+Ov409Ob1BNHcbvq5sjUlu2xjTDVj3SfZYbzNao5ufNCR+VZNfCDt5HP9De3C0w3AA5nBNfbrHgb
KN/S2jiYw6CmhGQP5FXuEWh6VtRaztEqGwJno4ZomqoDfsJBEc1rhiGtbF2y1WeReFQDUShsX2tz
HOSCOrxSV4gnENKaJx1WpTo2hxHgAz1a6cUC13Z4Z4O72eqjMjB3tIa53vyiGwSDWOyCRmXowvtI
NBMe5nEvUjEjRzSCTCotnDqJZ8JXsANdtVB55y2aCXNas69wi5ppT6weDtdxzJNMYvRr68+e7O3R
BHKto8/anVrgiJ3X6++9QYPoVCSG7R2HxCAPNbplqKNTtfCAJXf63/+932dI2WG+o2PVTcTPUizH
x8Dxrlb1iOPGI9HfxdM+/OIdIZXT4t1GF+72LrAr/rGbcYTU8wDDxvYX/sG8vqQjJfU4AQ26GmoZ
r61yR5G8ZQefJM9zog7eWxH/TaCyTODNMxFdMKUuc0J3XetwXeXFA9Q5ZrT+4A4OwmijH/gaYWiZ
Ul/ZKUC6SOYnvcDZdwtngu8j45AvHVYAzBFr+SgtX0om5WQkdsJRvyx5THWwdTOk+ok4pt8Tbrnd
zVSvSXhBpVSaEvXKNo+Jvw41BNiit9S8VHlFavsbhV70jvvSrUE9xGh1g0d7uDjrHWTbQslELD0O
9D+K3iwEjfi4gk9U8So7sW+eeV1Pta7B/2fABfLm6A874RSFtH8VMZd8D24400GceURdrsl1GObu
X8eLeTMMDHfRbbdrDDtrix6F5hEcrFmeGOrH4XptHuULNddedoYUoRHJk8J8vFVKhBoiL3C1g/BG
rfpjP+s0x75HADAb9FyzYQzT/ekob4FBhHOwMY/TiZuV4FNHJeKvRToNgiB42ko5VELRt2ZZbm4S
wiMOIKquqaSqhAe2F250Mp+1lIDM+QcjwLKDFwyFF4IYprtpZa7u7OIw35X8V5rQGIFKLeOkhrVt
rPABBB8AgoP3h0j6ZNCqWECoVGvooXjXWTeUqgMrpz4nroiAr55XSUu5g8m6r6KmTiicC7Tp21Ad
YA95m3MJ3PrIvQF0m+EQ0uEqS1Sj7JLP1c1K9yr1Of7bSswUmYauQLYVPPKyAROFaVM6UiMfzU5C
xHnO70qK0Jm3RY9TvmJ4PN5hPPELdw7leFEspx6HbhbTC9Of0CYFewtd/nPc0jKSWrpU5qKRMee4
g3L0Vo3pOa6MtdmUZhNrHt/SazPgx6cUIK8aQu/gNbfdKgbNyT/Kx5A1LgssZe2V35okJZ2fld4X
/TVSPIcSTKxuHDFXL4gCMoa2AySHvNGp7bDYP8sa6YPr08tlVcHzN+9kEFK+F46Czl1eWkpNjApT
grIF8GE9/HcoFd26JEfmWUJ4j9ASG45e0BZ674uYh9HFhF/2dQnvsfKm7Y1C+1wwudGeNH52oFVV
S/QnRp2MSgouLo5QDeM8cOxsi3FQ1FPD2pzWM6FLL+LjpV+KJEFfQr6qZHso0toB3LvXUWc7fmfs
cMoES+y9ABGaKWOJ1WePapzHGAkeHutkK5QU8scMCEekAznA5kXp6vqbBS8jJSEH7j2buTbUYxEq
8rojlOl6+brAsStnTNBBs3S4fsMc7fTNy79NPFcrkGHBav9lfanwxwotbpwb71FrI+28IzprSKZd
L8QykoaMclDAzjvneKPI+AmlgfNs4sB9/EvKuup9bmKxO/EYqxP9IyVZE+WSNGn6FcBrZn7lr1vE
vWLb1fZXGyp+MCg0V/+e6vmXk63puKQcIAl4aXL+C2xd6hW20HXTspW6AGbvRPY8Gfk1evlN7K7A
2VO6C2GFsyuB8LFEQ7crEv71e++GGm+A6tnuFOLpwn4gvkNI+5j1OYC/zqHqRZFr59EPt3TxD+wh
/qm4/2BOc+QBrSRq9leNPMjQAdko6VZtJ+TUmdh5qnjgQqZW7JHcJalh5oJvt0xvEtNKzhd2S7UM
ll768W8rsMVcdOTlwMukTDbklyoJDyEiuku2YImFhbNP13ZgSR/vhNTSC2PGWd0kkdL68x5Foylr
SQIkk0pJ9XjTI3dMhZOfYRll4i5dDT14oYogG3efY0hMujvs6lZgkZFeJ4cy2wg+Kfnxxs1O9OOr
9GXt2IVUQV9eBLb6h+UjTE7aVBoBCza7+8SxOz1qJ5jHUvhYSufpVkm/85UuW8VBkhYKpAOjkan0
v3/QegufWLchU2Iq4xJX2ekJBT0c6F/PeASFCk2UQNwIhuD/MekcRcOFQPyCWOjOn6zWAfVFbYme
yb6hWDaBKBSz1v6P2kepAC4kQRngzNnqHc6fVa/XAjsZ8TPgT4NQtCrO/Ch368ZvUzrOaAreq2yI
58aHEc2erVaBUV/IuLWCuYfnn5EWiOvAC5G5dfjojUaafRVfvF6AfKraDIsNP0oH39QLoT0JxXkH
1nOGjqv6kyn25EfQlsGjoFXQwnfvm0g30esov/xyE09Z3S61N8Fn/rqpuGPM5RMFTZ8nTOR+BqJ4
qpxNkR7QFM1ceOiY1n41J1VMzPvojN4vlJJaiB40N1MhfixXC0IGVo2VrOGofeVljsfgR9H6aoFD
OSOlFKSU1z0fEAbs3tEPR3XJV7dbaDe6D56dm6C1RdBawXmEFa/qLaWaxXPniA9WormJKnH9b15R
DADMN5Bk15vCUlT/FKGoerJfXCEFhPLwcWei3GpYzxR/0SRPoGqzLuA1YSiD7JfMegy6AOblWpby
wwu5Kj2uBnz8Cfw+wik2V4XFTpExxxolfBVFd99toFdnCbp/B8peNkv77NBYgJar+p+JuG43qAfv
x+9BRQTA5mh5HyZ3argCv216QaYhKW/go7LHkGB1C0ItoVkkx9ekYZQyyySlThnLwLsIrJEbkwsq
9txZ2S56AJzjPu96E8drZDV9SKEwW3Kh4x9PKR1HNFpXTURoSgdmq6XpXwHRiX2slueUP2RErgsc
L59Q/jaT65lKv1csMK7EeYtkXKUrBdNNQv0S0EMOPwN3eb6OqFz7WdUq5vDJ5WugDjMQ8hEjPkjG
FBUWj7t+uyAFU634+gi+SiSmsGvzuwxG/X5K1yL4DynZUa2HpKpr1tm52h17l6HZmBJ4oiqGQ8t7
RLPshduDuEP+1Fi/YrgmR8dHWJGFfAWfatcispd6d+fy4uRqVz3t+U/hIdFjORZDtk9n5jk9G0Mq
nX5n4HCoVxWivOEIhRsS0cLlV8mwvc+mS7L7Pf2HbdZTXCKkvZmp4bO+kDIOYtqfH0jg34WC7QeH
af8q9iDFK4/ml35eK0Jc852ClhAWYpCaAI7rhTwV4+na+PoYI20MiwUvETedpCMH5G42N7wPmpxY
cLmDHUUh2KuKaGbVeqbOS1fxSZrwfYwB1kLVqLAumnsZ2PPxfSIyXmGrAvoKlq7CXPv2nAsux8XC
ORAzCtHnmU4oxZERz1mTSpjWcPIgv/o+GWNW8cR8lD+MMXQbTc2YVnQMJ3xHjMRoT4+64InZRXyE
/KPTjxs6hm8wq7/ajDmlbI3GgzC3mq/zagU5X8BLdUPOG6l0Dm8wZiq1OSSQOh0ZUCK6JfSxgK9C
IuhFuX9l8YQUT0/S1axt1EX3z1QaAte7lnNiYd6nqDYHjDxHTXIr9qmTDn0z0axV1WG80RK1eRdf
cKzMrmIqH9+0TRg1o+iBrWDhla+kYL3FTY0ZmOj28vyd1awGVQXOda0Hp7sLoTisWIS48fH4aF7G
/SjOdo7+g3Kn6CUOsUnQdZEA5XjI9XWWzOS4R73jSld8i9wifP2Moi4NFmZMrraSSNRb2oovulNn
B0ViKTw4w+JVhnAW3cKQExuT7eXKbqIO1HYjH4qWs5vrVg7h4Q9EpHl6ZOTS53ApNOef6qqC5T2g
z7n1CmP5BVJqABYYK1L+ScO6Pir9x1y3Y2/I0i/jjdw3ci7oerX28EOUTTIeFqYtV3TfouOyUDI/
Ut+Mez02aWlOhEnWCtw+9Eo0pqSkmty/js73afi9yqAsWf5aLGdLWEWvIurlD3ivFhDzsyc9iSVJ
EaBCC03XHaaa+Ek5WuwAdd6SRESvM+N9i58dt9BImDF0CwMBv9+O3/zqMdqzvTcJwYaDR22QPFi7
NswBKQ0Ng/kWDcnMI1XKscc3zk1UGPPxs5uLQs3jETk1DgDqTFTfkceQ1RueLEP2wCcwNyDHEG0N
D2dGAQxBv3o1NK5OhM4i8CVM2i1xHA58O5pthp7VruoZO8i/WowCvgUH6UyXoyzTGrFsArKGdYva
EGsBhQ99COIpTdABYpequTXwETVFFk8DF9+aPrjRXgbODsduaVGheAMqQFQou6uaeGW66errKtug
XVkakRC4Gciy8Gawf2RhMMH/Lt1xJ4yNrOReq5VAsBGDYwVqiAJ3Jsg3qY+lPQSH8PwcXrzpM6Uv
pNB1zF/Sj9pnOY3Qzh5ewAYU9M/EVMMb+p5ldPehHMKQgYqbvHgiAawREAx8rs89/4yLyIMxCENj
+ZUIxNr1GqjfGokp1xSSZHyKmaFH/h83S7N9vweWTNk/fTrAPQLzhunzAsX2tP7/LIU+f7ZrIIHE
wCZJK4beqgc57j8wiC7HEHoHH/t2OM120Gyvzngc7UBXR9ku0YilfrE6imnjqicQbOLTwNUkJwjE
VHBoSygrsmTqdGVBU/Xr+XGxFYL89baFEyW8Apa1WL63Rl0xjJPWED5qFs3zfyVZZqCzPia4G4Dc
qi+Rv/Hh1IM+QMJbboII4gfTDfCWpI3loX4NANHCez26yYFaN8wfcUR298a9QB9uketZQaX2z3Dj
i+zCT2Q+aN0Ns8pHwVqj/9QZnvDIuad80auBTLE5sVbfu9YAg4xyJWwbniRI4tgU1+gykHK4+pbI
oVYBFTXf5BCiObaIZMk/ntqVVb5DLJHRtnO6un6EZbzAFvg+6nROiupEmQDBOoodHaSzRd8ijK53
44lXlrt4FG0wpnOlmjM7oPkgk1XoYzFfi9wg3fo0SDq3t+xYEmDvEomWwa1Zbai9GJLjg/HLIXXV
iH2XW9DUULMZfJBoeQKsocrqjwFJ6AkekibihnQCj8xbjt6++jp9islclBzfs0Epetid5Qa848Xm
p8FVl+jEMxN+rA/zlT5LFpO0mIhMN0wse7oP491rtiWCsB92aD4tNBpKydoHJp1ILeMpRFRKnxVF
HLvdAMpqt1q+EWimhU0q1XSm1ZCaCrwxNElNMIKio/66c1npTwLxQQB2O01My/8JVOSyWfZlDXjg
L5JDvhib9PRog8UDnxHip3FjziBb8ioO2Et12oqOofbGl6Cv0wi+AdDRQLqmO4mC7qHY5F+cc399
OKZ64eI7YN2UH8kS8V9VR8k3xyfkUgqeQnPLmnkoKUUltB31jsDZsBaeB+X/19jb/1Zkiuk79VoT
I7NS+kUCvpnhgF71OjT3mVGcp+IHylZN02S+N9yf3WIb1VjXK75V2rw8rPkwgvLzTHKtpTL0+eBS
sLKk2FyfBV7vemU4fjBqRChxbp8F7k5q6t38F2eDGakwLlMZ7c2nqIx0Hk6Nw/K4yffnwenUX9Jh
x+aumwuMWsm/IprjBJcodK37XjYit314vloS4Ujp+FVKCQcWvRgy0pjtQ2hDFWUC+I+nnH9vqkYV
U+qkv33BTtXKJyEcLworLW79PdaracPtoh1fH8ddPVNAJxsDvkuevM8Usv5sLAhawZBazkJIacFA
eYY0dLlgs/6V8Lio/MKphU8ceB7rr98M8/D+lSybE+TMAi98drb9jdYy0P5MLQXz7FoqpIw7UzzU
V4ljglqjZc4EIWLkQmeX6LKYuqVIWnQ40vyU9y8ROeGeMdQaPCf0YJ938i6bj4D+F5mIEpyieAay
BeLRALzZ5Z/LGqXvDjZFD3/uhvJeMKZeAIQadT48hYZ5xNZC8HVMdMTiI98EKNmYiKY+AQ+udmB9
75OPiPdcIQNzua1DMYPNvImc783yYooda27ldd59rHg7jivN5CriFilIdnDDhcW9qU49b7HOroyT
6rnyeMzGC7dAehyMRGOfa6yyh2WWMLz0wsJoCaIJgqjL0raoYeFw5LBHGMa+dgO02LzrSYAAHKYH
zCGdv7RFRae2zsnA34Wh6HTOfd3zouY/aeykOv3QVAQLycXm7xUKDtyVxaeEG+cVW2stFkZAn9Lk
joAFqaiMQOD8wXDtlrcaQoj33OjhH9IGeMKAtEY4ILM0xYKkDGC6kSWb0D5+fKNSBGXNNrrqV3df
RahPD5jndR8/rZPpunR1e1CyeOl7nPNflzsPrms83E7mAcmkwB4OXo/1IA3WyQV937DZttcpgLzz
QC2SqEwhZ1dXs8jqRAYo5JPhF7NYBHzvo9InnAK0mAdtlh+7w0fF5BpKlqWjdYySkxIEW1TX5jpQ
HDL13Oh1lmeG2gYxOXkl4CjcXKtwokO2D5fMVrWlOarbbqjHUFR4pGperY67erWNaUJf2PhZAvQr
+DbjI+Aea8ckfBk3GEKeg5mNZD2DhQQI5CCYrIFm6nCGPdGYh6R9EW0BExkuvkhslL4Usc3toV5w
yYcxz1PdGSCxYjE2IDrAVSHuwc4eB8+0D2IPGDEFdwA2EJ4dqUucyjMmUb87wJmpRMjHDCkAN5a/
wbo+j36KfBlBz0q6mrqPoykbZn/9ae1hYAtTsvIm9hxbDN5OYZbx79axooxyttmIb6Deqrfuiulw
ceQjSzdPkoG69FYHffLQkYi5lZc09kB/lw4qiztQRE0sEmgH6eStUj9BDXZDU/QUv/2coN5k93o8
bFHUrmEolmNcP4r6M0vErBOp8OqF5xifRFFHFFAdaNpF0pR6/X9XGy3g2mnto8sqYWTt+3dUZArp
TlYLnB1zcr1tQjDI8CCzHhmratWAxe9DPNCGG9kRZYnqOXWz4uJZ6lgUYu9bRv6/t3ksMBY9RiJv
ZhdikJVCyjqGKqwaNjyX/Hiu06W3my8olk6bl0ZXjU7t/urhNgkdIpwW/qEnjRI3rf1jl4dKvMU6
LfCvOHoicarDJRoGG9MJY0FqdBBVSBSgPWnU/rIBM03KLfvDn0uMOO+Of7C+NMqgWzbI+WVydvgp
izIMqxQteaklRAu8YodcIgibDYof+64bui2Ytclc9T4ur7rsQxbWS3ZBBB4cIGDf10/kuNn8jWUI
dMrHsqzz92ATz+O8MNP3r+2257VCJBeXLqkQ9BvmjZ/AXoSH7qC9yTn5lO/8nrQyuSa8JOGf/ehJ
LPWWoB9UyWAfkcEiC/Ju8S1ulJ+yMyeYuj5tAaFbRa3RSDv5NtNxqLFFo/y1cKdCZI5kwOtUzrTz
9kSpLb/tGa2zbAMxX/ctCmRMrMCJbK9g/3AO2TKH8QVHrMxVV//dfYMN4Yll2eF+FzQZJeAikguE
afvsSaSAIPyu1R376AJ2gNz/V2qlVNffMIaaK/fDK7OEV0+vyx4XGQDm7lqeiOmun8tvEoqVDAdj
a0FLkjeUIEdOd1dB1ObV2mkdMRmQV1gXbk8Uqx77/iI0pkHB+AxIoQOAemX/Lf15017ByVhNssCf
/q1DLMJZiNCUXQs7sdR4Won/NIIFsR59KxqJcyeGftHgk3sRdawuhpFhMbbsGHOr6C2ndbTqiI53
AHaI38BSaQfOLlh0FqOHaMLW0XALR9t7oiVPoIcf6ogdZEWf6sRqP6mpnjEnk1hBZcXdfJc/APIq
AKPRWl+NBWU2MXaG5CvFvAJkI3QgdPmOUG0T10ZClBX5jh6FnAepbN+BJBeUmYFNQSzGBTVJiNyY
j24kmaW5ZVVyyBGbGvouPreoeRMYOe6yMLfccDGfTGaXcAPjS90eXDINRqlbhY+5q+apL1hrovZH
vsNP2OwyGWxD1CwFhpKeJFiCSyR7alBTmNaF+RDDrBZ3H7FjH0tW4M/IP+l65WweLp1u6hi4swtL
5mcDuVZHgdZDSTRuj1uFK0PDYk/ckQoLVVw7/N5YP4ZbMXmYvPOINUMGnpyC7awTkl79qRJmNegw
OX49w2OZmJT0O5UHLte6BgbQDI5f03F0HMaB9A7m9ICTSe6LFIUgul85DUm5OPO/T2+IFxlAA6wm
oKLDm0WYocjn56FBmyCnyycwG3Sf06wwEvoF9T7VBMSdyzG4Umx67xXTUvzdAB+Pmorl8meTjxmU
85J0wuuGo/sSP1T06Jas3NsL35l/u9IX78PqSgD6iQH0x4PiSnxiZ504Eo28m+aDTzbCCeLtQs2J
QCSFMb8Xvy6smWgqS00cdjJ7+4g2LumVaoAwSXsThjg20X65yurm6JcqVBvIJtuy6CLrW11M6qh8
ww2nEkc8CsvBEhy8RFlmag88mQWzonjeep7Mi1WjwcgeCMMZgy3G84TAZhqp8RPzRAPvEuRcEpaL
RYuSwodqX+Wzi4dTlyTSlhMc4o4aa0uBjS0WuY959r2EigdmywR0KPEmptUtmXAzwqQ0NV2HJ40Y
L2ucWHI00R/BgNWFMaX98aF+9V9k16Zw5GSIqMQGD+g90OiY+Lg6mSLlqqcHeQQJmlC318pAGgt0
SYNab96GsygbzscDVrvztJygsDnVcurnwPoQah6YSDs61rxxBQt4YfcwZpEw1w88Szwry7fi/mow
hD9K9PINlUQpa9ZLlVffjH5/8Aay2uOo6dsJc2TaUvWUN8irGfHnmteKzoVjtJgHIcGJlNNZ4lxy
7cdHNYRi5ySOqwLHlI9ir7JV3o9DneujAx28t4qiUPFWiKtvziDLkPSmK424QCzbhgC1EscN8/3H
yoEeaO5p2XqDOIMfnVMLHu9TAgBaGvA9SCLpsquPpuy2kaE4iVUH9Q0rytHB9imDxyCYlJPxiyoc
re/Req/YHhxdfiTpm3GebX2CHgZcs71R8hcyj+30Bj6LEFvjB3gu5rcXiB/Rfljyg/oGbzPQfazK
j+pmWW0AY6nEML5jUKc+V9C/q+nStcWnOFv8iJpuihu2BXeINr0vx5BjpciGJPuZ1dBHt7cCU/TT
hd1gO36Fp1we2rnrwJ6kp8NFASQ9ab8HfXY9CzvZudJo2DNclePFlMWyzd4mbcKFEZwa8BmBLOjG
De8HmG3HUoFGwNUXjjvXjdKGkrKTtCrbsFOIRPmkK66MQdfFN6M5I/W2Ih9przkKfDl/SS9CDJ50
lgHY5+E3XR6yAIYDoSl3IuunM8xvjZ1L7yTgAbCVDl5wC3KuU72JcT5JUt7Yb2OKPzSwTaH0rZCv
8mqYzSGRUn+DGd14WS1iXAM2I5rUEOvbevh2WKbu0Tr5D8qhxzIwZVMt+MQXkETPDoFGK10E3sMo
iDViIEPv0FcPl9gez04dnTcJ+wJTrEVUGF+SC47D7FyNAwTXa7s5sQ/z6StFp/eCBhNSlprPVrKE
i2BwTAv9UXZY4KrQbZJHvdKatpAEqt5uJExXcoLLPS1VTKdIzd+T2Z+DmCM8qiSYL16xgIr/G3Qv
644Yd3qTfG8NPjtCIRlMK2Oqr+k3BBn7oqVR45fb4H8/DzJVlzOO00BPOEXhEzamS3TjMr6yTaDW
D5RUCEnBcbd4Cm1yZKicWefBu456tiinRdFoPy9JMtQOdV3dWK6NVYURx0W7yVQARo4+o82NOSnU
zFL7vJKBsymvF/I8VxDW67LTciXpQpOm2MF3XPco4Je/o8uOQ/O1Q5K9xNnGGK/ePRtkYg4LAFrj
23LMWIHJMAbNY9gKno8/X4FicvnwOxhfucQyvg0QudNjmMTyTbYIRJfngfxo95GNVHp0uO2CRokp
pqOT/Cl29VeGDGjDKt0mnSNvFt6QswIiyutwI8OYlgK7dVnioNmg2CwQ8YQVPFm6WuTMZMCY7K9I
YJYRjuYaZ+EO89yzo4jFDSUfCDgd9YooEONyxszqD3TqtjYQqC1CSiJR3HkX+D3VebPPJSmX4gGl
bZ8b5HkVNB904tPjQrD5O6MJlUqK7f1oPWDak1AuoNR1DgWFq+m3xbXZsC18PhUht+yRmUqEJ+e3
Fwv4t7Tw/Y6s3bEevl0EibmSe9WyQHlU8n5O5JP3u/fXY1AHOrZeiF6cD9KILBF4ng+ggE3RCBhO
hKFNsNo2ErudW0GFugY0NyToHH/2Nfl4Qx5bNbaKc5FsyZ6pULS1ZPUfYwNfw9vvkEODpWkrpCPY
8WB0kUCZWy2HmvUMDWnMrgOdKrBUhe9RBrG03gjNPKjTBiOyDsggmgiYYbN9EpQZ7AqYQvl9PpS3
gYdFrRMPTMzvOoeZemDW9YVxbHMO8j02/aXg4lxqthp43YzL8N45yNVpC7DH19wBr/KRbBoaWoQm
gehVz6KGEiNyCK44rRk4xtzan0NesRiZ8C8b+6yL5rO99E86FXI1Dnr+nsukIvN9F152kcmMJpAN
nnw7mDjgINbAMtDpA/odHjpsd/0ys1pAP6DqaAtzXp3tgq9LMJxsGe3kkfl4koWDfL+C3vv/LkCE
aKVE0GPpQcpDMdyjS+gDm7/4lo5JBDPunSdKckVZMQwmjspp1gX5IX7JlL8fVRqgfJz/CJLmKF3y
1iYvDzSf1fxLkQFs5BGF88vvb3onV7mhn+MGYYdLyWkuh36ov+73cPqqhJqB4zn/Zm3ewVzEboQN
+80g47qCyoJYGRiycteqDjNbNQYsecnOfnnyuaZEjQa3sqhcB5D6ryPZKJAa8AjRz/+Vd63ZabvJ
aNpJ1UDDQzrAKcisq0IN4uTMP0yL7/bni4SkMzYoBkXDpwQtHL5R+zghzm3GXYhUtJdsNAzjIIAy
a6+mD7Oj+2nIP9GYHLfpvVoCmw3WiqMh/ZlBroBbB6sAXKdjQEuNoItK+J38cnhM+O2cf0GObmTx
DUvNsWWY5YL3Airyy3IboRkxqqxd4OYAWSEo1rL6x15jJ83uq2fOHjsLcvereZe04CGd94GeI0EB
VStTjiJsLOeODIATyfXJGYR73KmNsG9skmXWuJob6zpHqGhhFD71HMB9OsH8jSmtNt/k/EZziv2w
b84ajntIZ8THjUqq5GX7DqS8QMoySU/TvU/r48By0JV89mCwJCWoCZNaPQA5l8rUTPAHX/4keImi
inrjqfC15jIoFFjFzzQHKMWb3nD6GZFG7Bsghf8lf25YYEAJ717ampxMnZJefaIheE3I4ckDOq2s
aOq1CZRFV7LUCOwgecXnlsl790qmjH9g1V5mzMBd+wqXMAAWb/CPO9HeULHiNYZvHkvSRmgEaO9y
y5X/OKVjjnKuujXblHLfEBSwYRPEN7LzPiqiYB5hb0HPBoZS+q1zRgwmju72l2swVdUsg37A7V93
+7MzAtobvMx+7+j/tOMB8ysg6ZlgAEZZRQN4NAyaXZNIt1l+9ZjZtSDnn2VaS0WP3po02I2NjYXl
Wx48/C7lCZbbiMyH4xVCVcFmjReJRjDZY8wx0KI0R80a+z+9rldOXT6mGtCts+TBfL8a3SiZAN0Z
iaZTI3n6mdTNO5x99tfJXZu6QRs6iVjV8caLWQCaudlAU2SGkENflKTLzQcCPCKd40Y1DA0DA+GL
pV+7Ppbh8rayufQfecboNFb5liSZjjRsA/4aEsl6oai8dAsrIWkldUXOf60yAkhtOs1kObNSpXRB
Co2JcOfapmRJE8UBEiSzk44b7qHOkuwlibiGRKATf0aNz9K3RoQ67g9t6JN5RZYhwqK9Me785OP/
458KrFHabc+XOddMiz25epqVGduSNOWbHMJjzSDoQ/R6lZqgjlEarGuOQOg9qAMbhHTsPr00IHd8
qyEGX6O321wNCzRdzI1jLr81HLdpERdQpXGIV+MuydG0wG7bWKpyeFA9uD48r6vU21mXpnaPyL7j
6cCTg1hWgZihZHeQm4OpDyWH97PIndmjWuP8bdudMM8vjrzQdBOIrM90b0gl+flqKDsvlHvRpk0i
kA/ZpjfEcEK5TeaBBGh+B8w07hXfRIanyKZGwCkfDIf3wPGuCcLNNdj8qZx7yur7Lv/kBBcaHoxP
SzzNZkFeRxJg3EN9OKIczKKdVAD+5L4+cbi/XvmFU0LuNhMM252u134oAsCe35gWOL92qQZAEAWu
hV0soXpeM5IGSLo402SvOcQeBai2F33cBSO8FQlWN23Egg1lBFr+ym2iaJ9hpdfUOvouVLDR3NQL
wLiQ90ozPJHA12XHtx0y4Z6ALjMBccPHK5qYjrgONddmgAqikFfZGVZB1YIp+jIq0GXodTJf/1oc
vs8fzKun4kIaqW+wG6mk3RtMqk72PqZGdWPs5JPfEuM3o2KB2tmj8iHnXtYVGwG85m8unBqSbwVa
1buYO+ZouYRCSMdwWBhHqBm2BV5INaRc5dXvQp0Hb4+exmAEbpQVTQULapk45KUOAs6/cao9Q6id
e8N+03miC1ApZku+kBXOfmMZecReD8M9WnTpqXCisnMxWJD/8zQjF3LDi4k5CUy944QAVFOwU/FP
uPBwKBlVomTbvEnDHBTHglhQtWfDwugUB1beJzx9yeAQPCdLvzPSYqCmhJHWgayZVhLNK22evCIc
ZsL/z3LSCqqQm/3p68Q708zZaaLTOEDqH1VbYOv+0U1E2IPqPrz9Vb4J1ZmERC3E6AxfR5tyGDsh
ohxFAMTCY8pkwIoGp/69iF+xhRb61ow4tPy5bQpZecay3GaBtBPCh7RaQBiGMKDIlv2GvUI1a1ct
6gpMum71w8Q4RilF64wX02kiqPk4EqeaIkWbsFZDXw3acZZaJiyMlulAmufYwdgVUBx8Vttdu/u5
7cNRu4HFwirPCar6pRr6br9Mml5tQrC4IAkKvT4vcZYRVvRoAEE55g8mEbk+I4mLec51GsnV7Uk3
dg6Seo7tC2fljytEWvYrQvM/keuvFgdAZ5QujrddJ7PMk1P+CofjnjSrQu2NbDovJHJfiW6mKe7w
zHJITrMSThi9e34VqaBBQ6JJx96DQp9VwLvzMsaL+tXtNYiTaTx3U331FPQOfsvwYVcvF7qEWhJc
g4fpGfgae+xk9vc4XikqgCzR2XnnmxDu4hc1Zj6yCN1Ugx+1X0ikxWOf0Z4eHWB/83x8JVUi0x4F
1m9XLWBqzlz24aOTDjKbo7c/0wm61WpwEa2k+x9MaSBcECaMZ20jK0p3hf0fPLp2SkEwo1MOLIAm
PkwS4N9m0TceRWTqmr4wsK3XyfHmFHEHkIHS+SPETp0v+YEH24Dlll25cq6IBDYDpEuztUW9qnFO
Srb662vUlBluGov8FDtBWM3XOwZ7vfIF38Af4vbnNkkjKl+sPRjcYWGF3IvH+bCfmK7OJQvPmV0R
LmT8u8FX+jqroN7+hAKGXdWwmmqRoV/71pXszqa0qJ9PFtjjccL949XCa8/SYRpHntY+fU/ifzTU
vXLdwsuGLTVqMTBudlCoctAuTTn6DVz2HLSL3GM2Ly3vnY5iN51X/jDfmMU0n/8/cSqH/IdxqYKK
u4yi1xFbrq6k2OOk+xKiO7xyu0AEt7VwHgC9xTtr3KizhunDmeBo+zru6wZL0Dcv/rATQrGUzTF7
7R0G5jjnaK2oRhg4QZcu86eNbbfZcWFKD3T+ENAMbMB+RElhz4od5DeQxCE9o6uZgaUO0uuzjQp3
yFafU5bjDqKs9ewGEz5GK+gDNe+eABAXZpzFDBDJSVO4TMOVU8pGdBwt7XCSLHj34fw0ti3kwTGv
tBai02e76ItLPqwh+CbU5eNuAHc8t+tljpxO1OOgje2xRhB+Lt/VC88FxPoGkfr5ujq8P330CgnG
cLa5zTX1lJEZObyeS17UDwn+PiShvLIbmB1XgaWsIDnZTN66jj5avz6tTqFLRfZDkpyU9x/aEdSt
MHxb2OjTWEuF1MTHeXajGxk78ZkK0FfVOb80KaCMtO9qRacJuGdRSLW11kCbq2EKZX4/Vvhicx3q
isODt/r4tBHTKo85uQCBv11rMx9jT1Aq66o23tRnjmXQmgWVX6We3EKabb9ZC6ffPCj6sWiPtxC+
Ev08vLjlcRjE9JaGXN0W9QkNOZMKWje5mz/SrJIWd7l2sz3acrUOsBQSNdEf+UKKvy4K5z6/24NP
SIY5ktGCKjEra1rZrJvsUG59v+6SpGX1kbfa4FrfqD9PleWOIIu5NX7csSIMXhN5tro2I1aVeVBq
2ZWkhqAuYHxeg9BowyYefuyvJ+upgAmnjQ4zox59EdQa0rbuGumnZ/EhpJFmYum5ZmA1CB9LowXw
X3vLydwh63iyDG+jw6XT45S1PQDGem7Nar2p9Oj63h/zQh7OQcsI+qsIkTcmQ/gjQP0th/1s7VfP
r0lRbzj2YJs+wB9To/o8D7fs+TQ2s/pqYgv0E1qlcs5dadOD0BalTugosUBl2RzM5V72dEYMRqlO
MpDsbuWo0SX270dgLV0CKLu6y4lfKM4foyNtFd/Rs4s1epgwYEejf88IjtIMYSUfOMTTX/F/IS5s
AKUCbaA1056YLQGZXxExg9L7OUo4HeE2/YZB4FCSR3GckqcGJi8cHSW1ismACzBbV0i0WiY7LKir
E/y9bmQVfGcFjseY7GMAgOdFLlZpeibF58HVVNlI5Ooy71m3xM+x3W2HOETIDRHIyyHUU0ZI6Lng
1l16wyG7wchagRprPeuP08olpmHGxIYQqLR5cpAPgiqE+Rwr+xekOnMTuM5JuHdyfFD+P7pCnyPz
0jTrKDSza2DXoO1ddlRSUOJU1T84U49Mobylx4KpuGXDi4PQUozVkFZOSeOvddK5TFcWSGZpl/AC
L0sTf3C9oJzwxqoWDCG6gbhg87IC64DQnEFUPwT+JflReSZuGSs+n8CwxPmcqrHyUOh9RSlBtwFj
KVO6L6qtY5Y9xSQMO3I731rFNxqhAdDg79Vldz9J2/uxiIBzxV9smZQifSDC30cGT1zRANGi3864
22ttGsnxBDP2C1UuyZdkH1PU/SqQGu3l58wicz1mks2q0I9pzIhunzimrS1MJSEkQGmjS+Vbql4y
CCfIbudSBuk3/YI24eAa+8BK5SQB5jGDmHiuFPFBXhs9VbYV/chNLZjyiqt8NutBkke26YUARvkf
mZ0FaBC0Hvl5X1JWta/vrfTNuWP6WIb+WhNgmlFA426QDv5x9EysP1dFwBl+ckVE88MLmQR2/l4M
58yjDIa1iyJaRwKz0B+7xzIMeVH3F6iawv4/gUV7+nZRFj5ISX4ConvIl7bBahohTyTZo1y752QP
2zEoS+PohQA3HdRHqSGx+hrI60zP2dYuXSsDJOqCNburV9zgNyPrITN4CYZyujqs7W3FJMEB+lba
5K0hT/9DWkSenftjUwzo0ZFsSKUIDzBBGbO7UhW+6ykcJtbY1/NE0mOZP5HSbv62J9Qbh7otklMn
/dvmcDMIMkB5P+Uippqf2wmZbybYOz0d+a46cZkv0iDCStKAnot7EHgDbIGSGTE21KGH9NmJugkQ
LCsvkiMP0Jk86EQrKSW8LDBFTQYZMeiWq05eZ94A2qsf8HuE8gtPL6Aw6KEs2b+IObZsyTtom4ix
cKnmhxwn5QpllZDEVHAwdyDWBhjWkv5BCnKxN7ix6O+LWCpa3kR3TQvEjFjUi1zaT1RLRbXJDHD8
2xV7JpIhJheHirRgzyieeyP9/gHpMviI4U90VtVrWtLAD7GO5H1cUyCSf9ke1wSsLxMm0dM5h5NC
/xEevuK3X544MtjRRmKEzsJB+Q0uMAThfcEE2pJmW664BxD1jF77zP5IxTcG1CU1Uqdd9ui8S/Lk
YHRULMz/E+FGeeltQe8y94vlqELsBgQ+OIpj7YPW8JrcZGkpDggZ7cugGr51ktVg3Oxb/Xnpvq17
ZZNDlcesgtrbqA4CNc8z144T5+yu02ENaoUDMixeIfWBVD+yiMAvqgTKopEJIlUCZ6/KwO6jW0sO
MtilG0ZbSHQNsYFnGO9hwRjELEojXVvI4tX7SRhx9qHCy3cIiAUhtlKr2d7kO343pG1wjVGMSRxs
lcTuXwsEjRjx3c+QIECmXnhdp4AZXTrmcSua930b0wP8MhySl7fv78kiF86srPf+xh0WhivqREnV
Y0I3J2GklXBWhCFRqDinNKnP90/Dj3CbCBIXOv6V2k1vcw3sdhuxLUv92uMXFTCa3k9SoUGeYUA7
AL0GKI1yS6ZYL/X0/c7X8a6q7UuJ8LtPq8XW+skwQ8qoghO/elDrP7huq6UQegMZQ4Da77j8avG7
3zjBoIu+9mSpw8EXkdWBzEk5p4KT00ebTmvu7hsR6JpzKnmGhcWWZZ+8VfBQCY8jUGWzBaDuqYH8
U34wRSMNxzUppsZTmtEuOrTFUarLaHGSqIUWfxiiVU7rsclYlSSyGkF0Paq8r/a+vV1PJVhsCFs3
OTz7o0TqJFyVlZ85jFyr7nh578zqZzxR21ZFQ2gtclx1qbGT0O+1ohpTTNGmID3syjMREXnsu8pm
zU4LMTNLdEnXr26oWcML8gfSy3pXyoX0/JK8wfvNY080x4xdSBMop6cj/+u7m0HOw+hkboZM3Ikx
PvLtNBPryDIuJZOvrz2T+VLBJxSLxBA+9cBOwM+7Agr2kGkYUsNN9GiM+PnqrAdLaGB5Ml7u0TiJ
OuKC+uIDzvZIqGpn3qe5Uz1hFFK4bhj1wmSbuz9jrbrduihwhx8J2nYnFYEzFSVBsHcne4yo1R/I
j/ZfHj248V9jepUIMmIbM1rr8NljpPkUbZ5hYS/jKGFpg7nnGhO5u8WGvHCCe+cJ6iOA7894Hr0+
irzJ61+6k3AwkJI2EWfLFIQ9ELNw16Ka44dp1Jf6YCrluYTW0Fk6dq27wj8S8G+5MPEbpaL8QEvP
4f7VbCLHMbByxkEnCkJig+oQvYjzLAoVkbZfpb0oJRc8tmgLtwaMeQLZNS905qhLmvLsVg6mUdxD
sGH6yxcJMpcyxp1Lf/nsdXdGrILuImXa3FNvKbTgh2vKY1uhlmTDFeTXfcCcV1sVL0hz7ykNqV4b
xz5HgHdmG9IQfpbMkKY124rEV7JVd+blCpoAqngD+3kLmAP8y2TLikCF2X5oKH7RAS6ODmSXCE/8
DxRiJ96ZrXnMzWJBtiRl3BUHaNAoCxq/TzKD2YbGbYr4Qytnl0JhoJt6eLCNGPVsz1mh9DJW+5T/
i/AxHA9nSDNpBfneV6KLKX5qL4HQJhNnorSHNWb+xGeXoL1Z1nrg/2Cegfrbcc3wOeiXFrrmUOLV
5OxSgFud+IgvKgOULL1tLIV5/iKVy8yRY3jnT0jMLygiqYqtzLFcLaPT0lE9+w2Io/l++zz4X9Vs
bKkxPX6qZ51FptKgaaCgyfzxvFPP1fJPzm7EIkdZbzTRcxJl92L/dqXmIs8Jp405yap0Mob/S0FP
yC+gKWxZcmorTi4TbDogldVK1btKkM8Z9S/OP4TXPzfr5XsL6tLwln17aMer0VnstpK9+nzfQT3j
9NqaOsA84916WL9eO4XHpDcEzQuxt0YCROiJrhYwSv+9P41NoHGt5u7wSLnP8lD/BB5bikCH/pFg
AYolJ6uQP3aygBMHMPoZBer/iQryk+QXsNwOnq8Pf1BSkltTAlbQcGW6VuFViEzF1ubS8N0R2U15
z0PxjhNbi2YiwSTMv8oduibDHGACCv/FoDx44rIA4XSUlGYuKW2DUpDnOQUdHvevXoRaAvVERmBJ
WORaCvQE4kHZDxWcH+XeUke2rxKjw8p9rq+2uTxfW8JEBvrkEjt3CI4+Va6rHCYvpyGXpFE3caVR
qspo3urcoNxZQd1ADKEUjiiAOcir+kx7fCEOk1nrDDzmphao+8y30h9EC8N8X4Tl2+QSJBSiZwaI
Xbvy1LBlYwy4wWW/ZrHRz2rKdc0fujOzF900Xy6YzGwzdNJ2sgNC1NOyGFc4VW7+Kdk7CEpGhR6n
voMw+iniN6LQUksL5HSUjulmvIzhs0LXa+DjnPaLVA1T9j/w/dsAjXHyIUHyqHqYX2M43PnhumXK
VRw0mUJKkJkjvdQHrsYcMJ42c6P5rkVKP4HfYVTNdYLrhfkdzTY/ON0gLoC+DDWaXcrepyyLIGf4
BN9UOmEu8qvrnt9YHuN8jrMRSezAN5bngRdqyl3Poh2xaU6td9X9tCv3B3I6wZ4g/oDpXuPqxjoy
AKUNQC8POYWRxKJ7ShfP/RtSmm+OnSV/AIrtEK9r4SfEdbHQpqzByTwqKamWwZ4NH6DJlZ7nEFcs
6uAI1J6cOpWPqh/RngUk6ISic1RUM+QXHLBqA0Shw06cegpgLcq1ZlPaRX5v6QP5zSpJBwUZLyAm
04h3tC6W3N5KYy+lVw8QAiwx8meCr3et2ghVXikiyyr4bkgLNz59Qq4LUbOCckxB2uN3SPmskJSW
NrkoRNJhgoaiDtszcbpHu/xkRSX5EM/2321XJMf14eJuf7rj88vYRle44y3/QVoQWWhxFyMyrwuU
yc/tmy8j3OfcmHAjmdQg99fn7b2p1z0HSB1LntNyJFon3QhsCurrO4c4Hq1wYE1+lK7xiDR0JxmT
4rGKG3vwJEl7d06rLN7UD6cGmMykQAviS8NtYSU270JH5qojN9lgbWHWK+xYl/8XYKztlj7Aymqw
s9ZzAWUlsviN8ZISLPITUREzsF1BbGnfffa6WTKv04SAAZ4xI06jmbYdGLgJ0jY8s6d6MUKKc780
NG1so3IeZ1QMcB0meDcjnl2XJuphVN1j4LOVBG7i3x36R0qzMans7jWJuu2z7090CkNh6RN5Otfa
tVg6DwtvOzbvGRzispZZyvvxKadlbffnI8vhjIC5Q8uz5oF+QH6j/K+QynbhBth6cwJrVzb0lr5A
uy+qvi4NoVB7x/bpFdIzy7gvfReSo7TLO/m8O/f+X8A7jr2x2IitveFD7raEZQrqkeq/VGH0IVOW
kKm2xotHfaQr8AZ5evXdMm9Rx9AdIFM7Ws9oHzmVsruDeMeNeRsj0IJ/WfgIXwfLlxwyq9TZ0uoA
UfS8IZ9fEO7UpWCawkqryqHVQ2C++RXSE1NqW2bPm67mOxePD0NJ+VInqIG9A9DjLYPq1Ntzp13f
QqfKR9J0ztP2VPc1js7nl8RaxVLHbBgrXQ+Ruz7w6uOJLZeQsvdxc6XdnYju6f8GhUzbcw4jBNMv
uTTQ4NlgB8CBqe54Tg64213B46pUmCPH30Q7A/JaFHbXpnzXCRL/KXJbu4991uNyegD41ybmtBpY
C/ScLL5H1pXt9t2cgwJKK5ej8bnrljULdRPLaQr+D1IzLQJV9r68z1szGx7wq1uav/koBBUhQUFY
fkNLZWqIsfdFyFPARhclZZmxA3wIB6d+zqb3MKjHLKv+PTr/eIPsK1jNP0ohi/BNRB8iqdGk5NZ5
UjjS+NAD/k/OyLj26B0e+VDu1QqPXPemJACzviFFaqsfXXwNwqmwxFKsYBLTjhhqC+6tH1pe1XTT
ILdYgvm9qJBMp4v/mBta2wxXvhBxiBcNJaXBtI1iIQ1WfcjapdVvPpyfwQC4ZvhhzxeTCGMunpRL
eF+2UrTWOQUrPPLsZwxN6H6o9OX5536fsVWJpq1BjXVF7Hcq3LNc61HAfPP1OwW5TWPSl7jlcOsu
/9fBOqYhwzs63qSTB9scRq2ry2R2lwWJGLGSs/qxoOso8+4dMbqzAYXTANou/YY0rM6AL4bHH7aP
J0kEP0TUCHC0CO13283RYkgnYrX404tEaa7XlLg3gmYEZVgOkUpVkkRTX4y9AC1F6OQFCjIt1DuB
DRKKa8HNl11hmQkHFG+w5k1YZhIRbF/hPy+I2VvsPSLDI/EiJl8pOXcqeY76DmjOMB9VqqYBXDBz
9gtzgojYQEP1H9FKyAn6bqGDk5o433uNsgf3eVlpJvW+sjyKxFndujTrGoXZG0Nqa1lvESr7kmeR
xDRmha9JlSEBXu1+2163lfKT9vO/plz172yECijm5XV08sl5zuANxARzuZF6DP46GWyQKmDb3OYG
HlInmNVyHPv3oXK6yMc9XpL9G7a6a+i8BEKDzpJWdLmvj3+8Zu9dHhvbHDjpa9QJDLhpzw0kbx+e
Geb/MoXIomINx3lk/iJhempuINdYazGjQqYpblrB8Ms+FrLNf0Kw0hbtUYimVuNPjhCY02ZZkk6J
RsIXLdkGzsWKY7rkUdn+7fkMoz+c1vpGJYlrnCv2JCEj2vBnfe9SltirO0+EgmRj9OYTs2ov2A/V
qkHzl7xJFwhan6qsi5jcFfugaVzwb0WBtw59prfHITz3lo48SSs9jy3dN3DkivzejTgS2uNrKmoe
3aS7vjuVLn3oQbHSpAzS7IoU4Yib+0CmgjRAQYXm297G6IelB5NFHki73piWd2RgEHtDd/ux/B29
cGUILpXqqqtKSPWT8lu/aq6eXFM8bKGYSQ9a6zWwxgfUN1iKvRjXSsyLaaD8rn+7NtGNWq/HuI7O
49yY0kHq5Fmjakabtr9n2JwvjjIN0vKDYyEwnV1V2waPuG+9N2IBIMdKDNJrcn1ODvwu8DJn71+h
gUrfOQGQP/HFKSuwPisfBg/stBfi1miSQcwyIvszH9CR3Ht/I/9u5wxTdLDPcsjOHO5XXf0Yi3Q+
fh58rvBGxbirGmq8wwikXtHhV8OsdAxO7kdAjI49vU702dyRuTA7mCt4otKRRdgATwpjNvkbUqQE
WVFCQEO8ydfejfzdNWcP/ivhHqniicDuYR21SS9VpxOseNTpdoY8wRUzjNNKnZgTctW8JCUtLFMO
2ipYEAjThjO8k2CldZ+J7WIzSPBCmQtYKOByiDSl4wTKDnYSpSlVICBqcwTU22WO+9efh0S7Q6G+
X7D0/xjnXj0z8MRAHtqdMRkT1PD8kwgLbSxAAOTrSPw3MmReysY8zJiZtI+fwGeCih3j9g8u+U3c
oAHYBkJVSwhGvUXhMcFH2m1XYWwUbTI4kH8jlMCDznXwD3BSCTKEQchbSBNQtqZ47JAavD8UvQq2
vNI+tr4omQta3puxabpHKTvLxjrTQXugYc67ZpHr4HTSgyK87s6ckmakxFj2zmKYlvg+Z+39lrHd
AMjWXweSLWCrGDKhARIsDQBOS8Q9U5hPGWdXGtA0m/4CD9xq9bjlKGNnFHNWwfg5haQ5A/ymD7U5
Lr9tkv7tQStRrxTafnb58712AQVPW/WIqcbZU5r+2uCjFUNpiy272RFIaybvANCxqKJ0KH8QIDs3
JrZiTVJv6s6x9beFxT9S/FPXtHURlgOVCvUJA230t8xJ1T+k1xG81HvJxu+MBI83RwwgptvGChBG
q7h8jL64HCs8uO/dfaYECLSn8GhOwyQEsreCrj0KTcdcjDbHJ8n7aNx7JlYYijr1Ju4mW+Mj+ndN
THSyRdpGAO1Gv+2K1QZLseTqRfTfXzxYGW9m2LHQ/rr48citzfXrBm20SshJCvYkL6aRBmXJylqe
d1UHUSF2oBem7yLFOcq5jlAMin9F109m355QO2IOYCyikpYaEy1TpVCuK9BGvTy1O8ZibAvnRZ8i
WwmSn2DtGWid9KKbafEFo55Em7VUKiQnOS2SQq56ORbSa16PKRVOV9NPqQtBMUYAfAFb9ueb6Xzn
stuX1VOkh09aIwa/C5ks8XsIIXoRL6IEpkImZxvIV6Ln/Im7Wdbd+M6SMZ/2baVfvCf5zPuxvDDs
Sv5ZY4pksKs42dAvRUtR0yoMvObgQu5v65YzpEyUbUySUaa6vHYuf0HYdNxsD2l8lAHPWyRKYsIe
Ljah3kV+ks5tWbFEGzDF2S+gVIiXN2XqkkoJSV+v36rAacbZGatTM2JaMfF+6V/gs0UjdAiyElZl
YNmE66bNDhS2LPdjvq4CsOa3SAp6C4gJAyPsfeuM8hz/TQ6g89+WdSYldfehJUzCpPLuH3zWroBN
OfuSpQ0VojATBjS4DyABYa/PH+N3s3S9k5GdtQJIL5ddlEv/QwtUrmyQQVPu7Q1LjOFybcrmzrY2
1v0T+rzZ10022mrMIRbIbsYkB0GQ86MRkpMZEpaYHOWBokiuq1Dc2Qoy4Zeuw2GGLtAw/wa7F1Zh
jrLpY+2iIj7We61pMVHx0JnEpj7bIcI88jI4TcDW9CLso+rul5FL7DQX723nQ9KWazKyHw4Dxx+h
6eCd1XBNW7KzBe2d6fYvnyoqfQiXKbKoltOHa+da7qAOjCC6+bGX8VNHNhlpwBFTRLpchDQ+aBXU
sYckReHudyxoUEdyuIyujISxVX0RQXXlSd5aR8qXpXAuDTUMounJi4q6GuA5NHypb8+k8uFHNBlA
vRUOCo4QQMbg8WDnc+nvzMsD8slAk22GlJE/bwNcrOupPR1+UjfYz82djltoA1+0u9yIM/euOp82
E3zw5kVcaVWgnsW9ieFf32wFAsV6H69sWxLPxFLSm40zsIu8DVA9uVViciNZ3VaAGx8OzN2BEFSv
Ki2STdWKYyymQbaxSVPUjPVBvfu1psrLCnwhfohIyklJBr3FekbeflbBg527IO24BZrxVQK0nFgy
ZjLW/CSmWouruwT5jGm8GrPxjok3rJnGrcQrYPqBhsocPSrzZAqo5BCzcv5vt52bqk5D3rAfVpJq
QkeSAUTyxrWg5CPOqoLv7a3s5xtOsvc3yAHllsvUXPGHFQgq/dyU8/ptbkxd3P7R4VdIHXx/2Ktf
j+mg6102KJBWk/2dvC9yYow+tzvEOdAO3TlvMmbywpqPgP2Mu8g5boKh764aWVuKY9BQ7fHHPXSF
agvL6ByNah7NTbEItKzFfBr96iAb6fhuw6HGd0sxU5tjvj4+sgvlk9+GYwdIsZkoCNPXyX2nnuPy
IPX6KGiN8lNz9wm6SXa/Cpv59DGqYA4TUjFVASUQQwqViYG3x8bLXQuslPfHiqaLwt1CT4h1i2AR
YK4Qdy0aFGZMKb/E8d9ONk5+Pg5W3BlwK/KzkOYFPn34JuAYPgZkJiC4D3pwUScRQSvYHJq9fv+j
glEStnA2OAnPrakDkiw69JwGWiwmlqa0V3DRhsVnQ4GnfP7XqDGmgBJfbEMoMQyIUh6QcDrKjnQa
5JGeUWibbPcNoarotMcWNC3etUfGdo8mvVek5eMu66Z8gi7bxriz0uca6wTj7dcb+sF7OlAaFxQ9
1HeEyPekVO2OV5N4/FlOXR4TFiKhkxEulKeHs3M+jL6G+BoGEO5ir5lo+3DWQakzF1J7kr0w9NSc
WIIDTSL3ndHr65varlfGT/ssiSi0Aa7Uv7Vf1r8woqeUarVDuTkF/YZgPo1Fr63ROk8MW5noj7EC
21shgy28oPzECG01y5lEF49eh/0aDHKdEQrLClFOY4W1zFisRw9NXwev5OTFi0U4uCPSyi1m3atr
mlliZe4G3ia0uA8E42hzsNk9wlss50E5BFzEojKVHdoMSv636e2cd/pcqrxW6RBmfGuN/sMXy7++
4stBYKuvq6DoSiRKjnqCeQk87IqJ8zGgUO/RrcxlmU8OzPt7l1Q0/xJt/2kJb9Qpy21BFXhjKPik
DFTnerI4cS07APwPPT2cQZrFFePKp+xrDF4tSL1GDuq730iFzmS/9CCNCZ8wjJRGHItsxxljr3Z8
CSpljAL+Flb3mF7dZfUFI55b4vjFpdBduRGTVxQlHfDhnUzBoCv2tVUXXWMZcXpJGw/KGi3h4u2r
BgN+C5VRzr1ZmVRPNJlM+4UIvaLZ8L5YmzAGDNpulhbfewrLFqxy3BVOg0cijSCskv/fh6ALLPcm
Q6z2XLXoeOIgghPkeFWj2DK9yr0UBt7GVTd0cdjGxRe2dZ6MON2ILdXCLtTxn7QhKoHmB4iLxbg4
8YqEIzpZRduqzFCSIsYbD5koMBOInqu9LScBH2gxwCHCVVxGWWrIOqp0xGG5bQvnZtJ9w/pL11G7
+jjRcvXA0xYWsTrCvQnDM6eXPeI5UiDoAThlIkpPK1tyNEDiEcjXnG4pT+RcG85KCTDu9z6PmWU9
KsQ9J3fVL0qaB4xDdikAsHD4I29W4aoMolwIAzevFqB+/49qJohTMwty0n/d3/AtmbWmStDsFKR3
a5I2fsTPuMbsbip5YgkSAWyQBgcGemt2WrGNQsbfHVqUT5uw+sARaCKyfCwnDjeLkF56KF8fX6TY
NhrCqbSLTG2N9RMEjnnI6p+QkLZVUlLXGEhloko/izstcgEH0Bm0iIJnVFDkhcYnAZu/7sAsBYQb
bPLrt+ivWRdsrdconinaTP9tqba3BOu92iw/k4pGPTiwilEX6ZaZRNvM68iOobJ16YP97HvoZCWa
f5CGMYzddprpdCVL/A2qvcovaB3MHDUTlTxOpPBIc6VKcn8nuRaq1ceoCPAe+HCxNaurJICmlSBM
WJCH3GR79VR67b+NBZuIXHKCMFVrwGkTGbdmt9oI56vdVvGnWUXFDhIqYafbHsbzaZbm/vhmHWTP
Jkg+YVlc1qSE5KsP6kKXBDrG7givXHdGnZZ8Yt1zGO1Zp4HIY9rYV/B8RsmL1+JAKEOdQ/lueJ4j
x6tCTN72716/J/lqKXH6/pUejhQ4RFf1UwDCWB4xPYsDp59LVDTAV43TyLU5y+z+5v638AUzn1Z4
G1M0zuTFyWG8f9LhGNJRNQPbljaqTVlEqEvg1S3Vt4bmSpLX57eiMmqjZOfIhdG5tE/ecM/xFk72
aDz/craSXPI6ecthuYmV2FTrDbDu7jGIoN3YbznJrRTOM+mfzfS0EocvecKCaVpANTCt6uZ8f6vP
ty4/sP4404akmf6xJ+8ODSOprTbkUVdnCZ3rlx597e2UVcpO2hPSJE6YONF5Oe/8i4LytUcDG/NW
IeRxC0xwE6q1B8Jqvjpx1TlrEINfsU3pGOanIzUv+SPme1sXEswUFcYtpfjIDGdEhMPcKuETSRph
Vm/FibSxj2YCW+UaFoIvCVBV5DWjeyQ7G2iB52ThJbbxMyz1RzHboUObx/caCmrwWNKXirtLZRcw
MxoL4tltAFNNprk6C6cMeITs2cylM39Pq6UL2X2s5FslkWpEr8V+SgimTv9mAanT+D3zXt3nKGhJ
b/q8n4n/H9slCm6tRdXD0F0Y04XMP+4MIB5t9KtlWrmPP9RrDMKubwaKfFuOjHoa8ndUrx5yICR3
mxwoKUP4vRPPr/Ra/psX/DEB/S676OSyH67AbcURswoQqxSO0Nnw6bcDs/+zpx0+TeKNWmC50v6W
MVUNKr4ujLUw9PUmW1V/NvrL2KVMCkYxQnK90U/MyqfV2ByDq/lTo8/FPZ1PzuEJ/2GWtX8MqeoQ
ddr1rjtMfBy8jqdPtQb8aIxeSta4x2lQRa2hnoh2Xx3Z3aR77N9TSBk+lri6bqgxcuUS3qmIZJMn
L0qkaREsmzdJ39XxeCN5VH6AlWQfNOS8qYgDyngmzPvVnTqiUkvR+WiElkfW7PsYPX0+btvPjcXW
UTVMALhCuxGWBfGMbtOULL5AwKxvYIdpYP04NGiPnE1dfNfRaSbQuD0gKCL3uScJrr2m2WfwLLVV
GO9pWKkWi4FVg/2XihHiq93xNxVNAhMR+VfOnd31N+QeXLq6Zv1E2fWrDinPxcr7UYLS+UF4ISmM
5wVM7OyQuFUYO/yvdNcZ4K9/ZtboFC0vqZgdVv4KDlsn1YwSc411qSNCHhj0kCCddtudKs+5y2tW
+iElRxYOqyC4LqWCTgJP0DA/x7zeMv5Yuy1cK1sQXiyKhMsbdQnUBqbyli9OPa3O4ai8nYLYSFyL
5lHRZAohUjnaTGQG9EmOQ3yKCf4QPzp+/EvI9c/EW1P5AhA6e8KKPP50nw9CUjlYiYrCKnSSgQ71
bw8UXAkAH+S1n4SngQfnU+COBMIL3LZ9nFnz1SHH6Yvrjfq5QsRZtWAO8b5sHC05O8fX7pvY17CJ
Nq8yT9UtQE9O92J4xPSYG7kT9xoED57ASPR9cmSofiXT3+68jfEaTH4LfvLLp6jbMlW2qBB6cOFV
GtYUcwHYWwTsVkT2VjH66SZ64n4IX1JAn3AC11SperiTxWrHDJF9N6XjUNY9HOEuDmjIJAAunKL9
/CHh4gLcW7ZWUdgGXe/KqMgh4yXqlfz3XtExfe4GBDz/qcRkXBGICbrzVGpl4sgv/XBSIB7SN0/w
3aK6Z581Nb0ZjnXXbt3jYsk2VXRS0EZxz6aohW7aHHx77EnzTVCHCX3AbzR9XD1L5b7NxHrDYApx
64rOykxdDBr4CKJ7hBGAVHjt9QBLV7fC2t9LIzT88lAIJWHzD57FwFMdc2/pJtiq2sOalfY3jTc+
YTSWLPy55iBprK+CfV6yD4fFW9/gHU5cR0tu8bhlT6pnEsOKRtjK0CbQx+Dn/Xs8B4thtUZTHSpj
0G+YnPv1MJ+xzWPN6bqEWUJD1l0e9I2clz4VzwBCW4cVLI1T9ap4MFJ6meU3t8tiPiDUFbSmARqM
Nw9mRtgZXOwOZzrdPy3qv4+wlbdZp6yOHnr1TenkrN6ON7gN6WVPj6byEOKToBDZ4RT/+LKZcRpZ
VqEFKx9PopuxSNpRFqZ4F40wLtxakjkdU8Of+4RhwFjRJXcigRrFfXkW6N3WmNCpkD+NtTDZmDn5
e6skeX/PZsUbVcxjxzWaHoiwbzauEf/pck4jZQyt+2e70THhLrQV0D17vRmNsXcZEWFmvYmRDbSi
Aph/hnbs1DF4Rlh2H676Fq6ka/PhZsxPFjtNuhWjnpGli/TxeFHyLVnN/3Bqw6/+rFug/234POiG
PTw19S5vbrQuOAp7hycgvUJnVxsShXwjYOG9tCHXuyqDwRWBoqOqbpIoclKLEdyCoyPacd1ykhBC
zkrPTRi+H5sQXXUcMcuLWhfxFPys3f5Z2dr9dSKyHSgi3whrGYzFrMZT16NFct/TUE+F5yZNgXcS
l65VyHAecR1umtcu9u0DDxSh5kp8Wnthhsez0TzaXctJQ5BtfjsJ1MD+KJO3Sh1IHddwjIi+vFd8
a3e1MJocp9kMcBbBgOIPejcRAbE5lJlWVu8w3XYTFW+hjyWCU9MwQAxZLb5zkMQv//vUcQ1FfUJb
5K96bh05VyliCK2XpoWOUSXrje+EpgWTi7VgR/KBqs8ZQceh7k6zvwZjRSyDDDJdbEYcm5ytAk6y
O2uYxcQWo9a3wGsPao35zTC30tAbi9S0YryY09hyqzVTyW7SjoC5vNp0Thr9rTrn3ILL+54YJcdu
Ckma84bZXvVHD55gl/VLxl/vmuoOHXWSqQQrrRNMTuaKSlte4CCUfQ4Q1HPOQjArhxliPpee+DEX
yddtbsDLm0Fj/WePjBOzadtW/g0OqMoms8D5qG392GFmJOlpuDCLpQrpWTQHx/TjfVNoPbSp/6lq
Ae+upEcPdtAkfq0pITFIrgCjqEc3JVKjZ5TLrpsthaU5XzojdtE/BPKNfbUjI2uTEoPaGvLfqeEf
LdzE3a9GPP7oIzFysWfvoNRrvwOkIFmR9fSwv1Z45m171IBJ0pmmSn3+M1tnjQxearkItYg9UFd7
ZtoaZGDY8hTfkcM0tpaxU+Xd6InpO7doV5gTIVNkH4kIXefu4jTEcnFKaTKgxP4UL9dmnkj413wD
6UATvVAzGE2D4Ym36Aj/E1rdo3jaIFBbrdM4/u6lZlk7fh8JxxQaNm2ZVWbVKymhymv1wymINv37
dxwPh+QukXYZjZsyGfk31/Nyk+pKy7fVkSIitlwLZXDXUEi9if/+R+irVNBMpNXyABoW7a2sJu5r
XI2/cxEihnEnvE8I53W3aUT8UYIyrU4nlEs5hpEtUANW4qyucIpUrDl+N1pzBcBi2sdOM7cuwXiT
QLivlBS2+lzR0ztgEb8NNE7XPgeD79UQ8nmLoeGWST1BvBrpEXtkBmLROHJ+Ma2kiPh6yaUBwUx8
GWOPu6KyMW0eQowxeVq9enbyWn7mJQX/evKIu/HuwCFLGgkGcFmd1wcb9vOSULqSx4x8bZWYa4uX
c6peRy32RXrq0ula4aBcEdqzx+wRn+UBozYkJIiWCt+fhUnadvgb70HurY2ByP/9JIlFXLr5be96
jp7BafllWdd7dh8Ud9lvC5lQynJMXTgfnBiulrjcNjgfKBjmqRDrR6OZgIuO5hfLNygizHM821Sl
L0i7bfPsMZZ68uFKHota/URJHymQzL3rfctscyoa8O5yLnN3HtV3W+lf1kdwclQ50rAnFyHrzpof
ZTqBLjJ77ytb5zHYZO6QoAPjoYuS9vvQdgYiWy2xvMtjk+CH1H4gGxz79tOXcvPT9I+T3oPClkxO
jXCN8cc77PdtzPj8PYptZWcYdXeWbpdneox7daWSsoS0EBx0THSRG4M1N8kOXJtVwQNKbLqtZQpV
zDs7PZ1q91V/NY4Y4J4O8yz8f8GFaRdtTfP/v5GA0vyBBq/PPSiaAFP/irqf053DLsX9G1436tsR
F2iP8/qYjpLCgtyPViED0ixiYhC35GZ2nP7jvKYjpoXSaS2aZqiHN903UjikSswDtQ/JVwPRuT0K
us+0jPaWrEsu8L0XjlKPHCCguh91sqd4EszZHtpYIG0r9kQfdlSf3otD3BJeLVPDngiLz28d+8ko
RzE0+yhqJ01eVfQafn/a3WwsaWCi9qAaUr3tv2pzyIijO1Y9y9XO7VIfqVGiNOa3BlqjhfO4FWoj
c15zgBxEGdyX8pRfCIvy5R1t9AKSEYIoXnQi8xD1VSAC5R2W2csBCz4iwWOslMaDtkjcbu5BNRzC
kU1QX2jjW6xGLRROVHOUp6vMcxOwwoCY/MsTq24fsmW08GyuxgnfSIwWn2xFMLF/LbS26mlJ5xqe
8uB7qqoNRSTfE5YWoNBogdaEUJmyzbJrOKr6Vztzy9lPfnTYLwKtcW/X6Fj92uXCuiJK5QPtrizT
uhRnVRQod/qm2CQ547yM397Cfk8+ZOnJig3d+3s9InQ5d6nBVGQrCtixzgODzN4g8FfSPOkNZ0ZE
z9dfXKCfFHICTtzFmm4dlO/2YN4fx06ZiRLmAH9C+oLzbq1IrTPf17usEkjA/YVx6efcSe9hrWfG
LMeM3gQzjQ9gudVR16PI4BBu2ymgnzaLwUH49ZYSH0bAHC1cM1N5YULh08tJHMJzli5VGIr4dvru
mNnjmcR0dWoBvi8NNhjR2Ad7/N1a3hQ8329EMHsVud1h/DURMXU8U3EykBbobAp2TYSaDoLOHMRJ
9rzjyG7VGLnhAdVA4FeG8g8xS6QcWGgcIcx7NWK7Itr3cXl7XpKRPuMLbWTD8DRzoOQieG984f2Y
c5S+cWZGoHYU+ZC+ah6eEnfu/Cr6MScaGqBQRAGScpMK7QF54QSplHdsvXcBvxA8ZlAaiVSxBSur
PaWNvkDVIx9pq4wPQxfhIAjS4tTfidbnqbddjUR9qSxVB45JykF4zHJGlZqA1J6FcwHkYZih/Uex
uEfosf/WIbTUGJUV7is9/biTVInEuIbx1ZlQupNf5LstmFQK+7PzJpJ6mqKSZRvpWnO8KcfhRUN8
o74lC2pN6kaKteD1+si17FEdvP49Db6chzTEpA63Sc8nAYaZX9oau0zeb05pmUclfnk5pf9kR8dT
5r33nrntOYQxfuKsfbe/5dtmWUY7aW02Tk3mhlU0l0IT5sWJhIR2c+hbN3YAglcCqv1lAR23tOBi
ybCgxKmNTdO6TGpAVIzgZhaUY9eTooTGKMNe5zJWBRIFWmLdzLNr47KglT4v1oEFL8TbzJR9uk3P
oLqheUXgfZwtDcrbx0qnni64u/b845GOF9LEhjjb4GFAP/96xLtamH9odFAS5oKFrD0MhFjqTqIZ
qo4EJQ8OKGjFcydKxqgd1gutCLTleNBZ0NIbG78s0Ju3DeLlLlIHlVEFS/1gNZHNWAN7Gj6UcK9s
B4ADN7nKQZPAPoEWKMmtTlpf6dzSGGbtun3Zk5MlFXNqaMz4qPs6TfxAWX1tDRqqDXlpaZLk4rjt
JvMF+31YYffZMrWkZydmRH/801DrgOYJKM5w7Utrh4AdCdIGdI42JOegIwOySWoonbsRI3IeGv01
q1NaUgzfokkv0rFvu4uRyYeUr0XiVxeLzN4MOX0uPt7/e8bkhopmI8y+vPi1kkEZHS0HuM2aAloh
4VmVkQESJzIOihlAihONei7LEOSVrD2lzRKKqsQ0psKA+7yuQIQYAP8CVYx5iPVz8AOl+nR2Dixf
4ik4W0aE3Zqyeeo3gk4t/KVyPJ2n04rdSJzKY1WiJMnKSO18sN4mr4lRjQA0aj6Mbjpg08OxiQC3
JulJcSbsLlROo9S0glQ2Gh+hKHI3pLlfpHspaPczSFbe8SlKXfkn0XRmZ3EcBKQjF+UWw4MhyhS2
LKyEiJaXv+hozzaqfIdvm2is8iQLGnizn//xXMDO1NmsNqwHS78uT4Zwb+ICWi411I0cnjetgjaL
pHhievjZrFvHWKs8XwMmB5ucvSKlgCTjEiCWgqZHWbb/XiUWTtOhbR+XazzZwEBokwQDDwiRfMOg
ZFwYT/NCvqehujGJXCCtIcDrZ0e3s4in8gN0qKZfsAjEi5wj3X8GlHD3V02HgL35U7DV7reQeDgd
eBZhl9C8h7WWDRi6i9sCI6yjs3iMPfRyUgeoxrE8UBdUut3o3qjzAgBztx6JtHIDxjioHwwJqC02
aInb7iFNewlog/lAaZn2CF3gMAEkKT9kZctsZhANAwYUDZUbPKTExykjmjueR+FHDRmxvbb0iNYq
j1jl6svu0rIQmj7Lv12cQWZTbVySb7volH/5Fk5JWgSzwWO79a4cJ/EVm9tkaVBS+75VWJ2qJ4AW
/9xMMuUCPJPCRsA4lCByXSJajmzja9R63Nq9CtQ1WKkNv8Ga0PIcmWcPXpTMLu4sJ1GpijEEQCcu
cBX161v4n1AvRtE7ZYeZawFpgP0XNRZNQSJkiYZkZQ4gEqPmcdt17qcfdDKxyOnFVwaY6246gscs
5M1zuW6zMQ6omlXmv/JmzJv8re+qiZBh5rbDE/vneFAvqVUIMLQXGNTI+Bd5wXdHAkzCLsYEG3Y4
S/Mz0mnVSpaKg7EakxwgI9tBU7DaYj7luxIqTZzpQCdv1CiYXF7WiFhuvkqx1INCZSSRUqz2jEL/
n95gRucK5jCRtPzy+ouSQtA4lTwe8BdPXSdFGOvFPIkCsy1kSrH5G2X5j4t7ER1iJW74oOBtvSJO
0TyCBnklTtm2SzsUI6rm7kZciP03MqfA/8s6G9/MIkmvu7P6CvkovYN5sWXXkIu9sPF9Y/q2ppvI
6RUZmV0B8WRWa0SWyTn7w+X4yJckDZAdfosOf4IzblhoGbXUIlRx7iuZWt0fz8WfoqO0/ETlUJBj
OxGdDP/9QiPwlPJe0jMKUMmTi7glMkJ8ngnY/Kt8FjGqOpXo1G2iRT2uaBntj7AMgfOnRTl9YL1e
OYOCfJ7rzevnpv1VPWp19rXryS7XSWMVWT/g943xJwdJ7jcQQ0mkT6NmxWjY1goRNPMyZ2F01sVw
Ln0VJMOnYdm7eQ+79BVIVjI1n2zJ08sMCkLAGj00WSK8ivRPJiv3R9RQ7yqND5rHws80VbNlzh9q
CjGAN31g43GYBjtLZzjCaudn74lMW2WghOHYZS+ERkqPuEBs4qXk8wd/nqWhuNcRReH2tfzy4ScN
6PRfMoCcLNt0D8tZQByDAY9H04Q/EjhNlbzIENOLJ1OUmdWjvYzI2dpA8242oFWY3s1wbDforrnj
8Q10/KQkNMDy9OCZuaeHFZ97tkJzM9wz9bBff+QiKBEmgcb/ncQh41Dky8uEV+FHmZk+gj2/1qBh
lV8r50WL5RpkllB7ru6+EhL3upma0NPGe4qFDNmB5PmIJhwtaB+cl3VH3YpMn/rP0dBfh49GVqix
t8kDVAOpZN56dNynkdVt88C9oC+GOb/3aCwCfVjPOHy2mWH+ire0AiUr759S5BZLTvqIscSVR/tE
qTq3YZZNjKcUMmRSDHJvZHhnC4EdGJZnWBQyNfaNa5wm/PBZVKTq1RNxj+X4EfO3/ISEhhdKHsgI
GachlyLuUukj1SDS5WDRw5dvRcsq2KwBx0/O42ceElmk9oASJ+6Fvm1bNfPK4ulTpXIZItuTbrDn
Lw5mY5/uPonFK/WdBZYrjkhB1qYNw/WfpcfwgVZMKHgPQ//5cuqBCwF+OkVu0vZByQwh1SvL0Mfx
aKl94leN8Nm/oIkV4qeUSY+RH86Wp5MI73CzdKETHnEO8CyTwkQQApuDROjI/9Xln/nHFZuEARkF
ZTfP+Uc7pDMAu1zCpc5S+++yq4HXOs2OIAKeUFrNDu8ZpGgNYH3QITvZry8QXilHmgbYcBAVGrUR
By2vq01XnI6sOfD+k6gLOmfYAeWCnnE5HH4vdDqWXJHyDZATRt3Aw6KW1ZkIPHGOpg/KT0tnPbdQ
gmQUPNzLC9+1BDYVnhHsmJ1B+ypFVZUrbzdOLk3p4yn08JwR33O8UbKYqCJmySiHoLzW72bA62PW
s6pTFQj/zjjfzTWN1phRQsoOsZmn0e4zC1AL+AnYGoU2mu59FsTEl3r/KxMuzQF6yycsNYs/YyOA
sv+Novf1ovVGRrr/SvTfBPsznFd8JbNivJmU+rm1WiTr/m4kNQUzn9B54Qi9tN8COWSfL5UyMfN8
E/Fti3IhIW48HoswupX+VZPuDYrWaZHHb6f/P3INCQH4lN057degODxBfApZsbJJot0yrOgJ6TTf
7BVq8eSsfRYyWAzpht8PovgcnhCn7pdI5yCrXu5KQ4dhvYY0r9sBQctg1E26hFdIX4+/yJ3qYvNE
4xVr9t96GzH/AvkrcI86/5ual6+LY8voyTbQ5G/p065Oh71zGosEuqcT6JroUmoBCrki9JD5pKnc
cGg5wEUKywWJih9PdrCuJFflgI2xf+oIu4r9wsYRCqXxQxCnaW8QMHONhmBQtvRlB+750XJT1frb
ZpFevOWMdZrMwqMfl1Px977wQynM/7EwoqRL48GReOzvEJV5Iz7DTnGZltWb6IW3CdF0TntGd7OW
yudpVFqH4knB2R9pljGb9glkDpRMMqD6hcPFv9n9qqRAu1OjY9VD2DplvC7A2PFZoqPR+44dxk4D
JtE5GTMtVNGPJ/q0y6QRnodQZHdbDE/JDlfCH4IvRI/yAkFYBR8by2/aq2FKc4zPNtL6jT3RZH5m
YKWEVc20uriRwOxXSEXv76qfFQ60eMXT/t/hSwk64G8xE/yP6r6NPYCUZNot6yLEEkU9PYylEpbI
BNBHq42ILTZdGrmLI+HJ+TrwRs5JW7hmsd/zgraOtGamICr5K6F+iKIc9G3cvjnDs8j3axedy9Us
xvXRXnjGIcDrlN3PPVN/oW0q9TASMQhIZpTx9n0rBsA9M3FpA3oRQYWIHuS4GPxdWLX8x9+Tbr+l
NSgvdtnNkIFJl2EJsSmzmN6o1YcH2Z5JjBcnW8C7dhWEwXoRXT+VoZ+AtTxN5syaslAVNG1g6KDp
o9MXMEOzRc298OQSaQsKTbYXcF6oRlSOyo1X8ma2zcP7CNPYveg/Pzf1X2MO/TiaqmrDKilnruMT
31xnA/uzEtJFlFBEsfWjfkzmCVAO4gAWQOaBgRXLxnMFYMiyNsIJYC5W7nHxLFosAz6AuRl3Arl9
f7u4IEopB3CtAvu3/6bIk9V7G4kzQ71V4doIMZL2ynYi5+uj5G25MEqArJEcHfWM506474p7WbTT
pSyFgYRKfcfIfpNODlUMxrPrlz8Fo6RVn0HHba01lk9UaRx5jd4ShAihyx0Z1ATk83zTIKqVX51C
imIq0HD60YOJlCT5AAnawEdd05EdLKqG7LJ6lHd7AbP5+nbY4fr3lrNeTBuwF3y8uhotRVKUtlON
g/66pUfUmQL4y1ISK+iFWhpX+BU5kHBFQCwaC4mLdW+5o3QQwx9wmHL3SAwPVcR4O7+nXF1tDtW3
UNSv3ovB7f47mRsTNwmJZUA73GjDOEQ0J9h9K5dwFG2qSWrJhRt0Fp//MvUkrO89UkoJZFvixMKu
4SJW8BYl2Mcd2CyPti0/1UfSh2wym3Db+zl3Me5rkqLQ0nQaKeiQqaP0n0TrcAuJTobk4jWKL8No
rDDg6IAi0Q39d7UUaiMQVqaBtFK9qJb9ru1u2Xy/FWGcqhRLRSFDlmgaW+ds6q/JawnpDu/s2STK
XA/UX9pdxZoIR3ax/Nc6IhEsloXYFqwmeKPsdv6fGP0pGLktnycmV7n/K8KUCSFxGRuKtbojmrvp
Sx10FCMDw1eRrvSBdLC45QN/xO1wgbM/Z36jg5ydr5di7g+xp90gMnbGQHQptVgxwpPfRHap9dY+
77LygllSXBD/qheSAnoFFhA8qVL2Iy8Nr+oMPSfnXYAaD3XCzMQW38XoS8h6XtDTiNVvDexCtLvk
8N1+q9tsFzXbbR9RvngH6C7c9MUGuYu1czSkPYwjZQXHvK6qFEnovE5RNcpsVEk97C7M7gnb/eCx
SCwiIiWauYAXyxUaMbWFEdWhmvAOdRxwCPxUV/CcakzfsSSwl553MlCN5MVQC6O0ospCrG/Q6bUg
nrMDtcJelaaqG4GMz31clCPrmh/HpenRwwIL+x3Bmj/4GFD97SqKFi49n/KGyfrBVgYsZTqdeMBR
KZTBVhkjo48sXxD+X1koFtCPyuXBLvKgbNC3HGR4KnswAua8wNtWAd6dG3xkMi32d3hafoOYSoq5
e+iE2iQK+UL0h6tz/GtCspt6QLpsSXieNtvca5NqJuRufylImcibvkBE7VWDpZVgYsaYlC63XQJd
VM5F9xXPlpPNDlytoyrhGXXdkCpEs5FAA7HcUcOS1eP0Bdxj40Bf9hLoqDumQx1OYc1MFmvPTFUz
c+HHpBKCWgboJHmbqqJC8DhLfWjnWz0AAJk2u3BVi4v8rLTQztHGpirs1nAYl/tFCRZBnccvB8hA
vdUW1FymCIN0DChXfhbvlVGx89DacINuvKuUg7rnqPMCjQ7Ua0o5jRV3GK5VDxJEVi8gaw1jffhj
itGgWxgEJT9nzqKXJ3x+DM/8dy1vUTUvlbk5VDjF5biWPCOxTwNkmxilJCdf6y0HuFbIFf0n/ipg
DT5TwcNnxLlwTVuWbFDqPPrpJ2tmi23B48yN1er3tgqKcMeqeajsvS6LlEEy9UrMZiPLijV1dI/0
4u6WFFBVfiORZQM4J3KmPpLeHl2WXz6DcTIf8TCba8iRlFso5Shxc3fawi29ozUgcgaaYiMnWFrm
TGVfPKuGUw2knjtOnh0JET5bzH1uGWMK6FciCadZIV+PnkpW+g0o07/vHJ1WRmcxcg3hlrNUN7RT
e/L7tUItRzG6zoZ2HhbF+OW1x5Vb+0+nxwyoNm7upUnKgptkJwW64fVmnuRnSym/yewXUdormRHp
M9W3+x5k0ZLqvzl5ptiyGEntwoyFSvkz5foOjy36+0GOY/50qNCoz7+ZoL2iM4+ctK22KZppkXKd
UzItJkR5n6ZCle2uJgfgcvISCrcxRZ5cbEl4bSZwZO19st8NIpM5oDgTCYsHGAdzznjgl6yoLW/d
sOg9v8cs3iWw3QrqO2t0NBcp/6w1lAzid3r0jiSlXwBH5rWNrfZjNd+CuV7ub/BbPalUrYz8wX+i
jaHZJHpJ8u9fPCNH240Xa5dzaxFuii3E5HQtzzb+QL1A+jVFNXZg6SN9nWlGP11xg/vSv7LGKPGi
zfSjH7p0acoMHNGbLhLM+adSmnMcjhIIAwDw7WBS2zNloYAuMbmIPARKrOLVcq9IsQIJO+XHGVeY
T322fe5nXhNztmEuk++EXksWQIBgF8NWNqts0oKOJwsqMSGkD3GTJ/yEKH9wHfDUjqMcGJyBsETl
/jb0c0kPpiaMWnZ/+PTM/VHH3kBxZmQO/92pQukbGU4OLLi4vf3FMo+nX5lA3EAx9r2CWrmBrzsn
1MarUX93jpc6Mde1a5HhrMGCymE5MyS5XwxGDhgswZyWPVJuPQBR3ogs6avdnXcNuXnOo02bP7P0
CxH2WPVFCpxliAqlXc9kQ5kTf4n0ckKSdFHezTaJ3CyMckDewdjdRcdwqz+gu4KUuukhH6dzp2aH
fcoWNVDaj/QkMC9Tg4bKjmOK5DGQRu/HNznfj69NnzXk43UMBAO8w78TcPlVk9ZO2VFB3kCIVEN0
FUYz/FrIw619E3gW09zNYcx9SmwrMCJCbeYsscTrTkuZKMXSApME7RS+ytMgfREQhaKcCFILLOmj
6tiVXpiGUZ5Az3rFEfOlrLMf/jIVngWIrhbtCOelytJS5nfzOeZl2cDIa/uM18l/Tbh6kzqdH7s3
ELmoa0IU9S7w4rYbZq/BzgpOOmBFnhr+1Xwk14MNse5HCPtP5oYmPqJd2Widn3Ljf2TxvB5oHb7+
oe+DnjezYvWVrQBQmzKxNLOcFThicKaG9GM0b3bRM4/GJ+46BHxcOhsCWR2nL9TV98DqvW57VCc2
60xuArile/GWdeiq1RxnRgwWO3DbhkObFBWFKtf2tU5rHdxxj9z8DcExqpxz96CFBvAo57P0IHxw
Ygy5Uktq8CHwau5vR1I2ZyGSb3rlSmhd74pv53Q71dZugKs8xNpZX2On7f7uDzJAbSN3ZfWb2jtj
LuriQznPxdtKAznvzR6a+7Q1jrZ6JxMcRcBB2YZvBtqUs23dfZseCIuFByD/EgJ/QhorXezgKLt2
ZyUujnYWpkaS7cz4fgGoppCizFMYP3o/raqsC4vNmhRxyvZ/rMReJkBNNhXgUscSO1fPxNCe8zUo
nENv7hqukq85BXZi5IPYLQueL2Xkc/jNs5azP1jfWYJhAuHW78vEWCC6yztknIUlE4DQeUTs4YMR
+Z8mEoDXJD445nBzkp5tly8RQxBWuKqYN6a/AJvzH+DYKF45juDu/kWutc1HPdY+oAF8AckVpPEo
uC2BV/7qQoEs6GINJgKPTZqe2dGMG9PzjIRDelXHQlKOrecmKmDFTGKafT0m1s9whbD2S47Z+5k8
WuhVKyC3oEnkYPBWPU8UchttPyjEiakB/lQ1EFavyNO1ywRGm+DXdBLkBXLey4As9IoggqoPxxUS
ZOtYPLdLLBrWlLNO7EFXVO5JoayHoaHLjWYuiBBsn3HFjp4OQruXdn775AiezM/2B8Q1nfl16Fm6
4fYotMbEQ1lWLlpH7zVqNuLXr4LlktTeHRQ6MFPD2mqPP0DuMFA3EGuDxOtQoPW57p+gepfjsw5c
NFGq/o8CkxAsYC/a0iL2pc3hVhn4Xg6WyntRt7tFg8MFkU92I1sCSfFkdXJcDcoAU5o7v/AP5L8R
uS5KThmEIM1sLBFaVbEYZT0N9GXjK7oFnq0cXv6/Tv0Gxr+oUfEC90fhoCj/IeB7fwmMnKQUPSeq
ndbXDdFrbBudE/i/uo/n/eMR1W7ESvQFcqLrMgZBRLVh/2Ba+Z/PqAUUrrM+v/PprAvSMV6dozIw
SXxdXLN1k2cYyZc3sA7LunME9NeY8QSRALylQFtdq2s8nISwNJmnXUck3aB11b7VTcNWiWEBT9bB
DTzqX2KjagMWQ/dQZyp7wkH+6cSHGJAdj2GM1vuiQ/21SZJVqa4xQhS1bUhUbpT6N11minXUtMAz
wNtLCdypFaOoPCYKGHG9d/sBoNBlsXfmDqJxqkA1OStP5wV3E2Y9omwRorYvXCnlAEmAM3XGJYex
ZXJKztbG05TejYtZUWaOPcKEZAN3SJ5KOxo3IGqgUwf8HF7/h6QYiGGmyONKAFj7SONr6Vo9MLd/
G9sQzojHnnjIdEdmHEuJW4o0HvPr1PtE9pUdUADwP5HVKDGTqHukLTe4xwHC9T0wdo1KymIjtYkf
1fpXlFWlfW5D0q5pJHP+C7Xn4XIZfMb2uDhK7b7O3bZWj6mNptXUjkQiu3iBZW9EKVcmVOF2Dfgl
/JuaEYMWmj2SF1V3li6iwOAlfDp6w5C1CGQ+QTLxB5aM0u3DuxOxxoAP/tc4YeM1HTPv1UFWZX3Y
ZW3yl2QgflJkSkgp7RWmN/zJfwWnHP18cFUn/d41Av2DhTrSKvI1gxMsKUo490nNCumr5HPXEQ1U
Y6algMkGbXsxcME2cE7V2SAdPawPuMzoFlJXhPZGE4hidyBRnOSJGlhBJgZGiyfSdyPxvX6PyD/V
sECf1hVTtWXVDSuxZN1FQ6dvujgcbIvuiMbJbd+nWmbooYC00syTIcYPAjf4ypIlAa1YDnHuVTAx
Jv4SB+CgcFV1dYSTOPkHQWEpbO8Weesim3HCA2J9PyWJLgQrmoVmbRQrPH83apiVYVEsrb2s2JA8
oA1nTKp/xiPjOeeI7JNFUzkgoqkDLGAYUechYLjLbHpv2PnlwobcA6o7aF4Vw3PBwmD6/qqb0Xzu
HHYpB9z5VB6OCd9A2xwUaqgrhmCOuStROMlpJ1NP2YGiuS+WnpSuzeqEGvoPoMIMaowiDgx/gCW2
NWYFI6syBud1MHxJFQVvuHful9jhYaPZ5A7D5ZnGjsvpMiMlh4Fr4PruSsHDHGFBLig2ezP1sEvt
3MHgxTZIRdjuKh4nVvh0pD5hat+SDjUCHcxvNR4ROSXhtfith+IC2EfpwNLUI2mki0Ge8YqNL+3F
A5ROLO40mXh320pSsgKyajWgpQ8BpqgIJThDZbR1TQZjGF0tzWzVC9Eqz1Bwq3btJYsic6qhrqvi
TdiUcImIJUKZqJc7BlqFW29RyQoKZ8p/I0EQp59mR0qTy/WXa9H9Nu6Oq1tzbTwzD9xpfPGv6ufh
UPIRh4JhaGurKbQXSb8Au4sn/SZhBjAoaMXDI1d6og2NhyAZu68jbEFmBtaOWP6Bk3pu5NVRnTjj
TMMgleibvUdNfDgFj3VSyWJU+0jBf1fV8t3tyIhRx9U1PFqdzVNy8BkjakD2FZrWLCjSObMYk0ST
rCxdG5GFZFYs5Tfa5UNt3OOSG5GvLpSWielyuchCGU2FWaErKkfAsY2v8yLL9Qp3kxl4xgybzaXg
ZYHEhYH5ocEGbR2/vYKELy+YhQcFDVw78uZeK/pla0CwMp+s/sKk4zSqoDQ8wsiHYIrTqLcuWsfO
L017JqZYEJsF93rl6HZmBvsMta4HhEfUu8IDqkM8D46VL6vxCdXf0By/oPaKZzx913+jowvIf3EP
4BlpW0iYuWuVw34Icyy40w2uMQqIWO2ARAX48nT8TAOU2ZgM6AZC1DzUCHPFQPUJ5hPVq2HrxV4A
MAmcf7jNgF7djG8a6nnHEgG6vFaXryr6qhtEuKh1WbvkAUZRA2soBkAt6sS1OUmCudyfemNNVKXf
fj2k/2LVQlHQZpbj9lDUarGssgso9kjBZkn/vQXfmwMa+I6vI/h8SSOfSRWhWXOViNl7zlm0Prgj
Blo+DU04udwQjCgJh9DCFbCRn196bVTYvk+Wx9sr8YATt9sXJD2eAredK16XxwRT7mpobUau+OFz
v3C6atsVY0g8I1xcDwqfcVSWieQ4H8QIuREcXFyTV1pH30oOoqUHUqn4NCT5Ei/eC6Igtw96q8w4
JGjf+ePPnAj3jSsde/IWP2TnUCDJBLerIFmRUll974MRHkKbne+9OkZCLYjCgSO1McsPlsC1Th+r
JXj3hR4P+QzIFm5LsG5DtlWyeZ4Sgff5QoKUPskhxydhbSuPF2fcDpOcmG9VMW61b+0eAjgqv0kV
mk8iBkn9WV9eOZVKFehD3nY9QaTt274/2kw12XkZmHV2SuSgKPdgRYO993UrmdI53G2p+MKyozwY
Z92FioXt+GSU0CInrofxpTQXKkUOZHUjFOl2R2qTZGIjy7v+jyPUPZ9KMhai23z4cUufGpM/yXFI
RX4P1dtqCenyatfJVeqcuQ/TecKmfiQOEY6UHNSuChIMY5rhGuc1XVEPAjw4g7Sb4J1t2bUsWrIa
Dj0Y1bi4zAnWMn3u2lN/khQo1tpNrr8mLsJZWLMkUrbyi8ySNa1t1EqTBTk3w2HWDQ5ilAK+BGsI
/v7LwBL4YfOBIz5FkDFl4mmU/lRqW/0YBUZgFCzvy5KVT6K8yID+zLHWFOoYd8flvhOfRXKKAz8N
48tVL8LzZlZmYotg1I6cdWtyDPZ09UP+8oGJUYRPaNfmYDE97LPQNpmRawHwTGMFo1csPjkGBKli
vMHlHEaO9mcFz0euhPoIq/AUmBgYl93/hbNimKN/DqMPoDS2mKV8/MY7LIoGxV2klPJjT6UIv1wa
kFtyIWVzD3Y2cFWWkbqGihNKL2ymuTOU8P8ZNI8FQNXrwC2ShD+jRWkAfHh+cfyB1uzIxk4OthjH
90sWuP8m67QVxrSbfTRFB2OuIX+j+0DXB2LEFbGIPlI0AKEnm+xvanbBQGzLnsOe9VnC8ooKcB8h
MngpmnhWFqZCGwBS9r6gBTUTT5ii2HF/lMmHRb0zY6ovB8S6tCW455aUBFMzIc6ys0Og0EUwaUuZ
LjTIdenJbZXuF3mgiVTp2+4zVeAFDFjT8LreEvt5dlLbvU/826LmtIpaU7l+W6Ldx8khNIgtdktG
eVddOHRiqnDV4TV+EF4v+X+EPlpl2YyX3UxOtHcnstYryoPvWXodsgAUvVXf8hFqfW/bx9CDT8l4
GZM0d8YxkOcTkPhVxyNrC55WG65GV7ADsexsWs0GdsgcPja91MP3Xr4OjcIus30/kXQDdob0Itj4
oZgllDnpP0M8cmARg/n7yrbWx/M7vv0iyL1RCdkDj+QLw7W9cKT234/aXFnQi0S5hiFQ21GqS5KA
/24zdcQr5Q6AphuEP2Xci5DahciRYEf3OzP3dD9p+X7ietVXnJ66PX50AKqB8tjvrPphebxPpe8f
X9/HbgFncw6oSfxcRS+IRRwtq/rm7cHBkRrsUeELdszhvG9kls0XBh6liYLRl7nDxssdRdDJd17L
QqGo8T/8iHxIaczleI2Oyw2dyhb1Df43qk8b+X5VNUOSUeWBuD13jXsymLGRzBd5QT7zfUImYTqm
dQCvJXf7H6P99eGEtB0XyGLvcsScGEsMZuu9pyOrXllxzbqMrTGbe7hRWC7hzvtW24FawLdu4Vct
KyVSRWPEq/yVFpcLjaveNh9iUP9AtzZZsv4xZmYLuwMsTDWOwkQ7K6x7xpcoYLgfzpgNZJzYTiOc
56+k0Gm5G425kymfPYTfKAIKJIsa7LtwBi3/+cXxsibhJX3yqaYAc6vUTFSDTxYbpV/o+Pt5/gEY
3biIh455z3Q8lfk9vdBkrTrjj8h7SxNShKCF7FQt7xrUfF6t+hQBC9FTgEPtAJIjOI2I4hUcajzJ
Gjb7UugTtMKu/L30q0OlOS1HeXpREQAgb7bKIct6hWJ8268JTygQkW8AjAkDqYoNNtuRMXAYWVs+
nDtOqEHcer0/9ZhjGTo9lcPIojR9U4/M7fLeSNYVVnzov0Lc0UKzh8NnRY9Be6CMEk2/VhMiNdh/
u06UkVRk5VjzU049B61AaIxoNrPoiXT8409VV8hmQMf5733j2Mkp7x++0PYXX+eriHDv1DMutshg
HR8uZ6WYu3PPw8hM/VlynbQjSzF3XeSsxVGFmeHzUZcfJKqPv+8BMj0iQxPHpk7cUaL3kidq0MNL
sLgFFqkOGMd0DrvFbepoGqXZporF/ETeBOMwpeRjPOO3SsMmkPDNVU0qIMocqnmjIjn5pkMzue9Y
ZhMY+t9slT0D266M/LLJX2L6l0sHKOBjlNNUYccGV6p4FFSSVjzXT9iLnLMhQHoveN4zKuXsYjHV
MUqWWGXXEGFIYlXtsdO+DeKoKTmmJmu2Hrp/DlbAXmJ9BSgHrGCIHF5BGj29seCh5pDIf0PAv1XC
kS6sekLxxtkWDNt4fV01JIBIAxi0SMcK3OIUhaXKSU29i1EhlW1C0kRnqGVP2i1hdwbZO86vIpHn
/jYB0IEuQmYzUnfMcKDdNEqmrMCpxGjfVFUzyU8IyJ3s6fp4WZ5hMT8MlP0iaoVvRUHD0F/MDqUW
rNhS2XrzFidjinw9kLMrqpI0UgYmShyXOGEG6bXJiMshbdVPHvuHUb4yUQFWth5BWaIQI6GK2wdO
KwpSydnXqJiuxBgpyxZEfiIvk2h6qtXWLhGxxQBAqu4ZQcu9qNawGRHZuyiTYdsS8FhykthGlDeH
CD+HkF4ms8Cy/LyNUQ/WTPv8TBlzkeFzBigaKW5a/fWZ/FXEUhrqfgL+//LJvagD6xxUmTL3Rwbd
WFuuPRe78TpkHWeWSiE5fBY6AMRa8BcMa/BOsJ3a8O2PBiXqBGFrvoVCWFUrraNkFkeYHzdvDHa0
VF6elYvdboEAZYVKVLQLIcIFW4nsKvW2l6T7M1aB4wsZ2dt3tYd4O6C8J1AjUmhDDnZ0KcX5N9w8
/ZkkcggsPejlgT1lhJ8IEoNetnG9KH1dxeQseh9dHEkf7hoFxyq+8iqn4B7cYimpFSV0O5s/jh1l
xr99pI7wdjIRC6dOXihPzQB9Luoy0uM6ZPBKjjDUw7IzsfUwvGKHxjRh7qxi5Ar+1prDynPopBjC
MX/aqoJaQ46VpKQzryvcAeunhAml+MNrVpQ67dMqse6R6RImmdKPLyQoFSrJeGpX+632Wzlke7Of
Mo9F9cU8VgbxWnkDdlGEiOiRF777xQ1RoCNGo3IP4XJMvaY4WckvB2W6jBUywrm6pFyXmiYiK1JX
FO4qonwlKpUTfpvAyr5aP+pU4adtfsmnGg5KxPnHetUw/qJeLEA0hL2VEX23+rZOAqMAtn2w6uSh
+eNwBMFVFugXk5bVwbe36LDYUtnlE7cdvEwvi+OPjzWnPGPBgk2o2wcskKvFp3JLWeEV6Xwu6KC7
JBY89pDJQH/LDAI8qmm0uK9O64uHuNnEqO0gk90m/D/icgXeMr43Ao7DQ9HXvuIUFBIX8iccw4rx
oo38bnxa0LgSBlhi/3qqZk0oIQxWMHE8XGqPX9y1jy6FlmmqiHJgub3fZG/ixpzvbZ1WiHtS5b7N
mC59b93Ceu61bakVgYktqAQW64cFrAo++VkOlazdk4OK0TZJP1NpnDRNuK5wB6bqYoa/uCxvrmCQ
Mi5tuUeD+yYOJ8KOeyCZxjxzCtK+Ztl0CGPCp6T6GfXodOBD4+ivRCKb3Id4YpT/vnIzfshwnTpk
uUY6cu4wFNugLuNhJBkZih4F8AJf6oiwMnUai18HHcQzUPIueM+7O9ZkRg8Xi/+BDjlWYVaHkBK/
Hru2wqexIIe63TZOYjPbczQdpst6CG14z2vwFMvER9heG10n+aO9JWfE+R/8gRK9kxOxaa4LBttu
rLvma0IwMifQzxeBG4rqTK4jOdcUmLtPd9fWgORQj8J8pRRT3Ee9f+SDMFO1IYGhFB7u37kLOsFd
HhrguHDM762opapimo86WE5YXUo2+VglU910AIICO0U8YnuXfWvCwwhnFQxtYipSRoFGQIHA4Bgz
nyToIczRjrKP8lgFa5/g3qdhAJXCbLE046inB4Q8BUV/6brSvq/dMYp9ahPTkWJlHGsydq5okQ5U
9lh8zIp7BBE4kK7cTLpzrRGZk49cuiV4+wRJPimgIDqr9H6xIleRpsEksLUFjb4pM7VW9r+Wsy49
Am3AI2aOJNBzh41kCR3+d32fjbRlamVC+I/uMzzogaC4ui6oYjkq2CD4+KOG0tPqlfGLhZ9VbaTw
Ke5sT4O52htHWmz+5Xf2BFsgq6Jk73DchR8WHarm27DzoK+anzgVvbSQfnfHbEPolWUUhRWJCnly
qfNEN+EiBJdmhoy8hbntWBC+a8gNmAKhEqAnyhcMUlhPKealR9//0WTvnasRm2kjLGjXjO97divd
XDEDWE3D4zAi2SjC5Nv+37tZQfHX5lrDipib53rOp3rX2Yd+PYQOj4pqTSnyRhj4yc3KBs+3Thl0
922NlzZDvZ26s9fI6f2JPP+8MkWNiI5xIac9rYsZG9ogCpjJ3uJU67z1+pQa60Tv2thEwiB42xaj
qJMTTbLvEWcF8UlMx0MovMwBjRg7ZxZ/qvziLGj+HI5lKdMrXWQlkxK12OMrnhGHyj8R0UJBqoHW
uS/RXauhL8K0WOs/UIhfjpMSdEXQ+nkEsLNboDfiB8atB922Dtd/BJUtk2aLObHonEnRaymt3lLf
8Hi73/hJWJQBvE+tCvYt2OpL9ZPvh2eVXFVBwrTag+ZOeQ1U6vh0q09yH62pGFJiw0llyxsGQ7O9
JOtafHS+k9dxR2H/H+uTfEEsRbymQKUfiTzLNtO6HBmvOgF5LaGH+4dZafUq7O4iyL6ejPW56qm3
9/N90SGt4gZsVUfjCbvhoaFMktukkI8l2WVNoXFMXY5wjU/5YLpgblfrPotbF6zTfFuP3W7KHTt1
/jVMB4MZ+hbrvfVL2ZBN/nMM9uvinrG9W5Stlj91DOH/ujjfLnPs1D1pqJSgLndjRO6LqRC5Ui9v
Jrh4cIllwUgYC1uuCMTMdFMPittdEQSCSIihCrDv4TWH8EV5KYn70JCxuDTjUb994Pkd6fbsZ6kg
GTYmaTR35/f17wfxeAEjQ58tv5vwYk43yS8cvdVvJ8wVWgcDPg2lRE2XVtiLNkTfUPSSU3y30LZs
wLRw2431LkZDePuznSu385xQ3xIvp55f2dPpWCXGYAQQy/X0CQS2QZFhds0bGmKbNu+0g+EJM9kL
MvebGBWUpBFaHdShXg9HJKKWeB9CnXzczYBKPZW6KkYhReunuvC+YSZGkuxtaZyZfiQlYFVi11tB
Qq3LYwM0nzboSi6SriyGUibVBPzq6+tVnK2ni8IcY19NjbMIKFjruur92oOK9DT/D9jabgHzXwhU
Kv+bpPNOyuNVd+Ch2FbrBjt1Iw3L4QprVa0pGVc0lOQOfH1A6EKQ9QZ8TgEqOqq/SQwQGdwCSkGF
1HWqBO2yOOYuvV8Mx2u/910oD/AgmvHkr11T96C7upy0M1l2QT6WrG+iY6OnS7VL9MCvJyYOE/xI
VncGtYpDZR69l9NlEsf7ayYmokPA9TcHvrzqwFH4Gjh4ojhqbbawrybkjirIROPuIRhGN2Jx74au
GkXFt0XiGa3ju0KY0ishBuoy+7DGffzsqbQSV//2F/qUg+sYZ0gfOlNV8V5KLMfn9f+zZkBMXsrV
8t757Dcqt6/gjGUIdjPcmSBGr+ZYk+d1h/tdttAx5iiaGUUg+S37To1//am3oZG2RJsp/mttEP63
iO0iVpSxJ4H8h0dvtyCPtZjC1JHlavKeZLEJIb4BCFqLuu8oCtNNUNnkKZwbpbV56llxaF2UT7Mo
/FFpyOSm98xiQ502KHOp+n/YaDBDd01myDLtzH8uifwLT3h7gjsJAe2ZQaM4+bIb30O30jED5Efo
0k5jQEcUUDlwOa8bYDACuzlp71EtKJbl70ifAmSgtScZG2rcZmgoVn5AiG5Y1XON/pwDG0TOfEqQ
PZOuufXmzIIf1Uh7WDwzoJS9Rjolk2JI9Le1cqNEyQE5FyUIN94h6qPeHW2OdyFMtyGNiGwqiBFp
pvC6OGzO0NqkKJjBz/u/rvOQPLaZBC61254OUN/wGfOMGXi81UIB/BAxu+qGwTbfDph2RSslwpa/
U/SBGbwfVbmmeF0jxUltpXbWDa+hQ0UpemQvz42tAK8DCJc+zzV6SzeY/xXmxy3IGH3AA0Fssz3w
pknClOATHn8xKqgRWFLVm+A9xqOV7kw5zuOP5FwXx2uFZ1Y+fc5xPGuU0uFHfoKXIwP/w5S7xPQm
rtP2EjUYzxQyx2EUXnmgiRC3drH6f+H2RVjXlAXto/ilIUH0AhZQzFBx/gnFeHZqlBNkC9cfnGnh
6tHV4IUSElwDzt8OKPyNRpjbu5qRpzMDGQBv52DiEX3SNBLguCN6X7ukGBIdIO2SRdovV/ang2nl
YRswLaxi3AwMFh5C52wLeBeLGtk8Y3Hs6IUHD1JmMxUtfg58jFZ603k7kGj15ua9VXk1rvz5pzqI
zeXsCjbZ8DBGkEZYp6/ZUshNVEdhosDwYwiBE2SyQ4xcc595LfD1t8XFccOWWpb4GbDDrYm9TiI5
ymB1+tx0/Brbse78+3gAoAxPdPM8nhbHDNbAENwWQXRLk4gkj/IZ3XL76bDjTWiEleX+BePM/30o
5tHRQDH5s0qSuk5mAs0VNedp3mUeorh1FAkgGRhZsYJvtRVmPnjhS87KAOqDvqRTW/SxMtqxz1lg
5w6fV6LOM8tHFHzvQdt2OL1xJuoWnAfzCOUn2ckSwPBL5yBP4cJoiz/ENSa2f6DMYSRIVhUHpCXv
AUmL5DI8xxeGgkoBo/NN5VdMgUxuOwmvXh5CpzpxxD5XmN2C5Nit1AewZ8Q6RYmTA9Pe1mkb3/XF
Xf9QW7ff6lWqFRdb80fKf0sOqHLLpE8clXkd5e6+TuMu230RkB6IHQAQ7mwvaLIIUPWa+3MVHkhM
4BNqzm3r0vBFcZ15Wy1CYua442ukWmPxFqII+afxDNUwKMwx1NFC/NbagddLQEypX+sVMxODzLka
uMz5SpjnRvXi1y27CbrKGETvixdGxyPMjaX+ZXHliG+5aUTRIKFATG31oJk/8/55b1oamy7fgfvQ
Hkb/LDPnibOKU4wuuWcXuit1rvP5Ltj+QbE2cU/zdsiSh29dc3eLFxEfd+gvBZBpPxm/1LZi3J9D
Kzx+nCR1Lsyzpe1rDRiXe0jRuRvzFMuchY7cc4vmsCDYIQwEf54on2e92N0Q7KGra7x0YmGOA8Ld
UzG8pact/UkcqfV4BUQx3ZvD+UqXlchA7NlX31jMh6mgCBLBSJffmOuCWs2wz9ubvDUiiy6oc8w6
oz9GqM9mUgMTjiWBWHw+X2F+ii7WPwN0M1eqq/LiRrc6WzvVj9rcFjneNoJULmu9ZLXIDTIRTylb
Y6lAAUE+dAu1s7ThxdaCyfzy7RckehM9sMQweAAVZxiVatWNmJTzN4TszsBNSQJ6F5A0cokGUXr6
G8JKIQI0PXMf5ulSsYXKCLJxpg6C9wjjphjjRCvTR8XURpQyw8RCjOJsGte1f4f+CkYtLRwSHUaw
QNOvJPJjSVtbc6cRSlGqyiIxPdPfd5dHUm1y8wb/SSkciPfvFN7fdh9ITGksECBtpV/vX6OY9UXk
knM2Sx6d4qv3WFjBa2/TKKc6SjJHqmzbhC9sKxPda3GEeNb21oKsnPI/owarMLALpvHxUE6AYQDf
hUX+tCDBg8IaZfNDVFCQ9c0aEpXAVSBiQfWfAO1ZRNfzjtjd+VYmQmvcGUZaS+OUV6s2xJVaLXBz
6Mug9bYr7w64tUPOr7y9Y8RibS+omx+xosT+JsIAZe1hpzs8B7r7/fB6AAtMxL4iixxJNs5W1qRG
3kot+y0mG7W4eyF884lUaUFJ+JGuL+u6qBgTD2QiU0Rc1Ax+KHhqQ2zy8/QmscWKo1vMKUAnEhIq
zMFyv7S8BbXKiwCrR8UFYc9EFW7z9YXPk1M/8EMqfDswiJEQxSnNnmaw8lh9cjYAyW+GK4nrkxrb
8xCIw7dIzyCqaw/ozp2icVQeeRUnZgvrx5gl/euNEq2CwOhzoU0u7+EgQBLTUq856w08MCCKxi8t
vZn/FIjWxh6TSAaZTIkKIfSlGSmxtv89GouU7o/XVdS+dpfIF0B9Q5PoehsRyI1+KPP0lQrN0U65
ABK3aVFCZDW2Bbcn0NfoU6txPkDkM3O0/SKTYDB4H7HLMFmK2DhZVur2ET8B9ODlyPgKSwBm4+Wt
EF/J6ML7T8v9f/iV4QvqYNw1raFBjuLSWAfv8p2XTg/7tErE0lQb19aace1DOB+bUo0K64KcT6tf
YKAjAAZfGYhT9E0EtAKmUMwPLNi/i2QYj98GT94fy3GpfycSYeTG/0QV79iM8+wx3X6BrFqOAY4h
lbdj7DijoOrSmU84JdWpDPB1GAhIFJe9R6ZIVAKCoxWm4ezG+eqeXrJR9d11akKc+v3LwRYSPYKX
oxz7nJLNniJqyDxqlyGmGh2SeQTfjLZ3L+ld4pKl8XW+3mINPPN9yIvUYAQqEL66So4RAN+ZQsgv
YV83uipnpqeATpWlGFXVGHA/1DZpjUCed+EGWwLHilKQuOD3V+YdOlIHnZUWncK70pax8T2THZXb
HdFgWA1imbC5FjqtPkzjMip2ofz311PTWjkrKltc7TKM30TOX7yApiNcZu8KilkAjSiqBOea17hy
KK39URShHPkJuvEVH/21BzVRxIDOZ14BhGI1WMBWBQpqj9UClXA56IpI0aIwhYEzRa9gUczZfqq8
C5Hk5SR3KyGXRqlraksSxNfM9J7CI/9YPWor+FpfwkDBtGCeiOYUIDS+IFxTeZN3SYu6SCQ2socQ
O0tAN/pwQ4geaXDwGx7GvbJMrIKwiGQX/pFaisCYnGhC0a6Fpyf9z5rxq7z0Uw0WI40Do9r8fQvp
boruvMfIK/ffu4J+6zApBNAJpP3JW5NSLAyYdkscjjIAsJQxeL9EaA0e/5wCFtyNh+x6QYHIhnV2
pE0VYxbP3OV3F34cGQ0juH655RBfc4n26kC6XjqXt4RwjAH5H5bJAnaffhYjNqOWeuCTg2mmiqfR
B6aH5hbFC1jJFFGlxeG8Msu4c1Hq/6ZI+RnPGHdcZc3xMLjogxwZ0peuFiz3DFLp3pHoZvR7+h5s
4t7NNEQtEBnjwSEBrisjRzMySixRgdGF0W1Cck0GTaj2QdIpHPgV3XtbJVIDkqIWYWSa/xwb48Uk
1lwDwdiLTy8i2m5dUG/drxc9H1PLZoDgyMlIyIvZb0XoqKPqk9rPEaX2dXsC3OUEYPL5WOgzuqFy
TiumrNnQLfn6P3+Rg1fNUSMcdPU6u14tYilUQ4ENnZrI8Ga/Y8TEj/+4eujiD2gSKctkD9R53SxG
a0Xw3uzYuCnHtRVUnGu4uecetrRhkJfLLqGDy9cNUVDqM4ffyV51ATajX5qlSgWTCCvDJvCCelAx
96GE7J+tYSq4afb1nT2yTQZgGph4nnbo0DBwRKbUV4jzVbAiSBPgH00Ea4jQuueGU2uyqMjafT7r
546+xPcSCeztv0TwNiSbvU8xr/Yyovs1i+YjhZmVWm25SSZoddOmYCpuobcyFEDEPaXadMv7AE/f
AjCZpiR6seEA1LhqJKvAROV0rOlOURFUhEJyEGYAo/JmGVOuFesmjMHvsJT7h3hgabyDMF3jfZff
ZAhBTsphhePko/C+CKsuyOScvb1/iIY+hdIYsw78nga/xn0K4tjhX9YG31QhV1Uo4Bvwv/75Ebmf
icGqKXdLhp+GliR1ZqRnJD4AsFVJoAoVWNLVEaahBtb83NJTyqAs3v0ndDuMWTF4jnUq1WkD9W7O
raLn195bcshyh19UNw5qo7fcgwDct+mYp36TBO4T5dHks7C7ZYLdhh+ytvoHZ7h5E0U8eov1qBTs
SZvnbK4++F8NqRx1wUJ/z68GANwHq7LLeGjrxstDkdlEqz85k1i7jlWBlxi349MHv5482Ygt6DXK
j4vRyrlPwlPXEGSf4zC1Cc24Jvp6YMT35trVnBmZNITklDAhT2cMRfM0bRcQSyfuXuGWIM7vKUL+
gbdZvg8Uvxm/iqJ4abBl5N1IG7S1FKXgBtTCM5NCy5QKJGzwbSrR2Dc188g1NawQj8fIyk+vT4MX
o1N13Ru1dtuckKvH2P/p4HwbK5KRDiv4L/X5vtfiCU343oFRBdf1taz8GvUXRgJiEJp7ER24zM4r
rBuO6p/fCr3SiG+IAdbjO0j6UryHKoocBFaO1CBBQSRMEi8dhsmJ8R7yGWHpqc0oj4TBTQ0Ge75v
NBOZXZFBSRQtcXe5RrbUucnfO5DzsPHFrTrIhttdbY3oeupxRvQdive/g30N6shF0IEDxof49tAE
ciN6wrfEZ5LYEbmXjssFccBJrjYzDMPUFOqpOIzCIpzQDxDdfhIWztoLKr88Bwi4Sa4Zk4hU5XRh
SWRirMH3/BVZEjg/o/mjQ3eeS8ixe/pteclxugNWNfY+s7uV56HVXdOpWyhlHTpOmuWX01QtFMul
EcJvib+ozJwUD0YhLGH8e5S1NZBZFNz6eDpdG+dEGZaJrHaw7iqbbc/BqiauCeTkS+8P86N7HjmI
5FN5CI/YBeLqSSdk9uqlIb569k+Mc64JJ78udvyXTI4/egM9rc5oGJnr7o2/kPz1nHuYfe44+L/W
OQjAE3RMTkbQ9hdaiBVvuV1brDSp3nroQkcSWTxeFkg0an99BFeQynu7nQwpZrxW5EFvQLVWIeR4
M0LFzu3KZXCrDOROwEKyOR7m4aZwD1du9xqF0s4Dvs/3kFoL5S+AxxaqTFlww16pQEKQ52RKlHEJ
JnrJNv+3aQRVCd0Xs4KM1lIm3TW2sSoZUpHHWqwtjcq9AeI2LAUyBxIBX9EjXxSV6XrMh2Ow/7ek
DHTH16HYnVcEM9OxCS4niq76H1V8WP3B1JYc0kVGzq0v1cUmplz4r3isb3phnbSrzbhbwQQ53GvO
Kf+hR75HUM0Qxe7h3WJb57CAb6n41OjMU7q7zFd1p05k4CkzWo/JqyGMhSzP9/E0Nnybv6CpNv0I
/R9Rk+0UUm2gCnNqwGLz0E/Z62TihO9u3fXRKaKlaIUPbrFbr0ccy5R7HhrHLqogOjosUUT0kUh6
/jHOV6eDCOo94oiOKHO13UjoUHSi5S6robISvuZgbUL3WTHlcZoIfBIwktEohXuR0k6gvYxW9LYp
T3S8/NOLQVVudzNOHVGBdebNMd2vHAfgs7Qqo2p7LiN9Z4j6QhyO5smyFO9MiRO4oNZ+hQw15S55
Xmwb0c2Av59BX1dTWUJqQzXda7zN/XozYso508K8DQGsWg5nIOFmsd+aDNUkzsp0hv8idj0rS5oT
3hFUjzyG2yFqKjzHMa3yPN4NxSdyUCbPurvyitpbBqOHQAK4Zy58c7Hrpaex0Ij+oF0HknUJz2iZ
bj/7O3BCyHqs+0NiK6RlTRbmUen5egz6i0EIwhNW2HNRbCpUjH+91ik66H3+ZYZIw/F1LfhVsCYP
Gl7W6oXwY/BHrv6gJWkISwjJeIHCSbsK4eeWDcc5rpAX8LSSU05cM9zm6y0tEoktuGUnawkXc4AI
tFfHn+GKQqglgm83L2GbLgR4/3oZ6S5TyjJmXLQBnH0QX0pi5JB4WB78z6YAWt0UZya9uoRyhECO
itJcCC9plWWYtzJsiR8qp9F9QxoRRnzhH5csew3C4Pl2UkXCHMzXOfG+zAG6H56cbG9dcG5dvjyZ
353qmI/Ajx71RADSsb9yGZQmSnP6TBKJiQrOpPLXuKUsIeAnoH0bMQ2FfOHR5r96uovWdzcWT3A4
nkpOY9PNxsUu5YW9d+JNNxIeaQWGyq4SAs4mR4cO4uyJbbZfuHl5EqbL708rReJSrMEGSJmE/BY4
EEa0KWMa8W/XQ7ygjKuedPPgC0onyhndq209CkucllQd7GocW4R0UzlOGphM1hfAKPbTcZ2tbepy
Ha+r9EC8Gpc+65Um5+ORnr5NZVH8VBXj9d78YGp2/hBw0BTQ7b5E9NJZ7Ps0cOAw7KnOUKtJSpwR
uVcvcNRjMaAlerjn5VrPbqSn6gdHZqxmquuJfiOGVfYeauooej3/Wh3L2gcpvq+XMU41MXLAHVEc
aOu0cCZ5LiffaIaz1ztdRX/2JpiRsOAaEXDsxSTEQJAAk7iF5uCfyvIC8ndPO0ykZeXHzNnO6kCH
beNxyND8ADPkTWkpxJqBg23plHMOkpERoy7lpHFCiTVDf+TSUTkqsHYGs8GAaX9V0XLC7cY/fIrh
TilwyZLxmbu8sdapYHWbHMUb893byRjD0R9BrvnQfJ2rnNTVJMj7RIZ9ZiKgmDRhWf132SxFvhp1
6pigUpp4BsAqksmH/4XRLpshLw5+2oGf2IsRIJCQeceoLhsKWGrUyOXdmBM7ciLBQmQiwTR8VZKb
NHSnTFy4QzTOsAj87DIOp1asSVcB2VWpQlc4oMndr17J2YNVQZCQ4X6UXia5g+RmQoZAiilZFx4P
IJ8sEAyIqXxPVBkdrLbhctfrsdcPZOGK74eU3cthrCN12scHKepBBskZkq5PH+sH4IlAPZUImQh8
D6MFeRabjiKM1ID5Y1fMecgYwPZkW0kD0h5yEhKsnU10iKD0qsL/XaSuClINihEwV62CpQDYyNWT
oSgU+rUHmorBX/ZAicS+eLTFn3KrnnJxnt3b+XfYVndz1NUl0v/nnd8a4d2P9ZcDThXdzJ5Ga3oA
WVJTE3NfALDzDvYBX3fJddckhHoVACEHboOug9k/ohJmLGL9FSLGgJaluQ+W6vijTv2PpYOpVrSN
0t91mX1KtTQFI9orsxwki98df1gj5fmefZAoKP/6ED2Y1NGp/lEkXUCewjOauvOd0EeB1n1FPOpC
hXr0pFlUqRyNZtwXXOxuR76QJVsHL4Tk7525r1jXH1B6CgX73kZXiD2VQH81sS0xguu11UX7kwzG
oy9goDnhmh9x7cduYEtNcg3l5jd9ZeQVr+ktpOpD7x8/rrbi5KiCU/l9s3Vh+xlWzmCQQkvqMRZJ
4pOw1ULtswXif6vFURKHclyWIfL04ay+A7coi/Z9TJyW1b+t5kIxzTWJ0SSfyJGk6SQHF8g620qC
0UP4+IlB3cvho3wrEQ0v1TUrVuRNy1Nebz0jrcWAuxZraCziJu+xybbNI+5827XJhxlC/73aj3b7
eR2xEQxvGH7SGE9+lfImNYsFs4KepNex1APfMiKad6W3T4T8QkzJ+C9PyZtJCilYUJWz+j7FJsYZ
Efd6BOLDTO6NXa5ltY4zTohRkrUBLqtsdoXLrBvw39wqAgbsBdH5yplX6sM3f9I3eMJEPinq2GlL
uOHtGAOJ63IZFWbEO+AdKQSVfVAvhwKQSFlSmZSHUW6ql0Y4YVw0brE+BaB2tllxvAdG39y15igO
s+OivHfEFbjiGcjZ8j0BQ24ta17wkyyd6a8epDU1Tqn5PD+qCyX0y1IrOEQG6lbIkixK34lDVx0R
VgR6w6FjgdV3NLtJs8x5bf22peymI0uog/8RvmXQdGJQC7BujqKrFwtmfQ1bcpFi06jcG1tBZX/g
4Ud7kGJC2ZpoD1pln3A3z+wSmzrCrfpRdbYTQ5xgB4iNd9l21s3tM0OVLFm+5ffyqilvjWqRAiD0
Wz+y7VO3k4LSQ8TPTeGweKjCuxHj7bQEMFuIOQWsutx+U00RHVWIrR0p6X2uF6o2+h39UG8762AJ
XQM7WCbH4PbyDTLNjvKKnNuvcsB6RHOaCOH5wXbXUyk8rPxcvngrTSHsB+IsUJu41W27nbVLIrs1
qa2bp0ozYEBSD8v6zttQYJAcV2PZm1mFXL1mhjJzfMsHsfW5O2/H/f69Jb3U1Ve+Du3bvJ1a/7H9
pGuLcRbtLVkrXfaeyBa+WY3MF4DZdfwqXTGYjqHPwVHGAX/hWaX5LaZ7nT7UvzIxiHhMtNnoad+e
tOTjxDZysz6+rMQX+P4qXPzmIgs4wjV6jN/eLuZK+rJQdNrOAG7TUjmwX3DjBD5RGn37TnW7bzUx
wyN2qaYRuQYJYV77KzcZQtM2s4vg2mi/ON2tRadvCv6ztrJ7u7lmFky7l1Tx/o2tfPq3HIbcx7XB
yHbwHIvyE9wpwwNZlRg2g8utYyg+VaWhO6VqkpcRtG7x66QauYxaqvKhFAmOhWkGplmjeRPeGJF+
GCuHYkRRFm9q+pGRhWyNMP3oB6dhZQ7D5wI4a0QjShFKtL5IvO7CZDfmYDHc2q8vyK3TaClSC5jU
lEsjYa3TURa2p7/xt+2LZ74krjHMnFqJgMXrKgRA4pFe0xKeYzRl/wtle2eFEUlWrVfdZ/cup37S
sa4oQY0askHsBYjj0ugjTC3jr6ukSSrLShZKtiOIM+vJsEQgVRiN9coy0s+RjNkaV6bM//bxJP0l
ThyYL/y44mf4dKlMjO6JhrcZrf29oE6yainZhXGQxl+t48DbjmHYR8iaKstmkVQ8GJigRmd6Hhv/
RtzMTg2feX2XJTXoZkoE0usW6CDUVTi6NYhpmwVqO1WAGVLG7KHw4rO7Tjh4TLS8Y/Y5O6PJWXD4
GdBjNfze94e2hq9BlZjCw9BTILQN+O5T3ocuqHjGtf/Wc4FNf9zgFKOJOeQ4n+JlXzv9USyMltPp
4txpGx3WOqLxFDp8wi0WevnlinwOq0g+j5/kf6xa22c5O35Cf3uellZCorVwDoc9i/a0HNUP59Ub
pIoK0EzzK/sFE+DctVD1ec7TheOy15nuKUMzq7kqK+ccGXfLQJyIteroEQew2xzPMfTb4NtN5qM6
RanUV2eFYrTKx39F99szmT9lW0AJJxUGlzks4RJOVYxX1HBrmtji7jPKZfFNKmJt6fwaODEYqNYY
KzM40x4tovEjf9T5jkgKxBNkk4RtsqNCD2SPtPpksZJF71EtSu0DGVqofis1kjm+sX082qqHHKds
wQ5PrLT0Qr0DQPSZ0P5XPfHMKzVAbvaA/FQgcU9r9txozHGRlpYOWlcZFIoPpa0PcvOb6dJqWmff
flKhFTFgXmFPc8qAgMOdS74GtGsHYFt2tY0ITbvbn/NNHEpAZZdbdSzuurDSNtfWHsIiX3L7+a8C
LUU6WCrGOg25pzkrKq78iw94Lb34lSPmJNmzpI49YRR/kIw+ScJLgeI9O0cZkTsRyl/mS0P1IJ30
HMzzB12GAreV8l3ZznrhcZBxw3nqLaY70PSU8noEX1hrfQXGxlt1EMtv3LtP+zp6Jjnc8i7w5yvh
cjQenmPCosbsSSNQMPkZf2QRmDK7LrZplPr0tJRpsKLFBseYa+6rhsLakSdlElTdPFqKjQHIscyp
ozry1DbSO7PVTPALj1xX9by+82pVVZnmGQDyTj5wvga9YOqAD96MzX+RswQI4CZI6TqZ6r8KYN1T
Fpm1PfsBlzn9K72t67OpOdsR+jwRS0F8smyWZEY7TVfKbZ4jYnEvsRLR43xD6DnYOw0sL/gVPGvQ
u8T2EtuL6ju1IWdbSWgze6qWpnGYlDClUB9KrccaURQIhk46UFvBQNJmXfjvnb7nIAp/wJi3rpVu
MT3o0zwZlWpX+nT4iaWLVQWCIgiep5UoG/HH/qatbLD4RjZ8LK6pZofeCUoKyEr1jC96fQZEx5yq
xBPdVEa1kQ6P9A91ewyOK59KdDQxmMiC9AXrNq5Ebw+N58RrG/XiX6xYCg60un2a6g5VwQwuhCHl
Elo+aj/BdEnK5dDR59UYAtAcAA1CF8iemHmoVIeBRLMOa71hiT3Ow4oYHIdqj3c+AtROvyG518CV
+k2Ww1Dh5JceH+fugWK4av9PNnCT0i6jb6qd7xdk+HzpO8mRjrqJcAsqg/nXxKOFcmTfBWpM/h7Y
mlBRzK2Zc8xg9wxwKosUxkNs/n0tfRrrdBnK7WUznMLq6VVdEw3nxBiHdTuyylFbYAytZl/cIfQ1
V9FUbHXmi7jUAXOJfBKXFtDl2CmjUmxs9eblcXeDcpAi4AGqWnTgt1T3vD0N5QOlk4J9kDbD7XBG
3Gh9DJ8sSWHOnTch7Ue+qTW5LA6IbfwMevARbSxNoRbM/SZNeOtze8rnW4WFpHAYaosQSjE+RGLC
6rvtNnKnf4AfQBYNbexKZ3LpP4ajCVhd/XByI3T3mbo7w9xgMj3qGcsVsowexawjhlETheeE4GYc
z6IMzHQWQGLlvNXB4tIXwZ69Wxs84x3ePNb40o92IFz9qGpYzsbNcb2KXAVVqoBCociE69vxpN9t
oIZrOJMt84Kp3F/uMl7LqBZ6EFOjSvSIqp7kPFHCnY5UeRxUK/Yio0SH5KqRz3RgQui3ScXxx1Vn
UoOgvEPtBdBrERFXh4Ob9ISR0LXcSy4ajcrrUNZ+8Zc3RdbPPsR+1fFerzk2wbGaeazyeta8ullX
Dq+5GZrkHqBKSu92sLAMymPO2fpUBSitjs6yux0TwcoZqd/hag7ZdqsQebtPXb903uCk8zwBO7jy
SW6l8nvH3gEpo8oR9scMlcETiBtLQBaonWtE2/ATLH2sCXi4qAO2vHykD+2tSzOvRnOEnGxHbOCq
1Len/iWr062utQUtn3pD//khHd3Hh08/YVJIuLUCqXmVHRk4YdwcMNKPIXraKcVL9vTQF9S2sh7O
2+m/CeHmaZzqWR8zYPQJlzGTiig7v2giNnFGHpuGr9FmH9X4n1YEYHswBBBnoXLAlS2dLTrR7BX0
9tTF0/7gH0DEodxBdI30ycRnqC0KLcuVcLy/r01xMj9iuQcaZ0zlCtMvsxIMBjdL9KfKIwsmAzFu
hK1ETBldnNw823ZibTg8RRsSSQq2fPrUHicijaq5q3qu+9IM7MGGazYzy1waSF0tQNXOoJ12MqND
rxrQl1mOK919TbHOtP94DetrFnZ9MX3mVsGUPxGbI4FDB+8TUkmDD8VMrDOYPClAnbqmPiQlu2Wy
6sLtF3+2uV1Fq38xznMLHxHyUVO/g2esWGN35nHf+nApbL7nD0KWhK32v78xsHwd0YZZI52SMfmd
1AFRSD0Yj50h2WnXNdZOHb8zUSevb/2lzEphxVio4v8wPSsUClS9jvfBQiwAtTtFHyesMdISRUiI
k16VT+hkp4VsT+0zxOPZiuOBVBpxkp2UDuzgzPmTROgCEJRXCHzHhqM1zbG2rO8z+C/Pfwv3cYo8
WtXlBQu5VfRxcBY+3n/JB1DMHoXIpUi9mXyq6+qsuxLBkMxyghQzo/cOcIKq6R/lD98BpmExhZgU
Wr14xg8SDqYUkKexm1r6FCcSRL+QUf+qB+64tzf9GprwfENiNVT5/8oxTBzRf9TnHf1EHYg+W6KB
DjbhS0Z0nb/JHmVlzfU4P3Lp2yHFJ5c77cKkgzmWxNqzFVeoOcMWV37cbLn8X3/WfiIET8Y62cMD
kesV7kyZXAtdpAzhjknqg9t8+3e8bA7qs/dROZRsz+m69G7kSp30WgzSf8c0EPqgB8ugL+EZsRb7
uoz53/fJofUudsXPQzDcbVQKwl+/3RXDWOjrv1XvS2BaOHemLGtv9lkjjXHIRa+gO0VxdMl3FUnf
X0PI7MKruc70KxUY5NJdnMe8Xo2kmwDUwq9SNoBByzfaCHeF31F1VOm/NEmE1pQ7kjHboWUKiSZy
5SHXWqeLz9+Jhod6+T+ETvyIahYf6s3jEZ5mtxK0ELf+pEtt0JzMvoF2VaOYXm3r0/8Bnf7sYLVL
Cd7qNYRSBiZSnNijfyaIFdc6KtHMx8Iyj6juzXClrjw6AY5AKUG1n2CvEGy4NGPz/nlNEAUvLpxv
Q6/OwoDzKQ2En5Cnd872HZ7+xDHCMT3uqB8SfwAODQj5ytQmPO21JGEWMBaE2lno4zumCsCXkBkW
vfKi+1E6hsxXxytzPb4g98czOSHNnv0hnPENOyToNpP+eK2l6LkqkKltvNSbWz6kzk20NHZF24Sx
rQM1xjFUoMt/r63PGNTz//eOIB7tcIsBG2UnHZxoJhxwioKF+wVtqdByOqMtOErHfcVu53cYI20/
SRu9SrzGBJsl8CtoI1kglJK9dn1PAOt1AoKL+UYQSlmRobAw+I2iTkZCobzo7/4QoqfrGHRrSEyT
WX+rGILJko2lTTqukDpaV+cnIgoJQ+k2XJvf9QyhuqL2gcEjkEaKxnEgnU/cK9AGK1WvRPQ4eXsJ
uc8/LkgH4v5Y2VQkPW3kxYqefiPF5r4KEyVw3xlCrQ/mIAAykDqg7peI1VHUetAMeQ3K8eJHNW6D
yOidSYfj4LNTOAop/Fw3IYiWfGXBWPhaGWe4eqe4uwTiTRh8+WokZoEJu1j0fQErIXTn4HfhRQnq
CP1iQBBK5zvAtxoW6J/zzEobwY58vDH+ChpfHVL5j5p1ngUiaK027dVfW7lbiUjIkz+6Nhz0YndG
zaWUOntaO8wjcQKe+XOGe4wX3gxfGiWWDJYXCdCqocylFOv5zxePdN+HXweTguTmxSE68DrwtRRw
fOQgkZfjOmRVb4JoNNrlHCrulEcXbhq1z3oonj6ZcLJZx4eyNL8Mh1S5zlfGptRUR0BeSEQsDh8Y
gkWzJ6H4Knf99/kUThwp58nETTPbWPsvD4f02ruc035vqEhwoTDTUnkK1MDQp2PPvpY/WPy7hub3
Er2WE/wKuDJmTSH/5PhLdwxYfdYPjHxaLiNSo9NAE1mDUjRqe46L428HCTX8jM9RFd4GBsZ5rELD
fybU2QxQqHNZY0N0T0eXBRIQmyybz5aoqupAXg0KropVblOfsvW1UyA99ARv79ZzvLp48MDNUtYH
0zsV2XORQdkdWJceq3KGxkxlciA4eZzcTQ53lt4GmTIeULsVsO8PG0RP8dCLI6UNCC7823gCedLM
ARHUFPLwozrwDNCsWZzSNl3DRD03ZiVE3kcMAUBzYaCuT5DS0SkcjeF+GSU377svgz2Q/w9RBeOR
VL2zciKzUi/+lmjAzWgIVF0csY+YRkGOJScDSZ0g1DXa45izU48q/DMPwNsKtGmzfnfCQi2iQEMW
NcIq748KviguKqSlmMZt+MeVKuNxdNUu8q2/njuZYy2YHWldTlb7d7OvTt4Lcpg8HwLxaaO3+OmH
9yvxkr4eUI5LniMg0dnrpBWZWm2hgKfoshBMd6wC2GqHWL1hf34EyiF8nTFT1C4aWvY8Ip5Ufp+1
Ffx8OfO/HLEIKE+IonxlfcomwnkYH2LcKdt2knxbYlR5Pill5SK9igL+3S9F4uq61bnyFmAr0Wnx
xUqWLEvsTVU0pkWVcLl/6fTQ+zusws3Kah+MoLJaIdFsCNj34kHtll78BgNtaHqw0JJ26GHYqC8R
/gihFuLOLX1s6+XyY1vxrPZYWOQUgv3wkXIayW7mBz4foYXhGhS8Q7+tJPjqIcisX+AqTCAPo4UI
zDmfUctWlVyVTrt2VG0lzgQtI+NB2Cbv9fgDfZ1fjq/e9EaFacgHCUyYuclb1bVNkDR77U3xwnei
MxrGS8tSVoNa8IZ4ix4/ZhZzVtxVI3u+L4yB4Nl1PE1V5f/KZ5y/4TixtOER/FKrLzLKXtn2tDYK
WdbwyVm2+Opnup8dEaDLGgWCvWJ5ZhzZ8ZX5odWxoCU5ihQyU6QCMpEJM9oKs0OUeaxwWDidNOQF
KH6LyKCYJWWPthDkGEvqmDTd8jqip/pXW8TQcjq95/kKvqZ8oQQRh5ArU80WbamlSnjvoTA8u6kR
vZ2/iMwV5hu5TFFGyj888OlF8n7uVd5np+3GmkNoaIuXLzwXojbwf6t6V/wKqdwkhZV8OsVHeXWt
EqvGFq7ot+cm9HLICPOPjt7a3vNm3XLkaQ93DG+zpPexM/7fzJAHcSJxENQl+yF6becnz0LCNfvj
/wK8up5w3xkaXceZC4xS1rLrtUWNBIhbTSyZGscaKl9tpeGcf1lJdkOSVJmNbUjLrF8Gcotmsqe0
rgsKE5k4fjASA+vh1Xfl+n7BaHJnkGViGoljxaTjBjp3Rs/dsEr9cU3xm1Wa5+fbGdGQr8mqIvf5
TlyDbd3bkhJjBLlZsUREx00QpUX8xKCaWXJvNG92tnmZz5UibZF8Rz07aJU3giMAGrgq7J2FFzs2
jsSxYjyxruf6YsMHxBX8/euQ74+GW0WXeMft5gFIonjIkntevWbZh938rquyFl6vn2tnyuF7+uoE
HBIJImpUajMBROsoZTxvu6I/TDvrX1mJ/8fS5Qc2jAjhZyxrMrTnKvo4h7b75+yoZmS8Pg2tjxRn
1tIhfAxkUfsFBEG8cNHhVEWpfmt4EcMJJH0lP/uFQq4Fvo8UQMbLM2vmn1UmsnWHkW1h+vzDHOsD
2nv3odegJc5vuGOuacTcOxW1rxEHL+lDErcHgJtLeb3RhDH9yYko7Lj2NqtJrz4jcw12KO9QBdao
z5eUxF2+PnBAFNLAaGYNKZeJCe2yS3UPa/b1EXSWawxh3FY3RE7tzV4W6j75hrXtss+SF41u2sk8
MprUTGtEwD73MTnDNKL7+wxIQt4CsuO//kmZhCRutxjQY314mHHJr8xjy854n/Ql7gjCqz0nUJD6
niS+tCNkUvUegZGEhzUH5k4zL7nED0JdBBE23n5juKKuZiLdAf9wjdKAIGPUfsxkm0OGNjWEiwiS
gxmAQTonDY09IkUMnHgSdnEH5Osc1gE7JuHnpuzn0n+6Jo9h1sjUr4s/itUryPPFmQkfj5oNbJji
xO0vRgvRUEdD5Q8IWgbC09VfuVwoQfwu1d36JHgle18LMfSckOHbOtRRLgy8b91+WKbd7vSBAsuY
mll5b67zoMUAjhk3++D3CSSPqXY+s+8LcgmoQ0vjFdnUDCgACAqVMGO/rgXwBDGr9MOs5M7w6Yf+
RKP6UvtUzrFrTmj89il/2UoO+KxlEqqvxrm65sVfbAS6y1T2NBH8ojWSnxhW38Dl7N377GltA62I
yRW0CxUf8gH3pUY9ses6hcOZjm/IXk16u6ZZiOOGleqlDo8NoboZ70j8C2tJak9pwu2fTjv5Kj+w
Pn21prrsNS43mvLX6a1mn/ezRT/cSkx5vpXmaskmXsPTItkHEPyzycyvVoRRamkboQlnqKFibT0O
XD5kjDmDPB8tE6rqfVepmC+zJxFspgZm+43KNMDQ7qxIGIoC+o6BpcPicP4j0ChhJwN7B4NE0n0Y
nrULctA6f8N4Ccq4yp4AiQgDUQwXDQLIlm+UmY3HQZT9fDMOH6jMvIhfTX+vuSJVCRE8XdtsHeLP
N02l/Ng93Ht1xYueMVGi5w8PwDQ40+j7GXqw9rndM5KMfBYqsgHJb+t/iyHh87J1G9O4E8pFReP6
fYxEJWUVfoT7VNWrC1oYyLAcTnJkhfmSZuV1BxraEOCpXPsSBVatehsV2oFxqiPFhUHyVq6cdzgf
AA+L4Wge9EN9e+9bYMw4rIsSSb4vPLn5d/ailalsg+coV5mLSfsATlSSqgIBUQtn//htTgr8OQKw
vClL/qVjzMa7Qxi/qR/IRyJUb4i10t2mO9qrwsI1VnpZtwjMTwp2vHxSXQeC042lNjtwcTDC5q//
DX0ODVgS+5RUZUuAbQcfGsHh1SnejOT41IBxp01xS4jM1NimCH71/2L3RWErPItekNy43Xps8ZJ2
HyxgLfogBpTb3zUrV7ounlDX2J6Vmp/JsiHuMfuyP4HaeDSt6vDlLqePPvML4HJBid2XQJioch5d
fwudMBUihnMeSRlgQ/OcEumcs/QxxnZhJ0tUz2P1bw4J+y4JtEdLWV9phiFc5oZWEJOKI2OTUycf
diaMc7TVvXWLu+uk/GixVoAum851zc3sLEb8G2AdKFbsyS994FEz6zgPW6BEEBZYeDk3njXLI9vB
Do76Xi/qTP4mwGjrFkcmo5/tIeYxbIvwuFdqJWwH/P+1sAOGU5eImj3Clz78Xx/QrdThq+daIDOH
AzE/Fl7Ly5yi2aqfXbaSXfekREzn03WErkIYIYyNPVMLila8FselG49Uoinn7QuHulD6ZSvNkn2u
p2DLE/puEVKvIo0fUFKrwuGKAEBG0ucwbi8C4ULlfCcGZmo1GkmeQm0XZcqqianwuB+rj8Mp3D+r
xB7EUrjgpZGG/ZeHQJvEG+e/mT6m+FtdVuSAaPw1p05FNQuxP4oJSK72+ZIjqzghHepcB0+lcPxU
SIwxJ3ZIbMtO79aYsKs+c4puU/u6zKwZp1RKAEFoBJAW91VrudLQaRYBwlptitBxC8X3spnJty0K
SDxR40f2cB/hzpVBKSA+bef4snSF5AkuVxBeG/hLQle3gqvxp8Pwfg6f3Y4zfCC5TzV7CdrDUqTA
Ktsb6IKWX5vaTRHFDffLlMPMBO+KQyGDAkS+c+UrVB+nSEFEdI0DEkYEHLkOPQVNt5fRBwoWXb93
XqmnmidkNIjLSdbbEZ/PcZk2YcFAhwpy0MCKt5CF+3peuWDFDvuwPbnOCrsNkuds+PhbJ98SmCSC
KV8TxaE0NRLCbas7wOGIjwyxYWp0eXlmUo00KUJk/LQ9BFydowB1YokqG9Q8c66E2Yn6fkr5l5Xl
JKZBUQAOW2IUp9O4E1qCgEtOjOwoSFYtD0JrMg/JZaB8fbhI1JLWGcXp/gF4/D/1VREyFxXZD9HQ
4RXop+RBqewA6NBUZFRTA0sPFBJUu4VYZ2hM4XF4/NFYm65I/oJZrytawoEl2qj/5N7lIkUnVppN
wDcVCplR6nkqOijb58YTBb0tQfJVrGXdNpkh+jkk/YFQkQcSmSUmx7B/Z4560COnOJzi9MP/cjSv
D36fEQWlzKwzX6c2NS+F+lv/0R0kOAnk1vrfyso0Jy5Ch2gQs+y/6qsedFQBBSC5uI+8CiNxwCKA
Zj5xPe8q+YkBFX9Ed+tzWVd4L5YrCCe4zmp8I83tfxTqS7hyVOSq38sSge7KyTtTWwhvF4W7lzFu
x2Ra16mlYRyvenPH3EUfAr/P2/NCRtSYYYA8cR1mAaLgLCLO8iVikeC4kgNLidFW3HLpmJUoYJoE
vaQwLruXrFeaJMoz7CPc73n3/9wI8ZzWgnLI8obAIsoSN3WXR1L51WvJb2XfXWmsn45prbLbZfyp
E0SPN/wI4KjbxVHrC7L4psWfNKmtWffnNUDyBPHYL18YRHsVZZH9ckCletItJecVsoGGhs45Q+mi
F8MMoqxbqaiNZONv1KN6mVFp+YQcrMMN2ntP1oEJU4nrFjb2/VJnfCux/vgVHRHeQqKuAOCLxAc+
ctnecH5E20KgdQS3BwOXeBd4M5daT3dIuLWLW1jsT/KacgqYgjdQr+3VsOOipj+kPV2Hzye/cIwB
6+5c8oT0F4OvDR4/3hOrOsJXnZ/xGU8A5QwFmBYAtKw4V4PZmYtI5j/H+ZJ2wZMHD/tlQ3g4hOLf
/Yn+RZJ3Sr5uw/sS1XBDiTq+hYD6c6x7JWx7sw5wBrEU3rRZ4hLumeot+XxOinFhvZ8vzwJRMAKM
kKofyUsEgJwpyZAMy+IemM6lUTFwflYzacJ9+KF9azmntu1eMxajGEpMFcj2dVfdvwX7IwQEPIN8
4fOnT8gC2QwKn57Ra3p+WOitptRYD2Aka868ZTCQ4tOtUHsxkw/YcXilG+NI1psO8DZQSyqKAG82
nFRLTpllCP0O2ka3rQhwe+B6sTbI0xFwQomH4uKvuOGHQX3wdm1l1sOoh8UN5K7R8uoOJvn48eGR
DCHoHpHSwFv/yM8ls8j4bpzoljtqfnnbemriVIWy7TB5he8GByDdCYforHv2zqI85D34tmv7Fg9M
9uM9SPU3mrzeHMfwtx0Q3sXieqi8Asss+Pq+/JreJCrrDEYN5yZ1kdyT9TtklegtiDgAtBuGNb5B
9cZ4nPvsIf9Y7GxfWqDH3QuTympeeh3K2ey3VMoL2GuW0/yyorO10Y+zCTcYs3a3Ap1w5uh1hv79
EKX6f4LeJ0tj4xlcUgue6QSBmUQv5D43NlnE+GPWdYH3xhBfzhu3RJcAuAnZdAMBhhUMlxCLA8ER
R5ZN5Ou/brQdYBElObtWFz0sJe+0X58I49buxZZ/MuhLi8bcpongTNPe8INbv5lyioh1gY6pKOtV
AD5IDSDwQB4nlL5DAVtnk+iFM1+bEvEUAHz5s0CrsmM1BZeSFy7tOQQND6wuFxhiMW1lpyDi0472
VGHBvCO7Ljvqt3Fbil1T45P1UbOsGVJSp6wL6RQN1GA1Smkw2Fc1hlDP1k3NRLuT1gYf1hrFDrws
JGaTYnQUW5x5xM3sLK6qYvt37ox7maPMNH2CXF3ZT2vnmupOYdAodb3fN9y1cWqWrFrVlkUIZvbs
L/w8dCrMvB9sg5GIoUqlRkLFSreJj7PJmFY6CYFQAidxf2NKhJoLIGAxd/H724bzv8XOkSfHi+7P
pFU/FbrmhRjR/JboL1V0jP8Vt/hXt/M6tNS083ZuA7dQCZNuUs+JAgwdh+4sVjxAIjXrWzUhtRjQ
1ZCMYuW4HsX1tpk7X1SIMeyUcknttxmOs0qtvtTPjZI0ZD6oMnyGeQZ7/4xfAu3X9rl3vU6R8mpM
7kOQYk8QddyGDYmTVZbZU+w3U1HLZ/L//EQatMh0wznf5F1BKNFXyJPGqf2PW3+9lGYABPVkjSQg
c+cvhyrt+1YkmPYhT55Rz6Zzjz3h2bJ+R1x7JMiiBWvLGeprJvnJwLnNkRoO+hRLYv+AV+LsEce8
xK4OCpPO1hWAqfr1En3tgKuubdG7MSQ4KeAd17UM0YmsXnO2oziFizFnZs/9gzN3cnG0k6a6AubQ
xW7Rf+4rxqrvvNPM/AP8U/VmNehtkj0nUXbhvZpM/eBJUSrAL8k9GfvywMWSNVX0KSYJTU1wEDtd
rn0i2fPtOJTFLB+xVU7qaUBOectSRtdPvi99lUrqS8MlAHgD7gcw1KT0r7fdIjfGcbaVn+Fds18z
j93ms54NIkhfur44elG25n6UVx8LOZ2w/PAJMRYFTv1mrR3r1uk6FFAI3EUOT/HkhG5EGUgOs9fV
VDGIf3qGZVsK6CtXyJJajuP3Lhbe1614j/6hgdnQoSpOS+6KTJnCDkoOzb3vUpqA374ON0KaFGtV
q5rxNagN7dWYQ4f2ENqtSc0fT1MW6eusNkz8axo28hBY+tHaopNuTH+cpCFEFV34+PBc4ayTNSMI
X8mPh3REmy5UMurMEqiaGCVdLs8a4BkqRvJh0Thv/hz3AbEVqppKOjONxyLHiZR+pnXL08s+wPdq
loUREez+cBYZiTG+KjG+pmt+9NhTxMODMHYLjDrPqqXXdeybXMv9rXYkfKEmgkWgzRiVZHHvyeL6
D/GJc5MWIyZpT33NdE31czyuTvkEElocgZxLq1dOedevcKpqcEZcFXkEPdjpE3JpJt0NInsoThHN
eIe35xhLsx4ZXDLVfVRmwsZe0BIWr3x0Q93nRoCdOWKGcN3a+BVNsSYbreHTrNc03UnqyHcxWedH
BouYOsE+PvlSEiUrUtVAMhpHj0YlFwbDwf5sGE950O2oBrOdqmSkf+cLQifuomrueDkJCpQS8FyK
QeznB9qufLJwjPXaRh1MxKOwaM4qC/sXyje5tAJ9kiAsWIgazrQe3lcUBsmPutL5muvXe7luc+Fb
xSNOXXtSKCsVzOIgPCLCR8ZuxWpRvSj5//itvCP3H+oh4auBomlHSJUHAl6lWKaErz1YS/vThIQR
j2n3i0SdgWu+Xb3s5lEkOFoGNf2fwQqKKH1L+tQqzKc5VCCvEAPWLpBEwcMcTaaWMBDDRiZBqHnB
PjTzVb4bhmpbZ6VI1dnMVCaGOvNy/QGmOk9jRF1XLVCVoobiw0WU1F7Nhvf+R/2rC32P8QYvgmcD
kyuqvCfY3B64iWqdY6mWpXhMhALPXNWYaCD/cmbkIU/yjo3MX+I3w4YSr1Z3TlScXN8QOH0Jn6js
D2HFJcUDF+2f8QnoNqz79Eo6URHWUObeh4zzQdAX6y7s7Igs0qhjnc7MmL38O7J21JGhC++DFQP5
e3Hyg+86Wx8UBK32Tq3hq4ATCGKJDPYeTGGjW+Gkx4BisXalHlB0+A6D2/XLkD/kB4M589me+S3z
/y3BVc2Ha9SlosLRmH/TsprpAteAddFYNTdzoyCSCga/JHt/Hx1L+O3YsxbBssAOXxpuy+gcNFJV
oV07cTXG7m8r93sDLTY9/bwt2tOyvM9H4nIeegOh8axWHZVNsUtbYIz6HRn+Qh1JYPQxgzbQl8/s
c5vEOSz8ir/XsYwE6nZggia8A8KjGRRdZS9xsJRNnaaOGL+l31eFTAdSuUCbCrKeHRY8mUC0Dq0d
yMTkVQPSAXbdVk6THQgxLHCm55VtU+wzdqM9epQoSdejmZ3tlHlU5XX+isRU6P1AXPH4RdspEZIs
w75tyGSr3GQbxT5H5xaYQBiSLPI5bKBu4AW+y6AUI3xDBVLJYuTyH4ASRkhl9zBWBMVgS+AaBKKs
+84HGShDwhNaKigIWekHNv5hLilupaibl6MaKuPtdxNP7nzygnxmQsKW/RjHEK8IN4/UJq+Ma9GM
j8UoZ2Kn222A6+ygI5SjEMzitsOUaJKTCmnWBI6ROGIH2SS6/Lz699GU17dVBbQUlMoJaNiQPHqC
t76oORjwj1zUFJyC5zpCsQKMkHnj34/zdjapShtI6sKuZbPBvVOkIBrh3yYkuL+PnPIiQ+UHJ15l
huK9diCS55soXc48umEZ/5pKo1GFNKJZsFJ+VY44MiuXPAQIj2iaMTjg8g2a9+zSxOlgqvtyeo/Q
6eubovM3L7GpHPJAC4y1oSbKfe7ecnsjtKs+swNKLfaUOf7vtc1/Bo+sVue4s3A4P7HBLQArToQg
f0OuBaIz/9S2Lp0ghb+uaqZM100NKA1tWAGxGLFZu/9Q77zkGpAoBkqz6hjS4hBTEVLJBr/iIKru
G3n2YMJytJOxHz8sD0Cn/GbqobL0T2Ck42Gga7slsyDrihb6OF4uoUOrnWdrG0rIoGFS2NkyxHgk
EHtCwhMOivLy9kH6lIYXhCQ9ILdSbyW7Md9qbgWfan+rWCvOCv0Z3lWcykdysUQjZ3K5GBDrMsti
eG8fWkdZVFk/W3Zy1BqxdxzGeYJ9QqPhLsQ0liULq6/XsdJ7WHlCK7g6UwR5LkXl460aPTHb0a2P
DHZ9Z4a2WKdeESFCGoctEsCK1Vvct8tkkJIP+Ssuy6EHsCD/s+d6KjjBl/WJiTNPF4FIHeEM8bbI
yqhASAZ0bP73e7uo9gf3V5hBGMT+2rzhrpnVVNNCguVOlFtclhtBY6nXw/JK3uMwQZF6NuCaLOQn
j0SMh2zXWFMZeP1hI+UDHMb5hsRB/+T9q6lPTl9MdKfBMg9Zwe6CnpM0q6V0dyR3YbmFPzjRqLii
2nu0Ujr//jqjaYE/f9D5RVn8pWr4z+xHYVW5iDXVef6smwIjiIiDT7lJ1cx9R+WiON/3FKzS2+kC
EgiAts5MjfZ0Zf6Q92qL7LKrHXoy/wyQvuNgKDThca86yIL4OKlWZGTN6MOjiGbyqxHMGzg5cT3v
0AyDdT3ib4tyn15YHBMlN0EPASbsfCPT0f210FAMRYMRtUfarTy60yUou1evtAtZeyaJ6CDAbgiy
GjhMDGl5LC7WyltC/LqjJ6tsT6EUfwIN50nJsXS2eQeLR1MyBosQtXLqoG4VQfXdPWJHVXGjlki2
AJ5Hr+vcH0BpwhzA2Zfpyvr8x37gzTQKSHfJ2+NXJCAWC7ncQQZnK/NNmpQ0tmvE6+rk0lePUHh5
qR1xEfJt5+HDdbXBWIkvQvb2VP2TbjuW0B3Ju+XNL9famm+hy/BYQpJU3euyL56JvxtfgObcJHBM
PjrpFWIjc9NHHiM49MPl4mNfpfAYY+O8u2pxGBDJxxhOBzeakloxpZnHYN5GtoOhooIXrUYi/IPT
MqmghN6BZjtdNJXkCwhrVUyskbs+G7yomofctAPp0dvbmOmdzu0a5SvicKNFThh6VmqQhwI9ws1/
53qmTptCINUxwWSNkxEXqOcFr612Yoq2BAQhKPAOOMbWkoTlCbrq7zZZv3t/iMhP6/AuFkUJoSxj
NAi3344SrdmfB8pnbW4Idli6GNHCx7/vRODBAjmWZ92ZxygpHWuhkJUEYeeid+2Inc6/qmKFlJ6Q
atNhQVd/Kf/6BEjCKa3IX/r3CfNWR7v8MrQiJuNesfJSOLcgNoo1Lq7ceYwcA4TUQ20faK7q66Bx
zGLo3sddKnIbVmTpX2G13RRsu7kQzb9dGs86bZmHP6JDBWhdE9+5Z2Qda1R2T1/1WKtNVSojwpzo
Gjf+9Z7TE+WIV+FyGArcj6jIGS5EP4n1K+eBkZNOsndWtyzNKJZoKoyqkV/rx62peSDKLOo/nGls
UkC3BvIoWQ9YSnSXQvMyKYnUIljIdIdAkn5Lltf77DIyT9h3PtPWlr4aWtZDF0wpuoVmc93Gyrk5
4hC5Q6xSK0LHGoxPrLfhMBrANFpDoFEL5UeQn5ZhekRCO70urNk7hKXL3eUCGhBJWj8Cb0QHy0Gw
Yz7ZUL8UupeH57QyLkJlmQdgZ0UW2rMCfXg4XOL0PLAGIMn4wF7vXOfuk+NhVNapcg3jmaUGmA+6
gzephSiCzj0/P/Y3c5R6aIAnQWbyU0a0zGBARcWOQqxaOPtnisCEgI8ThadKCJAvoKhrlaNjtog3
NVMPnme0+A9n7IC/FwWp6UQ4PGxisTciIv3wUKc3+iji4n3NHiYxmRwE2ZQYSdsqNYLhQKUh9B79
UlQyZ7ig1ag7G37pmUJHhUESah4JZavsorD7RkBgOIZpa4hikAZaJGhAUqzWvQFH5rOPh9WbFluD
IAocInME1AmLVeBQxP/iKAi7IdfRVPhu+Uc6HcEy/ZUFe8/1pv9icPp6g+c2976IR55ZGpWUCanR
med8xow7ZcdyH3hvTya5kkX0ffwkQd0XEUcaEPigkBh66xV+SacCZ4P8B8qHtoZf8DxJAt3TH181
wTP3VDWeL4VPGeq45Kz/kWfK65jemT6MKM4PYfdxFIpg/fsK0BxLim3Uh63LqocRQTsPwgUJtSKE
6vchegsFMPcprAHZOh/WncvPrtxSv/0hDX/1PnMJpievgUhsc2LG2ImPD4QpkEhk260GOxKtGPaV
e29i/VFP9Zc9Q4jr8PUTFAKUVQrY+BSeJR6Dgzn7Timrv68/5nhzzWrNvjdXexLSBLuR4aRP+wxb
0I/oK6LI/0RtyiVFz4m2t/rFHwjY2+qNJF8KMF3z49usriPXcEOlpRCOjTik+HbCCSLgB9nzSeVY
kUZDHdoTGMCMrlpaPK6oYlz0LAYP5jDROF1i9mcsJYu4/vXzPx4XJilxE71omr2Lk2j8K2HjqZWv
ShEzg3MAdncBbltvDBJkhYhI0AiRbT+PsrDI8SaNA4XvnenvJw0v3widfUQvZpg0c46fp+TG04uG
wqTkJGsnRvhVDhQW3XvwrypDezHt2xGh5uAe6gEnOI2KnzwLJMRREhnR/aUYSgIjOADph+pVOcVX
GTF+BbS8xnATU2M+cEA6L0yNwAFUD7dBEY51DWj17veWEz8HeiNgmnABMjCSChKy/QxoFBDY+sk7
MnaM6oXWhQGl5HnBNetVywyykq8cjfqCSKn8ahS8U2tSZUf6mBGtEJvdF+AU9dh3F3yJ+cXI1A23
hzOsPx4vk8tj8K+6KXmgQTOHWNeEffuEbaOSP/P1JmBmMhUf7lwl2ZJd7s6dsEoWYFCqGVYs6fAp
C8Qaocxv1x+2Ixft6k7PFce5KPgBeIo6NQtZHMvBmtZrqsKx8iZFWVN6Dm5iIn/sqrFY0eI2fB/5
pRLmZfo1UVvuKV/JFLInp62RbqOGCWCzbLQvuvy00mLS1PG6xjRcGfU357asps0beB7xON4+uz1K
ELLk+kHekrBVohC0qAJZKiEIGP6V7Fw2IXCSEP9Gnc3PFqWGG73ROr/EbiHmC76+W97q4bLGj4My
H355niWs1M33T60QLXA8vrOYgeym/vmSuS8p1rkSHkcExoRknHDIf0iJFjvleyUVc3+UI5M/o4Id
OweJal7jV4nIRzVqWW6yxaZo/PlyS1+pskJPgDiN9/kPFE2RUW5LIjYwV9GKIZvlmK5XBsIsET+5
8WCbhe5uNZmTw0bB6jCTf/OoBlN3zWGifZUPZyS9A8Yng9iUBie6oXDxlxBvd4ySCRb+mvFddP2r
LsjjP83YtfTocNVlSoiSQOSs8TzX30L4B1/wB2YOXzAD2FOZKJwRf4Qz6C9o6ktLw+UNA0fiDXK8
rUsIrwAYUSBqJ1JS9rqMFWuIPD4ZuwSssNV/SmpFKkEwo0hF4Rkh35HRh4AgpsS3nzQAY/nf6Gaw
sUCE6mu0DFDhx1LA6RO9l/5jLBHufs5Ze+QNQAkvaoTx8S3nPx+4iJxKn2TzETF6CGPvwrs7OaF0
y+ekTzDf4g774PFZgNHgn4pFvJNZgqjIk9XYQzDSXv1ZXJKKnGm1qF/UM2sm0k2Ft2I9oZWRtZbw
yOt2DbkxKmMC1ekxstDyIbXOqI1Iuf1RIQB0H0BgL051/gba5iXCuSyF8TbZ15OMuS//h3/LToap
72Fj5c1MA8uHdWaj4FEjqR1sJCNN19CENSpcpN0pQ7HBb3E5zDP2JzrIyUAGBgPFWN7smzlwPlcg
steHYrqafnTJGW6bqgS5yLVujbABuUSe99YUk7Z1W02JHcZdHsvWsAflX3XuzDFZAjO2B2UpXjwH
Zk8+mC4OBbgRKdnmcqOYng0ibX1WegxiUBbzf/PT9PFPFojiQtlVprch5tBk5ntspdRbmSRjVrqw
hp9OAfShTaHel4GelFb+CUvxmTtfn5df13CdoHYCwP/OHI7UMADskwap3G7m6TFm2cbkGLWfquf2
T8IJJO2EfgJAgxrNY8x4eWFquVXuW4DfYqnErgw9+BgqjXxXW7JoWyJ7rNy5Qjc/JaTWEOJZRMPt
lcI6nATzydlmCEHwCs7F3yISypB5Ve15oZmWKI6GmEsYc53QBPwDniR5aIUgM4Yvac2qqXAJaOta
8ff/IuIlvV8GsGInCdYbBMJAHe6Rl6POW/fTJ4BKW+9v0+uoXqiN/JCJZXmMhD5kts3JviuUtsJV
xffOW3WzlcWm+iUVd6rVouJpyXZ3mcAWz+xuogEWkKJZEkRLFrxL8ma2vl/drsPb9+5Mr6LVDCY5
11AKUCU3N5O9YREhCQehGcOrKourhpSgiMijZ7LwTdpv/kxxdGTT3MspyWV7kArNEQQw2DOQblei
2iU7l0DahyGGt1rRqAFDdDvVB0P8eAgZdjUFzmphBNpx+Li5lcYlb/Jkmxf+DePBeQJIXiwcOi2i
rtZ20RqVIw0ZmfDNfYba2t+IoyQKOKJA40ouFpEO+9uNsOJ8N69pw8U1ultK010Nu0K2ejeYj6Di
OTJ/eeAi+FMsqHLm1Zf9J51JiM6lrMtlMPsaqI/XUSlHjHTgQPdVTY8c5fTuqbZ1eiKCeWI0VnEO
3T2GAvbJqyQzEHO0MVfnR3N2i7CrXXKI5wMLZqaursGXFR2qd3l7Bf59XAM1zR70XOi1whq5ovz+
6XGQb9n6JODb3Z9UC/4FO3bMX1ULuslWHqVRCNkVDdNEzJChjT2dwQtPGbf8mDzmAqNwWtr3RD4v
0P0hGIhglBw0uHeSGHx1E2kJAKLWlR7YAvTYHICeX9JEDL9bS8dzvmrsIt5ptTCPNo0x7MLUIlHx
hAEqMiZB/rRHG55Lm0YC02I9aAekCeWX+QsEWclrXildy+tZdnCRLNY02xzC9UxLrVf8yUpCEbtr
cHfPfiLatHvB3kxgr7jEXhZVSuU0p39tSuQakTRi0DxReUDKGXYpDs5Gdix3edeafhHXpWLkc26q
rS47amF/Acb69a9/bT7OmzAAoYis03UyAmVA0b6oES8rXO7nNfa8GPYFwfyVWMnF43soBYg7yZBQ
OlJKdAnI6q40swLvWL7KNfgzw7Mjj49Kj3U/ZoIOc2XACBn3ilOazfZwY3YRvQ9R1pC5bLKnwPkM
XjDIzDDSAq+gmiubAJxi9cI8ta/u1sv2EF/eZbBs02LLmj8xzsIi9kwQ6Pwi6O+CAp3dYvvd1MJz
cadGI/pGH3CfiZr1DQgVZ1LAQ9VaJKOsEuSmhmbvQ43XR/t5wQCvfQwAl26M9taFUFGkzkIrJ+Ua
+OxdisLiNK/6CDYadsXAIcnPgZQAin6e2FvXr7YQr5d3uJuRTYwZ5jADjbliFik1/gpCOXo3v37H
UINLpz6qWXVUq8FwiIEwpgXzIO77z7bv13vaih28sxwm8FO2TbK/Q6zTEPCYhq0y1S/Bm6bAzbMo
S6LZkEGk/bJcS8Pua+j2cSrISmXSR99qk+OSE6ZwiCCKKN2/J5Nr2knKF+6xljijhho+wIb73YbN
xn+Cb811K4nL8eEwAvcCVHarbm+jD/FAX/y0ox542ud7z3QPDPLdTzKV9Z7Mzxea35hhPX4q2Hpp
GmttGTo/SJfWsvvd8S3rTao5/QA808t5PxeBDSJnkW4voFEPdh0IAZ2aBHhdMf+iUk856u+Ddi/p
CIBjnwhEght2YiQLIQfAqQktz3at7g1eLylZiO62jHd5VFwHMlLhgtp0cHJhlMt2Ts3W+5lTW3Jo
SjquHlbzQSn4rLEmOZvlA0ogYMqJgPwmLROB8lVDtJs32kRWSiDHW6OWOyCoX6wLUvVN3/ffBA9M
M7LHygbylc1cYtxw1eZn8OXsA0azsJIK4dOUzZleKZ3qmFCRRNPLqQWeyiSKHMS9TM4KU2C79/+5
d9phBbN1vahIZF+JbFHcEPp3LfcdwX+be7W1yIYuwPOdpN7514eLrI+pBXKeKtjiK/g3nvemd6Ck
qe9CVVuyknowqKtNwAS/mPMCSSiLgKRZxdpuRyTHRB3ZAMtoPoetg81Z2bcdmbrSzFj1YXhOcSkZ
2KHJzjRLIyTwr5oHYaPE+Po4W2c8q0TA878/0T/kEHDdIJvjKo3AmpZgrPHO65C3w3NY9O70fV9V
10UqCSSrZ9h6bt4Ladf8gWhiG+0hGxjAS41RzP/hZ8kB3IuO8I2GzYxUH6jqpAbBoyHp87lCGZIW
l4shizEfs8+cmDjPxJtxml3mUMusIn4UQAwLrHP07LGWh6jz1XdXvbmhh+Y/eiHjBWVwOVNWkIAP
GC+nmTGLFSaotH7oleIzWD6Dapklj1uO7F7QQLupCT+VAVgrnhELsIQersSuLgrUOQylIaIxL0ID
uVvExEt9eyHBtWC8tNTcYDeDJ2sGqDTVzlrf63MoUASjLp0YYXItiir2VJcABSu03exvhMm81wHQ
LnvV78tKi601aQ/esDe/y/O5SxQJQqvQG5dLhUv3Rd4iKLMKLWVzdw+GO95yefbupStoczdJQ2Jo
4ax+tmudtzKqnEhzb5jHvYb2xsSh/41rp+ByexrR7GLeorby/5wNADC7Pk/QB73BnGn4NHSsomaV
6OIm+OUbUD6UizOONVagLa25Lffu3nu+IUjfdsTb+6VdiXvc/HK2OfcQ3EXZ4c/IwytRkefatsOu
DfCASwioi3TQkHVKtnY0Ujyy6X9qGWizxBG1eSZTwvBFgF4Baj+Yp9r7JJYtq2p+dXMy9UddW3QS
S7nExHSYI55qunoxTtBYX6DUomMzf2cxdvlzveT9/A+jhI01H+QgU+3d+PVAN1on9FxulxoJFfmn
7r6mExkAK2zfn18bLCnMqkcUj9CwAkxiu/0oLJ9xn3SAK5nHeQrmn3ECKm8p5KacqUit+hEta3Od
O7QLEJpS9KM5oM66nDKSq3s7Bd3VNK+dWFQDuIJtQDuQPNl0kUMvJWRocZ9CSBLXNsulfwI1Siaz
OqJEIA7NIrtCKX1+uCvJBki+fIJpg5ye08jkdV7fj3zAKexOhMhazG47Jvtrc3yQMSLFg+z6R1T4
sQQ7nqwRVpORLOciNipbUsORhZdlSU3eh/V3cQLTUXp9ma0RXCYfn5BB9xb1V5QBDsJ6e0Cjw67R
9OfnH9yyPNv2W7LYE7pdLR3DpiI9+fJ4EdLO5AwlP76R+ZdnC9000Hc9BW/yh8saLCxuAkK7kxen
csdmscjcMZS98iwjrzY37Hs71Sx+JKpHeKkyOm1J/RSv7yRuO6ycyI6JSQBh3NV7bwFWi4r1DBEL
SeqIhDnNJw3Chb5Wod/XwELra5wdKkoF/aV3WfgPY+J4S8xDWnz8or3yEe41230zAAP+RI/Xig3F
cHcGNx9olKJS9QhQwYd7qoIGVV6R3HJimiFC/U7BOc7hD2cROK4Y7YGSdIWtAwtrmPFruN3qT/Gy
V3Y/gV5OWfRg/jJhcKaKWiWaiX99utFMkr6e5qGtJktST2SMR56uVeHsXWG7OUeVwKudQh5fG9MI
hqrsYS5G370Beb0ejDTZtZv5buBy0+h2rl+xwbqhXuRR0Y46z/61QymHV+Wr02QPa47sD5/RJm1V
1ZEecYgAGMlZaRybod2IPcgPSHdI7tg/mVlygITMukHwZqRbPc54Q4d5sLPyWVfwsaTlROKtXD2m
5LDPl8xuClpkSzV3Nzrz7PuOT8VaN/rc635ij8R0EUKZ6N8zoRuI46SJioXVLLg61HZ4lnIrXTCa
wYDyYsN0tM7JHxqVh8D8mKm3E+japjb3DwEki1hdYxYe2GEp/G5Ve3IAdbkS+kq8miRifs54PnSd
RASpqHn8ZnabQQ1Mzo2UzpAo98WqTxKtx52jGQWrM37pfjr6gsMLoI2nEUUL/NI+QfDgIVn9In94
zQIb2ENyyuks3iOmxyZvKvQ8lBSAUkhXQIyq56vVRB7hLddfQz2zjrv57tRIvlp6QEQoCTsRICkK
iUhbrU4jEoAyfvhWPsSeXEXGwRMbU32lEKjCv2JFU+OJqRjyDO/GYIVYi0hqvxZvvqThCnIn4cLE
186gXvBp51qrel6DuPBACOAlnAdjGNqYPRtzYTd9dHSKxudq0gcz+f0n2ecIpnLaIZJ7ieuOOnd4
eQr9bpcr9ravEnYNdR8cg/QcwdtJOdFfDQbjnsPkg/n82sTA34Iwgvm1vqR902+FE8OXXN3s2HWG
LOVueOscS+9jgk9vEWETjAetb+8FEVYlzwK71meU9RRPWHp99SYVAlIMgVjboDgDoDu7rAZx/Ea3
GDXj1io1rzh7P+WDZiW8BjNV1ZuKGej8JcUVji429mn89fgnNF616J7GJuQqV364+ebzG33HoWeC
938QCmGMiJKtgUzieIW1c9wMk42Z1jyzxhAx6R8rtb1Ky2j/Gb9tVsEG2s0CVZjzG/xERL9dZObY
yfyOR+/wed3hBQn+iJd9v0hAJxJ3RCBG6qpo5PclEVtbqcA3gs8FrAdyNl0JnZ1UJjDTOZgxrR5k
q5KM4WJY3xon4OyBV/fffkttpKP7yMwUtbc+WjCVVk1fGfwHoc9qw1G4YMEf394Y5qJJwM9sDmAh
lAboB9VmIach4X9syYIOeQtzkX89njW8nwrUgyHa3gCP2BLdscLJqhUfurKNpsIl4A1YM1u31KaT
QkAaSjb0yuDAsCXle3oH53RZuinzQbTwChp1qz6AXTSo5Q3v5P6m558qNczg5diJb2MCYid4+tic
jdSFn05NrLgOResxsTHiu9Hr9SVnJ5yjbpPum4xwbzasTih+MnWwSAoUMCHmumYPNJgwjUOx5K+6
ut0ZgnxzItu8DWb5WX/ezKf3Wj53oUWtWUgqmQWgxHSSJIFLDlURW2+n8yJNp7FYAXZ1jwR41E1G
pGxRHKWKyRJU0JqlqDGI+RM2t8PA1d7QjZJ9lvEQkzGg5W/HeAL/FjY9ihMP9YldBw696ZM6iPqH
ajd+48v1/P61E/bU+BwyXDtuPgOSdUXc2hz5Bbwr3jw496i5poiuStqT4HTBtdcWYtkPve+sVQ6s
CSBr0g3KSKOyVA1bFDEAkVCiT3DL6/MLyKeg4DDW4gZ866SQ5/TJZgLfjObY/JTKV3UWMBN9ue/7
2V2qZoaTHNuInxneviLQT5i1BejToOu1G0+uXOLrdhc6DQYKXCEujw5u4515jv+PYbbyyFSjvvgJ
hi3VvB7Qm2lM9N1yUIugmUfUZcR5lDy2xPSZAdaFiAZDE9jtzWSueDuFMV1KPmZWrRhMGtHL+Q7p
x9Av8/YORQAtOv5opfoM+ITa+6gijTBOcFFZKP4IT4li0Gwwc1qz8SF89alXR032kBpZ6a2OSuJ/
+6s8CikgXfFGEhfFUWvzfWre+RNpeRqm+7E/8NvjWkfv6Zfb8fFg21s3Dt8DpeZ+sRCwn1PX7q0X
/jwmY27yuDgTV7AplsawihGaeswdekwuF+0TkIuekAqd7GnbvqXF4DUwYeZMMuDcWdneVr6hWmRz
3k0fwecklfn385DNWNAGr3CQlhMewBaQWvpmQp7wU1eJG/bqqdnKK9z6LgCrVkIEWcL+u6icE18v
crulEM6NiPQR9L/Yoig70FQhRE3rNDlkZSWP3viZJz+qE5oT7GkaaYX7jjSxH6ERzlffmz+0zRVT
nrLt+gOzDqgmGe+czc3H6DFhoD+nrlPex9+m5WD0wvbXkTIMunsrbiyczDFu6Vh+ul+dxBjP6NnL
NzpMoz1VhPVx2mVlRbg9v9NAp1jR2lNlXBBwec4xYkDKr2EpU47/0Z+EDItGvUdeTvFiJiuXSTA6
C1XeVzaZ0tWKCgfIAE2qVwIGbTWNl9isjaJTb2xWsrDdqjjCWr+GLOFYmU9+GBeHP3VftwX7/J8B
idF09Kw1JiKyBSJ+m6zAhOHDuK6vAnk6wGWmjcjm24bJaK7RzZXBeBqCuICMQd0x9HaJunlCmtif
E044F91sqVXNHx4tFZ5AgyDtN0Um3X/YzsEFMxaEF30O3we/uUwanQBDb0DyXVBLBDwObUog45fi
/2Qw32HaJSdJJh7UKPJCK7JA+5Uf8Lk9MOtfWos9BnsdlOudh7/cIQNG9zAiV/xvqzqaqy3osCA6
iJ7/zS00T3vn0dp+b59N564RDUiUGwATWueap+6FQbLpKDTNSvvD4AZpnUvDVBRTfxc45/R9I3xq
Rqx/WXnSgBzuHTKhZP1FQBKRR8EjvX7/XId3wxXVIzsUZ8ixuVCtfIBhsHyg7aUXu1rKOHP5Gjp0
nGanpqR1JgglYS1wc2Aqe3o2H9rotbyoe60VDy8UfYcQbgJ/0Hf9V+Ah7mg8X7cmVe6zloYQE6yf
ASjx1JQFOyL5027QaDeFuwFlsXma8nOD/28gYhEynzx/AOLpLR2t8FeTkw/iXARCAxU1GnA2JIMv
t7squMW66LfqOYxMRawSpKm8Vu/IpZB6tDqG/mcZdwjDkt8Oi+LoG4GcU7luSIUHs/8F0HjoRC/V
xGYB6IENqnSuA8XR4lCxLutQEKYLv0F+c2u68BaNcgCuhszT/U7Iwah+fkw/tFyu4aQxfFaX+Mk3
4OvhfmQ02w2EPT+0n077kfluSC2np7WnPPxRitiWhJD/IpQtNubB4/OQnFKvcEXyVdAflwubhjCq
fGHPl75oK1cJm7NLC7nphQbrzV9TRfL4cS83qFNkjRdCHO1EM2c1l6EequgrVbbBhlKmtYdYuww6
y7I+r+OLjwzIJCw8ro4U7yevhu9fMAKuRJOax16U6mYQ8kPEG9+zHoDuA9bQoB9YhmzInPlSVBBy
QnObBfqeUIOPfCwtPf77G3d2mmil527Xr/3/ApUwAjMw0lmLOEKLxb5AYG62AQ88nzS8nOYR8NNx
FYo0mBsQ0NbU8GBT8KKBfgJN0kf+JXo/fLgnlG/PcQewCpsN+WtGzyEI8wREBTgsQ01f5CWYqlHo
N1VUpfWxIi05whCi5yYtQ+1EpGJ4eu81Nw7gWmvnSMaBu32C8fDEZukXZ5IdvJqLeCR7H2KG6RNs
Tm98yhau0RLZWP1+1txuznMZYKlNrejd6ru0kV6TGUDY7uhUGbnINFvQrtWVPY/RoIa/CY8ZH0is
qN1On6jFBVnv6TmJoAVc9fPUUptzGlfzOELp0vrzUZkb1hRvO1QgZ0gCToOYzYVBEgmrRRmSOduN
IrijwVLyWT0+szrGKZ7/fmQLePW3CFZW2W0P6eUNkO3EWpRrNvB6OIlTq1H/63Zvs00lkSDYkz5u
KOFl3oxLStNTiVQqySxq2VharrY+PqoM3eATHyBL9e2jCq8ZciGIMEMFsgk+Zq+0e5lQFpnrnPqz
8+mTxQVyMS7VmcO4WzsKg9BTZxGBJaxaIAzI/kj6zvHpVqmT/E35dyaya4iHQJHg0RvmqDxh1w1o
8f3NUvQBdNcchnxzAUbRyBYQ19wsm8/mPy1vMTF/aashxijBAKoUASct6Qqa9OYoBJRKp7pQvEP/
P/x0Y/csoX3+Emix5lb5zAfw7QNxdTZtYXRNymNLTu98Sc44S1jn/YA2tyJwHJJD61Uq5D02P6/Q
/o/svc7LsaNe/8KBExp7pRPlQS4KFavlEGXbSFmoSqVxUeKdU7gIGJEj09T5GfqtO/00xdbPbj2p
GDMpGv3BhMyLd+9msnWk5HDXaBpxTF2H2ReOa1+Dxhtmwxb2dAotzudOn0e0lQ1h5FKdYMuBiam8
KF1YRmN+BO+Sl/iPRYNMwuQaXFx/48WHRT6h/K8pOJQVyQjaWDdriXatG+k8yT3wyP4gx5jF1Okn
i0/ks1wQZhjF0VclpylPwBn3QHe4FUyCx2CDR+H0JD/4Y2nm1M8dEGtuMvwZvQ+7yht0t2PnsmPW
X2pkNdcjbdIz8NBiTI+jJR3CcuK0kv6U2kQLgIdsX/IxQlk5eIRpL/WG0h7qayGH+/8W6Em1EEFE
iBGN8XeZ/iB7hMSgnPysexFj9q+ibIMicy3q9XApCZIIFWeEBsSgBwKSDTqiWP5pRxCkkYOFgF0R
2UTJJ55vHfVuVs9/URKwFQd9lNU22z2ZmnoBBEOYM2nztnUGG9UDjMJ6D5Zo2T2LenZR+OR9tzGW
V4lvwBNoV1ytCLslmNdRfNWp38JWZeC/3ehI63CVX5w/O3JPGP1Bzy1kSXglLum9eqfYELu0IyD9
Llaxpc9yVRvehhg7RLETbHAdDQccKQQLT/B42+sPTfv4cAn4UqAJEWXneruJ+dAIjpmNxSwsiHdG
yx/1VvYlWUnSd/u/PQxki99T4zFQDTH5us37t0DaZtjHdTm7wTbmUJDZjDIScuFzkYcmtaty3tql
KhqC6X7HuwO/2JY1Q/XAHiJAyR1A+2e7dYepKifkNajAK2HYtbgd6J2gYkLlxQiuGj7gQQP+H4Ui
PlWl+sbEmI3JjUxB2YdyB/XlZxkjU5hOIpVty7A2JR8YtSnA+ZrpmUblaGDv5kAuss+qhmHk63SH
IPlIVA1Icraf9iWxQUFqHUVO6L+KFoL+iRAo9H4ovRaC8JjPVocBLzsYgYSArECIIVQBQlZsKxm+
TQ5wvakVRpmwet5ylBV0I6VuPoTn2SeMVedtsG270MSD3O4uPzKs0fkrYBb3uSad9iYK8YEprrjX
X4rya9tf+O04wVcilntNlGAw5ONrT4uikbD5gSkoIuBDa5XBnoHbj3u51bE2FR369iFEsBc9Rs4b
PaZ2PAD+uVD/D36tUXJkgRTVcuL0t3ccc+Z5yPYqcBLfUOVXzhIWuuuWLCmnprW8dXvd0ojkqsIB
cyqOlx/odAUfTekTUTlT3m6xNkPpc0odeT1+6n9S/X8zDdl8ldi7Ig8xRmQsbZq5SjUhR39oF6Wz
PfWKCCtSYsan0CDkeqEwp1iUCFJ2TCuWPRj0BwijeyMTfHi0xPLLU2kqmxfYgfmKeYVfNdN9MIGI
y2MkpMsIuBJBXwOH2F1bfxhXGtygZ3BsUHF0AH1TgIXyVFkIHHf0rgkHyzFMWe5zjCZavRsjAXDL
4dm6q+/3dPpiqFMcjsd2aJVmFN1VAEZ5fThPcNZMF30Myrnly1qQQMhO4OUe3hd5NNsaNq1Zhj50
5diXOOxC1mLFmckO2lAQU+/wk58CaEmMb4y7ge8VFcylpP/WvHrrxW8nda60rLAINp/MjPC1VzBS
YighFlf7CeDysmgbWLZSg+dbq4Q54/U6on/bORSzWvULnVdR3aJs3XmdnxmV/YygGkXM8qcNjQun
7oVWGEWDjK5vxzXb7xU9IPwf4kzMqqs1n44plZQ2XtgItQ/F6dwPcBYy9CZbl24JjX77aUeAkXCT
BPeCAd+RU6TBQkWuCaa+pR/mkqZc3RRPyo4GgWWnSxidpPuqCjhfqU4E3RyFNX4CyhHIKSn70TwR
8U2rLvFDum9j9/HirgBX66GqUcJeSqqv3ZhjlriyvIeXCSZR3I5UU3b/fEqLZ1fnuw5IpWcYp13p
F73E65Ey6f2U3HWAYkYNpBWljergkIaNP67koYkjuUZAtVESQwnYcYQOjgJ738qJOOFvF57djqnu
d8jQWmSDL1MMH8bA67IRC/1PtRZVJRrnWje45fqvYnrJypv87vISTiVLPBgI4TZ4wtjr/JPID3gf
0vUVW08Iu5KcTIxb0VWnlM63h2rRCpR6Yd0azuoi2Oq0A4m2vZBN//76j0dc1c/ZtYLSise5dNvI
DE9ztItHX9CRIAHB2Vd1MW4POwDlPc3NNqLPlfgGJBSbL3X6IgrBPZE5a1j3/R8e27X2QAK+4caQ
jMpQfo9Tt3bb+WkTHIAkXv4FnJ0JQAV1jFUYj8lgCWhPAT+0VihzF7WbBdtyk5qFmWTrjxdlZPSf
I1Lms06VIWQyyP3axmEBTZK45d8GWVIBpwCqL5NLR4EFPK6FA4JzzCSQhKui9qzlrT8WqrwO/tpz
ChPa383CZ6/02PIyofoKXHkJsRsMFzsiFYYF3hzNRQDRjpBgNZEq965WQJfxRrapaZuaqvwnhBRA
4sBxmlI4VWMAc4KY78emg7VzDxM0m9HHH5X/QlSz2hi/GfTQhkHiCTYOVvvfBisQXxLayO12D5TA
cRJpsybf3QkUoNdrYcp21p+G1hOH1eDfSNMaDudq1e1ZoyibOhZ/XZhs9yF0YPWo1aV7gKbdqZJa
o25xCyrr4eA1h6/YZ/Be2ayOOHedK8ACSfpBJ+kK/mCuLe9TMG9FnFNRzHseAH1Csg05e3wdEZLl
ryXEC5XSZM0rSs5g61llcSt8DJTCQKwWC9G3hb1Q5Ht/vJfTdzgQ0kGDns7z0jBqGkx+2IB7QxJE
5T/Vor/3NrkUOb6v6xWpq4hClvCPqPmqSIfEgUFEicII0THXLvqoL9M7XK1xn35B6FLWHRlZHt80
Td7UfcqSKw1ylJRMBQ9aD5x0nzGnmLaldcnJ4KBA3uZNiBD4VucYaeOptRHe7AeMFM4CF16PBTkW
XMVK4/jKTmFGeb2Pq94DoTpQPMAJaQ0bExcNspuGMJEzMp7VsHlLSxgp9PE6AGX328GsCsYmKoFT
YO6KrrdUcxEw7rvlWR0gPzXmbGtgxtFjEOCW+JQxYI0/Gj5RNIx/F+a8LdfjryPhQHNBoAo4IhTc
eK0eH+TH9yBatrzj8kncCPynJ1FVi29ZVUhcwji4iUHbmZfDLUtKkAici+5WZrlNHii0yd0Y4BFF
Gnx4F+je6gabVMxqdP8tMhKx+gteme/qwocIwgZZ9klJ0mnKwSvOUPeaBUeI9TkmTPBWiqKutq5B
fV0hRXCQlkTtjtkwTHPkXSuV26u4dXHrypO04JiK8RQHLyQvJvlRd3BDaHgE/ceFz4sIvE28P3Ai
fv5t+JNxrNZt63xmlcm3S7YW/cdjomexxKYqd8SRXbjjKRbge0boW6N+MoxXIitq4J7z/xnYTNaA
du6wiYrWgsi1vB4hogAXx1+sV7hfeppp/sTN7AHWFbyVTNY6ep5YbCoVmcGTvzr1z4q1FAlEFFpZ
TvP9BurQtsoT5b8s2FEO8V3HycwD7vZYK5Bqajkrrg2Hbeuk8vtifFGJ548kHXUwhE3E+RGven+x
d9scEklEsmrKjyb2iMq2kAi+b72NPMIpTlw+IX8Nu7ySXO7cYqO9KT97OdoSM+pNJpfvKH6eMYRu
t7YoB7QhMko8cwBZbi3FFianPEI6jQ10h4zZkQYowILXzNNA0JKwgKtoZCoXDQLigxLoa2IAtPP/
rpgvAL8gZGa1fPH5ZmZgLuQaW2XDXD17LnY8NRdCrIV4F1ERoU2xZqqr2Eu8Aj26IADXzWaUpHaZ
FG8wqwmYEAxi3IDR7myvLgw4M3SplOErv/W0bzQ7pDHxUlkdfVBeEAbKKWk1ndxPOqXzDyYNzHxo
OvmM4MxtOP/EjPtmt9iApQpS2pVjQOSS2iRvWqRCO+HCaAnhzQ4Fh9bL45uPkQgyKjovBa0/MA54
k9i/ZEV+C5+GQhYJR09Mvo/PdxBF9nLFbcReFzN1rAL6sS/vPXCeGe8PZQXLOh+mXGU7Uez0wb/i
aKXplJOd5gPjxLx14LAapsU7vpgecYgCtuP+fLWnMjiYeX2r9lEvWfKlq9OuJs2JEolBdP0lMwHu
ywBNVGRrdCtIo0TQNwa2Nqa+DywiLa90edCl4xiLuYtKcvjh2cChKRyK31hxwuDwLpLHX/3572V+
jxFdk2wTTHjlvq82fYpxroehfmtGeqq785ksQGxNF6hDU49HC9nztdUMnL2ST3rnP+KQv+5aOixh
udMUnyI6tYXA24kxWeYkGgLM5IBwe3Ui1xlTO3cBMbSLHxThWDv/k8kTB/GiJ1InHVpKKJtfA56g
aLuzxkpv2gxSymFNFQ3pcH5n1/zVINkCmDeEi749EVX+HLeHMflGWoAg5DROCg2u2Ixs27WDWZY9
kblfs4vch0IbPhExLrpqY8WoHf/vX123pK1GHRXE6mfVt6Bs/gaReL2EURq+jn+E6ZuqT2wd+pgj
FdokkYnsPv/aJO1c6cRIUcbLS26cfUzQBt5AhAYlRYETNo1LzokBo9IirmHLTS0oV55aug9eFqza
Rq58xC7vYL9d3i5wwMwHtJIrhNaPVcGCQNBjOmbs9FqFEAUAcxJVA9wgLWLYEIv2VVcQwdIM0eC4
6SxP0JxmqVABoFy5fnK35FDvWNyfmyG4/zMjXw+k4db0ZFUrxVBUgXHAG5V4FHvuOI3iyr/nsgGv
Qn3tMvrtUmw62yL6hRrZ+3VswrIKIxAJ8/q7fQTkFBvJMk6YGPIl/XaGPiTGBknJ+pmsSVN/h6bR
M//1PFyln48CngD7ucuC/g5qh/+4k1JaSHUqnI9Wt8jQR8Xgxg/E9M9sn0XglWNHcWMgu8I5/czP
Ut90ftUClKjKCK3veb0l58WNCrjo91rCEjDPP06pIBwzOGwY0xd2SbeVog8I8sC/RHY8729P5A8a
H5BteOhVPCzZpqTwgTFmI4m7K77qLF+5/gZSPGFqWyWUl0nd/YKY7XGyHHH3XlHAORjODDNRux79
eqo3BXdX6GU0uTQcn87VHKaSe89H9+5g+6/0abheC0wI3EA1PKablOoLb7n/VfC0dfa4uUPyhz3c
1d2l+JZRbCwIEYfBgmsAx1bF6F6ctWDVGUZ8N9aZn8+0bJdTXKAEzRx8w/PIbRBdxdh7LBaL5FpO
ifRmQXVEgFiG474gzTNoWkvhxEyy7EOULAbtXT+q0X62kNqCYL+7dagF4No/9WccYjih32qhGEvk
OZAsa52osQQJl4rYA95fwF1uuubglWyq9HpFIjDIuZO4qAEuTGxW1xRK6Yy85TR6ly+Kr3q/XAgd
uj+B8m7IkvHVFLteGRlP5qUEZ9YB0wH1B0UWqMfvabSV9TiZPw6RpkRbLn2cFkW8EMDR5KIzZ4VL
dNMlcLKv75GOLi8By4mbH9G6Yp8wy1StafrZnmNhBEaahi6amglQURGxF4R8PBBcQiqsd2DopAH8
vU8XoCznI5ZTVLgggswGUdH0lBkrdU8LqzU+CEmxr8xC3sZSFcdbRSgJYWmykSdpwYC/drJHsp0S
YLMFhsqK15gmNmgWhIvNvQ+KQXZ0n+E6SR3PMS5+behlUdzN2uqFs0Tn2M2XzeUmBQGgyAzRxgWV
fgo6aedmG4382g11r4v/oHsorBFIYf29eKz9qZGS1hnVrwqxYFjAKHzVlFh6mvD4saWzsqwsdjkZ
JdzdVEHATApq5H7m96KbjFXZbBtcBLhN7O7hiRgLDG/t7AlsnoUOElPXs1mgL6+FOOtnOkGz4U6f
9lLw8/uybIl4FqbvsMAKoylmN0n23k4ilAnoE22N+oyaH3eWRTZ+phzTPAprkqQtJaYIw2JCPyOl
2WibXTARiV9yioik4ANGsaMskwsRMxpWYCa3E+kHou2lQlLSpBDiJw9mDRpIfulk9K1AjvmexdON
4hFxJl/xYvlrEOLr3i/FvsCRn0hf9N706H9qkIL1T94byTZt+4qG4TyOzx5OWOgJ+ltvtzqSUpIs
W5RcotIP4IvH70Acsfa/2h10Zxm3CuA8Qr+a5Pi01sMi542ygn7zyH8Zl8aNKkUZ/WlA17ajRwa0
lk5VN2KeGIdcjf/aA7ZFov/rJz/Apx6Y1JiXlSk+5WGbwxAO+GRgD7AkdmgTHqMiqgeo7T17H+dz
+Bx4IFy3dlk5GYJVbpyYSsnLq5oRVQpBIzSb8JJ3Pp5eXAoSRyl3z7wQcH3SUZt/7fJjyJp6r9FB
0peR51dwQsZk0XtjzjMKAXzk/cke+UN2L8KS2B+mspHlgv3Yrk/7NLX+2ME7RemCQvEhrEU/2P1g
g9fbhuDU4dxrQoZJaYRp2WzMkEgw6VbOIIJ/4cFOdcqWK9QdI7ZXiwmzfBoAhdvjLyxMyTU98Wls
8JCD5YY1/iWP+xOns+wiI58qZv0vjy6t8uV+IHpDfwr7EazX+Zw9D0M8M2zGWdw6CjURO4qNktF9
7E/rRLw9PtaSjkbdqzz2KBjC4rAO260vlfu4Zx/co9NTJF7tlDmd1TcXkGirnCdUGmcN8mHZtCwk
fzPSyHM9ViG+eZDfSnwJ5tcajPBscJZjFjEyk5fTWvHIqSdp+xc2VjvMes66XPtBRn+j3j3T76He
abuwlzMsallqMWCLtZw6lIazlY2yD0dGY00GBzkrYJbwdAe+AnuQouAu69zdPIBRLvnURSv4vLTi
P1XvREeR0kHyAlXyZUOkD64PySN/QeSkhJwLQHKXJ8uGk9pySb/e3prIBvCdCkgeo/ZW0o/hsanb
BCXwz7dOx6gzjTVJ7+/y84yXoELWYadSJJrCdKjFCO2IBsVtfLE6uIXrCO53VpN+hw4TjjwCvyLo
Ktw5PMiglWq0zbfRHh3a9LAcJI2LohqgXd02Z5OUdJtKpOYsHbEw+98VnkzobOltTlKfO9qsYkyu
R6O9Au2bzcOVKs0hjR+jn2RBjTGzn67qlhev1hNNNFAHl0r526W0oN2wA5HsHG1vG9/nLslb9/RR
KA1dY5mHMD+NxvbDnjN/Xl6vwhFD6ftXj1IUFkSrTjrlYb+Qqe8Al//+LZL7qdzqZWOHg4BtrYuV
g+PUnsT+d6700Zr64lWzo/3eKo+ntapS9MzCT9F/5o9zI4Tpzj7oJf7RKohKCi6qse8KfaYo7cfH
Mg1xDWdhgdnfOWSumw8eCxG3Js2mp8hlPRILhEHw2jFCKvRMujyNPTMhQ7826EzlEtXrC2xM+pDZ
Ymy9k7+rZx+cIOzmctLhSTdrE4Eb0urC+LUf6Dw5S2AKK0vC7UMMoFEXCXmQrktrrxifjsPudTA0
1VwkInxmrfGn496Hr+MAfY2FyXKFsu0iYDN+vW3wEdSFe64ZqspEKtLqzrTyA1cQORHhIS1ygj1A
7UQZCBfFzF3pWGW+4fgBC1QObxhVKcCOhtdYtX+hpTZO2dBCbMfnjWxV4voicIB0pMTUcq3cukNi
S/PgVWm4gjCjJ4Q+q9x1ZEcopiFBwipOWZAdsOxU5KUVltrR3vK35gXsfxuIAsaku4EP1uHM6+v0
GLLXDFeBPjY97/gJyQhtsQkeZGuqtAR9yG4N33UNyx+CDKve7+NqxzbNnKRj+y5GtNtVnAHvNT7N
+2DUD6iDQ4HSfxjP7Wc97qPOnlDzPk/ET27wpmkxirfgniVxSKusOV9y5LgLruGtphQsmtBykW0y
7yMLLPuG0xwWr1US1lFe43x2Ju898yq+r+Sngr3YUyVxbSd3Kyu5T6x7WXKBkTEQA3XSeIWZJ9m1
Z1D4/+Ck+ljyOByHhEwQqw6tckZFrVEW0ThDrO52SZrEa49jIZ0uGuC2jBFYrwkjapLQhU2O0leB
qTSnoFUPHZlOcQ0tw90ND2R+UtkmSEUFxA1V0EHeWnT2L7GRt2JGRrrce7Y3/Iy79TReGy7eR3Df
C8w5SdoLUtx6+3FMFeY0wOfh7I7zzvqmh1kSbXjQFmwJ2cFHqkj1tgRRjwwUio42gCF3j9WOjfal
Yp7BlnC1cP16kWLypVsxCMh+mNpisrjIDepjaZNrmUDADxXTQaYfa3sHw/pg/ZEGd101bdY5vkCN
KCxbcXtLsfcRs9Eiv6iVlroCYGNWO9w9Czj1wlvi8ND65eBFeZD6tGQP0k7RMNrqarDAoBn8ROY2
RBBK7wbU1Yznp8Ji72vFw5bFBfqTAP6rD0839ZOpR9JIRCRxvBeVIioUMN0LXKBWMtly6UzEMoDe
kLayd+SMJm05ro/xsEfnl++hq6YswAqlZ9c4LhLR+INH/giP85dHg3Oj5/63uUlLoN0BeZDy3vV/
6VdbQXmlR+TPB9NNpcYmi8Brc46I/C+11LUZtCV5wAhU7tuEFtCEkmUlop2omDXpS6dit7gJRyMK
RN7vCzLSQUiHIihj6hdSPxMno9ztp22sOYwDFDDzl40Z6lENGQGq5/TiwrCtKuZvIAPVHbyMzEIi
agXHF48uVjKWiPrBNZO0BrcysnOrIf5s0ajIl2gJDwdNwhBGpAh1WCTMbadL4Ax8c/xx7ulGmAqm
41cxEp8V9yK8DKdMDjgm5Kh9hn6pniQfSqyQ0fXAkG9cDs2yVcv47/R/XIacugkqCxD/CxbMc4tK
2kEE6Tu9D8rtxozU/FBe2tPdHWp+8d9hNHpAsgn0zeXv+6rSfZ6/gfP971t77F/QrGz73GuUIWf3
5znwEFdf/Oqqb+yOldpn8H1B1fXLFOzix3GpieTDr468pUKmP0GKYwXSh7Dp85nhZ8Wmqr8mW4wR
bR6bEctW2XvuvuoBYkmWm1+TKBEmGqarr8imSKnNrMO+QLlxiSuDMrG6hL6OXsel/bghQo6hJEAW
5K+djVbh5OzojqqCFpfgut91b0LMvRpbpj/hpEqZ/7Ei87l6h2RqM/8C/DS6p8vi+/HHzQ9Pjlwu
nP4gsBj1VfJb8BG1ItVAMa6UsO1G7cl5iPgON+4xWrNo3yfX8sAiB8TdytrxoDb7mgVI8Gu8woXe
VZx0TWC0Conv5YKin2VtSSgNoyzy3YI5Rj8aURKwadq80DinyC4EM5a6552AihnWIjZtdHGKUXWb
VMLrV5HYXhND+4b3FigRv24rpZbtpu+526oQlt7GjwDcB5BWhMzfQu8sNBhJynKEyPLMaM2f0m9e
rmgEig2LHxISUlCZVkAET4ru2Yy8O9+sOtImTB9Zr3OJ2vC0yozJ9D9AVy4tCmBnVC+vuWLs15ZX
NXBiRwXoX72s93MzAVZdtRJBZPFHtWdF0RBwIvGm4EVCsETomipv3m1drpCt5C86nTVJrMCIqYbL
pF1vW/BYVocaPfSoiMalnZ/D8Y2LB5evpI+jCAlUjYvJ+hogmrGn+Fddld9oy3k43X6H4zquSp2Y
K3Maa122gyKEwLAP8V0t8Mbo7kZeXlWuHRRx9GGqnEbt8rgvyZCyLinMVJvx7L3wpcpvxQ+opHKv
rjvXclZKyb23TKBV+B12ICQbRuMbgiPTm7MZJPlOxnFon0ZG/ZOS1GOfKHXalZN2wYuJE4cQTuyu
azfGYfn81Nel+z+RgR1LYD6zcjmPC6vod7f5IeTa84l6WxIO56ppqQkgXu05WLQDeKsFcEE0Noc2
mQTago9V0JigzQvy6X08yDTv8teQZGjZ2uzPlqqlC1s5zfyGvdYJl4K/3XmWQDdWEHvnIPXO7Yj6
1g3uNwY/TXxLDrhHv91ZKmd6YJMnWnwz9vPpuczcezV2zr58JFQPe5jo6KTro+Z1MRW9/GL7QZxA
Np8wINwNJTLVGd7ScTl6rN25vfPlB1rFYp2ihO9PVD7AwYmElFOU9pSjS3UJrrUtxtu3Tjx7gMw4
hbBKOF72dq02EzxrrRr8OF8WNAmSCaARH4N3OpIm4UD12hxCtwAN/OHqXfbMRFTeTJhfFlqyHx9I
EC5U4GxN3yhlcuzK5k44IHdROyRRs50pFhNHrQEldwPIIJ+8x3ZPmAejXuf4qwJxEuEZU4zyfyRU
sRu7dlgAUchsKdEoHKnuLz45yRJgwb8Kq+6MSmApU+yRgK6yZtFsg53bBwxCQZ7UjA6f1krVIEZ0
ejoM1gXSdXKSgowOASmvDPFn4cghZ71Gc0HoyvBY9BDyCbZzu9ffBSgMMOrIlpBESENVR+7c3VC8
hhoguopCplS4w/C9hXNC4z8LIMjxHqQ8daPzMKukXmz3zBckDPRzDNFljM/qTUETSWlTutmfV4/O
uMDLsqKz9JL0pF7LdUpgFsvU50dWNGECBWKKuz8yCONQK5dxCgAKXZTczIvGYZlk4jg+4GhLch/J
fzJ2YSHn1BungCE6T2kmNXEf7DCl3nKepeqnCFehh8AnCcBhc78PW28SzfZzSZoVVpyxBKWBdrtc
6JmS4/fxcA3rnLnk9TVeC/399QN4G0dfdpJISHN717d9RaG39ZxjoTEvtb6EwkH7uunM7O++21YJ
1laY643rqA7j7VEmPdyIf3kJ6AXvg2PA/u9u3N5+VgC0rSk/Y4FrRLdjBKR03kubZ6HM2mGJK9hw
ak/kBQvl2H8tz646yLh46VrcNlvJ8JJ1YJqjFbTBOHdPoyK2Hx7ZzUHZxhNV0nG7AQ3WvAueA4W7
NOH4+nywgv84m9W5m8nvAOuOcgELfafzd4pU8EhkmlrLsS8MoNBxW49NkVspJqcnEXz5zLkoIg9f
NAwR1pMo0ll14rEdDY2K2KCySYrTFsOuVHQgE6HXv1zz7V5DMF+8HxdNHsk+S+6f8XLqtBNh+dKd
EV6GKNvL0ykDtJtu9ZwO6B84gcMggJRwOia1x16dzSfCOhshwz22GUfJg0brxKLJl+LtNi4tE2vH
49I0ukUFlU/xjXhyeg5aTf7UpsD13mCzG94kRbisUJtdFMR7QVQZX0c/6FgyUPqYaKexs8BoskQE
okk45gZ7/sf/6Lo2RfgKcbcJ9RxPG65CxOewyzghdc57JKCR3M6pnS55CVDE/JxBroc2boVa6UKe
hSbtzfWS2ETum/2UdNyzeEOxK33Pfu9dFuzbxKHN75rBjzLUD6cQ9+xaWt433iphzTPuszUsk6oe
ZuIIrC//KZ7W0i/T35gx8gWKCf0wliFcwpgaNzVvkoLhA2qCSDh9SH37grRiOX1zj9WRGFi7l5nx
oRB5n8Q0BWLMTzv0lpCOBMtGkqF77f5mUQ4+PcLMPOWnxA2f8XFLYY3HQIUOoHikdzPBD6N5Sb7d
JM5hs1kl2kInuvZv3ed4M6GJ3o9nxj0X+KH6lB8TkN9xKdmG7UaHi3Kac5Y+lGcvCXDWDoYr1eau
Ecy1i8/+vSeJB9N8GRABc+pPPixijt97hyxzApYJYnEkFLK9EfE07U0OTJil1CQ9s1JCTlCiCbJ1
wJogEcAUXM4I22pfckz7D1dmADOqgfcOrDKfyE2PoRFVeHtXNaPawDYVM8yGgYuT6PuHs0JWKLVz
n6FECH5pFEoU0yCkclOBJUsvg9RO83yAn1ae9KU1uiMSTZbT3w3YjQWJPfpo76JxW/gEXEAXAQIg
8GFL+aXWN/FKG6B48rp5zhZJSaxaByaZ5Y2QW8u4deaHFahx6zdWNFSYZeXP5X9htmL+RJV3z9ZN
/lQcHjNmn7va+POuxFjZxsoeAlsCFXLzjs54glwrU6l2Lc9C1jmBkWdE9cVxZrLy1J1srxkzjdmD
TdKzUyJg7lp6Qg5vDhl8lEOLyP44Yatl+IVBoABzYIaWWejeYcUHpIe6XPfxQK326V2VyocFex5Y
S9zNPilS6i9Qo3snJ8wFpdmcimvOZwn3s+J0Xve0ROQ5sEE2FYnZn7fFblHhDjsgEvm8KnXFjmo8
ylCLTm3KNwvGQyJ4B2gH4XjT9ar6Z9bsyXaM+eEPCeNtoj6a5GBnCzph/WzWphDcA4vPzhSVKj4G
PHAKroMVGj9FftMUFlIAaoN7NG6StVexemu0DpTrW8ePKTwhzABwxsS/zRB4yN0GJvAPpYwNSNcR
2PZwU98k6ablnK03RdlV3XFqK6AkCAH6lb3XZZtB9rqFdXV/cyeqJAzcMe9fcUqLem1pkRtd3GV/
32YCOArzXT0IrD/1eiR7VRxIYCkqlsXxJpZTkdrdJDYGM7tQRvfpKR8CfXSVmlE3SeABK+ShcFDV
QT7oE7ziC6D4Ykc8e1OP+vJUc0VJoIVl70lsADpMNT1OaZx+wz4dthT0wMmeM/2LOfJ+d9t7z/dY
75jRwIfUdghjkSbhjKLhYi2rEy6L6AuzE5tPedhvjTLpnlcsnq5UCVqNPBlHcxqBYHaks/s4Z2zo
wFuGCU3ePmS112ULMlmwZKM8jkIQiwKGQXqQiM4j0xkiepiLt1u7Dn1TZ+yKskPUoMSJWmgUaKgA
cxFhrAfVBN0KPtHsn3/UoVLhriespKWMMLhbfogLNHxlgXpTa10ECXlQf+tLzeD7jyBV5I1Mz0Ie
H9YPxcKdwhFI+5DuIeSHH3qZuFzYH0W2Z3ZfetJPz7iWXMpTtRKEFiY07sXpiDeH1Fa/EoIScyA6
OzlARjolD7PjjSOSHXwEEcCzRvx1+q5CbngLrLT4Dcrh13sIv8konusP4VNcAEFGLOYGuNRDzTUe
ylKUwY8ck4hM03nBsWs6jhTlzMFcwoVu/0rQuouLd0Hte/mUT0xEbl7ADKAfVO1bFqgYlkXc4rws
g7o9f2DhgOX8f5S0HQ9h/eqG/Z0uJca+0UJijscXPe6fv3Chnw1l5Vj6J5u9gs4Xd0fbDxoSs7ub
6u9LNZKKyOXq3FZtMOPMd9l4BIj+U05d8hqyJX3PhnCfxaWospnXOifrBu52UmsxSG71vHwSXH7k
+3hy0puoKsEDs34OHM+RdzUc4KjWsRCiWJKKFUpncU37gyRV1NHxujlR0aHeJUXIU4rdcAccYPvN
G2xmcDb6zV4QOHuIVFDVDYomb5ogvwtHUM51egwUqhqQXKseKOd8oQx4dO3jFMEzkrfzhq8hK8Qv
lTqL+WH8e9V53y4EP8Z9bUilAB4aM1KdKUPTeD9LNmmV8zD7StjSDgqcRwRx8gyP/KITjC2tdSmo
aY1p5B9Jui0D3XshCy/MkxicaTkraFZ/pTP7LWfNAu/kcFCx92mV5UdCo4WQE/LFaALXY2TtKR8g
vVWTv02AiLU0KDVYXAA0aTJFE1+fFshVI8aGW7A15puezCyavM+UVrBJfcDc1D8aBGNstQboDQkX
PmGNp+Jnndn3MKG/+1ZYo1iPpOGxAFm6lZ74CUGO73JpkLpoPDxikpbat8iZccuYjOWCqqX3Df6w
oDj9Orhd6V/lqVRzclqit3mUyluBWiHZ0q4ZdsDGzWiHm4jIWJ/zNMaDoASgJ+mq16icWEDYK/ys
eWpk4XRHCeIzgrltMObEgrkyuuA8MKDl/D8vuVrQNH5CA4eX1fnR0/ZAgqYinEJWftSWanHAPD0M
/Zh880klGoAausQyeuHBKuza77+CngQ3eVmmrr9/YiO6QeGEYjpJvadsU3RLpoIuIE7NFF48IG0q
j3Zm6cmgV503tG/Nc3uOS42258ocf3ZVRunnC7ujEor2KB8/OjZERQbkfR0KWl3A77uIojpS8Iaj
U66wCOPJjRp7EJ9iZwLeOGz37if3S0ZBrxgROZCt3NRdemAgJhb4AYcOnYsYpgJrE1sc4t+n6mj7
QU2IwG40lKyDJHZc3IDXXx3HRPb31s1PT1J0nJcL2blcpApEXJIDpF7eu7X6WApLRtSa097WVL3l
zSsAC/uGjw+5eY8SXmSYcCEvxWz4q8g2+uMOG4rDaX4YYbT9eGy9uyWZfeXxNRheK5tpL+pvmjXL
Vo6eHW9WFS4TD5THhXjWpnxqtXZ6gOsChiFyz51VQpwz4hj1S4wjMyK37FMl7n8FBDOjHR+YS8Iu
/vCdvsx1vsxF7UJ30t+y8RUo3Kym9mRoOkc482uOui1RVGioiTejpmPvw412y4rWlVSDZ4xh2ehB
HPnX4pnE5+E+1SD7jneV2ikfgSUkYlTZpXEuX4bzyyP1LvQehDJTWD9hoDVm1G+7myjlzURXHErd
t6T8QVzHECAbXrtDuSdSbd9hJOhvjElzjPTBBYVIkYqdxugROEbByTNkVdhW3zW4tmB62bJ4ECeE
SKDgPlRUOclHEKVK9+A4ywJLslK9jsUT+NZOu+nBs/7LykppeSxQnLxlfH+IBVDq/d3UyHktYZ+e
DuqatKX2zvFkDhriLC73WtVn2ObS1n5UG0zU/mXJtxkXy/BoqC4X0JgsZeufR+hhlOZ0DEevE55s
18dJ6Tl3QxpI+Dw7fvhq0K4/FntR/mJY+lEOA6rJFNGMOsIKYnc0co/kb8zfHDOG3nlufpt6uys6
Gb4N2+V9q2BKr6SFfe/fqtcL3NHCy4nWkQt72m3iOzyEfHAsG63zeUm0gvt5hn6mjlgUqSGazfAH
Cg4jc5o4HZ201Do8g9J6AARX+I2z99bwfIQb5IYaZi6Wiyx+C36LWuBuUMs5LuMWQWEbg/xSIN58
anUrbgZf15MHD3NZWKRMFMZkPqV/+TAk6RPszmKXEhpuL7mx7t/nyFrZ5iqQux3TPDavPP8ze/bN
/IgnINalfuHaCkXO1BLMR0Xmzh92Z1tgwrjeE8kT0qIWM9DmWoGbK2q3zpwIhfTL+Xj8W/hNySTX
sNKWnXZiXbPtRQjppS/aqb92nxW5axb5HdZYkolyV0t0yCp9SJKNpbBY8UB31SvQ44PenqMNijZ5
7ejS4SWjXFr+2rBRQgJ1oIlsgeX3llSSbVErEpJtjKghSbGuDtTbwfeVECVKqUpP8e5KC0EDmkEM
jkoPvQhkeVdUT6tprNeKZ9ykkJ2fxiqnxbMZFqR0bxiO3yTzpNrmYc6pVu2tnctl4O2F0qFDRGWw
kb0nVrOO6KMYFYHLEabk2GCItwCSGxQJQ4EzDFmf/PAZ1qqy0wt8wAp6UB9h8a5z0Nf7LJ3q6PNZ
BaIHS4t/uIv+9BeCuTUuyOH490c0PABDQIBEfVAIcVFJv97c+hMXH7KEphdHfJEnnYplqOUoc1ET
zSCHtMbseLqrEQgk4/fIW4jMxhZUnxX6GtepAe26q+pFWM+PpSa7nQmTe8mpeMBfgvJCZdw+n2xJ
+lSlGViR9/d5aQD1plLsSZZnGzp+sxV/GQPecYMEbTVjqaK5ybiBY87ALijPbGAz5A5x9pb9eRMV
3KIlZpSzjXhQy8AUOB0lzXBuvh6sxTiq7gQoG+mS7MK5ZDc1jkJK98dajqatj3FjpBUfHov6JDZY
ucS+pe83cEjodUlGPfKGNPCLgiZs+up+1zDPP9cLC6AoK5nMXWNvFp3vQdtlbbScta856i4nw+Rh
AOi9PddptVUd+4pIsXkrYPaSeDD9WKZLYPBXjy77gyQkUeW1irMnnzNO2j5ZxQpQsrA/WRgzsq5h
x7wBYb3UJcoggrPA4j5n9fyhvPBlRwY4XoNUhTs9N2g9hmY+geP220pOei0BPN3fjA4R6rWbkA6e
AUR9t/PGRUzpCYYhgjaER4R698q5MtImdYBMTZ/XWJyCalgxXmwpAgIDT7wtD7Tz3cGR6NDPV07a
QERQO/7buhZ9CPq0fm9xyzG4GPRsdpA0s+E4vgQO/29+CrjvGYIKWqJHuUo6W9V4MB2ukco2JDwx
ltxxFyZ/IFztKcUSb45CpZLvJafCHRd2PzvrQXH607xrrHp/hr+eLGDus+GKJdnccNW+7NITmLtA
cUi3UF32kA+SW4GFpyvFLuxZL/UwCPpfrz8Eh3U/rIOpzZ76qNoipOVt9FwrWtmkC35sxgMkfHCn
aNBkj4rkM3tBw9EHds0dXV6M6xMzHJGxymQM+bmzu4xe60ExxRWtsCKrV8v1LCWD7Sz9Vz1x8hqt
tn4ieknRyFLA45keUwUWH3jv0UQ36eYuXBB16WhcW6g7M1Fow1+u+dZDlP7HPJmZu9ARrEGOsMJv
sujBcwCPQe+IrDo7YAbSDt1mRa/Mbn8qT3ozpINbOtx8U76SyrOf9nhyeOFaOlLez2s4CI0iQctc
9/nb/o5iTqZ6kHKFuPcOQALrwPwFgMDwQ+zK1UgJiLlGks5Y+pJXm0PpLbUSQB5hDzLjIDs3cDDu
24gafJl+cDpjibxC37iFFJrD+LPmbeTz1X5xzdONCRxlGE+sUMZEu2Gi8Ui1oD4ubnCQTICHT6uv
GaPZbZ+3Fi7d0roWHY4OYbFHJHX2APgD1qewIqVTKQLk2wiuoZcppGLq7qzpysNKGXR+Fvo0qC78
6yffkBGY/yW1ziy+q4tGm7q6QctMQo2B9+gOychROVPkV3DIJZXoGvhJGtyYbP9xUPLOxcdBfmaK
Gw2HHQxkbVh+FF7AbP0JqLm0DE8XLUDupWoIk3z7UjFCHukvZu3rahrs6zGUc9SHCD/WI1cjy1mg
a3zivpm2xWl6DhD1G7O59l3H4ff9RYhlRleLGrjlC1GiFGCNA3KUFml8Pfaumf07s8E0iDR8NVKd
8uQmI4psjbgLrA7+hGmtxQA1fyc+ht8so+LIxfifMqq/D7X/D+krq2wZIVObVBomnnlZojLRWmCc
j8tstHazfOSIcCcbyVbXWQOuU4ezUuhb8PBraSeoRFqwX9fTeuAaggNO9xeX6RYuNyfhBMurDMG8
GeIn3W+30PR3+/6NQFi1J7RgNzITLA6ZLVHcepMd7bovLHakFv4LpmFVL+mOKTVtagPHX1gChdxt
5hVvZNHnngQzmX+vv5CtJNBWD3joRAhvvj/4Ovy2C1WXF7HDBswTH84nUKktpbrxPYVK7OwkYj4C
rokFpHRQNXD992DLIjT+YbkGE6iNqSBXKRTyJzVnhreVlazQk2uS+kwv0iY53gn3LDVNTTXZCM/o
owXnskkT5lmyPC4829yFfA3QX0iilUL0fOmjLzaz3RsQGDMhVqzprvXR4bSg9A2y99yu4ZN7EIAp
cYKQG6NNxaPfPWSuaDijnounn+MsK3JWrxYygUovrA+sZrtX3WUlA34HJcMNKMKZpWsxNGqy7o34
vrvhKbgiJns2ZNORHJKGR1VMTYN/xtxMsPXXvzZtFoXtxtVrOD3hoKQ399pxc4Cw3PyuJDs+4lFR
/6SFK6kWzrG/FGLBgLNEwvNwg5EZdhfcj1aHFlosHaogRgCBLTEH6aegW+bXnUsEORer2XEyGSOd
97sinao/RX4BqIt53yd6fcxeSpso+vhsIRNEingcwD1ox/bTKeL0fpSJm6F4XIksYklcG+foPa8C
dnQc9tFnW1rmKD1Myf+8n9Bg/QPlxJBbmtZeVIDAQ4l73prkrPntHVzu8G6Rv4bb4QOvnK3qfpdp
+EKoRIyDEre4h/Ki/wIDyJ+femIC98hcbewmAoM+hxexxofaqlqnuydqxdtYgZQNDGoyIGTKkCT4
V7vM/4b59nKzX+nCYu8XTkStiv7FMQxiBKTYToBovuzK66wkbz+VT08cFjWIrLRuRJrQ75TKOb/a
05OAoZ+NDQrBLNw5JFbcCjWwLkVr6nxNStU3zWwfV9CDE6jOH2hEQAX+VXKgXlmo9/Bl+JfmOVOP
yeX5Y3aR38hwKaV+AWHGxCRIr0OXAzM9WpDXj8aKhtGBPKX3h3lVofe1XM19o+mlgmaqIMn1P8pT
shvDBgHVsGSBgTioujYJe9x0Wp7eWMOg+vBaXmFJ13nYLvMvD0ndwjF2UnPuNz/J43GZ8MJ4uflS
AZPiSHnvztaIlaTJ7QBDHCHlEpFLksQsu+EA3wc2yqy2lljQHuSrriI4mgRI/+GDLq2mJp0i2thB
U6sojE4zuO3Bwlvk8mLNlhEKqIwaSHTgvqR1SVFrU8xv1CDRECqfItfZaI2rGDjXcAvWL2FyHfwZ
OUUBd0ONPRNiZ+VDdQ9tw04W2KOjPbP6MR1Kx07u46D5U7zC/0kbjOq9GiJm9bkSTk36vB95+b/U
ViIw/cVc32nak2uhWjK7OokMDJwHm75eDr7xXuA2IVuA5bjvmejbLppMJKQ/GXI2nWTPxSwhh2+v
P8wcwNkTeQNCOMjZ0P/kZCUyblXjMBisePIp8/wQkHWudDMgKmkrZaMnJG4RhQsq9bjEM35vrLPk
WyTNptgi3qLE6sY1WwqddxS89rSYy7Fkxw07Ytl1vIKOzUdmfJ+kRJuu1htv/CBMl3IknixE/uMM
fiiZ3VSQBd1AC2IBuHI4nzXXdU/Wr6RzRTs+ALdWKA+xMuh3BzZF7fhqoHPEodg3MNLnFDYL9VBu
kLSkQxGDP+fLlKaDwHKiL4HPnUrELXxVOhN4/nYxLY5dmwk0TpHpO1746W0h2z2y50eQct3HjrPN
60SskCu0RRDiUNxYkOhSNYZkzMvuaKzfAKeWUZTBMNFr9jpKD8wqZWdJDyHwnP74YcewN6C4Gs9d
JWOaAfO1b6tBI70ANgFTQq1vg9mcIv9yTgtMk9yZtHlmU1W4lmdpXrwdzlKMA8HuoqVLqfy8t9B2
rA4C3oQWdHP6OkgCWw2GEqCFht+sJQuq/RZtMKPbWecLqGRQIa1Dwl64qIT7FPySEgoVnCKeeS1S
B9cdmiLPrB02pfShuIvF3KZiorM9X5/lerDGk0bg/nEvlYKDnyIShlFGkH1QOJufJB8SqJox/i1I
wY+VOnyczJVs3tSCvntr7908jkCNUX0VJ2nXHg0OEPupyRFR7T7UZgsN+k42WmF1mHKgEPZR33A9
VxwRJgCR726YNjCfLZRvHL1vy4NXPDPJkJW34khNBBnO+N6XszjEkTA3XKD58ckPK2plLh9C69nF
LicmGF/CaV9x+RcSllIxpr6RmUKVWoa1W2QDIOiOC5G9bVHEaHw6XRdB5RLmRxKOf9dUGq+H762Q
hzD0vXOFR3YwwBwchQ9clxtlDHgLjTplPnilL7DiAvVe8jT6EvWF6Lgh6YgECS425Kif/2BKyFJ8
rRnjcZS+wr2qo0Oifm7X8CDMew2cVpCWAc1MGGBWMvs9FQZGMROjdeHhd5XojKGVj5QHSwNYJ2RD
y7t2jOZq6fLMB45dkSd3KGivbPefd0VLHjNeG+Kn3FJ0Va1WPQAk+u9FtCmRqggLYBxtdepPrlg+
pehz1QZy7Y720OBhk8GYVR/wk17C4jssoJJ5H0h6cjkkLMdatlJdYv9rAIKknlCaQx+NC7Z0t+3c
Pcr1wWrE+8JGgUPyaxtz1Cxp1I2Cogf6nI5CKPdaVSz2wHeIb7CSq7RKqkFlrnPtsUtpq6bCtFGa
O/F32GdKQH6yIHb0TZXh01WLY4Q7YnZCeAWUoo4Hgc1sJ7TXPwjcVCpedCCTaAZ6mOHt2OT7aMSr
XlLShf27QCmnHP3Du0+Pmxi5ADWIyBHpjbX7Jx6UvVBNicyEfsHc0RPyBqeHe0f69NRAS7Ud01li
ErH7t0bTLad1gh27Fsh1FkHRYmoV78YK+Hk7YMWKX7g4d1lZ+5v/cpr/pWuZYDzQEE7Tw0KMy1L2
LXSgfHpr1sHeOwxIZh9wvDT9QX9M8v3r8uMSdnAZAk5wHT9FU0uSkYjAvgF63/tuU4wjdgeQBs5l
qrQifLL2t+U3DMpWIIVF2L8eXtaTwCLm9nufoX+7GESJp/4vycIrrMsycDxOFCgmj3SMyy6WJBy9
Y9y44yn6tptntMcfWt8TratRvnXTecd3kCZyfIQ1gcnCy3O8djCKYdxsfX9KJ/nX0DoG6Ifzjd4z
mxpaUPR0HF9S/TSfY5fUjzTOxrvFFbttuXRN0M5TGiMScUZ4kG7f2Yy+kHf+FTA2m6VUSLnBgnB9
2relK6pJY0MrTnErThwqucVvxEFlfnBYhsW+5JVa2Pt6Es80IkjUzAeQOs0Qw/eTqbAQ0JNHtBJL
h07MfyuEZj8JVYRAlQP/yqqjpi41ThQrxytg9znHu1bTe9UQ8ZoMZulyvJ90O9aWLZFq0cAfDQvG
fRRFqdjmAmmgfapGGwDFdkHHNVyzZdd+ZWXe3pGrvP/hXOE7j8EuloaETKYqKEznyT/X4VgEu6zq
JCX/pb0wHZCc5h35XBGpMMhmjJjci29iUc8jfiSrsnm3UomX3X6WXO7M28CyrZOCMk3x7vR/yJHi
RJ9Hy9Iu8BLkJBqGooEA7yf9rOyLqblEE02GyMxf+TbV7B/nIre72GATZ/9314VXcGoPnF62F5jW
hFXmQCafGSj5HRAAXrCPQhP1CTpY5gE9MjPqghLSC4uQHRSuovKqz5LScPU/tneiIZm14VyR5k7o
aqiyVHo9oIetw65595bAWCFCpGY6NdfT0IyxUmzSmvPzNK/gT5AHFx3WYt4U1CNA3xHUxd4ZbNcg
JFkuQnvrDUPkuonjPYEjqUTrKX6qjpSuVlImlDFmDR+xCgNb3rh5oZyO3r9IHT6O+U9xEO0KHqNc
7TsaVAMMKGTJtxQVI7+LjWGPcgcZRv3TBLQMaev6ni30Ht6POghmU/3s15UVSuNOJqTVWPMSRAoA
JT6dQp3e8OhYzPmg4gWP5sQHAFR5Z2RD05MbTgfCdLMFf3jZi0RPbutbaTDx3SAzNifAGu15AtZ+
Kr8cWy5U27yPjOHLnnM/4CJ+cCyunqEhJhcNEw21g4rtWJA14HW0+Y7h6pxOmvhMdWr4w6lDCICo
5/Fvqx6OXlrjeIiwMEUFM35PO/ENHr/AM0zDlqxgcl0ITPRjHuFn3XwjfE2Z0Ku14G0/ybhNBKPD
5mYxWO2OjwP2JjiRgRL4vz2KaC+EWOmvzjqjKo89rSpVmSJE57TRsDZYzA6W65cyibusPIODHq93
A73BnOTsoZP42mRITA7PzRao1FMHMU01kUnMCE4CKaVdjgQZrptB62BtOzbyvXcktM6/kz+aqIuQ
d95Ly/3yolhe24TfGq9dDSFNZFLSjV+B3cOZ2nJwT23dMS4dPNIT1kHoUNdb5vx9GRmvgNzRrFWH
HhEAe+8E/57u/pBc5H37330k4T6WCIQs6Mrl9H6TALATMggfIlJUquXWGUVffFSukQp1c+M1NBlH
4BORz/AMk/81O2/9LCqXVgFZ9J8WvjJMGxPIPT0arbqAjnycVjGncZIytq63klAuSUphtQSjP5Do
CwIIpzn05knsSEQW/hevmFIqClUwQbt5XoBG/WDINAjCz7YtumlSeGe6ZxREXA8PvmmfoDdXJEGL
4Dr5Uhg2/UQhnt3RwXSe16ssCbS0CgPq0DbMxI0jtNuLX7asV46dLDVkWcfYElIoCHY/I1bfsaIz
JljjBoihln9k960IGkuaY4LggzYYdFmKptZdngz3z2pwS3+6qKWoxOtGWaygDv+QExNvtEYVc1xD
cgsT/wVIJDzjNMzkLU80tcNg93rSAWq/OqUhXa+w+K2Wpebx/Rld82y5mmXn+NY0jl45TApmzoSJ
AwteEDDT4jSyBFQ6UrR+yustpDEpFD44o2plnqSEOnNn3OTMLuQf/QyDkidPgyYw2JfiK/LNI3R8
QgajOT2WdmU+UOkrpJeTb0U2alCSp8kSGTmhW6Pmz5um4xvJh8GaorBYqoJ5bxVro0X1oj9C3vlP
qWv3LNRxwNg5idXbjIO6QbPufWeBtHmH5W0FrPeYzN9g1UZcWSk4wL2xtVikkbyoxbZkkclEcnYx
1kyaUsDC6ty/2O8Ao+MT13x/1aRav98TjZLgqMw3NU3A9Z6U4sBcd67zdAj6VZFtwX76JRivVXlK
dP7lYQuFdJQJ/FG4FvnaAWVtQEQ4fhU97HEqK1n4RmYNKsY9upT2hKnoto6KVkMzgCgWvTOngxzq
uN6JGKA6Ud67qNmFEzclRs9/JPvEKxOvz2g27OXiVvLi9/HWIQK5d5JfbhTtrbNwc7EWheSthXRd
752/JQ+PfM+uz7JpZvpCPiuTcnKhiKgBOljjwLm7ZKc1hbZAxZ4cEAvLnPN3WNjR0Y8RxiKMXBIW
Y88Eeu8K/YvFrC5WKhs7AVX0C/wD3OeypYzJe9mPkirVWPoMaYkUS0sM4XAKNVrIRdwDo/LYW5BB
ZVV1ko900GEnv+49ZcDPT95I+J/pqitSdDo8xcOUedIF8BSW2Xge5kUj7vssEOJCnfoc1ROOg3Rb
BPYOrsqwJhYbsdbLSvZH8EcVWLT+JVNqlumL1Y+zpdr61/adRRSkYIfepMzC6IEc2V0JTK6XLd5h
Ni4AlluMT4cC0j+N72vQ43nAkTH6TCDvCuPg9zUHWzPCntrq08miaSmbou23jbabVqJ0H8dd6JT5
3R+9IZRxpamqvxj3UsK24k5ZYLFiRmjF9UxEQXBjmlSpWJMmlXj+SpMpoMNwqOSe4slLi+bWLBNa
HrZvFuP7aWi4P2H9DskMY3Otq2QUoi9S5L/UqjHYRu8mbJyP5qPVUJoWjWuP/cE94CarH9FgjMJi
S3eCMc/QtJFAHtFRVN82feSgh40sQd8Aq78YxfLQvxCL5ohJHxhbg5yMGrL+k7N+AnozwQNaUpe8
6KKwsKberoCivYFVZHui/f4B/ywk+KL4zJFeSxlyttyy5vvy8Hw/X5tBOaPDWBBMy7MflZ1G7V9b
lH6c3q9HOY8IyC+FBErcfdWRhcYkqS2Q4ue9xTQHKuz/jl3a5PrzZ7yPEIaSuI9vRa/OGEnzCxfD
zvSv85fNEbrCEKPdAwvZjosmWMhw4ROL7w5w+y0miEIFWDaJmOiaxlcJnl++p+CfqQgOO54Qu8U3
uwnjtjln5Kj+AoZLJ9xzN1YP3xVNyC0k+7NCeW1KBREYOY8yoJtqz/KI05Jhz+eTBnqv8lQw3iXT
gXqvH3VXBIsa88TRmSbBbeDeAG8CeAEx+Cz57DVHzctGsOoeruG9cw6gT3cysth/9DWhfk3GU0lc
0fnRy1uAFEFdHDuw2ciflgMylcQHn9G7v95E5D+qfiHeWqNU2O+qegK7kZxS6eAoWsU8mCsLdmd2
iURjKqf7fYQXOhcchRUaiNqkPByZmaEwWyDf6dDk0QR1liiT1zoNqkle+ISfD5/GMAkXBg9+EOa/
TwOHyCffMRk++tSnY2h5dpquE5Q+o8NhGMT67eYchVGxZXk53ac1HqW7pUl5T25TkTHP0PBRs1cV
J3xwz+IQGYr4701YK4AhskzTmXsdpdpm7pTZFSrMc5/TqUWA3rmLH+O6ci0rP2oVUIJa99PQybay
CCFuHO5qisuclWR5ggn+c4R9Zv6Mdn0u+a451MXjTduQTzCUJfLbx+8duu/UnAU1MzkVzJip0bv7
1FAW1vcLF5ftQzfqFbI+LqNFWS+KECeCYY8W23krs/Sb5raoz0vj6bf8ejUe6D7H/IztRa/CWUMF
n61MgcDhF9mOe/Sj4ASIqzmPqxMDKMKjdT/7jsZvFrGBZVoHUmbD+dWJIizdg2QjfwDNoQYTO0up
o1L6rFnfzon8zAtFi0GyBPaOQrIUVH6jQJs3ZoqCq+zZ7EyrhxRFYRsJf04TbJ/xVsnBfPqgDLWl
mJiCdhLmGyqlUIdQvCtcIuaFuBe5+he6ImHuRvqijFBadPKQRvBpC0TmL7W4fqOMW1fCdbCxZfOS
wuE1OS5Ua5jWwk5PT9XTv/DVv2Cm8YnpKdc7M3dECG80jZ5DpmHHqBbZqYyZ2/UjFVaYH+QoH7b+
yF8XkqXtqu5IBopZAEVR66BlLBN4LCiLNJ8zu7MqSMEK86UPV1KjFrTb33NMyWk9lBTcCZiUFoju
IloXHPTX0VIyx5zyZpkus78C8Jnb8HmBD1Y95CAEpSkfUxlGLY3LynJGp1zd819C40n/38dJ0ruF
OffapEY0podHa0OVbEiK9lqj+F/wp8TKLxH8jeXyO7IAHoIRK42c/+FzpLfJ2AmkOXQhz8GfOCty
MC7jYk112aojkNfvNTChfhuoFkfPtUL55hUveXr8OXrPuF7MWT8NPnq1IDVpoWyhcrR55Mypau4x
xWMJS66FRl5DS2IVwA5aYboXLPHTtS8GjySnYmmq8C6Wp4YcjDjWlBi3IeOfooG+vSQh4Ex8izuF
Smtc/P5EGq2KaRUePP4TNsowiJSsiKXB+l5YN+budmX1T/7cOqk8GspdauPSb5vqiZuClUGapTiC
XYrSDwZt5ayjPnGjB7qBAxIL3BSQWrnlV9uLxc0Qj0+PhaszfpZCu4brCRNrX1T2ZltT/C/48OSO
gkQUYynqFvHQIwyQGa1PqDc0yHmSDXQ0ttb4/UWzqro8kmcR0J9NMEDx/bWsULDn9WmNY1H+HibN
uqYUqY70FaJ1wE/6uBMYGMJaAhHg0G6BX91Zprt02KIBGn9IZs/z6Jo1HI6AwMyp8VVIXfjNHLzQ
QoAyFoZU37joSrTVBrgIypsgfhNqrKKWmonWFR5Or99UPkma4AD3YqPGVPswDfIcAjMu5F01nhx2
AGPahlhMi+JKP7fNhISS+DAyMNTyf7jAGiR5TNAYrFnMh0VzXUijrz+bGRehyMsru+HBYGblT6zC
AVLmfb7eAxS9iX9mIZjfMNUIYJrzeHAj5KDHUEvIFaBTZSmIOXe/eqDZIit46o4QQ/sN6Vvn+vbt
kDKVepnVofu9rzqVdLNTFJofOqXdkD49azaC9nyxL//yjONqlySYGDx36KCGiGRBRyzRoIVkvJpG
U6WtEm2OUsE/VWzZVdoZn6JgMc7kB4h5rDc0BjoMPdjorBa/+z0iTDOFdKms1FOmzF09nmyytEzC
CuPRRtI+qCsKWflurAPwG3INcIUmKBtwjDU5Xcn+7f4yxd5KPM7NAwoX0ylCjby2u7DKJ6r6y4iF
9k9hqMosHG9yInnYfszsEx5Cx7nZOJpCG2biXhDj5169CDdwWjrK3ZtSPsp0rfF+xwzgcmsPcoCU
ZLfAwUagPSmmFNGcU2QHeEaVECuoN6PA2nFqpBCgDWAoJ/ZRBvUZYpBT/0BIndhxbymLDyklAN/E
rHrVHjnZ2oF5Nbad9QccDO3m3viPxyJBz5emvvbTgHANYQsBvsR3z8KBS9UyMfP4ItweDya+nW8Z
IqnScfElRC8n3SoVATN/8gRnoeePhUi1VkwyvRf0B7qEFzemjA43kjKKXzlY+oQlF7F9yIXq2Zqu
BGm1HpJgwA5AukIbW280mkr+lrim2wYDISxuGyhNKEOM6mOAHfj7IG/MnedrWJWJnHABy2yTiPap
z0D1SC46o3GXyyQ/cNhlpo3zv1AEuEOtDbz6sV5PYkxjVjzbPTMXjZPnb576tfnSdOl4n43RFitz
hMxsx67H9l04JPEG93GLddT9ngUT+RpgfJ1JqeIK0/B99GSFkbQ5ldVa1sR5NQ0+SjBQYzods/Tu
/Araji+SdHUO91zJ5X5NXF204aY/RuIoRbJo9lEv97m55WPKkTAgH4PmpL4CGRvfFeNq6Pwd54LS
WcEeafiTu2DGW2DEpccu+VN1ocfZAwdZ5oCihq7UAhCnBilZAqCNrzJ3w7Fv9fB79MQeksxgWJsO
6ywSIqUHd9rpHUrIxaKUkSOL2l+ED9aOB5CASiZpIil+T8O7iPMJcotIJcwdjrEUcAiNRKj53ejO
3l9h0yWoMBXGxAEKM497Bp3x9hAqVD7MsVINpVzoWA156AMdZDUWpV1sA55/owmwSNQV/dgEBZwc
YAsxQvzrUroTQOgIPw4QPd+HSsO2GYkx6sKz92YMaPt81/ONngVueNSbFV6QBFEFkk3wz/+mJpjL
GNaf2jA9R/IHMbdwCtosdtSUhq6fTH0FEg/KsEg3FBFW9lCiy2tswHuCum1HTUx8qtguOFoKYGGn
ZOkWvhelLMhP+jUL1syRuQxvYWhSOgJR3ezCqAQMcmG/4DZRLzGBqbjD4+oVKXBDdQ33fmGcJKnw
WyhN5Iup0yUrlIMVBFuMfhYVygxsnocALscxyH8iJP5c3hEbg3a5bYwjDU5F/Y4JiB66mCg/OqeX
/olMr/1FXQy0SOSQu6oxXiMV0mUf9VlyYQRrp1ryhskNAHBfPvDlToAxmN7uODAChrY2BjLas59e
EuLEQMNGnYqqqRcmIGt3QM585chObKNuiO4ZyKL+RA7S0w5NDSLsdupqFcWypjpiQXlN5A14UMEN
k05Hk4p5Kc8EfMBqsV/7b67kJl1fqRLwSm3xacG0gv7cnEwjDqbPnOcPT43RFgXgDUHbGn2zbszx
75WPNj/d9GY1WeXv0XHJTVNR3b9aD8X80uPQgrdsJA9Vi8662+7mZ7rcCC4Z0b8cyCtAiXYsP+Cq
SKT68KZ6GQssEuKxt+VXVblNCgqPmnuxkWzpq1N1eF+gcJHJ7ZzwksfIVLc7kkpg6rfxosfYjRUc
Rs0DFoh6Ghk8/25nM/OpICQrAPfNm607GAFAHJFJk3kRPm9x+ZDV26Acy4uueMSj0D07fsdV9QF4
nWcfck4Vh5k+ekZDVCCuTASf3n72jNyq985EO4GaZ3ub5PYEaVU1fWF7NY/cA02Q1X0PiyRs96Mu
E8Qp5LBCEKrznyqDI+szGjH5TrFsbXj7PdWkGNxuAlbMwrFTeGhyHBUfcOEZIkxsR6dDgL+hdyGA
g6SIiM0lJO5fBtA0FW+F9ggZvfypwTj/XsvvhDmtrmeAVqT4pfmftLVD+1RMGZOHsXB3xvPyZXIm
vNwSREin0MV4QVsfnxQ+tImOzd+2KTAVQqgbIIaly47LeeHT27aiyXVIy3TaovdBn55DsRaetDcy
mP0sBuHuqvXogQTAWBbA8tqZvHh0zK8BhXf5vCCbNmFu3F9tYcib6/MshUO6sJJbvZoGN7q6GZVf
TUYZmE88GF4XG+uL5z7WhbwDRRP9gsGdq6FECVtV0sxcuW0pE2Ib4hAxCmmRMamzxgQgt75dtkSm
cqREZrLmyo5ayMyffrZtbPxnGzaQSo3i6CYpFUqbeA0DqxBMXDa4+VLo4EO3yrV1f8erLLLi8jW2
+TjBkF8bDjir4RGVpbFIB3g6c7cicMdbS0ugtJpNsux/DW6rA08PrFkSORmlPC/JfK123peWFNA5
g0B0De45aX2Djmj2cRFHnS8ZMTv+ppbljIqDWEwsBkU4Udz2YysDifAc352O7NrR8cOj5TEY7Ktd
oiBnwv0PlrnZSjF/Mf8QwpOLwIAanaOzQYIsUEY3+7TrBp7krvrfXawsrlpTMir0lIV8QD9cF8wt
yS04Q+V+uMKoqB+QVm5SvXJuUFxMnPD3wiFjoW0l4w3OZYAjdAvYG6kBWlYWh3ugHfHK0DsApnyU
MyL6+EOee+oKgm/egI50vlsudb1cxZ2Q2DPnt+VB0cXA7JfT3+1QCI4ODV5nn7CPhO6PDxVYdV8M
TJCA2IqDIEoLGBZyxAUPA7Wsd6n+Zd5uuE/2kvWkNHzBJXcSPYn6Fsg54B5iHGag/Sni7R7XpryF
ZsJihW3kRga9e03x1A6Qv7wg00RlfWuuh60b01428sbzFy3KnGOqc1RfZuCaJX4qdQGSnn6S7VIE
76H0mXZjG+SU/NlVn2DkJo0DrD9SnrC5wcGBbnHJrlix+jJZZZ8pmpuEk8CsXIG1CeJogDE8sR4D
a+xYI8qarXGrPJDNpdmmz0+mz9cE57y5ZDT9A430TRUdE1+4m8FAYd9fHz+q2X8E++PVxTEN0tgm
yeBU7Mm7lY2eNd+0KUl2Xz7twD/jBEQmz0m0+IPnFbyt1o+pNBARHUTLzrYYCYHF8SvaPGW+PIwj
UyuZJ+l7hSSGEzOPTlXEPC794A8CP1a8aXoWUA3Dnc/RRDkifbu8DVC+J9ihqMfV6NIb9rg28N1f
gg7cB/QdUkBxB7CAGA9xEYXipHLNgteOGQTcmsf0dgr6weazdoRg2Voos8zJwyWYRrxZhTqppBa7
XNub6b3Wr6bRY7ugfYHSC4xJkHRVb/75eiXopsjj6Jp7Ki3pyFWgG4Bnte7RnIrvKrObU2sMiUqY
UHJllwdlAaxT7bz5XMbg58A9ZQnuW0NEJugF63LSjBzydWMx9zgAi7KPoFjH2ewo1W/HYZYqnnnB
Avjlgv+SlXiFwdLE+uEPDiWIaaq5gDEG9dg/81EivIOILoXPOztlkIunIPLqvDDKmbisvTfrXoUQ
IJh/CnlxVtvh/eYo3EDrKbcV3OPHotLZ5jextYh12F252bOkBo3FtMqpT9wkciZIg9+5Y34AcWPG
hiDP/cKvq22YUJSBzYb8IQip/IiSh3UHmTc4knLKzwlIEKIDljHtV8GXpmQPu0n/jF7dXqJATB6r
A2xzAtm+jZIYa2DOU8PAOcabUqs+Dwa174K6Lx1ugJyOqJqKkTpRmXXcJK1blmxSksb/e3ySlppT
okHbq+xoX5eJ5JkgjKXb3B7SzMg7MnR/E2htvc2VwZaLwH4Qji4XyYfYYllckbgfeKIAWesNaX/X
osdJKS1J+GzkngtVVWY7+3cpBWXvkDoTDLne6ViPnc8zfUCUmMbqV+JEq5tWJK7c+XvvsHYQxG2a
GC8TDTfrn8YL03zHAYFfWhr9uSBCFbdUD3BHlj6hy76s6yCAB5S9vvzma41Fz/Q9ZxJzi7x3/BbG
GWj/XVbRDEC0XXMKdo0VStfcCQ/zUQQsFX3pY4ahFj2VOJ2zJXfV9WIUgR42eDbHv5yX0DGvah/M
eYa9xHPTg6UbUYV16npZp0jz+PZq5XWTrq9ii4mHYLS7biySLdAhf01uThi0YYt/nIjSzGD0MYX8
q7UKla09sO9WuuyE4HLB4bsHsfOb0aBULINmYrR5qYYl8z9Q6GuJ7P3Y/XpLOAjI2o4H594EmaFB
0eRZ65JozqKgz9uEbNDZMBb4twZ4rM/vYK/zT+6rUgLL9xSWGpQAqv9H0VFNFJDfUMQJ839dJjJ2
w+AoQCFE/mix7LGXVnvG19EJbt4tpldMAbZ0AMTJSMmoAcMqbaHAsYJQLgb3GFrtMVquxWrlTe/L
On+kfUqPVcy+BluwioZrLh4prE/6eQVlZYf7d2WOPZjcS/IXy+WDGtO6bnEF6HeNHsxemoo8C6Q1
Mrefpb8cXVMH3z8kZzg5qqYHQJQefQrxgvC/v/SP0SiaPUFxFUpWf/m6Fw4KkfZQFakaEWehqJfs
Cbbssg9ZbA81GYARoJQca9PS3iIfMsirA7oohjhMJvgkrtsuiyK3sSgF71Z0Vptt1W9cop/Vv6rp
dPNvyH8lAyslmHquqwLir7SjUB8xeyEr/TgVNsPhpR3Nf715BF4NI3xquxNasL79ptPSoiKivCTJ
M+l+QXaaLgqrvHP95EyKYOO9v6DBbVeaCCK4thp5oDYWAVz91zpnMrilwFB2I4NcWMC7TtIfmtm0
zqympATl/EZAZKXSxC7ARaxXjX4erpjRCshPwjJ36rJ/tpETSNPDUDgitJn+xuCfugG0GeM/kzrL
OIfxbmobBXRX2oZYGf42rimVv82+BuxyuSDT7wBSlCoRG7QzbFBXM4deYxfHE3L1dGNbNnY67MJ3
xNFQB40qhoo2HYdJek0w5AVEni3JVfZfzZ6+wn2CU5eJnC5T+p7ZJbl3z4iLP6jF3bQCkA4Yxu+P
0Y6DSScXDohV2uMHMEPbcpdrAloz6Wd196Sww51n2v6h9fUvPe6e8Wa3n/LEf8bqtvdxVOvUfaBC
nyvrYlKET0Gbohix+yU9lBEVTwyEkuSE8zecMx/zPk/FbOhkFaddf0fTKonznYXczdfyJA9Z1DMr
v9g49xH1XdjfsmusV43zLNciGsvjNhWwNNzSJZDBsL/jBY8/pcRKgSPVtuR0+jIiUDVIhMHyROBj
GxMNYzJ9sXqh5lW3yY/PV6AcjQtFzxg7EfS1ou4E4/QFeQeIcq75w99MJWJxttSdmyMicv3ZEGha
q7mVRP9swv91tCmo39YF3zD96a1kfXDrsFQ3xefIzY6gTfWm06X+rWnDYNaeXK2C0ujIARbtvgoC
a8WpQ1mngbnAzV6Oi/NotJ5t3AtaR9Xtwx7HRd1uEer9H8dHcU+ga2yREvrHgm9VDN9JyNyzd9Re
WnfRDeH3zsmEcbhNIewBApAzY0ZzSWkcY/7B5fCQdTaCSBwX9a5eFxPlvjBdIKrBq87pmdFpU0L3
uEtE2iml4vtjMfDuYs1bqvERj4NhlSnKrj26Pf2iYWbEIuaueT4RWeqoGbF9ih14p4P2mEiifNVB
mQCLkwvi5XdO4wqsVEi7LktDZCdJLCpYdazVHjltp7nMraSCJs6E6oIc1qB8uWunTXF3uEGV+tAv
JeTnoJd62USmo81oAxrNUWSIHcy3KmUv7SNZ3Et0/kz/1R9kB1Ie7m/tshOpHYYwd8TwrMoPwo7Q
uK9JyYqPQqlVxnd41DggpEskyJFCwpZXV3EuR+ysQlL4N3Dwo3eV7m0LV+Y1HCbWUj0Y5GES/OYG
AOGEnA5mz2gaV9Y/rvHlHl5anzU2TBzD4rIufunzbmZah09J30jA9VFS5b29dIFvnI8Vdyc4myEg
S3YpvF4/BUbBNbneLoGy1Ekid3O2IIhshRLyNuqDroyM+W9ChXrjSBM9/9nXorE+NipM0uG/nSjt
krDz2Z7GzN2VzWnGKTfiJVbDaKO/E/Kc+rjJki+L7XQ9/jNNYvFeAHLL42E5TNM7+6i6Tw4h3xD7
Zb+ng/oi2z46HLaNQLCGlkH49vA0Yta/t7Oho31f1HdYSLkVqZvfz35QACPfgNgQI/nrc+eCH4LQ
gmOAJJnCSnbCBjvw7urq31b0rRVHUFUhh62DKq9+kFIJM+c0lzaxOIlMXv4TQmO6USLI5ApoX6FX
TXcn62pM0jCaHWYfoP7jQRjFSryTE0sqa+3zFnmsuU86TN0K0bu0WcSUq0FsbfQJVHnASp1lOm6d
6z+j4JB5jF37bdDxjMJKVAx12qW+Vw5NYbDP/lFMGl3lTeaPWGPHWl1EqMDubu2u/Xq0qqfsmLQh
1tFI/ndiLyclbISHhoQDnJmISrqrlAAGGE8ziseuyD9fVAMSSD8UXZX/02H8Ol9CE8TwAPIIxAq3
ZOxOhc/FmBLPGUmFSCdTFxD3OqMjZMFF9cCUboYA4CAlokyK1EPTlKCZ2l9qBcgfr53yk/HDPJoo
pK46TzcoarqYynBrjcOu2NFOL1Oo8fBVR2BFHDW4vTIvKF1Zp7y/fSQWQKKYMzeRk42IcAWmX64s
M3NwLuHUs66IlO4JLCUIkEKbqLyp9KnpfxpUO1DgZBET9PEj2SilxlOxX/06XYRUlJ1hBQbzmtZ+
Z68GfTjoPFA+ns8GE5FX4ViS6NtLkK8g7/wW6miuchNZZxdV2A7oAAmIpa/yWxwF0eEk35pq4NFc
+7ChjeaDzdoZn/lHR5WmfMrdRnndhFM8+Rgx7VzKIAfFcgse/R0jvoZahsLtscsffUPseBkGoV2d
Z0+g/ZiQN0+Z72/5dAGWYQFzvjrvXQRK1KXG6cKi1vDmpEepVFqNxst2Z7S81BP8sD93sXZ7NGJM
uIyab5xnQbmkgymr0xQO2Wc9NgYnAFsXI5xc9gRF1Aas+cPFFhkz5DvWDvyrbdJHR7gIlrypsKAE
eVUgHQIqWgvYKQE6bdFUX3G1VhaOB73fz65ooumrv0OLHXZDeZ6IWO2LNl+Efxh6oeZdXbCKiJMY
tGf6RX/ItD/k8P4R2TyJfZCngL7r2MBhvBab3Lw/0ujW7T8/bAzrO9DB7WQ9wf11/NO1WWlxyUpO
Vv4tQvsiV3cLYg/khmAeFvzNEKqEDxg7aD/Mljr/uLL4EohlCkmlUrjtKHa5MVQBwoULI0PbA3LV
WMqyz5oD6A9TZvi8OQoGtdIR+2tL5yjQI/AGCdTvZPvckX6Ie5hFDD9cx1JGmSPhiP0QSuOQH8Nt
IJXZBHR9kSO8Z9UhKb9U9R4+rQASk5TCMqt2DI+iHvzkIurWFzK0nYcUVnR4XgkZHc9b27yajvd7
fY/vTPIQAZu4bcf+oiQgM7z/GVrz2TA6lEy0U7m8ssMK90jN8fh/eq8OZbUIXBVo/WZmFcoITDR2
IM/TsupXhS2sJLW+FgGhw0kgRKjPMYmgFfBQkXruehFemlrKJvcfYCB0f9zJHpY6iFXbeEFD30IJ
BLGwBxLDgLx/X2QWY3AI62JYF8VbsG5BCyC9P2cMxZbqX4n2jcA+td6zn9N0LRAX9J2BQF9MvWxt
LWg4JZ2cQImp5nwT8E5VNoD32LRVZ0OAGzVp6Sqa1tMBQZ+jSIkIE32dmt8wT3CQtvCgDcIt5Ih/
oxcfSpFTrA2Nrxk7DLRZDT076ZGP62qkSH/hK2Rwq6N54ROcHyBRiUqZLjJkpyeX/LhbqeoAAkSl
YBdv4heYIo0E71Exwg7AV9SSnvdIlFVDFbudmHwHqDq46VIyWbPCMZ8LHvbkFUuk2ykUyKLu9uLL
CtcwFGSKJyszoyGTEPRSnkEcai3VaQXrgAlVB1uVx15vkKKMdl4SXZc62BrVMETepdvgsaJ1eX8b
IhuE5Jp1GAdwlUIpeGKD18bZ870JdF0/rDDkIJKQHAAcu3tbMNCTMvUx92AEJuEuMT6qeq3/Oeyb
DBtWwlppUU4Zd1aylDryKLKsWSjYYpqOetJT0kmTlir2I07rpa7fMXyeRsR+d8vq3ZkIDQVKqrzc
vpSghoRd+HnpgqTaj28S/CHhThsLR5TlvtkikacdipbgDmLcx3bEyWBmEhYPaWV500SOM92huPqk
vA2Kf8VooVP1N0l26PU5KB/Jle/GlHzjN+e+cFqNlOoAljP9s8hYpsrc+KPZIf/AUQZwp6ycdQSa
o2OqJ3EcH7/UVAnMXEh/6RuF6Q09XKl323gOhpWHbb2tOWXsXC7u96r7NN+MHXkruXHeutOC5dlo
rqqPBmeKn/pZv4WFFXlfjNpwbS1ACnTNTqYqXgrJyFMIL7/+QQGS1ZxiDX24KTjeNYZL/7MJvjEw
/5KDfJ0ioqgLuKZvDqXmPm5kdJYn1GltBllKe1OiXPOF06O8lY9HTkdamwn7IRuHuNfIhd2Tx7Yw
9Af84BeCaDmnzhaEFQhaZvi4PupOauaJ+h3Ovx1S0s+eoyRUCVEaFT8+ELCMSsEmwy2rVkH/0H0D
jDV8MgmCz/0MbYrZD1YguEZ9qNUACEbPaeXBSHUopHh/uu2TkF99DTvIZwtC4l2yTnDpb1+MNCaw
q3f7Pax1v8/t+4bmdBrvIrYkPsttKoCZ9/UL4mHCVKzDjluYhsvvh314mGYbGGx8ASOI1fDDoTBR
y6muUzeOL8L6fHlV0IIWkdcPPijdTAgL3xJaThRtY9WjvUN0yqqsLTTkTy9HOlcd7Y/wfFuRKMZ/
QsBrJfK9yOPpxoohYmeF+GZKK6xpPiNGs2gUWVjQ2IiUp/v8HXNzWI6T3tLoQ2kBE1e+B/dhlGoW
t4/T6pJasS8Hn6dCP12vr5lTfrO3JusDnkls9TwmjFA+zBE3JdYP8+xEUUNCUjpGyktT5WBhEv8w
P7QT0fziIIgvT1Q3LGhcnmnrjX5inMpYCNO2scbgoRMM7fevBd3hN+gTbRDng5NPhyzVie81ysj+
Uu9EsmDGj/dpJonSgMezblq76j9ANRsPN1++c2k2BQLwAfMlw9WNQXaPPEKtPYkSqDVB0fzK2CCx
EkwsVeX3kyGv7HYRQsmWq53bZBErIkGBoCr6wQJQoqqADuZ6e3Q8/uEQ+Dv5/VgalS4Dc5BOPGnJ
XFOzZuekSYLtPCqtSzFB2IWkhcOHESn5OjgQnvJu/y2iG1SBqaG+5jNKbxlNfUSHDWWIbXUctW5o
Y9NWRHRzDec7I4Uo9dZx7jPyt8foU/WwDor1Ord/vapQafn0KmiHNfB9W1DsGwwgwAs6MPVfTTpn
xUKfkHkG1XnHAs5+fY3FEvw6sm+raksfAl8K6Bi39kUZfgazXPyuAixw04Gdiym6QFCL6T5v0FF9
51oO1m2Tp+ihljdECe5yH47MVnKe35nyViQXkH2tR2x40L6qalypuAB6XwreoPFJLgKZoUYVlj43
xapvJ20VavRh2WgbY/O3U0eEkN35NL8D37uZsAIvqvEIsVc4KeZy0TDGlIsNigdoTd0nFnVLnsH5
FQe8iCBDzBqTeZlJ0AG5sv4eSAEVG2s1Z9SRIu/zDE3Bs7lJyyduMW1APNQuGFzLoOzVpDkyL3b+
9AxinP96xNzTjBUn5mQe8zOYWh/6btF7wwvIAokhtBBcqAcX5wGZaeNxQsp/PMQJWJPGX9XlYV1F
HBbHpogdmrDH6RZgoiINPHL/BZoy69ul7EBAI/d5ko9SR+3LWfWhCiezwO7KHqlKdxW1iPx8n2GK
96FMc0aaJeDoEkhTuMe7bbKR0fuKbRe5mX0aMPl51OSbof7hmUCoBJnnwO36ZC0RsKRrI3ngG+MT
BUOFfpS9+hQRky44PHwCAc1uywp4Lw9mERQ5NAtmhqnDQjtOUWOUPhiA4e6cjV57DNCeJRvc1iFZ
gl9JUToVPSFj9UDfU6xyYE85jTGm/dKRrNByzFdyeHKTQCVg2jxvZa4qJO77aKvfvgL5yuLbJSIL
0vzX3ncdOAJ8hS9vqsMP4ohHHgaOsV5g1hp/AlK6hayc6il3gLMpiEwEfWBIlHrZL/wjBtAhWhUO
ICjMGMJG9m9Unp7tO/vL1gWNdprjQdP8+ybQHdcipllnaSWBYZaVlslCWpGdxbCAROO7p6rFUByQ
vRQhOf41G6SjFUgrNgDAsCKjp8tdEN9qfs5Ksi0iCAxJCYjkd9CK7vHdoTUddM69upkrbEbN5Inz
wuF/NTqtya805D56moOam9UHGHDrv3kLYXCBOSE11XTaXvhAQs2QoB+XrqRb36G3Dgsb+7lpR5s8
EG5+5oHwB4oo4+lLRtIbVJqcl+kFd+ET1epQje3sHAkjzsYlZgOX5ABOrkq/CL09h0Wyza8ccK+A
3eW9E0S7X8WSujdMqVqew8cMQuqhGyd0c3BMI+YbOH5yQFF0Np+lYzC9mGboqLK1KCXmnTVtmXO9
X0U+FafW8jsg6xc+QdV58TNqj363Z3pO0xosAjTcQmkERGJsNNqnHZ7JLjrNlE5s9IFg29yX9hNx
MLUtZlZfgPf4pEH4shhdit6u7pLQ50JsGzJ7iegPYiav1qqNRZzotjajocRzE65uLsho7PlmfW5l
wYTBvXzC7w3Kbx/38vD5zyUJrUuHM4dQyFV/eEPWP3PLDswY/grCSPi/xqcGsYqFIFkxOvJ49jbk
zQXqMI2Vm4gNsxqxhrNtxtk1ip92z68BeYUSnE/sFTQchqY09ODxTAItnrDg+gt/D93e0hFrlD0c
yhSHs0+u1IkpQyWksKXEbQ14jx5lwiBCZZ34zQZFcEbX/Ik6LPYPoIrQ2ClckfSrgfN8DxQbdiEj
kfo6wsmVoQMZDQuvLUPxRwMCF3fG019+4WJWfaJOK2bEMl07MjL441LEAQy9DyEu2+iOSydfEf9M
eHLMe6b706dgtzn122cYBtAs4D0PKQPLH0amsFqBQ/sF2FYU375+zXjqx5X61v5At1ImzIE9ku46
S2lwbmf0l/SKBkah7GNWdWr/6JcMsLGTOSxyiEc+hTT5JxZVq5NVb8IM8X7/M8U5lIZVfGTGp3L4
Bm8IEftnkpLfohWGTkiRR4ZaN3PQRYThW8ac6apVKXYQKSxkzVED77nT+yeN2QDFckNyGZgjIzRJ
weMbS2Z6nuaKvFEXZlPOp7teON9TpTmWNtkPYdMCfqDCAyHzcXHIzH5r5RA8Xe6j/sNeEMbGz3La
qw6GNgKSAcRaxT4CHLIZtNG5ef/T1mumXkc5hq5vYHLNrSwlndkzDr83ZZOW8XkLXhUxbMzSiHyC
dwRNSJpuQ/+whoUDAtivVQH07GO78ogOkdGU1DVtg0zf09mZjgwtpIC9+DExjR2dON678YnNRQee
ceNRFkUYiU8NB39PEiMGcsvtIclWX2aasRzDLCAz0fH39lKlia7wy1NQ1q+EV969Bqd4BkMVxrPU
xaW7iUGPF6XkD1f/gke9xCzlcXC7MgT1rCnLZ7UT7N05yMO6qAnyDHpPb3NEYaebXG5E5iYSZwya
Bi9MEROUjYkhEm3J1P3DKV91rUj7km0aULRAPKuv/bRjBac1Vbp1uvMpdFV/ILXXlsO7q1R9YbZ0
OFW+1vzfpV9I6kD2o2PUvP4QJhct23oyrjGmb5GsXjHIeF9Gdrja3s3OOV3gC8y1qfRx61SJAumu
Oa45e8y9K7brREi6MWt2tqc2r7uriVz3cP9c21fcwzILCbhz/hmezEL98u6bVhUvQ0fSj8OaVDkL
rbzhHXvUncqNIk0KExwc9LRMdHhRwe23/qSPwLDE2lR/MiA6vTmlIhEL2ymvnPKB8zvspJOCsz8H
WDFNqa2Qh/uksiPgEPTCuRu1vB/j1eMSxb3t+rWB9trzRQL1BIF6o0iTM8FdOQ3Up8rmDInH+mtf
w/h0up7FIBWJAsaaVRU/9bGb5jv7qtBWj31OPbtcSAA2LhUrxpRXIlNHLWY5RMf56snTWVNKzJcy
QmOA1xa9aYvE/H0tB6zNpTGN2fZc36q6tHzLdAJJMd44/k/+d8wd7SkrgB7Iku74drdyBdUONi7x
MvgqdTUxXM9Bu5N0G1Cmi2K0oaie5rUZu5bkddjZnaIZpjzFf0O7s27nkqR1t80xVF/cp93aS7xX
3VngHqiIO/kTm6xwjjncGCkDX2dnzWaggJt2kvCHJoFE13w3Ek2lUOjozpjRaIvMxAypt9nvgBNV
OyM+T6uhi1pzQGl1C8vl2Nk5O15I3IDQQ2GIgiWAPBjaQBmM4EVBqazZVgo3ostA3oh2HN1OjNhn
Lr2CQYVAyDbO0yt3Cek4wDm4xK8AEp4yjmzyPzqo3K3uroOFII3CHMaggTdb80YiPvo48csrrQTP
mEZgsCNKTWgTZrNbJFsF4APZ+XO4gdmwoEehIBnuz5WzP+fT2HXliHqHUbtcbQ2aJRR0z65wjupj
hDNu7w3EACTMPk5w2Y2dhf8adwi4uNHrQYLc/G2o+XS8tvlCAMRvoQ2O0bO0pGjRSzfG9k1VAeYp
bEmGEkLbY2b9lbLZ67ScSJoYTelW0sx6ulUmVriIp3s+moXyH/pveav9sVeqFZWBtC04Qvy4QNxe
7LtXRP60g27kElPMVSUfZoq1iPOnQNurXLdYPc3sgaahGPlxR0xjGSkp4a1n2e8UIPwEFpIu3FjX
Uw298EjpQ1bz9idd/wRyIwhYdOrVMF+unt5oot7+rL5omO+auPUTwVwjKqEGu+2XSXV1/Eb0bgFD
CGKtMR53jbGatGVOQ2soMotYdPOKWuV3dfdcrOPSqa+RWDMw4NaJacVJuf4Y/hiLoWmkV9U+W5oi
MFxWe4bIgm3q3bcnmmuwIf6GcC2W7x5skyT/tviTkT87EQTlb5ST0xuZXPLl8Yb30bg2cg4nkLuD
DE4Jv7C7dCEJxjph7/6KdiaIN/okibpodftnSPbIdbMq/5Dq32BuMtNCyJlBP27HUxizCNUq7GBY
lGhZ3W7qBacGQ6tQnXHLcEaTHHrefzukkXIt6ionxvL2HS/m7S+2a2WjUZQpk4IZDchcyzwg4027
WBYoUEtn9Qp1ctDNCTaS4EqT/eP/Yn9bn+X7MNruDqHgXgKmv7G+BsoZWmHQov+0ZF9n3JvF9Mnw
2n+sgeywpFLWdRNO6hsi/OSgo7Ms2fN/tFaAkkqUpv1UtN/S45lVBgVGXyaTRVhOgMvJXIYnRNcK
zin5nrnYf9kBBbPdCVshntsmTxXSZAsg3dO2/UF/oNpcb5oiX4k8GHDdbwiBUiAS2fuU0e6an4Tx
AZz4e84S+0GVHVUvI1jBD6iOngRIjtZwGlbSVMXd0mr8s5BVpUmc5OaPqcXDeCtuSiftzcDC252F
+VeVBgFbkcVE+g8DmtoL7F8mi/NBQmpJ8F7J4PEsjqo6ZpzlhOYtMEZKBjiw9HwcMoByolZ/sipA
I3Z9EFarsQuAd2QFPgYu3IiNrwHGSkWqTo75JMW7fMzNNyweBZz5QTMF+RKM4IdBxZhI4nQzC2Oe
kmrGm5R3a2BnxoxJoVVjqfTr8WiIsMJHcyFBZkt0XU8/5o0o1G8xNNCLwixFZgboOYW0Wp39PV3z
5LeUIqef+b127oUZSe2cUt4L9KSUkHDynraaWo0rzvQF35ol7lz8eq///H30Vamno1KnPEr7roSz
sob2hrmX85MbntkMat5/mv6eMm640YkPsnIMXMFi5+u1HP01KBSCfuuQNheA3cvcpYG7jYU//OeJ
RGkDh7Kad9UvKBEnQ1kgo2CgzoGlpC6vERc+aQCIm273TTIL+yQJW+L40k3V1UBV9bTQU1Fe88jo
W8BVRL5jjwBjB8cIgdRn5g/AlQOSXcr8hmbxGmlrvkNLa0N+UjuX3SizMNCxL/XzxpNFdkKHdVAX
b7mmdd6QJWogkVoG+8I6M2ARsnomxPjsZ314+B59CIYD7jiKPcFTs9+lYKk3dSvy0fKGcHBNmvVv
fn56P7P4RVckXgSHUGR5xGYwDQQyjSQU3rZ64UpiaKTg9m2bHGDqobsa1YWGI3qmDfXQBOCriCYR
2hjZvVuT6FmHSOBAV/f5D0qtBVcdFChRXuzvpECqoUsGGidMyKtoCUk5FPV+uoW1vTuexPge7AG1
+hXbss3pxqS+YQrqmuWrZ0uwsS+Uy8/op+ouFUU1MBkpwdvUfMWw2fXiw8yiF0MUY0XdRJnEp+uw
oApfTUbcXX9e/Bvv/ghyQO7boeyAvwvlUt5/xqaXyOIyEC1LX9zgjB174AsuURMZRX8lCFiAgRBu
sDk6CyXQeiFMgvitE8BPV9corOFUvQDyzKdro1iPcd/MEVH25W6/j7fFlNpudU07B5YMmHMvu0Js
1VrqScKq29kyFnYZKD66g5LS2GMgnGtfxJK5wnyr3ridVuq42kurX2JTr9w7v8HsL+SWmi7Ar5AJ
q9sKczgAwyXpv8JTaksNv0ataQ1v71KrO2kYCC/Be7hLgR0aQWVOPXKgXoLKDxrboizHySJhjLLU
maBLjfUKMuR6+VpOjX3KUvWreoYJg0SP1FukCzSpjBGGgbn9D96op/sYJlktSfOtDy9IncuGTknQ
Xx0wLmqXH4w8sFf0kQ/MHSrzkB0Ma1iGAfHOmFDUwLvBmbOGixkgP0XVt3ecuNQYTIPoNBNIlPK0
wPkZq5B6S3sbnjIf+sX5BjYc4NYhwQCHv03W1KgmvwDI4yraRJYyzJ5aaVI/iser5WdTmX7HTYZq
xe4pZx1O9Bo5v4EVPsdyfsYBdM7eA4r/8qasDeYh2UrGLRfJmBMQG5dhLZUEnm8voxx1b53BmbyV
m+eho4Hy98/HNrz2Y270SCWUlPNHGMzYFUDxRLRyTeq9ikdOwibaerTbdYTXZcAO7RS5s3vQ88gR
p2alMHEnhehS1RXZwvmjlQXe6yGG3F/PyPO2NfmRlmv2Vx2jg1RinhyTPeyeAOf9LSoZjsHPEn3Z
LUip0H7llIaTfbs9rw9WUOwoUWAuMDIgUBM/Ji86fvAYeyoCScNoOkK/LIVJvoJo3uwcVNhpfhH1
3ckwAf9Agejt7oA0TPoMaFEo7jABV8zMUg8JfIQV7Q90sxBprLm0vkd5d6FOJrIkm/8ks4g+RdgL
3Qc99zm6wReZVrlGgy16cmW3E94le2UF2YLCOElblAKwk/gzMVcixsBWu5SCLzpLEoiVHnD3SfUf
lvAH5H6QW4TN7DvKrf5BFT0P65WdsSdxn4AGArC2O4BiT7VLuVq6JX/fwLIcRXIV17+lbHkzU3mX
tkQeSqyU1juPFWpFF5TxD7WTgfZRKW+278cFmW0kcEQwcmLFH++RIUEDfOUauwEskq6SFbNH2rS3
2oiguNbwMOnfJ2vLme1bKU5BjzuKYimoon8yBjIkI3VOedBTYpgxALBTAHOvHty2Kkv5VgESOA0j
xghVFLTMJ7HKecffvMa2+QqEIoEIDoYmLq6fSFv4Zw30NPh8+20RrWIGC2p++Ae+gWKMJtCHKMon
x0MjAzgwrru2ilUX0rs6yGGNoEib6nBZeilR3Z1sdMK6pAD/xes7xg4S3OVlsgjelnPSeoQEfPxt
IDhAD816u+TlNyfWQNTGW2vPM8Hcz8n/dqxwqQfQSdgxi60wgAY48C5Vi350U6Dj0LUpIkNWUasf
02u3XQRXQ7J5G4FF3iIosDXqMU65sZwHK5jkljofIeYbEmysmN9rVJS4zersBviNlIKPJE/hknUM
nHLvyYhcwPO341WblhIfsRTOWSHyAesIIqruReflQ9MlOndZxYGjR/6ozfQf7jPsWWwIYuSTAc6/
fUMneZGByHzH/urtRjRtxtz5pBFuBpUlcGAZ9saD37+LWQzdWFsGqdH1//nmkFVaSqoglqiQNlu5
P96Dhwg0i1DiCN7lei5lJfmSpUO4X8g+2gqGxrkMY4BPTZg9rRwq35pMtMzxPVcXez0DsF+2Vbq3
POQmP3i6u6NnrtV4c0Sz8P9VCxjNvw926fTY9azMXant+nkskcijs7Kws+cf38dMsOOESkY0byDJ
QBYysxB2FuFjPH2HzlBix4dnb3GlaJgJKjcW2wTWaeSvaRCzTcBPHfaxjtPm2DF2taKsUJOzDf1k
KsRtRxv4gRIQJzJCIyyo8m8t6f4jOEScHAUwb6usci14P4CWu0Fqcx3dCx4XiTnnUBFO0UuDjFu5
gIC/yHqwsKE5nlmXZDfLeP/gdl549kKopPqhaj25HXSuWdLL/DmS0yaO4ypKlQ76P86lNAJKPoC8
KwY9qzN7GoeA/GcjPZGTTaBnef8vm242onWHJj5FYVLiD9w2ZpZfRusjmC65m4EEE/UnwDIdnewv
4C1nF5FGtBDhAOyUlVKxBgXgYqc3p3Pyw6hPGXbb1FKax8HFAKskuTi41rn9yroEZElzXNvZJJVu
3rKhib4z0GFlk9KfUCrJJS3uCPdxCxF0y+6G/ZKdZBOgYDQBTVwdv0shCKljMJNzvsOO/nYSus5N
fP5cPfpTUu+hLI/bomu4mc/BN53rcO5kPRVcq/tnTnVGLSp1KYR0jFi55o7kzU9pK6TH5G0RKthE
RrmptU7yPAP/5qKF9T+uarDqVV94TQJS7zHUGQoBVDbeAc6Bksv9O183VdjTLMc/JQJAGqAkfawZ
KL0+ArcSajVK0LDHA5Kn/c1GyNxlFxgX6YR7Joe4gpCjQGuQnvYJjdhA5lgjuKKUznZm9fU+BZl5
Wvp9XZUNqPnN+iioxpk7/OejNb7aNA7pZ946zxW1Pd/WB0OentakL13qFQ0FvHXXJ5ZsEZgvz6W4
2zWqM4z33akGToq/WVMMg7Zh0YgEaj/wTbo219i3DCfXcE+pyKeudPwOFXWw0ZzLqwChQpu/zN9G
TxweALPNvdIFblwQoa2an7XGIAOwFIh1tk6GGHkxOcqoK2UAqlec9Uz8kiytbcg4TvP+ah2PFAiD
91J1v1v909CZf1MMwzTw5+1q0SE7brvdHvyZvf9MRUF/sG5yeJtAH+wAQl4qpqU/FyOv1BJ2dEkw
sByDN2LUiPHeo9QibEoCv0q9tNiG62EbMdaC2I8xFqKIl6rzkC3sEH2T+xKVypLT9Uvc1Ti3pRaV
F8jk1OtZJqET/v22IML68jlUI5CBE7PxwuqUKN6CyeVOlXLZx6OXUrY4S2lmGC44b3UpcX7hfCab
V7/1BTZjeoSv96usAYCAa0r3N04Rs0MQkyLfqXZXtUIYmokpQc+WzFD0hohMU53DdrnDsk7EIRF3
YXO7qYXVFvwuP+7tgVj7oQtuRQXOIESzWtSllYyEWdtDhBiV2INP5p7e8tqYtQL1D9dQmUoYitNJ
Oc7NGHs2RYIfbHqRzaqD1xZtZBOSdlXxukaRDdEfm3j1NVFf3gkYMNLo4SslpiNzdaSI2fhW10XW
jlnmo4ZsT37vPp4+xDV9b4st3jg6YGJbZ9N5KPp9yknoITFg5ggsKO+8Xufk3ikdOhWtqmGj5IFB
DoaN9uuUq1tEwo50f24KbUEhuMrAM1s0OxLd24saUmaVs+iwrVF2A6lQLA7QfqAxMvj2/oU0ocUw
QY8NRN+rC9r9lulm8Uw1AweaMxufLJO6MbhEE8P//rDK2XfgByY4+mdxP41qLIbndkgP+Ls9p03Y
E7iWOPmPFl0igCqrRnI7rpIuZdclSD8yWsiK5VXlt7VdkqQNEtOa70Cxyd41ZFvFON4ZJL/Qth0x
a7+rqsa0IbNPGwTIH/sSJqYbJhF0G1xHv5bcxJPydmJsiuZecnU6T1ThV4O9myGGYiS7fZDeObWG
cmZekPZJ39bifd3pnlgT1CEeLp0L6r7VTAuqjAPPQGp9lBH8vxnjbJWizHQgSseBbGYc6F60xiC1
3HfQkPBEqmH9vb+L04DyXbWgE/TgG7p92MssdBVH7mieI1hxe/Gie7GHc9K87hPLtgA+AVlYetxo
n7fGXUAIvMJG6uQSniyqgchIYWKhl+V017odexvOIdsMCth76HCug159QY/0f+tQRpqAHmCPygdS
YX6cnLNHwuaj/8S7jNBvTLiudYwyUNadsu5Op1eC0DrCsfExwkM2gwD9grEvzJ2Kvv3Pn4aPsSAQ
fhO41Jg9jJ6YHVFhrI0/QUoAMjeNS1fSfacjXxTeu34R44h7gSsXxucBamoTRQKIzQDiVt7Rn7tD
8iXc1jOUrXfjT9RY4clvk/6bEcIq6K0eayMZckATm3ycGyeMKhT1lytf9CWlamyJSRK86jsbj7Vh
Ge94IOpXINlPXL14K9Pq5BSA3Ywv6OyTW5/84yBFfHxJ4o1nMR5QQK9bAD0XHq5Ge83ssUG9S+sb
1n3kAjq/BNBAiGRgLzRSWYg/JuMbjyMykBP8ManK/tRUYWu1QMUMZsdVpK7vaP9FmCDxgaIEx6qF
x7sSojr8wpbSrZqwzgTJAEn+jkYGYuQpvL5poZLhVReVUowhsfOq1ls7yy8070t8JWsDWPhfBdBp
6OljbN777s6kSu92h3D1SJ1X7s/AJkbxR1o2Jajhbju6RzZ6sL8SIMZMS7IV5v+LRtnxtv1okjjg
56C3QqIkg2vpYqfhbAHCfZY291F4JnXsbW7lIR5/jP+YLuEzAE/2UOaW6WCLhrzDazqhabbVRb0e
WdY/TQPg+XOULNFILo/xo+AoXjCSol5FrL/U4enM0aYekhm75AiWMcYvoP3uq7dr1WeZGwjZo8UC
KDmNKx4deNhrinPGj9P9AMPBS6kqyT5pgHqW5XG/H3yLjulQOsWWWIxXy9vvFW5UIsWcccA48SKQ
GU6cRuxKf79jU3h+AGoCF1JUI8ri8PidpBGgF6YM5aGvL4tbvxsyEx7ceDiMBU8AZHHXUvFD38yF
jKKeZBpTwFFKjoH0s67zys9iHbfiqkqZDsJ4JzLtffD7xEV1jTw0DH2kkzseukfSCwUno0aEOnbp
aXESAZv/Bsow4Twd5gOrQm+m5Wg6rtsfeuiHTiv1FmQ6QDZ3YSwhHo14lzw5aj/GTsUNHlkzN4fB
xA9v/w0lOhDZUVYGAHHjfuzp47T0sO0rHmlkYK0oE+lUNIBmp6OAqJtNgsKXLegiGv7/e+AI2SXD
4rO3RjJI2uPR6NuGv8QqG3ZMPKvaAmBAXxK9Rmbv1TKOWeP+tk3X+mwxLNxitbsylGRPVGy/5V3M
MHB1v8XyIbQ8XrB9Aabx/SfcGPbB2Aw9A2fwJqnR0NcH+a1rCYaugFnF16AWdDOF3MOXK9MWoXJj
qbRGyRZPNzOsOek4P/ADZoGuwbTVDFL0KIH9fGx77SKOeI+rRISKA3p8boA6vLj5ncINc73va7c9
LLt5Tm1QvT9IT7XwOUn/1/wrBW/q2VflEaGHx+RKCuoeloWuwPhejX5wlcV29n3KEzim7ESEZmmj
E8zhCgBdN8hJP4QFJJMCGwRGOa+nYYDK3d5Lr3tp0IYiiTFD1bJ0EtZzhBCk7ypN2pbHURyNC+HS
P5xRIFPzSzByGonnmcq1YGI/lbM5rI3CAJXebFNSXyZ3fzR2wIdxtDZIVYfbv6KLR39Ubwkqn5W2
4INvSGc0DdeskgMtJVIo7sCtzBoU+wLHIG41kphrsNWP3wfho92kE9DzcQ9iEdeirKWG44fHHCFh
jx4oLOnySGVUaUUdOg2WkGd7bSfKMUX5SXx9upFvFANwoP0erX9Dwxlctq67G80t/SbKSCstXpPH
3grl5Rhw/pnLDOVrJjnPP5IKY7bM2oY24o6PgHDd1jqTLoycdDtmV1GDlcpvJ6tRVimccBPGtJdT
eUFG8GsZ0G4U8VDbp+snCl9QsebuUk2ZRVnTPKyo+xK6F7yxWqX7BdeaMJo4o75NbrkF+jx6yeTV
CDSouL1mnndnRU6pviFDm3rTiq41DJ/CMnFiRBPgapk/OGsmFjUCk39Qr7OIMQAECKZkuFyYzO1H
Up+a5D9av+6HbUhY4bWMC6W/Tzq1VGLABOpQXDIkrr4ceInDXq6GFLQB5FjpmrWvynH7DXLetUO4
+ki6dvbeuHxy6N9xIkf/GFDRWH/AoYVM59jRkUx/4QZ4xvwXdXnmEg+Vu0MHTw2LPnmxFOZSLnYe
bbHqhdFt4v/35T1Lx2yPTIyhgwFvxJpWvN6ApFi+WjIn6YTqwfydNxNVtPvJXIJdnF00is957EM6
Hl3r0rR2619ztMss+Itnm59jPaL75Z7UlbZbh2Op+ATXbJjffmb1Z+yxU0YQDikMngNxkJjHUK9U
2x7uiFsm8K002teyhOeyx29TeOFnQ88ILB8mjglT18XvJ0GBEVtaWkpfPYi7FPKb7055XQxL1FbA
aE1dditRNrzU3MThhb309Q38eAO1F1P8HaDrKFLL7nPOoLgM1QstHjX38iBUpUqhRLIJ8BL+WXOu
vbQO9b7SwsWBbA2VsGxqnbLryAEBlQAcyeDwoZndi24zqFkOHgGrcvkkcMUP/4iC8l48JU8RFQVy
9lbdP7w7qcCQvp7g4ooAHB/HaZCusgtz3neTvNzSn5T6dHPnjPCZ9dLvWRvD/tdNHE8JNisLCjpZ
KNLHg6BEI24BwFRYDo0gGNyUf1maLyh70+PA4du6weicIjTNerpEBSXLlcG0E8iezfhjay5nXN7j
StJd4ncxEk796LWvrYp7ahvgz43+BGx1rRyg/l+ktguNcfRwzFnpE24vVDa5Pop7txULsF0Fei8F
V2hQFqqlFMbVC9S2g0wMklZcgXSfkHiuk7n3mrrcKcYgbZ19ja83TB3ZoSElHsPsO2tCgRqL60ii
JJNXxODadsH5qWiS0UU5BxKghxRL0hTp5OHEufICRUFhXJpwkABaLokTp4oGBwCryGS/CzthkR6C
B0XWDFyLMqjpI9xKY+nyoRqFNhBN/Jc4plrUrqJz9mHncbLIs50AqaVOIl140apjOhJZCfBYjlap
HtN4ftN3etdhBZn4+pSP5yk/UTTg7J1Tgnze+jI5Ibqmxxow4Fcy5Z5J/UpiY9b2pEo3I1RKE7Ed
1O9DK2ERxSDMFU6DcaAv6Hxm5rHwcG4UjRDmhIavyxy9Qle3k5OLIM8h9bbe0hAkZIZSvDW9d/7j
4M/KZlr3hmFZsEmhqSt6KEDzapEXXk+xINoBB+kv5q9Yg9sNnpPsQdA/Z7AjGXLpD/Ame7aijC6D
fozThZdfWX7xJdeIM9eWIkp5M0h/8W8g9bXwDLZyYExxOYemdrXeapFraI1Hxz0aRws8ohTYNnmG
EI5C0oYOHRT8zbJ+q0Nv48Z6VNZy5Yyzlnxd4tiUjI6LjSTJbWn9GYq6pOJ5EO8LcQVSCuXbLs6M
ZLQ6K3uYHd6L5eBLLk6LT7fTzYqHvYARl0VPKmGKFv8uCsaMBYtR5blW9dixk2jrlemESexK8c8u
7jUP/l5ITeIyZ7gt8lNb+H8eL19+usC7egL6M3UMwkY88r+xA2I+5M2LluS0m2U0PBbrRrOjiSw7
2d4B1JPN4SdH0Eh0hCg+IvoXzoCrsqxqaCMXrVIOH1P80CxXpkWbdkY6nj7nYIT7hffG3m90XsZU
9kJ6bOP7qnMZjOITz9z6jx21PnV1tfym2Vz8ryRsr4Kv1/KKDRJ1cgqwS+qx81EaBlL9SbB7kvGY
QhIXLIsuW3l4wUDQj9HUidsWr/JKCRzlfqJ8Miz4CEyCpN9T3cWSnClq65KKdVQ4QTe4i2lxCbJd
dQNobY9Pt4bOXWkr/2LQ62p4X64Xm5u4XaUvZtAVcTRt8j1qRvKKPZr3TPFsrw/CkBAniEE3qxOx
UpgwoXd1rOmFZ3IW0l9jwxuo7t4F5br7bB4LuSmj9hmno7ntrzDI9xEdx02uflkLYd1O1rKc4qMg
LbIGi/s4lEldCeaiRuxwKGuKGGrI0HTAoHprEjrKYRHtlrhWCTEEOIiE660mLrUUEzdQQ2Tvb0xz
ev6OTsbjP1zwtaYLGkicHThhSNHSWq22LDVBksCanOvRPxXdBMJoN4FPpQcaqzKhDy2aKL1sbM9B
cZfE3g7sxj+T/VIySMdVb27R6uhojxOtukkKkqBT8nRhNshvpWfcQYTj81WXmduQUI04Xb8hdpsY
QQ85F6p0GcY4Q2cuJ3kEG5PFllphap+nxM/ehSAAxTAshWxnNtp5nLArp//NqtU89BdgeuhYG6Z6
ifKKTKlcaz5Bz6KRFUR3OWTzbyYhxQh+6b2MYvCY0p9dzTJ8HT+wGfZ6wl5AHDUL+/OTt85RGuyA
DPLjbp33r7H2xGLJwnYmeN2QFRiUNjVgVERntF7aXy1K8rw3sNSuYvPgM9/6NDLEMuZhIZPJDbJ8
bcVOW81+sDh7m9ON5WuPteAPudp3pU+sk68NlUZiuPKSG2P8TEukNwvvPUYYbc7AdutJYMlGC6pG
aFbqSy4FVlcWK1JuEFLFD+TU+yQ4tzLvmNqhLHHRO9PbbdXP8QY/kDcmywMkpiZzM5fBkf2NUh2e
JRt3Kxt8PP7DWtUiSdL7gZEyOJUGTIkP0j0PQiKSZk75VFgidQh/suK7DRXhGCC1qzCaHnrguqGP
pECbGbS9OUk/aUEmkwcyDN63z79rcYSoqCaFmA1cASzW1cYBLLCOvVCQU8uplWK4KV+ldTtbnGf7
8o/dm0fQwPxAiw2Fo48NtdDI5lW/yhYwpUx7SaMx1wVLo2L6x22f67ZoNerDOul82NhcpjwV4SBq
LGgYtdYMwBkihk0l0BKauK/fQ4f0sAOVIko+BN5/Anshef6VoFxxTQdlJxaq0rZCuWcIE7wTU1Dh
/BC38qkprSJ9taUQCSS7F1k5Dkp8tx5TqfVeBeUq2SnG84esN2PHZebRQJ81UFY/sHVm45cLM9L3
lJb8itc1M0OLT0XYLelPtU4PDnjibKd4J6FXsfcIGdw0Lfwm7eXySolQI+sgLNC6+hFq3uap9LWi
TjuE6b70SIL6LBK/w5XpDOPvwIUU7jc+xokTK7+42szHyzVnzkoJAtn9ur6jWhtnbIbJn35NEUeM
8lKU0kgIhs4xCmoVg5W1Xc4Q2CFWpr2zGcqd3ROWRNpADLePo0Q1lJN0p5ifaZVWOPQcL8tsPjQZ
tCInJ+MIdxhWJovAvlAt7odpVn407m6NMrif8PkBM1lqqY5+QdnR/OkYbW/8LKlu5GaI9fMLRmfm
dAKHWnV+TsiWF1eceY5CdhC7zdfb/ZrTWBKXimbsb527AR4/AUAme61acyLD5El+ufUJgs3kEPYr
RlbM6F1UsGCpSB0lU5Gbn12YdvKW3k6ZEqfuyPXQX0XlseDwTwo8lt2hDZFHE3kVqghiSz8iQghK
y/fnnL01ytZnIVd7EnAE/Q+eslwsdruFwzORMyFoRdjXI2e4EttUOAAperXGvIqlpFDhwrVbXzw6
UzvS5qZvWOIo8ftU5ennAm8MRQoDIEwO1T6cxSjrCFqQhC7Z2asNQPxwNQMTI3VoaCvReMzsP+4V
y+/J8D5HgqyG99VMGnCnrLE72nEB50KhzpAoY2AKzMftOXrS72CIOM8vgHB7T6oIC9xHMZ9pG9Jx
C2r7QqaUFO7IutnyhReztZ97JTib7WqE+ll8njs1CbwzVrxKzA7fYqbuaRuO9mY5JyTFwseAtjpc
cVEjCreXxm6vyMR0SXkMZu4Lr3fJG1q/AvWDdIA6Fg3gYVA3aItbXkmljtcDcep2g7DQ/f/rYrjm
wW1reIPbL+SGgeHKa8cai4BH7/KDOpErfLLmiWBOh2rVrK2jliAZpJwROc9G4Nrp4oUwW17qjA6O
/JqjMVrLyRbltxC+J2fDKfO4tA7wSWHtmByG76DmVgJldHX9AGoYxh1v8vGqgz9YkL++wTpIJ2Yy
E4UljjjyZQn69oeYOX9FLvvnwxQmDK/zjD/FkIu+ZNHeJFPlq94aX5FlXmoCeHJ1sxsdJFUWNfpG
9b/o2c7vus7Iqzp0WUSQXmWbwz9laJ24uooPOqp3nxPt9VEIJhTAaQT/JrP1g/SVNBp6dEXQQCxs
r7F1Ypf9noHBbnaAjXZp19HUYKveRt6cbB2CFOKQ8ioscl9fFoLl9Y+TDijq+kBCdEszn69jJNQ0
nTz7YhaXW8BwsEVpQr2Ih4TkpYOpq8ihQOMfoBuobnZmYi5MOBmeqqCSo9berzJJ/YpJOff/z+ec
ZOTg0OIfa+QZRNs4l/eZyYbr8E8aUzx7lTtapXRl5YoXEP241OyhDFpMtPsDOe+X0NupEm+xBUOs
2ZLmbMZogsxpIl1mM0HQhq+XTg6l0tuTf7wN5lMawa6wCtGCO2J0QlTZxfwGFbGrz+WNJ6vkFgsh
WaJ6FSFj+wdt6goyTM4v2kVJYTA1VbsK4vuUa8jJ50w2cWAjW1LKSwfEqiOW9Ov+8xURM3CGOP3A
SEX2QojcF7wIdQQdcCP56QVp6VaXDfoVrt4HTpjoF5MYdwCV0JU5MjoG50swnShzfCHZ5vdG2Xpr
7ZMDDUoBdTGz+K8wDD4KGtXVf8fa77LI0LNIHXN7HS4ZF7fpAegfgL5JikWQsJxuJAh6/Pwo+h+r
OOLhx8m8Xahvp3zYESc18yDLhopyWlpW7rprqNcVUHZDOtXOm+4jYFB7ynrgVR5HoRU0EpAkSURI
AX+wrNOqRK/iIrxcjAjGTXCRRhIfub3qmgchW8Khd0J3jsawPTzZOrYTWvPocn3sG2+ZP/cfing0
f30bCPE3dMaOp6ZfxJdDHzddBVrxcoO+hwPCyn1HwsXlMN+g1mKJrcA2/lmzBkVKNBhZTfnVfHgZ
xM2WHR1gs9VNV7cH6PLq/szizhnlY3hrqWZG98TPi7D/eLq5mtbTvOmEjNYZqBOqeyp9yVitRJE3
ac6eo7IFYz2wsgcv0Inwtjk9qkRMRMrdE91+ovTErBSh1ChXKuat/TF8HUMyDLdXzcHL+Nro6uKR
SLmwwEsMb9Vm2DIijfI8ILx01WMx44DYKfKvJNfZWPtlJmFukdKx/Uzx4GlJjs+gbHuH7i+KnCX9
1UsRTa0yDhLCYqL3qjIHViLB6K6FidJf9Tloh8dEUzMJa5mh0tbHUMLIvIHN94Yyghwmoo9IGzr9
gbL5dboDYcGVGEMzB9YAfYUOEZFtbVdPl+Ki8eX89DTMK/GOV9kENnhwzVyntJtGDU3qQSVqgZgU
7CF3FZT0Xaz2NE+XiQYerqm+WR3onkqnDavoIWF8dd4Jdhg/fIpkeGUiYhO9qtSKpFvSTunj4CRK
oID6iTnwiGjHFkqE6YPe7gBnDqHzV9slTfg/dtEqrTVQPb4LQRo5MDH9XDNzUs+V0gHYkvL2knj2
hqqd5VrsGIjAq0q4XrbQ+klsH0hibSMCcDb0/CxQ08TvxNP5gECQU09KgQJxpBqfx7eTMq0lzr9I
0GJ5liTx5LbuPPUVbrXFNDO5X/3rMR/qHCW5uSBAxKISVnfK99oy+KszVMNAzdZPWOyAhZCSKHko
7+iahfMyAKfKOQv12fcJ9BtKFTX1Uu45OkiEwWm02BxxvctA7PcsK+ItZLpdN8XOcclVIZEviy1i
EDbpYm8lFySlYImbV6QKbD4/s8xNwuBzZK6+Vn2Adgch9mQ8GH+4BWQG/cH/ZyQN+PdjE9mWJgAB
c2Uvi9MtNVu7IsEpuK3xJ154ZKNy6Y0ZQzGGbbIw9svY34BVle1unJmeX9V5nnED8dw3uzPd9Law
QT0lKJCMvSKVpSCgQLHR6XGNaGLjFr0a1Ki48+TLjS308ZoXhT7aA0F0CpVoN+fZpif0hTV5Slft
DCqNfPenk4t1FqrRpg2FmxaI0dHdFUje2ADn04/yhtkYCsLz8Inr0AUEfCPHa3yZ0mgTSS6FAuSU
7nlV0ULjh7oPS9ngY/dGr0WWmxjwYbiZUD2f2fGEmRyH8TBatqrgTU0S6af19aQ8uw48VGc2RlGz
XUb4RFnyrSVW2RssMVkMYWnK8Hy9ggDW+nesS3wlnw/MwuD0hrFu256FuKpGYzY4dPB8eouoABN/
Clvo2cdFguEi8wsXX8D9Pdq10lX9KRhKwSl8SjlG+yOc3yZe0LLAM1aZdm4MX3DsX9/kC2H/7kAl
JdAD9t+BlyOV4yUvGiziRV5QEz/qXmE19Y8gVT0bdZfNr0XUUtUqYU0tekgiUCCGZcfvboB6EDek
mcFImCYDYIfUWGzaqcgRixyvWWuxk1KsnQyQrXu/Wlsb0UPzDwbd3CzoeTUiF8cf4J8uuLF39hX6
DqN3RJq3RGd1P10Q3TLqAd7/VZJ1WYLmE3ptLDpbaZfz+nnSQ+evNJyzZdE4mvIZyaz08LeDOiyP
LqNEP9JP1UoLMx1BAhxrSDuqcpOKYVO9AzCYs+zUmVsVpZDmdFlyj/DuYecR0nh+mqBdJnA1L70W
2V96MUIMiLizha6Efz0E7KiQAkZOghMijQl8x5UI7mIrA4BFsAZiTAngiyaCM4IXKzDZHg7Dbz4Q
A/Fanrz6Ww3zoSY1q4E9CI/yBut4lifbeaB6hJQCQw9VnSs8rxEp9+9IyHSQxNq6DDmNGvm5pNq5
kJo8zqj/o7a+oE1ghzKbtYTjIzpMayvLaz6BU+pLj849qs+sR2i4fQZzKSc2/BsfxU/y5jWNZ1sk
jbT9FMcAux2zMHLxogoGr+mrj2D6mNCx9ssFyPAuK3ED2I7BtCbXqVY+8dBTbZdIC2cipcD43Lh2
4dFnRgbe29Yg8v8bH8JNh0mpCnN2qgi+8t2RjuKQ7L1BezWHOMJQlLCj8zC7FdXMexT42Z/9ZPOq
TqaTM8HVfF4Oc/sYS+27vo4N4RH7mZoMtYXvheOwe1p9nf3tzuXglVWxwLPYvp4JAumnMnmVeS3g
L8+qEL2vznWYp1h3y1ElBCP6AQ03RSDHcf9hzHOs73X/w81/9nFyiLJnmlOzTT98Q0FvNmpqOWb0
PQzGg6HNpzsxGGfU57xyNrXeXREEwUf85jmFNYDb5Ip+Gn2Ia7E5t8yH2fpCeTJ7hRx6BdhI9by5
aeaT3TrIQ8qtX0tR5wud/qg94hXtKAbZtEnuwBZE2kWZwkbNDchVJD3GjAZryvvbxysowDQBONpv
pkxnuOPtuOcUH8o/5vIx4OFdc5NRtfxqUx59cxGoEhz1ebY/UczdCodldu+usgHQ7QEDGhleRKuP
dRfMawAsVn7mEKDheuNAEfPE8Po1GSBdPi+dpkq7OlPi9Ja2KPC/38RtxRuayO2d5PqEknl1MdtO
emCv/J5tRKWtfLbOTlhMZjVUigeeuv/H8DNqXbkrN661rqHU3ec3+7saH5OUh9lFSnhAg+jcsp16
vKKuh5+tk4Ha/ZmmYD1BvR0Gh1bzN8+JNDyXW2iEJVG7Scmpl6a5hbkIXdEWYiZ2h3omA3wMaI6p
PIYsxXVlERsZjXZZEBdFX2FEL0y8LKSiUUN5//krW12kgt/Ctke93tJ/Bhf3kE641kimcJemPUL7
aQaHn9v2Hn/QPgjseIj8LPfBDeO3b+Hk/A83ubwz7Hdf7I60PguO+h+ek6l2fU7CZdbHVHaVifxQ
Jx0S7XXf6o7+xg3YhpsROHyG9PmpQrRzSIP8EkaqmSoHo8DR92jL1r0TeJjtPpYdCgVLslYHzFCI
mFkR/baI1vEfFkacrKu/147MuXOwEwUIVinRuqqnBeDE6RmZwO09kdYDyJl7C2YuGPfr+PGQA/N7
YOA25VD+YIh25dnsTGK47jLfr/os4vojGlo/+aNfUeZbRmAuh+Q6TmAIk7G/4kdXkh2EHwVcghoO
DgfYiWSryCGkm7V8dff1ji7BNpeq/o3utwRT/6ZM76GlSSAZrFwyPVpQg7DjRKZRsz1YCBAYCtgw
Ridj0HdHuC1a9VsxIsuxHKm+tLn+oLoiea3HfFHcxV4fT8M5C7WrQK7IH33z164OUjGQeTBBQpRM
q61518L2oOIgSmKrVF6LJ7hzft2PULAqAXcQ8baZKy/rTaQP4Ijdpy0JHd3ISiX5K2QyusGBT2c9
ep7RAK3G4jv9v6mA4t4wr7jOQ6gKLyIVjR3MREZRNgEflSqz1k3k0y2BHuKmx+vDxn++6fDxLSdl
ZwL+lYxThNC7Q058niee7aytusdwa2RCaTboXisSH9HLT9HeZcZYot+11a8lV+m2LKlHHYEbB9Wl
jocG1ZZj6x6ZCM5yQc9/C+hb4RDVDZ7vZ/bJBRwHIaMDFlH4sbCQWxdLOtZQgqBp1jOuLF6QztQQ
BL8dHY5KXrf0OlS69oZ81xsCmcOn3MY8q7s3ul1nvpleSKbg/0aaNaqdBLZtFlVYJM2yMaUEUvyV
aa7fwp+as8wcBNaNnVoFIRHTp22i0QGe7E7A0Gavn9no2wuE076GccuRnJLmqZQ09YX01p+Yk2xm
CNWRT6pSKwSlTWeRx9qn48xZGlznfc+FWvKAMOKpTc3nnMYOY39fK3NTvfHy0ZQegbGthUMpTOrD
um61kOjS+nvXv1Vg+ZmqW6gxCElY6T322O6GeivV7Qu6T/BmkfM2UKg87kntC033DhlvyQfLSGXn
whPs11YWCl19duit0Vi6w/lZ6slDuFg+jZ/eDb1bF09Z1X5p1PV2DhubeLqDDVAY//pRDI3UtHZl
0o5j+me2+2oAyCIws7vmbucE83Q2nLoougWk9OCRH7KpfYywDCGvwMcZZbCaP+FMG74fHjMSEn9K
JPrNd/3d+fKHnfDijkCmxLMKfLerb6Zyu3NjmBhfXC2FOnLRhNh1wbcE9AqgW93kncLgGyF/8GEK
9rQV2Yzk5b7uVgG0j1Qk1APVSMuEYqMSersZfFMRJZcDHug5LELEu5nrIWdngyiCCuRa7dNX/yJJ
MDD4Dt3prrtq9F0BTsOiE+EQ1f7+8WqRRIWRJk9MQaoy1AJGIVtIEnd/F8l7N9fi2iiJCscLeRCm
5GFr2lY+0MWzQ+2BNGSDxs5XGK23M27gPys25PwLu3uJb6bj7cbd6xK9inmEy8jRaD1J7j3Zf7di
17w0/I8H1NyiW2XW7BLOL+tIp/zBMnl7B8L+ysNUuBawjMM/KGHJJLDDVlz61HpxrFRDQzLXyhGt
x1kR5pA3mlcU50TCeifX0eYUy2/FuABydt+lgiWzyZT0BqPu6gKYTzOB31k4SGRLz4XVDNSrsiGf
AeIcv5lxf8pQ/D9cT6OqUKdRHfpqqmgN3oKV0uWoZDRY/Q0wjj1SybnKbBK2qTRawkFi+4Hpluyu
vDliZtAkizYvh2vT4WfY6B3H90uLE8mdakwJGEhi5nq/2gNJa0LvaZiXHHg+1CUDAtYjqG1I4KmO
edYdslFE2vsOb7j4tZ2Itgn56tZKF8MjSiYsy/8pOoyWkfN8+oupbC9A68bpcA2WHxzI5TTukR/B
X1/KBYfZziyQzBtt5Jr0cltBd5QB3h2NAPKk9gfsi7bsFYEWDPKj6YK4KQqz7OkJjwbhy0QkSx4J
fAdTRhhWmlsGUb+rSB5BWksl3tg9Z0vASKkjzGtsFXPpoTo1fBeiMw7HQ0Iss9G7GPSlzsmiaSOF
D2uPIkYBsx2YShnJeIPQ/fXWj5zGJoVQS3CG+rjV8ZyH5sIgRYzdXbja5qj7lfZED5Kty83+m+tQ
IW20w+QZ+QfAlUG5Z5Qnav5YPNdjF6X/X5OoP84mxJNhA1aox9UOlze4jD4fR6rH4+xiqNO1xw+r
Tj1yl4TzNmhEEzBzCr1XULzMXUTNiRvB/85Ey12ZZbbux1glnRyb9n0Q16uVU43ks9DBUqfN2OOu
pg5uPf6EqbKzFAm1NrluO+DvQtA9xZa+tj85amj0F7h4d5GcHOzki2o2EiT93FDw15WeYmmnEwm3
VKh643x3oMqliY9aYYn8pQtMLjUBjhRC9UUqcIpFdKfEN2a50FCDJF05cuoXcevrXx30tHRD4mPs
RJ4idh1qxE6QzicSeqDHFFAwLD4WA0lUbudVd/G5A/8YFwA5+6j4Nn6mDK+i3P3X5y2vak5NZBId
4uEbV+uAZOogQjKsC9xrzblXjfP9D1iJ6lmOgtaXoCRmJIse1kARvyQTHwATU6s3t9ElHjVCuTjO
21Xbj+ma1+Hp2YM0Ct3X1nz38uG6SPzI+ibAEYee7RoBL8PmC1I4dcXCtM4hnGkqURU5X1175DlG
0YaKm7w4tPJDzWlyvaCkGQ7xQnMxvLvFNHLomzi60G3wLPDg8IZtqJONsNm0zVmZwF8eHXF4IB+t
AMIth/SoluN7B6x39GKcsoxhrxkn0iH5UqIc/NK58PAJYF+skcmh0xqMnfXx98eyKQCU9RKvULOQ
aDmqCjyi6uLwUpay4X58X+7RI6EtYztdZRJBk6+LMgptEQPvAPT0TrcLTsVrhcPnBEx/UBTdcN9/
U1GRJV1IB+R9fh5p5/VCDy7UaWirzhKCN/XXGGzLHPhnn7D/3jZmwdX+3XD+o5WCSWJO1oRvfWBm
ELdaWgwMuQSJhum1joSJjyIkk3P/DZ6V0RibIoDXJRn0DSCitk2fqqwkKhGWEbHoinA+9tibWzFi
BbeAVFPg7nXJpTFjGT0OA1YsP1d2xwnsfKLTRt9Mvs2P1YNN27+EiQCMVc/SCLqM/WkGh8wS8NDu
oalGNyWtvnPnY2npFTufklEWjGtAKE+0q48dMmY5TLRRHKL/YHZceFasROEEPlnddlCP29nGugFh
0dG5W5XKeXFSlM+WT2wgrqL66KxChWX4sqk7CcadQ0qN3FuYXUaboc2LP2IE1ZcgVcEsi/gmUamx
Uidpnco/igLWbT9eDsG5kPzmanwKupdkorgz4Hj5wzfr1Uecqw1wWGMOXOoDS3/dg7ZNKmpjyUgj
+VWpuHeGSL98EWbznQj9YOarIOU2K10MPjft4peFnDNU8P3dlYGxiAUikHxBbAhf3N8fved7O11x
Slb0Fyw15R0arMKBrhENgzluvfOKxMi1vIBK1teXWW/5HHSFkx+O35PicIYKP+zcLA1frX+S8IKg
1kS1DUDyuv3zrcW78IOdA/4e+5SMjFP4rtec5qERmMG/TobDPGXPDPRKJrc1fD/leJmqKL12eIgp
8yNRIU7cbEphcdzug4LceZu44M5lWFnyMfazKIqQRQMDbiOzrGHKOsFr8BuY37MCng/J1MdT7VEy
g/vEhVnWlogLVhK5iTYbYjbBZHMf4KI2w3fFY6LiW51Bbf5uzWzb2O4uvhlHf5Zw8glYWatXKGbr
nYl28pvCAshq/RpGeh85DxVBCdVxO/OB32yX04izlq1UDGDw8xBFzsueyDlM6mYHw2OS44YJnzaT
u3AOyQNJQIfi8OzDYY7UnWVhI92U1q7gZXdU+W6LujoPOtKk5BI28azK9f/BJ1WgZiyANvsFRjpS
/V2Ky43ZaBAzd1IfWxfec7wASbWbFjTuAEH/lQceqDxMkjpTzRrxinJAT3LMxk2qHZGlFnrvgG6X
JWxeg1cqMYTGj8HsX4lbNDucG+7xMYwSx07hxGwYXZg75dLPm0KFZm6/Ofwtwf1AMkenKMacbQny
G4AmZL7Qg8Zwoktrrp68RMmkNxHMN3gkcDvup+tiIrk9YjpF5r0niCwkjNX7YKnBpPo3qXgJot63
wgULa6Y0cBQxu+yCi78o7mIFatcredwNGl+ggoPX9Zl0iKwlW6MZIauLW8pKSCoVP5+9QhgjwrWy
X1Veuw0ZBCuATsssSxoCVnO/z4qcCydpSJtAdov5jr4cCCDr5HBqPVQrsknYaZfFpGPGhVlEvtQL
o8QkJI2ImDEDXQqIXL5xI3VDqaVhkWca4iwxz8FrnD9Ymk4qfKv4IqAx7eCIDOB6XYS2+80Fnbx/
RfMr0FfdFH6nfbcw7I1incbfK225qbkwKyAJDXs/uF4uEcsQui73gSupWlBxVzEQFEYoe/2ObR4p
iq4IVqJ3/OF1Meob+2dqL3QzoQjU/s9oSV8eUXPJ8yz/ZAgJQBaLOjDi7U7RCedY/Gwq8WbKJnVL
DV5Cktd6IkrHzMFvyQtaJioEHYZNjXVIA9fpRZ0zObOx6fLVGRYQHrL5mqnvTkJyNp9R1tUovmmW
Ib4Zw7d0s8CXEh0KK5QwgZKQPAsKzeJPCpaL/wVQP/u0nd89IHc34ic6DkmTU+YjAqEkWM9UA3Hr
N7AdTiPJ7rzMiwhtD653D1APQyq5VNBxv77bCIyJdr+rdcDqp+EQeLU/EHgrxhz//gTxB0Ch7p3c
uZoLKExqy1FqV8TJhXmXP1mOilGlzD4b0+8B+ME0ja2v0bP9jpTnmBJ0ECb/SXajOShKeTh1pi5P
gL1xhY5XASUPRkudDNj6KbZ4SjZvvPOvGuAxzRGrafXoJ0Ush2AxMOkg5jrYhfFaRmnUEYQOgSgA
sFrZwH/AVbdWoAsYM7y5Dwtw8sKKDLtqe+DtnVWXFhF+PSeXxcZ8mGPeBMAJXgE2exKYbVSIPwfG
AfiIAF3yXYdGak9h/TpGF21tuoZbt66Sgbzg3O5SLqV1OBnQJRKF4feht7Dp36OVBHydUB709nqu
gHPJY6ZlMH3OF+fDhmR6eHUbJYw6Z00Yy3wrzqHlmjEbGQx6B7vkyI0DBd8tWfGZoACqDDB2bZXF
YsldapbQ1VWsvPOEPAo6j5kdUDXS3Ravk78Q/cGOceem/hvflzvkJWJzOTMhslGnCq5JAFyZXY1h
JQPt5zA5R6uG7L8QW2aDqhvNo54lJ+y6p+D7Zp7WTdMF27mQoMW1bzsnuQlxOhg3xtkSyRM3qORp
9NXs4UiDcmGbhCvWFPoPSFTwMlSCeQLkrgrWekugnPxISUw6tVI8oDGnbhsE3wVlvqMVRpQbAWEi
PfqcTaGfR4NJZpay27ViKMCRVQrJWMvt7bgc420dVB3IjgkjO1C12DSRgZMSP/lEZ6wgmUsiVndg
vmXYh8SW0kAH56o3aoUTzHm39f8jEQSew7xOPKLblZajt7L8iAdrH0wJk/iS5/F5uGFerwi2Ou/n
dQs0KdaSusSQYeuO/CDygu+lhAhCUHwSbDp9R4J7s9ls7ns7dwEpWGtbOmA7oIujnRUftDWxbMGZ
QwV06M+IwuvnXot+MCsNVnkSNKG/aEL+m3Zf7/r3yXCwbJn3eDCTGjI3IlAiwDCaAMFuMzc6AosT
XCxXs/DwQN1lnLgRDmAVhk9X0J4oED1ElS8Jn8AvqU+30DALOyX36F1rNcJwhTaJ7/ARNqVidB4Z
OYX7JCOqZKUdVigyep+3T/rU242FS6cHpJ1A4RPfIqv5sfDffNMoHEokUDBS0nBzLvA6XhlmOg+C
IojbjTkBGs/6+QpEAgCHiNdtU4MMrYNKoe5PB+x222hhy0ks42K3wKxbZXaevzS4fadX2Go6sBb1
4GJ4TVQJS5EnQp8vQ9lW50zUwI0keBIg+g1TXlL0XLeYcER+TlnsD5FDWC3UnEjEQAynQYGkcDty
F4dCtNzxnTxaIxvWu1IXnfAa9r4SJw0g6vFirfonFp6Xm2d1NN1VbWXK1ffPbG0VzgT3UOfbwhFv
h0cpdQ9cQsD21ce7EhsKXSyGuxBo10KO8oOwL/mc8KjrnwebQkImAApXoK4W+4jKNPO6E8nWYPSQ
CFpKncT91S40+nKdJUhV3EzBk4aHSHG46CXOjeL/y5xlpIhnDFfWimqns88enCd5e3yux1jzYy8a
KgV0mcSy2ruMKCeEMRLUztQNGQJyDgGFLOZfnHB6DR99UIBj38I2+25QNYqKj9g2Lfz7b84gC552
FyIyaIa0tPiFULQcntYnRfNzXlC8hK/nL1IcU+Pr2WqE6cKhrntUxBrPelNLyFNZFwsvjlSbdoB/
oqdvBODHVz1b7THetMqgN7JVulQ53icefzipI5GvAw/JXsn5sjQzoozBaGO9uMht4j3Zm7BfITo/
zM3XBO3ncEjMiA15n4EzW6SwaUEOsTPGqeNB2sF+LNRHMJ6jA3bgZXUjvWBf6IzKdi7cE3FKLfhJ
rhuaGZBVTGtIR05Uu5xwEia8sk/B6Ttyo2LYMy5N+CPoCV6YZGR++5Gsx2adqgoErwgN6j3sxt3K
BEoujQeDucZA66udfdxudvHVrMjwq11/mVp7TPNRknGfg9mwiQbnUJzE0iXndJuERrI+kYIwZ+SZ
XhmW9h5SKFRoOStF2kg5ZJQ7RyUKeDCaJFN+WlgmuRd95B+7QfPduVa0e1lggsrA5ztW9EO30rQX
MKuO+Fv2UIHE6L5LJs8IquqgU6Wj4Z7ulZqUNwF4q0Hdz+QaXu0aFpHdGHlx9QXxg6ipaPR8dk5H
svVsFTrFOdBZQEPVc/hK0uN3y3+mEXwTNJSQtb2v7685fOc+Zn/yCgRigtcklI5pU5lJCvzD3+sP
FYZBVj8qHeRyaJy27OJ0WU/uhUrSknC/QCqpAtXL/0o2JiLBTXRetDCbCNj9qyeGZFh1OAbsit2U
p//AfZiiFmgU9oMQGRINqXma0C0a3pqDhcvCCpDiNZaqdgQP6TYs35vaVzA086E46rkeajQIMITj
QZNBiRdPK5qnsWJwEMKCpKfvckHxvtGmJVYKmcTyb9xfTYjeuRuf62GjFD9OK00V6XsgE+t6cEj9
Q+CVpW9GFqYCd5yyu0S0472N9OgClGi8WEJI/WryBc1wdtNo2ePHAZxmQYNJeItfUdimG5kpG5+H
BpPTOLW+iGUu1EXfIczSnjqHJiJUQ9PlqULqbVzwUhm+VUQJHN1yLoSN+vBoFsi2zRZe19En6MzH
mGQBGi64ue1xnhDLf578sIjunTG/sYEapKZuaCqzgCPxwuBkybgPHCJ3ldYQ25bLM+GNTIZzY09A
94UnPRFJiZ05fVPxojIlW1gzxAyvk760VXl2WXGVsphi2zwTuuRiFUs/lEWqCCkkdladJtTM5W/x
wm5w58sXRJEoT57lTNVY/CvLrJkHGkQOq/tA6zGzImTi5s8jBnnogCYSYZKMEjP+ldUbgVJ8xD6U
+/MTHsAYUlz8ZAEPm3awo+PAci0ImJibsxytOHJEVdDx5EPzkEwz4P4VK5wf+NgPMahnITmu7rIJ
L9EwqdTIG2HZnh/0rNZC33jpdcsbtWKAg7DfG0QIrMvIr6nOj96JqwTFc1RhNpYNXsj52ECCl0Hl
IOhttrJF0MbXUkTf2nQTKmj14/pgNJ5+UbCDrP5R4eITKIibMKzNZBmSGsn4C5HO9E7IBBZLNVwr
C6/uOy2TL5jJ2zJSxi1OMQlixuIFG/9IVcqGFcSNvBeDPB4ZX6lQtkn+O5I9GAocvMcX5djf5g5y
U3X+dP3MqIasEynoCMMgYcdieOxWkpPSjuVfKq0vYTyKOIjEM/PxMA4Mje9TsjqKhcE9mU2aLeRk
cEIrND9ls72HL7lrMD5CoA94kX+JHekuVkOWOL/FyfMWhgvJabUTKdvuZYcNYG2EAFOS3BgxqzF7
DYh/k80aq9jk0F8qjg9L+CVjWNBMl492J348swk8MoFsAb8ogSYPcXbGmhk4bWTLZkwjDUAenqZj
KHXowhCZU1HO2kFiByAn0VSM/3bY+16o9usySKlNx0qt8ZO13CAzXfls8cPo1axtactkVWyErKir
IdfgwJZdT7dRAtyOTABR+CLzjOZYA6E+bRnGSHH+zrAFU3fw4LXSlsH4v7AAPYcuLye+b754+VnZ
nD/2vOuSOVsfY4F0qJvdI5cftXJ+WLstw4E0k9ypyRsnj+Rvw+j9wWUFATfrnb0WmFKPrAMYtwRD
NppUKovSEOk9w15WvsX/EWGW5zw74tWDJVEmSlcM9xJNhA1AmTWqc+Qrqo4NFGShmSf+i18Z0J0i
IiZ3xZRiGKXZDLT/OjGMF+DqVhEzGXl6tCA8yuqW8f4El6F7X5w6Xj+oRVCFhQdgyJ4nMh4d0xYR
Xznpx8qcGUwnsfRPvATovdMS4pI/9E8NZcB/3tdUVd6HMURNN/w+Q/u0GFG+4AvNbUjVaqWbZoRc
IRvoCOn2IJ/QJ1rOuNEXkXiHKZi7nFrNAvbGtIhmCMrp1mjqj35Bb8p5lioWQgTyYqYrI+ZU5G/h
0LCbZpTpLHRPeyvELeTwz/QaekTpxoxYPirNcl0KlQQUpfdlzc8dVbNFR84uZ240Rdqg+JuDb+iQ
MQXfLazUs48impFmqtEpNOMujzRBOWhiDvjKB4Pa+BeNyI6y/gz41h7M3eWEw87M1Tjjbq/2b2yp
YihK20nSguXcJJ/8YGYVAodC05GDLRFh/1ZHNq4CfD+8fxmzHi8okcuVOn0iLrQAbz3ZYXLd0H7S
YsrqychgB1bkQgx8UWyjWu7qzdWgo3UMY1cNj5jWElOuTrLqE/QE/dokXBVmwvzk+WOoOxMutbzI
ytGDghuxylzvtaa2m8pgx3Ee9FmP5YmjsdZi5ScetQgsn04yDTbcUagNr+ngECsr3PaJ1ufdFKqB
3j2Ykt7rlkkBKcqichyIXf7uUSyYA1I3GN+rGFU7bLDgLgZvaq/xGH0FSAHFFocAcC1SwsRGend2
0Ro9XDFt//IZrYjuJXre3ziCdr2ZR9ISQ3ZRUih8iEFH005avvPmfN05+Ba/vc1R477Yo7QPrTpL
K9WPxVmtxhZR5exMDhINKUdL+pD5sBEYAdOArpoY3CP3iByBK9F+lFIr7EqNugnpoZcere44/ZvU
xopl2Ci3nH8ShxBLSCkIJ/0vTdJfthxRlWAXBg7n8LyKm7edJ0FU4VgjdapGn0X8NUVk3JjaHJIS
53nA2wURcZOxm1IZPbscIsOefumZrh16fv3oLW2RrbJGkA0rnPinw3uy+JrqSBAA6MOybiTIcnjE
GlZG+tcNCa2Ji4nGOw1sRZnKmcs13aSHRjCXuN6mfJhtxGB1D1ph3J2fnZfXFiLLjhw82vdQs7aX
i/HBcbqmL2agidoj6pib0KKUWNGJc9Zfye9ZsBBcg1pE5aHJsk4XdTDb0NuhTX3vmk5z8PuSF0ms
WxrmrJxFW6Swoy5IGoqtQvNZ/62kpzqguvGCxxb5oZaeqgs2d6NXwiey3ZGIVeafIMgeFj/B0q5h
U7s1xwwrZUq+P+PrTZbEi6layDCAu3wmqcVorWdO9ODKxW5BD+0wQL9NHMgKt/tUwrbJLlUOS36D
EZfzc23k6YqHTRDVLQCgNp9WZmTcwZet5dP1mE3CItHRQ305tISsBLy6eEvLSbeMjofY4Bv0EP8r
dOSV80OxFHS5nnBJMi0s854+JwLzArFHK4PutIVQwxMp2w/1wQ90la+XNl6Qp/AMowWjMMYh6tma
yMDaFJ/kcLAEpP83EjjLMVsKPi4O3gPDuYpM1hFk7rNSwPxH5TIuKLuaFbIa2mesLNyctlkNwqHz
cO7petQUOBoLkWR5oB4OaDkbPBX8YruBxlaxjMTPLR44F++n+wMgzAOREpn53yKQsPFAKLuUz4Dk
z0e0GfZ2bocsJFeFF98eNsFnTrnVEM3ZG4yY3WSyS4v/rIIaYV+TRK9kZIzBYWQ9N/L0UfdYaUsX
FDRD0/D12Sqhp2AOvJv80E+T0qumWHrdjkz5tJcv2yi4F1O9jtocCG00cI6AuSjAYxd863winUTx
nokHETmMXgJfIidJAlcE70NmvRD+mUxge3UDJff0BNnAR7H1YpKTnZsaEepyz8p9bQKL7TfM0EUK
cxcOoY94p0pjNZ5m38Wi8Zz/F2xipAjQ+6kQC9gKwccUQRHK52xHt4/9c2PC6ym7+6MN3u19CXU7
jZWdA8VyB3kgVl9nf48K4jUuLvjuPZqSfXIiIE8gFJLG+3jTzYJh0iumwFcvliFVHaa3JK31ujyV
BnuDODY5JRId5iV1wj54fE0vjqiFH7ZXaPGWwEnzFkV0fpM5+7ucNyR0X4Iu4zj5JxxZBl2hhSG9
RO/8Xl4v1+xNDEB0VfLk54lOzXXxSUXnts5Iz8KoSl+p0gp4lMzRdlxUJPbyT2iEnYQj9Mg0QGAB
oooNgOzeXGQMw2TVCzi+ZIJYRj97Axf5R42hiFCLiok+q8QkAlLviL6/9NIv52JzZTBiHp1/6fbf
DDaVg6UUO9kXCkQjqN7NNcp6MhNTS6Ay2MRJ5b68JhnjbuBCqzBbeBrjB76Se7d+bB+Te/M1kjNE
cJ8azXfNN3ruugCgAjeaqsr/dDZq8CwkpTo0J7BCdrCDCXE7KhP8Ls1pyqqirhwUr7hrWYau0KVl
g+sQ00Pm1jV4cy6fHSS+xTMRI5C8VhKUSkSaWaFvo21xFNKrnTMJ+z+DSgbC86/ogF1VR9BCIB0+
PNQkk+2DxK7QYK9D+/xE7ijB9LJHnvf7T37mLSUljbwD1h8sDYvfn7ptbkEhUH0OydLMDBfsvMp7
i1nJAn4DKqx7tQWGls2xcwN4dZoUJ87rS6AQDRNB0m4iIm/jZPokbv3o1sNMygOWBjqV7zqgqJZc
7SLgASbkjh7TyOkUDV+Ap+lAyNtrWBEMw3NUibqQqQ9hxcGiLM99CQzNG8d6D8Kek62O3Y5giO8D
PWRgqGhNcAmU1sJoLr3/qKusinx7c/QuKCvlfcw+fRJGYfeVAXQHYbAjoeKd4/Jo0lxMfWX0BDwy
xg/vhxYOEy4pKFwTPLWxKSkM8K4hD6PzGxyGG1fzgqfvvtLr2Jhfh7ARVWNZA681nq0pu5Mje3uC
7+2CPVocuN1IuDQQ/tPRJPxPrXo2iHMUYfscGnSWe/fFdlIDBZlMKF9hzmjcDqT/RUQm4Nq/VwIv
ZtZOaj3bDzawI3zymkoTTIEl3tRhBWYej1EJmkilIv2+A1qE0K9fAvqPzqJgo0cCcW88V/t63rn+
w+Xm4bT/AjOPsHHpew/BKvDVmgNWbYGJl5sfsLFy4YJo9ULXqjN04WUbkmKn7L+22g7Ooj0T+OoZ
1p/ozVaKwI0nKbB3S36AdXMwmKpKPvhgm/oGTOn1PIJdT5DUQov+ePsZEHqGvWy3wJxX+NFg0+c8
hT52T3+kiH8Q+MPxPhTducARQhzqZBAfYiJUA5lfiQJqCEewpkJs3ddT8DCNoxgJf3W+flqlgWr1
NsRt2VY0nH7jnqj4vWbGGqcP+hsgpQDoFgaU0oNF7Rb8IfkOw6eVioUpwReeqxF22cdA4xAIOsYd
xvJF+fkZaOSCITjAtMjigLQj63J6pGzukoKiKLxrhy0MzeRFEKmvxkJEWqiFaVU6VMSmrXYSzPm2
25srfy98j510zMrwmYw6N3nCecybBoT8wQdOFqFfnAlgxMjyIhV6Pf9lJw1I3n+69n7/suB8u+gC
/6S4GJE0Lb/72iXNMkSNUseIRxvD2tYE7vcY0ju3SOO6e3GeXEd6wEqFGKXZ/qXJxG4/sErSQCMS
3l/Gd10SUZ17LitqzbfFoOE3eWda6MJxemJ3eJp9wNv3aUhV/oaLRii4oTSSh1GZg23mvWRFZdwt
0aqpFqT/9C+11pjvOkn+38Q52ZKWAkJMTjggNUpajwslF4MjaUb1XF2ZMyB879+swuDBsa8hYCOr
zk48m8dLXsjwgNBRleFTbCOjCQy5kHNsJp32K3IDSxeSrE7oqpHg4IVRyjLgDkAd4xyfPXqfP7vT
9hqcracNcqdmPtIF7Kdz1oYEHcxt5WGuyODOiRThl4gulUP/UUfKmAv6Ja533NqSrk/rtVpJHD25
bKpmGXIxZENa/HNhrq7B6OK1vxSWubOSJ8t/I0DUVio1uIiaQf2Y+XAIVv5rM7qBw0fzxtpwrxJh
MbWoqO1ci9N9dzA6cAX9u48qP8yqaET8PnCT8jqpaIgSZ61JKTgpFHJDe6gP2tdRQdruxKUoq6vA
Y8Lwl1EGdigpZwNLD7VV0SdBj5CDj9hvRL1gLKAW2wmS2N4rMdFPzcIXbDxzwxOQ9ALmbsrhZGIi
OBTtd7ZorGX3cByFftL/3f5V7ABfhD8fB9wHIE6vIHPwArbyltKc76C3jeQ3uvLiger10KHoC0uL
uwnw4Prgr+/S2Yz+SYRKH2zhcU++Mp6ZWOlCpCCLi5gLA2cQt+s/WXMCYkqboZUyEobI6JTt99JC
IU1iP7ufN3bcefssqpqO5lFT7WPgE8FV0RjsJ0h35YQ1INbIkKDJP1m79+wPLGjTAVWT6XJAgpts
T672rjhxMH8bzAv+y33OFI0KRrO4Q07cu0nbADmWUEJbcJyjoqqTQZ+2wwvFJuk/F8Pr1VAcDmSh
Q0LxTu1ZgDZniDT+ABDXX83ZdfDNtT9K0Hjv5nsFqmvrTcE8p9fQdgORlw8AqNYgwu2CQXsB53d6
TEwBObWQjoHn/DPvWaoP1wOKBH0Qbj38Tf2jLXA+dDb23nmtZV7hMP/IoR1NctwWv3e32hYPb+Uf
7r5QuID+lRus1vngyYbtWGnDEwKlw/pGNk0W7vGxCqJgBpORgMn6iLUbDOLsuVfiX18agT+D1Gp3
WsKAIkKBo96VAues9AyPgjmH+ll5TCo3ll9WuHQ+pIdFrzVka3fV7LGY9oxu6wKFYX38eT3tHmrX
viISnk6jxHwAPnOiWj4hMjTPlY2mgYqdL72xj4BAvnlx3hoCMZYnNFLWJKKxeVEs5T9c83nw5Lfx
tdWEW5du9FoJCNQaxYXEEI1tEL1ejeIg5Qf/BgRQgOPnS1GO0oOl0gLeI8cQk+1XlrPFHjyOEh7/
XXiJAcgxEQiCi0MrVdG+HntQAoclLiOqjGbEPtUOw7/i9h5piPjlnpRjSL2bx5fhtz1TjyJ0+FER
raOTXmADJXIWnrx5euPNmm9asFYUSjcUL0KtOynM6JbloaxwbnfyTi4EYNyE6bnggVhZ4ssubBBN
pauA6bWDBue1H6Scai87giNakcVKwGZtCxuP2Wbz05oWj44e1xaxpPMQ/bNLvfJKDL8vBssOizBy
qN3MHdZdh9cntAVGFi1Phx3/5n89kuG1BLT6FWzN8jcOFCyr7bNlzaNkrTUATO7LnadaPPgDNDce
m13yGk591jvquXMHHwcXmXX2Ndrk05UU5nPOKRopBI071UFWPHc7BLdhh2mnjxtsqJfsBrnuJTA5
EG2HHjkrGqcJJY6AsgeDzMghbo+U/GAJsQgHdGvMEwWXosHqUhO3lO5TISRZZS+zlT9aOxPkYiRl
sy8WAvU4Li+q32pPVa7VEIylviwJMnG+m3tqo8qWb6fsq5OxK+qoPdAbHycA18afbFixPkfEew4R
ZpilmeptzzELlwi6KFWKndOh8exRH5CgdEkTtDVFrqA1GMAf2v/8SX0bvDdMQm0Z1Le7ok4ToBCO
iZz7jf45u4sPZ4DJQ0QiS6Dj4yccXuEm08Rz50KkPwLZr2xmACQxK7szzeYVS/vXX2+Edb/MGnEb
/GofVYhoAeKi0dQW553Ry5ROWfSW9o1TboFXoMJCcSypHTKiQoqMQE/JUuzy3QiE+t6GLjAH5NDY
3mPuMaTlRSOa2ssxqSgAGCEeo5eipsL8AW8QXCgzTSXSTgVpYNyNShV4xvEe9aiQ4US07H3uE8jL
5snr+o8ikLtCRWCyt0lsHmMTiRA2iEQVnZiSsPZ8esYXNQ4v6zdOOZI9izuR7gvylozQuyGA3/+Y
PQjQ9w1Z2Xu7p7GMmVECTUJk1FlVkxXRaqXUAENN8vjbaaZcfrvTzl4TFjOIZxOmLn+mIpodhf6F
6T23Y8b2t2OgnbOlCx0MjaXbgktnAGeYeBLaE3oJqwfg0VVUJ3OOG8OkhH61CF5kG09NwVDQfHLo
JzIv6tVeNtroJEs+wDsetB/S+/3Wib/cGfTow9fOlk+D0f6SAK9+l+i1nwB/fDoKwO7kjD0rY/Cl
thD3f2u0zIzJk5iWOrGtV35NUXS3QPwJu7DuI0UD09CM7CgaAm9xoxK3kzt0ApCeb4BXuj1xFUUo
gWif4E/YU+UEC3yfI7lI+CXA+5mRAmUogjsYBApst6L5tH+RZV1slzcPXjY4t9qCHl5aU1DCmW6E
+jO46N3BYFnrNO6hocdnjpcy+VnIRbDCzdVasJGF+qhdzdd/UFKDv0WQSS0s/py/nwiMFb58t9iD
6KE0OwhiC5EFGXF9bJ6lqLoq23S1Q3BPT5FmdMuRSImoszJDwv64wgh7nrxftaMjxnrws+Gc+ZEY
lToKgoL5qrrnXVmo0onCvXX2pl84Maowveccv8Tk5IAVaLX0K9gSjNcBeItJHdTYNav5bb1WRbTr
x5t9deos8tbvdKrYYfpgr8a1ZRVTrBZ4nMkqlH1xFBa5nPAPFk7a8LTiUvpVqpP6izXReZ6VdzJE
h52uXJuhj6yeI7QnXbhc7464L0AHM1aXsq5AtY6+gAiqL+c+5A+7NIpsz9WoK1BZCmw/6Xd18uP3
IfmtW6ESqxWhcWnBf0shpRtZZWQvyLDUE07WBPOjnbWutDezZGj6vsdrfa/VXVhwHsbNAskT1t0I
Dnvrtjz9Kx8gFR2SPIKVUkfQewWAiTqQhoxr4SrIojc4RdteF71Z8mE2+Mjps9f0rukWLtVsy9U7
1CePgnGGGMXnpG1Slcs0d48ww0TG/xL3/H3ypAX969sFUkEWSU2ITR78+G6DYRXuNnrpXmbEQIQ3
Ogyc3Atxwf6Njkzq5ivCBP1IljhvZQc0S+AOYV5OrKg0UVsdjTuK1m9Hybfcq+omOtQ7p3o3+aMB
h8rISliD1ElUeKazjMBWMMHQaIyFNaX4Z21hWMHEjUkiGa1W820ZEGA0RXVvM34gc/kKS2S+CxoF
bjNvDYkMKG7VNPFTJj44eWwB0c0c0UDzcdls2TeFW3Snzdgn28uS5sd1d3g0aUzmeY9nRqhdd2ba
FopqSZYEOiMRfuI9610eh40PjdHbLVGf76QwzhU39NCKMh4fMjkUceV7dxO9WGOvlzGgFAGaukTA
jyfma+Vs0hVvHC/Kjk9xY5pFywxqm2wRtCWxoxF8bBAvY8gYsv7Ze/RGsUWMN03g4pHIC9qpdkbH
Amiuwb69RRYruEOLhOJL+J5uiHDrCareP+vA/WN2EX2pDrE5MnpkW8Lbmqy+lbStJll3ufKZqyJ0
dQ2FBhEmJ8NBZnGzw0xQgDUgcMgOvKZP4SA0eMNZ2yU7zucbEe/WkjnEo/aoOq1AaYpUVh1VQ9nH
urWaobhH8ddDf4SPzCbVEzudsXEDNKeh4v6vENsn91B3VybXLPlkzNEfXELR3Pgbt9o5Fm14bhFN
ZVB4FNV800LPvVLCCHHFWq52kGMFydOv7UQ5uEo9ySckw1lxe2ouTEm/c10sWLqCGhLZRxMOVGc4
ZPgaskW1MErrMo83TBHA0SOkmEQGxILPvL7GZw33ZEx/KXxtUeA9OeGdHxxIeWRdy0WBDLwWhR/N
6f4wmiHBY2UYkfOLtgNHeVsLdi73YMB95U13ev+1Rne41uRRtLmfJHlaSocyHefpI5oaVPK8mYHz
SilmgAnFP7AVRGNporgn14TbmysUCBf0UTNXl5hR45H0+HMrlcMPqgx/FwhRfRXg3wlhDRLWV/BK
nv+KSV+ckaKkvbS7hdmcghJB73f/fcp2Vdf5y1W/k30FPT9AlhROp4zOXk2RSsqzS6xRNjGe9IA7
spw/tWtVI0c4W1ZmfoprYWNJR+JhkFRINkawqF8/WuqkNsi2YJQNzmZ0IxOvIm8GREsV+09znLvb
xK31QEUMqs91yhwcwia4Zmzjabr3YELs7eZNIsgEZvsURYFuNturz7hIp5d7nYeAc9yEXxZ7jRSO
y6bPwVfvtoXRzKRlICElv1MHPw7kbAR7zv0Y5ps9pP4XL0y8hMo5Q9Zn95eFIUKi6F2IkSMyfeV3
RC511tDdQ33w/8IskHeDyGKk0GTKEaJJ0nJr6sXB2mm+LPk9dyn1MhPORedMrZ7IOy/EkKXzzhXK
aUMXkHkiBELGOAP7cel2jCcrSmRdlyGyM3Rz/GNpKy5XxPkYln7uJ3iKRjbvr9F+B1QavaE4IXLG
pkY9SMICyNO519jXOnk3MQiEWFtvsKFKqjFWZ4FKtMz5hyJ0tuZNqoig/3z0hKA143YLS7tTzBTt
Qt1TRbAIzX3ID1MpOIkXdi+PNKp2bnpU7AMBIj7GwLmuszjXFlO/Aez//7yF5kgKQ8IlkMB0rKqn
GwL50Yl6ks7V5Wou34J0pG2ZTNjHtrOpo1hsFsNPruD7DKuzFrkA3Rk4HKuQ7qfATz4uVof+zLVf
/MjPMhSQw2Zk/hjnBDH7E5u3tEaBZ5lYGvq2yUMHgt2ujlNNJoCKOdL/1nj4ZvcjQf0GwfU3Z/04
rc/m87mNK3cpM8aVvcYoWQUl44nCbvBiPuahi86pf/H2jX360sPzq+5F2KE9A1ZgTA6n3morgEk2
BHchQUM1Se3cYWK97sWCPyx2C41yfByqq867CvEGUa+WD4SpkQl+4XqztwWnXPIJZpaNEGfYNEmi
ZOorIuonxxnWWl+IVlxj5m4Iv/P9mxVBLlC1OhJVyQeCZsc7zWuRtEvkawlUoCW7d0UjRibu5O+7
4HRzYO8QWnf/kd9IMjuvzsj1+r2IbacNM77uA3mI6TlNBSYgRkjg6wX0suoFj9Ss5cbCOgVxhKLZ
G1U7m6j+gT6zrKDiiPo00MeslAH3wBhJgfQ31jAI/+nDSSiHSoOdy30I90h8Qkre34n++tbKUC4I
JFpwmd543eAO/fT0WtNaLksxSWwv0LHNcHnV7m3kRwq7Y4rNP9C+5IDxVRkA9vvgwkHUuI6V6gwE
ArdtN5CpGI/XChWG2elYNUovynaL3mucTAmHT6j3IF2iPYlFP+rVhqhpWB+ruGXiFsrRMe5a7bcl
SJ08rMUvpBemjbLa/gBjvrmvi6v2ct+s0bH9Ua45LwQf51HTn+tKH5qZin0n6zRBacmoFnDybkOF
6T/Oe9AkeIL2tFKhsKBBAsCAnjBQY2OzrqKoZhj1QR16+c3bf3K6Im1Hfu+rPAuj468AEpLVtvUr
w5T/ziaKqmA5beQ540sIuoY2b/QokBYTxZV2+wRlOtUDdUZcO9rKWEBUPXj9nhIFodAQJ01Z+Hr5
UjAvskGsn0gyuBsg65i9FMzr7l1oXLpSFD4PoxZ2ZsO9jlmNXvOHdGRySlLC864swowOqfvlS7yg
bVflbFu3DHk4KyqHJ9z+KRcX4jjxI5taneBZ1SPHGptFGrggnNeKHTGeZ7M25pk0QOT7hyFQ8SxH
bK7tvbBXr2NUhL1IvrNUqlQ0wX9E1vI8LSNvxOYxewUn2Amo2nACcKe1ZbNdXvqvHMN6XNJ2KaTm
Xbmz/HIn/3WJqwNRegestbXs0Z+2dYmokgYPZ+Pt8ONSvr6a1MG/6C+bWHrGSxU40eWYdCrUStFU
KpA5fhlduQJZuH0XPybH9/4mTgTUotSOobQ8yEUhH0b5fjctAjcWFyCvVjDbNC5XIqgNjMfOIYlQ
W3uClZsh1t8MSvINnu7dehENUHeY2P2Ise4gppXiGTsCTCOaClflfEFfHWazgtRLM7DQ0C9Epfb0
xAvGp6gPJn93mCg85QDP73jXUfQ8EKFrvG15ImTFXRlncF7TsWKofuQ7NSMlixvn/XNqxBDH3d79
jee2kdk23ETT1nukrD9nVDgoQl47LR21S5t0cGVkyw8w8jHiMuq90i4IgFDHNf23PTJyEeU9L/JK
kHV0zl5tJpO6XX1p2d2RI2a9LHMZerqOWbwf9MdiarCng+KZBzt2fcNPpcJ208ARlHy+ar6a7Bwk
Xnegj/2TeVga3lDm25EaZK5CIOHiEySorjub4oB7Jf6s5Z4geTk+zsEhv3TpoeCLJ+nsuQ/3DioP
urbL6B6UXdd8IdbrT39WIE3T101snfVngUqeyMGqPYg7JyOUzJ4dqT9KSCz/ssqC54H9pyK/miMW
EasiXUoqlcAHNyPgHV/kxaTHmI0cC4yCThRZ9wsu5fYP34lKszfz/kn0Voy05vleYgHDGkRtzSj8
87evceTakR6P1zWZzPhStQmtbSHkJstV7AFMS4cW6oGso0u42IRAE4wgxFXmFACQ54Ev2Pe2KO3D
1CPmHTJSsx5ZYjveaEexOe44DGNcqY1B4BarmNIOJb2hcs58/Y9FzEZO+0HU8oEq5A5gZE2W8MT4
sCHPrtAsL9A44QFDyvl3anWpfOOMRODgLy/qK7Aq5URvoUfbGVlHdh+XpmnlGdBjqaIxgLLwiCN8
QV/+daRxTg7FfJ/Ehdj/1UUYnkR0XrKfRClNJg6Iv4uRrzrM5gJRMDCViDC+arR5NeVmmiQKcI0Z
G0gLJf0bxHeifyi+7bluo8OBwtNaqP55/vslFsav6h32dAP0325tr/Uahd4ClkTEAHYMVb0exo5L
KL2B72Yvh1kcbBZOk5FrupGOq14ArQbra7y7C3LskkIK6Yepv0p7oArXVFn2Y3EBcbLMBOwD31Gy
3tOL7tgU1OayMGGZPDp0CJV3QRd69VK0J401qYdmHPzsknoILtK/9jdBoGF4CQs98X9O8FuOevzw
O5wNp202AlkG5p16AdF/I66ynALHknxC7M0fsa9Nif0NYbfEm7dJBVo5LmR5rapdjZz4hclHalos
k9HUwf8KDcKYiWtE9c1EPzMNt9G+bJQE/54rsbkYkd1pHguPOBYZYAQ793gbxa1hK2teoa5N+uUA
WoKl3scNeoSwY0Rw67oQBaXDpUvaU2uwy+VWep9iMETU95ou9nq7zZsTcUv419ENHs7pI1hn5dHt
i3fqy8QDkJIcYvVbyuyB+u8o7dYhQo/zAKFxSelFM+8TtriJhRfhioixXQEmv9u5KAIWFwPiX0PU
LmLD6ioF6pfWQ8XIbp1Q8h+sJA28p/BdphPM8I4h0IOxjhhGLPYfFJ8CHRXbChi75U7d51ka0LBu
PWR9dgrYAlxOLDAoW1mZxthwO/SbErfYKlalFkTruFTIVFdcawOAHu1lB5R/nJMwvtRn0vNBET1B
0qy41wjLUGqsd2ngfzwGDMO7rBcEDinDBDJFSXrQvgLlSQ58tBDE8PuRde7fwLu6Ue5ouMRYHbfp
kPFuI/iY8F+mIjuvjacMjgkY19Ocin5ooPJ6YQk1846+00ZGBJ5YtPuClcaH+/dzuZ3Z36zP0KW5
UJ2WbNHD4DZlRg6Fw6NdGxWabUw5RcF3aSk4N0seHcgWF+f7Gq+dasZiUE72x+XS0xGxRT0PIwed
spWwxcvwWkXp4yY8AcA+xLskcRZgYnx/2r8Arz4WdxlJ6IfEogOYrP+PfCw0qrIzxwPtSv/dQTgh
FG7lR7b8yWNLg857/qlesaDD83ULmt4Xvur44PadkxAfYh52qTOCs5d5haiGhn5AlLuigqW1WT0I
gUmuqYNR3whmHZpQEVD4rWK9wjgkTrPEQhLvCi8v4ubfOyFDha1FoVyGpa7PiwZPlvpH2aPs/b+A
i2FvU1b1UqlcrljcAX1BrwSu1fERKuM00w+Sovt8qD2i5oc5AzciGpbLprDXPlGrEN7yXukxX6XD
LlEkd+tSOzFc4NnbVrMSbaI92u0UIKbcBdjApFwkMVlDvzLcczy0rGk61TIenDwvu96zqJlaL/cc
8Gk6oql1xeGON0Iq74UghikQQx0ysB7uVmMOez4i9dic6sEiFRt+A2cwCdaLK53QF81cWlGEm+wh
2P6zgQyg5UcgwzEQe2Kfd5Cn9PeMKPbZ9G3lJnQv9cq1rSksu/8c6TmxrAbdrKvBek5RiM7XySF+
5L7KfoCflt0IFNReGv3sQcDmSYgyUMDwtaiuDujzmI/vwzWomodFaVcp91hs2Nz26kTjTKWQlT8H
Vh2N87j4eAboXs/57sy6EoPwHbeKpTwh50uT8McQntWJ/nSTVPq0AUWmTRQHGdaxEhvT4+6Ij6wA
eb2MAwXxMk2L4O2bVBK1ue9e78Gc+fc0Wc4WeclwuP1u3J/rP5u/F5lMS2xEZopiXn+bfOuuINSp
zjLMp5JRmxD51pSC2a2xX4EIaMyyxfk7/LC4QmJp9YiAZ3NzCaRpMAunTWzPRjbxs+QjdvcBgCTA
24pMO1vcIISBXHxYZNaklqNQrVwUfLDZbG4ZBNvoLt9bs3nEv+U72R7LFLsL159fAw0G3/ybXxdk
mYtpr/yZScKWi3mWhmZVVglLMPLNJiFS4wlSeAomYJ1lYVGgW6CLT9+Up/+YTqQWjx6lGPYi6CC+
JeMAY0BJ0ifrrrb7i2GNhQgcMqjhSlMXCqmYwgVaM72+FHarQHqxWXbw2WRdGW9DTA/sOXHoOnC/
bCs1XUsoGz6s6PylEI1yhyIkNnjlenHq8yuYlUg+5VjvrDzBMleqL9JfCv+BKjDEThV7J6e6H0Ov
8yqoZlmXIWOFH2bdaDmTHEi6vRuWGs7HuFODUpwKuV7HAkwdHNk68aoZYSL6B+2hgotLF+aa0aQC
J5VFPpxS5eXkmFGJQWM1cAh2ek7fqK3tgJ35QNqomHUR2Od3Uqn0Jx+2s6oYNSmyg9n7mHzTHfmo
UWYc5pTYNskEr78d09D9yR4E9X4+l4BfsvpTc/CKkMplIRMDP0iHSXeQlsSMTzvpMyiZtGBCxug/
xkWDpl2DlCIhwpqZHrt6v2UjHIkRSoieQIiwz6dPhQM9f0Deee1Lqr73JuutFMSEkCrpyRuRe2PZ
/rFZ3McQ4VU5FAMcr1Vbb0PhesGBhhIHqSdH6F31/HbJ9/9aVGMqrLlK86jjqp3PDXMbi4ZUTftt
7O+IlL3Gev+wL+P4PU4ogkIXwKt30b0e01n3D1SO7Jd3ZjZHn/CVK2t2S1Or95X+dQ80us0wxCcn
evWty3+4mhkT2gyX/C8Rep8yu9wCCIxGRnM38UiDwS1XIFXC/8zui0Ft8ADaZQOfMy3MdabeZbS/
3RJB9Uaskzpw0cKPMnLtUydsdQY68k3pEdvwvavu1xV28/ltF1LJbEz0W8qZ+pHRPOp+xUmOyaoc
BwqBwsGghN7cwX1qc5w1hkgI51T/cbk/TAly4PSk/m6q3HndwC66m5tXCBTsyXF+ec+R+hFA3Nnr
TLFf0kwiI2oFtE1KpVHUQG1lv4/x7Jj8gOFZzvAEUdS93VrpmZwU5SFmBcLxDDCyR9z7eMM/1lBm
+FAJt7OP4Hj7mwdWK0Xbk1457tLmj+aXL1ihWasz8KBNXlyk5mpL6EACQAWMpWfu0vrbj1MU0Dl/
L/UpcR9gIxF+n21K3ECei+sOovbFYMPDyvjiUzxcZ56u6bltpkXBXyL2eQ2Wj0pqpb7Qw6D17m9j
3TXxkEQ0f4nsxRUwjqDcqBclAzqlmeVsRCmkjIkrzZk6/RZyWOLtTvEpncRqmNo8sXAUr4hbqEk5
rKZzi1nJbBw+GLpTg7lP5HknZQwOecpJFP5IyKPEnc4Y8qDgHdshK5Vp+WDju0DxWYypNAlZVfmA
YS4x4b1APKLiklVr4RGKDkU+zDjxsVvLDJ2cGci1smQXS2GM2rWC+plgoa9hL0YtT+zDsCvdl0vE
+FSWdyjIlhBp/MKwuI4dZJ9C/sFr/iB8f1H/VMCgwTxdqTLe4FxOhBvAfNDZ5YoXr0Ij1r9+fix/
qTGuaeEEfHYQ85jMAi58YjctQrXM9DDqLl2yAntKPWt1zB6Q2EV8gvcpt8D6x1jDhLV2CZl9y8jx
pNxGUcY4SFJFDE6ggiq+msxDwBJdeAXB1hZgLSxqKUhEdsKye7+FobLhbyhemtb/jhXOzPCqosKz
TW6pISj1cPS5R8w76fO+mcrT8CaLpsAKaZnVE4nSXDcLsgsO/A2aA9hxw9VZqYklIezNgT5+/l/0
sKuJPRjORtjB42ij9qaaJVlz3ZCI91GErbGWuiT7mD5xGNXI7y4mLsgzZMnVyfzKQZWPwoqRiiGs
lB/J1HZZCAG4Ia0gxEm7SVHgIrMTT8qOHHkYVFsKnBg6v7lfvcEKAmFRkoghu8LY33ZHp6PG+ZVM
gfwTUDppb0X37mtUIvtKaCuJEhlZy4Z750Tsln845QkRdcgjJsoSa9X9ZrZA7B/1igZNFHuV1Sj7
ekprDpMmaYSvWZwwT0vLtGoRGrcyrQXb4tRYRHVmjXLHapsQBD+CcAhXM/z+jB/31jq0qzVD8rku
8EKLcxb5EuiLnjaSeEqRIlGgANWYskzK6EbtUfWB1BeQlGCrXx3Wj+T3M3xABwhKBt2p+KfmBBXD
d1lAOy1dhLtpWzAE37eU1He4P7g+MkR1vNgGYZe5u4OnYYhZZ04zccqgM5BTFKhMpERXCzEwo0KZ
qzlJAZIl2kOrt79H/iBiQx0HecQyLJOs3O7YXjmrwckTFBzTPGerrP2fvUG8GU4VNmAd0BvNLl51
DV7hGIbiMzcKEl4WWrflxlqSS4lW+NWSfSwAJQKbyHC8uSVO1/FBXq4ipdJQM7tRu7kQAK59Gfye
Twoojlo0ftILmDr564VrcaKEBZzBRZ7jq4SfnL0F0KiGZy4GMNaAsUdZGeyMU6IAfyd3lpORArKI
rPbh3J/kzk8lcvSNlPBVaWZ5SMFnsrERMAZY+T21/u1kPxPBMr3AcnawQTMm/bfDkQyD2XkzshJt
PMlG7sxR3SKVsX0k0HauDvK5NUbSa8AlXhfPESHuoeIk8usNRjEdKrCFfIf8dmtDp4EF4FQ6slr1
Kvd6SQA9IMZgIKtfvmeKfDpMpnEHJdJ90qatII8EPPWYTk2VrT3MpOoSa3CrTk7WSGoSl66rN8jQ
TGQrR1N1LegsdkWTqadJslkzTQQIPzAKWmjp94eGqTswNXY1fN8iR6R0zxvSQTcbCrvSueYeAzPd
AJasQMyoP3PedgjBHOLDUQsHonIg/d2tm13OYNy1ukuXKJy5/27YxedHxbPFSC1tntT8Qq22yhbP
LFaqn3neF7A+Dzq9EBtXDnO28Nms3FHof0P942vH/Q0vsJu9/vLfxg0Y9Q/KUDSSgMUeP/9rI4JM
VD5HOYMnjeYUd2IIzelsvGkKYGfwYKsAAV6FhaeuKmbRgPGRdfFyXmVeQQnFTDh9hNwrQdDyHrJS
P4OwR0mXhQnCBtXXkRyaYJZ14oqcXsXxQf58vvUjDgyx70J4W+yfrX4fVK/UPPTNS3jtVoe2ouGG
7ZN9pWm/anCKWqQYlDVIowtHT9bkcBOJWbiu15iQ5Gy6iD6Qnq8Su+3oGSyHVFJlTTeaZpON0fGZ
ycnFMOM1Zg2FM2dDkN4Z61NYk6icqw1Fx98s22APRD0xGGF40/4lU6f5edfUzP7zku0WNXbT5Ae/
o8RckPqpt+43Xpb5LlDPRbwNkkYoGhroEjja5krXbIVMcP/xX9kPS+e85AZliV8cjh8TVh0oy3WK
erj8L6CSIsx60A1Pbc9gNl1n9B03pCLi0P9znyLsmCT/03eArjsBCBJl/0fi8+KtIpnsdwkiv2wS
XW6g2qaLHqLbO27CSLynDRxXJplZ/s8qizYIIKyH4hK8XwTHX0/EpOw9FF8KfpFj6C03V2WrgucD
qImNDEljp5NaGxrq4PAcjs7RzcC3ApOKIdRkgOWknE+ndKrS7HmA1JjfZattk5qIpeBEdLHF9Y4Y
5zMVlRbH30PwqLrOrM4X/fFVGrUIXcL5bmwBis1ZQ6A2zpKtuR58Uq0LmiuZFIb0ctKmQ+b+2ltA
O9dXHqlS0d5PCdzMBzf9AYPjxW6xOD2mXtKZPuE92WQBM4JEbmfkvvjdyFy6+5xfW8Q2Fzx33nBi
JiRjWyarnC2Pjz82mWigUfSlKsMbWbAb8tVGMbHka4YMLo51IEsst/9HsIfvnflbx5YFOIlMU1JD
PcXYhyckZKtit9+8Zb7VK3R5JE1BQ7OqZ99yRGtAYfEmHzdBLp0vajnXyq9X0dP0aCVE1rLIIpvG
5YA0iKWaSQSau3PA0LyvZAKb9Dr6WG32iT0SlfofhAQoi8EitJp3rqDBJQ+FoNQ7ik44JKQdp3J7
y155D4jj71q8PSR4drE6eY8/nez6cdygFQrFWbWvKJHqQ2Q/LnikvCnZqpE+sCI6IdoincpOInAQ
Rvf77y/GGwZGC9/QhQCxfEvtj4D4v7uw821HLkKiLKlmjhs+XV2MuU52N1qBK48Ciwbo8cS096D6
1l8f9Z1LmxHk4OfIOI3wt2ErHxPyhAQ1c+yCkUSisQf+3LD/jslxX1S5VHdj2ybhETQNU3QoT1Hm
dj2E3Ur7ysI2GwYtEWX9AHowvuy2YsdOb4Hy7f4qsphGHYni16xORNUYvdU8P7i/5ool8E73UWg1
6QUBT4vFIspszbphHKM8twHmZhjHnijk5W8cq6cVwyIlIvZiHKaiHauStbR0eNMdpAaDPAhwHlUr
yluXL/2sEcpCJnnOBOV9erual0UgJZn0BfzkwfNY00ze2WF9IDQSbxfr1PpBBwqXap2izH0fNl1L
7n6HvgLgVf8tY1ITAELycF1Jr9zyNp/ebA7EwWUjvxazfi/Bzv5y424DdmfWBClhojAa5KUHQvRZ
qqH/pxlLoC8xmPvlNmLxwnVmOSaCaOkEK9BBWL+pYCZtqhbaOH62F34SfZOYAtq8U4sB5bQ8D+Or
3ILL28BwQNhSuGyUqbCsDhBm72N44bu336271IhiEV9aWg1EALQhDUgYZsLFT8DMppMvmffA/q/H
RvxIVx10DbmFrMdvMDk4SDRg12GGjDSDI9PN3BhbDYyGjXl5vYaOYD9D5bwpStzMY5LhiT5HkZ33
EiaP9JNN2S+dSMHIfR3xHxfIET2TGa55RFdz568gc4I5Wx2AVD7fE2EOksEVvglCzdZ/0DhmBb5t
3mjtrZdCRizDgKiY/viGdSWdxF7jOKL0nFfQoQOxHq7/R9D9Qs6NNoRsUlxg4eLkjkKe7Et7CHW2
Ubxoj7rl9I+DUhlHahi40uqRbr+WnCX7fKG5GKe1mRSZIRjzWU397oA4kEl+xRvzca1BlWfTdkl2
dTpT6omCAQENzYMY41oEa4OiCbH+c/DBlJp6E0WRwnMzltS4dDdUo/p27O0pCrhI1jluvtKgreDy
Lpa8HW7NZ9rPU1sA3OO1IMJeGlo7dsfvGeY6sPaEq4LAuyh2IZ4NmBMisAVRrgKUy39UTa+gObKb
P5sIf57K+9ZJzER24lZ53ZPwbNEPzaUr1izTJWbJD1ICKwEfSo27IjonS+1p26btLEJ5d+5cgMxw
4k1/lI7ndnnIVLCkBvIh/JmX862X7grGSmxdYLLeBf2ANsT35iq0/bX24uVtkxnerWJj3H1qpBMx
33BtNK+tkCygJzqXOZoRd9zRPaFz8/yZC6N4axj4uvblDHStJC4c9DraRP7TLOio+H6c3mqJ9Ej/
MfyW21zyc4cG3lwsFJD1iPfK8fG2kwFQUe1fi6s0u+KF54nljTgS9WPmWxnXosrab0wSEdAB+xoQ
V137WkBd/QHJofE017Bq8vdkYUr+bpMXS+BgbKtWt6DNfhEZreLXbaOcm/VTJfVz4RHpeiRB0rMA
fQogLVGwStF6bbgqVJkhhHfFFfFxl1/WafsEMnI4j1GjZiCm640qYvyhtJPUZs/xA3hMVRbX+ZUI
y3MwRuD/kPSb3mAjXYMrWx6KBtcR8fXrFPddY0Q5CkXTMJ9+T0zdW8cXn3+PgvMatK3p5srsT4AL
47PEMHn5PzVsUTke9yTz99w0Z/r+ibzDmDOarmpldcxH8vDYlM/4Y5Np0cX7kboSN1mmVQ/Mo3QI
XuAkaQgKSoANVHUcTeBGK+ad0ZxdE/t3AeWi+86diC50OZ3+De9XXFVmedilpfGMlyVXNvxQJdsS
7GSndbTOUyRFcal9/G9KPkoFGQ7dC9pUJjsKsQQQhyk+cqq3wYjXJ9QxHb8AtZlXe3WLIPHhF4we
A5j4vAGN3Wv2ggeDousUA/eXxT/nvIn2PojPypZsePz5vhFp8fccHQrKgiYEQyL7Rese+hUAnNCw
KpFxa2uptAiwdHHf6wB02sqH98RWQaxRjH3mF5rYczbg+rg7cWBXg26yPTq03MVg3WsEzs1Oa9PP
Tt0q4VS2mLShkRwZfc49uSzOF9+xjSYeMt/hJT4xDYN8l8Oty+DiGoLAfKqg3GCEoHV+1MXSN2GF
xkseWt9S6LbUSR6xoeDXRtcXnD2fIEZrC+Po5a2ZOx2z47FsecMu0grXcBVXZ2IkSyJEiLpVnitN
k5nS26Rlo+iI/RMccJbae1PdWyWFurykr+PLBvknJIH5EQFCi4YLtilOgnK5TulYU6szWdeAmWFy
Q5IHopySuILK515GyZ5SqbI8msoHqcAlDc+rK3Qnb71eQrE9WGUmedtCL5/XbjjqGLvG464/wk7p
4ifEzneEFN6sIrCFA0+Qo9mLBYhqHr4n+HmLJUM/eGMvRGtQMZH0nYzAW4+0U+LSP4kGHkVZQULB
1aMX2ysCT9ec/rdioMIrtIu5u0lk86u2uvmpwm5MOhy8LfWYwtJkBcKlqTYA/TcDxyTt6d5dv4qD
6hYJRlzQB64ldRbjBig+HZxc5AMZ31OBoaMbnK0LDVjIUxUL/hZdrqKS1cNiSd5ndBd08q9vV67u
RQ2f1zr7m5tZHyQVk0CbVu2W4YsoseQd1B0wsNIkEQpXduParftiyspTW9b1vlylsUb0dcNlMuv7
IS+U99g/1HNfyiBUENHUL4WiH1e9PZrK6jXlGVsLJ4yHN0fJzp9+SiG/nj5Hi0s8pKoO7ntlBQ7l
9FpdWuKLgjGYhYGBTcrVf0aS50456EQehThgoFU0clK/a6RP7u32rPKw3v7G7aE9yJljYyM5CzUB
5QO8dEvlk9dRNZG4+km87y5kArOkFzuDmnOCyA+TtNstVEBLt2n9g6/VdTS5jw5Zz+F/r/kSp7JJ
EEL9B4Pbade07J45YNCZTzBwl4NSxDqh/WXQW8bv7EELSYkn2w2TnQNz1Ej6GAx/nQThxZXg5nXn
Dqro7ESICXZl5OoJeaFIV2C91cc6LvHnvVLh1tbDAC511D3Fn/rdZzoy58SlCBJQUTQFnIhOMll7
efIxpNxB+kVmVP3NhS7bXBHSVDbbpDviPs9KpZRyhzLjG4F2KpfswqXn5vPrAzGrLRq8LAzXt+rV
5/flZwmETURgmZec2pBCjm2r9+qK21bqbONkb+5Ko+ZoSFM0l2lh36FLA54hvRAcSYbggHVv0Iea
6ATLX1AI+QaHGJhTZnhBMLU7ICrHKILg8y6Y/KsKqaQJSeEimMEKEr6su2xjaLm8AXwBFx05lK2t
OgzX9nIyA1ECB8VW60cRxVGu4BpyIHTiMCQz6gxX5WKvo8DIWKrqoVdazmvRizZqLZfGGMFT4RjE
nIi/+1cLLuldGnGYKBcWyKEE95JBn04yYdOyrCjM28TjsoLMnwAKIwm7fIZwVdnWZ+JDZY2F7Tal
XmcRPskEtLLqW6Fz1e6pLqf/pLPUO7BLdnwxC9I+hpjOnn8DoUEz+sk7n2IJ2UQk47PL4it1kDqG
jcNflzO/D6tGh23BDzKYxtlaOU3Pxrqp0xtV7VW1Sm7R5Pc5McP/FLd4jDJg/0DQuYHOrZI3yjwP
xDn6F/yLHELGO8Fvfh3GYo4Wqiu6ennPMj/XqsH0ZYAVbMsETRORIY6Lvz2gl1K5o5qfAQt15JLf
+hJ+VO7CPklydyqwfLuE+NL63pI4inPWUOJB+6EQ/wzwgeiWr/RzB+vN2O+CBByixcH52w6PN7l2
xYafjxUdlD8sc6T59r6Z9xl3afLs8pLG3t/xBCraxzGgoQ91tY1cD4HcIcJv2o9UIZdTZ9MxfAS1
p0eJfRVzjfq8vHC6z2LBTm6lIEzia429uUfoAb8G1JL4QJX15q0FSDYajey8LiJw5uGiRtLeq1lW
+6BCgr/oIgQCzENKxV0THNC6jwIwzvfwbGltJHJ39OTG62pBOtTS17tQBRoKZV43Xm9Grcc9gyRf
5hpR7h6NUaCT+qXXVs/mZeXL5ih56Ox1oUW/h+0zs0ej3RFNJXCf1Vu5uRh9rIkNoNM319glKnZx
MsIjXm/IxcozXA4+Ngqv/7MZTV6TgQTXeBihghP/98bkg41/hrpXQYenJ4RkvDTlktiDWeyj4RXa
62pB6Zjp7z45LRCM6meuwn7Ukqz7K0/m6NfFJ1N2LNktNWZWWGiHCCvsKQYVuo7qb9LE0CKLF3ku
pHSNHYA7ZIQTzIcZvoB/ES5o5nPUbckZa0snLxecJ+1FeLM3VQ6RCK2xMHWawSha7UlkAg+z0yZb
qPmewQsWJypT7UG/MOqeEkimO/sXxAQYy/wkKYsgk7ds7FkalIkMOn9FPIhNoQMK66311Ohulfd6
F9uj//sIHdHSjDV+GoCx47/MSdkb5sReYjQXMdtTCGqAL+0JS/Hr7GkrYmf1gN+y2cMFFpvTMUto
m3kusI03qoQv5/Sccc84A0STnaAwNR2pT5XFp9r16yFDXrQO4UHv/5t/pJjDM+cjp/mCG4GmEjrN
CIFPQpMzi5Mk0NaCcCFbex7TTQ7LwaKH5cQ2i5BZWku5Nb8M8cgAbyWfsK/nep5uDgJ+uj70wo/d
Zc7bD7l4nrFgvvtzztDJQc8nQ1ibl5uH14/xAGXyJuv6j6vDCFh7KXb+QqlI24RPll5yevRRnduX
8zte9uCa7kf2p8Abr1Zp8IwbFpVruM2g0RuV2fH0eSlc29dOlKXCmvO+LbbnWq4/7GBYkoEMIx/y
4FsvtDOBatGSv6aAWmbtww13/Z+j9touMgipan9GwAkmGwHR3oNUqzIuQf/UqaCnu5Iy1+tGGI2F
heSVwW8yK6dea+IsdXtNJWr8jXOD0CE4G6Kal5w00JepvUnxLB9swerRX+vvyPAcXJt46cAs8nP3
2U+J1mY66rmRPVpBtzi5OjxCmpPaGxJ1y3so38AZ5ex96DmFNs0aQT30lhotcnnylr6RO9g4wwpB
uziUcRq1BlUFK5DXQ/H6sb4540V9xUHqEhyBlAp2BnGYCjOhlr5lQdKGbx64d/YKyCLTQnwfDzAC
hriIgF9gWdhdS1h5a+R/mpinopaEOC1BiThlciN8gAvP2QSkRDGLxX06foJZs93Zn8LZKrsp2Isu
OOwYjqVWV0gk1CoVodhmW2ornkgH2fCEytmigDb+wL6t3TrkmpsQu16uawAfbldVrBGgGtNF1/A/
ZyeAjr3BiLGHZYF/QbGS8uZWQxbkhlYMOdLWx7GQCrvOFHZpirOn/ykao4idxaCZ+gl/Zell3dxq
m66TEeGqwWxV8G2FJihX4YTwWUsXew6bzp0ca4b6t7eVJ32YzLKAJEMGZ+06ZY9QceWBu/+o4sv5
mR/9acq2e8cnzNK8BTnnlpZiH/rf/+wxvvw1Gy50+2M6id1d9lSHZzblxbn9F7hd4upz+xg14yN9
IlW7ihrI2jUr91SB+l7Ao7s2laeMlLoQPyzX9Yofh2rG30q13wr87BtKRv/NrIqQRnCL8V14b+ok
4UGY92uNn9kNb1zBImL5eQmX7Jopy7cWHXTBChutsPxrpE/p4jcSgLFa/Bu6ZXunVLS1YXN5AVDg
mhxIB+HksxenElTQJa2oEYI+76/rcc60LhWxnnBdYU9App3hHjD3aII7gjZD2rPgfIeJ6tkwr5/x
a0N4QjWYeDJdiRTggN9oLh+KgOA5TAPJSXMb3AU6BbXMSM4ucGVcS2z7wakJRll4Jg/X3eW3poWd
LVSdzu7nBqN0SGTwXJh616Y9I2GuYv18p3BVCl3WwystotrwvktxHggmH6pq9BLeqyuI7jpkwzTG
V1C4CNNDbiAFoAtqapyb/9l86qArhG9K6wTIPUFfObb1SCRFuEgJow1+c7rV9MsCMu7YkLhjMQRl
JnmW+PmtFiOx+VoIyxvYc4RzaJwavID4BA7h6LrqViw0CA9B9ZY9J80MVnQoDlOSFdCh2BQqE5a6
ftq6cMT4TZlpCyaR+qcqzzAma1xz+khI6S7rChCh5btT7P9HSNAs+o30Wt3FTig0Pzx8MrHLSyoT
gPYVv7HIHlnPxwg8V+b4exUls2vC3YiUm/6r6LMzx2ztSJJI2AhSPireoZq3F+NdItWw432VPI0j
7nx47Npj2qpW+KEfFVOW7u9LCOGKWrfq+U43KnNv6OItqEspMx45tkVF+R9PlnNL0cmOrZqAhqJn
e0JTHI25WWHU5nA/7EQvDL+uk+sSBClFQAUQwzzCysp5rz9wuSTxSdQ8IL1x25w6OXjGsd8+mjMx
VzZ/lnzFFO2JZ1ihdSgn/3oJrSlRXf+/1IFliWGCSEDwFRoHTNoWnKf34Sfjgpr2MlfvHPi6F93z
Vg/oKQM7JJ8C62HwbqhMNiOV3+cmlo3zdN+d5u21zsZVn+vpg7WSpsLpoLuT+DHhF4Q0h6xCpRjW
+9C0e7Tq5lK4m2UT6RR0caiRxTym6xUECAgREeNv2jH7FH4htMH5WsDaNxxd9RMoggX9u/BMVcOX
5YEChfJh2jvlScqPCrHShKAnGTFyBqQPoK5okvrFE46/Xa1b/UshKNLJQqApLz+AtLemz5RGkVD4
QV7RZiph43iTriGrlBNwrnUN026KzeZUdjaE8YhsNQyoGNPoC8OOmz2ZOmUdSkEBtQ6Gca5FwnI1
58yR0Eno4qEhv+X1mez3cBkjMAG0rAPBNlw0lqBpe6zFD8dbzwFqo7VYiJ9+pTPRKPmfecNk88aH
4sJxQurJSS9kaFtDVe/gXqqskG1rS3srD1bA8KLUoXIELuNlILjscgPOctP/6l8i5N+mNJeTMNri
uQXvECZcbs+fEb1tQZ+f3/MtSjKpqAKpuWfYdrt+N8mmjlaz8v4D7GHzHO5W3boduaJt2FbMBSDa
lbES81CcOzsoiou2bEkknt8GmvcTH9ZqOspKUnhUSs8hMkLkF+XSX94eXDpsN7MLNtopCFOcwp8G
8fCoM7LngsP/Kd6z5/XnV5yOkht3hRZHgCCGo28kazSfoOtrrSBPr+08rIYrtQzK2TLQ3xwUhqFg
YLRMxAB06B23pdPYgSct/1NYnHBFuzqrGTY8zCHHsKBd67beILQklw+b7e3bk9hn4IAUJrHO+ySV
cc3+q9PZ0iTx4GJbxEUJyAzR8Q22TzR/v9Mv8CbbMgUuqYhn/pQCS/E4EpaW4lOYwVdQy6d7w31V
mhKXnoIuRFZwWNH5EcN61R27MV9cnnkm8lYe80QkJyrnuKPIb38iMUd8qx5R97XSk691KWaL3PIo
aHGsvLuH8JARc/l/DmqEvhtyIcdTecY3XxJCjsiNXiYXNA4nazw1PIE0SYWJjXtu+cdhP9V2dDf5
xd+/msigf/X2f2330Y0iEMGgV54ezE6zUoHICbi67uObTtKQ6+iQh2suz0shDTBLyq3fpVvh3sbI
IzYwxEO0BRM5brI6Uh/60iH2J7FCHa/jK221hhVFgGFBSMM71J8ZtECKHcILdbSgajLAIqxNbr3l
tbcRjQMcbLYkILw/LIRriAjodLG7rUNiVZdK4OW75NvMewB0XIz7IGdANiXyCuapk2BmmzGKwNz2
V+KPkNVfN/P+5uEO8hyJ8dUsnd3UnZPHqXBNCyNRgB36oOdm3Y+QnsGTdXCRJSlW/iQZUeqf0gJr
s9tTf+jHzOveqBFVa2fEGYP/4uNXtZJmASdz8Oqg9RtglvNwSvfx6t1aaDgMlbIdNyc73c99420K
A71bDWRNHLTyWbxQBZNcmnLIAYnbb6RpT13bE3dk9bBOftECiE4rHdnnQZ8zRXdk1kkUzhXCS0sr
ogPnNknSFbe1j27qXAaTfLnfZ8T+H4pzhduh7dHudlLDzyUxmd0wOv8we+AR9yu9UeVyjQlVeeu8
sXJeQzDwRgiUl0SlFHW3lUzGFT6WfHOlWBwzMpVfVRBBJTh6Qu+GYnKZWUqXwVZUEvUdIEmP0s5J
izUlpfm8UaxOeXmNYnmhFjjcHngW/MuqbrnJZRWEujG07B0d81cirdkX5B5pbA3wiifeUj51LVSM
+7W8+uwUC/LpQ/ZNHqzowonhVWIqRxAZKt1v+c44U1HA6a10I57MRY/a0o1QMf2NniZFIv1t4/88
w8Ut05WXPxLXOrH2rr90iaL8zmjxoPvT6tLAvm3TmMSl7aasVi8TLZa4Lx+SnQaIox1vmg4vlb81
SzP8ZF+2ltbYX4EBy4nWNzFu6679BSvkeRpJyomnMP6paVsnSD3nv95fEyWztDrAHWcSsM5/3lf9
B7kHWr81Xy1R7F/jfQyTGHyX+kBjPvI5z8GDuq+5GnuMgomo4oA6khbSErO8Q6TKmGNJzQeDlyJX
Jxpl8qpHra4rWUrNNA7ysETfoVAhJ0y6YF6lccG+5834S16dNvxH0/+TqE8uoCzUZ5MS2bjrkK8g
BExl5/x+42MDQFOC3jbj5df7nCKJ5WoMp1mrHyzCanT46Z4SkEAP5YwpOoBI9cAPOVM0D72wG0xe
2ByUca3ie0VamN4qZ+5AUYJbBDq48zy7M+hLfnTKfeCVRPxlKviDm6I1YSi3hgtXkDHoSLVMkWt/
TVL7XPKiIjcCb9OTtOGKMw8u3HscX4i1d9fVMCOQ92uQwBDh3XUw3g8ukvWE07QcAvotdKpCPUXb
QIihrQkwbO0jcgZFk2ligPo+JHosypxoznrMSrC2Mwlx/mLW5rK7IdP0B5v5jkm1mFmlMxOrqFg5
9MQulGm1J5UYEkCv4p5lhOz7KXz9uC2hGZhGFGQGJCY54ZCgry5wXmRpbU1NnZTz7PGRqA1kz9ho
k6iKYF2+/Bt8mAvMwLF1rdZxpbKtgQzcK743CNOvvdAB34nnH2xA9eJNrILCmQ1bJhw2Ghgfb03Z
KvNUpxWDaFTzat72Rp4xvEK1y2GR1Ta70qyxS8VDcQGT+FcwUQ0TIodafwNg2MNOU4f0P7YylPnn
pP+/s93gYVFesb50G9lbkx2wxH7x1Un6NP4GceSu/pwbrH47/exV7YcyGQ/F/QDsW7otKBbF1wHZ
hq/ogVi5pPd2HOWJRBwXz9c4eDsCaE8JuyJt39wYKTQ1YROm9PYBw1itCcjtfYXj7B9i4JxdgsUr
666WMOPczq0mEx6vUGfKNSob/r31maKoCI3noOO1Xn8g5cOeyUfEjTO92ZqF/c+rdYuOYFMWWyig
P+CJsb0zjw9Rn3kVB2LR03Wk30wUcbxW747LUVAyFjxZBZfXhit1LoTcXYD14fUeiSekEjwX8nuw
RUxzYm8oB9y/kZxWZxIzPSH6yPJmAdQGEp1CBrYS8iBoEWVwNYTJz1gPAkM22m16JuPJu2DnoTpM
gD0daLviP7FHKxfhYlCRQBlY/ri7FGGrb9K0RdW0NK4Dz8dpgWIfqUyDh1v2YEuO28DCO8djXEgV
N4l6hUkIhEguJ4OKwMJf49h2Qp7l52BMVjCgmwKocjMd30aw2Cxcdn+g6cLNG/m47RASmXQt+x1g
0024YCayPAqtMEH9GCsgIYMzDe1Jefjzp2o6e0SPLAs1kdAeM8tSaTFRMTfP1Wc5bzqDj1RZkVnt
UqPE5bDTYsGSEGE3AtSrn3ie3gcgK2YrcdL3rzhssJ2bm+PWybIEuDDf5EXxy6y7JzeCCl+4moAZ
6p3QPOPHqkf71eURY2xZ17tJX8lERh2rikzh/Dpg+rhJAnLNx1DR8OFAtVbl4L1usbmWmhFxiJah
ZpL/BmdGJOiGA+5D26iVauPkOeLMpKZZVWfCIraWQPNYpgpj1Y2TfngrcIrLvbSzQZ9YCVpm6Vj+
+efiCqBypynVgCz4Db7x9t4gv/GYupbOhAep7QH7lS4HVS6iNOzakpLwj2vKMm7kNQmdBsx+JYuA
pYM3Y6Mf4+Msc6MxT33iUAAS+RYEb2chgT9xj+CwY/w2zr7pLwmJgI4uX5YSzOjNEq9Na7ZFOVrY
pGIAHecriKsU3y3Eil0M9Uvl9/7pBRmvemPOnyBFu//idJBwdReJHErElshgFrrATz/YgxEsNJPd
mK5SzoKYmDzbR/00u2hHDEUufGtRWkAuoDRslW0qZGQfYjnXUzOirSv9oBpNCbwU6+jUi2GSIgdD
meJKwUrEQEs/79XDEunbnwRx58EUi2HNLc8NI3rkAEAWo6R03CYKQ3XPx4MzdmaVoGgLv56q3lGs
xiYvKB/42Vidu02ECkppALzyJ3gv2FVyDCcnrBq2rgXHPXR8zTYOWNbSw+x7Cf3jGM/ajIPk1Imk
plEV6Z0ajcOOEinJ+lyecg2htS2uftBXqJMiWUeFKj9kOo3KdpWsb38oH9JMRMZunWO2CSVn+X2v
G9iH0rXchC3NBh9ZAx5A/HhMU1FU/S59WM/PP6u+/FKya3GILcZyY85xqcejmVgkyfAcVt5S3ZgL
iMcsEC8D/UE7ft9tXyFiC88yAmoD3UXXYv7+Cl04TjpRab9PbSQ+nBsW+PKt8Ag02sBwdVu55TT7
nILImoJc3nNO/rmHZFOkYJBH6qOMbTDUdzmuKw3w2GqVK0um0vFFKsRfRqvNCPalKN8YjkYY3aQU
Jvx3S2kro7W7PCmJR275uTS34dtmnxR7AolAGei7VInUfacL+2x/a3DZzXDGo6tWMf4Q21jV17pC
vpQyKoE8nKloVD34BEuWa6PtufwBJ8SZQn20Z4Y2b9HiH1AjPWwMR0hLcTYOy3fRhyVLaSziCx0b
4VVMxhPze/c/7G60sTlQpiBWrBeREEAhE3/6AXFOTW5v2oFWHqxTh0FY7uRi44TcoJI21z+R1rlL
/GJ5mvvts1RcbefCAT5R6MKA0m0pcfnOyf8iH57txhhoZeV6f2aOBsg1lL9HK0sZNnCW+GrQIheM
KzJ627SMIRza2/N6AX06Rl5PrMeFI6GVKosk8/1M82x7nLoEDOLc2u5NCa9aG9KY/RySJQaEpSQt
29FATNMhIq58eHEo7ykq/h/qi3zYT0P3K5Q0w0cA1/1ySL/F2Z+7+3l1ZAeRnOwgjnP85T8zVfC3
3k4IYsR7vPlC2wxLt/xGc/iH5bX/vkIj3uwVoQhVx6wdhoGbzJ6eRpMVSih8Wy8BTl/33S31/4Cb
TXcw6uOeCl9+N6qoG7BNWBpPA41gE+ANVmX1Rr6ruOzI9rtYevy5zA8h6W8m740ipOQcj92vcGP3
VjkbyA7vB2sW9EufcBXvGHelnCqhVFLIYPyfmD5KJd7bSSZeMONkNXurCMkw7TdL83fGtXpHwRZ4
rWm9Yabn1OfQGCb9qula4KDpGeeIkLFKlbpcvr6rRFvrmU0RUhC0M80Zjk9Nu/HAD4/cVrIx9Rav
+O3tMDzv/eVVXsr68er1cnZ/OKhDmEhaMKQvpxS3WCiRgFVL5wm1w1uVH3sKx1Iu8ktDK4h4Q7hR
zIFkqoxnmkhAPcgJcUVIQS0z3dNYkCXrgt1H/yZ5C16WA+NtfcLSfngTPrOgnDYqWcHwr4tX8rGy
PsUmEle3iOfcNIkWqHIFkJZ0Gwc/361jdsxULebN4YiIdt1TjIimveeNQ9xYsPeK+LsWeFjN2aa7
2tm6vG8hU0EYX7f85eh0Wr432+PPy7GrrUorZUwZ3hNrWvZ3KypEHqRNBCQPfPrg7fS3Ihbus9a4
yX2Ge7lnb3wF01D5IAFAsQbD/fhnmhnSoF/7YAHwv5tML6/F9NvgPlNqLag1Ryy7FmRNpnLUWwP8
oNRj08KeM2N5sXRc7EJw0YtbHEP/1KorB6MNcxUOq54eZTzk4L2OByRWgJUfyv49y44sEBPcGgnT
EayJKOrONV3NEbWasvV6mdAP1oYXioBQr6E7rVCw9bQGvj61NZLa1Ylkgv8Q34D+bDKayxycLLv5
Jkt5QF+Vt6uD8/Xl23a4VILGVLm/KV8A9izwk2e86vLlztfiGfb6ibDFkwKyXW4vKykDGD3hTgd0
jYCQ4GmKMRzlrO37/iSmGHa5gE7kLO1Iu8w381pdSDhv2NsHgYAiD9LpNsJbe2QjmaUkDT3pp3tN
lO4HiJpCwUyY15wMR9j1UIXuTTyxyCHT3cxQlQ3sTqImDsIyRc+43oMPWjvqLsYUCdz8gO8xCAPE
247WX02a0ehvxfdImE9oVDqtCwBzLqmdvSxsl6ocTw3AHNytikKeSuyWpFLmjzSCiP7i1iQteczD
MZdXpllxhONj0wkAhhJHuzqlTM1OoEw67oMjeV7UYYVV5MWsGEy4JVnOWHQSyoqHeRh3JFGuVJ4A
jPdhUp4iJYU1N7u53HK9x/8NIZBtT4e9jNrSV9rnnp1KGJzGtDSBc0THVHe8kk1+FgR1Bx3EIAS0
ssL3yEXYT/HPZOIVOf5h6y3Il+KFkmw9C/asWLIlU1kwInNBLWeutNdXeWs48mv4TH6CA6816r+n
a9Op+1q5dFJQI9m4CUcX8foGTHU1BHDZxOtZykp3atEUcNCSPhKZUpC7N8yeyZkWTaMy8+CmlQlH
ZoPSsc74mvB9YuNT/WVUO5J7tzAOlD9FzKnGxs5+OpvE3/NQHS/wp2gJtwqXPz7MipNyRv5gQsYc
vviSCfvGAkhaOKYstv+19jQM2Mzw/qxKITJg/WrClrlaIaewwM0ktrRSFQmXLgs1sC3bpb7wOZ6h
a/a5cig4gsI9VPU1FSMdHTXFK73Tv4BCSJhFZWyfCpm75c6q2aXwMj2nGWBV2E6aB3iwypGowM2D
/dP9nCruykTh+Q7TBIT/9oNgGg3c9GXs5XWiQD1GNIFujcQxKDSHp6OqBx2vCWrGZgm1tCzMsrCB
BB4PQ733Y4oWYM8pD7tDaHhxTqnygSNIFXWiOMhQuKSG7sE5zXozXsGZg9AA3Cyd5m1amQXqSOvy
Yy/uhX2O8nZmUbPN2a5hxKz7Vz8dU1qXchthludE58lXnbs3CfRMFKAyIUW+Y9uIU76beT0y30l8
P3cuf39/CNNru2DdZf3RoJGzFNKNKPw79iTxlzogFzo76zjqGEbnNctzmiDCjTJU7HnozBybFWfU
B7xtdHavQk/1elt7xkIlFJwOWTINd29APmHqshx69S/bk5fMRcMvObYx4MDl1St8pp1jev8UHN/T
wGHa3PnVt7OdEtAi9QaGLEuSpn4A1lgvyvlJBmz9llPwgaS83QGQDy4gvrC6CpUkL6sgpDFhEb1T
+3bCJAPp0WDrP1etvVuZrB/hLGWyKrCT3aRw1lYXDjlt/glbL7vaFWcQW9JpMUcRzkLFGHa3ydg5
iuNbLx01fXAVCVGP9mOoZG+XVRpUrNm5lgFs3BpbmbN0bpWGsfDUfxMUQzOhncd/h0dyk0ke9kHa
oMUJvgotJqlMD7Xp5+zP+K2BP+uZe/J5flYk9RyRhIkJms76YrCGe8cENFBCr8KYm/mX6ZKHGbYZ
Z2E5+ar2AJLb+2OdzZZ82jzcUrvz/ElkJErXMmEPR1FJoQmGknOyjlQrVaLe4nfxVxmrnF5kTUHs
FCxROADHD8m5j2gYJGiJWyxaAr0TBACdBHT1eGyNLZr+tyjuNh0xYnWDhs3qAfoWyCvLVK5T4tVO
u7H1nL0wvKfDftDCpc0OQdn5I/VHHAJ7f6hJyODw1sT+JJAIz69Ak//DZmXpp5sV4qrWqy0j34vx
IvJGSxnGd1nN9RlADj2Ye1pV9zX+j4244twK1fCJF9FIDYBMctaQIEHX1plDFVRs5YTCXviqRNrS
RFzf7BSWriGTYFRXwGxut6dA8oJLpNxXv7wmVow8igsJWHb0Nas9x1/H3tmuPLjxNiJs4kKImC0T
AXc3D2LaxJL5vdmrm6lMqmVu5wPJxjk20fdwbVxzNL5YD+2oiEwnRddYc/nae2tBX8v9FWTdwrxu
9w8Zk/4WO70ayBltF795LR8z8gNOp8eso18ZgsBCqV8Sw5R8To4A7QiXaFodlc5gtpMBJ1ZXaYEx
ZoVSz2O4Gan4xJRStlT3BdORPRB1wNfxVWHOjLCTok+lj0tchCwAGQ3WQhIX/Qq6uiR04GICZIEa
bo+pW72oPK+3GwHmj55ViYyBe25FSETbB8uB1EtbpnzOXgo3aT7gvvaU8u22Ps1b8+BTeXNprE13
StUSwkC73tMrS6RxnXyX9t3YvcH2khGp7TwvajktdhSWkhaW7khVzYXroHdBtM/xYhUPfpRWQRNf
kwsArig+Z1dAjRB3228RHXvKFYnKH3QPgYQ1lZpLmo0juEsknCfUvbE5eGsTWyhZv35J7Uc+F+Hz
XdMHcUVVfGu7tfEW28noMcdlHPKrRAPevKSlTQcxWiCKjWMGdWlBYNxihNJLp4xe6DKd+Ru8+dWr
naq0ns0PGrGXJ+0zWcd/cXOmwD3Bgk1fLgUguj48N1wlpvluGlcZQ81I1sZFdToI2aICuYmlBLcR
cUGGsuzNP87P0uRqzTPkqrDb8+sdRVOzKr3uVBERA7za2/OYk5LXSQuDKnyZfpecHdis5rg8BDCt
/VufG8u9iixgET4NazyO/vhO9QUCuDEkHyDYR50TTzJbL2U+USmNP2LwvwedvhGjoAKc32p/Lakq
j6VbJn/IzCE+dZfVk12BmJHS+cMRNQVree5JSKB1rLEXXdRMm7xnxeLHtu1mfn1jl0YRfiyzvVyS
hDck53k29Nht0xadPdIEEdJOtCix6v50GoxcIlHaOes2BiUVh8GtZlTjxutnmcja/PHdfQyFgT95
OR/bYdxUInTCifdybEy0OGtinssdjzAoxAgfrmMAYUqaNHHPkUm16NRreQx6R8Hzrqo7B7mYIixV
fYnGWh9oeS+LM1NP7ngFF/Wref5MuDVGYTM7ZobDEnCmvoQq8imNRPJSNWRJopxszaV91ikQsPNu
AG+/GIPr17tMDgnXbQyP3WgdPKlCRODaRMvVoHS/qL+bAUjUKu6c4JKnBD54MXG26Px07XvIad+T
QeEwQvgNDIso/nm3htW54ST5K2CKbvSXCqKs1kL3iNRe7JwbqN9/yzqB/vxOLtp3aKfPNeYmdcif
FIlHlPfpl5a7MLg8SOEW5Kms8Ev5T+vrGOcQCFAvIn2htJdqwOkT29WH4QmBxvnc97fjqg4cDfs9
uojXpUN/xOeuItqn16J5e5t9xZaF55gy0vjxpOaE+TRsNvfJ/5ZfgyjcFBP1UFCU1/LZR/gIqmyY
jcrDncdRLZQ26xfqJxhwS26IU6qQuVfNqL9NSSMDz+AVhtDfjiwBdXTF3XRMkEG7P/0eNiPEGgPS
WpmlJ44P4JGPEkShWHyu+1Z26iZUdWfwrgGct3oJvv2ZmPK0MpxxJDmD/ZqSEO9WdjVNvJfnInXH
svx1zsweqs1H3b8cx6HQLKqthyxh1YEHFjV+w05h9N+v9IZQBqWTbwHyYN0mT77KbGtiWoZJu0v6
9VbnQL+3R4dPn1JbgGtGYt7W7O3zNNpE6Ip2jpUAZW78PWsKChrvLKiBZS47DlTrH8cqSZ2ndhUQ
ooGb6kTO7u8id6XIxkDuteaOMxOGlLmi4iPKMxVDnxfCFyzZC1Pk+f25EB/dEgDlvPtzdUJRR2r+
DlanzVXqx+W6kIZBwzl7XIQUA6I+xTI3PR2gDwPukHhAXDq+rbYLfXhtI8v2u7Kux637iun4/liN
UwwiWrDgQg3Gud3fbP4bJCX641wOtcX9SFADFUwkpO9NqCLwW9TeHJ7vwLvKHzdkR5eGeFM7cLYF
ltf90AZvHtsHWzsSJ769buTN62Ls4+zvXvrLZrKymdLZUbhURrgmmXodU0ivmJlYvow6HyP6ZfAj
Xwj39isMSKJpqAeGCZKjQgaExnjSo4jTZCW4DyUUsU0LBTbS2GPTszzaCeCI0/KhiiW89BiVNdu5
nYBvahSx1qouXCYPxV/H2ZNca57jocpTg7lx9iFf22tRuGpuxnV3HT6FqTbLEjq3JXqcF6WTlU3z
pM0o8Y1MZqtLPZp+svm8+oqZvyXONcHdtTCRfRji5EgJOQf0KfXXxm0QJiWPJzr0LWzWkWYJqprR
4xPWgRdQmNiI+bKBhxcH2/U6JnXp+49jIBpVPdCpCHqD7qs9qiGdRPWIJ/PfJVzjs92HWMeUXBfs
DU11e8rchuXP1C/M3uY19G3mHLdU1yg/VBqq5n8Ol9tOKNiWsvk+8h3PwNi2/bh2j/Ef5eRCmJAN
3g4qu6D6voOdZvCcHQy8JlanILkT5zVRl/yL4s1HoPOm7e0cZCK/Rke+IqcNEjM9YxFOqDPzfAl8
dv00b7VYUzcJjHhS+cmM703HBCkDiSfXSSCfIL+A0Gthv8hT2dloGVMW6sUkQS7NsyokyG9gUDGd
rg0DJme4Os55l5clkgx8ToEC5JDtFrmRtisRg9MwxkDHc8oHPWDsSayyTxmAvYeJa80X/g+sonrk
T0Pjoi/X22OEW5uYdZBAczp4HtXnOBCkWq4sKSbHK+ORUHw7nnz80GeljVlii7yzwUcvUPCmGehE
FJBTYpSmihUITKd1JG9j91023HWO4WOGX7FWXq6px6swZ8EQ07y4d7n0MH04y56pKdDH4UVTInBO
93MOPoHK9b0+BvvyzCVZy3QJ1i1AXpqEFzgAJA6UAIU7zr5ztb6Wid/ytfgJcHTu53sw7/YTVkgr
s4GkXQ5o2SOgxruz6CyA2nS8f2q/6XuUoDNKgc/xsmWnOFe1vNqZpzJZBElP9+a/tK724jHN9zgW
/feA1Pnhfa4l008j2IV06zyv3Oo404TJtSZJXqEHDFEIFO5RUifbSDAXd63rPgMJVs7nVb0mJ8xb
mbTr0/6JZ4x0Q25v3Q64T/wV7OaYEl12PRUQ1b9zHntASF0vXZfdeAqov66WjiWNPDUMnpZgx19g
CZ4ZzwZ8llHNlzPCd9xjgfkL8MuUb5PuxR88BTLZq5rU5/Kmoop5SrQTUEUHaHUjuoO4B8JL2VBf
Cs2ygc/SaxSs2W3UHYXqS9ZQT47uRRbs37jJBxcasZvqJa9/w8OGM08/X6aRG6T/thY8xeGo0zkn
NLEx2mTYkd4N/4tkfwBGgEIrjcfNMa+zT/7OxdVBp2nGKq0g48oGzuEFCY49JlssZenDJUZEXEfw
fWRC6DYjUOMjhupZ5uJxuPRzcebhI2uLF1Ds//MU+HEdoOg2zz8s20L7hYxtKaQNDrh4PYLYi8ix
zV/Su/csxVpfmpUgryWL0wn5uWXC43/aXw/nDmEJMzvwEf0DH5BM5MrsUbKAbwsQ3e4TSR27lpw2
Gx7n0REkB0N8sj4J7ggygqRmr/rdJyYURX+cLRZv0NqIXhIuWHiVpeWLB20S1fJvBlZw8GU109JF
aT0tR+EsO3+yOE8blRKBvXBpNbWLk63Sd/OG6H/Y/ySHJnUM6pL/LbMwqDJxxJ++dX53/6LVrPOO
GLYtWG73zwk0zA69oRUIXz/naW32x7oDktK7jA4enDagxI5aatIvX6iSkHEN5EggwbSwNF/ebAvG
Nqa5luLNaHxnpbzMI1T0dg8Tf3ABbQLyFqiuTyv6VZPGcgUxiWvEqIpaSN4noYnF52QQ5bvfMaQL
ipmCaSsCgCEbopF6GuyEvwhAQNvUw1wCOJFbE/vKWLnKMsQyWEMUJ1BLwAe72A8iYUtp7+R2Glya
6rz4L0TlDMpdtS0UFSG6wr/wPEcM3zKPYa6+u5N6Ae5M9SISZdPy8wONI+QMrcL0s0gvRj3l5gBL
myHFBIxgFkdy2UCZ53dAl2Ub/gZTEJiu3IcIe4F4vdB8rpCDGSl+dv8Rl5SNf420kmtOpA/aeF6X
zDuRtRAxNy7g/JYC/fhVF0BeuRG3PnUXouu2nFcZ074As1OL6Fwl/d7mysZsGebSzb9fa4fywdGQ
un20j2+KSriGY4vA5GvgGVH//Mey4H2dVqpTcF4F6ySlWynpvZL/9CsxCTg9UYzGydrZBmtjJpui
gfWmwZJOR3uFy5oEt9lfsDZ/3TA02s9YjCzES5EFDlZj9k7Jw//CE7ZUeutXx7lmnG0wOpNK9LGO
LYXKuDCNYjPOIAT5pgEMwAF+G1inEh8wOvXswzcfeASfU+s+9rynnO1Il5ufWkYLenBxsVn58jI0
uqwXALG8k+Ibk6RCMOUTQSLNIjdWGtAwH3aucFtPw68LqFCC+rrYZvv0+0w1VOOMbGzjcsXgeOPR
7tnZh7zbpLCUTWPD0WOyQvOU2h3gp34R4UmlG28J8J6YpY2yea+JC9RDUphLAYAY6I2YcIMS5QxF
3n9Y4I+mxsePWuTOKVWB54HsHeBwKXuCgMt6fFtC0Ad7AB1k3DTzX4eJZLl2dcXmYm3U2qK8xpU7
VQ2HWu79F+355VvrD9Dq2ax1P5ubELOwVn+EfPh+pv0RAe6qRDAYMrm1kEFJlhaSiuN03AwbFoMW
bYZ5ULXFgyw1SzJtJfHGcS7WgpPUow9+Tr3gmQKVnVnG6Ba0hzLLJl5xi15gsJ9lrdkB67LCCFUC
FshUH2dMUb9O+K50/Grk8H4sl5pAqSgWX97kWrw22kxWeeG6fLwi8yxUxK541PcbMLqrO51MKRTQ
Dl8ntody9YWMm+oalPhjLrz7cqRa+IZ39HH2+wA+jGBn58tK8+8qCcFmZHvI+3yGLkbmBu+ybxKq
jZLQ2gmAZQxmE9VL1youqmqM97ylR91xQCI89+XBToIt064hssU+GQoy3ZzmATFt+W+yJui+7WUW
/12LbeGDCrPYR0VyfYpGKtCWZafnWdPYPr8zPVdL0cc0Ua1nzXnEr+YouFJGs/pWBwIlrSEXtCXv
JtD3wdLLdEEv/R2fk0eEVuE1CBYHsMRenGeYqtZYStMTUASZleQgEx7beKUuSBIy6YbxEt0c1Qn2
y2sUcmUSH/OURr/QfwkoOpfH8FKZ316Oi+rB6549ebiRlzsmFP2qDKrjTGJ440K79Wf3N6WOxVm9
ogztwdH7YLz93S4+68hQlGHxOPk58KLEYlvB8H0QHMt7Ln2WXgfwzJsAnwBq/g/mQklNS/Yq3TLk
t5DoatHiEE6JSPmCOY0oAFEh9LKy8kNcczIXugdhtwQOpW+v0UVdkXQ5ww0SzBDXWRV7rJznEXk2
gN47Wmae4PFYIStmBWDmBo0vKRA5vidH6bQlPqVGUtmCfVGlMdMvcK4kzXPBwNgmd8sZC6aRTg4B
WXFgCnVCWlqQZEhspQSEa7E7foonJNIkYzS524+UAfYD9lCmVEvQZtHNFGmhnT9/msd4EJ9vIhaE
m3xouVC0tnfqFJn6A2eYs6lj499SZBDCnd0yBisWMAPBgv1ESj2fFqSze43qY6Js9WOXkf/+9/y5
C8N5vlWVMaDhphGxW5LqC10KoM5we07PwMhSDPT3GnrdgRya6nWC55QjH4zxRNv8qWna1af5fZMv
yToG+p93326pH/m+sTtBmgoHnUMCdgs/0GNlHD2ZiEAcers6U0DQoy73fsySGHB5j/bGxTGzbyae
VPi/bMs7spzRCFuAHLiQnGJweXCBiwvkTYyXsXC9uXyiLOoOhlnxhXkuPKfl+8FBEmk5NOukkqp2
RHeYY9KJIpeZvSpSnJNHX0YUA2fIh0ByvhvpR2h2qwWRIBEqxjnu9ovJuy7yD5B3S58g5lAK/PgL
GsD5E6sQiAiYObTTEqfLf6axQjwZACgfr0Zl+50lcy12L4+JQzVzQPYwqSJ7cBb83RvNmEI6RzYt
qST5HmyPl3BxqWa7iJLeAcUP2OHfH597oaWYgdI9qqLE47Alg4KsrVVd5ke2fFxQtcMaHl8dY89X
+vs2E6VgM9FNc2MFiuyOm9Ez1CT/hajVzzbqAgT6kBCC5uaYPYuxXsMFdKodH92+PjKQqT+p2YQ9
skyRow82An6rkJxmqUrZ8R+D82C39uQSl6Pjb/uPmc+wafMvL6jBChkqHu9ftBPDnSohHADMB3Xw
9uv0sVQj8rAVXGL5eucuf0LQyjji0nMBOPU7bAsNd9pge3vu6g3LCxsXiqkw+cZhQk9GnFmHTX9w
GkqvCRZSxvpaqyEmKLm3GCPG7bNP8TWEGQH4YcoQtf0HFaWhSw9Zct/3j+FuwEPkLUTZhkr88th9
Ve7Nl/KkOfU25ZpfdHfrWK9LEJFlTEpMyDBAV3cktQFMuAXHG777c/AHJit8LvadjewNI61BFcwq
F1JtcghiTQhmyvDsPBRH9VHQoSe3BKGw7frR3zIZ1kihgbgLWj7vHd2t/UoKYLyV8uqXO6dOt3HT
Qu5rX18Oq9gIjT0hXxd3sOAZAX1FN6slr3ip1LMDn2JjI9kumKrM1izbjh0uhd4vAar+EajCiI2x
p+HxESILhzTQTKubDgLRp0exKO7rWshPncj+1PTSL96WMGTf7NTPu/orSClR25iEdA0FCknPgnHp
gr0ucxOl5IKCSgg1Ehykw9DKfpXwW9vCmHAD7fw8AB+0pMsa0F3E9onaq/MFilWylqe/iIftbHl6
FCA86e6L/n9he3hoMSxJvguxGl1nNwSHTpN2A7qBG28jkG8DUdrGwLDbE2MRANI8EWSj6hGkgPF2
31SjE/Ah4yYl08tmx37bsXfAqKDk4q7bOz+IbFZ9/SD4G2MyGJnainwUcK1n7YVh+SM4C/tkulpb
3FDOlHlUHkQoM4/rhPOAzXQkUJVnEf6GqIzkpwJ3Vhu9tEx14xA2hHcWOWEp95vDGE54hHVqDi4F
/vUWIkkqVtXKa5YuR5SSHuhfwCPkNdQYTGMz91QqBSq5HjjP5sRU04gQsIjzGKhk+0GdoYoDFf4z
4SH9xjMPKzz1BjE4SrZRxWJYZvDM28HhB3F4N9aRjYhUxLxFvHaeHFBHafQATh+4P8zIKYYT5OGB
5i67uqLjZqYZzJRaS79q1HJNttY85JVAVBAkfep8XLMstVwF7nq0ApAzQp7zYdV+sXFAVirS0tE2
qLiCrXG+TyH8LE0iLi0dRin7RSllRFo2h/yO4mDZgLSPHqr6CYJ7Dh1voof72u6YElEAJZTbOSgC
qtckRyWAN3xu+7/kPyHb8XiadHk8Ze01OuxU84tr/EZcdwkL5Ht+cWKKlJS7+ve9fUvW1UyhBRu9
Gd3ehN7OxF7Wr4N0uKppxir7t33mMSNQLvtg7L8tuYBUK+iZ4dBY8vdgG+ssJjaRuLgw+u0cuOHr
9pgRdUQ7nB8nNwFhQHs9LLiaEMPl89Q39lSCawmQoVvcBsVgRrW26gr8YLli15ZgWGLGSNYa03E2
WjFLw6hdRT00G74C58JSE0et/R3o1YN2kygR9A5PcHZmLC0OilJeyKY650AzeMLTmQDTH+HrlUeW
SlvJb5nbzilv/Oc+1P2bGQwlQ79ipusKngGT8eNOHHZk1Ig8PBh/8QmR6z9evUtOZhvtXZUfqg36
kHh5x2HmLS/jkYb+t+QOoErAlMLy+wFY5LNsRN4ARFRjTywXlEnb3A3D91pVv2uDktiigpY9ugjM
SO9rfVBL9A7ySbhcNKrC9PgtS2BMDejogKZIfAuxSgi09oStCelUUg3ntDN7Q2JNAf1KCQZWwaR5
J7cmYnQJFWJN2hJ1Xaay+JaPgOCG+R18xhbmgYoxrH3mG1PJXk3Q6zh/tXJi5aG0urwyKq3074yf
b87Juj5J//jcE3eP8xFc1l4b7+H8b2Bz8WseXNNrevnpiUH7PZDD9E9/z3yeXIYK50bGmHesYP/e
K02PUXDMn0hLU5QOAhfBJ9TWBtBfJDDWKtAOFLaTcg8rx1A86LpHlBE+hgE5sYWoPoYgy52+wMvC
xpEWa8Y1pRozs5Tu4YRJoynGfJ4JYQtdGuhOlNaAQiyYanwmWI4cohJ/bEJtEN/2LQUpVj6mBJGc
L3krjzgOC4FLi5tAzey8h34JlWVmjBda3EkGJ1X/yxt404hrJsX3HjJt6JzUoPm/49QNlOIbGz6A
pf2qcWpJZWAAdG0jm1W5j+QLovM7Kpbhu1DInms6dU2SuBrl2Jxlxnc/Y7Wcfm/9TJemMZQ9Q1nf
xTJW3vZvl+wUVxGNq8WYj1vMucMO2nAvvpdmQsBvzp/m/qgvUaXiCxd4vX9GtTkjIcMEIqGhBjNh
vlYl4DJu4LLoyxlcO3KP5r5NkrECaqBhOJvYddDl7Hgy4f7iycadOlII062X79c79otP3sQcVGVp
F5SiH60p4WmOWN/1vtUu10zQGhBcg7FwUacG+armd19PB/OQzoxv4y6XWWKQY0O7xBqY9LaKIpmi
i4AsQ3mgNVHnDSlBcLv4aRAcAlD7lvALGyPTbtaoK50Assu7/pqI2bIjJ3Gd+V4aKrIKqP+qsJpF
HVY7ONn+TT1rOJBdHS5eE6AvrsmUYBrIJaHU0L7VQxR2NslPF1aT55BrjG3vJ8xjF56Z824Ip6eI
5354rNmAfCigvEULdsxAh0SF81R5TG5atwjDWG+Cy+FrU3yR/XSkyRGbeSzp3dO0snAtne7rOCHm
MAcBovCWRffrcaXRZ72/4D8e+EAiRST8nU/yKL5gCbGAyvL1nKhoHDdkgUp7+n+uFvNo0JQBD9wT
OpHrAqhTdS++IKva7NH4KgoqxPxxuupzlfUoDZ0hfkGBTaIP1K5w94U2MeZfgDyFZK9QnKieTb3E
9yV127XoCD6NSXXsM4PLA6lZoymqRMMzmatSDy1hRTtFqF/6bRQijWWmVYCVVqTRgxfAuTobcHe5
AVBKynVlFdvesJIj9bkhgru0wQo7jTblmh4N2req7krvLDMWZCEMmfGN63RP6cMSWmKF3QH1ux61
M2PRJ5H2WxUHUbwnSdFwdOQi2V01FTyibDeQqAvZk8LQfUpNsxi49p8RfGoKzb8RKfdw06A7zM1M
gxdDhc7qoWC7XtO4/FOaOowW4ptLEXC+md+odj2JGdtxYkyQuTOcjEc6yI/Ju9zruAQlwYcjVSmb
6TJX8NKYF8zM2WybkbhAmRN9Pq3Ho8uBLQNhyGqTp602RCkba5xfwPvt1SLf1HQMeHTDwTQYkE8F
w/TYKbwiy4QevDJRlpWfZQGayrqczpHQQOjHjH415Nl9wX/GqBd3N6N9eyii28vL+OkgF79PlYYT
XyvzvYpqJruwDG7YVnIU7nj6tiCQxm7J2rYVFC6gylD3gDh43fX7BdAYkl636zJ9rnkbjG4URVyH
7o9x7NgVBJOb/eI6c8pu/Ho6lWQx7g/bosHI4NK5lp1npKpPOzzpO7L8VCMWhHrvpcCKaNEQqwyZ
jM5snK0wO6z6LWQ5lEr6z+74p82ajrDGUTWsXJ15upi1KheLPLeOGlQkkTOKrt5rK+vjHL1ZP0y1
LQtz7+c5dmJ6kj8/8w575u5qozHL58rmmjea+SpXFgAiPLL0GkcGvRYSkBeJOUEPTB6gRU5hWQ4E
O36Cd/ipFJhBYO6DqdwkGtjdg9WCZ/kN7VM+EjkI0XpilKs/1zf9twdGTau/hq6Ch0ogFXhxdbxR
1q1q2lUqVZ1bma8Ybj7bXeWd7+NW46JEjifoR2ssmATPGW9M/AK58SYjxOovlT3PzW/jrLNHR7F8
lHvGK/uAFy7nWYIzxy0qM7ZbqXu49B55rdrW9IhIM88KNmTBS5wuePToifItZ4pbMaVnLMAFAl9v
JjF+NKgoaDsaRoW4GVksRNhG+CdAgIqovhRt7stA5UeUPCzR56G2XhDKHh5cWTCqy5Go99uDj1kS
hfzeVSGE9sd7coLN32fUJC6xrNd4h2u5HuKIyNp2wb3pXZ6RMApuHP/CIf9RwjpuzfJKi9RiZ/xA
2sng9aX4DPUq1LzP96gS/sHV8544owMrhhykugSKF/POcSNKqMCj44Y7Be7LnDpnNQO9GHl3SNPb
riipxRqYKptRatMJ3pGT0zYRsQncRripvZh7GsUKBcen18+qp41cuzoJph4pmrMvBzlg2DHJazhQ
Ad9VFdnwic6t6NjG4NlX7DPhWOfzpSwG9hwKsWPh5tKl1xYN5ksZnZPD0qsr/Qh7QnmyO/dUB7xl
otyiO26z+OCLSxp9A2oo9+ic0t/SWZwU4x8cyYLu1u645rAaPGskHSm40udvP7FAO46oRdSx8bsy
8sR0SJ2RZo2IgAS3rSHc/8EsCilwFK/rnb+j6xdI/1Wlev8g6lMH02EViZICbbmV5424Eo8VBbAl
UTs1gmT9koxTLO81eL8QkMRnY3vpBtPwntKruJ3rGqkJY2SrCt9Da9UUQjKCV9AY5toI2WfBgKCU
Icdi+657/CHFjLAlZwATiHNksx3hDsk5vZiXsspKXoXN+STZnm3iFQEIVodwzCjKFb7uXbQih3UB
91QR4QwoMpf2yoh2mHqKYyJ2lnO6H0j/MnAS0K6P8d9xsZKxShX5ZpnN3jt9/OsifZypz3vusL8Y
H1TM5PD+I03bibQmCS21/ce2d0/CdRseOpkRH4cqFwy+5tvAnwI1JEJXyt9i6RiZawSGhLT6FjrP
cObcUoQ193/V3ecx+m66lzVh26o9aDTF0glVPmD9zm2B233Dv6hJIbOWyNz9LrVmNQk2IWkp/ctk
R4XvTvriGX0uPEgNzrQSaWtCWP7eResmyYFmo76fO4UE4aTfziQPjgYCyC1adoKvPJAFgHYKp6xE
YIuNIuxSkCJqSCl+Tzrppov/3MNNPvRGN7A/xAjxzu4QLVRmJAqgLaNGLigT6euX0N6VxbYsFDwY
ik4rhiGxw/u7YHnQ/V4X9g9WuLEoURqMa6TYrmCtSbzsu6zyuyTZNNOKr9DrHTvxk9fsm5yz9t8m
oEO4YnMFzVLsDcu38Zj55c1uINzt3CG+1yRprM5pHBi8igAgFJ3zBkB9ASjwhWPKYPYRbSC0t7np
e5YIBb400ZJ1I3T9KNz5AFiuVuRkWsrfDsL9GSMzFiZpUi44bR3VrwL9Flmx3M55/2T0jae6mlDg
q9VeqPEtUpxBmBAYqGy76p6H1lcmDzgdCca21/+KZ5UJUJs08Snx9iikslpUTIfpdvpI7wlrTrgf
HYY5vJgjoBpus4nM4/wX4Mxu88Qs7bN6VAFWvdKlI+7A2n9E1sheQSCLbD5zeqwkm4WPyG+m6iEV
swIWv3RHN4QG1Lsjf/if1outlraYdhkWkQbKe9bwSwxjoYOkH9aSpatI7RmpSZxbZXc2DyoM0kzA
Ed+i5YW8cfQnRwTXQA0MEBdmMuAmWQHXXzGNEO7/4ZI+DLZCmtRzEy0VB+dZX6+39cB8srlRw2fo
XAXYhsevJOlgb+aWL20TukGxkGJObgX717hKyjJj1o3j8UhNUxwCrtfVvcSdAUFr1cwtDarM+xC3
6gwvE3zpFH5Y0Czn62b4Bm8NI7PRP33N8PLXECCrpW8nnMuaRDNhLSAsB4eR809vDUkJEAx3bcET
f+Ffz6MfYJZ1wyt8y2yo1FYd6ryM3dwx6WCt9uXnfUBsvzzc53tnF9IGUuxqD9CH3m/QbP+c3Cmb
sNpJJ49DlVgD13BBQLk3JwfKGXoGmQccp5pwSjDsVH1cdbjH7aIohdrsalfW83p2tC/TERxTxZPp
z2qPFtpODOIag88qpLCSVv2lzHmymPF0p7MFl40mmUrGF98JF/jDkZgKzMvpDX2xSvJShI/I/efg
8Uugi+7WU6GJBkHihVsN/q7tfjo/JYTxtkTn13KJmW7J3RF1m65tC2f8w/p1HfP7TWcbS2KViKyV
WrevmZgG3beKsrJsY3hY3Y5M0V0uNCcaa6f6BM4AnM9PKJ2Q2RsueMBZJN9lptYH/5z+ZIPnakPS
nzkuotStJqOheh/eZPQESTDXpPb7phVyX3O4PTX/LIY/wS80F4qGYn4C4ElPwKgo2WeY0bzqe5mg
93SCW2OMFMTgWFeCDt2bAFeQG2FflkmkwKHLjgR8K5O/atctEu3qN1m3rNi4YdQg0LHNINbyCZX4
F+VaM7rM07nEaB2C5knhOFCpcVoG18qaVYjGglEpxTCFASR15myGw00KCFBIWChg2q/WijLY1dUV
yqyzkr0HvsZB/7ZsWxyaAycUphrnUVQRZWeWbxG3v0vEFzt5hrOKaXPdb4/WllQpDFOWSIlbzRND
NLnt3UT41hdpjMi83famROSsvh8+khEXSM/cOHylvjvoCz4QNH3WgQ7d4lQUU6/PeTwCBg7Jqg+F
8AohYfk+GFvt4IDI3EA7YgDf3OMkYDsNMaXqMS4VZOQtwj0EZXI5ZP31yg7DSsGGdYfLfRftoVpL
hsQFC16IIEusz4ggqqlp8UzgzO5uw+7rlck5OAr+J40muJWpgQxvTkt8MZL6hC7MYaiGOTdvkP6m
DPYWKDaTmU7PZi7n0q0fTvRUcYSu3yeQcbqgJq7YfEgtu+FZ3pJTQg9vCDuWP4ZR9kW2vuWivieY
MSN5UvinmagtV2bH5N1HI2YwdQvkTg5DB5+IjK9pRBiReI5fonM/Q9H1jELsJ03OEoH4UMvSWIcM
7v5O35R2S4qfMwLFHaiqpnSmUbmrEN0l/5NbsreooDqE40Y5q5/kDXKEFjgLW7XaGrCqEWO5Jh9Y
wLWC0/tqGwHvKXm9+HV/PPTNWZJxqbdCs3a0yIiCqbNz5avAVq1+WWYP1i0nQ0fU/wcCTaef4rN3
YIKCke2E/CVs0D2b5E1t4lnOjKL5oVgEmQenbzlbl/z5ukUZylnf8vyGaqDVcn6Z4uW9etocSbCJ
8EgEz3OBS8Erth/iWGlJILvVFiaEpFnAuZt+5RhPCag8jPUso2UFWLJcn1FA34rHluIiSsY57gBm
eOY+SZyyN9wwadZu96ES2GPBTioAGcHXl4xAwpAePby9thjiq5SjUUNgsD6+nCZQ1QRxVW1tN/vf
uClv0dO9Xmi8aat06/Vb5GDioIfX6RBsYO1kzLBt5Dx+3fA+RuSsu7Eo9BQ4IfFx3Uv10zu40AOM
T8MOOE8ld6ahDRjIeChS3mnUQP1Djipjvfa+3UaaWvx4zH+bUXvN08DJMni9+Bw0UUDpYYvVga+I
mWSEmGAdvzStYYVdzaRmKtCzW8D9SR8/kw53tDYgRerBnyrOIzL4W+rprwwDOY7g2jhv+aBZ2xSd
kGn2Sq2b8P0MHg20uBRYHeVFA/cbC95oabAiRY7WKQxgtSlT7CGJaLkOvZIAjKYTix26jzT9fCTx
aK0TOABCP/vYkQ7iqzi0REobSYqWFQujJ4TANEp9E6WqLXzZ753o7FjdmwdSfazoWxnk12AkOQzf
315Hi0imNTVJsJTtih+DnTQtaOmcRh5CJmlPBBycLq4XpbTTBp22K7ulFfOZDZsOt8gJnlElBtHf
rQCNGCWe+abXH+yF9uNPIsPgdCA8cUZF9LTun4ef8hr+6c7s3yGPYS8bR7ZgoGQ/v72swjrxwrU1
lk2s3cXMzkI+CKyKggxcJiBH1EPmOAylsgOZJNk9/H6MkBhp9kbYoPPNTqmw9mM7tsIH5LVE6RmL
Rgi4afvfdA36xlyX2EmtinDK5jC5KTPf7zekcv36XDvdvNT5pXDhckUx6nafB6qU4SPk65SMF8q6
nLBA9UJsnI0wTf5J4zdVDWwV3/gq0TNBijrQbjk+DQwSzIUH4tAQHU05/BbEqqHCyjy8szIZgpDr
iq9e/XD47Wb0uagaC5GdVqJUH9YkYNIoOugc++86EJ4R1b/uiQ0O0LKJFmY6klzm8KQbYRZgJm1K
HhsLpHN3LbdHYulfduUbpYQDXY0b2TI+wLYqwkUIwQsBXFb6XLy4Ba+pr8DzmSZZ3drSC/ojNwPN
TzOduNZkrTx5NXFWhFwp4T2cEW9Wb/3NwGXb6eU8KMRtUXiOtzsIpPvUMiHeQqOzCMKLGOchirMd
o13SX8QgWHodrS2RMLC3/xSy/wEpOnbSc6sBE68kA9x30/oMW1pOS++MGfubHRW7o3n2KE60zQem
78TmhyGRE2DTVRl+uzluZwf33mX5Bh02Efe9VmSOjO3Xch5jfwhg9G52qpMxiJ0/TnYW9Vnj25fT
Rvo8DDsOsiEud9Ss5dCnOygNJ/G6zTw58t0WkrGgAxDCipNRLWpYnxy7sm2QVMAWXuciuJvxtoLR
gqnN43TsGM8o/RNsv0lYeW7m4GcBV3pyWsXl9UIZ6oqIyXtGvctjT3H4Lv8lzQ8sEAyImgTn+cSa
foMpWBsk531v/7HoaUJDKQGqHY3kNr+DBrTFUaB8KnjnN5+7hqJEI5kAXCJN0z4z+DPnEL9wSWne
3uQnGwnpaKrMxlX4Ay2KKyLXzmQFP/2biPHesOwwiqJNnRNZ0aUdIv+BzqANMIHVFOpZ+tRtLr4K
ENLbkFXe5L7JVOhWFCMT/6F2nuf8Rho+n6MfC0pdNZEDQGxZejnRZL3k56HDOum2qPANHVuSl51G
2oL2Zj+GEtHYrCeVO+Ac7V1xdKFTiCeFwQxjOXezY2MBwEVx0g7LcZ8HvB8WquA5K6C6H5tt3La5
R8unToPLTPhpUMs4PVzjOHvssJ33Dd+NRb/d0xkK0Z2/H0KzkVZUkg/QgQMpVr6bHjeJcSZEvT/I
Dqqt+5o4PTTfXO/4ZRh+8rEFg/HkyIZ7p9oy7Ry0XsV63N/ZOQ4ernMa938L86PbCl7XYgS9cVr/
5TUA8ZW6idBP+iCjLISh/qkXRsRHJ3g5zT0eyg8an6q1XqOcWxhqX/xAdwbReD+dv1+dWFCUW/f2
05cKhZg8pMRaIui02EF0GJXUP0kWXqqoVjQS/bbRZA2tTKafciBlKDUOpELfbPtAcMbf+exk3I/u
5nppa9IR0xymnrewvddCU4Wjj0TnTPzxXu9GvnsGJ15vQ6dKHZX5XOraKOcqG5QFiOoZnlCY6crK
IFVUMvlukWC3XRLJzxDTNly1n4glmOx6Y8+CzaO8vv9OgkasWeKg5USriu6kFW/Tjz6qMZTEqqKf
gKxm9mt7HZaUoxUr+DGOLr2p8ypMJSzyrXbtcFxdAfzx5u8Ql5rFONGpGvMFe0UoMlFxMPtLeZcp
09uilHoNCgZSfGLjvfp9EKnPRjIh39wMVpTGuN5PNXXr7ks25+FmDLnEo9e80mooNTZaYQwB14vU
o20DgaM8i2xI1J0jwag6YBkvTu+FZq3R398P/wWihw66zahYrYWxDOfnFAZ2NWY7z1ciPRfDE65H
taE9473Uw9vJ+RLK370ki7YmibA5J4GwWuQ0rkHbNX8OBZ6I4ImM6PRhXQjR552dMHasRoa6Mq2E
7uRsaip8P60FeA2oe1fidvUrgAE+SOY03SElC1NJmdDnbXnKeAkrHgCg7u2EUIaiG5cmfSthXSVu
LcLiH+KPnaTQKz/BhsacmbMFw+ExrjYDA1lOx1vnDBvA7lXT52v/li5IXhkbpcQs6v7lmn4DTRYt
J2YznP4DDALPFKx9+UTiQRueuNjrneTeJr9Q4yAleZdgyipavG+MdQPSiJA7/dm3xkvtx6uIVUzg
IUnSWk7ZNiOa+wwATq2U9yaPfI5Hmccwu2Ttx78TJ1mlJSgN2JFiVmNdpy9LRFmAaiU36D8Th0Sm
1RXWy9P/rNrrtZ0B6h+6Tq43/z5EHWQBkt+4h1pz6MS6x9iNrc/RB/HaQmnULUd5RXKDOvgyEsl1
bvOoHrqArdIPxHaHcl8yrosqwwBwQagztNIOa3AhQOhVblEoqApiK4oMMfjZ8Mr1IEN+rMXaqr6K
qHT7C+gPmob4b1hCm4z5QivC9hm6tZyeiynRa8rhQhGKb9mQBONALS1As3nEwRlZ6pdkrTeR7QGQ
H1YaPAFEVt3N2Px3O4xsaPQxBXxea3jLHz5gg/ZnFiUnraSr3wAQ1UNSfW3JfjIitboDr9fYms2h
K+hR0eT25Y7lHK8UwD7hkLN9N5697H7CarDodbS5FFj7kxd7GBadOInOIwOFYAYKd/7bjbqjT416
STQ4oEC6SS59wlDHuNZ+3RWkhHzydA+S4iV0nMy2dAQKitm5Gx+hWphqdfty9Vc4T9xTj3fIZ0TV
YaQ2NLzDuTjFO85shLxP1cg1Ry2cThFsWV/E6ABAwOJfWD6ue+zrNvuV4NH0lb1fJiXq+iSQjOCb
nazA4SFWoo0N8Zvb2zIX3ArplmYyUC0m3F2Pu8Q1YDrQJWExCGFp5dY4RzHGjfO2klGEnpiBZwGe
GPht6FWiFB8RKUHvjMwpgZsqlMDHYkrcKpEQUGSuikXG30hwODGAOExx5z+pXJ8ytd4AwM1+AEgN
MbfS6R/BEPwRN4N8ol6g3TO6DOe3GQ/1eC90t3Twp03RnT7Jkl1rk9eM/YGYhkz0iRM1yYWhp9+L
IBudebvDpkBrRNTpbrxdddigXOq83zVOxCM6N1/+tM2xP2x2Z7Wqt8GenoHqAwtfEYYo6Lrgf0Et
P5fYYRzT9FFcltcZdRBPhNjPfOiaDAH4AbIGDpciOa4opHuQJwMyEKLsKTpMMxJn0l/liTyxQvYn
uFcqoVUK+jP5bqXFvFe6HsE8hZ7GHaa4gpwgPxfFSGnBH1OYZNrwhTqt0+bARIAzAecG94xEj/Y6
6UOSdKoqd+3lKA4N1qbjgNzeyk/UGhhLvZ9o67hKnI0rfX/d2Ji6LCJyJxrg03o5gqydhrep/8cx
Vpwi5Gnd8RouVAzu9I7LBASYUVklnN17PgPjwC2iIy55QyjYXuE6LO5T5QCW1C8+xb7QMmiBznXf
RhCZZd14/yWIv3ajc4hseZ+lK1/J9cGV4ogXOlXq4vATzGkmT2y+1ogEy+BZsoHujmSRk17jjEFT
9ARB64UfdiMakIGjCQ7AB1K73MivCJPm3Xia1TW1H0/+pMJlBwBB72J0OUVnBpvF6QRxpRAHTwvv
ojY4SM7bdWGiHNoByCsbmpGkGyr5QeqbL3xB4h76UNAP08OXnR5R8iL92u7tr1IJ7gQOioOqgIGN
7qtYoU9fEDkN8yNxogYBjQ2+NCde7NJErEXg7v2n0eT8aA3wykCEGo8nyVXvbeGv7Mnry7WASikx
sbBOIHZNn0/dy8Cna+li/GP46G1JKe9dLXIxOr+I9Zu2s0wX7f6xrKusUNief1Wfri+zdRBoT0Le
IFDNoeTBgch2h0UEelpTogr8crpHuztZ6EHYaxSxtSacjGU4eYZlr/Xei0dh/2yQXpp1YDU/HwIJ
DeTCpJ0hNocgMOc48uOB9TdwQQS0a1hvSSdJIScI0YHMR7tRKyh2HbT5SPdf/mTbmIV7Ob/v7VLv
pqA9GYqrDunVMCZi3WNX3XLHRj3R/cmR9IsOZtGIbC+7Is541QtjcQFAFvNaUSzJcrGr9L0rF9qW
GOZ+mEgC3xYTu1JU3+33VVhCnr2cb2E1ZNFWHjKZYPntRqQhcSOv8Pt5QKYnQ2gssrK84+eOhdwH
bHbnGyuRFPHSV/N8D4YaaX6KO40R/oOFlwBM7m1whPyI/uXYKcK3HcySGADkvWXNBUtC9j+f9RB/
osyWYA/FKzhYXtCZJLp1+0AHY69gMRCklMifsixoXCOA5+bDRC4GQCZKTlXAEUyP3y3m49Z1Jnhh
vLJUZaeq3xNC6V9nbs3nKidGsPvj7uEujnQp4VdD/mj0tvhYemjnHNqnnXUy7hRaAE+wUzds1RJO
MoLPhFsqBe+RH6O46deiK/PhpmflfHgXzhX6qxLiLPvSOhZFJnPz3Edwq1Hq7qRTC2c0ox1fdP81
96qJDaKw6EJyQ8uvBS79l5KFvn/cNs87Kq4PlwbGa7DDbs6wsq+MgQ5EGmNgokuVN09riWRpxHVS
gqbtozI5+abKWvTyJ21n+NbyKmkF/NqA/FwSxmMmCtI52y6eswObEkEm7kYe8vTKz4nq77Vliuk3
eMOZm1/uVTykBx6Nr2FhwUZeNgcql6D8zEZelevsaHCmSLb+TCkYF3PHZxYGeq92E3KcJH01vi+7
uP+4KB47AQEL+cqi/XrnkhRsAf2pHU/nO7Eoo+vNPM51fY7/j/f5+fWkdF/98rNlLkbAcGwkr/a5
Pk2XMNfAn3MCL4DVia1az+Tf1+CQASfllxcxT6b4VuNQz3GtuH9yKLw66+bZwbWouxc9aL/veprj
vhXUEuWjfZwRat2Feesb7rcA+pm3hAx2BUl3P9soekUDzxWzw43nKh6i3iHb7QInGFNid4gGou3i
1YS9C5KCfxA6vS2F896FDY1Cqb+YdIEy+1KAaF5TrKvYywy102i/UPR3gAST3YqX/0W9vrt2xI2H
npJf2FmI/U9gqXZ6Ttzt+IV22tiBeuv1PYkfvjLEQDXGbRicI60sB3HoVGJMlR7EJTcNxVyv8lQY
kMbAMTjuhiO/DftlDNnGmOhtuSdOo+YlINxAarfbi1t1FuDjx/77JlqsMGTknKoZmYrjU+YAzM/a
yI6ettl9bbgbOdTJy6mMmKAs5pmKS5ap5CBr9kA0mNo23m2Wo5YrDfpzAWIbnGXFc+OkO+uKKjrw
l5GvKtkkOmsByJHJs1VpS8lAmqUAviW625d/SfGIH9U+EP7hMnxawitS4YmCT3N55kASOAQ5VJo+
CW6G/Q958qsMV/DV3DJPOklTxUDrBj1JaBa5/P1Y5wmNoHw5SoGYnJhSfZjcg41/nWcH06trnxPW
mEeG43bL6JzAhizglWXaNSVTr4mF0YhC6ksogiUGz+juU8LiB0O3SVzctZNB/lLdoZ+Mxf1uhuJC
dRx5DcsHba+X6JwBTJ8AViB4dVOwDD/a5dohfziVbzH23EHgo0YtoHKgUoxRNjVsGgtXv6M7zyjb
QeXBI5ohLOtmkQFzGps6x0dP8OrwCq07MWOGf6SIZfn0Kw8KFJ+Ci+OVXsenNP9aSGyJdwvO04z5
Y5UhhKTgH3gm0mrNO85XlN5ecs/d7J3/omOlSo6fMjls0/km/PZuCE6otjZI7iZoOe1YCeYVNvEr
4JRnQzzC6kCh4JExIMR3CEyulCGDyjpgHx/QqoNhtW2lJorFoTiE3+eJw+6zXoTKoHU5GMYmkXXK
CCXtIIw1gAGMEGPdYWbsQI/IZ0AKYzrR5l8Kgju2JauCLOrarr3knBmcwBuwTxxhZKNUhdeqq2aV
rmkqEcfCRoLZCug3/KSOkd39TmAO5eFpv38zdi7xWWJGl01RPkPmUxDuW5RcUqGveylC1ExfRbBm
wWVQrb07omNKA59yKPV5p+6k8uVxYS48BDHgh5LpYonkQyxY9Y3FPrifCWOW32Ry2dDrpSx0Gv64
txpqZFWvQ0Uzq4jPHfHVN+qBZFOLxFNDQEkWa6Jcw+v2X1pzwtzCLhwBx9J+EoFHR2lmaBMROaHy
0EDkAj3fsbgIst7rFlk6t+hNI3p+E0BfucyjJg1pi5FKHJr+Kp2OOMLwtWlicQ8uxaLSMa57H/Dv
AK0eerlDdT35+uwiu8yG9eCfgyD6IgVpMaKNrVVXHrTpLWRFutezj9OTCj0oRNrSt6Ofo/fpNni9
H2Zv6KHlk6rli1BnPET30kgKeB/mTy6kmGRlz550RooFOaVBU5NoigZy9qC6YpNi/eVD3E6ZzqPA
IeDV2NdMHonWYAHihcExFqTqdNsXWtDgZPeV5V1zYYg1CYIu5pVGgSTFgIl/4JWn0Zb2xXDfxbUQ
1dOmY8ZZLka7seu/SqlGKjcRxJ0LcnSaXW3bjFk22boe0k4iEt4BqXjm5gTMFYE+Lr3cYck8UOMK
AEdrhblJ8a0pdrb88LHZnVWzb/NpG0HaTojRPvdSIM39XOxmxMwVLNmQz/E9PlF51xI0FDbPoC7d
1yidVXcwXAaRkny3/0qgbR56YacPGqByjHKvOuSwRE+VT2X0WKai4IS8xfXCjrR+WGx1ALxw3Hrz
SswOsJVH/ggI9X717mYQFpbd0nW45TlApc6wVDA6DEQkxJ67+r21v16ZNSPHCZyuunC/evpqvATL
YJFWfABHODbOACXgnAaVX9W4fd4/sz3hQwfsZc0+KI3YUpvglmk6C+sTpD0anJfrDb65o9qSkZ3U
q+yLN5McfgjXIC+J61mpfE3VtfQ+kS5U5IG9qvAbjuCdwVLBymY75dYuU6O3/WuFXVqEeZJn8n0Q
1qUOLdcUhYnfz3YRn6XK+1IFulj8tafwN8o7WTTizAQu7Z/XKuLPhWcrnYjsYFYoRIAzl8oFFdoK
7A7ScO9jrVjHQV5UNwGGp9sLcqg8XYeYkXEgKSQJbnvLjCJ/i4roXTB6S3u/WyWAlpTeqANH3hQS
8eop2uiTsnUa288rsoCmEkoA5yXYG2Myrgao6cxfK3uh0cJE0vLWP1MRLL2x5V5uiYIYSdivstpp
WRI8hR4TuFGN0u0++rY3HiO5SD/T3AAHlEyYTOFVSjZRwPCo+mQ3FawaMJEM4cgbUX0z4a2aIuqy
x7AafcOnqc1NW7wnCS9lamJiF8Wk7KbiIqrg06wHQVuuw4wG9OmmGL6xZnX3SNy4roF0vJUEEDxJ
GGtpM1i0I7RdD3H5mXsgpcJ+V7eLNBYvAfvDHSfOdPvmdRnMi11n1xXsV6X2l9WEbYPVOIbhgjWS
8/mBRwMHCQ0TP6Gz+QdocNWf08gfnPzDsFS8vVs+EUhmOHnpTXqizg/96mAJHGhLou2/nkWttq48
q4jMSRW8nZ8ZmTHFCtdGMDk9tVFmdB32s2d1nkHYSWCSIt0jYWJsufNa4V4QTV3DgYZRs8McOWdl
Xr/LONXnxQYfImg53UhxkXsBr8k6C2xoB1XKJ4eUkKIOCI2dd0ld/WXhR4NvOtQkv8p7B6Y6j8g3
ReCN1xG12d/VM4dgjftbUGpZ7eFSajlpJactJh30Oej11YdSpMHg1wtFevyldB5OMmtIIfJXhNP/
MNw11PpXisQexLpndc1vXZZPx2CNYRJbGwJDymja+sSawq67ssIc2Heb6MMM15J5WdVW7Y4X2PAv
EAwCy3ThGeiHqe4aFX6eGrJaeHAqb+TW3h/avsLKZ4BVotwz9eK8uLuHOSrBSTx2TBSG1h2AIY5m
0Ocw/vTdGPCfKONqIP6psY/AnnsAbYtAkmU/Vyi/7eueAP9W0RWN1/pFcQsmJHVdrw59bmqn6BG6
lXOa2dbhkyDhSFQVit6cjh6bWHa6vjD9t7zSbgu3Qo8HN24c3UB6y38PE4mFah7g4Ay2fq4vP2JI
RLERiPDyl4amaCSZEqHS7ei49X8+ZWd4WAlhpgu3A9PJ+v6zJObQiLcyUO2DDemPpKCkN8qoWEFl
Y82nxF6rUijLfB+7GK1lW1N34DAgGcNLK0JhIy5Vn3hiJDd7RKvnrtFmT5pXjT6wDfyX/OIZ5cQJ
WduA5kDVwd3vqcd9i/J3MIPtPuHibyE4pWDV/YnH+AhBdkMOW2C6evr7WYFR6vbhGW3I/zf293sh
TX+q34bzm0AowGoVrWGDIpLycJTIoW24vqw7wOA+EosrdPm6wfBoRGRjlUKs5i+LPHKH4vSeO+xf
CtwFlsD85ArBt6c/LdIVLbWqEV+Yf0sxlO90Vx9dhgyAp/Fy04QtrPUXee9lc9hEfnHOKd2ytcMw
fA0kfq0ETLA9SG1i3itg6aXzE66UAhz2++dI8LDVWribxSRBYGf6TGTqco65sVvqXnRU8gONpeiV
S88sZSFGWBiDz5CJrsqi725qZ7xcmMJvQ2t/QJNIGFIi+VvllFD9OdIORdWOSsc0nt2HCViJv8w8
jZQQXFbwbHLnuEB9WSr3WgZlDCkUFfSSHD7bl73LjA20YE6anyt7AFs1CX6T+cjc8X2sNNuZaX4m
5qgf4XEHSJCXvHc6pllYwXYn7gQ+M1nLpmY642rLRkQ0/kXcft46qIq3yjTZz/Dvsxh236sUrBGP
F3MXwOOthh6g9rkMB6YFSi/HX1buXMRdfKhc5hr64Ma9vbzqGy3PZM1HUaPg0kWh+vTURcwv5X9s
h6890j+yKcRwVbEX+26aKguLunmfOMC6JMFdA9EeHgSRiE8xL0ovjHEmKbtkUs8F735mPfZIGew2
FqIWunDq2sD4gLSCj6T60Rkwi1tKapiwQaV5sB01FapSjEx+SX0XPORrSKp+oHqge+rf2CK7n7HP
NHvWykygN9/I3MSsrWm9fl1dDUwh/6QqOcpwKekvxIqv09KFBE91T8r6o1+pTUXOb3ghyDGZts4L
HgUxw3MNh+qTB//WeTKKMaRfVKMjwlL0eeV8URbSi2OovpIWb1tlV1G6EaVcPMGmgl5LEw8cdjmg
+hdMFakAUl/8/1ArIb+daZu4zNmOx+E7jxIR9RUUK8NfVgFnD5h3xKDQz/446a0ZHsvoL/huOpCJ
szBRSJ9HCQfW5SPZBQdAUxGPXgiYU3NyoCzjQwL1+P9opd2+f/qt9vonM2XhRTA2Zi1hcz9o1fGi
C82l02jtQxOkPOupPBSoo1YDh9qvfWx8If8qJDQK4rQuzS6zvszSDyv1fGhRjlocmLDNeEtfwmFQ
dfTI/OPk2rug5pL70r2YueMzfxJuPT361TMftflbqlVQpULZczER1COWvmT6FaMcJnQO2RvE+G17
6ms9B3N9g+2dPzThJJfF/rgyq365ppphIhekXAsMawlzsS1wMn1pS4ttC6zVkYepnNmUnLovPkx0
4VKg6zEoE0O2+4tgzvGjdPM1y7EQVpspD1AMLtFNRMmPR3+lHRNme4uKx68YFM2Cibvmapw+suy4
Gd+r2dVcH0nhpAUYoVoNq2VaPC6nKbh7ZB6+BiIWDXAxlYa+eix9FwKE04hwoe5Ne5spdm+IEqAF
ennMOO9wdywjOC0+GQthyxEXxT9orxjcXcEKAPFWvicxuur0LBvsXXiMtMGTmjrrxaYDdmaoU1yQ
X1jrH0iZWMwFDa1uGI4LpzP8gpA5Dnet9pqePj3M7HwhFq5WKHQhYEtUXij9vsCvaQzf99QfyN6d
dwvZ1AGiab3rtEIrR34oqKB5y53jUc1rETVsGzMLVVQ3DroVX8q/EHePD2V+rUwCtrj1Kah5azHi
smeU+hgvmr2LL6f5a6th5X1J8gnNuMGVVq4Y7gAiYYZhGvH52geZQ5Ey19oZ/aC0sqwoGbstwtBl
D8l1N/Ja+fqVrvLaPc2vudg2JcIlX9/ZmrtXtN/zeCn9yaOyV6RNmg/YCEb00bnoRze0Xxf+9i60
4VrOp+llV2hp4JUUp6PwulQrCG/uRozPeRg7rm2DNusG/aF3DS+maFjY0RX22cs/kinIGCEzlVTT
13yoQ9J6Kd+yO38N51B9H4lPndhZJzj/x1yFiHN8cgUUpA+Aih/Yxj0W2MI1U6NCLmkqLuBq0+Zy
Or5pNu52Y6NFMyNTZgjUUtnQ8kF1aJg00wKpuS/++Zn9tzY5PhOaKZpzsidd/fzHxVfrEh2oi/hO
HtnlrIyHSz7egct81H1fCtMoTfmyyBV01gLigZPCRC59uAK1r/h+cbLnC65fWIge5S+1GVUxwijK
2l/30DjiQezQWjZerXzR3ESdtJfyvsTcV8rscXnNIzSAhGCcyQJwmNHT3pMiNf+WJh558dq8Eq13
57UPwVL/XxzjhSnRcbkT+6PEhkIVc2aNFtlOX25vlq+kvgK0voc+WLtlo/QqICo+mDhOnWN5MtvG
6M/wSwfDYfpzbV5tVJIc4LCXJGDArNQnOhqazq3//H9/UIyrQzOw4p4diUud+TmXwrTSJcQ3CXYq
xht5/comL/vgIKvc3/BoZ8n02fvOXb4n4Q7O2r+7lmbh77bO6YBy6o5XujxH1AXHOLXwvBZ2FY0Y
DWRoQif1ybyWbwRZg4Sq1rUlBf+E4geZ5x9qMC54DlTT+B1KdprOYAKnGBdrQgHpxEzv4K5lPr7q
JMt9fhzdcV2SJeFekhNzrZVAS5v6O2XDHjXuSCQ0A/YH8PuAueXmkyraoM+M69jIIXuuFbqnz/os
Jk90s2CkOE+btupZ5IpN4Z2OZfmrt/PTLX3LypiudviIcD4bVNzaHwUG6r81GyBc+NT0cCvIQDDS
eFIgzseBIXUxWgpYi9VFFpX0Q0qzg2PkgFRwlHU0QX7IwnzfWisswkARK1hshQpCHcU8HZpR81Zr
JGVCvbvhl5UqeozSal8joAPReix2c8sJ4Wj6k80v3oRVPz+VEDn9hTa+BV4ExBtJyRWXpA8YBrIj
irJ+YHjT1bQYSuHUr3Sw/ZySxv4IEfkfuEaTJDGaPJNMG1VlfwHB5PHUnvpPlYuCfoUxZp02ppm5
eJAIwfKK/YfC9V8DpYorR6T3QGKwqLI97a/KS6YCcj+B3Wzt3awEzvD0uvSN0wc4CJBLc0OEGHsT
JrlSrjDW96jEYxGJmDyzOiY2VzvSwyv1rAgtQ7kEaeCkhGJd/QksIGbSfiw2WUfrfIaRtN4XG7Dp
IBOiF+WPb/wbCLSjxPI84RLj0HnPFdMXAzzMP2hnPqdOclWc9SWGMdHzbVaokvo49rVT6TgCK7Gn
v+sSDm3AttviBxEt2M6FxAnixlIEU5lwObnzyzVDLNKUP6JUjv3i4wo/xdRLfbYLiWS4XD+DkWGm
MEAmhzHGO0UZR5SxAZ0u5PrTNCS9FAU1MOaykqp88p+ohpVb0xArv2zqW65vzYdg15jWV7g5U3LV
lYe86jhhMRQOGOvPb3diCLyiM9VCRVHDAjQSH5pj/19Dd4VsubL4SMsq5Xw0+63+PH6yDlnrwH0r
DZ5h4SiwypiOMUZb26HRNkmcXecr5RlQIKgCBuE4VARI1sW6jZ/IrVEL9oay6E5zDgpbbxyQbxuO
HqQGcIAH/2Znz73oG+D3ABfI+vKg9qtIcNJnFcgwoUerSZe1JjQ1mSSyLk8ML+eVwIeK04h9bLsD
HNMvpPlufihsqtOwcWVDV+NCOUEPHPJfghWcpsJvEyT5s/BRdpfGZ1a2oxZnBdDdioSm+hQejA+9
f7CzBdRBnWzpex8uomehMlraqRZcCShS6NFiQs21XdYTebDM505ieg8gcHT1itDLBBdqQWrvenhc
y/KEtqnSvJtBrCmQHVqVPiO4bKrK30ZP2G6dDY6bEet96lqj3/VwPMkUWg0CQ2ND70UlI/f/l0JN
pP9tYPkFXbdhTHm43VO7WyWTqxEOJQoR9G6Kyf+2P4jLumhWSJBZBrGii9BuM50D2DHYsOt/OYIH
GqP49zFaY+A3NN8T3IUOEZwfROFaEx2A7LJnke4GvQIwU8Sy2PhJRl1t0oqgbTzZfoB3FCLyBGUk
pntc2c08T/OqgdYKAc/5qhA5ghmSKpS0ejFKhWFDKf9J+EV9TBzryPAXTzmcUxnXAUQ87u+X/FNu
RKUWG19ttrqZbxai/J/wwhwxCMj7IJibqxjawgUH/zLVfWiXA4tWACqI0fZ690OlHmF1QA1h1lM/
rCfd30d5UwIwgyrmLxtOO/dUGZExTP2XXzLMiYLD+sTrDBKzITY+k/56e1nSq5mNolmjXI7VtnVk
XSPnH9UQi1FLEFb8eUDgpeuvVYZDuQ9mYrnf+B1z3BMirgqKglvpVLd03utGKGaF853hWuU8sDsy
836Bep9SaVYcNXSDZ2IJXjYHHJrBZrgfzcSPnilFAGCp3v3DjMXE/HSGwZzhI1HNYtcJ5jd6uCZO
fRt2ed4nP7vlulDp7tbafClQbqOlcNyh50OVc8XWRC+a/X82BYvpPKIVRzvwYU2Wci1DHvmavYs7
TYR7zMUuBXg3O+cSOvjFXLZUSV3lvacZfZIUiK2CraiMBpOZN+Yv+cjRptGT4ke2JgCmPJwL2zJ4
dbbdOKIWyNKzMLtf0Tu0wf5+HyBXSPEOMB3LE++WRu5AjKf0SEEGsM4flkINVoB4kd9cOFSdEsTn
e7RNN3BAbvpsCcGnVEMA8CdPiJwBDb+ARwo9JwCJxKJezWT6PiI5YpZiN+tLIGb6zWB2ALJDT46K
0SNlXqndyRNAigynbo6HKA1oiMTf90LLX100ufiWmgP3BIeusDfZpXFRiDxQLp6Q/X7H7JpM48jQ
8I+WtOGC03GcYsUCNcqF7CDgf8rHjcVLeAVCtWd9yBKv6q9iYbGbPQZOMo9/kk0e1wOV1gNPlLcs
RKf980XytnXPPuG79tDn580RKM91HovIVY2/mSOt1CVCxN2IKx4bULE9NuAN7mEfjLkLrIwGlJPC
Mpka9dsZ/hhsmZhDZ8yTtuuxVtdAPuyp/T6BEUSA+qrLZt8WwFkrHuyPJTdI2L5wzLY2wZSLvJwg
N3tOn/j43+6o+/AIqj61gHzRoRjF+QYPpQHhCcN8Z8j9wHK6REny8jrEsRXIyn3OzZ83bvDf1pfT
71q/rpSo0eaLIhMacwDMVDkRs56fzRan+/FA2oWh8FV5L/dTRRj+bsJCEPHW/uuCg17DFEC2NPWA
9/2IDGCzgiC0fe51GeU2dYa/trKLzHuqa83mdJY7iNwU9dIuMLngGsP/XNMmr2JEF3mjVWqwP3dG
LAHVVbBiptBsewf5omuaB1zbNi14Bwg6xqSvmhOfdRTA6Lwnin0Bb+tNwR+pZ1K5XGZNpqJfVksK
c3zONF3Vcad6G5QcUdwGaKS8RNT7t+VLFUeCWoWXWvhovM5lN7OGxldqceENwweqQOCb+8die5fi
DTl7EkbMhVpA/V4G0fBItpMURA5dg+PB5PYcRC37N/n1WcY/JTPJ+gGXns7fi4OCMedMYJLCQVBy
c77oUVMi3XCxL8ccbmLoIhanjlUhEjBwSf63OZ9HXQT1vCF6i/V5yZGcZwkkqosJ5t3M8fFQWKor
5ETrnE90LC2mFjoTu4SABdVvJem/1JQWVVnHjcvJeg036YCnU2orm+yfNldSLxmLnasDBdK/5mhF
bpL+IjERZUg8Q9EX4RJA2vSsGQ4EFqYb9iSlSvMTnSiGtEArusGNd79RZo81wMMDt4L/yWzMNX9T
Ao/2TkXeB2CI6JhrI1UVkLP0YLtfJRRG/cq09vdW7kHweCK86PH15ZBbfv61TSs8i+Tlqx5kVnWj
eWa+7VNAElIlpwTJIVkrN5RRKF80BDu/GRaFsPyTneQpt1oGeLqpf/9a05FT/EH3ExsUKd53Xbk8
7QO0w8tbBwBX6gnXsEhmbBpQNPIdDXIfzAFrNuwwuZ7s5SPD6mOZ2g3NTtbYYIJjxlgJ3ZHXLKZZ
9EJhDdKwUvjfty2UX3iJGcPLGzYXW6rsXcjCLBVeqBZCnBmABytu6mXxEhslIgdGVRBvgF+LTGyS
+cvqyiVRcZMzHYPkKgWo9i8tJadUoLiOVSNrIMaD54sdNcrq3ba4vCHWzSjbyEamRfUMbSsR9OUS
Kmp+qlYXsoEc0ws0utaaJGxzzF5lko+Qvur5Wx7ETBVmsR9YDuB3GqI7j5YZEgQ4YIL0zqq2IXQ1
ARzjqQBo7d+KLp+djLW3c2js/xWN/MDggJJAx07ccMj26K2jSIi1+fTNMw8YYOoaf2YBLSarfKQw
1A+FRdKeUlJT5UafSydQwcG1MXFzvULKyc594kXWiz5W2OjeftpnYS2xBcEqHL4XLnUrJ8uE/6/a
FLxCDisJmyA0DaquZuRJG5iFAMlRz6eKY1aGiQGieGCr5pI5BjCU5Cz/9SApg4TmS7hIGQYbKlT2
9tJ7yjEghHpPcodifFUpxv6wQMpNqNnvknPKe3YKXy1iukKz5JPLCU25FjSiVRDtWRxepTatM2gy
pz1c2M2Y+XnXNrZzHckfzajsRLYxt7PSSHB1M/rFraixR84RfjePBq3oZ/x0uaiyvDUXP+so7564
82qezQs2vafxo8F5h8b9CKzjRoQnr3N1uilGljM7IDvB4Aj97CNBsVXQnPE1kuzxEYU660tN8CBJ
qd0gs2ed7teSnCL4ooGNrGSOhfHZO+Z75Z6ZXqi9yKtfbq7AUkLctQwXRAkMwS0MUA9tyb41wxJb
5CcyVxM9mdcKFwgQEwWs+EOTfWV8AFUi5gPJYnv71alds0/W+0aB3vTdWIT0NtK73bZDJM9PNlqv
smwd+rWYSp4j5tfJYFrhQUoEm9XRgHRUcm7Z1qRDeg9KeJZoKi8baJiI8PCNS8sMcK5BoUZsLwz5
OA9O4ksYkHwblZxcjF7aK8gjggoH47rKNt0hlUt+xyKyppFzWDjs3ytjdteyCIesBXLv+L72xu4N
RrB2QkbI4ODTf3aq8BmgWjG5DlMUoHdZ5h7GfU7US1ItfHGbazs+IAsQg3/MUY+jEz4b5qg8UHp4
72evEiDHbxLuWKnXBBXpcOmD0wB/WCFy4YigcG1ZKbpw5LpwdiTXw8/UbDmfvehk1YfpZjRfwzlJ
JIQO4tl6I6vDhfBkE4KAW1ug2XDzB+OFZoQd44fTKSRlcn/74Pm7g/rC2zYjo1p3I81MGGkSE982
hmGDFZCb2Oud1KRITMLAwa4XpQcmWsnyxoKkPUTV4EMVurrsxnLjdhi2l9A1VAaU82liGbYSz861
Z3snWEPXjf5kiqGUXgHge8WAJNdg4vDn8DWZzMRlGyoR9iDOIUq9NLhZ6wm7jKthE+mCtDmLpH8W
reflmEsOtB/6R4XhJqt1dJgD13aGdHYiG5x78dY3j38lBVQT8iNE3RfMWvNRR2TtO3yqeuETovy2
dXpXCGEbq8JjnUiHXKJvGeG1lqpdHhCLneMYgJBN5nwp91xO3oJTPeySDyfHbvpwrmv7Bc1Nlqdn
q7QQOzE4ghVEtt1dLsFiSrunn583JrRiOoHa1frpI7hPGSIdgk9qIKGBVFqM4DkVJQweunQrquAq
8qqdGi6T3g/AI6Nb80Ht3BZiH+abU9+SzYtzzCB1g/j+knXlQKzP267E6UN5TZVNbKDmhUepVJSj
MGKzo0Znkeeye6wKSbTrCqkvdrB+wrKxfE56XQDAXdtWi89kjed+bVLWxJqJHUsjv9ywhgSV7kZE
hssT6Wjx5PjbNJgcMZSfLeUiHavI7oNoxKId3TVdOaAG3xV+EF8C3kEVMhh+pP4nzGCexCDbPRg5
GVxM/0C8nt6FrrUaequhDm5hOmkdfzocxqk5YETqqoVHbuQ5f3IhI7mu4adwKEg5FuBXWwmLfNSQ
zXCoh47OIvfaWXQYzhVSuzkkgxyG8hX02igGv5MGsTozOpd0mCzzEW04uCrVHYk3GCG4tU2xVpxw
lHFp3UdoFVJS3FhnsggV2pJ3qZjfguSzcj9xcoRy9PQJ7iXBNCG2Voo/E9oEUqiDIcjBTU9ba2fK
nN+JwepkWyE7oLpmXiT+A8XeQsSIH09aOIj4fAjmnQZHUpprmSsGEvmWFvcjoR4RH/TPbbfH9OzD
9FPROI70uxPoWTNJpMDhwXxP993PJ9EsM90jyl31pkv5lPLSRxUkyd1o9jbJFigPOzWGL7wA128V
YbsrN8kZbc0Nnmzb1iWxopFuNcopyEkKHZS8TroCBN+yfloUpbHepGjpDIlfzsh+2RBamHdQkm/o
MDhJ3vYL95q6x7C60JSbvjtuzOmFHt3txhhX0zDEfFBJwlf5ku9cMO+wdNQyVWAOWVpmDNbj9GA7
J8rBnvc93q84M6hpyLSpKVEdYDeXcGmD9NWibbFJoHK9dlch6be2HMKuTtJveIGbiz/F5ZyaCvSd
MJNTg4dMDJiisW4fv/vdTgehd1FdE9qRnly3ekYO3O8M0NBnkZaugz6VqGZF9foXGqZBy5aG8cl1
SVEcNONqFXd+tJQrmHhfyTYiD/ZsqI/7Pf1Hqb4eCpxjpw4DYHoXfBbflkDenjD8vbZ5yHEusF86
pSdnCnO2mQOOGPhm7qGbqNjT5rCtEEVLgxS1Yi3eSgr1uLCH82K0mqRs7U1WYGkF5BF2T/YbODle
Hv55wAdJCNAG3R5jLZagE8ftvbQl9esFH14jcJ86G3Lz3Ka+MufW1HjmkN5JNbfR2P8ofdP3eaos
gL+DnSurxesG46SypWalM/yA/vB75/iEhHfm4xDhhYJQU3uXxHq8SA87D4bb1BHsZNrqRFQMtewB
JnekkeP5olusT65GLxQ3ROE13+Z0Hj0qiJckcIzkugSHQxg7rFdXdIStaN8w40H5luSP4Y7GKB9A
MmCDxz9itY4pR/05x6owS4A04RNeAdIojMPIErJW/CwU/tAk1GelRbyHW/DmQ9xZevZHYHAXJNrs
iMR12ItN3Fry5BNGVCYp9j/MCeSpdO1MFkwxzeaFcCmS7tBazkDErYdZNRwW9An7Tz9sqfaRo8hN
UMfi4IngVo5vqa7j1c/OvWY92JttFl+6+CsDPp1HwevPWR/R0+UXmIRHW46zdCNzmSi7968oDSa4
zjMhE+N/BDb8drfnQjM1OgeaW72HGGnllIgPp+9Nnzg63hXqUv3OXk1+mVT4dwmLdgOnwGVb0JEM
yqWkmAiRXA1eaO70e478qfH/8pPSSDrjYf9xxCK1lX/AQYIPlX59SXc72OW+pEpcnG7PY9xZDeBs
qG7tkow6rEvOCnjKpM5kNY2X3OdcVlwUSb0jjgCDz0dgnSJjodQMUwrltIJc9043p2FlmF5jefOc
aAv75HdE7+xb74TYJkSPQKOPqIkN+jIja7I+kKWmqCEWm9Ey8KRieztnEbUqJdXnosGi4AoUUWM8
z98bJ61Aekk/8dPOh2U/4ihAZg3l513EO4Pd0cBvYCcqQ+xl6J8uTePP3RzOrhR7QQYj0PcaWnW4
CL3OhwXnuXdeUGkyXoFzt62ICIigUEYrSKf48oHB8fTinTxHo6Mh4r1s8yLgegIL+/cnoiLu8rGP
3/8+v2x/mjC6o0Is6k2e0TOMO10qvrpOSGRVepSEBQwuKPp/04wMFfRReTZkszZC0tcHYDqgTBE9
2jrQXFkcscAGumDzxc+uC7KX3d4qaYJDMtCeblzfYUrzlOY7P1Fy1n8KTkd+bVheacfgATox6nzr
ggdwydKDN7i678QauBi3BtMaWprqJ6MIO/aLkaqXTMem2CVp8/m52i/4Mstf1yiCFXmOMc2BaG1X
VHlRDrRSETvmC6Jl62oCXbFVVuNWQhW+m9D7hQ6NNCUBEWvteXWfnRFw7sxTQwLpbfrbQn/zjEnq
wd+i2oQdh4YH7/wWPRBfeIGhB1mhCOzKAg4WaY8R5yECg6tT8uE67uKrQ8ZpBWbKdcRARGRnLM7W
7BW6EQnjO7JyJS3WZcLYgJpDxbcn1QnwHcXCR1Tl6O8TzTCPZjES2HlKKrfBGmNaX33KfTl5/+i2
f3W4cyvdov7afIAK9kERJxm8NAqDRYqKqaW29y43LBcBDT1Dvy88VV4rLaz6PehWJ0APewOExVC9
NW9pCeFYgV3YBMRoiH+sucqFYcgGJKkFK8e1fYtIQ79fwME8U2BmJPINImdfvrzve7NtnApSu+Fo
InuxRtfECVEaP0mZNeZjr/zI5FFvfi7Ym+wTHluGeebH0CqNOpQ0ir5VwiQzms/ZpmMbHmDkosTK
xw/r5tL1erFm0hMQgWjfmdT78v6WqrxuOECOPSxXXLUyduIXX2T4lCI+Mg+0Uls/E9h+ErSs7NUw
9NJclQ17gv/ziK/WjdytwOW3g+krCGlbS78wvT1HB/4+x+CnAJ4CWHFL9KpzXlgFkWEnqyhCWatF
4IyE5/lgeL3p4H6cKqmPyhPOm2V+hdMiSsq6PlwC6fmHfIITbzlE9qRlLQpYNLEclCTu92TdRC+6
BNqgAqMH2UYYfNXwPlchTKBTjJQUPyUlfyJ9BzBIJmCgrUyh1lYtElqqkn1tZ5Z0dioB1S3e/vU4
Yzkdjnd5c1WbzNDNCaCcpVvEpmTpRxGWYgYQKJ9w7Dv1LXqHxQgDlpTnp2PrvQIOV188j24svnF6
ryIYZr2hyNz36D5fZPDNZLyKQuq1erWoiya+/xYGtQ9MD1/XcL/JQ2SApt+RiQKeT2y8jV9MYXPF
a8W2G2S2Pa3Up1V0iuaCHhxy1wn0n0UHbp1yHneVSJxMtI687pdF1soJQx4En1noaBxE2+aJfdXz
zE5xtI+bgr5gH5npyvC50Pv0ckOjUxEeVo2b/WGbuelJS1ZfKnPQoVJfy0NxoLUwtmMnHJTwwl/I
XAWevAensnPP/J9dQpgESfnE61ysRiDrZl/v+l538bK4eqOHgJ5J0eN+sV6h0mF7Sx9c/sY0dzRk
1jR6mSVDvLm1PahPwlOcu8bhgTw1YRuCxV/juKHCDMHYWdexkMOEZTYFrfyZQdSpkhZNNz95gLPd
XPibM3z3EV/Wp9bDnsOLpvh8KloEwWOxibBUAx16djoVzz3a6tlp9Oz+gagV2npx3njyXVU3D4jz
Mn1KRAS3aQevFwGzqKpMhv1JVGdNrq4ONBwSg6O2OgVYiSPs6jCIHiuRgtNG38CbPCg7KU9jI5Yp
qxJK/ZylOAfYw5sv+cRsDY6uRL+dAFxY28A+wo9DOeBH3VyF25mqLHuJRSoDkwaGgyt0onf+PTbb
USVx6tn9Un02AXsGW53oJTD3hi+bavufX5IgLHdI94K5R67nOSSWAuDmXXHH0Y8G55nMo42JHg3C
SuWP5hC5YD0t/expR+HSjYkGfXq4zpZ/ArdzZfRohpZqP+yJbOPntXhjapvws0Z+hROnTvc99XA1
fE9Jom+wMRn80NAX4WmeBO+k81yenBdEkiZ/ttY87y/Lz/4FfURjtJNIjmz3W0RK61BNUv7bcAnB
rZ924j5BZHTgfvaj28QX9xki5eCUmfYsx+lkXdlC/hzi6rHHAAPiscw/P4mS9RnRw33KVvYuZh7I
Um34JR39dfGqzFiB9LRPLj4DVmjTteR5MQHCFMbxenPx/KX+Z2gG8FrijTfN5vRFYb6X2aKrxZZF
rzt7AJyHocel9l+E+JITWCk8fflcIUAhXXi6TXxTMek06ModMqv8aRol1ErUk49TA0dzGI1M0YCq
+Zr2QBJoSkFG3OvzeiPLwFyRN4Dat7lb8WBIaoBuWb+7sEh7+QClI6snCYQiW064pfbPK6wRbUk0
qI3N8uc5dXcXmjd7MR9YtVqmFppp8pHj2OboTxQryJMSR/Yfjdq+VlbO6sq45xQawJS0xiyaHQXP
8hsT6dPGAha/9uHKA1+USbAu4moQ/3rfSZ2QokDNFxO+kyMvb/xTte8vOc3a8H1uW2dWyDsypKYf
3bT7HH27s1IqdrUHQAY6kO5uh/rjJ87ZnEAcwUn076c3Wp28pFHBlw/COJHDDxTxJ8iFkfr8/k9J
+MojjSlSVrq5s9z58cdukZrlB4LEbokPzVBkIt705na/NRhMWOyGz/XKXVrhaZsL0JTa6VM2M5bG
4N5NKmZwqVDzanQioLPcLTCZN9yxBXhXZtsCujMe2r+NMqsoPGiGeji4vqW+Th31t1GQUgdwVc+7
62YrWa6F+Bnr8yH/Fnvz4VumIpFN5cpDN5KNj2H24yrAgSeEfznQBSvXmZiHahCwRdmFDYkKdEEg
VOSH1QOloFSrKAShX3lwq970n54m6IgAc/7n2lj6tYvTqcnvSFC4VmJsucB3sQdm68pgnqgl2owy
/Gfrx97Q3XlcYFDYxfjuVPtDQ9DznDWlu4T1MsqFrZLKnxzdHqJg7mSkH/feTJV5HN2zqGXyoLIa
OFqcPpfJXxx74PQ+yfP+mO+13ZKR9Z0CufO6R0nOLOutQiSWBVFf5ult81AfDfOo+tml1rq41m43
7tnPTArrXL4StsO6FkbAoiNML+mqT2UwpsICLsX7/y/YsQcbiF148jTW9aWr9n8I1K2j2zJfWVJ4
gQQaL5D16T06+5ujxqF7g2Z8iXVVVlI+QJ6ZMRo8aFsVCSeSij0S9SAO6ryiUJRf9oExabPJbmZf
YC/oly2QsTtJ9zHInt/WDO9glRGgI8D5LNY5h3Fse+vdXznFaLkVuswtmMA2y33BvO2Sw1Ivf8x0
5jfy1J4gTRAIv+ny1tRBxLCa7zfXkBaQXk8vakcUEE/b3UN1o8Zzd0Nav58/c2PBtwKN2ZdxjGoT
ybk0xMOvbKAUdC8fjEQud26X4hoiQ+BULZ2ITuNr15tzZCUNp5nvhg+yZ1o7RS7ZR4Ds6VC4iX1Z
FEE4P1hx6xj1oLFt845nv4IBGgGcMujbjZKVJLhDYVrwMrMPXCKxNpuPRAAlBKR/Vks0+cR34nci
pfzatz2wgMtOqvZ5hoIQ3oLTOGKs//OUkRmUn3JlftwlDG+Xn9B8e4i0AMivmUSIc/Jw2BE2E+a8
4qdFx7vZypzUe1IMpA7BRWNY8m1Yalvmh/+rZ5I1//aqTeXdaCNrtnvFOL8DdWYONuVn9rfUrMw/
hBTaztcqo9j5+vxDyMRLwG084Tnw/Q9MZDoLUUmEJ+ae+t2JvGyqwOe/JOX7L4Zme1N0mjM6n16Y
pxMLZIcqLGRIPHIWy75EUZcGK/uFKS6JhC20oDJN4RFPW5kdCbyKgNgepwWgaoWDPSGqp1l2VYUf
xdfZmGHKuaKd2FOxvFr3r53OE7PsfmiM1+9EAfuzJqGR5DQ/KhCYi4erxiRKK6mhjGCxZX54AhqB
GgjMVbP0eG4oiThINZ4w6dUJigpoAPJipJ45EnyMgRtllcqboTUoBieIOiKt3ed6ub642/Zo86ar
YvbLwqCNpTTksV6wReFcedXijYCVO8+a8n1NRcu2ZuYs0evicrCEVmsqqpW9of+hbOG4XjhS2Qot
rSC7uaKeOvuNZ6BkQAnCaMZ1zKKWS7hevJUAezlAj0ajmxpIRYE9YzcaN5P7eyFRss3srahZHMbx
wz/lpLDjekCjsY3TLgVMifgn0bvlJNdKM4co1yqRihs19UJozc9gXinvlgCawHHvy1AZPWfLrfrk
vh0W3XSviBMu/RRjMfTvWblru2l1bpCe603AG8N6+wNv3SVcK8IZWzql/Kw97U4TMpCUfD1UacZ+
kFZHKlBM6Fg86kJ0n/wUALKdJGEXxT7d1Yg7Ou+kplJ9qIiSo2dhi0hLMax1AIIQAPhqOXjqufY3
G9jGIViVf+uhVYly5DS1NoDFJAVfGWPmRkyiGkOLvsBICGAyS9YzOlE+EDTPLeVByZtvtu/zdOXX
3sc7DuqE1f4zkfpgNo9ESTcWqfFomiF7ST8dCXcfNavPhS+egz3UyephGaN5M9TE4d18c5fmuC5/
YiACkCCzDbNPBBE3O7+6GonAb6xm9SDJ7tU7mZQ1zaturRHcoT/+j/Twbr0zWzcVRk6g9sHMMUEG
qq64OSZ9Se6UMns0kS322Wd7PKL5y43h4oGvgvAuRv0kXRWsbpCZ8STaHMwig54t71h90jS0OJ/U
W+Ayr0soqWvZmtvaeaGOYTZ1o/WK1ty0vpFEoEpBE4NS5zex2WUTYtvc/svZaJa2+KWDekOERwvX
g+D9hke/rmzorvNCHUcShkGeYEJmUyQBQz35c3iKjW7OPsKQkZujwMW9Auy3WLKzuHUr8rzC2Sda
SldegRdKE1/wPNAWlqCE2DYmQl1W/RRXG0qs+W2+QU0u5UY2lLACFRxXnztut/+t4OEQiXf1Yrx5
RBUjgG0djsHGQ3X+Fv6iI6raLxh+pYV7sgmoBxXPPsV9PB9QujLKcN0BG/aOYBlaLwumhJiTaNit
7LJnB39MtOJ0ND1oWo7OaB01uScphYguSFofhWPnOdVMtd8ASH3wn+EI8ADJNY+Oh1ovBc8xZLKI
dLMoHkpMrf8fHRvCG+8mbPIJTSGBxgXa+meDjBpqMBMPMX7C+0iQgJsfsjW9rjXi2kk7ZQ2U11vP
nBXpDY8TvBWdpLUxkmM6//+JCZ3fYw1mZXCq5HKatQU7F7yascomEU5DrMDmhpUkTZ1D1NvtRR6m
8Gvrf3Pu7+Q763OA3LPEXUCKUERGs+04YBfLcaFuha1lcQ0wTxcmL9DcFCF+5Np881edMptGaQ55
bmrMlErZ67X2TlR0tL+MT6XHuHV1EgDVVvPZG7C3O9dynuSI4qcot5kORYlnaUMvnQlwydW+CC7b
vPuVoYI0v4QqvCZ0dji8uihwnxGrIj5uwy9G0mz0IHHNIT1M1lABx3vJ+tibSEll4MAa3y3aYOR9
c1DDWj8o5SKVEktYZd2Cgo5tRjxwEKfLxAcNPgWCOQlaC+V65zkDhP/qa9CRk+yBt5gq0qflRJMh
g21IigMhdqlDAckqavARZEvQbfEP+yTz2y/zGayfhPLkmyHR10Ebz+PlEDDzb6wMXawS6pPI/Y/D
ffEcj1AtY9WKhx0gFIRdOjbAlOJJhT+wrJS3CRBpUstFebtTBolvaVSoXMiBxBRi3SQrL1Flw7uf
CzaFy3XH0QwTbMDwIbwknjUqPB4Vx5yZrpjJ4ortnejL9hd34ld5+4FDhLEl9ApOw+lUkHFc/k8n
g1uGMg+LM/DJBoAW436/7AH3zQ53sRtnsoguqhU9f+o/uRjQW4mfZzmfUyNk+D98wb7NleIWxZJC
hifGBCwa97AWVBPUou9Kq3e0jLlhHkNpSUFmLY68KSMXsF/3spIhUxQXRRsxN9XvtYZjKsDHJhsf
5j0G5jly51k72kuhYP0Vq6xAVpSVFs9sZxG9LVzNYnjy6aDJsRYHreRjoFNkC+3ES4bBPbANG6+a
3MPgIFdcd9plTjuDp7iK90P7asUKre8tgDQpsnFX41Q6JaAsc1hTM85YaHgKRvbZJ8Zpmp9LZSIV
MkOFCe5hD6/Rr/1Nt9soO5xEFdaYPbp6EAbM8CbrjZzJDubct55tCOjbaY+IdS1Xl11tdLA/3X9L
xic2MgVwgZKVXHlBgDKK411b7giOibyH2LmQSn474VmdqnHQdOx5HCLJpZAJIb4NrxXcSyyMc6pK
VDnu6HpI0LqTm/6OVg3WU1tqpyRGGxmbBwVBgISi3CN/j0qkZb8YxsQt3haQpGOzsr2JtaeUhBsL
evLG1MfT5RXP5q0t/gaPzoMjRVEJit+rdTfTIqnzjMW3Du7f2fC1XecinQfFpCc74cm3s9xmkHnm
fTV5u5o/PxrafeDINMrDVtxm4eiQDyN1zgx//5aUYRVUTg6gFIveXnmpxMD0o6vGM7Duj4oqUL0J
+9zDn+eBAznzse3D+L9zv9cy1Ylhr9cJfs0tIsUlN61CMcVr5l85jp3r4f3Z2ETmlTz+vw6Dy3To
TOTA7Zgh1xU/LlAcB+VoEb4HD6U0FhNCXBxeGGhnWqvzL0cjkIo8Gfrym7Vvrhvuitx3pQqCL+P2
xgEcUFuz8GhGl5bW8UffHLk6wUEG23M8dbaQysVklzjcHmpmE7SWVfq8a930vA+Et8xwfbo26wtI
s3fnl3e9R5BguSFmYAc7Gxg6uU/l3zDA2cRzXChKp0fkfXfSiERUxyBcvNqKPB/w+h85EDSxleTb
YNnxPfj9X8rNq1OHHDHO2mO66R+5zwcUk2Z1spveV6UxzxzuuMdBOwZ+ShahEUixmStxgNozUx+6
5Y3MPQJ5udFyma634s/co0itr/CQWhANbugTQeVWUTC3UxGNNK9Nz5bUgPqf/Q+Z3AOTqhosTwkk
KLF7tBddeQg0yuFHUnu/Y9vxk45Qf2/dVr9v0/eumkkUirYCiTsH1lpCA7Y/QSz3CL/+vm+ZxVbF
SnVbbfX03rMa6uFO/H8lgGw2iu5jfujMR7C/VpvTyFvIvN9pog0Gq/YOm+6k+P73llb2arlPNQ4z
xXGmZHfhrpn9Fatg0X26W4xijueT6axgJRwsMP4FeSTisYH7t0+asPX+7VVCjispbDj7uLgo5qpf
aaXKPgCvmVv4jckLmJHmwVko5WLknWznEtwNDKzF17+bb6dURFFDTIiTIYhtGCkZKlLqQ0QU/945
cFG+zeOfecbLkWcXzFNot0AhQPdn18XVxrLqgpKns5TIyOcsEjkeP5qrYhYfxgGQgtvXmhGZlwFq
ipuiCRUh3TkHnGMIpXMPCPV5hEt2buaubfw3ErErN2FyG15BnphuSOHswnZcyRj7zD7rf8/YnV18
Y6qRLE6kzEXvAkLldRddRgEpDM6oa2WpWupUFj5KnybgaxRDw0wnC1wVulXTc2CaQNHAq3kQvLz8
L+k7HlfMEAQMKOS67pokQSOkCQG7wQmX4veAuKHXmoXY/u1hFty2RpnCsrhWZL56dxNplzMbeapu
7bEjO9XMUicBWWyA7ahjDXKTSyI0rMKzlUcxLaf7Rc87cGJL+O7om863j8P9X4sKBcrfxU8mdZoO
l8WSf/M19pw6Tdt+vYMrAgjujBgz2OWAQIfg56rkZ5ApZ+RzGUsD156jcv72TUCuZ5UaCxpJeOip
DrFs00mhV01pRnyZwH88POCZrtf2tCgCvU7rsCT5sNA0HVAsyvz9B6tkFOhBhd09z3k0+gGilY5K
9/TtVxxOeGGqOPahLsNTS1ZzMkC1jMebgSORdgfH0G5aJoFzRhvyE1JWgTBPcikcisenPYsh+rp6
Ea6tuVb3xsgMkSELAZM7qJ4lqBgDDwVcybCrEe5RXlT9ZN8afUmEJPbWM9VDhOfJ23qbD7XvlgEi
ba/vXinyIr6Ezh++1L0v4NHKLpZWvXzbCR91mPHQVS6z6FRATCl2bu063deCUS/6szcW30WwTd8Z
8jiDQJgeZbOHalW4D+g6LiZjTlGU7gzd7dMIKFw6fiNgfW0WVg8kWfLRdIE9tASFs1mzt0C0Rvdk
Dr3eHJ5U7L59cAWFqJCZ1S2eSjgJB56xcS7cFVtiKtxXJecgK5BKXoro479+ljSGFjFxij4NV9mO
LjNRZuUdfe6tGl4m8CTCQfqiFWtC1YuiiCesNyO2nVn6IT4b6MsE7OdNLNhxkexlPEMDfOCpj/O2
FZvJf6g/ZvxDxTUVKJo8FonrertaaeB1N+ykGw3EWEDeM1QIqK2g9djO+uAJ+S/ylX2iBl2d5d1W
pcpJnp5eeRRXabRBm4UjSuDMKoJ4S4xztXKcDuKxAq7G+xQeLiwH7A4KqPJTbzkwrWm0/qAFWiKM
WiJCKSgpwrnMcOlFXLflSb3/Ve+9cCNiOZiQSHP/HEIHkzdfcV0Rf3HPUo59kLeETTkJ/P8AfplN
bs16J3zSBNhYx9WmosqcsuOvx3BZEv/nz3LaWLwHjXaymzUthSgfLW/1eow2/3Ranw+PIbshgH/S
lUCPZePGPgkNtGHZOBFcfHHNj985LIypMt2F/n9NNqMxOsHcIHqMAGg6b5ciyP2jYxjuUlJMyS3q
DbL4qjBu3yiR6HfITQbUyaUm9H+1BsN5O3Z2C4SGMI5ZUX9IYz0ilYHgZvKbarHp1735eu5DKL4t
yV8/hQsNPhrFhvrIjV+RJVwF6GGOrn8DszYbtjj5cQv9QzHMhLShE6LJmiukikFMBiLJVW2/ond+
f6BgNwpR7GEj9vZQlNrNd8Rt6eay/kgt9/iOD2mpHNJ7XRZQtjPGKblY7FnghYJwNwQEpyHSKosX
dSLLoGcfREO813Dx0JR59q916lA/L6GVyiwilmD++8HxHm4niohTwR9FsHnEtd6X0QUvjafHqv7K
btxxs3m1+5Yc8n0Pu/M83v5hYFQZxKaDKr3SkS88nUOs0x5nRo2+kS7apiN5GBD28LLyF82WGyLY
7zloBqesXg257XIAFPgPUsyjr3VnHNq3C5dsQJx7VhD6OwDo7PnxCv26Dbi6ZR8B4HIbjiF7zV7L
vMTOC58Mw/aot+WzdkESnwv+TnZXPUrqWOPFT7+/x1Yvo0YCRLvl3VTYb/kT3zwmZpH9jwGdevYV
Sps1KwTXqtnRVZahbIkoOJKQ1SGx6TTbwO1ZRgxXK2v8rH9xjityix0siWlkmhtwRyN8KXFJyRWt
1IVJ1Kt8N0FesBgwFP/SExn5o0cq1sH5MneYp7/XkW1m92CoJdaONC4TYdzBV4kOZ++ZaasZk2L0
H2zQRqF7BNV1nt3PSOq2i2y+uJubuPrLlx782fPM1XcNFAcaqFoV8ZDLtaojtCHQt7BJzv8yMirh
838acS1Qkqw3vX7IW6Gq3DG34qVezgmRbAv/nG0/3SO6caFsAaIV8xbQq/TlSxtB4as/4FXvae8O
eszhGAQsn9Q7zcgJDoSthG/y0d3V5TmhfwkfAvXxK8p90sAWKZlLB5V0+uvIV64j7dp8SrIUw+QB
eMkEobnu/pC5tS2mjGWYUR8gOokpagMyH1l5tt86tqe6EgYbW2+0rflWc6xC5BLWLbbe9dhFIqUF
156y5mVS445eUCUKAPCbeO+5hphZu7Yawkz0uqQgSCaXuBDdu0nBFjGC8ruiI94/M0fV777nJ/Q0
XD4IP1t46tAkafc+bXgcwlIEoVLGj/xByJg4PXdFzm21Z1KO1DWuWXlWKcsuIC+BPimxq9OdMmrV
Dhxtm0WF0O9EOh7xkPgs98Ffh0Pi1iefH+NCSJGtwACSgoYl+7+Ha540ork7WI12M/aKTxAUWsh/
hMArHylaTEKd9SEL/PukSxDzcc2T9R/95Do58oj1ak+gCuX1uU+NGJkhRlwnII2Sw61Y+Fouuhzt
w4h8EJ1G5zboHtMJELFVOEcUl/ux+u+vkazV/Tfk956kw3oMY87ZmMXSDSghEO/Si3u/OcFkx0DG
Prg6wCyb+4H44gUfuX/OLBs+15/faYoexAvvMwod/qUwC9H0t69E7nKQ7v6GAVh2+d9VUTtrBnGM
xg5sB/GmnK13kp/GAXonnK/Y9IdlY1V8+zmL7YgJ6aVQUH56hPEZ93EPVWtGwZZFfcy+lTnyH0Kh
hvzkqlYAcntCc5mMzaXFQhT9NDELal0fCrSwXV56adDdVg0jFwl6EzUNAdDBBlryRYvOSwST76AM
2TLHguqEZXpWx9YBIKKBVXV9DtVbHzYmg8cgDyb4QsDgSWP0V9YT0atUxFmw/CVBJPNRp/VgsU9S
/H119YyNsSmPwkkwZ8+6Rt44ANu926K2L/u8fxCpcZpKTwHN5Sql45Pv6ySHWyaRGtOBBGsCOSnP
BrTkntOCEfi5n0IWMcgpGffTJaaw9QzXp2dgWyRQZtYDYd+Pihu7c2GdNULs6ZSBRoWaMKmnyuaw
gTpD4ISaUnFLoSVWsPhAIBg1pB6eYVUE9SS4Tj9Lbs4TEo9UYR1RfQPeE0u4JK4jzSnCzmacdgrP
d35yQO9TUZ7PqtMQmN5L284+TKXDXyS0VNelbgDlmnviaPXN78RQvTtyxVlUA7gZZxXmj3HdQgEi
5lHFbZsKFBt02CneW9Z8LlCA/LKL/TMz4UM3VzqINH8mt1FV/JCcYzlvXm8MeNu4YWbjEeuo1bee
2Q9zB/JVv5x0vl3Mnh+v10wCODe19Bln3CyQ1mwSfcjslTqFOy7t5hqxYo5H9E0ECSqaO8OlrYAK
n3HH52pYX3hWfIvwwSYIw4D8MZyQB4KitD/FWOO7IlDzql8pzb/E5/cpQx8XoMYyOZ8jWn0KROI4
D8qs+AJ/lKL8u5xeurBgI+0D5qQc6kAtfKiXCpKvWRNRASQKIR3ZozSIFs1d/hP/U8EFQ6wA6oS1
VwMDuLH9F1zWSJkTz8ap7gWn43XDN2hY/X1+lsNGIJ1BB89otfBsgSOniuRR+ciJQyQHwT0WIi3x
NoRbZC8vB6SMzJcGQd9fB4rzV3bEVTPdVS61tFHcXTvNi+ICapbkTNNH7B+jFLdh/lIgZXtbAcpe
iGw3BdOXikR/YNEVPkVhyvUU6k4XHgYx7S41gyIzRUYag2KALWnP7i/v0jQKeAPx8BtI1wrKsMG/
SZ9P3yq1N0Q2rM+x1DTd05fQiv7JfY1B/EF/UJkW9IXYkdPjUVuWpYyfB2AuT9xKR048lqgcYx+y
XU8kafami64kThiAAQs19RmMf3Q3dITZfG3Q4xZBI55dRbhNRUUI0pqE234ONFlhW8Bf2jG/aDVU
TgX2POltNbAXYr732tg3vdgA3vVq46q6cWAawJj46BFP5+ZjH2BXzI8XS00LAhS7bTYE2jjpoI6f
Cv3rkQCujHnoruBWNVvyh1Dn+C4t7aOut0LzaaaygGchMw3EEEdSJWsybiOQRYvVLiLwpos2oOb3
wADSjMU4iZHoLe3vMxrET8QAG7gT/DHj6WJJAwYMpOWBgz74QIHWgT87iTkZ9cxm4+H4qIZnhBPg
IxInZ2sR2V7YNMrHRAGhxfcdWqkYD2GB50C48X/cl2B8FL7upb1SGYI/MjZSl43kmPbMoE2fSTpX
QNIRbYSsvjGXU83Nz2G7CtJr3qaBJdVBKREjeIOHjJBE+G8SMQ1NimvPybtKMUwNsOuPhMCxoJ1H
icdRID5gS/gq6PBJrENIJAKmD3Se9sUfAV/Xpld7NHWNbKDuLvgiUiv+H5hVUS69p1JxARas+372
qHToY4MgB+LwHoR57xUvE6jF7W7lNbH7X5S2w8gwRqGBrVl2xHd7GshNPpHUUwplmH4PtBtaNj7j
bSfaHpaFwIdVS5SiUznH+y9GLQ+SLDGgMijjmzW8C5K2GfNAQ+bWv87NYMy8btGWJvvi4gV4bao/
B7GRjLLWVgNYCD62DutqpQuABTJ2y7tRH93J57bX+o8yULUWeFJVAc3KLVR6Q+EMH7YKoPiqPbiI
+K2hRkBU7fb3XSXbrBDJwZG5iCrN5JAyU6xi3whde9jxXSabGcZvJCs9D86QfHfD7Hj9UEgtbPJa
gnAZrvuGjudhgAsuofZcsjg9bFje+YlQKoljRU2Ywm3u93yLcPxKKXfVXlPw4/MQXE0czAQ7SAdH
AlLBE5F9RH2d9HRokEMKAtZmuwM1AyOHPQaAUhGb559P5/2N7LMkHAAHojNGNVbbE07SBywoZs+N
wK2vV5m3nLvHWmAZZfAHnMy/wUYwgtqPtS0pOC82vdegc/cLo23n4nsqmIK7DGNTgQ7Ntey7UqX1
Pkz5X3IXeW5vo6gSnhFUIbFrbjsk4ShU0hR2bpYj7d7SNaoW7KulY6JN6dm8GMKg5iabqq8IzQIv
OoGrJT8osjjlIv5QETe/UYmVNSRt9mPqlp5sa7fyBbmtwdKOSaAgOeuc5Y3bMpmRyOs6cIkGvcsm
6DLu36NedaC91NH4y4HRuj5NFbS2UhY/W0jUU5QtjqguRoBZfrSNb5FCnXQwzX/bi1Xo16j9HlP5
5r6P2zcfX+cArH7dSCbTwsQ11zKgzf7Khv6FLYxzo5Rs653cU3O9cONd1cAF4pSIbGz2w+iIus1f
m6aqzv5hTqEJ9CjiwdV/2LhemysMEXnrC8TBRKtDz6qFKhtJnuN/SSsH9T3zbYgmV0sSrwIzVd7B
uOoT5wmHu/Bo5XeMhNP18jT3LOhUDp/AwHGtVrf39sh6x18sGQVP3WTUOSAjNPC3mjHNKJ0xfvcR
AgHJnhyrKtJmRgl1Lq5RX+ZUVj7EmKcvUISaS7Ed2/UVWj8hiV2vfsaWNG/DRcPxAH8tYrEbjVB/
Q9JsJxIshoIO3et/povbA9dJWglu/dFSFIw7z2u1gsPNZykqgOeDRlcNDBUlRTg0oZZAFdmktWNf
oJmaJWuq/M20r2iJzE6u4e1lMPRSil1WZ1NHVVy03W9EH+Y0KQEMRrjSHeCXoBgxvwT8XBLOev0S
yv/aVQSrx21mcVO9jpMJW47ogjvEynGsJ4NYc2oYsie2AkkL8NLjgg1xYz7/7+MpuusZZDTIhcAJ
R8pjwqBjjYsufU96td+e0sf8jhb+4HymyqWBGp6uKGoGhV6ixGWhlxeIDIRa3tg+N54p6B3yoAP5
3PY9e1ImaatOVWGJbHk3ulw+N0o4v3Bez4rY/9AXYKtiw97W50nGtF29CHCKeLEofjVKWwQatApR
T+CE9b0Y81JNUfmEBO2fV8MjpTEMN0zVIIxCjg2o206PMo/wdu636cV3E1Fmc81UnSnys4HN2qSH
NkbDja/13oZLj7fkKOERPRQkH8ijptnWO/FjMAz9BhcaxN7MCg6zcoeoT4FuivvUxVTK8BjkiURX
IcQZsKwXyx0A57Bq+jmZwMGEDUTBrUWwjKgFui6PVWvogYwFX88/1u1OlOhPS+uTg2bf/f6WC/Uw
Pd/VFFrYqsNuoMrYtTp3CvMW5lC6avFhwQa7jKiWtPcavse7mIR0adRDycWoRXDKUitU3n31Ypod
Rjx9ty567r2uutwL4g+NVcbPhlbAEw3DYLLwCml5oL75V5fuQ/uNYMZPrJgyfYo83f3J7+2Ch8RO
utQNxX7qq1cEnr+y6KC7HIIN8ZSyUxbVXIoPRgSXz2t/acbHs8SPVvPuuRKlDigaXBrjVxpRgHQc
NDk1+XtCHAMcNC0LIVX2OgAdiQwlgytXABm5n/1BsF+kRDhbFhE1a4gbkHqPc5d2zUN7L3D8Gpta
avw3qS3xxZwgtrENN8j2k8kfd3p4iYmDgxYc/bF7y1VsE6tgaqna5Z5EfAUd5eXv+DobTurDf5UQ
pdkPUVVMGHmExB7tvu1E6Et/mbvTbGtBtFf4EtZBkZ1GjZtS9Ad0SaiVksCdrpKjqU2Pj/vRCzT7
VX29XmyAC8G84Bwy6BSV2EbuWsU9OhZtesgnM1xiyyFgDfQlvQTmdFgtRwdaBWbruquv1KjiJqjX
s+ohBCyd2XuoTPeb+92GcXYlApY7h/yylJWu0BAlakOnihBrmSNPAAYfn7NogAlT3ndupVQuXTp8
sUxN4foMeuSXj1PLoSdQorZKWa4QpoRMZcs/Cwep5q6bK2GKXu6BOmaGzBQF//1mVz2/+eEsAw/v
Knmka2LTzaMb/44R8fRZ4GDC1ZrnCqlcEMnqKZ8vFflbMJwBOB3c/KIb/l860a3GrmHxt1Ds5ISQ
yjO2eEj/cfCd9rEESXkxqEIkTOjegHvXnYtBm6ADKRnQ93beRXlOEV9zXtcaBZT2Vc3qubWMLrSl
hBbatg711Egm3mQAjyg+xI5b1XXIEeAMVmLfcCziY7pbsbmH302SjiV346Y+uV3GdiPwYEllYo+y
CTudi5CFRJir/UMaW+dFIKYAx5E+zkUzXjrdX/AjS1mdFTg4wUH/9aSEB2zBNvU5/sCmKFMTZnKM
YAkN3VUp/6i07Mi1vRZhj8eAHzpOckb4iWNqCzPyhu1i+FxzQrL9Z22BtsphWAdRIKc6MQxCTcRm
qoirBnpWQv/BQD3u/27lzqfUi51bMnZqQj2ea8D7/hNFEt7h0yRA0iQHR0UQoZ0lQlh14l2TscrJ
RyDZVCOF/jlCk3m+Wy8e+e1aY6cbOxr6/WqIIIwdyMZ1/kz/jdZogyuS7f+yKqrhOoOxNHiq+u8l
0I0Av7S/fFEMIbZvP7hlWdC7IAxxjyxQQrL6/32MJf83kGcHT03m/wVoCgxSQAISd2joewKN6vbA
gXHlJfgJDeGXjzE6/mrvXXlfhPqMS7HiPx9GgxYflBeq6+KtgmJUo7NzphzcfQrYCeJQGCkyfznd
7X/rvrY6VoKI0tVNB7r7/93V8HsbKCOTkw21M8g29euVhuIaRxoOa4bVajQiBQlia4OQiK5UTREo
QcNNPOHR0gOCddp1FoQBd+UzaMOfDeLLuRdZ08rJYWV2Yh+wJZwSHo44Vx0VBJR2mmKGVZbEPuro
dK9GJbOZ6y4WMcGEMxq99vbnFptZcKKmvWxz3htn6NQDyhJ2eH9MwSNg0XFIVspslTnu8GEg3Jmf
xSsPbH6tZyPb+UDQBBb5OwOQWegWapBlDlIlIpY1PNHXYWKXQWq3wpAKmh79eUbSnlCmgXqk+3nE
vghDvr4E9x+8aV84ojYcDPZ+Tee/MD8ZIlpN3NPmWgTnTcAa+mvAESdnnSfVHkCvAC/7qf2uPTvx
enHK4//pet22cknTJRSFiW5fAhmYBfJBE4dSeq6oSVrdW6C/b+dUDlr7fKnyeVEeyFAHDYVn0kA9
LZOhXjW9iAIcOcG28qgQ29GkkLOmS133SLidwaseKA1Mj+6VhIdSQEglz7N4bS0SJ2PCcnP2sp8a
DyHpLNbk7cOvzfRf2pN9supml0EKH7zkwjks2Mk6Tyu+ASjt/avvf5vC8DReAOyhzkSPYhBh0r6M
E8rQ+xZgc8bIK3qvkVQwaeSZ6/m5FYA7JaUHTSs/1CL8dxy/YA2IcOMeOONITY9ezenInkZJ9qRl
N12ykO8Jkbwkto7goRUzFnY2LwmHdxAEEkwInYvT0sCkR2sb6EIjCCWXqMYMRByMyMfBay9gIujN
nKc/yJmCsw/8oDFfLWv8qabLTpEbdbGxIpK0v7TmGtZq1yfqgm4PW074yyfiKEYFKlBtYmYJ/HUy
NZWlxqKB5l5e2j5dwXZRIlSZdvsEvbpuGklQ96EzIrTmeyEFEZ8d8wLTdLJFuhx9Fvfe5z6Esf+9
S7FHnoBb5ASl8uMeRewXIx1jrIGza1h4RUFE0pQ7iV92wgAeqzn0wLQji36EJ03RB3sYN8zKnXT9
J8RF22YeTaH9sXEpR/iXuAd6AW5Aqv3Y+V6NCGPBM9nSnmhQTy9TJTj/1oqulaNleezw/QULdqQl
0vGiIvXI+9TZUhQSOTsn2DimhcyBikAhkbNDmEHytySVT12aIvB9+cbhZBoUeFkirKYA/V93CENk
q3aaMr6dViFA+GXGs7/fxPAuwFaCtimdZK9h5a3ef6n/2zitLyk7NAOFtdi8etEVwtpKwAb/+tul
XrDgNXsPzR9IqAQGX3xxBMgs7Oz83LlL9p/GA/c3yeGxlorlIoTFYWvruvYtFJoa3gXWmCKpbLBc
PmXBoRtZ0VP9dyRXn2JXvs/8C8miX4dJ2YJF17qdzSO735AX6ORR2ChYv5/jjOsHpqkLfW4r7e8+
/zr1BW+/ZeYvDmYItXCLXgAPRhBIocml60524kSX8eBaDdf7wTPo/8FQLCGgoFDcZaienoZxBlgT
FO1p15IXMHbtY2VdD2Uz2ccaYXKVC5VukmgxMDSxo9XylbdO5xDA8cW3PJ9YZfgAJNez4Wx/lrJ2
sLWnbeh+9705Ze0FtE5hAHvQ0aOlvJ4T5xyxmooEciAjCiWgNZBa23AWeGfe4tGxtlgb42d7ufKI
EccGR1UqHomdfCJa9UHX37ZBFsijRXXqEv27A93Ckn8uZmSWSczJpUAD6OV0GAos7awGT6r3cTPL
xrcUmcx7n939YsumQPtJXy2i73qUCb8T/IbYAj6b+XRrMEiudGw6VooslGaw8U/8L1A7VZJMnnca
6E4LV5UUT7k+RSp6vKlUgWSa1ucezHVcVDfROC1kRw1tbDw2HnatKTSZH7TS5dKs+brqfYBO3VIR
DmTtzm8taKsaguKX6+zo609UPT8wBnHf6NwL0bkB/H3hsYRBY+pPH9pQ0yoWSYzIfQt3Ti8XhQdO
Xpg1/CSr21HUrst6dUkRzakRQc9MVgr/Gi8ZYOIbkPZu/lzPbTiNcLLmwJaVMdHsTgMxjPva/xL6
HX3WUC1GXTPUP/H1WIx5+6AldDFDsKh0boalDGVFywPfbjTWfZ0pxfOtX+fWbzkwOhUTzixGKU0Y
6Q9kE4PJWfuFpOII1dnEDKlGK6WzfM1VcCFdZ36HVw0UiL+9FWThNsz1EZrkQCc/NlQxprNXZ+on
t1hTWRTXSqbsPOSe1K6Ps6uxWYr+pK7CM0McJC+9CWW/F85ibCS/T+miW0hdVuBQ+aQ40qu0ZAR0
WzC5F+TEhMdRmOaZ9eXTckv22DvI77gGUXasNor/P0MAgzn/cFMpFJhw3g6eWFr2iCPpIbgwCnGv
EcoAPK00eqRYejdDrxBqEoDyKrCfhpyn2RESazk08evxYcLYdPfeolKKbERv/tDNdS/G1vu66/xT
iplsXRIz8edbMtha9Kfq56i4DEgo8UL3TfiyxNKmHT/cyiqqEcDfJEqafwvxUsQkAzAgHiQNEimV
amUamLLA8lUutgvdx1SYfcedsTUIs7fMgWtBni335bMpSdWAaJqe3sxDBJ3HpnATKPsAKUTneDLE
RLnKG+wV9ZzrVV0suPrHCeEGenk6+GMmbkN2jO3HUquQHswHklm0yGmjHin5raUQ9PXd2IGa5nJ5
Whjrm4VHyz78IkwDUPz2v7gzUAs+RLbHVHoenCdV57w9FaPxwG1dRIKe4kdp15TQnayRSeNjvmeX
1aeSrePBG8nf9rbz6jtXF4wPmRcPt2fykG3h2vghN+ezBrkVoC3fNMqMJnqDD8QrRC2pPVU3owXv
CVcQ3Et9+Zq0WwaXSpcnkRkcQTWOeSVEasvYcfSSNB3rrE5S9TQFoz7p9xbBX7uAigLAaI1ISc9v
0FEgcSJ8iZxqj//Oco9c7FtT5OSNveZnY/qZiLVjfIa1SEBVRiEOkQn8je/itJgdmoxafdq1iexo
gyMg62PUr3NC5XqEHFdWkJ5pnkhnVP+WSG4tmwSPCtzZEJ2OBguC/5xUzrQ+8H0sQYV5BPD5FYuO
4Z2dH4XB0du1ucDAd2ibcH8NxOKGTowdUbwuOFlZ2MWFqHgh9csIq8VgnaxAnziQI7dNQZNOuVPo
OTMOcO4Zh2ct14Pc8rLH3/xo69wzr77UxdVZzhwptn5RrU2apDDTM7OEtRcCwIeUbvAn8b70tVg4
Cmw7CYl6aauKmWHTNfpOscby51he+V1STQiXU1Ecp2GNQV02fWnN7b7J9yCf/iKuUzR6mihuDNLt
NTx3TpsddH2IDHX3xTIRnpNQ6nwICxm+y+SCv9qlqbjfzlytdTZ0K3UczwnJDq/Yo6HmQ07lCAab
avWvkqQ0/0vblLOcnNinhNykzAlMvA7aOmoyapjRzVrOAy/gQjVxFxcYV/CbHZV0zecLLuHjV/b3
w48T5Kvs77J+ydqUpTMeE7v5r2grweA8NSOQgpxd6AmCmN/Fu/dgX2f5tmvaCrHLBoQmTALwXC6n
cz6vQgbF1Ul1P143gsib9UhIQ7O0u/FJu12VDcJwUDJ9B3hFggeOlqHMdnAB+GZ6j2Y/DGmu0zYT
9Az2QEUQRsG2xPI+XU5DfOhS8TCnrtvmETbXaNrVOBeYiTXsQBuvFzcoU9bCNnfONOx1QqL6WyAL
OmoFHtK602vqVg9Mh5r6O+5n4Cig3B/UXsOF0AFX0Sx6jeT9TmWS7fEdoYQx5HU6SjNQXPMaxC4n
Og7IkaUds0HAjzCj581+3nPJLbmJ794zlwvpPVof43nNGsvIZWKxgb/7usZ7AHtxq/SgQjZ2xTHK
iZlAKYEq8z7migRfimuzMPwdBrCjBI0XS7EH5Nrfv2umxRkjh+hc3+Mw0PfkxyhYoL80X+bqKH9w
4N2wqE+RoSDqRbLxvk8vJQHgvUnoBrc4YS2aQIOAfEZ3T4LuDQ6qLSrEkSXJYaokXTd2hyKuiTTH
OtsIv8EJdw0aSApSOBev++s/jJoCWfL+TSw6u3uQxC6rgqKy8BZiVM7m4JWujX9q8NFsPaPqjCID
cakic0tTUmzpN4ILzNr9GGavlOU0smn1M2gmRmox6N7KJRgvOV2H/MPMe/nP8xEWWmlHelbWAl4Z
WUcjPWcJTi25yHr/q8EN/j9eagVfgLJsZO4NktrqdbySkluGJ25HENXqFuKsmSiyj2j2SB/t3jxH
VryJVgeqVEplr3yM/u3mdcu1rKR3agQfQbotxxPlpj13MGeAji2AxPIaMdDizGRtZb6cD5qXtp8+
0I4Ki+l3zV30cTpVfdsqTQ9x0TS9WMSPMYVAsgw6wNP5J+fAJhZ+IyC1TXAc0BgQ51keHSCSY6+u
ihb3UEB/WhgSNUl2nSi0w+ONW86KLsx6tTYXYpVcRNBpTdmB1DGmJpcZqjFzLl2qw/4oOUELZH8D
Rorl+x9OmHaCpsDqktb/uzzfsnEsflE/yhbnHRceJHrSzCX7qmRb60pVFXdJ21lCppgre+g4hQQy
nbzB6PK8kuLAZ/V2M7FR3eXlOcnIIbu33jo4GPbvSyvu9mWbJaOBIH+DwNPz2swfcE4yB212dcd4
ODwUIrpOy24RUw1NgV3VXovs2XsCzAqEbwNL5e3yVweslD/KvQOWic6M7ZsSynkZ3MvZti6ICq6+
ajksTumnh6zQN+GRjrRJsDo1jkNhcIV2eBq+k2F9KZIr/n6ZpgfwwkcaxQ91KRsl9e86kun8GqJS
BZ1eyRrKybhGm3/v+lw0P6Ni0LxXc3IdpC+/ixy3wGLbFfCgDWDlBBLGCyig9SK5pwU58li53OiN
YiXH1v/w8O6ZrYRY6ckQDfwG/9Hu+878fq4EHRi02nNB/8Ytuw7lsG9UytwlbXhwMhoG+zNjRtop
eUdOX+lNw59iU4GnLZ7ut3LdpM0gl8jKYK2duQx8ecdfvvj1c+MbZoOdpHOL1oY+YI8sBfJZqlne
yG1kj/ptMdyxT790vfm8pngaAnE/neTlBOOiQs0e8smneBZ151jr/UwfBTwgfiJO3YlJ6+hGf1KD
bdnMt8lfE6JY9W9rgknC9cfQK46oyBYFbyAEHyMVzUR+HTawLRWvfFIKZO3fJjbB9F1HsgTPPOtb
qRmFt74LEUDCCsLGP0uRWrSla2G4gDf35blId9ENgqOTnG9qYjBN+cb14CWddQh8qtAEg6KqcPWA
iax3peBXQQUuMWYs+eKFVuXw1Fy5lsRwIUj/gOXWNxcKxT25/+lzXM10koPW+hwBvK71ukcK58T7
bET+6VcSN2Ddk81Q896B/XbEiBWHFlqV8XMRLhHDhEGm2YrZ88R0b2XSrtnOV+MVkW3KWjbh+Lcc
hqztUEA3DGNp00bVmlHeAMwAiSAs6crDncYN+lEOSpI1AZHUzjhva5WNgcmwdThcpy8mhWOxypBO
8XdLqh1pLZhzX9cq776H/IJHw3AP0XKAF5BNTObiTxKKLFUL5gwG5LbXxr8fb0eMCsJ09RcgGC6U
oVv+oy/9sQHju3LCLF6LWCC/n/Y2iFZfGQdHeJgi8HAw2J5nP0ZGxCcN4wUfNXBq+AGn66BxKL+h
SaJUx1xDI86lhiK4qktPsLcxqqDl/Z6W4Zv8vVt/RJic/6FIJmDwiaJ5OjMu7su1BuiH+fppcHuf
p0hs6JXY14E9s12h6v0c877akG3vITQ+OorIkQevE/zeIirwPAhc1XqWu11HOW1iQbcMut+egAFb
XR3LMUUYnJE8pPg9l6MtgwWpYWQ+RkN+bftKwaMG8/yez4cz9/YiETGqWet3005x0URoq9HZZLXM
/T4b3blfkKAGEPhQo7oT2yeq8Mm25x+kqS8Ab+FkhReZ/MB03Y/HD5l+kvEVd/zT07nnLgy5pHVr
NEBLxo7dOihdZbz3r7uHhqaSjknNs85U9u8CshdxZF6pvGKOAgryticsF0Tv+BJtyKOXUlyc3b8j
jRMiWUFojK5Tz3MbQeJB4n41MAff8vzKvystxgCHB0CAnnDcYNfi4Xmu4zgFGMKYEuRIFeCkuIyo
ZIbeGVK4q7PSc9P3f4leoPrMxIGNyQxGABhcQgAvMtpQfZKgkHAjHG6WGx9aQssShUPl4RiXmk6T
AcJpNHLjB31Wz4bDxZai6WLV0SThVNJcVD7+PtJbbhprCu1KTVBreu5QaW5JAXZVk0TabGsOXt33
PPDpe9dFb1suEHeDsYPF4HSzhjYKH2SgQMxPHI6r3hg287POVWKWjUf0aURou0mMDCSnpLkgvk/v
YBnzummJCOlgDALqFqyw0xAqnZ2q+SEoxkLdRzY/7Yfj/ebJiB+r+FoeTC98T2Rk6Ew06x8Ca4Ax
hIud68Hte7EpdFBfPg0XzWWSxECnXbSLtoD8n//p7K6Ffxfm4MX3d5N1gYD/A4DAWGD4pVrSJ0pX
LLc0JNvXG7IjnSG2kCgCTjTb5sSaAslTrQW1th3CNNp13k1spnESHLyC8v+gI4rJmDwDdMkqcS9v
3JtA933OwBIITIBPulwkKloKkAVqeAJIEsz3LVbrHIenmEfd6GfiOlNrls3uQEtPv8A4q6wg2GSv
VGl7dAdvYRtKDZkMMtH/HZQfv5Dltc6T1U9ZqlkOYHFY8Hpbyy0sPt+EiKNcIBC7r0Y4Le8a27kD
0I0WXqeAxoEG8bu0TNyQgBtZTomlK3tQZnzpoNhK7/HTwxTTCgBPFDdIogB6VoAzDxaUyK7reV/k
UJRRS+vVoU5M36pN6MjYBhG7qk6HZXfY3ftOm1D0t6RxUHB31CGSqiugan+Fqyrj4gkPqnDDlFgP
hEX9e0knbFJGU6QaZp0ysN/hz8Mbc3/drJ82CwjZ4CfXBoM4JH/c0TiH9iaRPVCYfcwOZwMmy7Rd
sTiAJVTecRCG7daNGZWP/eyPflglVuAv+1g0FXIktF77V1I7Qwxw7NiR3MuzA904Jhc5jKf87mE8
bF73rtiNTsCXl6hO4AMocHm0bznzC3qsWTEqMld3HB9rLhI7t9QEJI9W/l+aZC3obkUmXbDyyHzh
90sqKRxIcX6itSNI3+FPelR0C/HdgJzVHtGINuSBuFq6kg2APZx8dSX0RsqTa2HGiyjbo1aUkD1r
wlTI9bTeigC2kaBhX4ev1hZxBHScvBaJufoufRdUeLUd1ssX7tS9BiEf9ThudiLg8/jIhxJ83DNF
ME+BgrZ0wy4uYeAUGACW0QMVTf7/b+VkvkfJvCTDKsMQbNOqOJHAF/7QIX6u7aNMOZyUyBVTwWQ1
YUe5D6yySjH+2nQxJocjXSU6y4Rp7XBemCN5Qm3ziLyEXAkkTVRVneL5JNyu8mJppcG6zplEbE08
kNXuveCx6tcVuo0WfTzax0H18ez+RbZAen+GjpQdh7iGjAgH58vXqlzO9YvXAKSVLD66bQ5C19EL
jRFoF1kplmwxl44zNOV2+vv/YDvdx85O9v3tsjlqypl6URTwilpwS/6ll3rSlwbfK3ZaBjycwZWe
LQoD3tN4LDT8a/PkKv4kYa+5zyOajbnPIiAHvUZ477b56/WLdKdET7iht42fZ8qXVgTHANcp85sk
LoLGfK2lrlhHSnFZY8wsLL/33o4oxW4dYZ5F06IXodK2KTxzquNvzt/+yb8z3YB41RmI1O2ltNZF
ib0Z7ES/Xbui1hJInyBJzi9Ut+X7fdpV5vflMVRb+hWQDOzG1YBGh1eS35lJcOJgtmL1GKoVGG0F
N7MYow3n0o5omifT7f9FGBZ3HSrXX1mBdiG1t/0XbAMiXuQrCx+oKlt7wpFEIX26FhOnEcFKvAlj
WXZyn08JdLVMkE4RV8BmVvIfo3OgDTCB1NcJRXTo4FG40QUW09VYw9ooaJmdtq/1bFsqI7HU8Vro
Z7nODdsDXvkyHo2saoGeD7JgnhAHsMBTZkDT01agkpaisVy5MmjQBgyIPDFl52du0Eiv8rvARQ8l
Dh5bBcvM0D6TLWNOxjk56slB1/UL2K5LaYgYCffHBn0l5Xm23mwlPU57iDWZoSggnzExo4Jiaj7c
WcxKjUOWT4rwXBEG4MPPmdwO6kTiKfPdAWXu+Abf0Ml9hooEx1/YwLoYbGfK+s7dAKX37LR2X6wF
0qkxW+uen+3qud0590m0uFq1zVZ62EBbEoP+SZZhjhLyYoBJCopi0gbzjd8/Rrn5S6P9/OqEQNC+
5DmkcF/qRYaWNGPS/t6+6NMPsVinjicne4I08jIf0y2BVd2COJuODO64bw4FZMNBRDxiskBVwYPH
CnQgXoDRs+N8+SIXsuUcujDXrDHX2mRz3nf/qBDm9Fokd4taGVEP+63ynO6KBKiqaqpqkvivxc4g
H7VE+LHBnU0SF3hD2svhnFcBgApiI5EhMSBzdq9egj7IfVX6WAAY3c/FGaCk6HCPf63pqYvDQh5S
jWjbco+e+6k0lYegQwCJ8ijmtOMbbyWZPhAkyaKkvrSwq/wXB1Jxvtlqyh6IMy+bqn8ahWjxJFeu
+MzFjkiRYOJk5tn+qdSbRXNso90sfxzbQ+DD5Ercs//YpWvFXNxjwWVGmKq8FmFukQh0Xd0eMRmJ
zqVRO3pC6ywU4T9zBsMzUtdmbNsjtTrqH0tFUi2podmaJSwmkHEWbomG8dWfD3PqC+IpMnOzGI2C
F9OOd4/rGBAjrxXmww7rvT41cfWvP1LrCU9x51hk1Y+kfhAegO4RRhPOyN5474L/b9SvKqQS6q+Z
pe3i3t8tuw7ZuDB7c1no8U6J5lKGvZnQhiThUA8cSAOxHA08XkqOXs3Yp2BaoQmvEDLKIshIRrau
0hBSAuBd8XqWXkCOJ7wQv2aTg71d9QEfmlgx0AQvuMdA8OX2TOkLmyWyg1F8N4xbGR/jbiweLNiF
Nt4vRkWVL5I7LOzWyBltMB92y2taXeEjVMATSMaRBkYgIf/EXA00KWL0eGqWZqC7N6kPxBBBSAwV
5g/IAPzuvnCQA12HXMy3fu9Kf2M0dm8OuXNSfy9E2X/cauwUDjGPCytV0JYKQlVy8MU/OINSk8q5
x4TX/QN6KIS6/76Q5EqD9zH3TIX21w/OjTq1gIV4mPYc/rOOKTy2ppEvYO7JG7e68SioknKGesGR
rn96h0+wzEvoJvoWuWUDWfHgwhad27O9i1obw0flBVU8eRPCTfzHombJ07GNgiMuzaydyt21QJrh
rVaNnhLa9VqsOWbQtzzn3aQYFMtMUqniZKs/2yF+AYVzUv7v2/gjh90SXkRVLQp63RoZvjUh7++z
zRNJJVRSO/d+UaFXLv/B9KQqLTDU4VblweDbatRskL0yQsBcHnf8NvPomGqcOkHtZes2Z5Y9p3Yz
u0s/uwSV3uq7iuy1HSGVEcv1ZphXzrOyNTTzQMbCjlXyCwECvGUSYUJyfKKboSpaMWQ+cWGj3JOj
bADefjBqGnPG1bzbWakXaOWjF9qZw+nwDgIkTaEIA1XvvS5nfjB08vha3B22lYQ6ozqHGBwpGOhR
xxXkGCTB4ymPcop01Syyru7Bxxm8UKD5xhadJH1DF3Gr0pyIz38WlrByAvodiXeO+6pGhAz2ctuR
3k63taPqeWJIuAHYFZjaCrQj2pDjUQd6Ai2wyjeOqfazEkkVZ0fB1DLm7qWvHMKSxirhefQsDoGh
3JWhStHCzsWVRXme4EyS5ORMBx4GdeovAF+76Dv8X+uX6fOklYa0vuHDVKF+MbtkcaCYOVK1UBId
U1ScJISJejUUSrRihIrr2Zk0Y2gC4gjJ9bBeyKwRFVGFmTjLFylIwth3WQJWXXHaWahTvw7bwznQ
Gdp3g5KgytSDfHcEYeFFqscKFqjjuF7Dv/emcLUsWfJjU8H1EQQApv3C7JqLSkckKFpsMFfrPsmX
iAnFRHUmAsVnm+LoAfiMSsYMQ3tTSHZco7az2k2PfKMt0VRnuxLfmVECeMbYZZGnyPqMQXqnCqDa
BlivIdtyAnGjZ6MX9FhKoPrCLcvuNzfvEyx0dHZVgu4kb71h7qL0rQxxtBLKmlk+MZ5h2bP1r1Na
1JGTBfgwz2gYjasotcBZoIgcULOy4sYVw47LUpPcSpjRis2SpHoBbLvuvfDN9ekm36xVSlHL237d
Q2FwSMVG+ccGuTmuyEegTXFdPupjetNMaclUjfawMj4IGbWSptJ8kfuM9Q9GFDlDz6YsZFG2dQDW
wRmhUuM5MEagD4vllgvXf3gAJ6H/3gR28KbxkhnNLUsQ5/wkzUWBmQYvL40debZ83FeHCKxSiMNz
Ia/tuhNFNFudcookZpZ4CaKIx1VJ0iS6PPNvoBAsa5o8CefqB/RjSrDnPLyFKCcwWp6OpJ3TMLAD
7J1R8D4D9Eve3Wcq+bvewqPcf4oa1Ul3KpMBheNLOLwmP47aIZxhYMKCTjjHhLoyOuWOkvQl0SWE
3o7b/6jPDhIa1F3sXSvCOQpLTo5myLkyj+SaDpOUKSkdi9/1hjL+p295a4dvTofwRZCqkPfkuB1f
5csuQVjgqQrkiGtdqStkj23bD/gsbnqqAjw98uCXgUUwRrGjoFiy9Tmui9HlMT0QHh0zm5LXPGEG
T36+fa3dZIt96XF+6jNy0rmew86kJkpPsHZtJTIyMQA/cqaHUexheY9H5dCCn7gDURenFCs3dKIg
HBAoM6s5QeOCz0oU7aOv9Hej9/tYcEndEz9w+QwqgCWEPxT5hEjTpZfK5K8dYG9eENKRznQyWWr2
BxT7j/kSbHsKCcT3ju2OQZjh+FtE1XjUQsreBme1/PBXG6r0aJhhHE/OMV1uyoafRx1+j1PLYh3g
X+yhfaQOgfEkiBfiVLRqOTCah7o8W6hnu+NjUmtNDnx4/OEDt4Umw0Ri3qmdigeoesL58TJWxXFX
AHHuBU4pO0skVn2juDvelHOqn83UdU7kX45Wu3g1QwrIZ5CNWAj3LS3q5z5b0t/FBeFyrwvbCC7u
Kq+GSG5JcrO0vUI4cb09efg6Ut/v3Rn9IvrwFGLVqQqiB4FMQB0jBordODAig4MzKqzHnJy4NWXo
n54+Beq3Hyq6xKfJjah6/eBTefjnykxkMGvXZCPMv2Txj11jJYU5EB1SbS9xSEv3oBA/T7w9mx+u
pghqjE0JcliCzFhntHDV95ZzXGkYuyFAAs3dqovl5RXklC4rE6PUMPK25w2fR/TEVeE/XUgiy8xE
mDn2b/jaXwPIsz6DXPFHHLgH2WdQPN+PGa3+Shg0qrcuB3n9wD8p+XP1+EIt8T3YdEVpBLSEzj+9
3YnX4WuCStjSsn+TEwsBIGQOashAu4X6IWZBUb0pnT0vhMDMS52G/gxOBlEtZFqQph2fk5LSTJds
/YPBtOsbf2rxLjjy9VBWe1G77lj257nABXgB8hw3FW1XObgnraPId6XHb4atwL5ZCI5ZrW1wlc5l
PyIws/bIz74qbI7cd/xv4XDEPVUmV6W6XcFUlpKlrKjbDabth/+W0uGQSV3FoHtd4VwUBWfs/DKQ
nCu00HsALA41kqOlTS/MTQac3Ee54nUs44gBgsDCJMkBSzSqKYtFfLGE+gYf/2DnK4OdK7/q4hUs
XOkXRQn6k2g2iCmXRxDdbfD0mqwtY3sJZyV7KSUL5ryRDRmW76YxusK6SCpcFJOZbb1IM2Nl/SV5
j3t55u6QTYgYKyT+OJQlYZcLH07up2oVYSLzdDbd/QQdAA68zyQfXw7zQMxCLOuUc7Xkj3Kftpdn
ytxP22lM4oTK59BHV/MtgOu+1Olr6q1qZYhLuGD7D222I7rsgyrQeIxtoSfca6QOj7UDhSNwvTD7
0WGSuGOFJNJb6dI31KH6v5BKbF/9vR4HRKyIcpwHJWpjmkinJ6Aw0bxPWD7UC/will0gVvGX7ViG
oT1udkf78mUAnGA/OKKMTTw2+3BTBJEyNcraRKivhln6c02MnoNIRxdSeuStjwjjIckSCGKTBSE1
UBjIERhGzkulEYcDbmIJpNCUseaKhK1YJPYuB+Dm7i4or+T/1IrjsAUIZ0mr4JbxmBdEy66JlO01
pMbt1JRmAxG0btJaUOYpdjV22/ZYLd7oSqUJBGDqD38UHvcPreL0MZqerbQ7fTHBSV+l469RPPDW
aOctcsLiAotC+YfL7r1R+WjMXEphFsnekA/epfghaaOz8dP/MJJf8BegsLJB0qtplYMejuYx2RaY
7Ag8mF5Swx+VtI50+V352nYzoMe2kLn6skMcNRQ4JNXhjXe0wnA6RhA0382BNlp7e2tYVQXTDgbF
xRHvA6blgeicggAwbRf1UyO1bjPNAQVgbc37tuotZJGmgWGFyoROl8zgLwAGd1pYNC30uuCMKVl4
tAmjHHd3EDGGdfPpJGJpzz45c2qyZfhXbbmNjotAQZRAIiZ3ZBGUp3oqaBjJSW7zgoVqed7WTjGQ
hS8vfVYKLTtFjPh16rPwUEpULOLkrAy4rYUagCJqKX/3IYt9Lo/WyMc54rraLsCZWpkLqE9bjClC
alS4A8HHeo/MmNyovPzO43fWNesLQbjJVPFqpRZOGa5izDNrgxdKsRgln5E/lsCkqYwSHEfP7hdq
X3gPpG7a958DzK/wVQmmds8v+CoO0xxcWrwHg0mUTw/JXV7TevnQlwGPDKkSKQ3vhynBYFTXZz2g
TMoC/1tBgaZFcD5JOdCMyMrxlA+H95VSVVXaHGu4qhGB0xGjTuXqcS13oD2uo9RZt/P/QA6OhBQV
+Gea5CdeyAAG7heAwOPZeWPEhSuUvnYCHeigx8BzrshrhOpdPFrBmFxH/bYc3mzgPwgfZjZOFX8g
duxZpbPw2xEHJGPFoEyHktjkdGmS3D4tU/Ve0r1n8T01SiKUjRTNmgPkhq6dsQGByvKjeLd/x7t9
w9LJLTCRaxZsfBMmCCV3iaDwXSymbAl2o1oQCPJvQ1au4jHfMHYHIdzcjNVGcgnTvQrk6zf68vVU
ETETPH/GmIfGZUckmyNijBiyY66yIibqQbj7+VFN8P0eNYy7QDmpVNHPw7tk3CKPcqiOpwK0Sary
y5Q9w22K3y/ITjIbXDIstaNp3EznRNLiEwfBsJTgfelPNHVuDZzAe7rqMfyDDcce/2qUV4ib9tod
8QxIKRNUTPrt1jqpTI1werzFNSedV7md3P1+MSx+rMf5MlFP8HC20chX9NNMmNEpgvkNxfsLQbpV
uadETdgWqEapkL4mnUiQSqOAekOD7itSE4rq3Z/jvWMwogGUOK0f1dOtvrpyfNu+9E4N1euloL39
5s5+TmpzkO2vjf6m9tnGhRcHrrnZY2c+UZY/FERStU3ASu4dcSgbmwzJH+7ylrWfpSdaTwkoQTaj
Ym/aa8neCbGfTNulJ3nXBNOJ7EGZts6YjESixX+OAWolmhjo04KVPqlNQKHNZRAjpEAB46dVO3JE
sMVLrDPQIvjt+MZKw4ouKKUs36rX3A91dsRReAvttW2sEu6bKSuE0xEUmh43jpAMDY6t/XouZ6+2
YBAF6o+EI4RChHEbMlId7+WMcmaZ11HmDu1Whpjdo1wrt7PG7DtwfhOVDGk47ibt6o56C7euTxVT
fUdBLX33XtEE2vFaAgyhC8iynpT8czhuwUfA25z27myipN7TzbYyFsCy3x/iR9UCxy/CoUE0xLwf
x0OhnRXqBrByV0G4BGKC/fhWHoXMS06Lz4RL4z8s11tBfhPrnALPR6xXJp22WBDTn5TysCBE5txD
CrlSGggbZ++PP3adyZF6oumcO8UXpe9OsFyVCEohmyNYpWp+HDOw1gFO54nYC7cXzJaSVcgC2ItI
2iRgrKvv4Zw6n2ZVgIJ546uVXSuy/XjkX291T8n3rNvH2nHvjXiqM6JuE0MMAZGL2dmaeAsKFxf3
zWLQ+tuAPLccVu6VqEZuLr841VHP1wqvm6l4N7bCZFcsUldzW1MbWgaEf989oZXQ9XKpb/L/YBK/
xgEGHiKnKDNuT24I1jcjGg7HnW7zSQ3iMnpgcXF7s3TYDx0vLKO6Km+kNOQxjuWGCu/SAehpfX9L
pEMmhPegJp6bYua48EFngIVATabKjUQIdWFQ8OEOZtcAAWGmTtL+dpo//CQBIez1g2N4ST6I25pS
l11g95luxruPMNJCRjvP1G3DQaq+a9Uciq//Kk0j8Ex1xSaBGwBqzaBfyUV+2qmMPK8Uwne6vUj+
i1g1GRY6+mo93ggKlPBTBW26Pla4Nl0kjT99m956dnKdj45EqaVJV+QURH9DepC9P7ql+RJH74le
unRnIvJY8TDyOtHpXD+hqhTZQVPTgWSAwGsFGykOVB/7Oy7rQXT+NmHBrBXSKI8rydzbX8LxeuCw
yScTsN71tFSfzByd79rgt/+qWgb3eBGeNb1vVkKPXHPeFFCkjQq1x6k0hxTb9qNgbswj3uaD9o3S
paMqHuHFlfPTf8josRiuclEDEQgosD6Q1SEzjfqhxLhkT5EBfIUs7M6Y9r9IHbN8rAt8bcqID7Yo
sQEojqgCAzH8gswpOw99FHgZcrOt7E2dFBQv2OYcYnMbawuv4ZiksVGkgiOz9ujNEZpIDbXBDccD
CDlsy313qbM4ij0hi0J03AgYtHSqhgnsoOLAgwMt2Lg7D17KFg73E/y5MUF0lEf0zxPMpflr0mmK
E1hM8Xw8ooZWU0wzhOBo/JQQvDqqMfeIGW6FsiRfk2o7OgflnRoAmT0l+WC8VOqH0D5f55PQSgfQ
AMLSOQMDzX32N8aAM+GdEsDffrWPxDCVV3swcSzg8gJ1OtXzQ2RZNrr6zikB8mHl/J388hmcShj7
70fCXrfMAn84iVtEIRCsTtJ/C6388IouMJ0Qm3+aq5CjchF6SRrGzf7PIhwq8XAjAfw5+pzwn86x
dyJXG/kv2O4sLZ4Y+2CUNBRwFMz787yYtV6vcVSlXjXMZNvK5YAj0VNwKRNFs9g/QlHZltxZaXbn
F2pVL6pCfdoRvcR0iHh9syoVgmPL4XXCX3pZ/8cUMmk4pmCFXK87gP/G0qjeCQOt1ZHUthuGtbeX
qmLOhDOJ+tpZQOjVMNoRnvSJ+DMDzDuOWFR0HjzG9DEc6SCKbK9aHAa5V09JUDISGVU9bXG3fg1b
h/ZSxDCwF11GHjKoaSDXG7KZTiP5jyuEvsOOf7wdN7Kq94cVRdfZvbqXkhYVuqmurAnr/1Cgb9qG
Etkcnt3+whto6BhFkBu7wu+VF6xAklWUPaLffUIJNADDmN8dcpVsibX5FN1w75U6L0TMzXlXq+Gh
fI0jo8HCKSteYfXUwreeFJp61dBi9S1PeawxYxueNubDtf1I987wQ+2YjxELXxugmv3zTSvKyBkP
c6Ox9Rydz43GKs0k9vARGYPuO43XeM2F66sKNdGRBvpqTcCWHsu8z03W7HXKsSpgOGtX/2dg4x8n
kgAfRN53NKFJ1mnxGaDXhl3cgc405Uq7e+ze06oarUCWwMIdSlNHMCIMi6EsLGiE03asZFT+DFdm
WL4PWNEVEAPXjCNRvN7IUJVpF415+VhgPz1OzZNqxOKlPgm/H1//klDSg1BPB7o9KGOfAqJ3FM5J
6nVhMLW5cypljmMFGPKFTYHlPVq6lhNbX0zbbr4seHPSZdBGgRBv6DDnp8KEQbb64lQGCBtnbdsV
Iby+mWXSB6aHbXIDpIGurhmwxL/L4VHX+xPatnSohBHe3CfoEY6OfEq2F6o2Ush7Ocztl48O/BiU
WxJ03dtFTIsHiRhbLv+b7WMEZlgvMCKFrAxJ9bOCaZA+YYdhayv3vjZ6CAKLtvNtVL89vZwlxUy0
hKZGmBQ2w8uFhcfdQ+t0KeDMwN1AXQLOfCe05Ju1y1hUplBLJA5J8j/Ke/3v8mNBscd9m7+JUv0m
zSmrxi4D+tMMQs2tdYy902IWQ4maDmXSwZQ/eMTC9pyXyxan0toNCnv9kOH1rKZ7JMT2C28vWPEg
hc/H1PodwPqWsDYJSBXa0OITGMkOOKEOsb7RgHXOcc7+ZFfwph9FMXO3afLvHplUnGCC6ITs8xfM
Co0uvFq0uuiO83Zpqt6RNfIFHjAb3zF2jotWN3m3xA/uT5GTCl3pZ3ISD8wgVA0l9/TF6ujc4w4h
r0mAw3t5HozWO2tOlADs9uurMSU7fnMdc8bdwFx3n0UtgJNZ1hfwSf1pLefSjo2zKoXYvyZ/8j4x
qhcsUmcxw1BzSX09eybidtbUEk1ShzS5Dlu7xCPsDvDFNkmqlF9ncKVHjvbdVPjQffcEDttRnddG
1s7cvhV1ZmbcldI8tJOpJZiE/RIF0Xl812bxh5JfEhnEpMASZ9rLTIrXFO7DkDgV0qsoFdzE1GHG
zky2ECJKTHm5oMp95GJvnyTtfhiwRIvFv8RFokdqxoHShNxp2SMesiKoAseBtTCtuDFHDKmXOKNR
G5zrTScyde6VUUNA/6iWMUDcJseEmQVnePTtREUOB4OYPMZuJa+DeN3ZZBLmqKZXca7hQUmRAQC8
D+/adpGtoFDZMYzYxfF/UMqsXPfbjt/HWSWhhrPQTqttFNaRdq9B5Pe50GtIwjbUTj2zVVmk3y+K
G2nFp/mGVRKTwM5c0zlY2QYQwUdjklrpapmYx9l1/td/CALGa4T5rBkI+cfI3FS92nbqb5NhK0Km
aBermbKOKgqDRTGhHNBWM1BiVAwOJFjBWKiSr3pPEcc7HXprZTrCJ7jVRd1f5+R6wGWqAHE8juDD
K3egZQLlQwKcebACv57SxWun9NdSTLc2V1BqJ9u5p9HaCdRbgJrRobOydXR9K+NMXtzq5X9K1GrH
kMMccYMkGUyNgsLBpGH/kL9ghE86LY6pDhIp/Wje/06hfUP4Q+kzXwB3IXtvLNtRC3TaHcqHW4MN
p5uF/7P4FsBOaMjlFe/EM5RZxz5VoEd2bJSs8eryi5RiTDj2ETSLF88Gn1RzdOVWU01Gsryg5moU
kdUG6KEVuY/m6wYEKWLCFbRLnxRe2ktVCzZLIEJ9B8v3PKOMCN7aAXsHZ02Jsvkf5Z4PDItr5280
5cYGVB7ccRsgKYL5o87Q+DaeetnBvvWAj9oyhd3mcAy4DLm7pDZFxBaTg1SEL6K5G9yLejAxmetW
QUWL0YA5D1G5/fFrvG5erzAqPgb0CpHUj/BG7SH3gOqtv6Ln+7GEZomsnkfpIFekqlr8P7Mp4TXp
yMFLLUamvUKQVspFx7Bpf553yqaKsrkLqccksF8Uy/LN9bKaIkv9FZGf4xVHm+SM3kMPIX1e9FH/
T/xRAE1txHUVFLAA5RCNg44IpDoX+rh+oVK++G36vhHnQbmGgia4JK42JxB2OpDED1Qtr+gVVdpX
eluH09BxIJKi7WBFcYuE1uPZsm/qXC70jO9D/hXLXkhqvsWuTGlo4zSQdDMCkHtJEG1TuHOXyuEE
dmqCSNbyayzFYYL1I74wKd1xALMLy3R+lCWjuWxWLDI4tSgcRF7WEa6Up/Ydfn6yTuYuJXUyxuwA
v/fT+NQyEr6/SkMZt21UleAzgXKb33cCeQ+s+TdZWQQZxmkw4zNzYjSeQotoGEM/r73ClY+qG7XT
KdE5nIqJ128GaeAnf9dvtM/YNOC81uN+xosgOGhSAb6NUHNwIs/A4yfq/mWCQOKjAkZCdwkyNKOq
1H95CeHphOuIpnexjdEIbAjB4BtaPON+YGYSgaTHJD1NJdwi5ntwSFd85k77+rX+i91Ebib3OO12
N2u/PmqWFi10jeV6L0GWlYE0XShk/T6kkFinuMgBh0T9SZoP2uTlw041Zrb+ulkndzgSwHNiGVXd
5FP55DDjGIel01BKcekgFXuAWPZaphulJqwuIZxqVWEIAU9L+AI+oAASl9S8eW/1wjInmT7WXGc6
uOwACYA84lk6IIuCMBW2sTzKlnYJSUCCN0w4cIuWqCL8wmPN0iFpBg8NFOOGl2M8UmaO0wqX409k
f8Pyh4mUsz0hVdCW/5sRUlzNRjpRrWI1L4GY29xIQig0VCevcmvXZE2uewnDGygZIkeCuAmlzlI7
z3zeCcLM+A4GmdIN+GhytCWXqv9f5xE1XHVvvFdUi8ValTTFLSO0nhHTjwhwRoGO99rAX2dE+746
T3+0k763s4pUb3KPFPjcmTbEX5oYJ7yR1hQLqRu4QeLQilPF5HVC8jt9kEGpCIA9iqgfSSrJWUIF
RhW2Ob0oeOLUrAgBRS/GjNwDyYb8MKSqSstIBjdenRH5S1i/rwCyDGVQrFFkASn/BS7J2iIBIrUF
ooG+RQlmk2r9+SDK9jelYayZGPaLwXQx4R2Dqsj4xg4Vgdk5VErqcMHv5Be43Ba5+L8uWnrVNIuF
Jo/qm428n3bpM99EOUO7wmy/nngV0rmIoWgKiwAZi8JesCJtPJ8NQAe7JwivLylb3jtdWZpeiB7e
ANBba6pfONks51CMdbaIDpbW78L0J5rWa/kg8arSC6Tav2qpmiRta33ts5Dk38McvAXS6QoI71mV
II3pdxF6gOunJQMEjrFgi70oj9Y40Pvrp+5BeWNJ+5Gigj+ynCt/OrctHjq3lebnLTOAp72VGKS/
d7IAm+/BSVeyJ3oQis2my1vaOBoy5zcSXgQqPNJfjlBih2vFjx5gK8gwtF4mC3Qd5vyp+pJuWbyh
HGsH0QikSG2KpCghKES0oaC9hENArox/wKtjkPtfzJcwsS+tcRi3m1oSOj6obJmalOZdOcEPladn
2h0eUQCCrU5QyXkVQOJ8oUJRops1ILX2blWk7fTVlRGbAEw0Gcpa+JNl5TYrnNLE4kzlYpc23tBY
G9pnoLHVyyXJVMuyjIdxfRyz/Ly38DgDh+zQGYTBbhuIyUf0rWptjH3jFngAdrx8/N1IMyLuKJgj
TJ6uTt2q3eMbI0xSwNo0MkM4GLuI8XL+ZSP946wO6ar+tvbybWsQIkt/dx+k+zpHXhSrVeTRl0Vi
FoaVnR0he3a8wmUyjlAUdLWGtxX22IZONlrkFWn2Ed7GfRSJaI2BsqU6JcpNqIo3KP4lfY4oMpvX
Mtu6HQ40DpMIHaTVxACdLq/lyZRWaeaKQMeXZkPFumegL2zAtAT2T2ZUNuAXEcki3y/I78UzyLLl
53Snl/9XCIJivClKt9JZdxTpPpteSTfFmSPOXtJsdj0r5wzzTDJXf1uNnRb00r5Xnc55Zw+EvG8P
gW/hTET1DXelSs/f03vnTZsShHLUv+BxTrTd7jaOGm8GwmtMlOAp0H27yeDsn6WbCDjnQDTO06DR
83iCdEO0jKzyC+3Zjfb7WuJKw2dF1rw9M3kfAUv3YvR8uGNrlo8pf1WhCbQAZCicOfHKh0DcApbN
2LdDGNR5gi8FKrMorUL5NK96OeOtD75h6ZpJC7QaJnND9suK8bUQGhgEdTlAUVyX3QtJKmmzVv9I
R3/0ePZHDisgIn4VHkiLMjhmUxUMMxF44wo/nmxy0LHvauLfxOcw+zIgX11IPvfB5GHtB1Y9Vqj3
XNPilak6qRsljI1ElI4Zay8wQKJMS1QnEFpcXNbv6K8eJde53v3Fn73Y8ABPHQP2VKJMDqq7l+mm
KrrhLp7M6ztIN48D1AjMEwPIcRFditk1kdUiKdDy4Chj5i1BUfy5AkeMEOmeDKAxV6DeENUUqgj1
vFKnyxpIQm75+uiWRTBWW8R48p9KQMKwsJj0ruOUZrCfUYd1LozGx9nr30bEQzgx15av4oSEi9q2
lzaQ+FGZmcNroJaIsmNRtgD2XE7YDCaELVUvsoic141UoQH7tHV4S59Hnk3qFN8RVy6wfyyBoflK
XbCgY5qd7P3SjJROW6E3fGAiAXL156eAjDKgjfuyui2vplcO4zthphQ6kpSljHK0owitltOjl5RZ
UZ9EmsdALtaaKh8SKsQTtmzSv1GIJ6WYtoMOa4H3XjzprsNp1mYpliGPPUB81VD4yOc0Yl3AmQvL
b4QU9MDg8+3kyfdxSihwHUuaY+wyGtqMOXZe7lKLbsseK4JeXxW7UpGtn5OtERHxxrs+5L0tRFkW
EnnbtjiUon/ftLnjDa6N+YfHKdsUcQmuqmEWemlE1WUzZP0CSUtVc3+r4cRSY2mZeMhydmh8EJqv
7neQ1p9eGaaxg4iCSRn1BBUOdUgJ8Eyi9nc1vhxbypB6r49MeZ7KxBcKED6hUuKYYHIyEx7cw+AI
J0c+Vf60dsUQnnhRi107SCjou+IkCHVpDDYJdm4zTWp1E2W2i5dC/sSNbPdHXO+ZdegULkZYoUMu
sCIpMRbpeF0KPgzkAXp0YDailcRCnWG7QfcFYvETU6zdzquQGPwNnld563zvVRZaotUXX+BPZuzP
23TLimKJdDxybozLQzo1iLbx9bZ9We03CAdmrscznf0lTqedPYi1fJrq60xxZSJfCUc9ii9hEFEX
rP047jBQz1UdFirfLUlAYgH5HG3ItX2Ogx3amsAJVDl0xq+lbWR1j89NLjUqm1H0Q5Ao64sdr2ty
c5CnPi/g9J7m0THnXtjze2YUbsu5MLqx4Ad0CA4eKPwuH5g1RcnY/vDtWN9UG5RmxDKKECoLhTgw
5TPxs/Eg+ohubw7t2YFc8KSSToZ7nvogdSptNRtSAt2xw4lMDpSsYKVNCR7JZuznxv7GNMD9G4aY
Qtki8La5x+5mr9/lcHWFFoqs+JVroWjF1qG6PmCWXNmsN8epyRsyOFUBwEAvb0M6bUZrqrG3vMh8
NpzxhPZAWrbavIKKyZCGGO3ZdpqvoD/KH4Gc9dQwJFGL5RkD37iefVCdvebb47PcMHzJlZb3i6HB
d2PwT56i/Wrkm5Zq1zXqH5YVjD4QrjqrIdhE5U25sERpgILhtX5PCor4RvFtyAg8l+F6tVAZoTrb
21vWnt9hI6gAIorxOTfG0yDOmOBEciygN7QB/RfMVa8QQJTQA8PRtA+ABmjarICuOGYPMfXNi9jA
qb9rU91igauicSuNYDWwdP627DHvErGqJlf3TymOT5nec18fYufnHhj9xjlLYMeG0GL9rlhw8qUv
aRZ6i4PcUnKiH9RqlZSs91aeGOOrArYD9NhXq5OsppFZLESqI+OG04Z5HeYntG3X0xegHJMK1zMf
nTiMHzkBY4Y9YEoR+ZP54C48657psmCM/qFmAvp/xqk7QhZkLfBDO79cWd2uBKZF9ypaspyMxWNZ
NvHzHP9gfd0AzRKz2mTZHZiAoTFGceYbcr78+EPfiWjun+93L0UoI80Ym1Pa6fikqxf2mA8dgFrt
EaqzVBHKK/61CdBAUqQ242VPR17ax1JCyWkYKyelPmY7kP0P8+RKb3kzBEJEYSgQT3sdboOsmDLq
/9XkxOljFcLpAUWcbXHvlJNPbTtcx4aJGqqabhlCz8suef3emM4Z/3FZNIc+wEU26bRDaZJvxw7m
CAVO9YnWi6pee7sJ8Gl8cqfcWwm42diJH/0480u/IMWxyEl0zWw/Xnpu0ytnqH89rgDIwRCfox3K
QAClUWyr0iHeMg1xdKyhxTZmRYC+opnXyEVHud8vL0uq13vNhwY6YkfUeeVbzpDHbzO3p36nrhc1
VfIMOOmJDSaQB5SzHKg+rSfnHaZjMayTftlR6ugK/hlbLLVSk1FGdvfDo+HeUBDspYVu2QqaHiH0
oLoxPUusOAwGG25d1e4OMZCIkkm1G3XTJZ9yEE1KGHLPBMZ0EULHu0FFw6TnawTpma7ioDBC7shR
eCyLx+hFsLrRQ+ywC54hwhI5ulHncqadgE/nG0brvfIHKvCKqGZecKoPvk0w0g65JkcQWHIWDsbM
HgaIEZrKxRgPcUp5px52W0sk/qle/uf7nnEqV/7X3V3H2AQ3SKK2Ka1EETR/jX9tXFdR6ZQCKbus
CZtYOpPM0mGY0bcbkrtLvie9bYSlSn+u7ThHWZ6tJgsMUK+nc0IoJnE3r7hkz93upZpBA9Ojs8dr
iVR387lwf1FBfHeYtHo4+gXJc+gkIoxoKE75PWpMmUAm3JJTTooR1qQy5MrbVPWaIujNycb4UPmo
YaLfL+lnousJX/bGKiOQP1oI7erfT9o+ztdEb3Fst7iL4x1CtxTexK6nkUxsQFxTPGk0pGexAaqf
Odi/pwkbp3K2tQTarxHI6n4eXYjferyTWlfWshT5O4/DDzsdT9DRwvYLyrUafaPCLo2KDGye4vev
5s38rQJ+VV++aJWxeja9Q/x0wobguq4kxkyMPGNSqJcEuVCSN2VZ8gKfnDRVxAPNUlwAs7a9JYOB
GDRjc3HW7HYcYxmZ3lvo1hzjPv60tTjhd4wT3AMbs+Vpgh0OWCRgnC30FuPBGDVWEWqvlNMiAfeW
AvrK3bojzY+5IfEpC/J9NdTYV0NdHcb1Hud2gOVbskT7YkEiAZTj7Id/iyCDKaW/Gl0xnxsVolIL
2wylglOggaWtMKsOEFYHr3M6faHMfNN2ybRLiSl2rePjYTNvJCmxnw1qaWYiVAKKZ/EoCBOnOBU7
WxkdsKeCyBCWCyTlFFm4ZygEve9DhU9Giv4HxO29U25EMRKUllPAGEAl+PjqGcvnhUNvUIF3wEW5
7tRO7O0IE6aYVGtEg6OgoifBfFGXqR0ba9aVkCGXPMkgA+zECDuJoPTJQELZsXGndgtz63Q29B5h
k0g6QKmBXFBElqbTVaB9UlDDt7QTL+KVdDlLAc2l+C7mZPg5fxqZTVZDUNPQsAe14OgQw8sQA0Gg
rhmOn0xor2pfSkHWAczz2qb9TRMJGNOEHE86QN8rlDOJS16ndecJ+4LC92/Wh2upDJvaGJUefpAs
mIXXhiIfbAyt24J9IVlP53zXijj7NPZmreI4I+SqcBahbds9kQHSviG0r+tR6iPhxfQspi9QhJLQ
2UASktUlfQj8kBhLNkcfXW3/6pLIa5AXWInJdVv1JS783G97dEC5/cp51Teh2e/qieVNfz6stTbc
zs48B3JlZB+0ksUhU+hTQcKo54slhoFtEYQ0kA7hu82V57xbko4smF1Hv6Ah1a4xdP0i7YxoruZM
yIhvxbv0LajrxJHwPkQAmWnO5/kFSdanBz/kN6Gt0SRaRrvF30EEyts/4lFoTbIBb0HgFZ/yIS//
HoKK0yIoGhwWvFEEemjf/dk9H5B/Xy5qUjunhVrB93rhGMpJQpbo1xvIBaB/4yyKDy25KTb+Rebx
LqjH6EXSpiFZi8sw8qnWbvbAKrxZkKuBFz0m8KW375q3VV+etdI/GwkDvN8m25XUx44CN5Iicl3l
Dlu7FPj6y3I4ElqUmHtOkhVvOSZ5IsnfFCm5KJK5ilkfIgbFXMufNDev6kXkGwTNejr6N9Rrqn30
IWr2hpilvrVmz9WX4KnWa5zEdUCoblIuZsQMUb+eCXoYD1blqXcxfCVaHkxpbaKhbwa2lMiLKQMz
2DHrMDRHDHC7FliX+h5G61HYH+vYbfMLMaXjmTEQrQ8+V2DdLxdR6EYlUZhkbYzoyrA45V8Dxqv8
SXNhg5fF2CAw7eDO9Z7URvovdv9UpotRm76hwx3tKJd3CjG7D6grjJjTG/9wXtFWhn6ft/nmjg6H
Gg8djeWfPbFGayR39dcwVqbCLFqwuS9RbomZ4MANFQiwlYcMSY+5h4+o+OVdpF1UkqDyk9ZMuKm+
FkhRk8P59BUc2lNGcLMa+JufJH4fdkVEVjpQTfs9Ok43W1wPi+pdl0jjUGqZrCFVdbJryhf5jFpI
XKf7r+73UbHlFmWDjUtMZgOicJa7KAxC/vKk6zJa4hERQR9HLxPKQc+gMPwm7zuwgMB+axADZJvE
Q/M71BoGwYD4YIWNwgRes0q/OVe5pF7D3GhOMXQO/bsLs/YMyTm+y4LzMDj0XHW1zYnwCEQgHTAB
NiXCeqeP8mQpOP42yZcGOSOx0sb7EsepwHQ2ggciJYaBB9e/n+TxbvO+zppPOAIqYDn83zJd9WIq
GxrRONl0CEvYUjjN5Qz0lQ4n+5db+gS1rxfIv4XUmD8l3GUGneK7XcF5o3N6UEk18OPpvSdqdI7Z
kPLwly9qjq55WEdzRkeqHfAJFOl4W2N34pWoOUQssVsYzeYlT6JomGuTFdDpyH2trlKho/ItGFkT
6U8aTVo1wzeua09V7ckXScIHI3Bz/bvRYFuQhNW3oar1xsPJItRo0oMr54KI3s1Geb/cC53I2sD/
4F32G6zL2IHBeRws2RsOJZcVwdzMjAO3yKJhtohCpfALN74NEGJxOgGF+1fbJi3moKGr4OV9CSgn
ebvJYF29BwyAiqhfmr8jgvOb4saC3IAWp2NcIaR/VuGLhlOghrHinCi+dKd4lgw/69Srwx0GJDZg
ykVXwC6ybd5iGuZJhVwQQFbWoMNlIXJ+SHzMRFNUYuC3IzHwuTn11+lIMzXvWoFRoube45l0++dC
hQUrghTmzHP9i/J5KV3xDNGfeMI3/Rs/BGn6LMy6g1Kq1OSapxXiA9c1J/FYaaerPH80M0OP/DV/
r6a+qrMu+wEfI4yhYgzjmFDDEP7fbcLVu/2N0kszSf+u40rpU3r37oEEaLqmbU3D5U7IePANrgPn
uUN9NAIGs7rr8XsO8+eARIXPRpkqMA5iqPkTRqll0aPHuPBTWqc1g5c7cfRl12aiUWwWRu8ZpykJ
CnbdKm/NZjVDGh8y5V/QUqagNMhRw2y7yXddhmRn0B+kuw4d3QGkeW6dnt9OnvCslO5YQARADdYn
XZtOBSixGhUbD6Ertlu/4RuBBKtXUD47aFNK7ZTNT/YuCoy+at4Ngm3ncPFIPx7J0ynIpUFTgTjy
T2nkEP72JmKK+wN4TzbLUDGgKzSeWwYOlgMCDZRXjUS8wqwBCohD4DG6CQP0h+RAL8CKuZJ5DijW
4N3BbsJfeMLYSmVaV/gn4xLiJKrF4rZYCh5aYaeNB1VxvE/pWhI/m0Lbj85vlS+3MpvwF+yO9z6P
PP6/SkMF4+lSZ9YzfYJ59sp2EvgDnPQYWGvBJbpGVmmXJPQByiL9yc/3q9UrN8y+vDRt7udJhaWy
11WfgJ5jreSmrzWcxyDkZ5Vb/4JYyVu/c2ppF/mFZySe3bfpwZuMdU5AsyPODcKca4jGyD6kt/05
BUQ+wIixXNspz3OdUDl2V2X/4vuGOVZpQoXeS1uk9UEMFU536utZpYPK38gXOoahykHV9iM+z2cr
7hHE2H63I0snaYyNR1e96tP/RpX98+yIVK4RVqQ9pQKY5CXnL0LHryaHY9hICuXdU34VSRe3hkkW
DbWz5ytXKF73mmxUA5A9T/aMumkF1+euqsPYl2pSwTozmZnV/HyRA5RwL7sMW/vjjghAQeeILC0z
SM6izxsBBdifKPhtXXHnPZBo03pHAQJeAH2WkmzwUaVjVEtI530ly/M/jHyYk0pPiHFzrZrNNgMq
ai+snkygsKG05+q06Zp8swfFDmTPBUxYqGmrpltTJ8waxLvfKL1vsKRBz7coM/pWB8nSNAyX+ba9
stSc0kYrSBvU7Xrhh7c+bOu9OuY2q454wr4o8Z+pRoUeJHTeO/GgOP8GBTvdiDo0gm0N48/EWrBV
Y5mYxigZFOU8PnPU1vrCvz2qkO/g+IgZ6F8hEVp5BufW1xSif91+PrjlZ068PTeoz4I7jXtLCEh/
UsjTIhO/a6es32Ev8F2edI/GMWJ54t1w8pZSsNbiePXx1B9B1ulWC9LqEXHg7bzo4eaA1VnEWlYe
VSjIkjtvcmJ79VuI+go9HuNHc6q5ODgbFm/hazcAeZKSlErVS4LMsoK0Ap6V6xGt6lRC1qRv+gj4
U24b2lmlvp69v6MItJpucp9xxzOSD5o8C5kyeJjT1v9mLYtjL/5M1qA5AXVolHQ/4Da2eHIzCwKE
WDv/bC6uquKkMr2LkzEIsTTb5KHDCp+/pngxOsIhzgHYLgLFR+JA/fY7nKUE9wX7//bSqWldc+qG
19x78j3P86cXYsiKcHhZVIop0XaQIPHwupmu9RT3oloOhOfjfNRWV5pPvOto9hkSDQxZs88RgURn
7NBVymJeEAWks5wafVVogdBcRBl694Xt1Qphl41fgE3CVbBAgUxFTCFWd6wxza4MtipKOrkx6WAI
8J8NLjyW5mMuOVn/TZ1gb7OnkZV2ysk3KivbasSjMHkBnrQBQAgfKRMcV9cy5paEoa8iO6bsmpBu
lEqywQyg8KMgSMes1jTGkofYHwAi/MLpYHORJ9xDbQfBECjBo82P8YTCFN8qHweUxY1xBe/+EiIi
YLf4r2+6E/iG49gPbzBVaPZBBQoyx+weJ8A6J6XvmeKRg5SzmYg99crMTE2XHHKH7xR/m0B3PkmW
zoHHqjcgpraOLgyyEmpY/PHC5JRQsWYo3vkajkH9eujXdDhNpwslPRLwOg6WUZ4s7zgxy4+AD0ZY
czvsYn3LBPqDLR3C2y0fxYr9QFoHodI9gxdjzU33g0+0GOOAUH7P3C4RxDJkV57EIsnxEJ1jPVjK
jQuW7Z3LISVEr+oYY4uZpKqMrMrxZgSohC0O10ssS+UV4OhDYqaxRUaYedTHwPKF4ow3PgXndCmI
jHgrutYE+Ccm6u3754KuwkJ3XF20ZeBlaApteV4OX9GW4Znw4suctuOqMmzl+KUR3xA6naOLz4a+
RjaxcerITVisTDR+Kbm3E7sr1kbYN0Rgb7I/Pvl/Laogo1+wWxQxf4+1SCSK3SpNhV/rB3q2oB7O
/xLiOvIX9GBlsWBLzUS+ChxzCpChwBT9PXLpXp5hk7+P638/uo8MqWA4fLnBTB+3gOHDOQULqthZ
BxYiXcotKnfZmDux4iFdjJdvln2V0921VHKYmdNQ2onEFc5vjZnA6gD+TzLeH+JyFFFkVq1TUWeC
c1W0r94bj5bV8cmhf8zuOSsjwuPc0ekUiukcSqCgN+axn0gtlNre12zW+VBkqfJKjZUFzfmYNo+E
kSEheVbqPocC2mW2VJURJspeVmwz/RbYOoEUboypEvGe3ztVaGDR+7QzBGtuKwCicXAArsdwBePI
DMiNyDthfPZVD8Bm89TzJnZWsNouKe3d1LyflvAuRb69D0O1XP6PgA3k1447XrmFkMTVvjKykvqG
ozOBK3Al/MFsis/C/H4Qa/+JDGTw+lwYUuV9nO/2d0oyRV+1SnlqK+uLWv+H9bj8aoBydY7SI1aC
4Np6PldceBNJ510hBJxA+8Np8ZR6j+hCj+yaHI4d8Y0cELm1M2dG7UuPG1gZPaVMfNhsnlc/PG/T
uPVXRuu6hJiK/Nt+Qz+va61Fm6tHfeZSViVhb5kBObTGC4H+BajoN9OCGbXjscVpPeK755RXmfPr
CHqzo4sbnB7XJiCEAJQDdg+30rsE0e4tEo2OE9I1BaRO5nvcmCpSXs67i6CuOwSnZKAuS1FS17TV
OOW/f5W4sMv6x1tVs9AXOnibo9bj7mrkY5xB0SjpSPq+eN1LRwSJFJeWDoHJy7+moeTFO0CfyF5N
V0oEfyZhr3FUoyWJzYeLeVXZ2gluRF5lnCYNDOgAKyQXlsJ08FLfo894Nf8yQOHlofBbc7KjiQJv
pgKeD+ijGPXia15xirjUkEhjP65wZvLRuS3N34SO1iBHOttT3pCB81O9zoq7CQeYZbDJlZ/kM/jd
wi8vwI+ksvHebNzLqxw3D/sCZmfZDdBBZwgETrPfiKSK3W7wsOtxL976qz3AOAw+/qbteXN1IPI3
1uXKhzDKsvn3WRUn0JDrN+efbfDdPBguIwMqF8yN+JvAvnw52KXt2mIAQTuWt1lzpFcltfyY+292
P4jl/4OMBVHZJG+2U/yjdlemFL3QhLxQnv3f8Fe51saDAisQV8S5x0aT2awND9VBprHyGDyk40bW
OF5Bzp+uTTQxHps40BzEfp/xfFECPmMne2wjo/wysBhHBWARgdEqm6KyxnfIluO/8owEQXYScuCr
6KdKyebmqPmTPOclQLnbZ6qCjC6YR8h4T/+eTGl8nw5P033ARZ5AKjuRPeUmGQBXIH27QhibavT0
JiykMD3Zdr+ynjayY20FHu284+7jiKHREwaFzvXX4o6fXvvyfg0HD88bAxzzP+9lvp0QH1G/3omH
BzSaq0LubGhWKow/E8vWeVDHpxRL08zF/+fbXOVR/nV+ONnDVPMFJaNStpbg/eFY38oQRGqlZIM/
sGwFhz7GPeXyTcf+88dBu/z11JF6K+3b92TPJeRS+Js6qZCS0X8gj6/6ypKBYfl6fw4V4L3cbRz8
bk2X5cnvAIi32khayOPE2iQNdcaPXvhxlKvuRAyVpviK6dwHznU66ECNtXJxNDllEohwwu3GXsbz
jpkTG6/NrPZh5LaZ31Xx7td0T+sCxLW0d2VRlaeGTDbfBAlExDPJTCpu4U2y8M/EJ8VWxQgBk46Z
HZvArcPLtH7ezoNPpob7pUtYWydEdl8BKgYZgFyVVBn4knCpzNsDQZooHNY8ze0K6s3TNkUh4Cvz
kOMiPGexKrpX9m04roCQBllUbeS0RDoJBs+PpEe9MdlsKWqZtQ1frCSBifpqG7/oL9ZYIJ+jthmq
L/1RjymRgbwXFQDk5T27ajxNJFc8KwH9PLcKJl+OXj8YFUJRaonZVRnDIuzJDPtsdpWPYlv/W9kP
J9Bs8rNK9yspANbL5IhAhfLk6ZCgBb7+Aat6KxtQHKhpMRJPe1sfn3EDJLf2S2EZwhyco1I5aXRc
Pk5P6zzqxWCuP41VQUs1Rksoa+PtQdxWUp4iLIuz/PY+DmCGuOAtZft3S++KlQkKSt9sWSZnWP14
bSYZuQjH++xtVQ6F3GKb5ikwR0T/CpWn64m6+2+G8JZc26ReY12QPr8P+6D6Ass57okykHjtVNdG
mMdi9OTAv9H+Mw4vNaKBGgqvCob1/xTQ/y9fcIq+AUI9d1GII5Pfjfn4L5LwylGR30YBLPy4J6hv
E/rUCkyb7Vgewq+2wsUhIJJKR7F4Ltns4pl7PNReeuoghBPeiUixiCslREDy9uBzm10MmsCh83pS
0pEjnTfgVtV3GFFDVrg2INL6IE3M5lTk1+3cpojQBTSyZeipRS8w77/hKun1Q5U6z5Jnxqyp8fHD
fsWuWza5ovIYha76RaAhddwW6CzuSZ+Gbuv6InntnvHjiSSGc1UN6wS8Mk4qnK0vr0GkXIpdaEM9
zqJr6jOjRJ4+Gew1bOCXBnKtZkq1MTYS4WRCxHi7GGKqmnTODbnAJusdWKkUHHDp1tZyu6TiSeVp
AUibXkEsAoHbubC9knCdlzpn8C1lT4NWnW86XUNczdObrIJd2ckfPPuCFfb+rJYE6G/8LMk3ARzE
+viT355Fk4BuVkSnq77YqryLEArM/PYCeuHoma/A0pVyIupSRODXuGb3hyaY+4Ie4v7j52PkLOxi
eL6Gn3AnZrOSlRkDPsYf1H+OP3xMjJCNrhFH9AXwRqN6/vao1WS6HJO8WqzvCQ9hw1V2dujQDxxj
+TvndA77QvAKYtv1YV0Lql56lTAko4Qjy/pX1jBrEcwQRwX3+2VEToX5ggc2NPjmsbY8BlbxGml+
5vWWS4EIVh4JKErT7X8KI9Zh1sx86sInVArTjYahNwB64vfMIikmr3PN9CIT211ACM1soj4juijg
lLwTxw0HJGqp0lzjDysHOkIT4325Q2odzCiC32vMPVESznGW+yjPp8bs+fv3XA+9UC+9Ez8s+46B
RC9GCL/oQBs5RKGy7jOzUk8ByLdwsqZPWNKnDn3PgTa7/NMN6A2WtwdHbV/SzeT9hNeoX5oIIV86
ENXkW6uJzVu18RZuiavKsaEikiuRCyel3yiVbRap1hp+Xhed5U/D2uHxrxYm9zihxr2ZY4wPHAzS
hhgzzaYTtwoVzpFGPjydhX0vBw2GLGyoK4n2wFG6epEp/SbkzPJKK3hwFXotEw56Y5D9ER8uGwtO
YjaNUI4lglCSPpabrrb4Qx4pfrlVPLt2Zq3KsILhjQpXQ8WrDsn4nJGj+N5tkdoczm1EybNmk9h7
ForoGqHPBrGpqmYzudkf2bJZn4opdZ+I62BfPztO23sAxHqrxDUMGHa0/QJ5HuZ3ucTU//N5YeCP
GrB48bSYNGQdSFCJty5cZfHHsDwuOFbPpzwQJ//7y/7Ky6qIVU5WO0hNRjEi0y5hx1Q9IWWKKMvN
8WSg9LOlNxP8HAYk3G/UK8Ht5q99Kah+WRzy5mFAeDEnHi4XWwWvgIZIfR2rhtMdnjlZPEjrHGzJ
3pokcgkLS6CLeCMMzUmaRHPcRt2S6CZMW3NRxCjY5EHsBQhUa3WR5IwPLxk7vzXE9EpvRbaVE2JT
VBbmzG9EYvXz6J+XcYIJ0hwKGElvf5t8zBwUfjHs/hNwHjnlZWP6CcLYxw9Sn26I0V2n46xSpW79
GWI6vHpivJVa3e50ka5CJgCQBhkBRadaHdZuXJ7yJdDBU5wEpYu41gN5HBlqSk+nOzN1ACYkZYD0
Prx4WgGbiJeDl4ByLBfGQjkj3u1QoKr5raLugnS5ZDZsNmsA/lLExabYBHYTF6+gFyauMmc5dFz5
VH6idBUc8Obm0tnNpHJ383VAtq52zP6u/VQI/2FIzuSAhAPShxz9Fn5eDpgRJTd1N9Yje6OD8tL8
WvhBHHEbNyn4+tV6djVflTXTCMxmySOcDseh7T3PgYOVjOHCPjzrLSjZRRwPPkMGIsykU/bwlcRf
As3zJwsN5WWQ8VB76wcuLxOg0FS/a6MV0qB1jqBdXxIj7WgtYj0q7DYCbeMbWFxl35zfgq8zdq0r
3Ov1a5+kxHZdMcMKkykoWx/ZNPposHK47I1tJP45koQbcDhswgh5TsbXGWwGuH/5fT+CAs8XBjWX
26i+gBNaxJkoCz0rHteUcebsxo5cTd7WV1SSEApfFBXMENRW80JJb3rH5pY4/Ib4BpXj/cdoT6si
brJi6mX9g0jyaq00tWYoIafu+6yATlZsiSYBUPzVxsKs4ro+mCjI0aGeW7LGltMyt0tih8Zvnxlx
RUuAeck3aSwHLypft8OJtEqlYNGddkrGVRMBxWUddutoShSrYLSWgEuHuG0ivenupah8t/p5c+cr
pTuVCYMmVX+AhTl8FcmUUCYX82OjJW5//G74A/b4KnStv56/Fj8EPwI3g3es5kBicYCZvuA5CvQ2
qZ4UpXv/3xu4aH5qcENcXtanNM7GsXByjaD+pdrz7pO3a5JRWv9D0VipTIvF6sELvX4v/ITYtD1o
O/S+Di0z6XyQnbjbcTjJOokyGT1JsMuurEz6qHCwTxZPalDlkpJGQtXr/MitdxS2y5kMgcf3WQ6H
dQ6ilqe93kUJa/+L7IOgabgT1MMXgHcfyzCg9OV/87g4RGvlBIzwA/Nw5bFUanGT4JhrSv3imoId
HMA91UA/Wp55GyLRGoyxHhUMRUJBXQftMV9KOuxQ3D+AHECzOHus9hI+4JemnjbBkxHEXh3dETYu
xBFsGEhTbb1LGs3QhfSenB+kt9FOoefcfGzzRLMKyeU6BgDsY6pRkdi2AYvUDyAtrQ4BGA5hNMUP
qyQHQxlCW8S6u/tjuW+vz5q3L29KU0NHKHgPZuZDKbbix+M4Ecj6y89xfvTGG7HyiCncVuOqC92S
6NEy6d+qV8JtBMEBoyrfzY6qsYW6JmC1Nb0b5rD7fRFg2Xym/9ALSW4NKw5YjxR9s2bwf9Kk+H5U
nGUZnHULdiEjTpt3Ns9dgIgXiQmXEyJlgRwX9jL2sXGqrIsm+i8ebRz1CtucXgx92siP24e8BB+o
CaVjA7AHKzH5/+2phQO+9AK551S0seU3jRbDXh7k1XMTCBZY/jPx0GXq6cPZA4Q1WFqChWi8cIvK
M6XtPEBQ4w3ZVIhsGFZlzmHGUpkSqHbNQNkLO4xKW2x/SlpwKYpQd8n+E8213jojs9TIQD3oq9gT
cgzj9huNUNTpIx++RCllA5p3yRE4H+9WyyD2yEsvdn1V5TUaf9jM19nJIbwjAvr6syAaEqGe9CpT
+dCMj+68bhfz6bysM195BeDa8zgznO9ZIOV50cOnnnHTvA0rzDNnVDMD+f4JUm1yDNTlq3cIP+kF
59eYSj19QChHSqdBYnAEyLEaIlLY+anZguC0xyVC3Y8Jnayrp17PsTRbEaiW46Dr/q8ng5DfGVDZ
y6VGYQnlxt3G3fs3Ea7t8q8VB1TaAkjwN/iPYmRVOCXgL6UMO7Tmf2gDGbvCZYcb144ZINeQaGnJ
qtqA7t5erX+MT0pA1qIAfp6JPdsg/OQgei3zqt5qyTJMQHWqh+gqaapWDx/6NTMJjvc17Yinu+mK
VwyPsILMiX6FonZ/HabNkJ4h5NtLp9STSWjFpBPw57Z5r/ylhd48AYRAVGQstoxW5Ov5qZrHTV8e
xcEFEq/CIhWBUxYX6KJTB+qSd7cUMFC+ph20fqsQPx9In/V+nA92IgyRq3RevdUMiJlv+dWpWcFD
T7PVQq9r+ldXyuuCTZ9pgieU7P5JvAqTKOYK4tq1hMg6wdyomGCS945BGjto4JTGx1wgrurGY9wA
Quow7JwLEZpAvyB/MkwchQfmxyLIOw0szc19/Gs58q5REVR4mvSypMwJPsBS6fMEzkUq9ANmQz4W
/X855JtbHd0MgyjTB6UU6/Nw5dvAlpTts5jHKriYD2Xy9mjq3h/sz7yG31zXfHrxyrNLzPtr5/Ru
cXN6gVRRXaQEsr52UI38iMdSLRpjPxXuJ7XkviZ2BgPyTJsL+cS6wp+uzYGq0ffwL3c6Am6RaNRR
Yz7X6ypa0qzgezORT2f/USyhvLeLcZoYEd/32MIRNUfe6HhpFukctWo1DsegT0zslGH2dZjQNKV+
aIO8trA3+nqC4hAuPBrGS497T/ySFyGvcY0AN5gmlnZhVDwet3YVVzCReSiH/Jo2cNiOY4gnVHCE
8XR5yyZClSOQMMlceK3eu5qvS5MC2I9waeyvbiBuOIDFqmJyEUYS33fLi29XqpWNWlN8AWnyYydV
DbC0WdEi1BuPcCCZCCrp/Eg9CS6AkmcLR8hWMKm4cj3jqNY9gSdDTUhZj+ntx1JX64gc4bwgF5m0
kzgNGiJSuOi+4LoQpNwm8zpONZE0S5CdkihQEFHPrxu7DBWe5DC6xLEx+8JHt1KJBCWdUyVit14c
4Wf1qQ5s+7x3iq13NtEbadM0F9YBp0SzURNNRE7ejhby/REpyHsS3Mb3eaTpGmmuESVIFYVtnvA4
JFyNGdKY4J2UkwofjNpXX+qyXyalu2yTyJQrhrr4O9m2ZWmrShfIapb/iuKTIoUZaQYc+xtUfzxl
8NifDcpH300cDW5zQ2N5JkOBgfqcbwp7G3QCg8trqufDJoXo0+uwOtJledVLOkw5Imue2ygOBrqu
cwq+7DLEAmlMwb3fpjdIwJICpy/W4wZlxgEtpRcE7xixRRvVgtMSbSN80lHIUcqgAVrUuSviBFFD
zaP+4pUPT12el+04i8g97CKLRDM6O0JxLq5mYrvkgVyawIPcOUePFgbJlgpjyhqattmHHCesDGU3
poEK/agV2dhGqvr32OpLMmitYCApTZf+k12L3EeQy2xQk/iL0rp2ATFJ8074NWW9pwew7+u74+iJ
c9l2qhiL6doG0aFssbWJzCWwymaSDD2/Io+0GYTiwm9lf3l0IvH93QexFnOR2Q4QZXwGVZnafpCJ
/1dfed37APtzSVc28qBtIm65tRCJXnoKyIMp0JhH/dpRgONmw0mfJtwbfHFKMvyKEL9qlUxCm/On
JO0NH/WKFnZNcv/Xk1gzVhAkmnIiwvkIYNWG442bj8a7cPtO9ZZelFfG/cnoiGLmRc1G59LOB608
AFzT08+UBmJaEb16gb952chzNQgNlTW0S6CTf1FdwfFv9WMb5Y69X4Sen7eBTJ5jQf1hL3sXCy4o
o1Uk6ZqNvvoXNjbeKLqLQwWxC14/QQ4KllbrfoD4ON6TZKwlah3nXf0JAfi+Gw3VNM65nM42dLOc
rPNRcyMkkhbNPDS7S7JS3b9zxiDZRujzJQiv4FQcci1bmbmWhmlgmwtegoXUmaeo47miizZW2kT1
BFBHZjkAmhz1uJWtGdLeQdCYDvIjC7fWu1JUbU/jI9OBVVOxCwGqOPGRsih+N8hEr+oH7jQODKR4
IMlUl9E/Fz78cNjGPugE14Uiw3HFO/U19yWCbkAwd9akN/VHWtFhLvUQkdI3cwzRfFZEGQuZkRq4
1jWbtBaoFX4xay+q1PPkwRDzAqONKi6SrAwrdqlWlGFZ9Pdec24ZQ5ieHhlU6lE/sFMbcMWbXMtK
p/7L5qanpNCZAixYSD+LjGGoDQQsDG1CKfAmPXv6Ifttld2rKONVRhE0cqboDDY6f6snv8C73Wi6
Yto2s1A706WleWN31GRpEzrciQJh3c4dt3Ct9Y8dyAYZXW3f5BFnWrQT/ICTuP9BpSrUNhZThnxK
1hiS1RmIGkpkj9lp+S2jLbYV7j7QQsqsHVlNBLOzvSU8SnYcqNWdcaY1vUxm2slmgU2xWd1PRvNE
PMP6yvHTNzExgmdp409i+4B2POYwu9pHDBKXN4z+PnmPWsF1z43fN35uXIo6DIP+ZXMUIj5tvArz
ecb93c+Yj8hE0Km/mGbkMBetGhCeyiqxskC0ZycYMr0fqXgDKNCrFXhEjBS0nZIDkFL0xCRmomM1
DvHkbOI+fmaybrGLiPl87cmFuan2IfWBYCvO8I6svz8o4wfE5OzyCtlAz1QDmVbxCX2vQojImego
8MNpPZrPZzGI/zg6jND2vfcPRT2sNU06GfnRtMn0car12xmZ1N7bj5a/816NPNTIc3qyINMc/Xe0
OlW3FJA0k00GAm+8QJr5UldmqPVKtx2C5jknmsdde+VYnmWQxXaJneKnuvxsPvAo6VBD5Wf6ASpE
/FPk+u+TQMH7ulzl9+Mo/OPIHN5Mw7lvA0uxLwN2XWhUARkMl2TaTq63k/V1FjCLZgbZ6oSCS0TC
nrf1yY9qMfbHUoqij108+1WBk9gWxYkEGqk5TCmJmEuNi5gvidP2/MmFuEW7NYwzoLxuQplyGVoy
SQGG+EcljNvEF2CZHcg3IHeZgQu/mfEw6fVKd6+B0IpjfaKA6cDQ7BEw6sX05ixK+pSFQ6ebPYro
aiK8Qt3nyuy2ZznOBRZJERfhH6lGUytI2pg2oDvwTRFSGFguuzFEYUuUxM0blaoSc7szYNdWosTQ
S4gmulTN5+NkcmtwrfJ2+SzHG7gqI1l0cP24t4EhubfT0qtupdTQ22+Y7UbwVYh3oU3uc2QNrn1M
mwLqzbyAwCsURm12/di6pb4UIGOM4AeqX0QI3l0TumH+QdfFWIeZ8HuMagpGs1TZtkrxiq+kBjcV
6VUBYIKzfnGHVY21x58B/9p8eywWVR/VwMmhxGadkQXY98MvdnDHnFqM8538/uRALkMmAckx96hr
TsMx9CNjG3kwiwAX9dpxEMJaIhVGOsQSV06SmsdLsAKBHPicyqs6aDzD33vgSApMA9kfTL2ujfC3
JCMqS0KhRA1El0TkSnOMjgHe12qF9xZ1gQFTSBq5rJxLxjm2uj3FKmDCVsgp+hKod5L+fLoQkAba
PDq+ZnAeVNWuYqO3PQBTWedNy31Yf/YmoHVicEPe7b5oDoK/GXQOGcLgu5w9EQ6Q4UF/yIuGPX0x
YiyLZCWAeWB6kv1qHeAQvqccu1oqeMpPmB4V0vhYf+wnTlmKjH4ZgDDMx6hL9DcvV+v40FdgRfQJ
qeNleZKKik0VIWAyGbND4kBrwvF+V6B8biI7Mi/715LH9Pt+Y4J4FHz9KfOrdjtl6HBNcHKvIc/t
07CUPas0fIBtd21yeONTBikRcmgHaZl9VYXIeBQBnxf49vtT7NpkdYmZ/D+LZ5OGQb2LuNpAbIVS
8Z41SkxaGzI0dEh39CQBXpUQEr6dimRTNfdOA1RNws4wQr+DE7UiEm8Ll+nbelGU6TveoYvkmFgS
UQKu6iKTx9Fy63RSPbbi/f70uklZKTjmnMZ4LGVaz62jI/OIYnigihPh0ooA7rav92eidPRjBAyJ
bsjrw32APvp3dOmZkRwrfPqIF5UCkWYrtl1IksPTGDv+Tbqnjnd5LAi58zqBJ3spsYvNt4tKjSi0
aYiQ7TJJxu4FAp1gBIpxpp9I0I0lCYdjV0dctw6+gsAnOiBFYOftJww77A16XoRCSaOUmLT+5PRJ
NWWyMDAPTR5H6yTvqtfBE0CNRIgula8UI9Z6vM/JW0yJF58esPSfwRedE+RcoWeJVkCE9S0l36ws
EqDygc7hR54bnGBWvqrmslUFN/kswiAez0nD2yqOAPAfaay+gzlEIG9KmlnJfrS60vJtQ30K9YNj
x67JxTRKk7T6Yer7AawowqbRSvogwG1rnP1INiiB4ANt7m0nxq2qAhB3KoFAzDv98m6GqBlK7dHJ
FlEw1rHxyzTrl/zJI6zN4WkiRMGM2DVMh7/7ESZzZk0ZeVNUSncfIbvyXf5xkBTKS1Qf1LlKvY/8
W0SqZm3T7X9KdlJ9T35H3WUCR1F9d3ZmBv3gDMrtsIe+h17+P2f9FjTZ+3NSzsVh1smcbtw+QNVC
hD+MRrK6SaTVD2ayhIX/BqK5ZGUSeJBQsSB6JwFC2PZPs3+WyTsy9dzCG9CqytcuKtopnRW50liW
dgmtMiA873rSbdqMBGNG7Iz1yKMlP2GkWI63wMuriUCGCM/wFMVqx6/tK244gWma3mrXG7xRPQYP
0KqUPLK++0JqEr9fqrJSI45ZAi+u5bwegAnK9xgKPed6fnCT0HiR9YMkQif9lRXiGuXhxinEQYBl
DVcElryX/+J74L3XLJogjxvxQqY22gyavMvBcCR0+GvRUF4JuhEypd/oU3uYRfoeG/3wRrZtJ6Xv
wzL+7pe0ODoXdQNdN8O5vFDz+C1E4EXroGH3iMxZ8lXj2YualrNQnqvf07xtxxZjFriwLTuTxObY
vHvDe1LCuZCpxXEXblN+gZFDZUDIt+Cf8yDP2c+OH+Nv1I4oKViYpaB991rTF8Kz/aJ3afY+qEqH
/eMkOTKUogj5Ztz0YZ13Qq7y+7mdqwJcEBNPN0T09C3avWVWFKMVjF9KMK6cvTFiTV173oXL1afT
QLsTgN6i2ldzFeefsj5C5UxCNfvWEygllum2MmcGDXqpIZWh0/tCUQaviQZbCXMu1Q6+PvT7LgOS
jq6PeqjIqET/sWi68eIBFLUkhdlXEb3zw+Tk5u9/kVa32vYzPOKk5RxNIfqSdAHZzt510YK+bnTI
akWC9j03ORo2XfloICsVV79wUhPTx+T6lkDJ5Z5vxxh1lM+DJxiSwV6LD34tv4XNYFzqc3Ml6L5q
NhItEQ3IVdsKQqe6kzC4FgH3011M2yOEgF8o/qx5Kh/wLexZMoBaqCWb3mKfBFJb0fAZQIL+V5Uk
FhCDvYvHSKe8FGKq++nY08bqsIzq1O9I+jE/8idmcvdvz06aVWnt1vogrHUgNCqBnBf00duL9gm5
pcNaMPs8Ne8eDSCsxVtnCPITthDAJtuhH9qUNmAdTrD6bhw8OtxF8M9gFF0var2QNZ3Jx2P5/4pc
BqW8FQUBw3XI0YQxPMtt+xcn/npkbpRebtmDyR4KuC7DJbglFWohVJa5iHjVNYBqbsqnIvcU08u1
LPrYuDJ7FM18FajMlY6uoxEq9Fjifgk2z+BwMu7S8zApzYor5wmiFu1TQAIrmpO7KFFs6je0h/nE
/qUv9WUPf5aYuDZexQEzwowfbzJiTT9CvuIteQCNQa9urHhJvx6V6Be3aCXYKIbR5piPdxvy8sXs
eOGr3trS4VVPNqUuRh3uhC6t+erf2BaQ2hEEw3i7sreTai1rqzZntTxwu6XnK4phTw20bocwykRD
oMnbOEK6NX6bwHh+FH4I98Z8/ALHMZAc/LlR7EZvixkFovJr9SpkQq+aT/++Rcvkz6+/kCwaIj2f
OHZAPn2UDl12ge+Ds3jgk6qReH1LBJfVTxd6UgP+RhaE+40v3hjG+QRBL7hgqCf305VnCF52qwc4
1CawrrzuocluZY8jF5tSE3cft+QKERpH0VhS32/zjl5jx8VipKLKkij1epMK3yLjE8KU6mKH7auI
lYtdbN7ctAWRGl4HE14LOm5XdLjmJUOOJMeXaJbXpqNylG2+kkDpkP5bq8g5D05XDzKknUlYOADq
n0GuMS3zkZJJjEjZBEmuvaBLqQ+FORGrBej8HlmHOaELjE+Neo0E1vDIxUymltc0U6kriRZn/tNS
yJCN83KZGdQsiVKRHM4t/OLnqqrlaZsVYC1cu11Tla/BisT8av4GWOPwXOmROwvpxjSkuUhyU2bX
j8CzgwI+e0VQayNfOYwBOXrGLW8HK18ndKWyxUM29oeByM5V0569GD0aUczd5H76xpeQWKC4YYlj
pacoyBgcqOeeN/XPZmmaXGl2UPZh/p5WyXl4ZQM1xcrtcUrJrvRxkN88tIh2HHuOn6bm1gcSt5db
0CEl8TGP71YzyTqY1kcz0qPQej3VEqZQ10enjsUQUOxNdQFEEvbvV4n3/QjBAcHhYagtbOxRKplX
HbWWRTMHezRLSi29EKYZEb8nNMUo4IGcmS4KBGzFugX/KTwhxQ4NVruOVyuNp7VZREoYFhMyM48a
yef5nx08YRR5jItyoALoPVZo57VU2e2lMUt06Q3ib/sYxNH71bvOAzv68rOXxEiES+O57il85Qcd
zob55RBCxjKjdOZDnoD89DHkE6NmzgKSXx610byiOq2puRTullhSKJ0zIz1fiSOYRzBCtZpmGRiH
J6+qV5BKRG6rAyM6xeoL5Dd43jvxh0YDRGKYILh8fxkYAwD8sCq/mpLE/b8lYTlCJ3Kh0p8AZZAY
/C8zjdyX8Ue6lNK8pwlpCl+FX2z/KPmg9tohtcRtPDrtysJF7StJ7UdY7iDkdjL5FsCs7TmvojSU
1X2q23d4zVTPSJnmu9tfVBCbKgHF6eztZh+vgf+ELEuLUOcz2rZ3l0QQH7c0+2Bxq2VZfKWkOG3S
FPPxDazw6Y6EjR7R9k8XWAuIidKwzg+AwI1+rKWzO1aLPip73devYiVs0Rwde5pIE6CNpBQrjo5k
o+sVzr6dtnyy3G9g2UTKaAbqa8D4R43pYMZcapDpftARbHnPPkY0m0cT8iSGGb9qbrAt2p+7nWnD
DvfSwxuC08mpms1vhDSDbi/+br7hWZ46vA9cPq9xv4L+5e/E5+dWuFnBOzPVw6jPw6dVz7OvZBP1
sFvuTEIQo/JPhx7CJpkqjpAXCq1kmPZDB/JrRyAWabrist494AtI6zxmOtklcuFe3qwV8UlHWv0K
xov6v7aPi2PYEUQ9VQ6GUU2QCadWHqclt5y9xNT1iIIf5nGUgKBIN8yVQq+45hcl86TTyGbTBvVh
a9rtTtH4JhuK39wPZrokWvMJ9b6Y83Pg/WAcJlcXzAf9fC7G61ETrKtLcao+j7uBEZE0KqUHqiH2
b6Ao0CpH7QCH/7Z/b8zIRzzAxON6BisHfsOpse+JquVDwLkzBdqTlhpFZoUUW8jXj/fqT7h6WLrJ
QZxFulX4ZR6P7UVI1fVoR3A12BRbKDDc4tnLwdlqZdZDTdWA8ddHcp0sKwyVVYCPtRUmU7LbbN3n
Pf4kLMV4wWREkA7oReNl0YKf07xTk+/k9Y0ACn2yjZF7PjCqzPwdCy5P02UbvnoRPeIu6UJJgW5/
n+HbMqrVOQP9yI1ATHO+YRh6uFAUoz7PZLwnEPdctJRUouzv3cicHJeLVpJ0rehheQPgVi+qVZ5B
sQi+pjAng+0YbsVNtP4ssubzQZcCTtXgWTKVgNML//5CbVMA/EiEpZTEIX2XXPWVWyh0NkTyyihv
k4EN0OrRuYCI9qXxLRUrJqnf9gvdpnE1wYubMDqHFoCm2+MLJVNoN86y3oMCZ8hoX+jCikyS3kG0
RZZDQKpZPuEwPn3fN0lzsxRD4R4Ne/gVAx4w+3+HcOZF+bYAcWYh7lMN1NsoJx5nZuKZXrw26gMu
BPvhqOmMnoW9Ws4hTLEfzec/eGIGkEVNn0R9CDfBSGBIeBmThLy5TO4pmJZTe8IkeOGBhNOOeaWW
IMp/nG75yqcsS/FGelSNrM7snYtJdR9mw46ytV46t3radtOGJKRrpKTuj1n06Kpdmf+K+Kavr/jz
Dhi0n8cF6GNAswycTl7bHW1asldEIi5Zzy7MB2v1A9nE+YPBsMzhwU8I2XIslKsBeHcfgrg9ExEf
ZuPAZ6uRabH1HYaK1nB/Mopt3RlTmPos+JJ0eFF0LfhmFuVDSZ2JkPDPSig567E1k/iYJNIewEta
W+UvuNlIzjNn4tOHi9mmQuuajeW2KAFFd6OdqLGGzM689eumOL4mRdfQlTu+OP1Y+6fT1U3vu3Zs
C9nO3Qwg3bot14WstF/QTVvX6WzMYUn9Jn01PpzKhjVdj1foPCngHMFmIHk4Iq/fPtwbwEzlfQLc
OCsl04WPR1g2uUDIcUl8xB74AWpDrxuJUn25bTmlOp//+wShg+4JK60WXeQ1GK8W0kvGEz75hTaN
rRjJ9X3uzLpoiiW+wv5lkL6cCFwv+IQWkdA4nuh/+6b3DY6F7SEUDZLwx6XiHIW1VqXRShK/HQFU
xFHEtpreQFLL73Ib54zZIGRTf4uZKvY9DpQ80iPAOtwyaV18SfwgYLeF6hYGiDlXAc+YY1K0FGXT
H7JY+fc0EGUCj3+G9Rvzbwy9VCvzOV6jiAN4PYM7PNWnBjDsVj59oM567K7abVziDL59vPhiJDt7
iLaL0ltfiaQWHY7g+F0oAzSR2328DpvHlDPAhImQHDHg95FDuVRJIj+LWt6RiclkWj2B2q9NK+3c
0wAkIB4JDhHzNCplrnSrNY7rkzGT6Wob9aotJFbC2vzAM/F0FGk2bEMaRj416BC26vzcMCaVerMc
uXlR0EIt+CV7ZZBr9azP3AFPtKToc+dcqh226mHAHq24gRAIg5VMV/QSIPxRjUpUylsxb3O0uvbN
0eKdgbkJ3EvDuxRJzsctgcS5HxTwAmvWf3v6/WouuppPMfFCiHE9KJAo8bFEIlcNLpl6uzXhawrY
HnVJQr6Mw8oaLeu+yHPtFo90fMr1ceVrXQrEzKgQZpdUJPT561s7RpoTQyMqH5+6hfzkIT9uWq3N
Su2Vm98mkCIrmZayWMmcRZOPvUgU08tHAgQE1rEazcTxHDqLM2c0CnTDGZOf32gBUBKnJ5+lS93B
gE+1P4zlrfUZsH3qbML3IQ/Wat+Elz55HM1K+1rhlm4VYHy4GJrjK2Gs9a2aBwyR+hutekEGPQ2z
xgsleS2/8j2BNIth9DWNE6Va5yWvnPDXFUoiI0mWK1dDZfJpdHjRETV90Wp2B+JcVxrlq8BYBdML
U69tqxS+e+L5SFp7NY/VASc/QXXAxiMjPcJeAHGSmTpgVltda8054oQXE+bWv7Y10Lt2aUAs6jqT
ubon7xfSRMJDT9iF2UqIHQbumJ/fUTcS8PgbljCLL3mgAwflq06UFWZs9OhuZdo/9sQg3E3Ot4dz
0OZkAkzFtBjeOdQZWgmI098mJa7zq+TT2ImGS8inslbjyykTLynhH2JI1YOzGnlgY1lWholi14YL
bqHT/EZ9YJFXSf+h08AdtDmfTQHPXCdVnPXixa7knR3cdU+irH+3Dlcip8+/tokcLy7MikMOEe/D
RwK+rYEuLVrHTxpS0r83spV8XR+u7NqSK9ja9QOsQxFw9gLkpwiMegwEz4XBZYGwX5HUz86AsVjb
5QMbisqEBBnHm1LEigPPCrhFBTUIIfqqeElPHTrG6fLb6FYqjKIIWsdiTQlndRJTfkUZ3MWpMx3z
oeJP/b4icFaNUdcvCksp1eE03hb7v9sJfesUFn89OuhvQUC7uKwwQjECrU4sU08Vp44Y2PVIny/q
YRZ4n8v/WCK3q4fRoadgj9ENcsSxrUvYKv3klfmFRgFSC+5DYWfzG8dWwlWbERhFEaeOqtLK5ovT
wA1HQGtq9uccUm+pnPLQ8QASMwnCDhHMY6T0DTS37SBgb1Oqg5ANF2wR2pa/xe4T9XifQruMjw2b
qjGFWrxWqqmOskP2L+i3IsVnO6ERJykWkwfhAwFx8qXv3plV8/c/19nLvzp+2Hmxs/kvPfG0fRQk
d2lviktdh++WoPl1CDvReWYcAiOhTVzS8jJtvsi3ksfNAO8xG7/M0NNQXu97+8Xrp1LRlqRcmUK1
sRA5QbJ4k6VgBphr/G1fBLuyPugWiOv10jxZK9oHmlSC/NFP8HrSA/hMjfWkO8ff0HH5I/DB2UNZ
GsrPYWgqS7jtOL9rkYBtGhR0KT5bF+Ow0hkulte1M34sVAcyWNjNutJaib31Qd0Uudxhsoz2TLhV
hpwglK3iCrgCsaFLyNbXM/8LGJNGalU8VSj1/0inEzZ6EgcZwNQSt6D+C1iQyaSrdbf+tiPcI78v
bQA5R7L2g3Zd2P9GjQFXoG1TdabMx3D/CEwpJfKfjvjDjrALrvLpmUw2HGFyucPhOBN1TetOWMDc
JCQx8uNzAmfpZlauD2ww1csd5TX0U3Ee5HOehVkZGqCQFlK5DG4qqhA2ofYTvDku024ihqmx1b0N
byl5EtcgjU4A2wGku85vH8gUoygaHREmdCeHN1x1T/wvwf2JAfTtFIX8IQG6okErTPjtYH77ssOO
V0XoWcU41KfC1CE0X3OXjg5dONzW5bQ5N+pa+YB5kGqp2PL0eJmMIZNZQRmJa16BjLBs8q2hvbHB
36V91OZHTiTBGdBj9not1omH8huZ/EcSSaNvG7SyFYMt83e+GNwxrylz353BkZS1vV7Hyf9/t3Ub
PXVOkZ9r4fQdzMwJz8i+Q0ddtwCFftPt37Tqv/7Le+MLbQMzS927q2xe2cI7vJNeQEN3qzwGByzM
zKeyTHIvRpWwK/mUWR0yTOqURPnAT9K5sso/cPq35lj+01JRFhXR9yWHf1UYUt2dzDnROk1FCRK5
Js5iGy2WGfYMdzoGVWtm81HhdJriBiF2Oxv9qDOb2f9KWPa9UybF8f5nAfoY3mpL8/0tkx1DtDtz
B6qMXEIZBW27koG3JdksI4QKeP2LgmZfU2RoTmLrI3X5E0mRuzlRt4Jp7fvClIDVMkWwpEkwxitC
dPXDvRt71GqjmSLRS+BCda+obeMmV9+CjoxAp6bXYngpIgH6lY8t5o6niABQ5P18065G2zITkHjy
ylKE3BUZ0yCjnfDZjXa0z5HZiO5MUX+6OxFiV5XZedQK4ybKRqtsSffUR4Yw+6H83Zv1OQvzxLXl
e+harxp3Q494o5Q5ajrFJSUld5bOk1+spw2pmbWAkSS4ZnmAlgFBJ0h/TrMGYZyqt9jmeNAiVsDj
ibDzQEslSYhvYrtionQY8YaUhuF9JXz2st3IcfHjRQ87Yc6kemo4j9eoydCpAz84q6W5pX7QcNtK
1uwYEFiQsapJWChkCUWk7fRAhE7TMUZnGO1DPKNPZwbyyjlx8t84KfF7XPWv/jgRDwBT9zqoKQL6
BBtjbGtdnCQOHzQx4qE8RsqfQ/D4QM9VCnvgz2+GTLxUHhZtmu41QV4cYYZu3i5Ap3sWmMsyCdCO
WF5OZJ1Cqrp8WNA6ZFa5D4aFZi8G1iyFzdBI6c5Tje2L63TfqeJm9Ycrf7crRZ/7VMYJGlda/e9l
FYSkYMj3xcnWAh8ol51pBh1OG2dIC5m0Xy7Xbws6LFjjlBoNaYZuAXG8jhS7HjbTPJBkReuVgCLq
Nl1kVBPX2qWT/GBqzLxgYnc9lvm4Gy8/n1PVgMx0Yum4gKjanVJWHXLJ0kupKE3Vot+mvuFSJBA9
aLrNWxfZ7P25+EPhVr6sKIOjtk6KfSTCJaH6vDtuQWyfTC8NwOigjj93JskROJXW7btKdjGfSayh
fo7PI84WaTknNdOmz2MMnmOviyV+af7F+zE+tGh3kll5a/q98SQc6sI0mguFeguM2MnT4Ojh3q5w
bBQAiI75je75UNfR2A8aDyeicAXH9kKCPgCV7tgJ2UNOAdy/KtPQiFNWPuGDF+NV8s20hOIxDUrb
E1MYJN0HGey2T/7R9bv8kbSwHxS43B4zmjVdB9k71yb6iDc7ZYSVXpGVDhc19agUqr7g/3x1Ka1Q
R8fOro1qQrdBXTU6z8R3V/M9oVMPcgk8jTMTy2JugX34D2tUDKhnIwUmnEkLiCTsQ2lT6xJYQkDN
whPDi1QN8dZOw0VO63qY2pslrzCfXOyYgUfV2F+JNahHzMDAnErsgjnwwt83zy4sAQMjJE5WWU9f
AuEyQ5MaJqYqd+umk57n/bmVAVojRnvHVGPtdXgSlUmC45bmdK6vYvx2CXQSDVDEQq0tOd9omioY
4DjhX7uZD9fQoz3ZEuj0QtDTQDiVcddlbLibSjjpfL/F6eSlNhbWcpSmsORBixInHSX7M1kQ2HPm
qXZk6IsepLtwplPLzBRlRWGS3ADG68VAJ//oCJRAHoOEX3ck3j8s/hll/IUWmmDB9/+fe//O3eB6
3ViYyBmXGsM7QjnkA+ckyMx3h+i9g3EykwlryJ+3ysqvOigqINBYCsdAf+53a9WTej3NkzbQVTZE
nulQ987rx1w31gEVTHMH5adLAsRRV3GpiHTDQdKx89DP5L1wxshbhzUDFg/X7ag99+cwTg9YLjnx
Lit3fREvSc256fiTh/82+kTtc0DKJ1UKBAK81UZZXlxOZ2tSpKaEGdY7FruO4i41oYjhHlquDI17
SsHuoEnmjkDWK4c2Bu3K7FRpR5uYFtwbY4hgec4ejYdd2PdkzoWa8AVZ2+ffaGO1NnT09sVBidHs
iIgem72qq7FXaJhEh85Sn4fo5EoNNMxhufoEgOsyibn5MBMWkFWfV04DG6WBw7XWJwWklkEWvjPp
Yv6Q7IeGPt3LDwclJ7y6DwGlRRkiPe3gTnTWMyTWmCg+lGh0kWetP01whRL0dM3ircyyu18MI213
yIpZkAkYcDvV1B4oGUnw7SN0tkKtAUYTHvDKDahu0nVySGRFwq0X0rzPcP1+OuaAFlsC5d3UGAA4
8PbqorrtnjStUg0Lkwh/bfUve32wkBaYqZFKRu/N0IFqFnPHGhW703WVgTXxXnaF+k+9KPHR+iZi
Q3AC0vCYN63EEEwT5bMPxxmapmbIzoY612qgVYqA5djiz0DUtDfU6WPy3uzjR363peGyNHOkZ8or
SOHPMQweQjQArO/sxQHBgg+cfo77alS7GX2ttPXZphnsMF0ye/Ql6emDz+0NAF5huNrIr4ag8cxW
KazFdMbYbR7Irq3L2gkVoAd5CYGoFH7YtxO0Rgh8/hC19U786PbwVAX179UQw4Aw0TRNS62t0tr4
01AuSxRiZ1X9WkDSdogr0lGfgKr2LsAy7I7VznjuMaozRk65QFhAa5rH+pQqjdtzhp1N1yWZhJbY
8qbBTArzws4M6rgAoFMnu642fbL542WLouU1zrkSJTTesX48FA3BTpfDJluk8fgdJc/sDUdHjkDf
UIqqZUIFZto1NkGs5TFedd2J/YC9yuc/ijqyP0kqjnXM1Hendtnz+oUerexE3wcXd6AM1LF5vSx5
54BJmVQQzZwTXxRODgDhEUepEjjuMRmE5a9SsS2fVrTmVx1pWQjXmXRK5ppZsXBBcsIkch8SRkfM
1cIX7xwa1qKMLo2woXQU1LOdSGzST0CMHFxSZWBCojXn5kKgk1FnAp+6S2tadhRrDRnTc8PGupcF
EQMsCSC+idFmoBPcWiHQutGrH5MbzmePgqGogpihSNDyWlgw0I4OWdvhvtyk4QB0KPSz3hFRriM8
cEdTSpDverTJcbEo84hYA1zn4JWdhSXFyN+DkqKEK53NDtT2b4uAvn3h/eFgKlmF7Px7ZxrQSWI3
1qnZzJsE8hPkkne4tcKNhgfKVMn0+K9VAt66bXv5eYWRGmg+glGedV9yrSanopZMB1tPpkes51lZ
/bYSdUgutdZLN50J847hx35yBZOzIU0GEqSjBMFOMTzCmh/8HdaiWnoRPxyjD3JfsWWZvQ7t8KPv
/rG2F0QrMX+HE4Zfzklo/alZOt6+2bHCPvRPHlTDurHUjkyBQ3FOXX00eEKeuzYOWDajdXqr9QF+
A+qHpg++ddnIYK5b3CqT1r/oPvoNeEswQ6sg71ulih9eDdZxfgVIxoFXspye1dDVTPKc1IvEz2bT
FrZBhqR1EEvPeYXDHDUtaTAdx93jyo93qbKF32/ytSEJC7Qalp995MKsNzm0EyA45bir5rGq8Njq
TNEnDoK23TgJY+5DswYuLBb3Q9z9wq1+Pjx+5r0Oe0+Yt5QB8hyEv+BFXuiPJ6umCxnff+7zHWrX
QJ8X3iLoLhKgaGQ+MD+VdNSbxZUObrjGSbThKfMeKwNpxl4MKhTfmy4jdAlmhjqGXInjKdf6bIj6
uFlD+psQAeRUiB3wDGQgU0Ln/B/SOQmUrC6ldltannOl63xCM+JHy4KJOHBhcNi8JLFiYXb4DPkL
srOv/lbToyBpY5D8xfzgmoN9+rp18G5TPnWog5heRO4S/mijvTKikxxm5SUgYFl9N5dGSJOrdQ+x
RnV0/AQ5hAN/H9hv6hSyn1EL7aN1Ed8vvOmkV2Mp/3+EPxJBeW7S3NKruL+KRPqt6whvtHTaJRWv
8t0CJcDIv4ysJfBU0dDBIoaiijUHYuAYtcMELeyDiObQSzAaWc2CpE7VXSdwK6OWNtxhDv2VsIMq
Wh75QuohHx+1fe9C+HoVbrdvQ4QE5grdyREVyRgitzjkdYnylHOQQAyJNSb8355pNHVWgUoOWjGc
pKbQ6un5vE82daYo07OpqbYe2A0WPKmR2udvFdN0fEjw2jD2I3RsbNZxdWkoMzg7zSQdP+3sxP4m
Oo9c9V9pMV5Ykxdarfr1oajqlnlJEyKfYuTDS0HhSbR4EyakhpRN2yLEV0m2cazdKXXO935RfZKu
GjQ0vPjw9618w+xc4f4jvS8EKkiG3xwntuIDSM6azywZwrtwp6fKAESmjeG7xOMJdnIRTG0Qq/lg
j3i3kUvjydZ5pCjFPeWleF1PAlTnyrbnmwc8VgZ51eoTQZdqCyGiJj+FiI4ZPTjDmPGFPwO+gQA7
2WCGAMm/5DM+TUnoqhvswVHHJXsbYjnlzSw4XqShBhXFPEhjrk4ApxmPNV3gMqeqFjDCWpdefz6F
HJRGeG9e75qRVvJpXGEsEYLLO0kyna9q3/pChuTQzWKWP97/Z0/g9RCqjUvCdXbe3A3kik2d8nRT
FFI7p5UPafmyEvnAL19td06uF19ld8COFz0zyXa8Nt5l5BrRNUY/fdmGXrxepZB6COgpexJZJ/4D
iSK/peCyCdRecyQtBkgyKtJs6e4ktAtQF42H7yY4zdS3+BhahV8ttRn255JbwUlt7rPDV8VVvsCB
VLep7AwKnkzJlCvSRX7FJ1JP18UHtv1QvA3aSGd3BEdssy9uGnYUzwVL7yEbsHpB2N/Y5OxverbV
3rlYpBl1GYv/mICJeFgyzRvuwRzmsiT+NwEwJKnSdYlqIuziJmaqWrV70ErxyOj4ztwf+G3GqlMh
HJzED994N8LmXEhVsRvYrolyX/BDBoqc5CYmrGnk27ci3ILquxRbyR2ROaKsucLjfXYN/yJWVKAL
s4EpBVLmCUDKgqmSl4KIWfHc4/LMLlDg8xWNoJWJuEwivwr6H+t7a1qplk3yAN3n3T27TPuhN+ct
B4g7/tj2MBEQDP6CXMQ8ayUgSYd0Fm5r2TV2Sq7vciJ00SJfY7vyakQJmj42NduLBlboGOkh6YTt
fMWLrKXstSRfe2giphJpAbs+v0QG8qgC481X2HK2zVDpjAVaOBiHr41x+wj65QrGRVcu2hzs6CZi
26PJb+iQ0QTnPuJaA8ANiXRXZN8VE0eMt03cNjdFFTHwNKcAImw9IptM01ygnx4gawew6LXbwirU
fCNVsPfw1zvq1jlbY1966b4hcUybZosDKGyfassxql3RTpP9kCTATwYqrt+Xz0qgzr1E3Z+mtQTT
PVoN1sM5k/2R1hOtcxlt+PTMoRE1gEYFU+v2TS1FYvHT81ktSjKDkQZgd7XMV0NHCPML291EYhae
YyNiFwIvvqTrLNXq+zJ/9GK3dNqvffe5J09/xMkYgwz/FoShyc4URZ8gFbkO0XwouMC8PH3V/YPZ
TN7L6rVsTSMAL3vFN3xg3NG9KUiQb9vj+9uS6QpdXqIHnFreCFeWFhmlPwzt8DPnta623ZqqkApU
f03c0Yh7d2ZNDPvgfROKTxsjl4QaUzkI0dhjbZ79CE4It5YYtyLdDEh5K3HMFhHOEJoS4bX+n1T2
sbNaOn6eFOnVeZXRObBo+GT0evqxX+zniCmB94y2HsbC6CoFbu3GYrDbPbXYEup1vm2RUnfJNk7s
slTDZxiYaTN9TCCFx7ReGECbFHDKvuOT7atzKXYdineRQxqy8q5lMIEtVccTFaEgE5eNMZxrDQ8X
tO+9sY2/t55Byai3grVgfIVCEPLU5+gCeQgxvpy+5PU5gQJ7zqeD5bDYDvqTEAYDJYxEuhsBp0IQ
Lc2mLl+Q8J54ZdQ349HEvm202PK3jjdnQQ4pqG+eATvOlzO1kr8k6SqDfExHRo8yMIV4aqm+kFeu
+OJkoOw2MmmSt4Kjk5CQzNSTAQEFjuV3g/Ut01nn3HuidDfuSWOObs5w1IVbyvC2PDEUUXBYH4DS
7lSiCufDNlEVtJ6AUpy5jyj+x6fOWJVbU1SEDAE1jSlMnOWJsP3LTd0g/DLAFVH1SYxCCA96N9SB
X48YDY7nwI0Rp6Z5EjYvFF9W/E8w70mFSB4gBKkmovw7fAjL9iKRoSAH58Ze2/SwebYPv8DsEo8L
n3RXGKLf/xahAj1Sv9BuRr+ehPmPDcHeUofk3H8ocd+zxAkn1dm/rDF4NYmrdedBwAsPAufaBnOy
68j40sFSo4cuDVwgPLFxdhMjyHu5aYySxOQVza0vshOtGFPAWjFb3jxNVD/FZuYx4cSPAmq2a//7
QHheiAMG9kqvRlYc4wzRCNdFAamz8aVGIVqPpkHUsYmwl9qRbVC9WLqvS08YIH2km0/DJRGzkDcN
j4euPGgJq4g3PqQkfLudHjeOLrkS5gYwGAafEaYvI1RZq7rbm4M8nkQXTOOWWwKkTiJ5q4BEH2vS
XeV+5LgVrfZ2wSqBeRkSOlb8YZCyTwxu36Irf6ktlnU3o4S2tTMb/JbVg/Qvdwi3hB+KBm0waf/i
lY4FuEQfdP7clTCRWH2N12Dra2v7h8RGsVtDKUBxLs8ArsZHybNS6v7RYML4pj2xo7z1exl2Q/3C
3gL0Zd8tadFKZBmN4/d2DQpIr1famYzKE8bGb56dpEr5brNgISL2vhxuuUv1opUfcY+OJoUyi+WX
8UedYcmaR7NrC6ztrhetIgJ9SNgSi47uhjCfT9LyGjATVUh4qE7ebSSDvjEs5LBQTDmf/h3m0Gsc
n8AVRtqshoppramwV1H9n2djVJeoRw/XvB5cCPygUtS/i4ix2lMdi0hpZd7BDOidrKoi1JsYjECw
cYL9dUZPiandpLAUduVXf1ak16G65yeptfKirse3EmZhOIhe9vlUa3CN9FJIBa20uTAJKjzojykp
raoq8p+bcW5RYFZbvl8peIBCpdQiunWelGEIu4h765urq4IlfS1m1akT8ROYZzYEbvHUFG+paj2J
WMMOe/X/45uetEeaOE+rHALv5T4LQnmZqe2JOp8iOymQwpav4JgEyGQF3OyrUiQfXtSBqre4RUT4
Q5sV7Njr4J9jOgVFJFDIRExzjT+aJbl+GzyFpwSjLudO9CEjJQcpjYnYz5i1lqbDdrXMi4He5izW
NIUJxmK+zsYi++4ZqqeK3M3MMDu9Hq8qvTEIIP6qyJwuWzTIdmHrTHRFo3t85ttp2TTjNrDPsx49
2O7x21E7pPGkWRk9rDSucVAJmvqn3epG1R/oOjRrowcVWi9BvV8MS0XWG8vkrPOYat/ic748yJMk
x3YvNUlJn4WwQnpsSkbQzLmT0n+pQ/7seL9wYuCkEhBXlUToBLhTOoiC8d46qfAfEB4h4Fo34qIR
aNjHkOIJPzfVFAzt5YHm0BMqlw9QTSEhFNIfpfod+2lZdLnWnk3OgN9YLpa6q/cqHgWqVrILCM0D
FTiEnvPP6rnmMMSwrukYqVjDpjg8WDaJreEF6NC4+1abEZLaKARkW1SWtyD7eR/7IVUtfiJf4M29
EJyhZLXQ+dvhbhvKGk8Q50Z0+mcG+iakrVctAwy5jB6Er92Z1By3PUvHgGp9bXlnSWEvgfnXypx3
ZqjnotgW79wqvp4pvo+lwui9M63cTHCuqVECXKxuUkXcPgpa0HlYDDNPOzSnXy0I5OUaE6GNvu4i
vg6LNKr0DRszSyj25My8iYdrs5xawxJZyyLRHUDxGNxmZ4+Lqs6Brgj+kArLOJ6sVDgba1mOXnu2
Ub3kb1qjdePcu/mt6CFfFgkkKS6es5tRdWYp5/pGqDTPvnLjw4Hxx5S+glPS7kuMS7uU31uWUCf9
HbEWOSdBYmMS4fOvi07odFUV74fmB587Q7sULBa5YSwUV/UHLTZCsLJW37Qi/xxO1FXs2rUxdppa
/Ll4YMq7bzrOktyhZEvv8/rvA76wc2Y3Ti4pG24wBHTpvEDR8hUK53jPqDUpSiIzTqud4+W2Sn58
ShJM/sQMOuRxjRGmhl/ICpcOGpmGivXmb8O3U2oT+ezHps4KQ5xws6JrZZEV6FRdqaCr/cMss1b9
/7WnylO2dPy2Oer4EIgRSyVwuaffXagCHBohOnd3Yi+7hfPEigS4NLQ1o7zimHyyIWOI1cm53Ca6
zpYfYNlGFIQD6MuRSizSU4Dl10yBCSjYvto9iuU1+zAERgMnEsfQVc6g55HWQCCUP4v5IvagaKM0
Rmqk6xWA1Fd8VaJP4W5VBxkjv+QPmn7tPCRP//r3vDcVsRyGVksvkdBsI8uN70Xi3faE/SMC6ujc
q3JbB91iUk2QdRI1VfZbUZ6Bn4Mf8AwRpF3nO//ZiowTMdggOb1KboYryc+mhs4SCR2qB7KA0j34
G/bW2sOMwwYTr8t412pD4qbSl/fLnfbQ7sUl6IiIcFEfDC53xoTfYIhsp8H7rLs2FleN95mv9COU
5jodb+2HPGlHMzGG2dHIWmxZpvOh/stMnSjLtuz+reStl3csLUWyXDtLryN7BoK21hNnp9nZ4eUU
MWNmU4mcnsPGs0jYh6rLh0qq7w4DdO4llmRX+M3hSy4ojeW/9iHpoyYrPxuyKCU/4Mui1nmQ9GN0
WYoEfDZKRAoVYrkIpwrcDH+Qn5Ev+nRRQnAOggR2tf1K2g1Hcw4J/CMzq45P4bMX2Q4eOcB4Ftt+
MlEzo6i85aOnLMSGw1kdO/QkOsivrLTcR7So/+Lb3vxJ9X5BPfW1s0DSJtnCaYuAn4enCgEw2XX8
+Dn59nB7tCZtTvAPuPksEHCi3UBHT0mGmjF4H77CQg59Zkwa3GJZ6cmMO+f+kFXs/q5rm1M+NWKQ
OfmehmEuumcMj3kH4SUkrRJYOoJITkj8RKzvJ30AUEdYT8X+73XR0TsIThEpM+4OMHVG4cUh1ObY
K0qgOC5NXLaFWgAcgeSu3epI4efKytJ3sv/Ly6ay1b4w7SgksP3D3F4j0yZmj5O7DV0SpuD8vWcT
DqbkOH7gI21IH+wLqX/3/Ps+DksNhfncot506ruPGLD1EuIrmuyDVpwpbbKtmiM40a+v/l9ifeYM
kJMk1xf1W0QcAh3G7ZqQg+zt+qvai8Wx+Q2DMbtG7UAfzrRaqI7v4uIw8KWn0lzvAIvi3RhZ65Jb
i2MbnVCEJRZzxBaKVbUJ69lIC941ohxOLN/BhmHX+4sKCf2pYk09XEYJ6xO1XoZKVkRPJMNmwu6M
uLUXA3QQbIJ09410wZD1LI+akOYBUUd7PWEtdT8x3NrbxcCpWOqMJsEafrdWrUw8K2n0ZCgxHMAQ
2OQmlNaLXLcYZcpBgP602fjbg95QQy6jt9cLpmGmUKDccGhUSV0eYJusVTzvQNwzscO5t9L+2MZj
wJG4XgPG9RK/a3FObqo2Datne0xG2m8RVPVpS8hBYPHScfRrz0URUY9ovZDgca8P66v6Lu9YuxJv
Gtr0oxeHAj+525C4mW+03eG9uJZZEgemGdRBXHLxQWwumYFwWubDQVvg2ax3GeBKtJ3tjBGtPNZM
Dm7eVAJ65nUSIKL5iiv9JknOIWeRTl+uHkNvX/cic3ExPfjuC8awPsWtbg+K9T2ettHhSavk/CX7
a/mOHgWpsk5ojsGPkUBYrBGqlJaV91piOIPoduvMu9jiZ/2O1O2LXPrnHCnVoECpld/SHyOmMZCJ
UeQD72TUcxaTVL1+irFMax7M63Z3Vtd2gUoyzj7fLJbDX16dB1m7XQFfw4dCu1GtYOg2CGWwfSw3
S9I9XWIsVGmXzq8Qo0rBiF2N7CF1qGzQTZW6sbUsx4zdGZGmuDy5dU6kQDTqDXVin9T3HCkgevs9
m1Lma0AAqyTQNvc+sxYU5sk+8gv01CRjcU9RkZGezFEUO4sEBe5aP3my2c9U96uxRKHdkuNZCYv8
OZWX4pAL12MppEe1HgUlHcA4f+OfxP04Mo8H+4fOxb6DQ6SRlS1YZTIsH8BwOPNBxx5BSROajC26
7nZdQOAO6OhHm5+H2k78zLSb88vyqU9oNMCetdaJbpWgqiOtSP1F3CvMkEygUuUkM0uz/VEt5/Ro
vpobPk+tNFwtxvdTbudfqhbBcw5oBoj7EgMS1glwnRowRfOeIBuCrZwtdomnsI3liJdAoUZEcde6
ok/i/JZRjeWi+6lkBuwVpFXWZvOcHRrW/DsggQTKDnzZtBTViGwpIY2397GH2bGx+raORO59woDo
nhSihshGugQfBzXOGQe2geVVX6YyhgGP8ARqNCq0XAw3fOvyE7K/y2kQ45eA8N3/tLdDGBqRHztq
LyZapz1NXnpfiHvfzmCtd4awqL+42qlUIUgM/QywzXTHUe48+L9NE8ZQxXP8RZkO70rHv4I9EbvQ
2iACqclxNwNlUoBV3ULL7pZwFLCOkWBaAJDlQHNSk+pCKpR5SaMKH9lJtYWtNj2tlPKDOVrPb+5F
5L0wLSfx3LR0lMxB1qgwTlzhG3O8P++Tq/3FoMEEdwO+3Gae1v+CsZkAhPdjGQxvRqG6KdOHM+zk
FusOFjzA1mnnH7pzKrkLHvq4I5fNziMbzXENKj8KnPX57m0vIMRj2DOmjYqFxMchVlO1Z6VyJhzl
mEWN82M2GXk9e183upFQ388cFbjbyI1nReyQX264OoueLUgINE0DX4g/inbenMMvUewrIr1hhO29
oFSd9CWVbZHIbhWE7HHBNxWWc20VFcJSusfdH5gJFjaG4xnsrqGictxgfQnQEOm1Y96iKo3o3l6L
bRDZsqU3od+mOdo9yiviUODaVE28ujcX7coaN/IkXj9FunJz9M2HCbk0UZpidLtz3GZDew+6Beg0
LXwbJ+fu5D1QRfvf4r9FoCTphPFx0i5WZqXwjB3IJnsNktrJbauPQX3T9NLUtrlSqZmPoPdZL+Ol
Q+E+T7tenhKIBi3qlGAhXU8LgXoDTHKwF9+c0BMgU9tM7co3vRFj9Yc71/epJQ2ppbsQiAvBNjeh
mzdWQizyrGgOo7uSAqwVMw3bOA1hBWBdq/uUejKzOKGIyNeMsGTr5twhTdXFhRHezNs1g3MXum4C
6haWyCgbAdssadmaoBHUFdnMerjuHp30GER/0ovE06eht+hygRIhRfefn/0RkY2XJ/nPfwu7Dw7v
CzOYjFyaD1FNzifemhwedljlyzCmdCP4/QXm99J6Wu0YsE1uUM+Dil1ZBzYYDUrwxi/Kq0Pspfnk
6ECV/9Z8ZTrY5VeTupemE5eMqRvk+xaNb3HJhe5g3Zh/sIyhguOZXMCYmooVdk5nIBQobJQZTMdX
SsNP8HE8oYwPh2B2wSUdjoW34NvarG1SlNVgvBQfRGSjmGKpVkqDmQsJSP6wnli750QPtyoKexKd
CQmdVZ8aqwhhsuvugJM5UYlfOWf6NDidmiDLh/blBkwvjSFcGLQLeMEUs8enwt8Y3qdTZgaqLXoX
KwN9zKaFlzvI5uXSAI7U3M24h96ilOHNqS1mRwKE/mnEmwgCWjSTXoKHjkT6JrTkl6NKaY1UWhvG
kGAznYoILbBYOWN5UMCipuK9J4Zeo/MEUWQ/RD/Uh7D6sBN4oD/62yER8q4jNSrYORAmwroJWzbT
cxkpZ4pxl3QVDB29NMCjpLpoQsLd2Ax4Tv30YKXPpLxCLOwVeE2FQP+FqOcR4sW4J2Q75kQu/e5W
rTzj+WYexPO1H/qAgUvXN+dnvPezBvQOM7P6A8l6vneUgpu+w6xtt1Gnm/jQfYQRU7qTcpDqfrpy
eVkOffcQDAAq+iFCussV9EHJcDpDhetnfPUMSaQPExLvruPwo5HIAneKtINvmC9LDtJFqNTJDod+
ZkrCRwOmxkVnw8f5uQPCsiZSaX1KjjpXEYO1+8lm6YKUSgoIPBH7Bw1eJnPYrN3wmOgKTptp1QH6
xpPS0yF/F14KnJWRtgkHYQsM0M/Ea5zyEV5JGzk4DLeqKpVfxCeZrpfVIOEw4zHgFEScYQqLqPeF
ZfgPo19qtnx42xqoXM9JgOzcf0LY11LcVfecyJMFHc+As8G8YW3RGpbfGUW0RU0t7Hjl8+ygMG6K
8axkiuqNYv3LZgq7vr6oPtpKfTp4vAABjxNlkLB6rlCfh+ntJVZR2tNaZ4yTkV+A+cRbSRv2Hfmw
kIzrTn4bhjO4siwR9T1bebp5Szpg3EyTCgGqfBYThaApNCpFHumL4wlwsKTzdXILz+TUB8IZT3pU
crC2gxBnQX9ky/MP4r69SmIPBXw6ZN8fzp/bRXV+smPzL/L97xYaeZQ4RikZx+Q+Po/lWQik72DY
Q2vuZ8d0VDdbORorPYtpzxp6rMEzu1cMX8GfQIxYs0TcYJ87ZPLd2vh/LD2OzGXiTPOuKMBJU1f6
ZC2pPfY61EfTR+hrrknhMCvILAyPFkTemqUoN9oPOF6bVKwo3NntaDLH+MioC9W0QVZ3c0nswCRk
aPi0d/OUnRMy4GGvjj9mWlhzgpwXuqiK7/bX35ZKZZCFAmyX5uelLipNwEPQhex/n1Fdjb4EyH1F
+RXf1kMhKR8iP+dmnJR9Nm/9U1pvm5SwjaqFgIlGqHb/JNFg1C69wg5/aJhZKO/nn1ymzbd9NSTs
LxSRKWcymSOwsc29b24EDL3idXKnDxAs4B07aRplVZZBy7vHv3ZTnDQ0T/1Q7ko/h1hdqYUUke9g
GEtJgcJ9LIi1RDOi/m9po70PGHkV0rvIIwwG+sVABLunpch+/Kjc1Q0bAPh1JwYj1Y4UT8rh3SSw
LfFID+ON4901FQeygxMBH71DjYGnRchRAlTqYLhcwka9HHzNQalh/QOFeO/S8Nw814nORASdhCwB
FYDn5y0GjcaG2+Y7KZ0Al65QF+TiCyz1/CHXLs/nYLSIXQ5AYqCOGa/wi0WF125HXTEbL5xA9W0g
V6yu6vNV83MVw5VeW19d9DVPVP4G1S3nMuJdjG/tWc6Rjv3S3p0i7JPdyAxYe8aLLkjCLIBUjGLq
E+9XqiZ4H0V7Zm8TdvYjSsU9DAYmhMdyl09bBDd1oAm+vww5QreGTX59ugbLCWKVz+3pRv75cKcJ
3wCsLTMjOkK9lqOZWCr/Mn199e60kb1a/1bWquYmmKlEKBV7IycSgJdoMZNWykQtfv6bCqSCDUqH
QAqQCXJ94EtHcsI874Zwo789Yn7tpcmEyTCsrc/Vz/AqY5EmC/ZmDH+da6Ii8ftkliIZcv+A11sk
NJTaGX6qoaUe0CLzYfGSQ1IFlQh3HZQpT1CphJDl3y+OKoG2dAqfN92bamS+IfQ9qu5ZSn4KXs31
1OhvMxnl7Fn9Dmdq5sIS9omcn+UNus3N4FI/m0l1qsrh1hto18vUAYfXOQTt63SCrdgB24wz6ZRi
ot9h23IOVOLdsvCJniBJN/uJEb5hpImcy/HEA6SDs83sQAtWpCdJB2Y7bzscIayXg6MnY+M3J3kf
5godqebmh+xWe0Vegs155zh4F1pD0uOnEAsX9a2uS4KdPORaKRDUfgyH8swaeHFdV9daxA0621QU
73Rw74WCpcbEZA+3frIYUoP9qa36QIawKRgdAoN9yYlWlYJz+AhyeQuR0gXG/k2NUTCLkNjhV5mi
Vya4Q1Vo2HKKBz04s6jWq5Wo2iZvzsfPiV3fcrJ/T/S+mEyFnW1lGDDE5oRqGBa0YSY619TWvvGh
APvJIfja4WJdfUn5rPcGl+NBmfW5k9ox+ldQVPxyYKjKxvxuLBFNuI9rHmUdjJcKnmxRBK7PHO51
7qQH0AayCmuZnavqkUT/8LMH3UokVkjD0hQes30KMjvfXsMbatq+WwAkhqCv/YMfyJ6wj0hrPDiv
LWUBGrX3i4HnsiUAprf6Ylu3wOvs5DHDUqT5mOdA4LhpSrAeAW+/enTOwoNtEH7S736ePv/ScEEr
7/QzunC3W790W8PhY0SRMbNTn/fsrlH4mqw8nqoAUBoVVPY/ni8gqpSoWVefm4zPjfEEuz2IREuV
jhAr+UMOCvIBOEG5ZjFLNSLyGGveMGVcyhtj/FeNBFTXyrdDHWAqrEh8IN/arFiOyi5Ek40AkJ5v
Qwq3L/tXmbf8kh5ah1+ZHPvsAcb+n3nstH8GGymm72arkoOKMh43uaHNymTHcKYHMVW+PoVrr+c2
0ogU6P/DK+NJm30lS9JRyDQWYqhN2iV7iyNCcjAMzLj3VYNy4gtQ5ZmFYrxNauGaIzCCDO9gyYbs
0kkNLOX0diLRJBoXjv/cQGLIogtZbFHQ9M0zsmE45QSK8wtheMH7TLr7HRRACHR68L8Ecg/hP8xy
biRAK9LAoq22jx6iiykaNF1IcLKUf0rjlxLUCcx49U/pyfAyFTpwqGnahCyDON0hIu2zxxH06wA6
v43I8B8xpOBAeikNySfwf00cTI0ajg/XX9+oCVw6k5nueStfFoLfq2miMr/tXxUmQzor8rfSEuDr
Ux1Ba9SFIC8g943y3NpMl2aKehMSuKRDgaXwz7Vn/RZRkXq5VzgvpAKUwYCxhmitA1u0M+nhLkmH
nM4v2NnQ29i8fKsiToDOo1cY2BzAPXtgwBQuTjIsUTyLrzVemcZjFbawuLVkeUkuiggEmwY6mo99
WgAzd0a5j2XOUZSE3B9vnaqaDBu1DdMnh3KS56ip/cCguTwhP9IqJpnfVfMVJrn27SYHa0n6ZeLi
Zf4TaI3tOI1NWcFxbapRc7eqm9NfJI5ModIUyak9iXQss3+ASyP9eVBLJ+3Y+TfcIGq7eurT1eSt
MVY7fACB5aXm2CcaPTd0i30zi9Rx/+uC/RACsqfwpp4x3ZcBF9nEPshYlQF/2yR2BoAP53OTteJq
Y/cYJnBzRtHvZhOvx1n7R/Jv8wCacNNMnG2AZDkHaHwSOCLrxk4JMOHTS717dduusJGIFNVkavcj
S5m9GpWyAxON3NoJ+M98SzriBGTAVZrt8f5Y5Llzn9jceJ2vKVYbHxa1WUhx9NutGFSF4DCkOKcF
7178BbB20/jPuWSdOC7d2bmG2vzJVpDQaBMeDGsaPNXg6rb06w/RqIbvuW6UddWFf6SwtvSc4IrY
+pBT8/IWmCADS8l+xCeelPKyubkkk+vKcz3/dSpAMEzQ61/bHBzZ2B9VjXWkeQCI8F4D34MT4S09
tS4RzTkzPZCZalmNIrkHWUDAmApg9388WFr8dTOlHNNJzIJNxftIFBjmcuIyEBluN0VqZkWtL2uA
4fbe2BE2GGle2wmB6TMSfE6ZDS1NcBhpjZGbVDpKXI62fvabqjAbYDiIOlKzM2wJ81YaLhcmyLIr
JCz2Yre6SbYn6JVijf5Jrlr0qNwC/C7v9FaIHJQ+93sLzaAcAJiGvZi31V6LxZJq16771MV62Eca
6ymlhMUpDpYIBdTdH204W4rlARugJumTdEP08a4DFH3tbE/WMPrYKEGn2eKmeubnFLr1gTqD0/PB
RSq6eqOKU8OV/bTi+eu4geGhTJQVPzvUjbGLpmXTinpu42ARQ8MCP2kGHIGmxbC9cScpjPXWJzaM
xfUngn+wHthHZYob+24uEaXiiC9vxtPZIrBUY1UVwPKVUZFbpzLrsuLpwje2PIw2RsgeN8EqhGvB
97zKWnRZqA4ln6td3Kd6S22vY1eEhWc563iylKHtJN2v4CTCBkfHsn6JVosViuVUpTKz6NrDs9KQ
y75a9dpZN7lfhI7nuP7RTeDQDPVzNH9iVrn2cGWafW5k3TOz7NXCx3CIpeIP1J4rCd5NKxoC918t
L4qrz0UIJfRgK0WplB1Ez/BDqCyqFZCrsviQ3yKBxYRB0/quZGoGna9Ts6rz6oI7dpTgAwsd89Ob
yw18Ceg08FBP8KvWPfFv1LenUdq/aTWvhHk5B1qBLX9xuwZXbxFqq+Pg99RJpoSKv1x0/fjSykse
uFFt/1dNL+I+mmM6pFc6uniOgcPLcWdb16xWCUK5bnhftb/ynsSRDPzQkrapE6c3gqNIk6Qklh+c
BpaFBYtggMG01SbIR4wpU8Q33Cb5XY8Ert+KWn02VB5R5jYjB/jiJndsYBIFJTKhHbySXEjuZSGj
b2PZCNkhI5MdoD16lWxlw9XtcR7HCFUVhbpxNL02A68ah3lVFvOBwm5AFAh8x2ZbjyMJECU+JKId
ndroAccPYaCAQPldgRHF+tyCi/knECH0cR8Y/gvL3yMBNN5C2txuT9vArXU81m9lGYibY4C+QN03
To2li1U3NsEAnw/VMQ+9Mc379YgldM/CSSifEDKBqP1p4pPKK18hrtsNaso6vlVLXD7nQNqkksVk
AFBV856GZvK50MO+QyYdg7k0Z6Yac+FSWuCc3U+AeMhZLfXeKyijCyD8ArdDo9LrZ+TciW94Hzou
3qF/WsXGZ8WdPh2U1e2opzZR9MOmautfz8ZedxlvnFucStvnvQWNT2hvXjrrzNN8IdcO5GGGvzXG
oAEopQlBz4VLC1SPV2J9tMe2jvrudjIJF6CD/FXoqbjGQTyUlVKT3/7SthblC01Mq4RJQuGKqoXd
XaJoYrqB1QtaRuZWhwHYMq/G8jykkZFvE6VR5BLl0bOT7NKVxpOf2iDj1fVWdjyASVOoWN2Qyen6
qi+2gx3jSmDDQXDWI/NGBWA7YJ9jXHmt8mof5QJToJP+2djcJ17C0YiZQg98IE9vTdRq65sDWlr9
31R6l0a2OxwFmbRN+ZRSM1X3HeKoeFVHlEBUqAFWuNb2FIEwCBLWXeLN2hBI8LMUiJ11znwUEAPO
s2k9juNx3lsCWJ0mIsB1ThBv6bp0ceikst/lf/+/MmZak64MzBNvamjm7t+Zi3UiSAeXLnxpG8cd
9Vi3XOtKK0gsf1r91IKK6qmMOJPsUcNVdQiq+duuseKecBSyEfzpYerEWZtsjuStVArrVBvNxFJM
tnHNIeQ8mAMTbtKbUZknut337mc95ek3jldUBmjmMFHOCNCU+9r/v8B19W7Q4DTr0OAHvVDSsM+V
C4enmqFqzE37+YpMHbpzKJV1Qklewg0V3rgcUyRIownE+keTWBQCjtKbfkYhlyawKRrxI6SAkkeS
Q0wrCEIoumRr3j2dVxHNiO3jQZpOdPz9It1fgpC45V1QUqE5GAgFLHPLFykWN8urdP5nPc0ib0Dh
wdk+aqpMTQ7rbW2SWTvF1P8+gRfMArWNGrDFUVsSu7VTqyvEMsQVRrzJ0d8aOT4+a/aoy0DsDDqN
TBCJKjmIXrhrNSDNRius1yHx/PhwgsozwnarUj2/eKB7/IykrD3Ptfpab9SXxXuQmL9A6JL6bLez
/QhMQfAkNj5fJZWSOegaFeLvrZFKUPQ1C6kNuRvf5bla1fhD1i90FzlcZyqvlgZ9WCGEbPWIDE9g
7wczQy/AkeAUgVoaKIlBeO45BzQwrQnnfkVSt+zqHplxj4hhCjyVVLD93HYh1Gc//iQ4ejS9GonD
cJDgJnM9LKPTUl/S/N6HVKyjOKQUFHkhetwRxH3zV4t1lgzRkSTC6izf1LoJgiAE3KuKqVd3x9LY
nb98fcMxTWd9cKG0gait79RANQma4KPoM+yTYR6WmIqrxv6NwwRHmckcdj0+b14DJEHVrVJq9dnP
lWFtKiGIdAiq3VsBpPF12SMKFClS+u3YGEObnhuXsaBs/vigyiH1Q/+KMBBd5LA/613AdrRBI4S3
qeNc0YYSZx+wJFggnUgyRwGTiJ8MIg4/bbXOa1l6v3B5AlAN6HiMh42HG3Srn80eI57lfblhyCH2
JoIt7RrKJ7OkBgxJC8h+ZeRdNZbHUjhZDHdTDw1l9zkYi6guqRoXcFsuCsfIVf2PBrKc+Uz9nKAY
twti29uatUA+E+HC4YPo3CX7mD12tRxrT5hBSfk+uru8fBlHIADCORVGHTlRYt90dejvvzzzw9BL
rJvFlTckNu9WC50m1ZoYVaXg8ccW85rJsmvpGLIyBJ5kOf02CDZS4p/RdazJh9zPTL/zJn7JeZWE
uU+CxHIooxhelDZQ+iKD5hC1yc7vYGP0guwVLzZu2gIUUcGtSyh9ZDpxDowHsvwT4e2w3krD0d9u
v6C8Hjz5M7w7vAIsmwwDHOnQDSqT/6/QzSkJR08Ivw3pfW2HlUvCDMf6i8V37heSmU9CJ0SzmmY4
xf+5NjSvmwvNq0YBDnWzM3SwjvC1yw1aZKd9o56/EGCTP0l5dGX1e0GsNBVnywiAqR+kg443mFVr
Jx/CE+z29lf6OYBDrVqyCyodMhvHGYk++doL7RvxpPyGu7LxrxV9pFF6ICG5HkA0q/Dq12OoGb8c
8yVUgiCm2Tc5P7PKytzv4spd5fiDwLq5ghZOAxBG0yYHwn+mCfnS9FdQ4ilCJWGAImoK/OiNCS7O
iE6jERBJMsTARmZrNbSMlzFSQ17mVpuKlKgRLvCNcI6QQTwaOtzstwmWRK+SpBfRJTMzXAi3wfz3
eCs4WYKpVjqAf66aOFxPm+wZcbc2K12TBScZMzIAns/5iNfTDImBQuP62l02U2eYLKZjLFTwlV7K
v4nf1UKrassXfuJGNnKPcGcQwkPTziNNkc/584uW2qkxaOTSVNUfREeyvzB3QWaw2bS2DPk9XlKd
wXdkYwrjfoRRu2MENKKCZqDeSXrZb2HQhtsS8Xqmt0kwGhErK6skKpvkpHBxO7qSrFV9RudM3Glh
Ft/Ucz7DBe+NQ16bfwjDgZYF072i1oILctVcYeM4l/KKCBDtjm3MBlx/X1vokZ85r4fvxOvz6b2+
V30Dg6rZa5E5dZLWFsQ7yx0hgtn+co2DJcEbC22dDHJbdA2W02PZZB+jrOS0DJLffPXFuOGiWPTR
SpvktzziOD6RJjFehavmiRNVAxco3EOOVG81wLsQSFOIjIuBwgsCsICxMRhoxRMaZ6LsaTQUuYoy
b+NaKj80t3uVCp+gVPEfV7v3DyFIljWtBD2PhN/cUe3U8g5f8zA06UNc5uUalCIP/OvxC4HgRrpW
M+cDbvECDrf17DMDYbEah1/wMHNVb2IbhS8LFSuntvEOBCA/tH6kosIFPQYSXIQM6SUenemfo0+Z
LPor8NaqZnD6JzvZ48U61NAWdOCaebKJ4t0cDeSGGl9InRrkJW1N+YFarMIC/ZwMHmByPY8cOsu0
WcV4VLALhtBw1qwnd5EXxlbELo00caG//sw7CVTWBWPF/WxTX6OggKbBjzpacK4vPio458zhnApp
UzwuGY01dQodFGSzhyt46kjwgsmvhqHO8dKlReCuQWXzfQV1XsVc5jIWV1vV5Jgxa9GAcJaNE9YU
hYZfQ+o0tzjie5R2+SG0LgKLvzj3o2mGu4dPmLdE++10t62wZmsgz44b2w18pQyZXOhJEs+wp6kz
bHBgj/oixHZ1zBLOgUR9pf9AkHZJM99gAvKZG3y+uWkSdBxURuUywHzLvOz2C5L4ZQ10WLG4CN4W
LK0tO4kLatMPs0WuXyNIJIrujA2gtCOEpIjPUTqGmIp7mviuhJeAIyCWUPM7Dumk3NxH6Yr3kVT/
NXsOSDyiZ+Y2zUUZ3HL40T8CpaMnkDwcOHmi8qk9ajSNVAEOXRtI2/Ex3nJSFHAFeqCZibXqy+eX
ytoXEWTkcp5ax/jQYdbNdU7siQyMM5IsPBMF2mPFblX7l8kY/zCffHIrIMRtFVP5CFjXWHSlMqAY
OfVDrBvsssC5HzSCNFoAvOrXCsE3nvl/WEtRR+BVEFp2QsOYGUHQkeulEtqNM+bJJwd8Lqb1lnhN
exAS6K7YMQ0keAC3T+ccziEnArNRjZBzCtT3EuhWjlqLBuiQxJrFGsYI4lUjNaStkZhM6cP7BuRL
7XpTJ7bv+U7geeqmsGnEfgzzZ9MMq6x0IY0xny0cPFWPpdpPXwlHyV+zHndT6jEAr73T+ZLf6j5Q
6U9SMkheGa+zwZfEXjQDeUARJTVle7/bPJvMUkViZXENrYSETHhFG/Wl8fLakLO0C25Rvp8XziPX
gUsgqODMEd4QqKonG0Xw5QzlQ60f0xc0xk8VuMbuXG59iexvZvJjT8cFAjV//vx3+EHaPZnQxjUv
3ZaAXYm2rY5vutJGLQUO6j6zwh7+xUZy4j0hovbcxrO1vcCqZuX05eCKzcCa0gB54pTpASycABTn
nuyFE7bKiqY+GFqy7WZBKwe7zxk2jyQqYFA6/dop3Fzylx7jSBpP/SjC2FLcPI/MmN77tme1vwJF
u+W6oS55/Ve1bvuouCqV2BRZint5o5rhp3nIkEgHICrL+Zl+S7ADIqENT2msYkSCC3BTMxYgkrQy
psRum4h5WdKk4DEXxGhYYZwqP8N855N/FXp/bezLdldMOrO60NuI5M29NXJDxkMdTpydrBzFbjVW
yDncp1v/DkvGAblOxgBFrROLShf7LszXbTXLm84OvjAdKQh5ld0xwbCyuWMymBvVFI/jSIJNw5o0
67/Hh2cOzIppWw3n49STVVJXT8YxESrvLaBcqKEyfnHOP+x1WpRReMwaYsI/PS/3UMFbZIiPsUGC
7ExwgnRABAjMpIBAZACzQ52Vmo9rX8FC48dZ4Q+47wOFtHxQ1pUP79oYtG/lmrCNactM/bTC8FPQ
FDRuss22CyOqhc/dl/jYNGUVfw0AXT1Cj5Ix5izcsy/h66b33djwB2pHSRS3Bt/itQAAaX0haNhu
Ha2TxeCtBB4IgbR3vng5R4M2X801dPcZvMXTZ1uQPM2hHfr8EpyqBZubqMJdZt8/b16/AhjEZ7tF
7JMDciRlIErtbzPmtvnMeMeo2+spQwMwKgSCHB5OwI3Jwub/cjUoePyIa6xs7VhD2IDZzMDvSrv8
jgmGT47hwRF79nxged7x8ciTQ+qnXqdNJG0dvf85pHfRg/hgt7Fp/Yt5UKS6XxIV0XCH3a6kVt4Z
m6/VS0oE9A49NWBwqbN+uM33HaHbKb3nWu/3hz/ydlvfFpxjvByYZ5Y28KXNRN07BgWfzeU7lzoA
0PXvcEJET5AJJYXxRTLkoZeH1NpB1NVcQfuGEDvraveiUVWhjXE97SsQRI//pOWN0+ozmEYKvM9k
CB5EREh0I2gRiCTbbBWe8quSXD0W0pryyR/f2JuGjQ54NyKH+rW4LSWSfMXqYxGThghG3y8T6y+1
hNTbiPVbQ2mXKsTMqpPDL3g4+lGvfFRWCWjDbLxdKFltZWfDdntexfQyIJ6KNUwEibc9XI5ao6Te
GJmsFerBPF2Ro0n/Wv6mJ5Cbv+X7Egx5G6kyLv5Sv2b+IZMp4X4JTFY6RVYHkSJIi5GtkPUXWLAR
taaAg1sZaKb95Cr8jI0wyTJmpkJ0QMTYuvb6/8AX5am2yxYFY1PJG9gYd7e3AglHQe+uezFqLEnO
TUfgVRYwBfAhniIb86w5Zt1Pv4ab76uJvgwZIHyYRwsFLrOMIP9BeGrmxGIVdDKPQgsMftwBpeBG
cZiFldhgi1viIb8s1ZtzfK0+82EzQ9RVTejIwkzrRkP0owEsMfWoQgX6R8S94hylVIEzYraNqZz1
eCTRocPIpQPqXAG9wXS7ov9h8WI9M0OuPwxbp7ceMmVUj5TfCk9YtTtGsAy+1jFUw5wzhq3/XBfD
o46/A6nzCtzjfu/IxxmebUr3bz4DiMO4KH6zV32ZfzUAIGiOQKhwCovXrNQbPEbLyKljBkWdiOHw
hsPIYVV35NjP7mb1PiKjz6zlfavNje0exWvcdyTRPwv87ji2JxETzBymbqV0avB1p/m50p6LEPhu
mFMWo/ov0c7ufQTJMWfd/upp0BXS8TymtYIGtBoBCND7+hgldQCceux0qCT0+yW9ptRR18H4STHH
46Oax1iwZQn1PxsREdiFT5+N0X6gw8edaL3q78+vLUG07JwA2vxq8wV00pgWk2ECtZCkzesYkvSS
0U/aaiiIf22H1o3tdIFov572FZLbswhEg5y0KjIHO3x7xYX5EPs/MaXbBMT/9j3I21QUjR9KrJlU
1EqtB2/GHinpIXfLkWGW9T23kywGeUw0JWQSSl7FXBpPjM+gA8vTUt8GJ+73F7OWYV2kbrw56zZC
h+7aE+gPoLaHNYW2Fjxj3tkqWVxLvcQU8C/XhdP1SzF3paHvMqBKdDDuKzNIY0CI9HSSRMkqoheZ
bwZiB1RXE8b2fpQX0+BikFj4QKHipyzGExjpKiSBdbswgTrgTDd41D/QPOPYztLY48prm+CRz5Yz
UmUknFNJDA4Z/BfSslI2rO+rbq1FBI/TIrwFbYJbciwTrbY8owSs8mXcQWehVo5ZW5d/nkadYCDu
/rZYucLJVRhp8bKIlV1YVqUXmBz3HbLYKE89XX807uHORjkE2U4B09CtKk4LrvCDlfT2njfniEeN
axX+4VtZSjJ1poVWyyvAHTok2laaCkFRsd1R9DsvqMxDkSdY/dZBcL2uePiHS0FWbmud/xggy9ES
x2BgqP9FCxTFhLMtjCLj4DnTlxUPT7eKkFcJ2+XI+Fqnr5hs72DZNRy5dKQzby3Zw6kKktCQQY6C
QjVkYM1mLyUZocB49UXKlmAbUY00ipKluRWkot6NlbOeQvPc+r8Z/Gdq5YMq9E8mtsf5hpnygofx
T9T83aGJO07ULbJf6g3Gs7DTQelvH/I4FRXdg8m6a8tSHk0TYS6nz5+/i3ON+RcH6mHA7rnr7r/G
XVKyDMbEKIEAdissyafGZ35DoI+TdAXvzwi7a1Al0rjkwfHOhLgjsw2ccMqTQcZpwLRiVWsbsqHg
InxzlFq1bHIUVmi19tM71x1pHjJfUWrKAWdYMhHZO3wG5L1VmnTJBirxRPHWtZohwQgyc83QaP+E
bYSl9AkVR7+ybh1l9nDHjUWHf3rBX08m3VWLxMSTRbUrxfKZlaZ7Hatq2gz0imZpfh85rEKEBosf
i+J8QjdbDz2o9ViJ3614ZJ1moX+eDrkNTQmCUlayk3YXxzzpWUD9kF7XbS9JhYlZdV3hw02mbzhA
Txu/kHH+EUC6HJ3Q32uWfcOTvo195CAuOarHppolOghP5u8rCavGWuIAaUzMzDCWHf6/gifZAoNh
L5Q1HzFIrx81aUM4+pJUKc0L7ZR73wBJyT3BntMYt0VnXbH5q78RMycnnkYaJnZV2cD4rFmWGc1J
nb4hD85+ftQ3jjqnp0pmepgQUBqh9K//3xAYK7cfTX5AsHY/OM/1UVOS0davwkwX40GO1xwvv9GN
cmURjL69M3hMF4T1uDnQvdyN3C7wm3WVnly2fP4uMawPjxw2d2hp5ckkmZpUVF3mHUX8oL7hFgy2
d245B037zGJCJ63cchv8DvnrnB82DYW2Oj7BIq5rbY25UVqV9z8kafmeosjMBTVcyrC17a/hY+lc
LcOefg/ZTe5Pky7K687khKbfiRRvWORMLXZwNzjOYhto1WLj+jORa6YTU45i3CU9OKVZBnYQokxs
nRpg1aTFUo//6oFiqPQ1gtgs0OV5XDiR2Ip/IieFpsagoRwSf9ekE4VzZgecogAfSgDIf/0Ol+KI
XsBRYcfdyXUHt/0pu+Me5moNgsaap3bYdSvfLb+7yBJKEKbPdltUFD22I606YnxhV+etaRG28xWD
CxHX2bzd5Ud23IVCrFcOXW41SnVFn87xLoIqEamT8jd/zXRUPH/KT+sUT0ecrI1DRLHbivM8cttv
H8zRKoYvAf+BWTaoJZBkq/p0cmBlKuabeMjHMNELHaPs1KzWkhR0hfTfjoRWK5G++raJ/zJWUzuC
nNY73lnSPjzstB7nYK5WAHD1rH2++GE+U1HUgUwmqaiSn2tbPatgWGhx+r3D9Q8hMv8YC2TSpKTp
T8IeUreZtLGObeggFAEyr+bq/EAgcvHAetkd3s3XkyIOz0/lf7oJ1NfOkjioIg4jOrsPBbOuTYPa
xgCXyV6WRqwCF9YvRX/19ucIiigU84+BuiZlK31QGfQRKOXYoAJnXQyzXiWbLwn+SVhC/4cPuoTJ
vSACuI2SYU08pPsxefbi7LK9vcLE8k46SLVSv/aGOmBChWGz4pWHUCSYfkDN1RBOlsBGC1DCYQid
grLvnaVIfy0QFGLnbY2bBkZRZMl1zkPu4sWcuqaF3JgEjMKoesp7nN7rlvIovDOg/zjX4N6z4rK2
nlQCd6X8wWf5GOsML0RAs52GtrdbQyTVHewoxr5nhBNeRCEVucX/xblHX2aikH6o4CYNOX+nOHkx
/9JbFV+qaVSM0iVCtEOB0r90NR3H+POXUrb1biZXCELo1IIadq9EsgAeLddNNeiQxNNAdsxWChCp
9u4PtnK0Hxt2fY1WCHJ3n0SUk79V/Z4kDJu8vK3nBm2wCNdj30SfkPYkdC3e+I1iCA76favFjlan
PYLDdr4IYuMCXoUGhGtfTXtikmeT0Nu1Ioy4AyZKZdjwakBUEFle6OiCvpy8eq306BYvQAnR73yK
FzDGQz1UiOnKpqpyZEHCCYUuKfg6NlmWoIDFIfTzZHZl+oT0gl/XEUCM9VR0CgV9FCh6GPaInTWD
NfYNxvP4wbHvWK5XXwray86st6g8JZGHsBVGsngL04inNWu7/tkdn4eu4k4V8fCyQumIJr4qlvpQ
9+Semt8iQb+Akx8ziye2pDdf4HJ+r/jN/0KKBMN93JwPq4LMSAq2FquJ6WPH8aqX5h62fhsoDOhZ
WVwxM4gqC7SZ9dYhUXwLmh/yZ9xrqqMdbCaZqqgYxSnIA0E199uqt1xlrcWhmSWPe+ssFjBsbvfJ
rq3ni94V8UOnG/Q111Bq7KEs0350r9gzbvAXOAJrqLXagSNGqkdNKoZmgxhaWz1BKwFkn6l6t1rr
+CdyMtVW6PuKSF9OcxLBz1ajye/yYHeGM/r9skcI+AGxeQ91PFvxHzmywASi4RNtIFr+mg2MQIW1
0M38JS+0610nOAHhAypJM4EM/qLVP6dGxNHi2bUUqKryDIDOXhQ+grJZrSJNT5WcbgcQ7vEaTDrM
Ky5O4ruLUuBKHwlFs+1jDymLDFK3MbGNHtHIBlJ9VOYCgmrVd07Xz4aUhDEM/ejJe3ECclRKdCXo
7K6MyqB8b1AIA0msaQ22ZJLLWnBhi42PMXRVmx9cJgxslwwilDLuPX/qVXYmDvIhP0s8Uuq1M7Up
qlAZiYdHDclxjZbKZdr4pOjSzirSWWjhPeRly5z8UA7Z7aKKq16sxOS8KAdHHoSq/ibL+PX5IviI
LpbEW8pmplSgA+irGPwqBGJo+3CqU6gUwt7hNbNzOEQ6VE4Rmq2nqL1EzQszIJ//1tbguh1BJ5cM
XgZk0WLQbNwgA9hbnCYXBXxN5VjSBMu5BqUkiz6roFZ7e33RJs9wzYEwWS0FOHoaLn3Ku8T4Ai96
8elJ8vH+X9jcxx7foVC9U3G5LjSjiM3oQkD14K12FnZURd91ST6xKBZj7KiSrFoXK0gl5qyJ3dpw
5HjWtymZNl/nfDOaVBHY7Jn1li3dPqIkotrGbjQaKH7eor4bwF8YTNTh3y5mP6B84oP4FhwqFwRP
PCAmy6D4BvPIAaR6yIpe7QtF2PuuNTor/ZVhQbZoGFy8+RZGnlHpLDzP50accFBpRWA8kwKDMj4Y
OhhQZKmkmz8Mh5AP3yvs3VMxPV9j6gI8NW2wxohmjDyDHCRchnBITjjK1MwysQXo7rgk5b5j87gv
vHibHjq0HXPHyq/JmdsvRub/26pyyK8fcwFSfuYeG5Wp4uKbdxZjfsiGNlpI+Fri41smd6H+Wi+/
WXLv+4SE4peg97uaFm3Q4oZlhTHVsJItHK/ix3qN5RG5ehu1B1HRuTQUIu8s7+6v1qWXuGoU4eDH
JQ7qyX0o4YIjB5cwoJ+vJ7ZGNLS548qdyQI/zbggVWxO9dGdsc6bqElBNTw+cb6twlA25GCN2Qwl
/fr0fjzP1ZTW2/MZHG+MsicuJ+J4FsiCvtlzT4iAw5M+p5EnMObCHYghGFqZmsjKgMQULreH0IBN
WK+s9Ac4/XqsKI8b71osk+QOfPjUgyxNlGMTCi05pEJdsnJCfHQcV5dRS2R372jaK72SAcugrfs2
bJOoBFiC8fJZZVazztUDwbyBGeTy5BjTqDEmRjb6VYz1qYf/vhbRKRVZegBZ8lrmRG56CMWsz956
aXesUv7ab8Rgl9JLP99OaHf42wSkS1p9KeyNAdRhS0yAKEIs3bz9WL8ZIH/C1ir2nvRM3W+wWHni
1IwooHOB5llLwE5Qr5R1T7ypOq7oZnxdJhH11n96yx6ALDXx7Y/LdXgWvD8DuS88W+3rtpnFagPM
qSRmiE3SsZbsIqMLd/M9l/kLjbKMM8leRAuJM3qXVq4pCV2WNGkCUSm3+AQ/Lordm9uYNXHicGRh
LooPDBaX3IakuZRDubtlo8Oo//sUngs1QZ3/j/J7K+ZNYpyPgcVJZRxZ+GH0qBl0AfFKrVMVPK6k
1P29UJU0XnLZ4S17CI8zsO5D9VE/ZMB6OAGByxVG1nx8wc+D0zLVEid+yfxIgSQoffcjqaIZBKR8
Pgc/30rDIr+BdvTro3V7CWBIoasQjJuvk0FhuKtFJOgx0InbkMlyhvZLpYJ8AObabfXYJRFbAaUF
IurS7Qq6/DWq9kmS1tuK2IUY/1KPjVR9oZY3j7sTiT057SN68cF3lZUCld+ISn06X3EQRe69IiLk
9kQF2bKFY4VLbLLpnmS9f899NyEH7RzJnODD2M9I249Uuq1AE26e+AIlPfz6BLnYVim52f61u6qy
56OaSc0GexdtC6sWU8r7cOBZYKglbluubveD+YCrKI18UV4T1Uydjp/xGYJaJ76FNO7xa11utHQ7
DpMjC+KHKqYc/zOk9NxehbnAJ3T8V41ZEuihoOoBl2MJ4Fy5B7o5ZdTelP2DqFrTjad4NMyQYRNo
cCC4H+rkk75o+rNUa9YRz5qgz6Ws0G04HdlDjKfm4SxJYQ2k0SRkMLyFrlqUlh+U0RB/PLh6XtUJ
EaixVGOJL+OIriWpyxdpdmq1kPJ7DQFYWdxlrAAvEfE50LfnDquW+SR2MUN2fZ+FEqdYBMWNGz6g
RW9OLxNKFbQyt/mhBzEqBjvDavJXfKj3zGbQnBhI5ztn2RUzn4qOAaGyibRqgBxQxc3xza7UlMcd
M3zaikOldeLbVR6bVuaux2t7LqTr0Ak8MKCSyyEKXdUzqxJp4Dyhr9A+j5/jqJZmLdA5IhjNEwAG
T1PTtgKflsbVQB3/W9wHyxoDaBk4QaS9y4vVjulNPx46486q6LUOdoV4sXS6Kps9J4y2lxHkUoIT
q+NX+0AntBPAUH7ClIInfZQ9Srb612YaWL8q4GJXLxQuqrmJsC560I18K/2YHfNhE2q/09atKxjs
ylzvuVaRbvfx3622hujx1l2h8STYjxvxf3ztD0GDXRNPj7BcT0msGTitohDG72Is/A21s9ircCuu
WSKfCXY1wHu8X9qZOe1PZSNwEQfaURxhr92/g0cm6PuHyMJcAVUIFcy01MfGGs8GLQ8sB2VuzDhc
CVpJ8DjJrqCyLdsBEJBu8yV0hJHnNza1ZeosJD3/eaqXpsUDswh8VUjvyBPxwOmhdXkI55xSSQ7S
d/FIwd7fEPHoL7Mb4v1mCt675+OPYVojKL3jR9G9odLhYkCZbDD8X8gBUq+mxJgxn32SkrYhgYKK
ZsYUQO2VbVfSc/9N4j4gbvOfvP4D+w1JO9abyxsT77CpBQ6IGabNJiHJnD5FPRSTVgtnaPV1DFWc
KsbEIQO0qp8RlAUekPqBpAP3LHC70jaojin7L2DhKkU2M2biwq+bIl+ZGfMJIAS+XGBoclIF4zrP
SIfRc/IZUebR17UJgUVqjzg65tY54gN7gX6ne9zcex5RSbQkKw3mpwtdoIj44DPePxSj6XdxZEz3
PS7j0atiiv79IIFoZ4DjDSXPL23zG2IL9vnOb/prKJ/xzgS/G5Qk4qzaXD667TGkyfUBvdpu9yVr
V34VpdMtdv/B76xP7SW1nFX8A66CRV1DXVBXLbkt1TJ1FQAdd1MCkjGwv9zvzBzkTC/Lo4UD/JPa
ZSRiWShGOPDvcKnHxChj+HIOnyA3Dr3yW9/j33d+rMqjdxr5yjo5RdFBGrzrdInzw4Fu86+W12FW
IGf7j/Dk5XIuCnvagsxOf9au6MwNY4kuG9xU8DsGHb6eUi3eZ5ROTsSGqezoI+5MFmguYoLTtVxw
TtlhqORSqUbB6WdREBGJ+GBOYMfZiQa+9D/rU9nEdn+/3V1YhACVMn8VItcHHgCKTzHsuA66x6cG
CvV/iE3pP7UwMuXZFZVIh+/xh7S3BonEDrNNEv4yYPLXzkQS17eA9TG5X+gf4XNb7W0bZaS/Jbt+
y9WfH1EOTv+X3Q/q/qPAEfZvUxW8We5bFHQG2CZ81uVo6nKj0XWISIhn55WXNXHQc1e3leY5NSnR
x2YCHvOD4F4w5BXuLeyxviDQg+nAC/abETLQ7AjwVNVUlVXtFj5lCAdneLOIE7wnSz0iEcNRig9X
x3IAJ65JtrejKfgd2eUXhyTp+6Kf4iZwTRWjJRYUCT5Lqmn+ZWLV8VO5/XA9+koboIvLWwZ/FM5k
w2If0A3OZur/YEwPRL26hIO/4D4pY4ucJV3pOhPksS26Te8MDL4kAcXQQYlvsojRP8Pd5OZhv0ji
V5dupqUnsbJSP+ilRlcHHxeMPi4SAyT6C/oTWPZ5HmUDSB+G7wje4U/eeLjxHoM/m8Ka8GWhCjbe
4FPVpNY3EGO3H5Ct28JWHyahwGCBoRH+9NbqjG7Z+Upau6RMyy+47Yh4fXO8NxSSgHIdCo9Uy/Zr
1v/TMj5guuZPMRY6rN/Cy7gh+Bdg4Zbh2JtL5nfM4scwLqKYBXYxKU+BotwrFWRJc+sjRYXvExTe
/vOYRmLUE8heSZWtBUPxT6WY0lI57kcUSS3sIbV7VhXgOZ11GPzQ8IGCktZH21bi38N6sn6i7k3D
JFjy9329NNmqh4Q4ZNdMcyn5MqJf8LYzl58eKRUp1n1/zCvjnDFc5XlwodKzA9tPFvzUe1pmmukv
xm/OysVX7mTn2VIoAVOJszSwUK3wNRCpeXqhOQccQKacxshrFWpyW4hlRjbuFsAbwCDoqy4WfgIT
T82AjN8m2KTqF3YsNUByli7x4SwFki18FSEeGsiJ7PFPRm7mQR2TV2Rj/PwLm8y9uYeReyRIwza2
ubGhEglyfbhwIImOpMDpqUP8eINeHGgIqSzSC3ARajamPpHskDYZsjWSoqUFtj9F5UsidCpb7MBi
m7n2AfpPEIO+GRzIggtxNrjPlDak3eLiGAOxmg0bPJAzGZU2LQDzDlfVThfPBs98SEXAsblhHV5B
0JTt71lmyC9tJW/Le1N4FDZR62+pvDDG5NvdPzt89dSKbr6MEUQ7y+snFjqaalBKs0ZHshHUfwbi
CMrZMvCRXFD9EA6ptBMxoKUVeP33xZmZ8cYAYVMTbFBM6GT0bhPdbRYvwV8P5dcNg2JEi6AJrK4b
/6gGa09jnUl14B61TN9KuUWRKVcPsYc1X7Ncu6Ry5u/KqRueLABmDo025G1EnQsW2dVB3EcdukKO
RgYQRbBwYSYHfclTNX+pTBHt7AnCGnKx3cz47fFL/3cSDFDrgUmSpIceIdG7GoINk6D6NGCnkx63
aUlsU+eFkFv/URkS9qCerhtCQaWsKkgP2sJzLSWEgHnLNJDInKcTNZofkzgLpxYZNqzrW2kq4HIk
BvAhUKw0fa/o7v9qVqhvk3Y/0+mn0Ma4yA8qt5BjjcS5VAKz4/h305QRshoRfR107ZkbN9N+Q89g
2hPaLRRDo+4sQ07L7R5q/nbEEqQ8dwjjZoLCY0rKAWKoqSvuUm/DL/Isrvs37++fCRZllQkn5I7V
OhOiGSm3X4kCp6eSPN5z3kSTFkxzrpWsxdozXOnMmz6wqYVtpOc60JMpMOZxrtQ5kTIc+4LooHKK
YvYdwP9xlZpBSM/9AtBnEan/9W+CErINKHEe9iRn50f87M6y6Z/J+0QQge/kejpJjO1aUMCspWVI
Wl3hTfYSeIYBh6cxCadWkMcIEDFwpOpXGYK4SniMOV+shz7Y92S9C0q4jLeb8h346WgOPtgDWUl7
i/Em/ZOjGu6pX5fQCLeftZMqx45w0iUUDvuexTc34yoxpklzWEbDhecGK3HcLBu3YRPaVcE/rQgG
Pw8eRSl0FMRjNuNIJIxNxQ+dz8ozciGM47DS61ZEzBZ9JebwBGjD+QmEQalDootYzOuVzWsCFDYm
2JiB4uXhKzzkMZ1ELgpx8qUEXkiHw7Y39VnEXbMu2brD9lLNBIoAP0F/0ryIt37/RIuXFHNcgzzR
OacsZ4xJ4hL9/yGT01BLqO+7XQAJulqn+Ch8pkSpk+L7drP7fu5roD9JTea0WitKSoncUOZOHksA
kNd1AudPnM3c6W8V3ux9s6Z/GWYSH2HQbx0cgMECnj7Acip+2PkBc4Fii2fFFs4F3Bjjf3DqCR3U
TUZhpgJbhZs/IY70wxYq4+SUa21cKmNrFg9wQDAt0OghbUySPc09X5nxU9Qb6yhXdcCFrmy4Bh0V
nMio5EueBmK7iTLVlne/a3hgD5vWIP6ElYvQK519iUX7PAlJfPp8WtiRpJMBqihw+rV6pPzRvRRE
xk3lKhlQ7DOlrGHSJzjkcsoZm2uru8o+hgZ50lSvZZq46fIW3wdfORdnCJnkDVJz0qxaef3qBfCv
Gn9qTsFrgJ0vcx84QBys/DCUwPK1Y6LsvHZVr47IqE3enbRUhXzlwDdlBdppzENiHC7EshOhu5pI
Jz4h90EqK9zWyRegxdMSI+vOPbjlMhoO+UMXfDsqziSkPki7tmTKqsnToBgD3hRjoH0AshD1WVMN
Q0jBIoNU+imWy2xcjG8tpLGM9gCdiER/9ba8KAD/UyWm7ph/Rm7aHHWfVpp9z60JyuRQw0dXeDS/
QDr6Ghn+nmlBFasvXPRM7byH6qZ15yAHqOMcFfTo2EIcdDye92wUgxsLzcA99bYfZvtbrudNlgCI
X/g4+PBnWcxK5CVekGkvn94lGMkpQq6xPzjL0DOEUHZ3JxEI+w1+ueSuPdLPo/CZSgyilafjpMgG
XtZJSlfZLt3iWrshGgvy1/w5Oj0N//Dnnq8MLkDEOvBP3oM80gbqmz+4w0lgHxG5KOG/TKMrNIB4
Ig99ZAXZ3tabSUpWl4wF8eogRnnDaj+H9hridW/BmAXHSzjOYqRWgyu3lhKF//zbgptBzSDixPZH
IOd/r3BzBB4d5u+I41C5NU+02iOY8nmtmWeBTGvQWH3SES6hKYplN4SiEYNgkibo2BkaWihqNFYq
q9eY17G+4hQjzMTh0JGcWFuaZLyf2MhFV+mKZy0eoYeK2S6VYANY2wSCt43uC9x5TPEZp16Xp7D0
I5KFdWVVuzUl/9VN3Qvx/zkwoKpbtNCC5zC+Jy7XYSC2OIF20Fa9CrGmyTEX+NxluC4B/CaMwNWp
87SxThVA2WM8MLt7r5noN6Lo0S79+XBvCoCaJdF4PTWNyNsvsK5XClfyCHltSQ930jZ8LY+ll02T
bqUfJJYU7+65wP9lQVsI9LNzZ+GoeryXYPwAldFcZVQ8YeL+N0bGkqLAS1bFPv8FwRZY9/PTIQZS
gEfwZ5LQe17LcehKw0Tu/QTKbV+YUGyUk6a1lAfvOHKHVfrrtVRxEi0cYyqYVILRS7q/FM1TukJG
xAHknk6o35IKKsTOIjeiM0GLHkXIDol2MC35t0puKr+VNwXswF041FgjDVgnKYVxRLBozR/28Vwc
saoCFDTUuEhrWQ2t8jhIuCDMXbtGcTG4vBNzUAhgf68rjlhEhvyT8XKiFQFztlS0EdXUhKSRC4DW
3t4F+HUhNlhYk8SOYdt8F3SQQ+VbndYXUWoX0v5sIU42JyfL+yBdeTNAaI2hMWCMCJcarMiapsW8
BsPdKbGynqb3B/6ML+j5pao4gL+O2T6eneWNhBtDWdqKYLZIvXyRSEDAXWros4bBTTa024RsvltP
horW/DkFFAJerJW1r4QOwzyvLEQSRSvatvEYcNBxWnRGYSOgtOjiOrVQ6gcUjO69BHbTbQHPkPmz
2jLy5Fb3Q3KVqpE6KRTWpta4hdUozXQ4nWpyrShFJL33644aPi3DHERteRIAhUwNjXZwg9S346+j
llw/TGrec+zeGEDjcDTGClEDIkXKGfA8a1ZLRmuogTRWB77F6xFu6BKm8A/OUoDZDihLkyh1jpA4
SHSa5srWlQizCvdOFw4yc3SXq5yMeGzdTdCpnuE9emRpSxTQzGrbdBl8eXsDa5IOi9Nx+ydSjKLG
WFRqPg6CVdFiSc3IxApHCD0rqEhgV39ySzC6EmzyLts1EY5JwsWDc0gijCK3eS948AxxRJpNbhkw
NRRR1zejpDKnS0bviIrYNKCCIqtaCnyEjPfNdzq5cnxK9PaU5oHTSVy+I7kwgZxjzLx1LGT2kukn
AvVDueYNzRAqOx8r7vBrnnqG8RJ6x6e4pfb9/cWYRCVdAXz48Vf2s4TOfvSyZDUqlSc4uNmNufld
3ImWsa+9u80Cm/l7B4kJXa5JxVPOqPI/0hw/JQdKo59FSemmoB0jQqVWkfoPvi+WHXqLb2XCtQ6N
C4WYW64mEkDv9zh2IDILXBrQftvQKP2L5FkT5xTbyI/qADiKf64YQih8fE8gNW/IDMCKYg+UF0zZ
NYz0dBmcEme3C5hOrIIZ4LSEcCSdwY6oP7L4deHAVXs45qdBQZJqt01zdkX5w+6voyjC/fX3eSET
NEF7MdEAAUYDb9tVi1qAoa/1HfjnWKfHzJCvhT6dzXfAyRz/RQvnTwfaVUEN8lXzYURb1U2Wo+DQ
bQsTMs1Hflykse2j8i3LmRkT2ox1Ys81VqdhF0e9GCB2yIo9+2/VSrBlHDraJIyVNJd/r4UPDWx5
+xgxui4LnLg0QWXxDa3Kug46ErZQrComxYyNa9EGCkEWe2M/55iDN94u1QyTtoN/6WcFCHcnjyyZ
F8um5sR7oTmMqERJ2nTvYMaXRiZ88DB1RLKUgY154uiiiFA6C/fq52jRhw4qWsWNqBRHoxQ4ua5t
lRvMTPois2YXYyDoa3AHxiM7zYi9axSqCU/83DuW53B3Y2par+qbMZdw073naxa2SeW3xwYGq+HA
3OlAgT3dpNdghhnegqnbQlGXiC8ozxYa1B6ixrWRbbLExK+jSvhNSzRYxalD7m1z7v/D8QGLlSs0
usbTSNU5diLkY4mvGmhORhpli6aSV7sSdOYm4wm/akNJOKREqdlRH7FCt6SuID5JR4WwHephsWKb
oMY7MIcjpywecFrqHVRSzVl8Zp3+dzUCHI0WYt1paqjmkSuVeqe9s/jziL3kTwUVH5j5Mmu0MKFd
PuIF6rDgG/ij4kyO676nrn1RlykeZ+TyAydamjVXT1+Fv5iIYzEn6O6a6S7LUXyREpSHJIJrJD52
jgW1pS3wBq7YTsjUITbzFz/wPbzZDaZtefihsjEuG9sxGtt2PG/a5d0HB0wzZT9OrdIVDkOa3zrB
kuGM0E2zLKSTLQwZlGDIOGkZ/OKuFEYtcKFaz2J/lSIw6P7oZRxK8RW0Pz2vmiUBSM/YQJxw3Qy/
WBnZMY5KtaF5ZnIACn4f90guI3HoCJAF6Xh4ABNdeYhtqbhxqTkPNI90lmAv4ost7pgaVCykC3zb
7KSU4fCCxaPOeJsJs5oZ/9CDVG7TF8z2KUrfmZp8F0GN6XwfF72JwHN6c65kuoLB5Zglx56MG8Qb
1MnB8Kp9Eq4E4VnUdUEeUv4XLiTSEc8RehJiVi1yY1cKoXk3DAluoAA7jHQthbwfVpptQo+SoJPv
kXa/zxD6mJxMjMl49InnNIXcnSWNeaaxkmXpB25EWMb4v30EB3AI+YaO05J8pTwrKCElP25IvARm
ZVsk/NAqpWQSsDkgauSUZQpwhqZmNaa/fsaa4OqGoL/YTe56ezlhzvJg8ihTXG2n/jbPEjZABGP6
1DejjBehGCL+VAmvLkkmjUfkxJhcH+4fFEONh8g9CmYY4OXN+xvs1YPjMpjyo4THuxgI4ttvCSLq
JH/3x4vesthiAToQ6JO9BnGPdQ8OIvTs8mXZj29FuimhuM9Fxofm7wLImPF9k8vEy9qENxWx+29n
pqNoWPhJsfg34GXr+L8HEKjwSDjbxfq5GTiFBpaCy/ewdC8r+jDKvoCdAgiTOSnjQxYpXzigIO2i
N2/pdSHsmsitRMTsgK/sJAyDIf7hjMm0R5O6xRWaxBDLQ+rVGAizuCynI0BGx3CGZyAb1HojmJg7
wVSqFyC4YtIiYdUsfuuiKFqTF4aC8iMnVqsfxJUFxceHreWx25F9q3qWx4uq5xO+vk5+R+6034By
ua1IVC5Ezit/JpuAB3t9wOEMSBbu+LiG9koyptbrKm5FbpIcGKtFozShCdH/cqDK4D2QItbGJCob
luA1xy4G3R8xe6XXikHab2Ns3pKT81ujze1TJBZo3S1khASSMshUaKroHtiEr9NZ1XyOODjiFriW
zrqYQ3Qs/iDNOr6onFUwzyMFUt4dgFv9pTNDD4VKnNUOMVfDIzO8i8PROEGVMqPcDRjmK0PAWMky
WsojLt1Mgrj1+PgWFdqVtN5tQ11uJ2OA3PR/uiITP7W0ccNzrdBWiH5CeFXSFhHCj5oskUu+epWO
gy7Po2DeD3mJ9xX4x9y4kehDdplV8bDBImPrvqmCx82eNDQ0AGqnAv0ZuqHPuTo80Xdk0+SNmOwN
K60qjU4i1wPJsT3Nky1p4NEvtTLy1JDqCiWiR7RMKR+zvNSxSBeUDAWe0patOu0VC8VcbtCzRXCi
Hj5bTTdJLIJ/+Gk+KgI+J3of+lAuStU4gb21XjUgAb6fELy8fu5fYH6+rFvCXPj1XL8ghwRFszE8
yPgq5xWuv+Aq31s+Gp/Zv6Z4gz7NHmUYnM8GBYaxYL/7tlfBpgM/JhxtxmAndR1FuslLVPCCKnqU
sSuRBVEff/p8t4SqZp7VS56/xPDlWhTrIGG5Grf3o3RXZoeMfTewB2DTo2pgnynlCD3jKQTJj9W4
qEhKKP4JZBH9FPh1mFB5frsLa4XuDu7t1/ENVnZRRYel7WvCZIbnWaAfhO2O/S7ICmaoePbDVwWK
6EqG2zGrdEKmwVq12+uNlT7X+GF/W6vx+ESnXrUzREGjGLtIUxya7giwXlR9F5ZVxlowUdof48hx
TpCujWffAFvgEpNCJWimO/eGZb6YtyxivWSgps91wUW+pRnr6W/cC0N2gmn2luJ9Pf+AZVzKBBtI
bmRrOswVMBILevEhDqnBfEfFvTtvTOqxnzWxxgKpcUeHom8HEYsvgj2DBNhGHnLzlL6kp9pZj1xQ
5TYDBCgUzfg5mCTZMQyToSJiQzL1TxIr8/T2wDWOPlneUuFeV11olgavb3IMJaBGCDfI4sEIEYBl
2yS3t5sT+5e2pw4oG1oGAowzO5fvHoZTb4qknkRzNleAT2oZr0yMXZGdm3JizqD5R1Nt4qu412yI
ttNeFRQlm1PCcGnZcDEo1EcBPdpdHt2egBa92RxVd3zzpejj/4YKiJbpcYpOgYd/D7KhnfFGezdw
Q+BjXlnCwSfvOOWQUUWCTF5coWlkE3zYItVRdSoJhjc6O9DRSpl3dHfWJzZwYohPs8Y6OkKhNxgw
P8L2qsyzIu0Us9+uLijvX/LgB4e2U4+7evubL8og28gBB/djZOn6D2smU3kl5hBfpVAihZ5BntbH
SclgaTp4BH3pHC3bO5QrFHly1pd4kwq6gc8syK/6k72H6xlY/1xbyvdVG0dKKZCGCo8T9CB7nVSE
QnyjFKhBH95r64GZbC3JbHf35lypCgP4/OZUPryOuZ5qATwaqhs8oRbJ127SfzHEHHsnRBHkZj9O
8V5J2/L/axeSQQ/JASsYBOzkQSvxm5TDRHzHZvMN0TvngENP9YNJTb9aKWx/QDZeUqQgrme8oSq6
cv/CTlYAmWVU+TGKLBiSECFtMkNa3BukIh2qajdHy/Zr3Uke5QDrUWMlr16J+3OX1kUxJe791Q5R
56ZcK+iYF0+OcmrEHdv/5XlPAAKIafF9Bm6FQ+Z20m6ycWUpgFbdGni/ez7HsCeebCeTd+Aav5B/
tXP6cT4fF81EzelzVIHfUbFvrr8sbQWP4Sj+GM3o4o/P+ypDoc5N+v0d4p02RSSyefrySnXvN+EW
Xy5/QfORqBsAGifM1nelLzgA8DcVpUxoUotoUsF/EB0jrQTiBlwDtTXlDVv+K/NZrZK/h442z9vh
d+xb2PgMTWIVfTomMb32kXSYIMLN38yWC4sE9V4S85wyKiW5+kC7zWdetTDP/tKYfZW415tAI1SV
V7pGNyFOHjCHHKoKM5P33YpH6WR/O+uOOw3FmfHWwn3Yo8Uh7TLUBCE2xiB8YL9skSJpNXnv62eB
4pPZw8qCop6gTDpIFpdtcquAONkAS7sCptgx20MQYGkwV3/Ia2SDbQ3qZ/hop184T0nJyI9hS06Z
yMcrtHqvQ60XKtS+Zu90+Ec7RLY359oH6fthYYuHwwiDHLxujhW3lx2qLOaNuD9cvvqdI9Pt/BZ7
5C/DLYknvRYkqzvnEdnfsJbfZRLMI9t9lMGWTUCWJAeNoxh6ndpZU/vBCPeAfYiCazKE2Wet5ekm
ojpgwhDbQu9p+k7BfclShS297ur+9cdFx/L1aK0xHeKFXv1SaadoqcBopya0ArFGoMhVeLcfbvqn
8Y7p2+JdnVrcnkO8+4Lv1IyiiLvUh9xur2VSUrwxD1EbA2ENbmGfrF2fXWRd+RCbwyMqwW0pze41
MMVzdgST8/IFz868uIoqcwapExv2YyiokcplvbwetkHqIHFSwKvp0jlJt9A+TeN4ZOB72UeL988V
ifeOIHWkuiXJm1G3Nv5fgmN7zIsWLIr7J1KyOYrQGjFT2fA/DqLC81xqzuvkAvytucg0YVuGl/OI
5gL22XuB5rl0uI2aqoiW/fRLsIQ2sKoCwBB/rOXYnZUCRXaOsQ0JgLzOiF7BOaQfctfwAk65ltV9
vRzuhg8JGQ1ebbh7O+HDfUzUT4KS+oxc077gWui4bThl9mRBf51FJt8bB9Oo3Ukiq8YK5OHlv909
eRQl72oOt5RwOhH9w9BmdiEJ/S2nZOoULV802YwsBmTMV42rY6B6zodGPoX8u4Vtzu+cowDq2J20
vp5qcp13427YSuYkX2IAhLp3ZRaRQig7Y5rv2vRepuh0TsmTk3rnbkR6kuJHjY7cBXdSj5CoN+ms
qpDtxDGTrG2RMdAZiguN7a2Ox/fsT5ooxTA605LHxKaK6I6JqekWRpTaapoJn6O3YWi5hIQ8twJR
kd71+C6iDbMOsQxxeqWx8BAH3r50DX6rEJVQuQnjBs3aCUXLau1WcFrc+WiPaK3JYN7kcUEns58u
caMdWiSe8xfXk11FSqHSoDPZhTvdUWa88DykQfPwwsXYJ/t3gPW4zIVe6xL4/n73PjpE0Wikuy+d
4udN8ln+r0P7iYSkRgGYIlrXDdzhLdn5pJfwQYrDfe5wrmbAzkla9XLeY7XfNSzA9l0bFDB/FliM
HsYy1CyWSp9M3M9vJHOxvfg4RDJSW9miaxqBsdfJUePjFBuYJVSHh3+o6XdXnZQZvdlQ2wiolMxg
Lj2evWf133HxPjpYO9/DGie8lyzZd5rCQQiJ7NCLMfiDHg18SuHeom2O24Af2bRG0U5GIGzjNzM5
hSBH4zqkzBZxSgLT+TbLVkXFp6xF6kENVjprxBywwaLih/gl5rsgZ2Gc5XYEG+tUzA8diG5IKeOH
vWTfABC4r1FS633vOq8EDZRlcwMk1m5AunPSK7zz0i009x0vbG8vNbi4xsC+yfOf0dd5UZxv/Cqg
rxPrpt9LamS58fWsit4yFhtlpPeH68BZZ/cuplp5DKFFFh+s2r3qtxv2rcJ1Q7H/ea3TNsXqSkVi
jNmktMem3Euipu8xyh9BOlqDUsBX2fEKsovYL9PQ4iYXP2PJOE9j0l0C+SCEpjRf6dstbmQHElUj
pzkwkuIuHE6GLwUkXLbmbxGlNzmEmcR72dTOe2gVHZHmfwpBt6MF8KipozrEVMqziwdB7l5WcbXk
7k3uHxdGOtjmOkSkQBDNds+5ZH2wwS1Y+GJL0zYvWfJxyjMtrX+0ymvk9+GLXtxDqytc0Ym5EYaL
90B2MJosqvLbDqg69gBZs6MGLkZvbLFD+xHq8FOWt6zLBCZBEhpsNlivldKW/+DUp5AlbY3AJvir
hfF2EvwF7QaVA2VcE/FmKtxHJ7JjjJMslQQeblIbfToD2nnyWwr/ZSIPRgF8Je4PLOmmA7W4kw+u
9YTZuSVmzoI/fck/l2WJetoTm9XCQUH0xFuV4P2sxnL5UPR9glQsbdXubbLC0nkBDH2jW5b4zPKK
//CY/blc9jFub2uTVEJf9p8oeSsVz8hZdIOJNAPD7diQQi3ukxBxGe1FRPIbloWwXE4gWiUbmvZM
ZVTu81RpczwVx84QvT/JslskjJrXNgH/rIqoxKqEzLo5tgbA1z5F98ZFOJFss1lyffV6fHAszW3m
OnMkbMiqAftjI6BDoOx0LCca1VbqpQC/881hM8LWAv2B0nfitnsDdKSmzO3bQOKhBHpiEeB36s+Y
F6xZxPucq0iS8BgrZJUi1V0BPUwOfygcyRYNslcuGBU5zobzmH7yAt2ux+Bcik5ljDWoc31EU06G
7XFhZIGtrUYj7Fb3+1xT4GT0lDoHi9N9ixfQXpXL+fH3XN7AZvRNxUdFQ6yGnx0SVeYDYDpS111X
zyZnDL3PZ1oN4EFgijBYksH2Yy8kq7j3n01ozzsf3HzaJvrWpytmFYlWk033y9mtF21f9KtHHgSN
t6D/n0fKbouCfsO9nvZ/aS8Ak+QmdFGe8/N/0Fi+2IhcQH0hkeGOWxzxk1S4fMCwF+ix+k5b2Tm7
nQ++iF3ki4hutcsXfrL5gRwaqqFsdxSLjJHOAG/R5HVqX3J331xFJn2aXd/h/jjZ10Zk9Tih2eIk
VleQUCAVhLYQ42R8cDEJc8ujAs3eQTlP3IBckksTQ336UCXDqaQaTcV/C9PlA44nr+6R9F0mbA1t
+CnNe7y+wpEbHK2kBN4soAMty83eCc894Q1YVYeNXXrXVHXwgck18M5dwwStvSBta0yELV5COJj7
CdoQYKfhkK+DmqH/+YlxjxNGd5psrN0okGxmYuz4PkXWVkvYDDLW7GeGhGIqUfG7V0t60dsVn/Wr
+gaX1uexAUQ0ULuiHExNSXAebMDbCtKoUKyvqE9kclNiSlQh7MWvpGXT7qY0RcTCwfYveVaPm6DC
ow7L+pvBd3KcFoxQmoZXocceRrO+kFqowgUjFWE5Pbq/0Nv6VfiofQgeKADx9nB6yEI6wFEcJSbb
9iu/ckuQ6coPiBlvjdTIjt3MnlXbtUkkAXnS55eZXe4zFe6r7oFGsu4zGM8OFaWvVCpxsWxlcLAo
PQsJvWJnGHEKDk8AgMue+zxBY6a0tOEbowgqnFWglZ8ByrWNlh0I21agbjGhycqGsBTsdmD0zRM2
QB+pvuGDibI7OS4TrufqW8YuketZ5BSbZQqlOh7YMxyUNI/ct2m4Ax0RsqJAO1VkQpLU5TwX+55a
f5RZYooDwZ1DXSbVBqyzgY2XWp3QMJLyYmd3F9slwa31c7MuweCB9Jqq8B0B6bfPNgNbm8PPpHGj
VeiTLucWqLSTW9NP8EWJHJ1L1i8AOz8v/DREIf0FLXI3KLy+5EJIOsYWuK2cPTNQkdIHrNXz0K/r
w0IJcV5M+Q6NjIuPozovH6Dh2IraTD/AnTM40//kFytdRb0eOmUNckpi7JQRXuEJndsZfjJ2DZ2v
igOREDKV1GteeXb9k/aPdL6WXoc0LYu7Ms1TB64et8eUYhmeO0dXPKkeAf/bE+njAyJSsxBiCxwx
JRRSmK8wTvo1kGZhl1asClr0MGGYJ5zYiCJFsYMr22dGefhIZJpLC8IhecyiOmSoDbbnWP5awtT4
j+yFfw6TR7SZVtuflU0Ma/i3yk8P4P9nQsJeK0bsh0FVvRZgo9mwKD/YhcugmcfdE4LBAWh0kt4w
i23QKcqkD65G2jnyKVZwDR2iCideUyZGF1f0O2plFF9fFg2RUIOr+UBlhcn8dvyFqnMwD9QtFOih
KE8CZwWauiKZO2olCjgt4AXcB8uPMFjR3x+Oq9v+RPMPIBx8TU+iInoLX+IxURel4MSU5dtG6tkV
XxJRqX9j42ycDgdsSNmNBlBGBMPY/XxLwbN7cxYDR/v4ugVaVGBxZPXPiLHbd0L4ZY9FJ4MrbAMY
Oj6KELuhIFSuxSwZc0PmYvf1FVXzUxL1VEbrjhc0nC3WB+Z9VMDO8FwAtK/NFxWcnrOCK+WbAiT8
qNBSAPx93jG4QR/hMjII+5GAO2MUmTZvL8a8QXCiGMA/hwL50QN9mdTPR3KqtUrksrcbPHcKI7kp
Msq95Gxe90qTzy9trnXSPyYyPG/97bbl4iNjoQAHMDgLtEGuMCL3jQm5JZ54jrdbcqN6HWdTu50T
s/AcpYdYM9F1eTEWP+JCijYI9kidcGVbrUxpuvUk/iQiKWdYneTY211KITj6S7Ot8GXFwILL9unW
gGoUZLFy4tNo77RzC4UnsWWo5+PyROE5Iut59fPPH6ePNbxWLFEjYlC8GfLuiTcZmUgDuFOS7i23
U86YbWDChRcBgQ8W4NhuKOZNPh3SqgtfChq8z9D34zVY4pBgtYef5Ffq7r0hF/xXhKTsDbZriQHW
fZJqT71AtJKou0v9t5P/yPgs8IpuoYTNllj68AMnd8Lm1KG8ht99l0AdWD2EkvYSabXd6oHbQ21J
sykOyd/k5a1eesm8fz30NjR5iGtB3ZpRhdcG9LhVcHGJ9wFtuTfO7tVuf+yIYnoEfh/0ktj+2sFi
6W3+NjdFua7O0d1Unv4ZdwwbLkIeC4EJdRLLxn4fJhwZyoQzOXkzzIBezFp4NXO2QdUJzH67gFhL
jXM7P9YNBVWyxUYkcOFXsqh6nN+HIGKk/kd/PtOU+A4CYes4KDRpYFFe5MyhODf3Hy7GidMCyCtz
CT+faE98g7Hfh7LZqQd8pBlNMGzagoYrXnePyWxkwrJG9SvVmyMWLBvQns5SEX3xqw7qeZpzcXsp
U1PI97abCp+cRMMpWb0r/LPrP+9VDmi/9BY5Ow8wq+7sZ2AgFEwOhTl/GIblbsOiQBB5Czx1xdwY
5LUVPeZLSuy6haWkGJf/NIXRU+e/A3JVbT2BDWYKh3nVdMBg4IM254fwnHHeqSO7+FiqvqUZ73gL
xkqKh5RIUQG8d81whWorAYceZxIomBfhq3ZSCLRKDUWywxX8OY0tvEMCxOOKqzR3x/p22jrFWRpX
BH9BotTssGcEtDzEKFAB9xLhX1dfiPJMg+yKDdn3/b0pee/4iOkhh04xLkFnU7rB1qbDUhTpg6oU
IBc/4Trr20Flf+oP2as78KTEtfxbVnJmNG0nXQSnxp3/BM+TrUSSGzsQbg/3S+sMVkl9KnG2drzW
o3uEw1F/prpflKrc9Tn1bOwu3oggNWuMl1jddPg3ala+497DEJcTM/1FVVv9msCZmA5B8TyLnstz
XPldEMQTavhIUurVPPvWPeBA33CzOyw7jBEEKNaK9sdgP7f3vkKAY+OiM1yozMMtP61fl7JYUqFq
TD9Esv8/qIPt4qCSxkwHty7yVXULjiKeoCdsq7eltudyBj/mzhTRQyCmc2ovCxYcNf5/5/9wfqWm
TpAsPnMEui3giesIIAKFqQYkIuWyELlcsMuWkC9jHdxiirB2MgfoNdHiHN7vzxMED4kIuKksCEwj
2yOoofkN6tPljaJX4lzUkP1rtMD/YoD+7wbVTspWJFgeYnWR7UgvQKiNGUqDRVkGYrZQQaaBm5DD
zRFofFkVpDwhi/J+ZOYsVGtmGj9OijAuIux3DwC1GYQpLdJXPmpmOYS504+YBbFsKF4K/SJ65Tx9
eJDKuADw3uUNewQ/vpHG9avKR8COz9tzbxnYK8YDKw/68osFqz4lpMfFmgvCfF4EkoR0iyFiICfC
4aS+zvi9DBXT3awAYlCNjiiS73m/JuSaWSIeHkNNrhtHrh6zhdgD95Zd6BWZPf6xT9szaCUEfldj
Gg1gCPrPwXjxXQ4hA4A1VNv9eVD+qheZl/ltwcQ4R+0LGAkexpNzRKtvJQ21d7Zex2cN2jnw9IBS
+U4HhEhtYl9oUQGL6Dwi34K97ovVWjdQkVfK/X2Bh7TE+NLQSS28ibV7b4dBbwtjWQIPFV2zPN39
1buRghhdlVDlgVAGFMVfxQ7jC7KkAaLOjnJS6C6vFyytY14EZBYeoHh7/o19j+7JYHXdAyj4vH43
3+uTxkFV+JUYj+5cn1UXjaArHUXUZ8LfQlrwheO65VXF9f/Eg4ugSWUtcG35VZ0iJTGCIT+ytSio
FInWYNiG5y6/QWqpscPAURuTqrOVr6+2MdgpV9dZtNw5nAEzrMQXtDV69fMO+5bL3DPVpSwLO90a
m84C3VII87AwuvBBqOnpqO5XA2zuOqP8AGfxgFRvNSgsHYlQ3xaCG2+KahrQFFc1Eq+njds4KGES
+qjhJA80bn8o1ZI7bGKVTlZ8f8XdftLex3gvMoj7xhBo5FkeG1Sq9XbwEx8SxhIBv7bQE5mu1txO
yh4DQNfASF7qxVLDVyajHDkGWEvadGa4YInuzh4LGxJ7wgAychNBGsa0yPC8BeRV+k4/QVUpxMjl
ulcDPFdy26/Uw+qQWr+nFh4oqRAcBvvmtJc+oCtbjiRUa1r5W4FFW+HP2IK/jvs+l8Vbeet3oDGz
WlAB3XOYWtcRgcVqvD8IR20JeCFS0KMmqkGdz7Cfxcb8GsRU59PUnJBdHCjvG/9LCC/HisHUTDUp
2/rHuwpvBVLimla8Z6zbj14gLYA/pKRAAaDJaVKlbg8nyWE2a3ilb62jgvh9HsXzhLANU6TTzIPf
bPFBKEaFxMgDODwoRXzpQVnTa1HdYBumOLUUr308CKq/782Z9Zji0eFpdEMdBnw3BJmzRrAor/EG
RzzS1Gt8d7MaQ5EYL6yU2ht3rsuSacZiYRy+l/uUjviR5aR/NHBx79Ke9Ud14Co6Y3meXJnaW/Tk
XMFfJXl4nQMgQUCuLoc8OJMw8VDuEpHSOmDnV0WJJosedgjCi07YsrkaHQOqanDwzh/wgVJdETAv
P23gI1ob0l2ks8rd5GwEZMFZbeP38WzSBfBU49H4FDVOGpMuqaXM7LjnuLEcdoXtJ06OcQlfrWf3
RucaIPGHB/cPfLAtS8fk9wstbRfe2kFlH2gl55FSgznCx5B8DkGkRAAYquCVthBC2STpQYQG9uqI
hhzrFH5sH9hBs3DH6c7GE1vHTuVv6xInD7xzwC73CVxLiRRZrWAOWKO3XAiBbYlGdCohuXv2JFNX
4MuISzIs0XAN8vN9sPgHtklL4iNQJXB17eU/9m5Q3sfr0aXpYHfIOqtcoS88GdZoDCOiHkNIfnLy
9m48iZLupaDQnpVHM8GJiqHl12tw0wIneZ6wsp9K+MGpAUxsBDuhX1FqaSRujQJMuS1hqsiEg+7u
s9BQwKMT7Aorph7EvTn/I6rHl2OKOx6dm8EUtmFGDoJTukQSfLSWhtV0VncV4qtbw8+BFpYj3CyR
soinB5WP0AQehzE/hORNdaSuFOpDyNsfGI6QXpD2MHGU/i4lI8nK4jHHHxJ1BnR3n11IocMnOFl6
jNFPgijhzJlUyMboSAZevg3hU8VYR9JAimcOtphw2jByrzyd8oYdh6jQukyGBQhoCLvRcISGOj06
qWc8UZyqfjNqGUWCy0q/CAnk3eklzqb/dnDPIqJdl7gmQgvJczVlnMlFU9+gBe9oSkKSc+wesa4s
Qcren3+5Tc6/sL0MIfEFY6eMqmnSWr+FaJn9UiUv5gRnHRIh69jcdaDpMLItBMjjxa7nezyYCVOc
Y+G0v7zYowIX+JFylA/N/nk1PVBdHYXauCpGINPPtenhPt0HZKfTonTV5dwro5QtXtE8Lkl5FdmJ
hj9CpYTrttbxlVc2EfZdMiwmRXGptezMd2PCk6H4lQfvMOtalDal46qQomK86hBqQnXbnrSdC1xk
narIf2bEoVpYCP8cKFK7xHjNSugYsDhMKL35eE4xHagff87GVMNQI1HSZiT+1XTl56/mr79DFv6V
+IsFInly/ssBjY1TYi9oRW6zhRNh05wUcmFFDy2EZlb2UgsGtPoXQ7IEgOkg2eNbYUv6F8TK5Fo7
cMl2D/0mh0le/AzHR6mX7oJv941cOHYx6niN4th45DtRQhut67F9rDNW3rzxy1WfWkpKBOOQrZmE
AIQAhcwRVB2bEZ5tQvPVpj1+5aYvzoVPehzKV4NpJIYE4dpsxkLptknlT9DMZyWzOcHR7f7eTzi7
rVQtqJ0pQSbN/mAxVaqoIxHZc8zjOSPoJNshva4k2DPd5srY6P6o2HdX256nR5HXyujuj8SMZxw9
YN9WnLG6hPHw/uLfk0i3vB4hYT1mftgJOG0RT8A+5M7+4sjc0IChFlkKAsI8rsAyGx5fPrH372yU
kEQ6Kc+Evdz0OzPHwqys5X08cmxisSlVa6n5lK9+4j5fh7l9NEvvIN4j9nzPsd7vQPOiDVNoxtkS
3FrUJSJGbpywXsbjC4k6mUHvkkwjGWrj8lTogimOhuV+rdCad5eWkXJXjIIMqTrXnczO/4Tsw8qj
S9Cri0aZl5rnzX28d2VDgNXsGDDK6iW8O3YrbyJfNLKtfVjQnrpT4c7iyt8h4VJ7GJQ0zjwEax6a
td7sKSgqwDJkh1DYXkyRnbG0FelkEb8EAwVcd1ijojj+8od57p7yj4ZIEAl04esvYo2jEUAxqZpq
We/WZLFy+3+JSHI7gMnfsasjNsrojOKPM5Co/xX+nMlpcfOzL77ZO3kx1P8Twe3PoJv/d/d0tEpF
XLgy59t8sPqzKmhQd+G7W8MSOTcgdUltkZ23KrgK2zXYIQS1hMaGJoyXADzm/4pN+Ilp0yLQX3Zs
cPy/OiDOnflV/0TwHlpd2ZeabzMBPP3cTRUfLKuOWxbSQXknmXqktJSCcfh0DQUmnQqPgBSBIZzX
6V7bmJuSfAaA008hHPtzGekxqUbItRafzLsjhoHmf/1VGaeWk5Yyly4I4fVjRfQ9CcYNzlmJb+Jt
ZDoZmt0G9nvZV6SktwWQyqZr7R8X1FPE/IsH2cutNiWx8GZdCKGyR/li5GC3cwD/FNLtSgk/NKX8
NVWdeyU+PDwMy833kt+ccbhq3CALKvhcWOrBk0zyHjMSQ4axXHzvz73b/0UlQg4thTPUhFthReOK
85wVPSVaWQsi8DXHvC16Z7BId+WLyuaJy/h44ospWbzJtJW8tK2FTQ+XtAc7qTMqTTB63DBqJHm3
z6JQjvoUsIKZgyNSkc5qhnfxjgEZHOchCP4ife4d7zH46VxF/MZoWqb98CgnXSfc11Wi7WC0AvnH
oVjM4/hMU68LLCdmn8z+M3C6zHk530sG8zUyPCrfXaR8PtkVK4B5Ib8tM6MzbSPvS8ob7DoXNta9
FnXat1so8OCSYtTSmv9uj1QONLxUhRSaLyGQfenCRakPQT0z5MPZP2HWw3Myvna0MvDP78/jgjhg
1bR/ecCYlKTFvxQYt54BBLRvwMiQRmHmZRZx1O3TEvDwkBMy7l1uZ6Zg/6fs6jDUOqdqawBbXEYN
bBSSQfU0+u5nxaZCw/5OEBqDPjWy4mRB9JPS8A0fT5AqYsJqam/7d5drjU9SBCn7sgh1XZAiAH2p
9SXz0zm0HkJfqhOOd9/pCYlveMXpLnYhGxktW+yDXMnPnzAlDhKiHF9D9FWG4MHHojK83dgNC1gA
3oIsB6/7AWz+0HBjbJAdCeyRrcFU6Gdo3owlZfEh+4H4SxBa8tXRqGarTM32ErsdDqcznfP1+lFj
thXkUjwRgkGi3ZGNqPrRUrSi8aiEOvUM4xUaRHjc6oDqJblm3j2bIftBpMWKVQjUgTs2Di5Uz55k
rhrEeBIsCgfCNmFYBXQVVDvzXhYJWwz8KXnpiiMoN8kK9jN2twrZFYUUQb4UVpHddT/0z8jPoZKo
oIDDyW/L568tz/48SSsAd6Cjzrd9z8a885az5oq62MI9LSWe/CazoMwzPi2bBt2vRnY9l1w8bPpS
4T8SJXPpNdUbyCUQS3ZA/AtkLWb5fdXmmmLN/bT8maEmwTilA/l7wrBatALDV5zatjiM4KywOGWz
cr+RYyTL95otmXRVIgkQD8bLXVvWlZSm9uU6g7dQ64B6rsWVyW1EQ+6vOhgd3KwOQHBOp/sN8c8+
YDSGxLrq/DDcXEk4TwejDRasNAd7LoL7j85TUB9ZTb41jow/LFOwmDN3+9ROvWLxxZFey+IGvBba
48tO8gzSP9bcEITG+1M/SNwqHqxpYaguJHSPFIOlAC1lHSin4qXNCBfMUcXRKPRl+xvr9Vq9OeOD
INWTXYHwBE2gIeETXBr7NiLhKUuRA7/0PLXjmCwaC7pVDw+UZhmsFSVqmFwDizZPltY+UuxzsCP6
Bpiy8yx7jYvmR+H91cgmQsy3HjUyDsm3Ll4T5/eT58gj46Awgrwqt3hZ9VBIdKKFNaaY58xHqxLg
Ws7GMgIhxd5Z4HhthjJAtrhQ5Nm5RSSLrQLQnNe02zxcf271AUCE9vSBw+CzZ9lDBOCADlS5sDQQ
BMokWWsQm1wJZ0u9nnVN5itTOTzPnkXOrJ1GMypUgCWZ3WB8zSXL6MPDW3GV3DKOR2Z2JMHW3Hkv
Wi2ArsP/YxeWscpD9xAAK9/dtIG2gNywwPKV8Q3ENPmYY89HeSQVxujOtzwo4DkHfTA/4hdEta61
3GzMcllJ3msmosGHV8ShjkDGSEV9GSgSLPhwZ+TL87WdmLIUjY12KU9BzLQq75gSV4OvxWBL9pJ1
xnrXXJSzXAf3hIY0r8DSLXFeEnzUO33LwhKye7DuJMjVv2E/gNWBcpXw7yXrzwWNkf5+i8E/RhCk
g0ye5bDpl5XFpbdzMLYuwsHH6Ymy+117okWQweowbcZSl3t8KkpAFBmWpCOzGQL2MchKDwicVRt0
4xxLDT2mypXfyxxB7XWg3mVnU0ljp+wzbDJobOWbNl96mOAkqeNFBqF1RcQjb6qD99hbwF8ZitTV
s5/QAPZfAlGUhzFYGLvfzugcjoGx8e05iQDJZZBm7XjyWCP9L6k9Gb7O0PmLyOQqVFTde7FKYUZj
eFVU9gXrETo8qU3cAMivZMdWuuT8MiQANWIeBUvwUPWfRLWBJob6JGgcNOCD+A6QviIPKdO8BY7+
0LiRugFebSj+492Lsx4tuNfJnoU4qRiS4+V9siOdj0nvjj4nEyC33slyB0jyCV2Oh9H81H1uv5DS
Y9oYX0RERsMXaD6oJzwtUFgVq24S8dxJuKpoSqJXOU207iHBljJRiMsU86vY58iWNdA14wHn5qOq
hvoPCgu46OCCOH1x9x2AYfea6lzg+PY2YefhhyMylk3sJzNzBXQM+h64uqtUXpHGxQnsqdl9O94j
0s6L7FMCbhhDhg7IfZCfXiNrLL5GReZugFPL2SyUw2fvUC3xu0tVK40h79yR5fPk9hoGappsAmrf
Flwitdq68NJYDH1CUIxiIrDKCJGEd8GqgC7V2WPHjzqBrtJWr63v2nqs+ioU4NB+KFp87yfdtxKP
tRBC/mEmOWLoBflrfENibJH6WWxWFzDNAi5PWgGGhQnugGDNBQMT5V7MDDdnwuDeofJl8QrQoxJw
aqoqeAicPSlE+Knt43gy5wg4fTKt0NNVpW5+zhXghU/Ff8L4IQ4oadv5FHABmHmXWlrnoXL9YlYR
uLAYa+33IGObyhCjtYjOKq/EJH4yaMHErCdcqoYgETt4o7cZuVD2NvB0x79CqmOLcqUP/kXQcoFh
51vorjXdE6kTzJfo41G0b6WVw0CpfFGvpZxghjZLe2ph5ZYwNpqtOrystnoS0R94RMlocGmaQ7E1
j5ShfBrygyr/oq7kIiSnVSCTlpPWK8auJdcmrB8HzZHxfbSaoT78wXX0wugeeYcqjgwFxgOb6uw+
WJFCVHXDOjW8yArThR5NsFA1bmU3HM6LOSrjmkQGPvs4DdgjmeOB4tM7QWuPWms8S83PX0FtDADG
3frQYI+hf6LsOcPljnusDVApjm7jVYGL+DYbIJydVNHyQg/NjbBvMWOxqxzJizXLH+obH0QMP8L3
SIcVYn7dND0/I3/awAdr2GxmhbiTA95Sz+5VFt0wtfNchmdmufDs23kVd2CSKkz3XdA4aPSDc2dF
fQvpyzmz4gb3pXpEf1u/s5jUaMszD07tJBQxBythrQbmrj4+2w8IPX7UOUSRCAXPwFkU+FqCaESz
t3aAQUwvhf2v5SEdNb61K3qFsKf2jyRCx5SqPkDN11LKMYnmNbGZUmDTl/HghorZaFu5B6d9rT6Y
VdyITm3o8+UyYpBYTNL2ma2MtM6IQ7F5pD7rj0NlFPbr3cyUeCY6HTAtyD8udqloWD9utkrbLzwo
GyUNSCpbwfxprpWCjj2Gyb50LT3HpWJwAMFeJVco2Ro+Mvi0C8YAvaZvg3+bvQgOTXYxXHrTxjMF
w0/wHCNX3+bDyXrINbkKWDBbx4hOx15Z+ZJ+ocG3tFAy8F+1s91ngzdvQ1xNj0TgyCU5pYXN6xlp
IlRTaGQfyQT0spNbihajJKh1tI6o6vQSbl1OXhqaQS0OnvScJsuT2YrqQJgXBRNwPVP4KlpI2/bY
NXo/1hjMwKktzZV75VpCaFkvpDnZoJezFyrdW13jUDclm+dekhf2f+LTfMpNnAbZ4uf6K3Qtv6Cp
Qlo/hsltvi9pe98is9Y+uH792Rn5il1Xdsp1FAGYSK8g3G7A3ROHcjr79oUtQjXYkb9zR0LGz2Wv
yvoAhvzkDD9gyM928eqkpG8NtctrakOUk+02W0/maQP9BXRGmXk3ik1bTr1Rnaf3x3O5XM48+tA5
jiT2hqtILErLK9AYDjNby01N+1Y0Ojcn7G9w2aEj51qTsHFh6TPAu9il09kSgG+6wH/RrEvx09PN
x/RmaDxVpuVf+Db9ePFVdd3zGSmczqzhc0YwAm4dlFhNrMHgGU5iDK4r3Ozv5h1Q3YOkLFztwppc
xgGRZbhvU3e46aAX8H4lsun/AEi5YzgK7kFmXtfcLCkTzK9QuSJul75qRdeeV8sHxVyDleJtrrZq
Ae7YZAxhXYSOeQTsMYSh7dYoDjQxVUzTJCKVb8AXC1jCdItFyP4yGmCiRQuFHbNEiBICAtvrUEul
y5I4a1PwqDj/4z7qAH5cYvnwz4k6BQLeUIrLkvcfCvfmmVdT68xvcpGSnDn4YeWtQWhxvgJ5UR43
t7emDv10yXaFj2ZW1CjXGjfjTOKsMBTaoRA+/fzOywNRDqaCDJ3P0vPjxKYQgYnHvzCphz6QJnws
hSghA+cLijgEWvCRjdu/WWU6Fx0vV783y+xQwQYlKppxkZJqMgnGUVxFDTQsZs55a60hsMRRyhGd
bMnUZrLUTTFQet4cZj3J3XEvGD0lTijSGHQg8LzfbrwPWhcYCHTH0DSaMKuQPwrYx2airc4D84tC
4DOam9SsvPzTQC9QO6okaarK/cukfqv2OsJpa0BSLtBCQWgfAWhH35MhT6gS6KELdfKkJJand+Nx
Kkc0JP3EJqx5mEIKESoymqFzkYhPGACI50vdmAtJF90APXHP4Fe9klpJWaKXsVyGM4AZh0zMEEFg
FuH0XhNOXb4D2ykoZbIptoJr8q8HtHaCk88DvIaZ7eRAnbEpyrz7vb4hpmYQ52al/LscwsyUV4NA
9qt+yNzGCkAAdd+bjo3D8lPH+H53zjd3UrKIEAD2x16dbpR4pkJUVlDaeSjBiFlqzUWXYxY8evhj
s5inQbFwsNfLeb0iPPj7phluzZ6DxPlmxV6dRLZTgMZI/e4Uv5G8wbewGCF6uiKTFHThD9Bcdvtx
3VaynIb5NVy812gTPkTgkusGxMVOnaS0Omcmy6msf6fYYmkj2A9uUJsZilO4B2Qc3zysqqJK1zER
wAcQRoagnjpAW+SCUVt2wL55Rar0ijGzbjDhMjhNVy1inFG2PaQpSEH2k0VOVQlXDbc0+2Gf4kxe
igAsoGJCe9W87Yy49kZ4aDTBWWhum5XnNYXEtRvY/CQBRftleUOW9XoASWtw4FPHXUVwYsk0S9AF
59uRXjT32MGs9m668Bfx08y4JApCYhKD2edCK3gHiwVUTIc4EV4nWzwZgZwFBnJ7olI9FrcxPTI9
45w4Vk2TpLtGosnrS5RuThwohWeTaDlOPhZWovoSw9H75Y7v/4yVD/KpKBXGsi5IOzPqUxlhbRBr
SXOsM4PqnyzS0vbXa2YUX2uAn2OimNyM4iS1PDDzhjkH2wxKZ0Pe/wwWYE02InJTO+cuftaO9k6r
pu2n55w0fW5vLIv4JwIRPFJXtbnIvq+54LNMA4P3NMl1tJ+lP85ehEYSmoFNHUkSG3Wx1Cxtl8uQ
lmoy85QXrfzkcGtJzlv8vBGp+pr05DY04SBWxXb66+Vai/TFxW8J+XgWTCgQqfcBXgGUE2S4nifv
euu4mRiPzf3QWlAbnXPE42usjwHvX11CI08bbwSJeVBHlOEnMttH8jpi4RDrdA51gNYkhaNRcg5l
mrnuSo9MIdDsl1Ueq9kuC5X3ICRTpcW9K3k0SzV0uaDvq3bbnslax720O2jKzfIEA08HvMBcKLdF
YuTWsuWUY47NX/5zEgAPNDCRKC60bV0JhoGnkkviB/Nll31LNSqwjq4PCag91XJUn97C5Dkhy9VR
DSy0ssk5brrteGm7xU5AzkRJ53ECFgDRo1eBczLajJAhVdcHolUQx1KybmeIVPDcWoUEQzy/BbTp
u3qyKPC4wGP1+4lhf9P3h8YS0ch+bQQIb+NDIxle7iL2rK1u3ldgs29yWcp2R3No0Tzwlk+xEys0
9JaZeg7+A9I/bKZjTKcG3a8N1c+JsJtnkw9E4AohlZy/UFNK+wqdsToq4/RB8uMXVG8FGTaAy/dn
YFgNsuy47eT4IvdgSMoHO6bN+Q+2aC/C5y47651Ol9Aq7BRC0yUPPz6f0zfdKeET2G+XaZ+9LbSZ
spJBZHIHWfznAgEpmIivGqvgbWtwb1uvU7ZW6y0tT3L8slgqZPgRNptJyKlpAz/efHi65ERVglCv
3aEz+B+G/f1Or/wUQtWMuRw55rAbavo6XOusvpb7MmPQTwKHeIOGtW1G+WqoHjR6eI73UBE9kFTa
+Kln5THYDrnE5RIFjkWQIfHcoP14LX0mSGo3dNjD1DhC/FGCvrXFltKgX3eXoW57/FGgNU+rgvQ6
k0joM5vvyGKJd256SMnJaEn15CXj7Z7ZBEkQGcySuLrjq6sVzxD+TA933rkTgCGtpumjz+FeLO3C
CNqNriJc+N6QW7TzYbZkJVV2FXWqjjAASSNjA54wezwsg6QUAsU+mknfrx6zjUR8d6Jn9udA3p5s
BGCL4bwMndx4LYGhfk71LxsqwpKlri1JCeD2jXLz7YsxPNOx9ICwWTuSIMBIpXOdhR+mlR1vJdPP
56WuMtHCF1frJFWWUH9vpNFRKFN/nCuqApKz4fpC/s8yVpvm5FLG3r3Xobdfpb2uo8X860jnNSwj
mGUWL09qDJhgAaurqi+UqFiysUH0mLu9gz/zXhjaqOOdSIKaZfeHG+7QCCFksIaZLwIrGQs50qi+
FKQiH1tK2tKF7eSGcuiD7gN7SPMztra0HYeZ+cFlW0OEH5N5lAElreKP4LFWucOqTCVuY1RJ6xwj
7OWVDhQYFwu7iFg0ehzKLx2DhPRS7RECMNODbPGFN++swvkM0RBNb5MahVj72bvhV7HHIoVZa0/s
mrUshFvbWBhMvbzhVJB0ImtgQDRXUaWA/KAUIZLQjVMHcDwqvF7TBAnlbtKH/D+zz++SNjj2Ra4j
YgvVXvXAqtCQDSIIHBLYg99BF3QXJ+hTtOrWeckEpPKeX1UZB3b26m1lCVnhilIkT3cu1lj+UOud
FeSEy0EzOZujuO0ExFXUafmcM3giycVkNMNNJQQnf8esKv8BhR4w8RFnSfKGKLkbiP5O2emrisRv
qqXo6vr3VCAQgTKswuLbUDQgZCn3mAye0+UC6DvrJKztCvl0zOW2B9TUVwJbDzdU+149sNqo9sC5
pZ9sXvuOwIra1Fk3jy6JS30Zw7I/EB5sKVTmuZWnb3HMdMYq2Po2BUNpQF/f/CZ5WXEbNPaceMzG
3dJRo1MaNU8AVmJv3ix0n5nq4bU1laTTHxnKT7NMGHlMmcGnHC7GOhHBY0xqHDopE1+AMomVLYX9
cHtuIqRgpk9r/cpzfxPJaakQUHbKRYKMTQwAeCnmfyKQTvpDJExLDKJfnTEjjGmaT0A8T/oVI1x7
rwNUqRpg17HTTCUlYRHpwjrdRPZOKTWevovgvLm0Qa3jJPRuj+e0WnyBv/slq74+rsFbM+HoL39e
qtGTA2+i18idgTNsbIwXUCYPMUvgI5WxJ8U3Y5/WSvOX1QrbsmnZZSuF9dWBvMFbTR8Vmkge/mfv
9Kr+f06dR+0p0taU9//kKTkxB7ZoikiSEWPUon32OehEgr52VWGgWwc+ukATIkjMhwQ+nMDL7kRS
cn0ERqsCw0fhuEWfMYGeD0DfuiPOaTPtHN6F62hZci6gXUQTh9ZUX8i85x+WwjFWl/VehKRJdFcA
64HNA5hjhIiLfsAuc8D3/XJNII02Y0i7VDeb2EZtEGfAM6c8Glqjpq0LX1q66gYg6DsrhW89UkY0
JowDlO1Th1xom/nw/KH60KENRUM1srmXyVXdbRPJLt5+zrpQMv8/LXHtUMWTnGpug/ErXR7VAF07
XL6L/ioPtwIzNLJ294rqFHqe5pPnu5hak/mXAQtiOXZqxiWCk2sm3JY6cU3Vb6+gJoyP41oymQ3O
dCzc5N2vRtG5G3E9AY6crcgHYT741AW84EfyTOHtqRKwaV3/UEtU1n3hOqXSYnqwWtDhbH9Oww1B
3l7MgsBcpC7C3ErB3tn8pP2w1AINEU/Z5li8j4JE46MYzuG6gy3XhmdRKRtNiM5VBRZ3cfzkhjbu
XKGu3duJKSdWDEUrbilxksM+2lr7cNshYjqAJ9BEjEGH5SUhDns1xvm3Ynzxm/OOr8H29sn9xh9e
VHNmAvcKP/xnLmxDCDWPxYXsIdHaOb2ctBlf1M0f15Q+eVmCg9UEbkmKfvNtbRe1sNyw8h5piLY6
5X5KwBQ054p3NdUhZj7lYAoWUbPhLQX/k25c11h67wRMEP1Qotp+S0/qb7/A6Ewjn/XaLHIOxlCy
DCzXQTuoLa8gJwl+u8o9Z2HBtNbUSuRZXCYZhvO8NIgIzV1uvU9VmOcc9ZxGs5tADYUI3FE4Bhmn
2hPLjvSAdeWPN+SVckoI/eEz7L382qTjp/1Wb3/kHio4SupAoynJtUVtjdUqonfjiwUumoJz7dm5
9O4QOy38KewtzCCkGiwRuvMzppwnzA9+rwoxS9FA/R/dSb6XKd+E/fJpmXP4MH5Iuh5saLOe0/4b
N9mdVmf15TT7WLTjjKjb9UDLrtWcSnBye1BLgRnAUZZtjml27MU4kxQuYVG+Noz308eLMsal5FDn
eK7P1CwxJTIJBCjwWmtkM863o1I11w7RUoOv2KR44n7e4CSumzvd8Es+fvIp0auI444OkIoGJkWy
nOpVaGvvsoYN1OE7IEd6j5OFz7GzVg7rs46RuDM8Xr8Ob2z0ZU+h5gRtTnTVKwslpKP8HDSp1JMR
OJuJLV0UAVZBk8WQTzD6m+ckzslby3oPOAyrgLYSC1SQII3BXTi8nG7Kt7jsS/CY0oRYfVDmrf89
J3dbAO1WVSOCThVUN19E2Wk0TDs3Bzkm3xtxbNF6TJzTg1mEoJ0/msATpNjtA78X5DD1S6plv1Qg
mi2RO1cyjGcTRtmAnLjPMqPfBQSBMujHDwAdYj++9fnkzx/0ZdH69fTyQ8q50kzy9ebUb2cgPb9E
hZkJZfb1QVg34twxWihyjkAf/kpfZ878kxmW3ujwsR7zfJDWgfSTQEB3PYHVLXxYsTxAc/pMSfZP
hwlbM8wERBu89gJeNScxiMKvSYr18OQzMp2jLlZeeL298Pj1uwnqFQtd6ASrCwaFjwTbe0YXXM+K
n+NaPVs7SYjtjEsuJhGO2WZ/sGbziJ+IHU5BbqqLEf4PPW8l7bGFDt3sMILDDxN1Vbtucx0y3TP2
5MH03+1TwueNNv3W+oS4oScQb9g9fTZeKxJga8g6RQFj2hMQ9KSi8AOQLvidH72RCvljR3luKVQc
4n9tmSimVsL9FkblNCD14fwU3g+GbcXDHs5iKFTXzG3czekpBGaV+uBQufuVVzKRZaJ5+Z+fMI5E
UbGnva3r3OrFyFYDcP/cFsd5AvxTbvzEg8UhJhEAZTRqqM7WCd8eOLvRg9mNNpsi7rg5o7iK/6Fp
z0P+1Bqzau2zu64EpDHPIQao9u8qFTJr2tO0YsFo7wnB4+N/HcPU783oMrxC9hWGTNZB8wTxByXz
uUP9I1LD8x9W4fuea+msMN+S2BN/dG55lzVZvNAyZH8NXdkWkeTjgt/7E6LI4Nafjq192+LQZgWM
XdkabdebLY5n7UkDN/aPUVUnbBckjWOAMq36cvBbazZUxdfgudE30tS6hOc5uySKrmhl/81VH2zn
ckGykcZz1Lugjzsf1Gw7wa0gme7zV1Mpug3qYCn3+i0Kj7/po8SkY1M/t7YVJ3uU2uq/hHsL0+Dp
1yjqYEgkq59iaFw9786aRYV4LnrFedbJxlqB1BXea+/3Mnh7XMjzvvsg0V2o9Nd75NBoOcweucMP
1YBRFg/GNckuNOdvo8C1zc1JvH3eY8Kn2T8w5emm3lgDoUCKRkzzN4vEsG3gNNu0SCxLT8ftRfdS
hLAKWzDS8MqsGVD7G0ccOfmzf0SO50C7952o67cwL512ubAVkzj/yUHqNqPoWjw9NuU+N+46ovN0
YcG5qyjM2q+D9f8o6jXkmr0WpVl/kxPp8UyfIyoD9ghnGmvCuEFLjmxQ5gyWdhJ0ZdtDM2WQFk8Y
3p5iGythwGejBKw0fgjp4uMNsZlisb5rGmhXYHVf4wuk0XyPONHTLLVv3AeDYc1zT83ftwLp0i0Y
v3xxpFFkDSc7fW1INFJ2TLZUsjJDkocXVv3wW19l4U3cPU5nCe7g0uUdF+CBERcCiOY2QuFzsoMh
cZZuRcPHbLJTMS6SGdKitnbFXWEwSm8327Va4+MpZOeKrh0tGqFdvwPQ3R2TJOkQ5a8iDjqHqgyv
ShNF3DrWSwnuIteCBzEDTNcBUIH4MHZjJr1RSMTJoBKXip8iC1jsIby0fI0F9RgG/hni7rxe3jHN
DB0FJA0F/3IE0K5DlXKztHyEbGCG/VDcp88ShVsFl7Tqa1+yoBb0MDOfMqTz5/oVlCanuhm83CtF
kuEex5oR8QK5vORXNMCYoKB0oFAAK45BfnrhyCy4BZEpIHFFX8E+9OoowJmNeCbWE8DA+CXzvGYF
WqBhQFC65GgIOLzi9IHprtfb1fVuYDeHm5wFG11bbCVR10I1GQM18+uHrQfrgOxishguM/1PAert
/IuwmCcyMuh0g7SuReV9iKBYL6XPvMRZ9Dwd80P+sl+UCsnq7Lhf5sxovZ/GuPUFaBgj0QhYoWXk
4dD0vJVuCFC42UjIiQ7rR7I04U4O52KhnzNII511yNsPRuROt1fNi7ap9U1hQXFpz50OYIGhniU4
Qttf6MXz0WWSFynnM3dE8TjRxj9/Qk6BYPk51bcUnFOmHE3OMRqVzWyegBPlrcVzoGJ97mN+oZDN
IOP7HMNlXVKY/yc57NC6GV0hfcVEd8PanZZaIwtKsHiRnFILFGO+vz5ZfzzPwLCYJBIDx1QHDfT2
l1GlfPHeZqaOAkPh0Psbl0qXZO1TOdzAgGD6mNH3mIHthrdGVsBoPZPbM1aMTHhXmFSWUD0p+dUG
p0Bk0KNkS9u1yR4AQFBk8WjdPC4HqJe5k+/LnMq1sIx2qOJd/86oSotpdeYPmikIYJuo1aoh8b0Y
KRMvMMI/6g3IwTUOyjJQPPuiyBzVl7As4KyFxzDc/8lSNMePpme7taaGEjpNFG8mETmjrB7jEdXJ
6GpmYZ9qSVpe2FqJ0mZxVGNs6hE6HPS6g9ThSe2mg+i9D7zvLilTMcyLwmMkGpLdu+pBPY0O9vei
MnmVw0SOiwLLlp5iG2m7awCGhb3VqzTD/XLUGLJdqnXiybGBFLrn4Emr7MZ8Zk/dCp0SBwWlis46
R3ySUlNNB+NHKYs1AH1YQn7F3GMlP6IW272g5kDaRb78wkghR8/U5UBMowTg6TJhnrdEZW07+oZ5
m3y1spslLtMGUyT1OKPQ+dk2GIgwymgdpNahWUqcyqIUZjBY1FawYmNxlr25hembrcTFkYSpXTvx
BUj3ujoDiScowml0eyL4lLhurRBL9deiM6v+lM3vAcnYiXlwKPy13eU/dL2Y177h+3aQ5r4LvYU+
QRkvyZKx90tPdov6YTIhTWo6rsRyjGkcclcb+mBeqR+vFlAGRYpZj0uE1lftZxhEgMEo8S0uIKGD
kELJn/fgsjq+rsbbziQ9eVqa88N+oSTfGMIA40PuKYRw7tK1PzEzJi9BZGxpWpztxryARR78aeVm
sm3GfYHoeNtTHKnJ5dwusv4AwRxhTkC+fMBubyGXZ4o2JLXTxifXseF2lDl7ZOgNXbG1mRn+K0Jp
a71nkZDZWBGhKbmDD5ww0Gn7+a0ZJlxkg+0cFOGAV3l9Jqz2YvJcV+LQwOYDZCfAdagT2W6TEaYM
ge4tbnYBff1TJk4OUtwutxPquQnOEeXMmicR7liibypOQ9PJCvraRBWz+1ahcykwFxPtu8mG4nCP
Rx4N3f5JckfCwmN9AyYK92NP4IDfhdoFvOs8UwL9C3Om7sKR03xy6vZXahRTlMLis4pK7+MTkWgU
F2ynXOWt/fvd8x25ZSyw9FU04u0SRqVRwqMtkbcKgvbDL/UctOeB8EE+COiBOjnju/eC+k6FdZBF
A62i3FYNCk/Xo4hlZpLVbkrpaiB7uGYe+osa3ejWZpsxWlrhmLMlWHh8srmzgt4vhsJShS8R6+s1
EV7r6BfpUIfKSd3OgtbY/FWxMGicdWH2LqurXpvF8Kxdwb2Rl8DbsDy5xO9BZgG8x1Ha+Nk7eobm
dNlhvhEvufVCo88557MPhXVNrCHITlww1L6MgGDvUz0+YzyjyICA7txvsrATUWWqqazn7u0mFIVV
U5bDOn+v8cmYQp+BRSBFKhz/y0kgaHy0ggZo+zkZUaAgWtzsRXDrX4HHUnjjFummFvrOtOfjuklX
oEcg27Rf6mhZfMQoXoXQQwC7tNrwewZHH1B/kRa/zPY7FdoHtXbBKOf9rNhRNkzONLEzWV/NusZi
jJDrItr7KyMdgaH902idiNxYDY15fG/d9VOM4OO7y2wEPIqN6gmrDB/b34o9JoxDktqj1NpH3rq3
4hvBHRdnID2pDp/Uh77XNlqU7zQmtMwrSDO1oLSs0kkGtOCX9nCZfnUGQkEBle8HE6xN34rMqi1H
eI1cQV5ayIW+PQwPkjvlnYG3KvcD0pSPq1RcX9r6noGasZL1T14ICoqpEHSqkWfoqPfYTI4tWcye
DOgHnxeSbgqNUGtwrrkgH/ycXeKl5vUPTen+cAwiMHqA0+gIp8fOL1v/GTBbg/7GiMPfZlcSk71X
2iFTC0UoCP3NqW425S9+861l9h/IlsE+Db3OgYndlDu4jwYf/2yh1TGXyuL9KTsstlTG53qfaBmH
VEpwVHGYK5kk+szRfoaLnuxPZlBy7U1FeRzv5EUihODcQy8FYx9Tg+IR3DdcJUaoSV9iKkm3GIKa
WuyMz6Fl/vlmUWnOtXOD7GKJUXVc0Kx5V7XVsxA2brWnJQQ0JiQw6lVmoNKmyCO6lOnRe9n/Klj9
+U4xvlLbksC1fyyVa/L/AHI8rnx28QGy7jAYJgfDvRzOPL2CZRdhlqUAMpKKbVQBBwAowRvdci9X
TJ8+j57YIVuY+EfvSVldNhDtNBvey0spk1BtJT8fAqphamtxxYXU0BWzOaES8QenygmMhKhXKDFe
ktDZfJI6Wu6nqpiU+7Lm0O7xnysAyqPBOkAicRjK6t3LMcY9mxGZnT7ZclenK9uhIOhCuzdOzcx/
3gR59zZF8hmLWHMnQBmMBOvoVbZNmHeDkL+ucHqtW0dPf5ep5D78oesZ3zj5FxhkOcq4MKL4u0Yr
HbX6UbJtRLTR9X8DfpxB5r3QJ86QLlwvaH00NVpiY9Z7XWaW5/xPk8vNb914daA9kkPe99K/WdUW
HaeoTgw43fn5DLHoucCXYPk5hc6jn5WaBi+diJIM0c2cOYn0T4f42yHYzv/8XWqTk9SYQdfrUpUk
9ztftXF/OgPxbZG0jOP+zwI5NkuQgfnnVAa2y+VQUbLA4yFkIoZan18urroyGnymWMkIP511ZY9V
BqXfRr4qPkCkCRVp4ajKWtjuVm1kUfBar+IqjW35xYlIH2gcGNtkzfs1aQNWyyzoBx56+cyVTBMu
G96ZVbsD8S3kkB7KDJLTQ27ZsVGFAW9k2Uxun5YOjgMIrdG8v6MPddjy86E6MNWE6S2w0KlJ5J/E
zBEaBNpOZyEZjvq189UWflcF/L33ajLAxbeyMQhOma/8Ck7UIBJrWUesjCT+qtF6ijYn+HxuwSg4
3eR8dhdKuEIckxIuCVF/QJ95zWkgGsWEAL6niJjO7ruN+SMGplLDHp4d5BQSp4/4tLGTx4zJ3nui
1BR8Yu0qZXO2Q87QBwA5KxJv6Mm6v8WEfNvNpM7YShMMeMINinpCXU9JWvFnFPZ9qdoxMUw9WfR8
AhBbJfuWwDF77uMfS8tZ70CopAR+oF+mXd9HRJ/k5u+G9sW4C9UHIAlcObBgQajQxHni/KvYeDhF
WYKlwmxSJagL22mtlFQKrCcA0V69E6HPL5xolsgFXC6NZo94V8+6Xk0rh7gvFybnI4Yz40ziEp1K
/YSmlLr0o18/xazLe9JSQ9vek+GEZ272TBv93KKgGNJlSdJ5sTASayWOqeATZQ6Bi71o8Jl14PtD
Vy9QVtmRMSMFpODWkLS7OXBOt+SPsQupzjmqg1zij5Lm+TT+DBDHNaNTuo0GaHCct3aTSxUW+Pvj
nKS3y74bqxQMOjzEa4CbSCj/SbVIJQARU8jkLzeBMp8OwJdMsjtBM3oBqfVuo5ZsSJFiQ2nK+7vX
qcn6eig1kX06vPMVIkKd+dlkObNZaUugrVOr7YF384g+7PCzcQDdMj6y2B+/Lf0OXOE+orWiOAO0
eew06J1xb0VXeUWluURijjzrXToUYAc8X7QXQpFPWPQAlhXbyPbY5L80TAU38IfQ5rI/dq+xbdl6
lrzfpc/q4TXRVlgVEqdagu6sh9At9h9tATJ/OK1eiv0jyO3hT4zqqBdPNH3i3LvtcYmpeFAObT6j
AI//CITRlL/rYN1fQkpiCHT4migfsQmJ2Nan6HBuBhEJtARz4ossotiyfiOCtQGX67qmbUrW4hY1
AroGyDaHmFJBOthdVrDYr66owi3KoeIKGKjRryWuum8AY2PLrIJtksACqmFg9NtDyqsbEtXOmk+b
KlEVDbKTBI4Rj8ZkJjHA9CzEcYz1OJeFautc+OF9+BVV96dtNs9RveBK8qejuqLH/GXiF25NhdpD
crTTDJWhJ18BmM4J6Ao/MP65PLlNrml5GbJPdOn5pTrpRSmIXUap0jixXMLECjFLbTS/t6H8Jtpp
mhuB5rPJS0qaht06paskvD5y9SI8Dx4O5q6gLbCsnsHyUxG5rVGd3fpjBpvitUvftuxIJjTWALf3
kmnz8dOcl9mR0E6DoomrR8wRz0LNNac6aKkbu8E39taAp3DPAvrCHWlqCVijC3g5NDggXPORNe0l
g+NviNvlqNmXuxphpCtiYjmVLmGNMA0uJ1mSnAP5XfpWkSQRl7Rfx4pLjMsjgcEjsFCcBwmX1OnB
53tWRQah0bI0rj+1G8/thjmvCCw9OkutIzQYY9ODqbHe9kvAHJM89peNENg935NFRViiwxA85vtv
jTVYXf5rtEWLg/0G/8w9ic7VE90P5Da3NFZxH9TBKzs97+8Am6nukWpo1Ip3QduztankcvzI+k24
CXDvtumU0uvxXinL9eFeEODsQ6jwMptFhjp3yvlcwXjY3Rg1hjM7nMVw2FDVp8UQQciduzaFI0Qv
3zfP+Noso5AaD6MLiO0kALUs/jjIECQhzFyBMdpHqp0yVP3uN8EdmTPkxhNbtrBbXp0QixqdX3/w
V/Qyx5NdwWWNfwP3sXwiqTxs1HoUole8CMVxJgioHNQmIINYCkZwKrSuraAQHHuiNQ9+i6fKRAHD
kl+RuyyN758e4IkP5meNfSjfeIQ04Jij9MujsXtGz+ZwW2qBPmeSuuWf7QfNWbLuOvbqf6KhAF/t
i9dqNsPhkK1tVkPr0HCsDLWUs1LR19eqNEU4j0M7+UcW05WG8C9fYyS1+0Mo1SXEJp2QNu1quTsS
y1yBQKQp0OMA4+qJ46GwmSihteJNRk3r+iGlez1eDVXGsCtBSLCIJrD0fXwrWqFdzrs81/JfCw4s
BdtErCH4lH6kth5qlTQZWbKxUgMYMA42crUWMwXDMa0N6siK5bPLn2yGUOb3OfG2ed998t7E/KNY
ZSX1jtiLT9Ke4Oy3mAMwL1kqIu0bwEuyuJkIUs96IfxKmN52vwnud3qF+1AY+wj1fzIz4OQA3zoU
eiGChtWv5ZsUwhkYSsW7NYbr6MZDyJwCPeOlCB3d1NVDyaSDu+E9xQeND4ao8yxPyvx5Z7OJTWk3
ylCGkO+aFIRSAhjmooc855gCvA4PX6Fa2lTsHkDwvsQU7WMywaEBgITytyfDYWqNVvVWTPknGajI
VB/1K4ZgMkTGPYRIA8+Nta5apEJnFhkUJQfWtWqQSfYUIfzqTRNgCJBkFIbFYqN3yG/D3i/yy1bc
ylgnP8C9Z46FWHtlsowT/DPeW3++hb/wj/+EQ6X9p/cZBWdzyTNFUq8772ChctnfoU8kPXE1MCi1
wvVMkrCvsntUkFUbLLRKJlWdzO19GcQPAzYP6397kKvVsWvNQMm3vIxf/wB3bJ29mh6j04biT5Cv
Ayo+dAudNKXLzKUHixf/ai1baSn9Dcl9Vnh8y8TC+/Hh4j6rRQUMAQTqyvV3kX2stAj+SLikMJc9
p17NhCpGkyCTa5y9hEYiSYjWgI8vhL+0s2xG7fBIsH5kR9nPCXi4L5MJrtJ+ETONaTLUC81Dxr+C
jGA4jTw0X4rhyr2lcgYLcGixu9lI3wn84EiqPLEpNtIDOiTnSg9MbhLDuiB01jTVXOl264JGJeEN
xYpqQJ3byhx4JQL7h7iZalI4XDlWzOkHlj7Ct4wDI1TKcXDOFalcoJzRHABiGm+sKPlmJ6WoTRhU
hF31haDwKdkv3DXgu3Brj+fwcwPs8QrPDzN6dO8kUuV8Gwh/ANBSpHaJLkJNtwkGoXj+ZwoZUOPe
u8xJba8NsSMRrobCwwBRmrYQ6uhzxMMXS13Inhf0eeA2rXojg/eIc58ukDGFURWwkOIL2xEH0aLF
r1Nr2lQA25SsJvBQEdu0nUyAZ2mM7yFxAkNfj81cKBUVga/lP+yuc98M15/Vidb2UN0C/iVPoYJJ
loHgEx5wRzidmWnJQazJyF0toL1f4A/n3HRn/Uog3qsynC/EmzRpyqhD+gdoZny8AzFAHpsywtI6
h5BlAibQM8Igz/E1maw81XbqUYbw1UQ/WsC3ov7SLkM4cJQg5vCAdMC8Vzfp/+0tUyzLwDCEiaoj
sZ/fy+F2KQTMBCVivhwXqjex9l1VC6fFzoR7uTxu68+nWxOWyKoZG8OM4Fe9YytePLX2BDQPakAU
YhzxsuUVZBZrQfK5HmiKeFCKFAK5NWZlXB80GYeLeOId/LajcxUpsNjx1E3dnJTwgL60dVV/HEwZ
b9kgSedMa1tiT455dnPgCMRBN/HOlfo4X6IOXOjtITCNViMRMhCDurhvlLwFMonGPMk4sthhj0vf
DJmH4ViGUF1dnwwhNsabbkBepoxAOB9bhKj7ogmK9vVr8MHqZ38yxDIyZlJiA+z40K1RMuqmgMbW
MANHxD5kApm9gAqvFDQj18Rn4AXpzYQqJnjDcJv97Rg+8OiwJE3LtQQJdk5XcwfEQ/yN+/HR/jBr
D4sRdJsAIo5rXLcNPW7i6YU99Mi/Rq9efPGEdkBYb4oK1zh5uS0ZC+TIccyAQ0F7hItDE+m/hMYq
6Qu7i/Ehzo3gtkNDd9ww4lY1gaGdb9wf2n/COFke+vFg0v+8qWAF8c0lZ/OBnPOlCcvIRn50kooD
jv7r2oS2B+NuXje2Jn/ikHoheJVuX70p1Wtbp+c2dnYann8svcabq/iyQ1LdPrD41z5FLHIONcGL
0O6XzbGqZVxhgkRBcVG/6m106wnZkAUEtZyIVYrnponbyeHW36WuRFDtfrHyumvqHrUX6oFx77kv
Di2UjZo5aGPJDRkQJiKhkB5YUB4jbn7C1Uk1tmGd6ezAKuzJLmzV8dEt7kMFK2J9yBILN0pr9XvW
DO0AWx3ALJ8Cv39kH4DgylhdVh2ioE/mA0jWh33Ta6fNKRUElcipOjielAkRN8bhAFQI2Qs5owAQ
yVNYnJJAGZwEiwV4AMaZ21495jIWbJvFk3nAGTMaCMYzQsxks/lGpgWOa+kViIdCp4eEA9VT/6Cg
3dhHVEDojhC5La/hHTUzsVVH7eLNzKm907C1TmvRY5eGp0iuBZZP/gUaEBMFlvpthOZOgHMk+qki
JD1sQDj3fTyAAbK/qKEcgff73tBvvSG6rAbZYPKXBKV6moUV03LZeRz06RkxQl/oKHxPI0NlclCN
pNaukk8p+0Wc0TLpOFv+icxfLh0IfZYYIIrLCgyMwLZEsYfKVcaz6wb4NGPwS1ciAYc32/qY0Sn4
8qt7S2A1jsbQcgdWZbROGDb5rEhpLAvha0Fcdms3Wi51RxPt7tL3IyvjPmRh7fJMVX17AdJ1pZ+I
0vG/I2TqHbqobdQ4aCVeBBFee2PTnVEJnSwiTilGLi7VUw1KX1cc9K1dpj3OgayER+++Mh68Tx1k
q6MNzxLbJdKteGBckwvgZAvMha050SKN4WZjtxzLJ25VYHGz/MQ+waP61M+gyxRCvTa5eC1RBruw
10cQ6FeylfTxza2OC+/RHbDVPmKgtWkQcF5IQMomrrHzyeQk7XT7/7hX4wHL4q9pvCn+fyGZm9W6
xvjXn9xniYThlJb1YSjhPW0R+z1N+70ht0Q7WuRr7FxlRKLEqJYBGRW+O5AuLbL/aDKNwJ7BEFfd
hrBZVDqIMP8Bijaer/xolIDQhb4vn84Io9Zwf6ZJLN1+P0xtPk1FM9261CHBhjaAcQBc2NvLNNck
NWCN81OZDTfRJixPaHVK1XMBSqPrBiu4bYsmQwiC4BHK0M2dS2PboffVQjXyELC0X9ZIvQ4Dc2ee
6gi4GwEAdKSKhMR/cIY3tuofqmgtFWfJfbT6ndZmndbRzyygHebBlmnsUFpLoh7TaXupdJbkKJeQ
1OPcFBLL98zP53AWYTMxZoeRgskxBQlBvOSGMagbtjbKKJ3GfjqenMYi336HtEw4b1CVIDNWRDU5
GGcdrDRltBKvRQFsVGloloCwGLZsu0DNF6ChuMdA3DFE0HTonUiYud7xXL4keg3dyw6ZwuMcM4EU
GStuVtuQLzhPlrPHwKVdPKFgKEa9P2cCLToKE7RNERvafawcsPRJ21jKUwTkge9DYhho0Tg8RK3N
Y39zyuTT0kBlF/xt2ZQCJ9GgM1ocLXPK8j81YHDBMnIo3Idol1M1yDbNFMxPknYlXCyzLBjDsEV6
8rfD5TGE6TWZKnj7xl4PGH85IhZlOkn/SAFQ4H4/KUuQoU+xMDBMoQr4S0lNDAm4NBioUu+bo++z
nMRzJ7ATyi/vx2U7VrkT0BON8jSZqToFtyPL8b8P9wwZmtZfGj3c4GdtbZLWVWAOrrbM1/dM/a1o
JypG6OVEel83e8z9RB++TulFRQ3KCAeW1/nGtwBGIgxVSmTTQCwpjaVH/D0QxaYajklisw4sHNoz
U4wLGQiRiCqexE3PJLDiW41LvPIIEa2Awqfp9vNqjdxstooaQcpKEvXh0wYJsLuYZNzps+Ysr8k4
MWpLzd7DGEqpMqtrLFUYZ8ek/9NLpRSjS+RG9yc5dpIcECVHRYMPG3QRYTzE3wHmiu1u512L2GSr
OWTz67RqlHQ44+kvR8EtKMkq6BRxhvmdPlBLoYDYZ5LJskL0kGZFs/L1I9ACd2x7vp6cbOPZcxyL
IxDC2VdvJmk+HlSqlOiNRxbftlIDA/a6OFxHX9fbPK3R4vURGJo4cIMfgN4AWAmL9owkdSGdmaEZ
JYV4wgPwq8NmzHRhicwjvSlKhGfivtoGRb3aY2j+kyiEYIJjnGP05+vn+M9pQ3zeZK0x7BmuPlAs
+Ga0GH6W2DSM9j0Qn4RrgzDN1MmXKxrRX9L2WVv6y33Vt+dKgGvoLzajTHm4zhaX41SW+mjUG22S
TMmA2mp538GMBmLU6MrfHEtteJQQ+hwe4h77TzQKM+wotT1Rg6v98844H+S/h1FKMIMykyG5X7+8
Y4J1cRzHh8Jdzj77lvMi+Wp/hJbqLRQ5qDLfK2j8/U09bbykuRE3xJyitG1RQmUt7MYM3L1CptEn
SHkoaxbXTqn+GpBYeHxIRImwROSTBpWekbaPj1nJScDNTm0UhT+DHfuJZXLr0WaR/yVTjYS9gVU0
WABDsMeRQ0QPKvLXV7/PUKlyAakTEBeOjbzSQNyb4E3X6k+2qJ/6GunaFy1rny2U9Df8oRCEPU6T
tpv76ehcPRhaRtCx/sMbjdZX+qmkSO6dJCV7YK5gzOsGXi9BoyiePERR3ujj87B9Zxk84vj2iRGY
RUmuwqMBJxVYFhCQbpt/8gV2lTAxPHk4f+nqUVCfW712dn0JLF1oFBbloy8WyL6aPuYj+6rEBQzS
bhYyORpeAah3pCZ3OC0kqUPJtK1qBne5ruAAZR2orVdkUE0qg58nO1e78e6fjdI9IEAQnh6IzLmt
g/A+qti65tM+u8S9bhA4zFNBt+FxEoMNxmc15neOPiNHSLQxTEqblI7zDEaop++O0ED9AhCz/XGK
Pb5hB4o5RucuGrW45ZCDtunNqAHFYIcvQ4P//P+1YSRVfCyzthRZwcvrI/EDU9b/f8U+ogY5Q64o
4YIvSuZ4ImQ1d/5DGWwGiEzpmsHakpREvUcjlu34KBJQ53WJWG/jHxCBqgiHYQ8CQWaWjPcf6CHi
FK3phS3YIZIsaiUIoJsnFChdvH5LLhAcyWk8G8fVBzAPJpAw5ZOfRHaqTZAaWHOUF78pMwPjpUH1
7lUSUOKZVeR4BZZdD5I3xrfXXanhvMFmPStE7dNeUfh9YDTW7ecb9ACFDPTVZVlfFSG0jt0J2gm4
0Eb+urOD3L1oETULV2+yGLP1GgVQrwIbDxjYG3swq19e3MPyrbVDcjmza/mLnFUFYOFG05SQzzzk
697dUQmBWRbW+J5YZqdLurx7iDXTKxdA4y+99DKe6JVcjeaBgDcI7TaSxAUu4MzmYTpqzo1/lXpV
V+tpSmF9oUWYe+Ruy8z+6P7dmI9/oLCuURcPA8KlExw1qnPq66G8+uqqk6EJ/hGP/WIbg+PZifso
t3Sj5Qv6LegE93VJX+utRLgIGZcpoz5QZalqD4eQoW11dIG14Ya2b94y6kuxtXBPeI5IbjXUS0XX
1yWGa0Po1vjyes/p2W6GcKZdda+19Nsn/UCR0H7V16ZK9OviDj2gZxyO0AzwMJHK836OurstT+iW
lGcRGB6VlT+KfrTzagaC/xkgtEVedT+ttW6HEvUamfzyUu7pHLajtdt8TOQkjadVj2CjtxTlsq5s
34aan2O5AP7G82msDC/jAoRfim5YwZCCzBkbhPaUQnv3Ce4ILrXvxZ/X7YQwiA0l5Ehrazs2Kii6
Txxb9JVfGox/wbyI6bzQVEx8QqK2Sv9TbW0lWZ48zXTabZZ5iIf5uGWFtSh4eGjvpTdtAHtdNPE0
A/yV7tVIhvXU6WEN4ucwaNyWUtETWYoMghanvbU7qd2mMIYRifLuTd5jFfXftHAhqxqLB7/+3JHC
DhgDmTKM+4IllA2UD1JvA3WTOCE5QfUsYXwVq7ycHdURMsgACP4auFNFWcaybgh+JqvdfJMsPtax
jSm4dxY/me4oXU1+8eWoAL4aq/Y43i4XKOrfKdryxfXGZvxE+pP+kYqsRKqPFqiOcE8Bzb8Tko/K
Hezf8rjDmFql971X/mT5o2V+D2WUHIM+1d/dBeWzEas9dV/TfkgqRxhJ4kqyvqdt9T7fALjLR5vO
EJrWySevFfv03BMKI0FGU8IlsCcMrJ57RaDtirLjkKQIoNCg4+aASAM0L6jESp1llmtSpwVYyxD2
uOt2ERD3NA76iyvJFNNdYjuE5CF9aMK/wsnlREKVObLTrQqPgX4aHoG/NDw/p9m/sGKSomXF55ws
dmSPEFefmBj3Q3hTP8D3zvAyGn/p0rVCdtDJ7om0jpsuRCIA141nsCT/6RejGle33VVRUpIi4bcX
STkobCYKSCsixpUfduR03XMiLtNZ5PvkaSlkgCMxiHZ59Q1EF4vg2YrfaaRiK44rchb7DBcAjNQp
UMIj6k/XjP0G5NsynhhOyrb6kj16toN4uKScFQr+2UaKrsX0DMkDNCxNJD0aStgu+8KpDiej3QbH
0cFOtSk3Uvw0hDHRMYH4qukFJSA9IxbYeEuXLVmei3l3YuzmQU7gB+lpz56/PK5yVYFPoA1VpI0Z
b14ZpYxX4wNuwsreItCQ+7R0J8wnFgMVt00VMxFNP73+qGCtbxRfxhuED/WPK9FGMID4ZaaAZVmi
ge1dSpKMTVl1hGWxmpIQ69r31EQZVcJiheTpLRJCq8CvlPYS4imfNi7u9CEUf/8E5JnYaUGGHJCw
j6zQSEiHHzj09KPTPAm528YaLFP7NyyUNCOvhzB1JftpxkMZUXRjkdtNI2Zi7wOzKGswbM2s86sG
IMjd/2yvjqOCvD0zacuaqJC9rX+hpGyUxMIeBa7CMK5oakK3T1N9Xh7TqMgJE1GT0U8A7a+M0yq7
hghdyL0pU8WS72WndvAqBkDs3kzlXTZVxoKtvHDcVo+/Th03KeT8wbUfmjCj3G7sFsDYzyWYW+QX
JmWtlT7xH+/MrKvliDuU+ZDpm5qgRIk1VvYMUGghXQFn2KU7EZ0dd3EIpdor4DtOJe86tDdthyMn
86zX+T70m/4ChsQ6BosgHStV/pChBKyhaKxlmWh6YSRTKc1x1dDuogVJxQHtYRTEGTaA5WSM07xJ
O2FQqJUcm+zr/21mTbkkZ1PaoS8kMqo5kYxOUI6WzFtoVIjU85CVVNjTwtjC+Zs3SAynb0gv4nMm
3CTqC5bo5boFQdvmucCa77JuR5doUQPqBiUu06c43XaVb3F/r0S/LB0Yy2rhW/dn1V7NERXbB3Bl
nuz3o2VKifnNZyaWPLd2slVQcpsIjEHo38TiSEqX0Fck3MGm49wrDGH8a4xyn5y5rkUbPOlBPser
XQcXcNu5WpQh6EY0NLUz2gjTeYLXq/uLGRkytgdL7wyGNw4E3rVbh5/HZBkTqFxoNZQp/a5IEMWt
fatyewFeqbrXMs3WPGtvJ/nlFdZACdNrPkJcq/H/HFv/ibqjnraEmAzl+UxQFlHeGIJudelogEJ1
DQCmAZ6waEjnx0DtN7uDCOnRfhzh5qR/HQ4+6cEMZ5Y3MFZ9uMPxfo9dMnXZ/gQCTF8be7jgbAfl
SM7tIj7n3WzBI6GHctaklBcEeiaGBvVhVWVQ8ZmxlD9PyXedQDR+NaEdlja6JWdCNJZVQJo+yGI1
R5++czPdNree+84gFYdxhZAMB9neVyok3CBCRliSgo+ZaYIwRAQ8Zg2fWOypO/MSQgus7TustwRS
gHe4bjCE9M2TsbYV4XqfzbQAHCzvQf+zgphBpTZu6cr2VgYYI6O5E66i568D7Z6/d/UuL8Pg76QO
qN/cy/yiiahJIOBEClwAlVcpRaT4LtXaUJgNhjsE6UnhZxVRm5F9BfgNzeJnZliG7YMBZjxBR3IN
9ZwaqBy/glz0zBkzK1PW3360HggCP74MadFbj5NsImdzCM/ekSwGFo5YyLeB4FvRToNb9f42KRGl
dI7OQA9GVlDllgmrFQ+NBiVlxnaxMrPqpEsFo40aBGAco71WLxAKEGwdhwiYrJSzfydlsgfmHTLd
n+RtxYO71olf7eS5l67acKDi6Ig1BqHdeYuFlwvj7WdFnqfYQlCdSozAATuBzdLsKW6NZOKdhQpN
PnNA6kOy9xLgXsvHChWYUNlfjmZSVKtg6CEP4cJInkxp3GMld1JTD0K0phoqxreURgGSijJnRCSi
BkWUXDpkZQs/7LyxL2+1JwJFmSO53qq4iqaUoB/n4XG/Gz25e700qPOSyY252neH4ABLiNjw5CjM
BAQ0LD5m8gAeGgMOwYjq4l6iF1JT6k8xJmWc0THfBEpRUKvn91LA8Fk1F+IehU/MYFy5AoM5tUvq
2EuInOzZg8gnmefHHbTmDZdT24bpxN/PxFDPR7luaRWaYCNjaOI9syUqbMFoEAFNwzWvWXIMTY7l
yAqOIC8gpSrmZ6BVeHOHTEvml5QM1kE5s0+izFRSYblroMCPtTq0ry+zq+Folsfbtsnl1FrdEKCR
ulkatclLl+qg6k8W3irMVQdDZpKf3hE8Fz3JkuADnFtf3CKTxedDQtW7Z5mx9TbZ4dEoyi+4vOVG
24rrHNbdwycXbASGoIbHgHDBTSPTgqkSQrTHfb57DO+4O6TpjDfke40Wi9W1kYCw1/lqnhEUukpu
2uPkD4v+IWlzO+Km1GYF9pMhdA4Mbs4m3tL3S3Af9AszuE5GsVfb9gP3eT5oCEcG1yklaH5xvk3/
mrUAOAlqBedtzNplKNcjCNI6MHveRSa6CbqcgemVhtmY1Hzb4nLXLUYgYV8wfnONVjuTX32ZYNIc
9ztiX0ApcLu9U4e8Hl6XZYiNW7IK46GtUTMVx+XE4sEb9cem967TqJ2mgqOzpwH7lUu/UvINVk6/
z0j6MaArY5wuP9m86Y5IOiKjR9csV9SkEOyaIQazR1GgSVLirYmzSD1R25d6mcCqTJxoAY4dYGiK
b8X1MJ6jOCrZWmajRWz/Ei37H641zIC/fUjr/xiOvrY77uEspN9GKjU0knJQYQWIJxKsihnsdvqY
QCOaTfhUNcAJMF3ldG6usx4oi36owOaPWtPNsGBVPBnhRJB1c3TVpGG0XiBmtCPR/ntXlDKUtu2t
BIlqGXf4obq/pDF4HEv4Ryks643intXuhlbcmc8f2ipVTgh5PrzwELXmbA0qza2/GXtkGR7MV7sB
uCjzGw6V5Pvh/wp0h7WcAtQCEGVOS6cbhIXOgZhXm/IZ6da5zIuo5KFjxM4KfA7ZaZDhbKV41jFc
jHNdRXdfGItBgBVx2nUUWHVNNaTxYR8eodCwVG7yl2kzxJ7cYr9I/UYy9tN85ZtSb6xNdyqF9pZP
Hi9o6dEq8FOqqHliH/aVtk0JgLUibiX2Y353encpGJNRH6beooiOCgMvAyVCEOGo9YyCJFWlGA+n
q17aytmb2hQPuvMOYATgNZ5YZVjCKO7A6RXVAJNqso+jC3Wx3lYKQhYX2yjtOssBj8014NZLTzRI
OAbIRGwp7qGoENNdmdpozxp65I1+Kegg1+SaYWIbvgSj2HyLRGXbDR6jqlEC2UdCBr5TsWo450OF
D+dwStyAasQoOIXB8bCykF7MgT+JAvoMfFPZn9UCbfypw0F/Xzg2L8Ktz8ZNUnpO6JtxLxI3P0EF
bPZ5EUqON66+j6tmKhi4ZC7nZKJgpch46hwqUw3MP6DYLbesZCdZ+aaUK1b1PN+xxfv9+QSNhoJR
w3f4AXdmSn/o0uir1JKt+xW9VjXNBYBWvJabfek3/7kRO7rQgC+3IBIEY4KRxqqae1w/4YGdWYXw
X2MstOouDGMnbFFsMTAd7Tb2XHnBWeTStPQ+XqBrb+jDNVsNgMs0VknbEqwsbRcWGyzmbD17PY1C
9p0kCV3Cd03+G0IiPKF/KnnPsOAJEbwHzCIbRucxO/931uGtwsE+rS6t5vwTdlgro8E1Bn9xDnXT
9X8NQUsLagpSHG5Ge4FPdl6Ne58ce9Qu1j5uuMw3epBYPe8wt3RnN+wyP/x+AAoQicW8NJlVHSap
Be2Bd/3ya9FL8fvmDSCmKUQJFFGyxxc7114pGQUWngGDoZZGzf/07SIZgIh7MgHyE+ft8I04XAj5
WxnIZofYCqUCOXw3OUlxezKoPM/brS0st7s0ehSVZxo2rwZh7hQX27phbWYpJzru4lvIBpnnSf0u
s3cREbKN1+khjh8yx0udlGQRuMsMrGOdOALT6f+kwDYUDOoQZfk0H1m92x4KWxe2Po7dRKr2xBEd
PXxKegD5rW3CoeFPZRnZASEnRwI21YUARQAsMX4rinMKSv2KFu+fgBUPxwAzmrG1NnNYj+vTjSBC
qvkCDeh6n4j8db0Yx+/sT2SCEBbsZJ5GMdahhJPmqDpVBdkZ8XBuQAXlz83x5vsHCLA6T/NiMhet
PP28rMTj7yd3yTdTMS8YzrL67XkKZuIiCrgcOJHc7PCBc3H2NmTNDFC4li7UqB00jcsA05YCvB0K
c/5DwmdqKfDozAEBRfnlOQ7Dt7AQVVx1gbs8lO6HfDIX6f5SXyS1PxweCn40+LiuXG3MM0DE9yZf
S62DxZ7F4v6ztRJLpdHtop4ADZyONlRZWiSX7nzM6/tw3Bryi4R8l5p4MfWEWxCrviOTSB95NiMT
Nifw37w1g4J/cFBWY+s4D9go6oSG6WFTf5wvSNmRK3TsDBfMLwGikhvo2eEn+JYzviP5oHnM5KBI
MICAhqLbv+vNk4v8qSHDv6CAXiXowr0UE0WPaqI/NGHVAE/rL5VtlZtAf3n3NHtMxKviEpzZHHuc
Nvr6INgfCCsBHJShdmpyOya3GoKQGi1fU7AhjqxZJkEtS3X1wzdspl/8oX/krAhG1MEASp/3Xeqw
igp0fcGzvB4gV//1OX2wBDNsZ/BwzahSH3eyaAR64wZvXUxw5wBtPNWLQvQXgMnbuxoVI8dcU0wL
v0ALlmKp/prkUXnu1VkKrT/YDlV3YQh1Q36eAX+RzArTR8kpOmkfg+7t0aCGUedv0U06nz5ns8cL
vaVQA0/y48T3mh6DqmmmupNs865LIDsZPERA3Tkl1tADFr4QnpaCGncS4nIZdTDVAqwwnYHMk5gK
QEyeN+D7YHph8OoXBWqQ61NQrQwyO6XL7HjYsp+1AvUQdlPq56SnEhLXpX4YjQFHU52IdK5D4UkW
SVo6z2XEdxVwSGU6V9ZTeO5X4VcK9ELpHFP+95vEDvQL5wCY+EERBzSwgOWMTNuEE8xA3TlJ6SDg
yICNFGonXyvnC8rVBQPm6DKSZL6LIWQLKqP9rwHul1tspLvK3/fuGSf7/SfabhCdep2jTPhsDgJq
JAtG+lSAmeYShMK4HnTmy9GURer/lhgHXLZNZmZVlYs4/AhKgMLrxbEM+2AIuA9sVRGztqiGf+hf
keXYsF8vyzV3Ax3eZIfYFWol6gHeQd/SmNfFNABfBuEO+KCkhw6D2DpsOWnJCklDp1sKxzP83bCX
TJZGqMzW1JsS9julm/d+bApl4qV/vahI9LUzyYrQ2WiCNzosaIbQhGLw2A48EDkQXChA601j+dTq
M3o5T+r9dHrrSbo+g3Wl7Ne/byhMLusnFfOrH/Nb84t78q/IlbAd73ZIVUMKRiI/9V+he+4MY/17
W95mrijoCxvoqRufbgA60ERsNHU8UAjpfKZq7h3gfQITNwuoCDPJc3abqLPrQ/vhuDaJw+8JrPWy
Y5sNYBQkY9nUGZfmRSdkZ8FuYJ83I1HUGqS6SHKXYwfywnVL4ZQ9NpK/VKgGzI4aEfB9swD5HzB4
w0OFTCUFIx01wG+oIryrnZcEFM/E+dsIMD6fApjpt1/JY+huLhHCoaITsLUPbdTKx2v7WgKpD/17
qLtKGS2w3SwpCnZlYq7tPfKwS5mNkAZNYtRz3NQ7g00jvPxKA0ipYzaQWgiC0WoanQDRb6+Ew6AD
cuBtzuyGbgfe3RIG4coVOXF/Fb7/z8kSeHt98hWJ4zhZRN7fKLiS05vN8Fh/63m5YLX9aWn+iRUi
bFcky5TBlZT/L5VizHgKrIhGU803y7Dxcpxzqg+8CNg2WkotpsTrq1AKJr/W/9MOncK85n7lhhPZ
scl/voNNoaKRrVJnd2mzgVPk+h9I6JrpTR5Yv+jq6/4BJDmqQoYPG+CPGs2tIq1pr+8vH4NiJwc5
EmkETWeYHAd6Fdhy8xv8GfM733dWf8jhIYhnNKH+najjrwFYqHhgE3f0VMzuEDMJCuydOrn5H73o
cZceqbSWm3QumHFXM0d+V5gJdUwNBQzvu++Ga13NlHTQxX4CF1XFCB+Z5UaUxY/hwETo1PjfQ80F
lsX9oWW7xf3NAL5kFusq7DRcv/pkaRHjmicdwe2PFml2lwLtt8hn5HSlUE9m5KoNAkXfZYdSB7yc
aEdJBl6vaEV702yhVZpNpXEaPxLqsFB05X6isEjmrzIyebRa7drIcVLAMH/svyMP9oehigiZ5HiN
6HVXwpR1mAOM1aygqBo6iyJ+rWcQiVc8aRKJ8+hCEHt9vJeRQsLzLp67aPJh4r8MwasWDp8pdfxZ
vtKBEU5Eu4iHqZa2JTHuTZbEMLzynRFoUbbnK/tSgv169szoIfiNNf3cNNy6Kcdkge6aYG3MCo0j
z0pHK8aGmrzMxrjfSQFP5QdI3S9ln/2AAp6aPQ5ft+Wj80h97uJF40ofOV9g9PEw1h2RNCmeS8uY
XFbRbrJi5d/eRlcZiZxsnsNAL+4yMYWYMyxa7iODz6AVVXt31w7jt/rVB9qyR+AzvqUmKVT5J/y4
h+Vfpta8RNka88BKisOWnxHaAgaECEVg3rDogXz+13oqG++7sX4fvGv9vkbFNsWGUNWMiOSrsvYf
gKSWaiScC0BaRcANOGoqcnjLXRLld9B3aFXe1aK1XahyCkruq3OZluhn/LbrV6qNXiUVrQ+GUSR1
+xJpZMAMUXxI+CRrwRZi35UxclqQ8Vm+ComUVW3rUdon4zNkiRjORCF073Cp0+m9YOnU4vlFeGfE
bp3eKPvqNtGNzuqw60BPplSQr2bFUQsEeivQJ7VJAoPzT2F51m5cNjcovoiNW1u5/K2XA2429U1X
pk+ApXCZ2DJ7N592AKRbbWoyzyVWCosUNnTi7f/2jmB95Xc2vER3e19JN08kNnb6ArjH1NIFWviP
2QlDXV4QWvnJUeLLY9i3QvIna2beeej0UNodwoFEOEoS3eZAab3Bk1DOK/+MioElkZZqekyIiYzp
2YQNFXIe9xXqsOWrFzW6G6WuTS6vPZrVbEZ6UdLZWsqX06NH9ByR2mhqkhNXUZE+PIGNio/6w1ru
FWPSdYVJ3qZNUmcRqG6qCbhoRMzSm74q0r+39BUSkh6O/PdlbAkE0q2XsR+nBel0/PwHRLOIpyM/
V5fIPxK3XkWplEB16Nhv+XhyQzfXBHg3dMWaG3zP4uEkD6V2V2Olpl8sosVhdv7tv9GA/fM7HIvk
yasNP61VHsiqCYOSc3NRRhbnGwMnbre2uVaKzhKbbXY2PjzIOYXMRZ8Z4ITfIsrQWqZ7yxwRuW+k
qDCbReUl659yf108w+fDOalFGeAZrFFCeHg0na+3z8vqo9X76Iaqveihz/Js/CN85HNxToGgCZzC
B8TF84zlkNbjeIooIg5Xhh9tjOQTe1YiM1vWbFwsJ7dcCaWm4TGNZrFDKAO0AlpnylZ8m1rJeGvj
uLaTHX+c+ZUF6amy0nGR4LI+Bpdcy6SwrseQcQLphiE0VNGCJi686Fa6KEnsQF1sG43Z7fm6p6pe
bHuSbbmBBcLs3L+X47YBsMAN8dKQThpmIx7qLGhB5zzzJL22exOq//Eh3qn7ZQ0hrKZY4kryR06R
dbrlS2afGfcnbegfTgYh6n9EVjnJcBFpTtnMFLWs+5eTuqvVrdKe7Q9JzHqJo0g7ng0goWE0VTi2
Hk5HCO5DIEJeTiUynUbnSC1jfWSl4AclR3wy2JJWm2jaQcMpSl+Au1v9CZeyb2x6LWQrayJhBJE7
Gr/AM/1Jg0hD/yn4wwP/DwBsn5eklFzhTcUQuyC2hQ2W7ROu3H5RILdeBlwX9J3zF5Es/RPDkLlJ
a7BhnBnHdCYTPahE4IZkXCNJQVDcjElezyCTKYyc/Xjp/FcP8dMnIC6OJrPDNCrn2q/m50/lJRd+
4lQBPJdFZF3Ut4bdqX4tiKUka1WGv4y4Ua+lZhXU2k6zAPoR//Bxl1h1N6Gdw4xSDi2QgQmPU/m0
UTLso1glf+Jp+Hd+Mq6bgfv05khUtXp7qfAUytNT74jfE9mdo5BoqvJr4LajCcHwtc+qhNNUMNqN
gQjd1BZqKLr9ZjWg9/2MNQkl0fpm5TSZW4Tj4H/IukM9KP/EO5CAnquCDX0f7ffDYRg/F9cJWgvM
2lI7T6DgUL3EpJic9pvObjmVapHC/utB7veNBzgn1qeBgaQzmB4S7RCsNSh4O24WEH0+eeB11y8o
eNsncqE3BYj81bsinGgnSo7/vlk4y48AkTu18Lb6M0PdUbxp/VpPK786fj8enly/zeqUZXHGqQnt
aEU0Ynsg8SoYAU/tkmfp2EGp84LnmaY2RmSerpSbdhon0vfwEIpVjjjgwaW889i0ncAEeO0Thtv1
HBkGs3Wf9ox83caJnY4ppa2U00Qk0U3sUIWiaU6y/XBl0kCboNFkVe/ksMecHfJcGHaUWGFaRTHS
b64FaYQtnhHB2YXpg5f96iV9mVCfJjToQ6pEZwHG5jr9FsBa2JvIHCxsfF471HjW2k33DpnGjAnE
y+PDZ+qvw342MmhiwTEwXWcli+uWivohAECCPxBM+QUZUWWd11Ok1Cc7NgWMkZVv3cATdp7igwrq
RnuxI4MGN2tCs0bklFq8CdWh72yiXnMIq67aBm081ln/+Gw2wfjkFux4xx5qEmnEAMlh2a5a6M0z
Oeh9mTqDDdWQc1OqIxysZdhKGUGSJ8Z+gh9lRoQknwaPwFxQhaiMJ2EZLY8wJVWfDjWGODMiXl1m
y64FkU6UXpCL90vYgnaxb3kBPM4t6VDh9oKi25u+iTKcP3tNA+NuMV2ZdW2aQHRRbsHpKtj98uiz
KOFZNHHhB4dXVlC/MYjB3guCPRK/PTqbW1krNUa8nh2ryuTz4wwj9XM+arqXHdFK00JmHH4XHWCU
OsFMaqe6+xKAmHF4SXT5Hu53PWE+PXDKZHmW3V2neCPvKURFH4sCffL1aFNVsWedAQ34hRXH7STN
zXFR3Q7yIV3kIeFaBEbc5ou7JQu1sHln9aGlA/ef4iZLzDQLR6+8dZY2/m+2hMm4CYwTIHJPQtUc
8nHtIeZD2p+VvljY8OlgXEMTpByZFEO5QK7luAPIurwJXoNfTTZbyHWanuskUS83axqTT5MfrQLf
W9FskKKtaZ1dPiMiIxt+JzzIPLmrDN2U5F2SvOKx6hhaa6FQdPHVbsqTY+/qCkEhatqfOoyCTk88
8I77nzouX7JVenVncCTr8IKgCX0HRWv+FzHqkgD2jViPCwZ8DZWenI5MCMsR5kAzc40peW7ONuWS
jkwuKPbdUJMlOMwl1+Qo8xfnQvhcV5rOmRRyoL3eGv2smCoGKuGdivC0yKou6MbOHzJ+QZKK2W0o
Ol1Yl/Ra3rZkcaNMkgdG2mWHdb6s1aPZBlCqLaUhch6BdGbItrUu3qjLUiXUHIcHPRf6T5pfbvpY
cVp67BH++echQSLVlEpgBzjFbDptsqKdN6Q66Ee+/2grCG2/pVaaXFEW16J8R9PrNBLR1vWhs4OE
BD+es9CEydjZFk7VmZ+pNzLW/4HklAj+566xma3eydy9wVmNzLoagacCFnMFL+ak/WYpzn3MKKyr
oO837sdr/AAc9xBxgUhHU3+h1hFsBHCayCgNxq58eiE/TQCGTc+SVytm96x6GwWRJCnSlqC1KS8Y
SmGp48NNCCT2p8E97fn8RrdlDSZlL/uE4lf/4op022VpFslNj1fOhPSdA5e+TmDfUKbGJ56pOcqr
67r6Z/rCH6SsdsvtPbtTlOJ7Q3r2r/v84n5OqSyyiRiwOc7JGQXdfFTWlwWP0a4mcbEJ6/hbPpO7
Frn8wOluq/5tZBhiVE2zpWkiajsI7l3tNupT/fE6HT5/gcDlw+vrH8NkjZjN0sWI2jKjw5Re33xW
MCVKeDLh6aSnHyRWzuOVF9H38dAF6oEooWop3iZz7iMIyLsoOMr57s0dN1p9op/mans4iaqpVEPm
Qxb2Yu3XHl0umhovHYPol3o+8hmbMcMeTxQvqIP14IVe1Xpj0bVRvAG/8baXy8epI0d1HNnEFRAy
ZRh3BTT8U/OAdGO2PwL8PUFJDLjETn1h6L48UOXMxyNnmi7ttoNttFhIYjgORsq+TDJAY2T+A9Jz
r6nm7q0MCBCo1SBNdET/14i0F9c8eB8dy7jps5mSv7X+RsLHwM9CicxFhnZGB6SStds6cK5Axisp
CPKfvf3zM11bzTFcyWMxHkWJVs5zjuM/Q83IWULSJLnfpogqbJGsBpFCedxMLm35usisMBJph8Fw
ERxIUjt/XMseke7xrhwN+mBIGueFJVO8zZo2w7G9EdlHwkBn9sZKgSJXhiAuxKnBmdKHyj1FT2yL
hbpV9nn+aKCcUH6QS3BDlHPSq2CAp/DOsUNPqbnUbZcKW2Z5jkuoK+5qxDQ9n8XDJZFrC/eszpC9
A1iBKTh1A4Qn0Eb9RD8Bk4kKV/s2meaNCcuktgJeq4v/zEAsMJaLUC/GlDrDjLeEsE0DZbHx7YZM
kqFQB31x7W6KuXZt+bry0a2WfdZqRgoYZi3sQ/CBwfglt8lU5U2mE7ypI/u9DMJbtkl8IE7HjnXk
JhdUtUIsRkjwbuFVk9wgy4EHirURRWKmVrqFclOapVrAW3TZ/s5R62ZpjMHRFzJ+hOn6/MWPcLD3
Icykosvw16kObwmNHbkbaLydl+LzxCr7UkA57xflLghfs/vW47zPEncNmc1SerQspOCkNepxAOeb
auMwXZILavaUJrRfdsNRxXKq/bScqxAENIx/ABpi/O7xolf8u5pf7G+VBzLTa/z7p8ofiVBTrwfJ
51umc3wBKP0GG+TdPVsjPNQQs6pxTp6xuwQw5BK6TWa09dbK6R+pGLujS+YL86l6mbQLAyEefI4r
4eTsi+EwLNCYg8+kIw/YYtQ0M+KBAeq1wR0BV2umiB+uLrz8h/97TGjUWlzWPMKilp8tAUAJrTIQ
GXynCkhgb5z0AgqZtcpDBIWgcyKYHRgg64A7S4yjTtAKiHj3wtztHhII+tj4Iwa+hjDMz3OGtMCQ
tGcoVi5sZ73EuP2YKyiWWIe6lT8ujtbQl9syOYvHufJxjUKvBMnq+T70ncUBKxIMNf5JyEJI9P1v
gUtpqR3gWCJYvmz2VNpsV5iW1uGoe69TFHIKzhkskHOdj3k2E9hMyHoRG4451oG21+1QFFQj6oPx
EecmlU0aP9UgbIL/gQ2hgog8pKS6wLwBRFvw/s7VcXb4dogmbMfJqbJmloQJXQAqFJ5q9C2AaJ0K
MMqvI3itJDMZO5qr6CFPvWIqtpPACUgOmZgEHcq9sPyhKdlBiMTFv81fRNX3SFYRus/1ZrWSpbp9
YtF6HTyr3kvjR0TaV0wsiX7we3NlG2pvOXSFePsZPGkDQ+4AnaGpG8YHFQzbXE9p4XHpbzUHR9wV
x/MHA6sYDigpQ1Xyg9+NU+xomFVdXl1nnvxEMqAMdPVsLt1bvjxLhdEL7FSXA2+eipwUP3zoDnlS
HTobe9aJ+NkxBy5tV061zjEsCRRB50XxAzTeinDQitXBb8VmxuS2qS5JbnrNxBwZRcT4ZPcVUXa+
y4S+71XRB3/uiRQWm7aRAtHlPnWbDkKQMQElqL937wIVJPhW1zL7vJkQsXzZgmHRNB42ZHnccdUz
edPN49k9pIoXp+wsYNlqe3WF/bLdFnD00OA2l91MzZAKFFoedNI2J0UkjxT+W7/ug26Gy0c/saW0
EeML8wT6moc0KavwlLBNFHGq0/QCuzHmHP7QDART+AROsVHc8Ve1g1dGfQ7FC26eLgelMFKfJ/Qm
bS8vJW1fvEgSI7QNfeCVu6PssMDGYAg1LNj9xcviCOkh4PXV+ysilgwUte+cteSxs2vJorobZiuG
tfi3iDcLDdkLiGZzL9fTMh7P6TBu7tfG6xw+cmfOKoulENKIbufhdh5mQuXcHyzsgw8PojL+UzFO
xVRIa/3wgtXLjWU3ujUUpv0hhjNADc9HL7GVEadKQ+E4swDCFcqw74UnPpZdy9LufsMTs5hCdBsf
ifSqVwrca42WEsHd204Q8cuqj//JddGUYLphz+vNFETUaOcnvLWCK9o1/DyuRuxUQ4iTnzrMDnmB
yFANtOK9hfq84Gg3Mb9MntEmiq0L28th4SXz2DDa5qhWgdCsACXvW8hYj+ce2lGxhvDIeS+6m9FH
8xQkW8d5x+/WWWmqpT51FCiemDh9zb+2UgZl619xihumWdDPSl2RQZFx8tfPSh3IsM15nUaLmZOT
+8KknfAz/t+ecisUJkGNC44MEWu3laAj2pQEEs/gihPRyRPfO/QSH597v8HB6JnFU8IEOHJYHwvC
wIEpRTWSQSkOGbNFUCySJhhKiSSCHQ2+ohPhKDsKQsVMC3uZsJOW3pMWESRO9MJnx2Pug/TSHVT7
gLmO7yKvEyc0iv0wc8XtKrU6A6NU4Hiie/oDPe6jIPst/GAU4Y1JS1rweOaJhduDfUNzVt3tVFne
roRQFoUnrvfrfYmXTBb44Y1Yokc21FYGhUnTk1vfTDtzRTTLcd1cjnoPrqsZjkqh9XOiV5nd0qj1
JPZM58pWYM41oDMxJ8AX/yULEmR50RWiQTukrnYb/uxkToEfC6iAMfRA9P18jmSmXw7t6oJ9b9B+
2LTULGO+/JqutIyhqZ6MA/I/jcs12dWnzTJ3cyNYdFsjFvk2aAHmRQppLTVa9Fj6v3QzoOlpojGc
WAR+HhQ9SRFU0MmByVbwd7Bwoq7nVIgYSNl4ICAioS95tARb8TITH03s1B+BNnoP4GWiJDFJAEjf
bz+S9yZS6QzM/LeExNZXh7Sch5lVqZvIQZZKSi6HMQeRVE3E6Hfb5QpAMCNIhtvf8iTaFvorMe6c
PO+JUdi0BAk3Niq+aGEOS/06v0DzVB3SHdNgGDGc+SGCpThCjqqB/Ifw533PZA63g3p+xKgnM4Qk
pjL1DVR3XdUdQI6ymKqI/dTUv57xvogdL+KLIrHQj3CJ9iDX3NH12vRdQUDCCR1pZf3ywatjgoAa
BB/zB3yx8Toem6335A2wHEzbcdUzC231kmJx+AkkL49QOTisu5dW5/bWWt5O5rSfHF/goD+UhbbG
83XmeOGRaN5EbKJJnEmuqV/o9Ve2OhAOU18NB2dd8y1EVPp1whg8eHvUxxI5XyIq020+nlr/Wb3c
q7FxXsmDk2GgMxEtT+M4wRirtQ2omT2CB569pwIk8r4aFxmHdCnp2dCJQDKgGu21+T38YaZYMXau
98aPYVYairRAm+3MI34I8s3du1QIwjzSjQjcFaEzEvnO83w8tT16NzL7KnOI0ADLep4mrnC4glnb
VH++9BWGiQ5T5ecxd1mWAdvsqR410hNdFAlsAJbazK6yZr0Mep8cLTai9eqaV3JcGM6+SmFK/VFL
Oxm8aVtsmdM343/U9W8il00nuD09Cs0ciaA56KrRDplQ7SyUm1MFb+xBWtui+LyBfR511+/3QXuz
KNWrGqOTnodfvHG2wzN5mAW/wX7xmQKRY5vFKTnk/dUK9oX4SA+tOUx4Ga23nFczMyYc55fJ6267
WkzZbttsLttCDWojW+jFxw1ORQq+dF6BVp3qU+jvCh5SVQceqRTadD4SYVKUuZNHWaLyvxj42hzZ
Dkz2gLsXtEBxCPZVTqhhWIXP2jblNMkFhegYi3Tl6M0PWHPWzjss06lv1QpYwKfRf959CFtqshrO
DhjnMUcwCkjJgeSexXt3KIW3onFpM0PyEy4vYYLew0YF6l1p/9ZrKsGOu4TDijlQ6F4qemsGm2iJ
qw+FsbG/v2nMw7NmJp/Zi37ax13XJ5HfBLCS5IFowiv2jWNxhBozK03v41BLqe+wDfsUyIlhzFom
5z96ZdM1xZiYla5m2GABGDFjvXlOARhHEOS1s7Pb3GkDZsSqYOljGYzqZc2pgLsY4sDhRhHFqy+h
t3GB6V2ZW68t2DvlsYH5uH+HKxf7FZQFjQGSj7gHsyXgjwIy/ui3rm2Kk5uwNp3MaxC4EfjR/l5/
SKUVUrkD+aqPXZQKInmDebgL4YmA5Hxf89f/l/dfLykVmvxn3fBp7HO/nQN+7UcYmSg/93CuPN2R
F3V7R0IyyGCTV7rIWJWUjkkrW8EmgMfxVoIVnVo3kheDvo0+GdKpf9aB4i+REQ3s8BAmnjh3WnSn
JTGiIc9H5DbBOHJO6mXw5MUaj93WJFLTWcWdSwHxwgbu641kKPgvuVsoxPvb2mJ2vjuRxYn+l0te
Jm0TXHZ4kcGGKBNS1tSccSFcXPvFfeycSUqFXo8eNJxL9QowbR+WP26Xodyi1D1dX0plWiqBjchn
1mWRTIdj79V/k+3vXLpy3h78AAKfiUcNXPGWwYFRxcoovE68UzgxQdxojdvAJilgfyi+v0oL+s1z
TTMl1xBW1xwmO4i55iqCyYSuGYxkyIrBzSUoDYm7QD4H9AeGf4fK2MI9gxJ4Ip3n0ngJWEjqpY8Z
T0kD+GaJhj7YLRwPoalHjREPI1YY2qQQf+RTrB/VJ22//WwvtK0/b7IYfzhOhdkoEfEaUs9dwxHw
o0kfZ0oGRdBxuoLgBESU1MMG2LHEg9LHqFnM1+g4RQCbFeL1CCBQ8PvcNswAq6itUNoMuRY35CrI
nfuEH87gGEWAVKD7J0YgDI7ALW8X7tG0MBRKtqRt8HGQrjXH79k+V+JLvyKAjR11xTaVwWzhii0+
WwAa9JwmX+LrCaPS8fbNDyDrD02k1DIztIAVxkta7GTNUYBR+UAjjLsx//FbJ4LOi9w2LbRX6BWS
tq2hilN073hO0AsW+VDup+y/6izV/joN88jkpiPdtgHkx967KuK9xJ///oT5THfLGcympujaCiXW
aNPkrbWGIABprfL6h6jkbHRnSonSCNxG5Athb9wtuRkIRbmqf4xLXu4z2rmH3+1yTCqwN1y6dJW3
QxuFo5Glh3F26C0S98pPxRui4nWzM++upEjH58GGZKblGvW4Z5YQbfd2hD2uI3lSymhNwbcKAAd+
6QL9kKC1rAaZlfYiN6vzCaXjJTXhHLL9gntGhIIj4k61Z+YLVBh4objNoImCdlYIJQpnnEboh+ly
DX4Qlds1uS0Q/7FAh3tUkpN2n1ZuOQDEdsBKqiN30yI9vmdx06yv0DsUIZ4mIo7W/yqYIYAFCUyz
yaItLLdGdt8a5E8HLNOe4ZqKsCKWOv4a/6bZbSBqJHfOxAozcL8Ba43fGt5OHaD6q5a+3J6odTHe
PdvpmPkyXtw5COOCUkSK3oXElt8Bc5ULs1sZdsuyBWwA/x3cmSkZ8ZByzQuGj5ATZ84ewOyfsijH
/lxh1psVS99FGOiA7fIP2B7Ew6nt7NNbSXysFrEx9cU1yTTglQnnrsNAauf1IZha2iXJl9WEJxGC
mKxWjB6lK90o0QmwlVW1WgjVRF3aMJEah0noTEWHoOHP/GwGifZBuPlLQRDA7fq4pxq3IYC2rPNB
CwyHMNJWiJaeMY2L0Nu9ugR1m06YGLz9c1Odo8HAgHsoK5NKcVkijaUiN1zhrmeiC8L+ed1mC2DJ
J0fGMVEgwOfkx7myD9V02H1t1PRXZ3IE2jIBo9CeJfBYBpQL7SwEsk7eps72RWgpvwcbHXpjToWb
tXB4yW+FaxAMkFsG3efc7p2YlHAX5ZpzlFCCY15I4OMML0YEwKNe+w9AyBY5gqLCjri7NOECiuUH
oqiMbJUKYb81M4lOYdJnSh4CAoylgCJA5PzliW+JPdFpV2OAp+wkdCTXLLQX0OCO1beG7pMRgQFj
T4AUdPpsBM6YYl1XaxW37hwT0cl/4xuAV4fZYBamGVSiFAajuvWO+X0gq91rG1jvFOUxpr52vJvg
YzPUIoOeuZGbLXfm8Y3sm2hdow5pWOrAc5fEbUGNupQGbQbgoDltNQFxEDCnDZeGz1MS5ljw8P3a
dm3PVBuflCmJLOu6SpvUX4wPL+Eb3/705fhBScwmiKLkgNFXiJOKYj2ySe1odjGDQWses8keKkUe
jmB5pVEGNsdnvMikTqUPxQRGSsFWB8l/FLEEXUnvq5RI/liIwc98YYjo0I9gP9gFVhKlGXcTJwie
yTl0mr+4KVUSiGiDI3z7rgJZt2Sbpno4BmtTNangNTm9Z9GLlw6oBp582Y6kZFuuRubLtYwRnRA2
fEE+0A1zhel/cba3TPBL8r00utYzSc3GPyVWNJowBiOOSTVSrC/4uYZqVTYinRZB2AFrvYLq6m/1
+iuBmT8s7hwvRgT8i9GxN4yHemEQZKPGbYZy69hmONssi5koR8PbjKdl2t34awiotz4imdQlRSFX
zb1qVyyeMxp309Jjw9z00flEIj73k80SeqPaLTQrP/Jw7MKxXImYhTMPP6CO3FxIfXQpCaxPfAgq
6NJZAmS+8Iknrbx+70a7FVWwXRwr9AdDVDi1Ij3AkOhJ6qFWFCvoEA27c8bZ+tjfSHWiJXGJhyGu
+vK+NPvupos8ju68LvZZH0sZ2qhaltOHkEgCNxeZ1rCPFlftn/e25gsSjcyB1KfodB/qFGKlUinA
B2dMFrvHrSlaFxjAUoL37im6E0aUBHxQWKKHz9y8j9wxq3084wKobr0aVNRnc8N4iU1c2PIOpNHk
Dv1xOAqyrtqEAHeGAqhbNWJdoicZxrV9sMAAsWVorgPopmekCfH8RMabdbFrT+f6kCjzP9wnR4sk
IH/hZ7tQZgdLCivY9YhgA11XoLOJp78K8DHKGqsC1OFDBbBCi3D2RVvYvDWKk8aDlg7GDIkpe3Xl
JkVjUDN4CYf+1OmQ7WTLwc5y+F43a4/KRMQY9jRUDXq8u7MPE6eP513RF9lfUtHylDNzr6BdfoYy
j2C8r4othJsf+ofo7KpDN7SWcvjmvn0MOs+Vg/X0yY2EIc1Tq0G6w1tJvMrpN8bsW0lQcVPFnp9B
UbVKV7TNh2pIVEFrPParGeMw2rVRwbTHiTnSjnt3zIhFGH/xvAhp9DrKd1kijv4CqrfAiHu21dTK
ypbqr9WBAH5oczNxNedEN4vh8L7aJk3m3aaof8AVnckEreQN1HQ983RAUtFuYIvDbBp8gKuevAlK
yCF5W+xO0dMSniUN5oxypz3QtdqxhkqyaaNdW1EnKpvOxLI949lPqBnmSWioO+p1+M8GZhSBO2dP
pdkVSnQtKpVFenHw9almFr+o+fQ0nqoHva0k1UZAEU/8OrVG8rM8shpQanXykt9KLr1D3Gitqx3R
AkxkHefeNnB0P4iQ9i1x3P7FDNFy9hNS3Y8DUg2DXb456Ami9xDCc23fTotjnUOSPQBZmRPvlVq5
nKsO7YbMIQLGby8FTyi5l8OzKU1ghPHwP4Q1QIXUF9gd9Be1jR90iJFhpaHLp+FmPfgtkBDfXN+g
TWBwgP2lN0ZJ3eKFQQGCMuDBV/xgmu0G1Or6EHukSJ6dA1mjjI6iz3hepVTAiSnrDywu9SAke+17
uRiq7YT9Wpd2Ws4mDcuC43w7b6BLYCs/BvWknx05L4rFwf8WCT+XlN/0WAotlnbYHDGjJaDeRspN
t6SDOPXFjcOYxexdb+ayOA2nBAcw9ltNCFMt18SCGvd+NT9DmfQqWiYEItcrOSmEFy4NO3cFU2SC
AG1O++dS1Kl3c94GGjRdjBPZtazbzHrVSImaYfslU5EBkMr9IFFEr8CKedGflEfzN5x40bN5/m8u
CiVm8FO2rBLIOJL/x5nU4TFf4BCAfLOmevq+bHEsRQIKA3Rcx35enhsxX1ehssioAnK9xkH6mNtP
6LZSzG1eCh2rn2unj5PuVVd2ribSHpR7YSbQTe91T0/2qYwTbLiuWOafDFqtLCkZOOOxktytXCRg
VCIn1xOI9/FKIDiuWiJ80Msfcz1QpvtmwQGeaWue2LhmDpjkzNRpzT5v8vMUXRzVzICQwhYY0uSN
MkFK1bgC+vdCRFIlKDqXnhgPB+OqMlLRne3n2DfvYdLfq7R5tkYdPzdltgSNt7Ds0At//xAJW+32
XNMSRhqinJwLP0EwOGOQ6dvWMrY+43H+xa7H/GTWUeygjeXTS4Rf2BE8Bvds8Uo1IcIETvuYsizn
oET7/1s91XeHwSkzRg3jhtV5noDeBw5MbDgKM5t+FDCV6Zw911NpPBkUX0Qkm8Y28LYweQkVBzEz
PEGSFNqpifCInBLBdEcAzzAb8GaFIr2BUK3kWcI5FInQ5lkn8zB7hM/G/LcZxPXsrMrhXEmmDAJg
2MvawlKZTofC+HHrP+TpbF/e+Tz+udK3g6lit1H5+A3tOwO3iCSJZ94YTaIooxftygqtYHz/+Cka
CcHCMxycJB2jhyXqMOhZ+mWAHrYPKXiiViBYRcAzOK4caP9EXNQt9ZztYKD17rOLxV3kCyk4T5Yh
mwJUGPgwgl21equoVI4gUt+8w9lyiOUcvJdtIIDMMffNMoPWiujXrRgEiKGd6N5t90y4mn0gpvJJ
sVOdf1ias7D6L5K9+GbUFyrqWlQd0zyas1G7vJ/vfNOqxJLp58LaRS9XeuE5OtV3pxJEB1g/PhfB
XBWZ09/XUciLA7/p2TGBUrlrGwoIMgM28OHIiDOIvI4B/g2VMeoFwVNTtvHqpZHj3+MPR1hzQOm8
OqMB3Zn2wVJob+WQpzX25cUcS8A/s88REJ3VuwVNaSGYDEoSLC4bV/gS7vYYBSHPsJZ/uxaP03eX
FWKNIASLc8FuW0cxafC2yuXuMMv861nV1K1AZLhurxlPMMSqSkKWwHgNW6KNbA0WObz1exUYbd5y
cZ+hkcxzb6z1UV+KT8TvLu3ypCc5XYkxEX7zIrpY7DIJPG79WkOt0/H5HvEkDwrdFF3yVE5c+DFw
/iVJ30vHDk3z454I0PCkmLU/deWF25oVHjdIrtiyF2IZ8MidW9NCz2c5QOFAkcbAziwH8z4PgaBE
KnQUjVbEW+e4JgW89cJO6+s3SdAgIN1o0QLygFAKRJiFLZsOpJh7XRTbm3flviryBWKb9kaoQM4O
P5hx0XcLopSFyEAKgddvp2IF1wTL6veEpuYrgqmC/4p5QHLixLmNDS/GGdnXLq3HD+r7zfbU1bU5
idtwFImwMsGIyyf7Xrj8xnQZeS0MQP9w9NW3W9I0BauRT2oT1lh0kcD6xQXTrP2x+GiMQi4crKyh
fbsPSXnasgNcSVkmutpGc3zWqpcZB48v3QX+YVlgFdTszciYzYWQt61wJnPnSO/XMZ1kch4ZA+AH
rTpMUrR0NsOPlVVMWDawXIi4evSQc42JcLWyFynhczC6FO6yOMfwqH9WA5c0JnA8LDDb0Wbs6Pm+
fp/1nTDlUq0JHenVmFC3EhuCJertCB7Wav3576KwRXQUtsYgeOkPwLxPWAcYaupoPoH2+h6GR3JK
lcaTW1pDzm3tlA+T3mXZNymlvDW48mnfKbPWvvxG6grl1PAusZjlIpzaOkMPyhPNSnG+mJboo/0x
eNCpseNfx65DEJt/pPbYjrFxDi4j6gJOP5xg5SVaOr+o7ug+9/0gQpM/L9+HKgYz0PfHB+500MJa
s9rD1QPn7LVMvvwcfbdq6J/oBQ506SPv4UbPE8og9inh/3liRG+e+rQQzmYoDs5UiX23yflgkRxK
wXm2vdXJPEUyr31y5/p2+Gcmpcfe9S77NAN9cjNftDA1NLv75KKzGx4bgfqQAdrG2ZMViF9Ht9qK
W3WS2sp1gYKLMaKuOhWud5wWCqULsSeL6iccJDKyjU8FiD6Nemv590Zem8XuPjJIWOs8WllxNV3F
NMn83GCztKngAAJYVVoMlcBIZ7CVUuC65Q2flRqT26zfWCa+IPYLSIaYS9ocxrH6UzsDK1XtNJbI
BcCh5Bc9I4U9BGeMS7eaUFqZWkzAx3aZqCP0fBEINnnB+7CPK+Y2attiU+Siu3AtelAuOfV2AG1J
6GYAfIIjPigfiBJnXMzeXgo47NAP+u+j24eVRuDVk/fzJvnaH52XZ6/5107vgsq4rDhBZp86hO61
Og6ck2PcDwVqY1c8pqlNspnIBR2NzIt0zSSFB3HLcbwBUPAGc47h+0l5dD1/SWINbNq2RWoEWAWH
IxPNeLBwdqAdTT3qzyLSzVFyhFW31bXtX9fKbZuPE7Wy9yqHcPoD6ZvMT6OYu6GGoTMuQMkdlwT8
l/hShYJbhzUgwGmuBMMKL1ySPSA7BWBRYS4DDQ5KHKOWds7pz+l2l5C9PIGPlvkFdXJF1isbBab3
jw6As3GBIX6gDOGSXdo3HdLG1MoXTs8i44KCijaOMZji4gf/zcC7i5FPlEJTGVNlVmy6eDeutaAz
L2uhEUdNyGA/MuUZwUc2mrIbF66isDUjXUxgv1q5xzq7mNk63resMPBVHViPpxunWyHZDvg8+2mp
XWo0HtcNOXWtZkqMUSft7NkiftzbDgh++ibWP6xaISZPr8N371KEJ6QZJYe1OZdGGaAW2tEbq7tn
SWcTYCjutnlcB9Ns1uHpfNrX1bSrS7v4113nBChYqsoZBxug8Kg3AjWTmAiu+f62tD0EmnQfv7sI
hAl5Ub5vDDD2DXnlg1bJQTNdkUeFJY63+SwkMhK6kl5A5oPxtTH60qoF2tTVNHlESXGb7GAwxLPl
Q2QB/8OkstjECY2t4CoF42rYuvIWEOszPy3mlY8UkX5KXjL7pd4sItUhFT9MFBc8tH2wu1U1DsRk
Lj8AoG8uPTtYCEZYSTVpypkkmD0DJ+XWU1+SNMMOTSVbXwMjVM4xTOVsRGc9RzYi3gz5drC5xVoe
D2kXhLL/UKPG4jErInvhhbtG3Cyai3koNtwuzNrAqyPDOZFxiSsAsRzkntcHVfuxTdX9JnhKDukb
FQ0VxxXKpPvA8jY7ko3Jw5ZhubiJeY5qp+BCG2aF03XyvgwdMKw/TdNX2LmPbGQF880/JoKh9+MO
B9VLbwyYhFeAFX8/aYHCurTlByry9s9Hafkzryti8hJbxmE33GdAqcyZ10rM48K/i9p7Vs9nOmZ+
Z76cMiUcPTCrm5idHzOLerteP0Im+Ad+CL3ku3cHReWrpyYAmmHU5ne38IZNC+rO9wwQJ3Fxd584
NMD4c+qHB8x+l2C+tEb6XCvXffbHYucV7kNR92Pvsd52rB24AoxzEgOJPzT0qzWB+gOw9s4qU7Yl
lBUHIyy7Na1SFGlIu4u9TiCK3nsS6/2xlCBVms6UoS0JKDf4LEgjhhXeC0NzK7o3+RYcxfiCl9UP
TXwO3NLhWr0LuXZlQI2S2t0uxAIoqfbYlZzKmLk3aysJsVIS/dBxXj2Tl/ymMJNDgJ/GJIsMOy5Y
MhEKwPWv3QoAWblpb1ziZgbyKpol2sES+iWzIf2IJvkn/cV2QGZ2Oq3BdZsaEAzdkcpfA1WoG/15
YnaYQzKOgh6aHqDRcbu5Fxuzxdwt9ulcU4cqNVW8cb7YWR4bEEVluszn/PJf1dUxiv60odAJN2Au
fkoKWlvAvRs+AWQ1WbuKDT0sHLQCKWhNjmB0G1fBN63spQWO3JpPWNrTjErZYrKqdQ1C2/9XAqOt
IqQ7FTl+Fu5VNYzrcZ545SOc/0oRREaM/4s0caY4fvU2ycgxh2EjjPdvdwetu1lo8do+QlyR9fTS
E8GwuEJcojQc0jwfYanBP7ek/k3DtSTphCoiJTNcHSFgSjf5FgoGd4hzVq+w+3ECIbBU3ecO1G5m
w6HERER4DCSy/5b4xdAaUATTcoNx8eVmNWD/sQ4HJk05WGYAp9zXMxnwhTXuCRc1BSHvfyt+PsWu
kBQMb2d5C7WsM9Wjs6b6KrnC0eC+E70AKIctxrG8/OUXuQC9A8l5z21RpgxRza6fmMp3XgUVt8Yr
6E03PXhwhbzRwjUc/AUhf6hG9neLpQ2YWxFHPIjNOFNSA9GLoeUG1BktmrSgENWOPjwBWvnazKoW
kn8j9o2jOaA6DTtuEoxbBXCqbCt2zv/Q2LpbwcC+E9q5DNfQk36+HZvYSuBxunUpo8/TyTEo5/4V
F1sc8R/6EXPE6Sa/daUh8BofrdJyY5bfv/YFI/spZlnmupQ00SUZNndSxMrZk0EmBdEtY1Y6Wxgf
GQ6Rv8XcOcvhERsQ5cbIQQu/V0/XwHC6+4Y2ZTRA1jTpwQzmPkfI0qtrpm8xIzZiTH+JUQDWaoei
SZgucbGifMx7Z0W7/V9nyC2i7uEe30mx1zHtesFknjhhXtGBjSXMvpQgCR401I5h62rp3Z2keaoN
L8vBMIJepHn1WMXd4Oy6/6npwK8j0hV7h7/awunutj9El58Yi58TiwtzOjHPFt+mtGh91HRZGr6B
UWdvleQmPr8EybIb6SimX51bn0asosJtNcBVvocTKSKsUWSQ6A/M4uSG8wPZe9ZlulZXPg3lQEzW
JkOp8BxWZgn1myUmFxQ3hEOrP2qDyFMF+di7g42davFl/mRNmEtKxVVKy8nYS4odWtiUoVj9lTd6
5UnsNwP+5pPhHBIlW/89g0CvyJrBlWmO62dHMeJ1N8Ggg4+eJntibPMr+8NxEj+M2jcOnTKDR721
iPLFKQzT/ZRWl1XtZ4iWUoJu50GPVb9tCbdI2S0PCSsZCCPDdYX5tMdathHdLcSNjMNnBTgCgO8l
y7SoE3GCysUv4lAAD8nsuXA59Pdnh4NlM7zymk00mUJj/4ncMFmEO7q8zrVdF8YOBQAN51lPSQ24
tUNF26kFWbFtsJi9HmYVrQZDheH91GCdcosCeC5G0LqHAEKExWbOHDoz7onUBpBZ0tX1boQh2VWo
xV/H0Pr6fTvnV3qASNWgfRk6a5Yo4K24RjRcgA/b5pbsx+sdHuaTOHFTnAIARHE/3jD0v+KUVedE
xRMtj3XnkakIYO5+9DJwPI6MPQRtbhCBVJGuRmT5JC82jZeRdNTjBOEkHBh2DNRCt+O0UC32k5r6
WTHd9BdggQ4id6HvoFKA3KyFAEmubvPKJHZdrAqDTV2Qr6bEJPL68bGyMC1W2sRjZc6tgzTGfd4d
r7jTfjLfvZfFmheXdNcEjD0YzsZqljB2yzRR+5mDFuYy6xfvzqXu8AVuKZpeAHCBPOUdWW5JPPyG
5lhj0OE+I47olsO6wXOQdtj2lISDzVpwgdGvP+YXVFXBtRoo6mj1ZavFXn2wvAr/ZoVfy7s0NwZb
8sleaPrPUpyCE+7DuKsG3aZAOLBrooo7lBspdtB9O0mWctF2T3QlrPvs0Y2rtfjlEhTdgLXN9W7I
J1Yoe6vDpTOgNxDni01BefDBfMqdjmWLI4JTRJZaQqpfdUeFE7N8EFy2krFb6cVMPiIFq+1bnJ7w
GT3RcF4XnDa7kTCLS8/V+L4yW6dHiz7BG6zjVDj84owpI5Xxj+xa0IO5BXmLliJt8T6iKj8aHCUS
g0DBqtKnt4jG9rFrOfcZRkmUVIdkWoI48gNqx2DFMc/fz9kB9CD9Y8DANYgFmP9y9pTkBLo3AvaG
NWusQghKbGuaYO5W3Q+K7Hp+SBqSoZH6sbVGY95GPcvM6Hy1TTJuLi6IadrO5jQo9CgstCnpY+Ll
PvhPS5XaFljaVfU5ea5XAvv0aByBy3PssHz/NpclyBzLv8uPicbhELnmLN2c8QKyxDZi1aId8l7T
laJsqUU2vI91jIccv69DhOgq8pa5Lb5gIv8z1BPU2/oeMR71XDYybgSY4nV+1XLNgurFLcfYfpw3
rVTdNTjGjC/KP0UH+QBNTsXoTn5E9QFX9W2DI1u6kgSA4QfsmIPQV+ztnnHlnKLZq629rsvuKrv8
x9iErySrpOW8kIn0a/498ZEVd21ckftDGSouuyzz98T09W6+FuqBxsSFN0DbuJLeg2itVbc6wwE2
k4Qbnkf6epEzHIpM3x3ABvPt8JFa6Rvk0gudxAMdPhcLtJdt9dj7CkTxBfi1BPTuCikOhftIgS1c
zqT3PBWiLsO61ySnxnLIcKinirXebnVqR6SXEXAGFuakS+AnmOyjKTCAsKyf0aelVTwJ3C+bpXus
yLFW6ZQqkZ3phebUNuqviytr1HkeINyb/vFVCyRzClTwQ0XZKds2hQiOGJhOAZhqkgivwyutxgRx
RmCe4+dMqx8mN8DUCUVy3yTC/RJ8xRMSgdz0Bg967R0R4eKP6hrOKMCms/BpayMn+CZE2K39zAlf
wl/68mj/hnITCoabsf0ZkGZtk5bh/lrYdEVK1jBCuPk9gqwZ0fRbtL/+yB55QlQ5VdV5O3NQksvT
9IKHZ7tPPRukXbLxhFHsacJV1AHSXczLn1ZLH8Awgv1L/B8zWpqEAAQhxJvCgtabYnfjJSZAKXpz
gBmHnMUALlefPM7Qs95ahniwkoBNWpHWmwYOJNxJbWzoVMbbHLalVew1JqqW5/2a5HuSdiKoMAhR
Mm9u1IfcYuEaT07+OhF0jX9S3uXTUT9dqOXIR5/ub7RRCf+4GVr9LrC4/97/ofQpuWLWcgPtTOLJ
2cwESnEdb2ynio/zgEnvvgQr3pnJbAY8nHdnhq/xVhM9vbV9yEwyOsb477UaTLXc98TeXRJCC5q2
qQ9yVdRJTW+Cbz7vFKR8GJn/D+3aO9z2zp9+fKxcAQ/wscHQEdQj0WO+buW2oh0ZVHqrP+oOQqGQ
cjGeUAmgmxx4Fif3a9kUIZWDiTmM5RJTVKuducPVJEqWRSkrP+E0w1PVMD0AwX16kM4A7c94RkOy
AQHJw76DIVdxWxPfxvpnaxGe1wOD6agWedpQa+aJhSUrDCZvQcUfkcpSgr0e+CmToA2RR0b1vYY+
BkF1CFnggvKo8GcmNepuKkHS/o3NGNbXE/SmiHq68MI2q9kIHlS4O1FifpIujfOvETo+3ag8h8qC
LM2KwG7p91To8aepVBMX7ls+TrgAnjGivJNZe41+giC9ooKTUOPcz8Ab8w3K2nC/fOr8/z7ZROSn
033Vuou+wa/ir+V3dw4K2RusMysR96XNthbBCseZJVxgkc9JPsob2eUtKegxrvIE0DLk0LjObUJT
gOLl14Pnd8QwkNhGjZ0KzALP7OoBA+pFNV0P2QdoqkIVTCkaeQGZar5zh443a2mYZ2Q6SXKSmJ79
cjg8ne1sa4tsLoD7LQ74n2Emz5Ch9xI2kJxnfnvfADQAA0W+b1xpfyYLVaRQ8BhRe4J42Eh+QTRX
6kj2qjnridPXm8hFYhOI9n4LjSjakxBqD8Nb/vQ5QaZtcl1/jPXupHCCBgbwAV/wf6PyNZoEVuP7
rlTYi5/ldFYMPXsv4wCCRiC+kTGx9biW+MjaR+MFpHzdW1J/mfClMFdJ7bobdJfYHmKTQ/7lrBTr
e7wK8fc+p6CSzyZS+9MTrSThEXq1+WZZb4DzudLodqbJ/dzSXiOfRasvYy1XC1xb3n5ytVZ8AVM9
AJ1Ao73VfATKVflCu3/xk7APVnYtwycW4Z4tUzciA/R7QeqCRp9bAhTQvrfk0neVpsJJlVbvLpA4
Nm4LIsc/SdqiKHGwrRrV9uzZB2j0JjTRulDnnzNZFMgmnjUiZTDo9d75ipPNw+LREIGRwslmRXAV
gSulOEah7D0roV4TcygDX2HB9BdIDkGwd9ZuUBNkDcH9cx/BN03c1PpQ09KCPgl4SgB4Tcgudhng
BW8KM3XzrKrLWYzhQPY6zsuJCURmTZ4hZ2DoUi/lcZsSTmB33cxF8yjoT7QYPyRQtJSUjwYmxEJo
ENwqJd+NPugaqngnvXg5v9JC7dpkGne83I47TmYzZfN4GgwO+rh0oX7YM6yqmjc8Hnu8bJSMfn8a
KLODPb0l8o/QOw51cTPCROlCn64NDE2+85MuJASGhugCgzhthvfPmHanzCO0RKKVFGAbZ+guxpdp
Ji216TkACkDFvxeZJe1o80sHGxxpexow/9Ps/zQGKWS2pU5/33v3tYRHEIOrr7t7009bWD2ry+BE
a9Hwz/a2QPBXRnMkhNt2od3pg36QJh7s/q+hIyAsRaz9ztorv9XtI8NNFf89qQqIUVop0gNOQPRx
U3zbBoUlomGQsDqgpfg98MoxEnvc8OSFrOqReTCCzaG+6pYRPCI8KUvY31UfQkLt8+tRwLhoDt1v
PLITHla7GsOn2cXGeQea8BSlkD2TTvIc3grHHhedbeiRJk+82hyJ32A6I+petjHqtkByoA/Qyzk8
UK05O8PavlPS1vZ7wfIIErbjZ2s+2t3qvr3K/IgOvjwYGWUOdh6rlqrc8yqJ/OFsQ21Tm1/iCmJO
0CNaz8g3K5xmrk3ZWfDDxBDPXnE6QPAD0KslU+QtudolQx/ZAq+/dh7Ufkii4zkWxHj9kE10ZNAd
v6nyvNfMN3zWkhGuHNs7c7wIWS9UCtAQ3hfeY7yUWVFHIc7a7VtIh3Uw/jqVl+R35+rLh03Psgsn
YJZkjLrv5Ygt5WsJ5srOAoo43HVpi0cgKJ/y+yFPfj997uXxb7K5sl4A8lrEguJRmX4FAHvpa8JJ
I415pwdna1yUQ6mZ91LeoXJ5MQlDBT4bJyIZuynPES8+ASx8T3xNzCjfgpmxpBZP3O8RW15hY93X
i/z40/4Fp5JVBi1/H6c9Y9Og9wkIccVbOZaqPhsAg08uGSRqF6CE+WOzx++H+qxB6+9nJYG+aZ0P
BkHMctXDguZLW5FQMQ+ZHx3T3Lesa6ea76N5LTjGZby8hhdjmsvd8JKPEJ/DoRi3lok2EYygxGqy
1H4GTsDZTnSoMoQuNgFAzCAg3upmGV4jmLSa+VJLd0U84vPrukInsLuvts4iwNHOdxZCaM1taRbu
j/hwqUQDWtIv4LK/cdF1mRiA/GbdJvkexaCNn71N/PYif6/b3aoAUD3xASuq8D+jhvOmeBL5wiCf
9JBz0Oh+Vw9PVOf+RInxuQe9iPU06xddG+fwnl7wE/8piEwiCqbJnEYPlVOqLvjgNS9mFAi1j0EH
wSDXpoNgMmvodiNAVCvpxlrELzifu0TeVpVUnsPLdXFV/Ne+56QbLy+P1ABhxs1qGtS3LYS/lBPZ
saHZ+X0G1TocOp0JCBGsvCGrW17QwUZA+77Yzz+U/4g3f61MJOqMIBZ5vwQnGOK6hrtHfkjY1IWP
ZiLvCPLetJsDD8GgjBfgmID5Nh3g1kpYsBSIhAnpgRljYSt5rEr6Pq1kun3y+6rQZFkmElokFTkR
U2+Bx09JkbLgjBQoBxF78n6VsC+U/joDLciOYX7sVGKeNo9IBo+37frc8x0zbAWSU6opX8CMLspk
uHtue63qPQ6gF/8RjgMBdkWV6MSSNN6OFU67ZgZX268S8jXYFENDGHRBy4AGsJ/N6mu1STE6gL71
bTY35LQXKLImghHyRuLySEX8a8ZszRq9Td+9sFpOMIKxAiuC1G6w1sD4H4lSAjuzfhxIOKCAjTU+
Y1hVbqX1qhtwzKLF89qv7IoR8SFx9YBTbzcdZ1J09mfYnPZyYkxDR0Z+k7D51chacMZ6mFKcegPn
gdAEjXOI1koID8V87YpsjfawauJLVgfloL799LSrsM2qnVW9vkWwIby9srAB+DmJzJ1Yd8ERIHO4
7KY30Ke+thKwlT5LvcvHHV+mtgDqDP5TO67vjSxr1ZC/1TdDge5dqgaU8k3SlztQqPT4Emm0qYsb
hj9+Ru3l6pYDuNU6621r4S62WU71uI+/j+YDFwHa7LzLNYTahBVEEJwnJ82XPGzrkPFEw+q6+Trk
m0V0Q8bWsnoLVz6Au3Pl2LhLHwKUKU9puwP6xrIPCiBzBu4iPIV8v6QHGVGg+hiWgpCB/+7+FP3W
MzmtPDCLqpeKcYTySZyWtUDj6MY9f/xy6DXWVgdBGEM5u22OYiZAfgDdaNgEk56GS8IfxGe1Ilk4
+JTMJ+iBiDuBOHD0FS9IzM1OzOOsLf0QB4484H3YkDqf0KJ9hMDC/l4nCsZaYUwWucERKHQNnR1c
w1ii5voBt2UqsZOd4RnHFZTj4MTRfTUMSrGXrJ7xtZmSpaXnTS1slrjddNoWeVBE/utW+8hzcw2t
whaDxU5e+QC6shDL7LDb3AUT/eOB5h0cpy7EoGnpGaX97052rJWfqYYJ/sevTlb1HaIesKWyMvg6
FK5kGuByR36YZxvkk/D9F8eNOiKC6tvBM7V2BllqTmpHgr9EAJV3gUBvXHTNgOcD5qdsJ44llg0/
R5LLomCVKuv/d/zYK89pI9qhKlY+UMm9fy3q1LFbiCtModvsyhIzT0OX5p8kGYPxUPhWfAw0kA6k
m5+l5sDfYZA225P2Vj1gEwzTDh0xstn+cMnr9a7sFw6W40TeiBe34oQP0mogKKQU35FuKqTMoVul
WCs0NkrBcbP8OxvIU8YlkIQiVMg1KVSl5zP9ocoRKDqpbL8sZ3StBqkb06vtM5978TkeDStGgTC9
7H2Qn7+YgUNlfgA9ee+oeSIj4mzo0LCAIUVMtbqXZXW4oNF0SHCoJqEJWygecDOfBBCLNrNyFS41
vEZUNf9MHyDO7/0duZrW6Y21S3PKHgKkqm/CqkdifH2Eni12LQwDNdVlMQkQakg39D11D6XdbeVi
lkRWdBAh7m4+wu9nzOYiq4OWbKgcJhfCJLPJrw4iiiaUL5bk3cM65QJg9XlcFhbmtE5XVGOlNknJ
xlJJO/ZbrUyZxQkLLnO/NDJ6i5PCHmppvIG4UBP8VJHLuOSuessyHu6xdHWSoyKgIFDai0DMoON/
eAi+ofH9AnAYF7zebyMONuu3XGmYzS8IswUDkSvXsh9u7sUAigcYA50a2QtaLXH5ZqyJzYx3uVqH
egkmHPgTr+ibOnqw8cZoBSxo+Zyi5svcPUaN9SnRI/fu52KsopvdL5paY8IeUXnAV8yyN+WQcUYS
JFyeNWzzluDK3izJs8l68muObG01YMxjeQPS7K/lhrmREeBOTxjbsh6YloCiIgZ3eiHyBN3CNmEi
ctcEXtjecIJT3XLSUnVVxx3ghRbBADcJRhRJ/19RMJy5exRNNnw5gO3uOcd4UxSP3lxYCw/MXclB
309EHLjXB5otahBbRSrqmx3PrlqTIEpefvURK3B9FKSpb3ebV8OTpL/b6VZ1gdigsSWHbjhToNGu
yR8ko/g12XnR5lKUdHl4Bn+XkdLNJpfho1UFxEObMVecVqODhgBsEJhqN634LdTzRtNKZ6fBotfj
VIRLHgd7Q8fJl8vVra+HGnRYgrR9HZyvmrFtRC9w4ohE81phKPKtYROxJEA1m44Un3yXAbDGS7lS
rqgT3MUIbgnCjelMBG2lrs3Xh1XavYzcNnEoLFHZv6/DrZEAGlMwBUxSQ3ZGDy+aT1rOUcWydVQg
6qZnUsYlNaWFg9vy98diOoIBamHK1SF68XRLcr+TibA4nJocbVXmZE/Vtyueoa3L2qmxAclNijlZ
1fHzJlVIuNr8hxLsJrTlejLPeuRwHGTaMDViLT23sdDlEGHdD3M82KXR+SlRw7WAUWjS7m8tzN9+
R2FN+eGkm04CBpqpGeTqufESZFSDNgjJjt7ml46UJ/rL2AkspiT0bGJD5wTr8CPFnZNo2FI0OSC8
Wnonb/S5hgyfTncuDZmLjDAYhG9bgyfZa0yiLFX27Yp9QotTCiFc4TYDkANkFuzkQ8PN6LWFaW0u
ZrgRqnirUbGcjpR0E178cNVPz04+7KfpHpUfdA6Me3bVH35oYE/44IDRuS4BFJwkxgRegVkyKcUR
+eURbOZFdN7SUAtKCWxYAi9Eb9QpvIcdy2h3uklzspQE4HsO7jkQ9j5LZvU0Tf56IIgNxsv2rQ67
jIuUkVB+WpKrLsNkTaSOGPwM1LRz7Q9aeI3FpEN54BE8Xt+6wINGo9LSpEtIIoS6i+ym6L3PuTYP
4bWEZZ2J8PERbntX2EKxAQoI97ecN/K4uSqJwt9bf6BKZWk1b1NSQcFqwbah5qth+bQetHeU4hIP
M5RZuTBNmhvXFZ09kcGk4HXKFesywUaphaieH3bN+3pVdxkqPxunv/FW/qyGdOBf+N2K/fgVnG5I
Qrj8oUVPNOoZBtdwuziUKlwGwiJmLVr2QxJoLeOIrpGM6Iuwc18CiVFnnvgPNrng1PHvTHcKWUY3
Lpzb94BY7r2GfCntVDhSD4HGb55G+14TRD1ly4k5m3HFS55Evl6jy51q3mSV/RYOwKrsHjZmWxMH
UokkM43LYCFWGHwVpFPVN+syFX/RpkJQmM19WynUd+6jxGDuYuZyVpPQRuTiLMkr6iSAymszvFDN
CFj0mKjtXer6Kb2n3vKcNwarDLndoU2Q9K/Rw2OQrtQDGFX3Vbh4/071sAPE6va81HfD2rcdu3Si
olyA/4F19LKIR74d6fDqPNNV666ELSbzZX12IzbFsVayfQBayw577f6P83uqri7sQVOXHjF6hF7Z
p9FylLA8s+reX4Difx5/ioZtHzKhushx7M/qzyglVNlGeOstSlMIREg75Evs17iraUs3pSJar+yN
PycJ2fbWOv55HccWA8FzRL6bRmLWnCx8rcW93x/Aiab+yD4x7CR74ADPKL+Q7sm1P2B+KoLk4/c8
JkXYH7Co7H+Y+qh/eQ2A+PO+MPsIO3ILA5auJ3w3fFHbTxDtOPbVZCLJEFCuflVyt4j0IJxDdwON
Skwt74a2q/ovkXe7GjR/7625AAOZShOx1qak6hNDQMw6QhOI6oFPH9rZZeSgLn6tIIEUX5MfQ6+9
z3xScq7CRvHCFmLnhxIOGn0NToLDpdeIvP+OxnYsCL+lXnzqAK7alfA/1bFqz3lkd3hD2Lau2aFB
qWHIZd/xED0Ywi3orBlQ3n45JaeFE30WoPOup2aLUMG6J0D71Dg25TyydylzAfzqescEEIkRwUJm
6YNpeoussc692tEro9VIJvCQO/sZnQdUbTqy1GrIPPzFmPWLIduK9QmVHnuWt/eHCnjvkjvrEkW7
dX3a5LjVw9iBLRcO5DxzYEDVarnikzvG3WGyr0TRVH2jBL3fo8m6oaRqDiOpzKKiP+ASgcxQKA2X
ZjAvqpAORQLIfc/fSMkLJpmi8KeA8tnPaHJJ8KPy1JmQKWIoKnYRHEadx0pM4WFnXseSuI+GlECB
EsngRjOnHe9c9Dt5gjSp6hyaxaEExDI3RAEP5Td6lp7pJ0xL9XHpsFOk/rWepsoLcauTxAMCLz/n
MxRa3R2zTQUZzOErw7LRTojlk6xRw75nAhwFqamrMEOOFLVJDl37T/zt9UIrWnUZEA+L55oqsCzA
Rrr8oNJgi7nhArdOPGEHzeOpa/zdVx7fPvAN3amSH63k9szjGhNDPdWi47SVzt6XDtU+k0Oj8LVB
QVNVXeGOCuCPVbWPeMm7FONKoNUbJU5pscfNx3ONr7WLUe9j2uDfl60t5ueQ0X7FTsTZWdzkQ/Rt
Q9UR+IeUiZfA0s+xKYHN4btSOeB0sXatIdUFDW2MAmu5+jnLB5ddbZE9sr5zn9hw63jrh0mmHrbH
wyZqG/Vkd6MisPDXGxw8W7LZzSACWoUl0BK4ZO6dH1BfylPzEGaUJQCSNSCDFUTdwLtL12ys+08f
F7+31h1dWdXWr05B2EmL4lDcPJZPLk1M/SVC5/5urIB/JW9FzKjipn2SWvmjeimMEHBR+jfGDz5Z
om8RawNnM1WyDsh/E3IuPQzJ3CRy7NMqn5ciLQfeHT5GeqEgouzEFEn+YC+mnqfHnpCLv4VK0Hzp
4bhAyExhrGmEzaX+lTkdXrVGIA3N4o/8FXAl+4wbjFNLg1wXrUWUiCJ8o9KtZRS31WawuJQs9WJQ
v+3SUpoyIIZwZEDqJIjwCuXUDwOH5W7ilsbfhEeKxpUEwkhAPWosb7RbeqJSNX4QKZRIw4DQka/9
ABQNloP4YmGQ2Co9B2NhytJOm5rU3ndd+jNyRNh3PThmRQV7xHr+fM6++zMzvKi8xm2TPUiOEPIb
SyHw+JRXqh3cnBFg4SC3YOdf/aMrsHMXbNEsl2+8PuNOSenaWcANs/JunZCmL20SCIvX47oU6JEB
evUTX9YmidXimOJZbbV1/qvCFIWoukwl70I972gsGZfbYvB6bW92x8pcjXqtiw9cv5y0RtNvE1AR
u3CFOfYPmWSXEy/0DtnkPEi6Op2Al0FoGam2wLFdeQB2vkYWHWkvBD5DQhLgZ4vXo46awBVABmD6
oxv6TjOLL2PF0iKbYtKrENzoLolavjrk6V41WFycWaFrff4nYhLsQLSXpRxn3TeDalKo5mnkT2Xr
GTegCdKbacIYJceX1kV142IrIuvs3+sUJJytezG8bOwDuh+1s90UPMy72L72hMHHxb4RecdG+xyT
wdO24L/ILPKXLK1ulvdFK4y2mpBK7kBvz2TlJ0E7t9KgJwxv7c6to8xY/8tbaWNnUTr2Zjp216lF
/eiesUEYjXA8QJmyHetsXJvNLqlhZRtvvq/hOVfuCspNBGYou9OUVoBVIRnlCQuMvxLp6p8+s+8a
L8SefhdgV7gpe4CWw5TmEawNU879NmikFogi4TtRsOjjW/7Knl5GhY35tkGKE3D25qrLCURv9Yh3
VAhPqZ6W8rpetPQekhzb8DBZdgk6afv+OtQOUb0nj303fi3fA3QiSEYNaEIIZm9TPm/cpFPc2LlO
a3EY8/eVzvwFUYOih9o/Ern1bNk9gDfHtupnaQuND7qsjnvPjNC6vLfTFXzIb5zkXqkc8v0o7BlG
1uPdx8mF2GSfoojGzyY6t2svyZRGFowI6nOW60D606I52xQ2rM/AKECLLs5Xn4HJXtiE94MO3nMo
PSKbxD1SCUIlFP4LPH4tJPlaH2y+6vmt/InHPESNT/E30hbROSl0rqcYp3Sde2Gz2cgNknJViSaB
4fHFr5MRoIEpdRwNGOBUgEugbX6qIQ8GvMtHeSZ1SFfz1XdQtRX5Q6aH7u+oK6NyP+zcX+SLWNos
VrHG48OYaVKTyuqCtiYFrNn4Ao/Qju95HbH7nvZmki7a3m5gm4LQorXwLtDY6w8p48eC1poJPcHB
WeMlxtJ5thyIsfHVp9iSKS4UcofOEalbbLwxwkhTYeCH6RgpxoPB0kayPcrW9IJixoHuK3TF6/kW
CCO0mT/gdXTj8i9xNZ/9bAFPoy6jAj6+aATCJYidXhKeBmuadUDtfWQUIazNJxmkBuQcthGX8L+C
GH6H2B19AKax9EmAwpFGrq7McYiCraF77A26Kov+Kph0B3G1aDPjiojUvGLlJpWcmq89ibH0rVcX
jX4To7DMuKz5bqPsqLIbmND7K1kMvpjh2zmgEuxcVEent87bGxdEO6YbCkyZXXG1gPbg9Qf4U7lG
M2VhODbpibWD85FLP8EwfFV3QTYY9hmOCnGBpqN42Y32pfsZXQ6OmttD0rT11vVMHUeIUg2H8FzT
71HYJTzTiq0xBMsc66/xB6Xh8gN0KbE8yU1LtE/4Yg7JvvVZLYENgoWz1r4RosSAW52lqKHfNCNs
aQhOHpdgnjxdQ6Mxp4UOmvz1JlG6RjA+KHTCwqcY+HLDy3bed0MD3Y2lsSTr6i1Q4g93yQYN2wd3
39Qr5qEhOthHv3Lw6f7vj1apoAMPEdbNqXq7xJXfFdxj70a4VHG3anoM850GW1ao0E1HcqOSiKQA
5dLOn9kvzRxk1gorhsT7NNu25Z1rdphY2YDJblNbXoiEWQX2DtWKtHDb3yMLDNvsgCxEQNCjIUfH
2h0h5Qi+q3KQd7r2QbmUoL3lNFPYmQ+Ao3eaZkZ14YKSJh/BOcnmTlKueYCQoccpWy99fAv9lswe
XFZoCCht/JiQqUuB+pPGWA8eB9VKD8pLiY5qn9RId34CvbzPylHZrLtoNyLinUzCg5/85dvn8QG2
b+visSk2U19jqYPLR2o6+MEvchUwhFFGLBJVBypdO8SGsQzeXhHSi8sfqGj5jo3p0Wnhj6NG6Fao
9wkupVhLVb0Re70ypaQkxfG0huEpgeZsuezm18EUPStkrvz8MetDavTtXpJupuvCjWbQwFj9wkHL
WzXMy8TfES8H92wrTPGhlXee3JjqShKrtWH2gRCpiTTdEhjlra8Y6BREas16jm68fwzLQYAkzdXL
nWTV9paoa9kQFFx03FOL+Yf//iaP0qbrd1HBAefJsKUBVjdeIRKgrV3Nn7ZfqjW78TvL/qVnBVeM
hnwfB4dJaP+N5QQHeFaKZJfFvGpYpDFI4oLt9nKGGvij2QBYe4pDzjPZUQuq6ov0/7c4pLddhonX
q7YvimFl7Lgv77Cylz/MTp7Qp86k+kyWKmIae3YWZKUONkDQ2wbKP4zgAm3sPbiYdvS04bwvFrWn
Hw3xsZ50OmOqRO2vU9xeGcK6v0q0BBJsrTYhHjN8z0ilRGm9GQ45P+LnD/uhyk8FMLmbYO+wXIi8
6WQySL55sKDZL16fz0rmzVmeBpvCowIwV24zGySTPaPfpd2KQKsKcAyP1Vyx0LII9C9JVbwYofh1
QPViZJslJq50cE1tzlD18FoFl06nV2VGaZwrIWoENBP68om3Ak6lGwU27IzX2sKsNTePNa8GLwCK
JhA6A3G4GCkyintq7p9DZB8+awei1o4VZqhqkCAPtWzG7ExjkoQ9rVZfFJ+ynnBWMdQ224qJ4q8m
AOjo8vPFlbPj6PAVz0TEyqwXGtS0z0v2+9nhunTj0sRjazNPB5g8SeMXIjHK5tFxrv+5z25YqWTi
C47dW9abj+8mnlWJpC+J73aHqzfB/v+2SU/7wOhl9UEL6k2q9J+HZSFnqPsH12IlUZRwBYecUMO3
vWR4rPm4ficAJslX9Q77awAbvsXXBOHdfQoOHFcF7b6GZmneCCKXe5GhkhQ+zqZu+t2+38j9Fjh9
5WJau62BNKJUlAaWCRL4IO+5gabcyNCDjQ9S4alGOevi8ksAHqRJsl6lQWjMprrAn7k1SrdUndIw
uQ/ZaBozate8GJko7JyD6Rf6kt17zlt95naky2H0SPxP7yQ3/FknT3dcNCtLnZCJaQfo1CMtXe2p
KiuqIXhH8VKk+b0loMgmecjttCTw/4BZIb1A25VDBZnaX/WF4dyQGBm3TVpTAx+dlCo0tc40zm+F
MahnxVm+tAR2bOTOfbU4InhLIKUa6LvJZsBINRikK4wjQCuGeIcBDMHMEbMvLiR/6WGDRlPk81J5
l7HhyDkk9UlCmweVlQKhryVJ/u6i8A3YdylqtrCrync0qqI690mONfOepPCzIEJzHosh1TG1mqz3
NC1z2ryLnnvPGwBxoUksNfKnBLBpcnInMfWEmj/jyuzCo45Xr0ud7WThgSzYV7+WPZtbv3stB7Hg
wcgE/pUxApGNYIAygMtdpe1FKZ0tWJYvS06lHPn7CVFrLD+TlQihD7FF7dET3XpXQZ9ZzkDSvem8
Vkv5XszmtmrdYFA+WO/CX05YQf4OjnSwnAHzwZdxbymwY9ZbfEAhkSEghvLMmntu49iGK17paEIO
Xk05cxAWFCpjP7iEC68c+pkW72FjK+o2M0HcBBQNfkx58p+eOhIb4I6jAVzhFX8YrlueECHY0IX0
7BALlDJaALLDysKwWEbCcjRei5IUYJtqgwu8/TizQIDo0tqUKzrnxA19M9n54MG9LM5b0oJo9gxv
3wT3aUMRlxnZyWPP7MGQD7TfVecjSc2HDh5/7z3VMYc4WPgMs6unziG4TBvTBG6/J2SpEnmvCCzy
DotlsiEBjzPo0IGubEM5NnEqMqwKzpqqfgiLL+v86PpsiyH59g9v7YsBgSvrI0jEJiMmS1HmJu+V
3YAnEx2OxoFFl+pZlbd+TP5p9xPp78DkALz2fIu0VKC0R/kw9pogciulfKNNMsSEifNo/kTLfhvH
5+ui9Nx20FK1ewaH7qUMLk19xX677KtKPNNwhaQj6bLK6ewIWwTpjXf2i5LZQI4q4FHdI7V9idk2
xVmeH3a1ha8qE6wOAiJdkpoR3GXo2MqruvSvxI+vCua+c+ZPOzcgRjBisV0Qdi0dJSyk/bKr/KjL
Xw3KWdE0U+BEqnSoa3DrxWs3WkLoQqFAy1EcNKVhBd0ej2j5GX/XpVI+m18mV4dYWMx3JhpTVVNH
f4MtmdsgFwQYOiKtI0vVrBX7a8BC8vuxmqRaQahssaJ3Byr93rSz1etTMZTcMkNfE259qtfAaYph
sN6bnB+TWPYlCXz/+CkQiCIHoc2ccrRaIJXbdRh+ghxbMFoMe4iVVHNSwOO/sXZ6wpnVeGXGpi6X
/rHmEN2AZLLdrk8HCqlc5Oj9QEjPDwdw6P7Lk15aFjSzFX5nQuZopLHk9VUmckf6HB6B5Kx+qXNz
qclrY5MZ5F6/m6xoRB10Y1sNvszTRK0wuK1BfXIN/uabj6rD4v8Ee5aEeCn5J52ucKZXqSMLZceL
X3SrIRrutFIykznQtYJUYqcrZOwTmxXLzREE4JFGr+PXmcXlSEaIsI8HfMJ7Qj0a0IMyFxE3NETN
5haQcicZ89AOmgwuQL4U0TiLzgdC5d8Pblc+nsiSgm5Mq3ighuHyqzL/GSDE8E9h3o+2U7RRuQzq
LCKDyCZufOPR6UnKg0nmNyvWg+p+Nyp+5m7e1+g70xv5bTDXHwGfVdto3uZ4CLO6pPn7aGNlYJKZ
bTnuF54Hx4p9/q62Bsq+eTgsGHHVzvZlxx7x7CXTv/VYj3DEZLYAe8IXeH0rTzWEL9frrBxutdiE
zj1Npo+4RWhcqqlw9RODkitDUmGwJgAx/uq2//uQv4CkLa3HuJ5JjPf1L11vLDCYjDwUIYEq9lEd
+dPHPIWCUzR9KTCcHqCzyLDQTAwJxEfkzzw+B3YinsnI9d7kWrbJOloHK4kJXkV4PhO2PWYfvJ4F
jpdXoRJs/C+gN7U0N1RXwx4jnkp8R8BQoAGsF3MBBi+clgUiHLS92lQySwkEfFIzigY9J1PHcMZy
Ez8v2byUlr7OqjL5XZQG8zYhGQhHEvcm2t0ieKyrnT9Qc/lu+gUJXFCxmEnKbFBP1zTI6F8w8X4t
kO3YP5IymwqD8o4DyiX7vl/CoGnd8X5oHaYBTxJiGmGSHvoAr9DBNlb0LrIq+K6s5gs3oM17edFR
5RqPT65JB3Fr6vGoNye+CM4HEHpSwDV5btcNf/Hb5CfAvtzpEtoDp8jOYpqJFO3Tx5/QCrVz2I1q
9OCfM8A9GAQaHbK5t0msrgn0etmBfHe71GNL0oVospBiW6UD+69FvlvOnm8vsHCnfzOkjtzW1I5M
4BHPGEYNBfrNcqA/fKzpMn6oJRv9vV4sK9342+/j1AJGTp3DRAekOugb4mn+HuU474/LXR+P7icb
+FQL6Tj1/Dk2BkFwAalEe7PsCKEExUe6AZM7uHEGGlSD6+L3XEjRBecli7jKSwM0fEJyURL0lqCE
7V3UcIjeD0ieDISnVp7JWWQ21elRHxnfltsLFIKjdXAGzpcqRixJKUtUiHM+gKds0KipbFIuxfmO
tMQtYHlTrkt0BRnMEDsGnx47iJuYhh75uPIBfCneMmdiKGWQXM9+2sOfe292qv43BG6RjASIc7nr
WLE+Im3PRPpmw6k/O/R8xp8Z1z23m5+bJxbuoOVJg7aIEFgfJWCtlV71z+mkon9TNLWfOl5npr1+
xcTKBuhwWdA/BN2H0BYR7KBdm1VDdczx757YxB9sg+PHb6wZ6jZTmiWEVaikTUwkt39bysYBIjSl
VWAze4VuBwO0+5OIQpqB+9E42iQMtdISzMIJWLfYl/9Y20WnIctvNtd9DaDeWwrVFMjrAFJ9dkqM
cpE/uhcm5KEyhcPKb1MxrtVdCNL0zsYFCh0z90g4lXkZbWEGVXqG/FhvPT0JoPTG9m4LEBtZZslm
go+Wnh7sYoTpU7/BfDodxz8gz8013E40WshEmGKY5BjBwzZYdZHicHGAF+2ni3XRpfRVW83IZ8M0
DfsTCozFLiyC35sKfmTCFCinuog2Uwa3ZuCKc7k2LO25uqrJFJbzOJFZfIhAxJ9DvNYyeLBmBixj
8OkO62ytAO/nWesQdoHLaixXn8Ai+OV9ETAgn10jZgz31oPBheiLJ7PsWEj+W1dUohlUhrjmQFjx
eeqQ1IHwzGwpBmJuKZXQGx5mzRXPGqNnASbeyigUDD+r5MlGYT8kkGUpOB/hOI2IJnGsigkaL2LD
ihAi6NMkEmBycYIIQcWmXxJW6qpUlWHjQqQJM6QwNQGGVpbg8Hy4wquR4In4CcvbqqBNof7q9NBO
iPKp+dPcTXuNxlEjORBo8/iTawa9pGdX9vRuHh8ydKbiqjQEgxUo+aMmTMKb5/GhTbMvj2cnIyrO
K8WW7zuBKBM2C2TqieYnQ8UCBlQ5MADN8CNlYmq62y9iAjLhZTlNNfDBOcq2hEwBfOVkiEPsheec
CMYWRYeYu3A69mjXl6ZR2C43R+N3Wtynx4Hq5g+5Ra/pmC3OtWe3Gu5ynXRL9n6GDjMT9baWmSuG
se7MoQp3WRb4GkV1G1WQBst1HG+oDtdGQmMe6n453I56ts50lEvYJotioxsR9qdk1lHQQEkeJdf5
JRWhf1z41bh/5I/CUA+Vfr2QuYryrnL+rV7nDd/i544slPbGQMs0v6Mg9HO3QQ8rEEvR8HbbLM+r
QUq+xoqUKo7gxlIrlBCccpTyVtDZcyTRDUYWkKFkSYp7MH61q+DbqGalwjyGrcSY6bo4ix4F+TB2
Nz4wrBNaqGc5ZxLmRcJQlMGGumSPrNKW7cujkSV78TSa9woEtYdIhMGcQxRMoRwgsSxkaHKkY3OQ
yVokpg2ZLQeJCx3Sdhze20rAVOzPDkisvL6yrHOZ2S3Qt8vf+b+CAEYCULrUJNP1r1KDQqFJ8N76
xgds/gw7Ys62fm4PKl6RrwC2IOywbBotY4LIwB1cz2+kMuOUFBcxRaz/e28CcXt/3mZXW0Z6QYn8
MP90nqw52g+RiJ+TlTqxxVvPuOVYFsET5Xd6WJ7xMwT5Pykgt8l53I2wGl6YmuF12tuAdxM8SBSA
5w5rUcaIoxDoJxkpySWK/dLZwOK4RjsAWK4n44/0XpH0v5LT4woPAmFRAn6SV55NRHXm6F6r/OiW
wEaY14kojj1N8hW4IDkOHIz6XZjm6L1xEURRfkwZBFyrQYjHhusV33wHSkymaJeR/KE8UHfczQdp
Q6HxshqMXkfVdK61lHuWUEgXweeD/fdBlYDZRXrSpGZ3Wz2ou3x/QTcGa6Jc7U8Rooxrnynzm5m7
0Egwn4YR8DxqQSVB/7LYpBWU2zqmUGwO+oHg06EGfR4JGn00is/F3hZdo51Y34NmZK/c4Y/dZTZe
f0b5lNEQPhj0W4SEnrhLi+3L7Nk/yP5q1B54Rns9cInxy6PqzQjGgHvQt9lP2OjzQzY6nTBSyp14
h45qdHlRJPWaBxrpc7fwvTXW+2Pnh83kSlH+7iAf/Y7vQD7wUn0QSsdXukDntkkdVBo5q2Y4SRS1
zmOo28Ls/vfiCkO2Ynd+DBBfKY4xpn0Wy04sy+YPonkwjO/tWN5mvDc8i71/jW5ZxJqxO5MQ05t0
oLge+cmz46qxOpwZ6AFbr9QCE/pRFYdBQ5DDEDxGZkSEOuQov84OJcQ9e/NY4rO5skov4IqtkRQd
idvRinyUZChke0F1OjPjgaKqegBBrhtFDSoeMdyvIJ25F9Vq49PcS4871pRnJOuKJnAXIUFgxdxX
p6S3RdAhv9L1wRunwA1BckGZCGUlJYh1HDylcCrr8h8gFAGignXdDbD73XaNk2uCdOYlUzX33U5S
gKUQJA08rmkJzLGaFCBoNZQQQcxJLqsoxsB+1suUGVOc1qTkOQ6ndW35PmmguLoh2YWhjqVTnW3A
8Cd6W0EFK0krZCFQrzfjxtlX3wRb39TLkoF6zjXffyD/ZG//Wj0zt/2yqrzfxslAksCjhcEkWQN9
zawnSNzQ+ZTlN+NjrrQwohsbQk4+eWiGCrIEnxCnF1X0UUlbVXQDq7jaTkI1h+u+VI9FIyqdp+/K
1vRIBboNkFXyIIea/ACSuDPd6rX7D+J0dIVtTwRiyaQQZ/o8CURj7S/xkNfix23t8/J0pK18VSVY
e5YVo+cchJr5mLC705vQs4sOqb8eD50RXf+dcAsefXF51VhDp7K3JI17n3L4/JaD5Io0hpTjMjB/
JoTAoDe3TmFy4WF42sGuWXtlC+cinnwEKvHAZl9NV1l9D7HCnYHidUUvSnXkuI5TsI99A2P8NHuo
4ypLil75MmROqudn3fKuCeVr3CRZ3hg1wJRfCuauf21zi/gdisj7E7+WLze1SSfxPhAg86i9YEIq
7u+tR7KtAS0oHrCDFM5F66vap0gOu92Zf1g2AOz6RajuVwGzUFr/zjJx56H72qlgY6fFBa9I2t8F
m1PrFTL4H5e7eS5dz2WaVP03F7pUicqwMBRi6h4Lav+ST0FdZrN4zqV/muO2ibYdQwNd7FEkfImC
lUSxkX6KLjRuH7weEthK0f7/EEKNqpz0huREIq585ybUkYBLJ0HGoNUaROF1MbNAoCw8TjVK4zOk
3Ytf9ytayeqVXLLlpC6J5CRN4lbKlr0FNm41nPTKj7eSEiQSa9haJI1O9vTSJPSgCE5o41bvwml9
fIYElPzj2bPWdnsPcikcfQJtOtXbBnX140onuh6RfMvQ3BNweDBvGwuqbYFVJFDOFXmfjHemsFYX
GYKvCDpymZrevjtkR8EpeICc3Rls+H7LhUdDoNFBeobipmBGgarjkYpFYRi+hC2SH5yovz8S61IW
F7Ga15vRlssUtFLXU9+LP58zhNQQY9IhuN1zDMlZTrLB8APj60Nr/hroXRfubuR/IqEFcgApv2sQ
PmYPvW5tawiN4fDB8Z+w2MeLUnMy/dIKml+SgVfQCvuxJeT2aAdu3x61YEMjKIi2z3rgf4mI4w9a
Hj/Ioor7ICFlsYK+N8HMZ56f/2Os1xTRBMq8ycD/c28wI+xP4DgXzsm9+YlSIL67HwHf/KtEV0DY
n2d163lgRcUlcLl++rBV6xs/+DEsOH+VZN5KMevx5B2LMuXjBqKHiJXQTilPjmig48PWOp5mSEHp
Uwln9/CjMnifvwcFjKzRb14e95J5dCTIcpGhsGXFZqAvyMUFt6L1Zf2u05k+TO0jJf+zbzW951eU
tRMhbhQaLRiY70DPZ5pHL7CsQTqSjoQJT4QU+FrXW9Q0AW8Ved68nWOrrA2Fjk3uRu5EwyWZdQHP
ANLavsHrzo4pozpZ2GR4RY51GfOmSzKodviHhrNHCawdjelwsxDoK8anxLC+iDHX0vMEfe609MAT
onbFkqhLmv9ISumTeZSojnNHHHXtTPABSViMxnz7Ku8IKYqG6ysBW1eWOBCdUo9qBR1LNgKXJId6
yMhc3HpYj18bjmhwYV6Dda4jPjzQRrueL9xmmamGcir5YIQx7jdwYneVml7PcxXaAdqTC/95lX13
wimUB8gJOTlnVF+WiwJkB8/ALsjBTqmpWZyg0Y12UtDWzKYTZvwPUANv4dpUGY5wm1zMR0UX2ur3
V2zLzCBfrAKvHUWBYQmkXPL9M0kgIpe1HbVnv3UmLCzwXEt6CVvnMrH4z9vHpzBV8X4CZGTIad78
49/6oDiHYX8CMyV4mbXdGhlTOt+hB5fTKSUcycqJVuy9/nlYaUPfRekl1qKEA8e8tShKQvXlIKex
I1RdQAjpAiFr5g7Yh2tllji8OxvN2OKRAB8HbIlycQh61Sx3kHrMXboKJSnS0vqt0rf/wCmpFImv
uXjFkPcvMoJFdshqIwX7iemm+/cKisPiDmFTGduMEpbvK0Fkb+/0ooEh8Qjy1eOdiyX5fbPoUSKB
wxoo1YVIhAg9GhGuuvFeugGCe5+gYLhYhJfqc4TzUiZ5dYDqzee5XrnSVAqnAo9U4Kwt8Sl+CSoa
txEwXAjgOnu7OBFr9+xhngzt10KsPoUIKCnEaiWwEvJ/T7jyy/1e+kZcXq0Cz/yzy4hdEni6VkHJ
KnMOZi96Aphd8aUP7xkc/hGlwuEM7YCgvkA4mpVcJxq0/XnLrdv4R+BbQs3y2csUNCl1VZA1D/GH
mCaL9IOBT2ytcZONBeX6XZ9lsunMUzlvTdLpbpIUN/ynAgfBkRissvhJIoehHhq8XBd+sXOGCg0i
H82r0UJIRYm6slKt/XVmezOfex3WSXzebi8C+ISDWK6tLKk+h7BlR1v57YwgyHvUOtQRpnRr+vgc
ryTr1e/UuWeHJ8JGFvxSvAZyKA1ZP5t57tA+ZxTJrR9odMpO22ETvQjLrr5glCMekBL+N3jKBx0A
JmJh9AaVA61Cuzia9IDXvtte19BKaRXRsX723lhbgovFdtYbJcNQGAnEfVLVtU9PXjWtTYG+vfIe
XvBr1OgyFDyni0nxbvXPCfnfT3MphwaxwQjdc0DNl7zXPsv4Bz2eVqXfRo1BqR49dCZbtfWWlkAZ
SpYFh6iUQFBn4zPWsWSYHA/DjYv+zDCKZCeO1kDpO2dImWxjA4uBqlS82nsjYubLMczbFqTvd6ti
eBTc4ZTDYeV4vRVet7Qn8NChsGpIlwbQVR39rXH4ztxm2BsWcAl9vYZgXtpSxZTpAAczEo6Akt/0
N1+132uwYPowr++D6tMVRYU9QQpkY5acMepzWUCLHiS5n/mDQx4RyqTFYG5OW0C+inwY9ntgDBlj
EtksSUYTJIC60+Qc1BaUyGVcMqguGDE2mJVAPhWoIEG7UUkl9x9FRUNxzfDjHmlegMIVqvfGRcBc
9vnVSUhEkXKHnE6etGyn6luUv7NLULbarVrbVqMWD3LRg6bdykDVafJgWgNMpxTwJT+Ty/ERpJE6
OIfqbwcGNnzBZfxYrSJCieH2ksoR1PryGSVLB3k/njAluvZTsBCpFluBKeU15iJcfCi0RPE0oTcs
4rluxoZIOrwVmJp+YCSq1fkJWkE9P0G7/694CqIZPP+6mULGttCTIFN8mNx0WgpPHa7UeRlX4qU7
bni3UpRFOSUQaz1MkOdxqx52OOMsE0Te4Tv02z/YN1CayasW5dv7oX7oMQJq4iG1svd3StLsn+uS
C7F3GDKy5ZTzozzhaT3JAQZKmf+Wv2//2CJYJTyFvwPtm2B/4VTsSbXByXUKCAD3Tx3vtFmR6YCs
Uu+dT0VxY8A+oVZq1d1ESSdUT+Biohavy+ojCA+2HtDbc0qCsNBzKdsUNwIPprvprvCeXj+Ojrl5
qFMiqoxWrJdVBZveucK5Ylm/csxpKlM9AIJBjdU+1WmHSF8UmwaB4GP/OdzIj/xWaeYCBnmhR5bl
2zhJufF4sSCOZyCBkpdpGW/VcR7Qu63kVt57Gludyz2Vq/xFU91+YYuYoroVsMPXCw6LE5JYf7vE
SUVPdihKvrj3CdsAnoj15RW7Az8nTcTIgT//FxA7S7Wg+//H/MM4C3WwSJbihzSKELYXRLJE2oGj
PXwpMqjry8+u32Mj+3eTqU2VusBbQvDf/FIYlfvU0lr3MNGiOYiOnDNiL7LROiirI/dWTsDuxRSs
solzmgNYcDsIkzla7r22svywDf2vI9acl3lVV9rsszLVVQ5SjvNaSYELufjIsHE1RiKJPARavFCu
z7ywfgR6u3CCIFRMa5Q6GOXtPze6YjQW2ta9mipdqhzt74tK/vKxv+irUebTPqDhL6wTpy9MTmFq
sFoi1s6hXMWorJVdYenDXcNqnvlThVGfIp5/Qo1dv202NcOb6JzqmfQM4ce0m/n7+f6dzyZ3su3t
94dk91OyOW97ZEE7Untlhuq38Y1wAz9UvNl9i0xXcAyotfrTTUpfATG9GXzM1eoqYFx2TkEiWQaW
QISTxQ+/IA9UWvNZGwdKG8O6PFGSAmEmv4l4TSMUTsfT0too+ytAtFZSmZgWVU475pwD/c+/MJzW
rvqD0nLhMzMcCEa+4fu5e1kBEW/ltg0J+YwkXwEBdxn/znBVVgpcKL2MWhR8fDBBTPdi0VlEKyJl
cHfPlig0UCG3Yssb+DA0wPKOubHFlJDx9a+BRjZ1cJnoFJycJnzXl7EHV3ANOi/LfnbYokpGSuV/
OlAmCRqYK3gTceLZyaVGNhkuQdFSAWuawjIbcLoqnOaKuC2fwGPG/+SWVoimv0nNBR0tgbxjeVYG
q1HuRE31ppI8iZpcHbUR13BgjkS+vSXa1JCJZEfOjYsV4hs5gs1Kn6UlQBRCURZDlWIqh9r80pl5
7vQ0eonPb+Mzl8TjeLlfeBZnXFtsjnHV93V9J2HAaBp+UuKAw5Cs1mx8donR2kcwO9SzLma5C+o4
6SFZb3yMMemrNjO1ASz6rIC39VFT4BikRSJtUEcNCynQ9VCODXYrG5dKYzrHM2WnCm+Tg62a/ZpD
VHsn5SKpTopHPaGQdRiiUqG1PzcMpV1V1A4T7IeKOyQQ7lygYNS/5RxyqIe+HxijyaP7oy5J5wmg
HtnMVNj7j54BhxVZE0W/Y+1Pu4pC5CFuheWxcngQuN2xsE1zGCMnjiJ8+swd4KiKgeofiQHBNg27
STlxYxfHIkRr23PqKOnInaMEwx1TFU/b4f8FUT1hkd+fyssDTweYZeRQlTOvqq9u2sQYCMAelVW3
yOO6j/BQwOxseZD5cQ/KuidaQmvOimDvd9krndBl6I9qrllnvH8myxffvnLwy1IjIzI3knYiS5E9
MJGeaRroEChxvwoab/GIxqUFW0Tb7FEtHOnJquJj5IkREAzxANODpmkNXVPLssPE9ODZdlzukWol
Ww2hWwtw5E2MU5UKeAnVsrN5YmWRxMHZjKRb9wCVwMP+JJg5zZ5itzHhCrXSYT03VICoeUk4feCN
4/+CRVrTmsGF+npX48qfabs815ADBBd7w7ydZXSXA6HvRQFMoikLOfrfdiQwyjMgcsaZ8a+Cb91G
zjRtSmYjwTusAB6ZDSmP07a8+H3hcWCpiRUbSxe1hzlj7Y6Y4sfqYQOUyLGxdCF1fnOOF6YoIa+z
UU8GAYFsbHEn5320LcXZM8gYXrMfTTm0grwEjUIhzWFkM1ztPIiihavHEhLczfIrgAJC8s48aT3f
Vj8yOQoGGDSOKNxLMc2M3TbqU2YKga1VNfz8Y6hyyru9QHuc5qt9URZAFbNvFNciiSMqX7SVx5a1
WaGAndsfY7Cur1QVIWO7t5BU5byE5lOWrexIW+voImzU24epwJGQ5VDaAAmnH2ecCXFshK+gW0+Q
CppajlJKuAfCO9SJbbFOt+v6NwbVOoJ0Ktq34maIFV+YEVNefnFZHV6JgLkbSHjprGI0gE8wOJsl
wXxG7n8s5iD+w8QmV8UScgVE9kNtuvH8V/UcOaap0hkF2UXvTm9OqoXqcVaERw4b4KTlki+dPca0
XD+bttGAUzBNHTWSvhVCeBWzzXxqZr0Bl90vASbBJ2AqB/6wZkUtg/Lo+MWXRaJAK6AmOXEeTGXG
P5hczvf90I5YUBji6JlQLVWfb8XNiShLEyt6aaUzvWhAxmS66Cau9R/dtyurTkFrtM8DAyjCQvyn
wDlyhCXzfD8BD65pMcMW3vtWXpXiGcZkSjY/Aom/Nz9Uh+S/AuDL/mZyJ2dhGpxyvDLwPju3Irrp
AFqzqeav9lyiRmfSf6EkX5H5HTvKAue3s63/r/gKd2bIVeYqpN5gPc7y3rQePkdfYuhnLl1vqA63
9zZl+ErpGBml1ZW0uAaFYFZtClEhD+rRBvncAGHWd/U5/ymPi7GxH1nXcWD1ZSHDu2yM4pKaeyRu
aQGT1B6qRMD2tKd6PMt3HTRgxgNdu3YX0l7QxkHqbZz3tv2Upq1mDhlE5oJvRnJPzWLBJvyH1kHS
q1H8hWMvsaVBMfS+XJnHFLDITH/et1cJgBIN5eigEYuWdnVwpDzxbEHTom/ruI3yA7gS4reNKUSN
toTGIVPzfjHRVWdrNUNO6wm6Y7ZCjvuMlffN7rB4UDQiG3SwghSX2thNZmZI5slFQ0VqsB9beYW/
MBhk0bFcqzwzT2KyKfh7Q2ZtdQYazUNg5jHLhmr0AmpMSr8HtEQYZm5Wmw/T+tVHmaRyyPBEih6w
8jbaG9UEPAu7UZn1nVB3lXz4IbKDkPTWMzKjyGilH8R0HJttS8AMY+FnnVPcvi0GUF6GM0XwnfFl
hj2hrNsixqobRIsGl1EajnYNxd83W6OTvBDNXtZiFEitxvHhIaL7QwPrcoIEfteyalYRsgWkjw+o
KbfQH/8eS4qcnvS2kaETm0n0T8zrWspd67boYLFJyIep5+rTEAER+r24qkuVC5iwAhHhpmBNoQ3D
plFtFHxh+xGm4r+LRlnj2IGCBQ1HmgdUc1Ka09VWXcQ/YA8sCQGMw2RmZYyTJ+FUL2+5C6ybPoLC
2lIUT3Ek78+2chD1ujGfcW0b2fk6lq26agN6lHUpxt8qJQECCCEmQ9NVpvljfgqtE5pZnrhSd2G+
4+fjyrKJfk4tBW8wND6bgsjMRGHxXpQvhkUuVXpDTc7c4N67wWW/e/yx29PuGpgkJWOjcaVyaYTW
9CDsJeovkFcsQPycXQ5NuWom1qRj4YqwUjgfYieJKaDSuS0s7FTLzUy53jK4ZNLJ+vIlzj8hKT3o
5fkhUdgz18qYeDZ5db6DtGXLHSsjSdkJQ8COIoXfDMYTTeYdmxXZSCT3NBOFSVQSw5840pp3JU4n
3igYRA+AxVkLQOrRYtCLfiBx10ga+Oh2Hhgpo8K33gkJUnz5z2rYRQO49qG9CL7ZfioFkhUMJ7ao
BoeIRD4y3cyZ2AVIomI6EoHGCM2jWbcytaEVPd0K/uTB3CPsX15XNyKRuZEWKZdoOsgXUtneJo3N
ZI+Jmq+c78t/BagM2DhwOlO6Fovdd0Cz75qqJlhCQR5+pWvT67n7LHDkxGcM6DwLJv83u3mbhEzg
dXyFdfw2GJ929tJQihC1bbD4YYktaTVu875EphYQBLnCar/Lk2u+MEFCb2D7VMAiae/BeDzUm4CR
UvQYc6l0/SlaPTBbCQWPuXcBMuzpTHeH3C9QUor7WFPjFnah4qaRYb/EuIPrFxuzF8Hjmh7BKt6g
0Ju/RbrEQJoz3FoveNI/bdgCnoDZng4pBt+s8cyD2ulB93JbjNCvSM//rHJxFP6CxjVxkukoXcH4
0wuaGZhu6mU2uft9tXPDucHURdBdzJZGgFCO5C/Yt/773a7zgOaebSIeDm+xtKJ+ScngKJIvTzDL
W5CG9fDxsJFvUiAOldnvGXBP/kRj9wGUlKlwEt85DbtlVErkdGRukUsaLJep5HweySssnmrByT9a
/4Vb2Kcf4/S51fKhAUsKhovHalbt2QVuSAcMqJ/DqFrlShoeHA/OTWxrkyGoIgQ3DUCqNSOMIPwI
gzFtPA/E6B1o7jv1qqus1fEgWX3iLI3geIPdrn8NY/ij+vc9TXigD/H27Dow0PWfbMg//aFkAZAJ
sLc6NhxOBbHdaS7RSz4f2sx48jSi4UJ0FQCONQ9NwAglPPdm5rLTz7YN6GEALBv9LZOmyqZTdM8k
f43Y/GxImyazg24fUee/Ks6bTm6Q8bF1OzDugYTIY2qExnR0uExSd7RtLu+XgOOusFauafb1PldR
ssYMzMQJT8JEC9fZm6HTyeXkDFwabbos0+z3sSQvFGaKhDyov0ipYKjWVsJDMJQEOfl/wCUlmwPJ
Mtq7eU8g+n7Tp9y8zyAlkna1XqMo4IZzwIV6q9JqjYSv3rSBsJ63JVz8azAzxahpmNlb2Kt+/dUq
qOQHR+R8IOxhM9BCQsAdqWHHPX7ntsq2yTaO8AhyaNgPl8Ec1n3Cs8gYhCZndmZ8tO7Z62zeu/pW
pUOoru21QvYeearDJbEyy8CDUh5N35EgbUhc5KLfnIgAqupba1O74PxWj8nUAKH80J+AYZJ3oQ93
3HNqdeUPdRva4JygFuW1KZQPmuO0n0tqONfktsSACsww9vdWjtaEg/zRxuTsCukwYUUsA6XYe6I9
4TeyMDmdJjiHsq29glKMRzJR8U0hp2DoCJDWB3B8oCVmtr6OOXroYO5VNdmBJ1j7iwrkpi0LIQGu
qwf1Qyb8+TDvbXrp2rJbmG1N7N4wTDmyaOGFbAIaXn/3bxzFTc2zgZsy/N/56FrW10okqahD8sgU
gW3MysyVsvmzYhHpZdRv7E/4lTtkKjKk+p9b6dDNXn+tpY7vmtUMrilqnNaaU2hPjy0LlLZLdMXp
KRR3DQoFQr/pK/cQ8OvS/KjaEYe/jpua9otb9F/b7q4wl2T3iStPVYF6UN0n0EmQGatyGbG7trHZ
Pxx0Owh4dKdLSKnyKa5pfxgmwWi5/jSIneZTyW6kR9KekVNLofrpJazPa1E34v5p94Z7V43KaCPQ
AT+/tuFq16oak0kVw96eD6VCd7a0/Vk/c+L/RyBjXt++aFeSJgIUo+0CaMzp0EAgldYapCz370AE
yvqj1s+to67Vfu/0GPBaGfpSluk4YHBCoCwvx+YLGx+HnMEclzydbeoL05fhG483IuSh9bjI5vd7
9V/BdQFBrelo7lSRqp3GojrBU7u534jRJMW/JYgTgGPGGucRHqVDSTIJrpKaYvI6xddDSyzX8A34
Sdt6jQbPShBR/DfLIUWgRb48OmlkrCry7EHyRiZ70Gn1irmaxt+Ekmfs517/cFiset8VnY10huN5
711zFBlUnhUSBKuGMcp1ZmHzeLNHY0BW3p704WNYYO66IlameokyYWC0dz2Anhie26YIN1kdJXtg
YLDjvJKdmM/v29P3HYUIWjAkq0+JGXUziHsDdvwisaqvkkfLL1e0T4aAP7AY+FzldA/5OhToHe0b
XngTOlRCmZ7KEXxm9U9c3sM/oiTDw/ilI8d/Qi4TmdwMF7kb+CmJIF+ip74BwJyM2xa3NmzccE8M
dW5kgbmbsWuI894VXAmzVS+pyvS2w7saeNkdJjO3c9Ky+/J17NgrdgqG2Re2sSzMZDw9PcNFVmu+
PBZmmZ207rCcWbbwX3TJ4QERSg9unncBKk8ADYgmazWQYGNt9Q7XmQtxbE1rIg/JzFutKOgnTPaC
t+lmRSOhk5n3rSK43PY7BfZJnunMuXpSoJ2SInvW6JzW2IEg/ihKJCOyEHYn4f0HU15VMjvzXgyi
HXWI/eTuOVLnsncE59nIcYRIImapOksT++ELSqlo6bPaBCu96/6oxBg+fKEIkZoNNmF4RfdjOuWi
cIk89EbPeVIUesPsZN6GvpiLdxIahFgaxAcAk7tGswI9PpeYpN2J+uBzDcL+QlMiPnhtdnwYFNzG
gn93wq8n252gE1BWKO7gQVvBGqo3XosXKI+3Tv9q/vc3PRRCi4oX2ZMzveTQ5/YL2d6cbPJs6jRF
Nf9jv/SrLOwmnVl9qeTeJLWmHRYrNY0MaYaxh7relW7Ukdsi4MySEaYbnqxMwgyaM261BZNogE2Z
jAi2zt/2fcOAY5ZbVo2M7Yq9AxsQJmJjatN+3ztOJ350MKNWH03/9v/SgBM1tH5sVTp5Kx5K+gLw
RvNsAoy9Tnx3uvwqxOVUlfPj30+IrYxWUATZqRMHTh6yPNvfhR4xrya4yYNZJ1TpJ2YkfOdVHMst
ZBoaSNbJ+8ZFWNUkEkLCj07/v3F+/fgz4C/3q8iGmAAMVa6jaqKOENIaY+8oJYjxfJKfXk+XZF43
pxingb6E5POILUDCcfkm3jaEjZOkzhCNTYhCoiXikVsZzikrq7BAFTA1Y3Vendg4nmaDXS+N7tvc
m0ZL+TiepUflCZB19dvWc/GsBtZEPN8DhpKUD1bKbfn9HFy+w5btbjD+eO7IVL+SgLdxptHpmueC
oQHLOpArbkRHOR69m0wN+aHRAFzi2IR/O6Zd/h16ed+O9VppsdQS78WZ9Siirm72icmn4XHLvmbF
gCnZpE4avbFY2TYYS/YC4eJeSgzvxcCgN+aHF5zxCsU+vNRNscUVdOqbEJ5CXiODbX6XYWO/DUQp
433YPx+/XvCA7pL6SJuYjCZG7ooUZX1vos0jkgb0b8MZ6lz5ydu4KdjzkeaFISVTPNqGs8CslUZb
DiX1fEIwXm0J8ru0nLVVqcaesNfslUQlw9VF1YReoKjNL+8RN+iVL6RiaJx2CekSt8IoNJjFFb3+
uwoQyeZz+FwtbRyvDEWNrYfOFzAVV+QpBC8ilp4e18v43Qxowj8tvkDbBCQUFbvMnMfb41JDBggQ
9KLtsjj9mOJQ6YW9ApuYtsTsaXtHnbJCMBFKFKzDLxgix339GS/CGRdgVnZyqbuc40fo2Sh2pato
pqwXENffYLftLtOHgMNa41ekJ2/ZcJkPFDtIVbpXeCJE9I1oAEnayT7uVOg6np023uwa8EQB6a2g
vS2P5QnZkp96G2wcZKdVTywGPbyaDrxHVVhTlbX1WqXAFxJ3AgNsAi+DVkLQUQb5LxwBEJ0ql2eW
QyTzIK5gEE0lXL0ycbylfb13aouVDOK045RzSsZ7PeiplpIn+yrBliTg4RhvZc/YjHPDOGvcf3QE
wS+Ju+IqYq7SMd9+RV2iX+72kZjs6o0abc1vtoFjrV540GbN5BLRxvVOGBjjjR/fvCj2ER3liQyq
cz8Ry72xmYFkFRXK32n20vqGFAK7xHMJeOnIC4KMhW0V29i017s6Q895+/HQB1A6Aq25Bo2WKzAJ
lazZpD3RlS6Ohl8WnyCrLz6JgkWtlC/Qz4APdFzN1jjU5uI3Fj04pTsNC73XgV6KD4IePpXHFsN8
LjCDz7M+XOxaO4N2gXC4I3M3JqlfQ3WKlDIQJ4QMRCPBAnnnScu2obgxKNUXBGUZnnlu8RaSq8oB
QNKJfkRMEgh3kcCWOK6WFjrzr8UiVxnRg37E+E5fO+XT+gCOxS4Et71DvNtL9QUadk+9rq2+BWc8
gVDD+H+Fx5Utrp+0J9hfXYeOWiO38/3iz9MwYYivCbP/1AWYFbFIWcW9DglCBlvPbM3OXpLBzMrk
3egUJk3YdgXfDfK5Hw7FG8K3NYmKnOfDDxvqRQVkOZG0tptIrlNyr2gr2AT3iBTc786WM5YqhFK+
iskE719xY38l3VPTOti9qf234HlQiEXP4yVqnwbNAyk4slzTls0VZ/yEuBVIV7vcYz9sT5KMCDdH
LF/qM54FUPGapHkEMvXc+Xt+e8V2+WUbNixi5Yk+aJLn086HSmnypF4jKr1HOhXSCS7M7poFtaHB
qyae56vpFllmE70CZHAR5V0JfsE7v+hY2EZsJMswpzvGVIim8jJCD4ElquIfBZ/DJYz1S5d35XK1
4wy8JXNr9HQL/+foJo68Uw9LScIhRWz0X/UR8JpSfekozLU0COiHj/oVLPb/VVRPUp3U7zSQ/6Lt
QKZ8jldCopz1CcOo14g/rqayj2ZAIAO63/hJAvrEbqADpQ3sv0eiMGE0ogCJVoicHb9SaMx/u3vW
XU00uRoBvqeiUlG0r6jGnoDZauNUGUaAc+FdTm/AJDYKkCopeqJwzTamzAVMHGww7QBHECqphe13
4PEoVOHq+DLBAOqmKev5gpwjnSj6XCZFoiVvmUPEK06JDJa98junxzghhy63QyaCx2ZhEkNDUCuE
ma/dk4405vOyNHe3I5H1oSRixzbmSj9w7asEjRTANIIB34UbwpMzawgzcZ0g+i+nWJcPKjNnaXpH
yB0JjtsYLeHGNvWNnRY0V9r7u8bf16vRzyQNnbiuhkMtHPi5M17Ve1r/VblZbZnUoB4/zoQ71SF9
apxHWLdqfQJ1mofBmWOLStXG+rmhJqS9lIqQNNf4aNgl3usfBy8Jmk8tWkG7mBlWgxu2x8TrBXeY
ZV441vaqbRIP6rIl+6+ICNP5s2h14sHSDJ9qTrY5aFGnhEVHx5/o7Hpfko0hq4tXJ45esB9hlqG3
63CigPvitaxRpXUX1AczYpQca7EbdHhMbBpJ/42X1IW4jX2ukSjVfNYDRrbYPgqTVf80FyCNIqdm
wTBi00Qh+BE0A25W8VANXXE6h/70nfYuWBIfDmOor8wzvvm5mr3Y+hkkfLn4HupHNzZb4CnyDLqx
0IkF7qjF0ANbYN+5Uv9aO/oda34doV8VLOIZlmC/t70KhiamQyTxp7GzK5fPH+k/dk3wNJ8KpHuV
Kr/gKtgTzVI/Ps+gXM0BjgyxtlvQ6r7mFpbZ6RiVNXJciWGwHwdLHQciFDH/R2Rx8n6fesdpUKOV
0Pwl6oclvC+3sIDhuRKEpmHxZhvgJNwkFNMZt8DBpN/uMkSSMmN0dwqkI9FR6IAYwEubacX6ZiTA
i3wuetubqLnvISlrTwRBXsQiJK7JebsfizH82TvgCRlgXQ6muSIJ68Wr6zP3PP0JYH7Y9wa+Yn2k
kPfOm2ZQDlqPM+LAxu1eHqDf+y8boA6xh/aR8751lmSx+mcw1vMNxDfMzqTHNph5h22weMkNnPap
9ycIs3L7eJynTYdFcBWf8o9mo67Q0RkHQ+5mHuHoVeg+t0Ku2d4gu/Z7l3nNjzp7/rMEQBs7sehY
ZLnVS4mB7E3fx1iykV19ow228y+IsuCPZsAK6B+B99af9CXD/4yaYiVXEjNpdlWXBMvCKgpKJVEW
fbZrpwfotkkqD/IxcGLFupJRzjecXho1smYYXIkf/Ef6sjuwG+luD0odzYJ5I3lJXN74cor4NGAl
5EwpNHeNdjZFtNog9PwZJmLpNXfXBrswkRdWuu10Cp6ab/SYYSDspaAu76j9gKZmvp1VuvF/OACB
eePh3YSuskqeQZjoi5IwPFv8Dkxd64atBENRqkWs1KDpcC2vMEKYzZ7pn4k44W0P8oVyZrjK/v8z
u+tpn/9ecXVDPGbkrCnkt9nuxvMQopzjS7Wffu66MwISER561u0jWpn4G6L7MQJR97mPFCdUzh12
r7aG100RaRtVEGhBENYVIPbeS9HRLag8EaAiDUI+BFIyvLnOys0JshQdbQMawdjcdoqxKKaXw9FN
qrUAnWCVszjQs6h28c94NxIYpE1X1HcVRDtukBc0AAs1lLWN3LRkKyd+R+X2oPn4cWeb7U/0z7El
LoEf+HBC1eWdHicXAAmeJnNpiMU8kX9UQdi/BdSelTZjTWHGdZWJN7PW9z/yHxVdP9mts8o2T9+v
pk5zVwPSmexRqTlmrFN4kZhdjAX4PPSzEsw91aJZHHuIxOkXtLPpJEWbJesG+d7DjQBN2nsM7bNN
SMVj34crzXaPjTbU93asgkfQ90BZ6wHMwLKt4ysXCiTJFUGnmwHcd0CByRwnCNGobVVd7ehySnSd
waVOO5+JauX68oJMb8rwnHesS2q1OENQJsD8C/Y9hNzi4CkqfS/3yX1B6Ia1CGJtxr0Y5jUYq1KE
JA2ZK9JyshSw7Rvz6EbTw1PjupT7wStfzsK22b72Onu1uwIuvaY/tgDVSzCuHXhWXJsbX+A2Hw4y
MBGixnTtrZkwaqi/g/J4vA4qu95dcCWoJGKE9DbsW3rr2/0851LjI+JxSqQwnv2r9QZimL20MLVU
EinCJASsCkJ+s1nocF/cLxoERtB6OFUcwgVL/5jjNuaPgx94vEq3O5xGh4oN9RTGtVSmYOv44RUA
H0fXbmHT6ZHQVGHLSmFDPvM8IcrTnbq5eDGwtu/b89efnJSBwUYUsS7ZcluFKjwJC/fZgIHLx7su
3v6hYLbSBxIu4NsHAn5etx036cSRCFJ4zH+A6Xp68ofjBzB3vYtUJotnz4Xeu9ROP9WP5DfUnV79
1C5LfgOH25BRRNn4SZ8jFftDc69nsgmxYcyZW5OTsWEWAQyWatai5NzolfXosCHo1yGbaKLqAR/M
XFcUhCYEvS/WTrxXfrK45gTg8HXZpLpFPOdZmQYBeBW8B2uX4FfSEKZdDt1OWEm+fMiJZCDxffz3
9kIgjgAQw5dh6ZombtJ1S1lIOnpCjS10X0Z5Ca50o9Dno6JOvRdirIsdr+Wx3ERD39LzaYS+p45N
9dazZO/rcIlN2iU/IWPx3egbxT10OzWyX5Ix2ggSmnwxPGt3+6Qm1HQPgqw0goD9kXx1eAP0AKsh
CI7HFvC6SulDQzrQNTsRsG43auvL2rqQq1mqIY5miyEmIB9nYR30cbE+dx8OKscP0HRq6NDjho8T
q/MaNfyw8vtBNaqQHQf275G8MB/zsVgB4V/ZpkrTgoxaa/7sle5FU/23Nu4jWU8kj2nRDuehV2Xf
Q4+KLCz3hTxzXYvaqLEr4rxHD7PwxJZkHC9LDUi3AP/KUmvPGLC7+hxn9fXsCfHNMJUqXr/8IQpP
BRYWuY7yw3B/Px++CPA/s/AfFW5NyYOnPX81/oaAxmczfc6yhFHCE7Zo/YD08/z45hvA2ZZAUYkS
iglL81AmKqbq5V5drwFyyZdBvM2xjEmNjzB6pV/YZ4FGPGn2qNEk22UauK0pXrJqguKrAueERcS8
NGUswwzH7uLdjjPcNrWAVq1dXOFE4L1b8hLLtEHWmUVHjRE027IRgK0OtgfwhrvWWd1RrdanIzui
5WZa0aGd25SSmlGKR/yJ/nBi2Fs1BBnayYk0f3a1G4gaFo5wFFSzZ6hxaUwt8rYMpmZBJbxZo2t5
iS6RJ5HO6QdHT/w9UnxU6+EEnW3JkY/1mFSkJZuPoOl7z6dZQ8Z2V5/pMsxD+I76VsHMe2EpiMq+
LgWySAFpjFG19R/+qRk3ptHx9hctKj8RdvwPOTND960E8w4dzUMOfwGbm3shRdSYt00SgRJvY524
ngB0gNqhifZBIcS9BB0Yu1wZeZhO4ERw356WT9gv3BuvWeAka0YdjHggBAg5c3IQZAT27zpNHpGt
focUQ0Wg6AoKvHcBVktBUey8PUfuSU3a9SaIouMp65ykXQIIiIoC85MnpDXfxtxmejESLCCU5hHW
NOJcd6ocsM+QBW9GIyo9+Y6ad5yi3Do+4bktEcSqk2YwOWVZxRd46mtNZBMre8B+iFT1yFm511U0
5SE2Rp/VsYnRRECwT4t6lMv/7fjxWjFGjl+MhjZwpdcHa+kXu4r/+1uuQzXZGJC/KILMTc5d2rsx
r2FaoN85OFufR9vf44qMOpdIW3reAL5RMRj5LPUkymkOj8pmrlWI5AEtUf6uzwnhiG3i6jsy24+Y
3NC3AerH8+vrIne0GgVd+JX6SLf07hfNHuBXKdXKMM+n/1EDx5Yd0qZTtW4bYAfk8MOo+T4yu3Pq
BHTC/p1bPj+AmfmFHMrYOiOOIb1wSb1vixdljuPTEER0vlNK9j38gy+AJSSlhBWY4wdl8RHq0g4G
Za8w4b4FchlDcCOXyJ2sF4LPoO05XvjOTu36flt+yygn+hduc6A5M9Q+B24nfmJq7nGUaFF7ibTL
ZLD4nwJtmiNFT8F1+HCQE0CyaDz9B4dxSZ6Tf6D1jLI6Qz/aBiuwcpYisxplWkGSkcmmQijRmfID
MThYkrH7R0JnwlTienScEzLC60tsF/U/KK7O9CGDhmU+V+ZFJAfKcN5XemhKi5GBanp8m7wkoIxh
kOL6EeTx/Qg/DIAR7ERAaQ9vZNcI6QiyWQgbzfLFpbIsBe2fKWWz+kBSG41NdQvEIZwkFEJzCfC1
amXt64Zme7ls9tV6fqZAquLXX0L8uW9YXnqApD/oE4vRL8e+OszEVCrd9Lu/UwWxDs9icZJK/33Q
DBoozkSmSEepfz1p77+hd7Qn0fGIeATamy62PgRbh4Ul8Tb9PikeGNfp6xfngEdlrZv2vj//M0Js
pr6GUqkxuyoQE6Ln/fc1U25ixa+9xAQIV6LKfIq6I6BZNn12V2V7glfsDZFqMDZRn40UqJiN3Fok
yg2NU43I3q79D53PQDAvTrppl6v6gfADzK4kndUblny0r5wOD83wAnp496HAtWQMRvlV4/C3dUaL
rHrK/WidvqJ5e62TWxee+xdtGbQUF3LJcMUZjO/hLKommdlLcGs2KbRlO8e7/4ajiVCXZnmyFc++
CkmAP4d7MTR0NrrXFjkyDxwkFyd5yX9XJfVrtcxxiXLgyV2oycWnl+t1GPJMI6nOcyizU1vOa3Ft
wTgCHbbhjNWmN/HkW9u7Qz6mDHwg5R3Qz1o3IWXw2KDKqW3AlT6QDx7EoWVIZ94m3SPAVQbXreiu
XcGGkBkE+JT03cvMu2P+75NKs6D8YifGZnpRK0jeaKvduWzgWfOgzLUbQrgcOvtbg/6m3mQaD4le
LpPgOzaWbyJGkjd4ONqpbXOs3WfAh7VzUKTdnZHc/lU2Zsd7Tv9e3GrymLHH7R3W2WVLpGUSmXJ0
kCYU8dTUz4dkC9GgbIOWDIJyw91Y4hMMFYYTp5PzwC2pBqT2NdnnK4ifgVpNItb1prP4xzXnIANg
sLn00q3o9wZ5rEq0ksDc1ARmDsJxQuDJYqz0/buCFOo8gv36DyiStMvf2ZcZyv1jOqsWRETS3unb
R3v7RTv+522jDhlAW8afmDXeUR6HQ9unOpLM71ygwPbwl8lIUO2CyzJnpWPNy9/agQg7vy5Ff6Kt
xGfS9NlNOlnkD2KLP1Y7SsOqHPrjNGU5o5B/auVseUFSl4JiBBtc9MNCRjmxDs0JiXGaU0/Sexmr
w7RsuzK28RU4esY54TqpELOsY23I5Ehzn11lKyy3cdwNY4hhruL4ntu5QFefKJnC8oQ4Ks1kHY7l
pSsaRr9K57hRSczAi84JcN9gzmC4Fz68Nkijs9lFC5yLDqmyoo0VBnwy+6uSRSDXXkKQKRkHsjoj
X1VKkFNAEgtFDSW+hxBH5FTJD542MRsHyfm8/2FSxjmpDwhCWmQwGjHXDgFtUzQQDrLNHP334vgh
I7zy+6+2r2rhksf/4/ojHyDWgzVDriSmwRN8Mc7s2Yw6VVB6e415ydgfak6SjvVpMbKY5ruj1n6B
X0jJu17OqeXZuREoUFqnfx1YQpqGmAI43/OS9312OLENsgL26P1aYGkgN8DLs35AAjofG/KQkuVu
Ssizr8qzL4x7ZV/7eomizsZdkXeJ3gCdkwR0Dgq2RxhrJ9c+fgpuAuWNqQbK1MYwqX0a6KLWqVE1
rTqS8lqnrH+M+bENVQt+XEtVf/UiZt8F2c3Pntlg8TMqNbBWE4AL4kuA3XW6PX0H/WDd3eaX6BvH
1WwVA5c8mcUHsJQ/I+x/r1GnJ/7yK6JsP6bbs7FYa4pBJFadyjRsLD+vb4CuUmrr5Fp8LPjqnkDP
P7ifE4D1bYsWMpSfEFWLzPQDk/HWPHrIuHMOJkung5G7iLOYLCnr+/ztTVys8IShniume9zkKisO
pbFTUVeoIZz4fJuIkt2aYA6T0YES0u5VF9upE3yfoXRyC8lLU0+7jcv5i8FTT4BI5c3qplI/iqA7
x8Tqdz8PXGTT1hBa+Vnnk1evGp05Mr6oaHvFcWbEGxwBbF73KA6PCs+C+tSTA5SrPk9P4H6urB3r
ZGlRYj5/OI5TBgjshkmGFQ1FsQqi9C0D/UJOTPgsRFSC2v4ujsLLLC6JouGgE4w9JNvmRKH/4l0u
njWhITfIuKAAJnF1yqG2pgGiRbEGuUIRhT51XuAjTnp+/49/WkfnC7KFjh5GlJVO/OBLzC7kFFHV
g3nTQIAxxJI+EnqPhwIl4Na3kGGgoC+XyRxMAY1hF8m46k19yuTaoKQm5XJLabIRoIj9TFPUYzeW
W/uJxT2EXq5Rn3LO7lOwMop2vl2owGKkNSZIqy3UcsI9a8CUu0p2adg/hGuwDjLwVgis+7Ho9Fr4
fgNf3mPBJaZmsvblCriLr8mkFyV/7MCiQ0sEpL93b7Cuqtk9XisE+6M3uZ/TPPstuZRUih/6qceh
7dB88KQgv82wTLU8RgrjENBRdSjPhw1H5KKSnztsV8lU1BzguFaoAl5QOT+vudHv3M0NXd2BRKvj
dzeJ00/vRj0y/0XEjMDqEUJuq+PX9K64MVfQlisxbFLvIizAhWxTXNzA19IlCsdSj5Ez0cQ42M+5
n0rMgF4iBsuuyEG511NqkoU6bx95IqnPTMbOXrvXwTga+2McAnh0D+ISnKz8hu2mYdgZ9GlvDiep
tru83Knjvs2u+t/GonKuxcgxg2KZoUOytriQDnteVY8RFyVxTaIxfhZMY4FYG+EMnDjzKba/sjGJ
eiYjXkPVfDigasc8QO9CJ3GkzGUTydBup/k724C2s3ABbWcztm01Ndfp5NjOcNTLiAJPBgpWZCjf
Dp8zx0DT8FZA5lrDP8hYUHbJoL/LVnuu15iypN56QHWM5IH6vus8GcsvjdIzgJb7ftGovUtksCPs
4YxNxExIuyoKfNr/kZmXOwjNYizTpPYgrWGr0/XL2fNHyCqTaIfLBFZ8LTZNW6MVrthB28eRWule
chbf8wyxEcEoEy4YFS1BpU9HYwxKpYW5PwOMvC8yuKTiO8fNeSa/CGA5JSE01p+hMxV0lQefe5jv
rVNtVxiqWfDwt6o95Jl+iR/8fpdfMxbuEKm+YnnYN7Zxc0EcKkKlxHawZTBn6raMJDIzgvWcEw+/
tqM3YBlfNAVvNTTQNmNoukfojEfV64tHvRe9tLQ5h67vxeXIUCN6IwGkpBHHBKME1GN+yys3kd1D
6N8GP2/Z6LteFjLTCrstz1uQhaDPAhemtUcMyqCYwOTbNW+lJ+WVRkfmajKSkhhLr1qg8SNUMBCL
cAaRyEjNbnQgmAd6JzDzSmZQ/FoG8qswb5iBDUiEmeF+I3bsIx28N1aURZtroIVSWi4UT93duqpH
dc3rH6h7Y7vhv+rt5hs35ezjUspC1BqmCy/WVzozZEekaVeR4WtQ7jDA34NFti/Z5xTltT4G31LO
aO4Eb76VxylKSl4WATTYXiCVK8vr6KGO9Lb03JWcz4fmaU+NbYhlEG8DFmJ+H5V1Qe2Ys8c63jKg
iMwYlc57cg7X0gQDC5f+VJUwwP5CqKSxBb1Gkr4rPxMb5UakAFM6V8Jj9E9yYkZ22toR3sM+rdSS
gb8fSLt+I2xp3gv0OFcXJjEDK4AZ2ULKHojz+5qPDdqCQwe+8huPLoy7qd04xxNhu2zs4JPha6sg
kL6yrdST0AKmALDjd9yAlldHo7G60D/wpLNByd7uWiKKd/Rlm71FsNCpOVj2KY11PDyblg88ZzEh
cru63C9nXgufRX2lmJr7bbpzG0ApSMauEsbCCpMGDKmEUZGPjR5rreNIzYPY+e1Ez9mYcbFS5gVy
iOV7NhbxZ6hU8RRkS63l8Dfc3nXU8UyRcyHtR6fIg5Erli9ucUmMpA5LXFaa2wjojQ1W8LneSN4J
jFyAF1vdJ9l3EYznDYkmn920bE6Y2wdcTZsKFVeNudA+rf54ZcQUsT0ITKS5qD2oOxwEevDaMsfa
rh8yq7Ev1zNTfe1zLO6vNp9eo/vV6phMYEmVmNRVVTWMNjXtfdafXlZxUbJIIW2pU0GmJX5JIdIy
tPhS62NEaJBoeuYQAVAmL6DjzYRLh8yChFCWZhx4eOxP87NkuIxak2XG4fAu7514QVFsjXVDbXUc
p/e25I4hcHK92nlmiqYAdvpsFzs4UBgUGLVfURO5rC9qt64N9AFA9zU0N6HKpgMEkqTebclrdsg7
mpieVWsVp+P+6lS7y9nZwdWm1lVh5nO1HU+zCWqLyadWFOR5gc5kF92EUqd6dnL3+aKK8EAoRNGO
OvhylRQH9htOgORmGIf+uSQ3zFPe6zCkUa6K5j8tHBor6oNxGRVqaM+D9ZYowkJ//c8RM2ihbKU0
ywAgFBXNKBKRVt+kuFltGszgMmasurK0By9FJ+yVz/Ido2P0CRkg4dyQMOMi7p+HoHqd3GoPZdAm
0eD40RlETLRDHYSyZGJOnkYoGb8yq2Ica0Ks10S/Ni0UkGa9SeqJULl5/eAdHbXL3SYaGuj9aLnX
s0eu4EPEYGpQavRzAOQW9j30jU8rJdjlwJQEQZxAcYHUFNBsUMwwwx8iTHp3aXWlIrY6Nzr9B2NG
ZugM3geD6Zm0Up3JoABTdyNEF6n+Bipcdk73EvfimEtXnfxre0ZTeHsl7AQFtwUk+uqbUkMOvpeQ
eFwTNwF4tlzLcmXK3dPdY0yyKqjgCjD9qqF35Vm5ZAEfMX6+2AywTWzPp9+feo3t/Dc40zg1oMAo
luNm6bddvY9/9rFBQVArqB31OwtOGlpo0kySo65UQ7c+gEvGDv9Dt3ti06cMtRci17o7nl9l7MPF
YyvvvaAKrj/tgZIu78ZRNyAQorsfkSGPGsYVf1NVF6iwQMgn74wi6bhLIJL1uyiYPq001VE4zQCy
q2B2SNo7SMhfKJCAT0VAF41YUwFVZwr/SIey7PXjY8ElS2ziXuNEa86ytrTyI5CYnuZVs9/xtf2b
GIeLq4C4U1y0owSJocXPOZEbM0HHDD6Fw4Jpz7RdxY/cMv+ruqBS/tnKmHR9hCZj9U6mpcUpYrXW
Bf4q1ndI5+0DZTo5gP3R8GxJzujEa9blwtbKjQsIcOmK1oatUjeTulMLEZqHMxn12hr2yi5UAqCP
HvIAuYEEm21vk0KaeqVMyhOsioy+dKQIHkz1QxE4QAWMxXVDJKwSNU0hI6Lyw83p4FkIB2ZJpMgw
CIunl0UdCODcFITUG0iuJ171VVZ0JdXNkCQWld8sENcxryrFWElj1iNLrjlRMrg0V/P8OKHP7Vuc
ZilX80THI3qZmKo72z8Dw1qQ1GT12gBgE6ZZYfe8PpHNXLKqazjBFFutg5GE0Cn3g66tSUZNfkDb
7+FxMLMIq4OwpOyoFCqSXJp5mTuAr4MqThWHAg9iRA1pTWdzCxD2Jhwbem3YWY+Lm+fp6ymfnx/c
7W+5xOCUeuE6ZJ//Jge/oTdqchkpBTlAgwY4CyCWPgRgYX90KgEIN9o+antu0icDeEPHY6ODtjR3
03ixdTMhWd1PJBIessHA/R5ACcjIf5iXgSoIpT9Os9t3R7mlLIshF0ChIOdnZaZEWMIBqmv/l6i7
3da2HmOywEk7mPTyX9Sggk98ggA++9jX2Vm0xr7dxOfXTjvfXZl83dxvBVukGYBwtrdvbU8retSK
ZjM6+z5ejOEAYPwrjS94o0P0fYwo15JfGeZ7keq+K1fP1YFknBR8XHsphS8ToFkdu7b0FUYyKwOz
I1hbP2ecbB5Dd1jTXxkRgntm+XTnP/XJVLJlAsFp38Wus2Uc8XoseAlAzBEaFEODGlKztqrFG9/i
sAY55ip7o5b3HGFfZVXrHTt12xWzrgNskEZPmkeUYgJJbLTxGSqi0XTL7XM2Nq1mac9Gpqnzr23U
xJRoz9DI0n8/LHItmU23MhyVyUMd9sA+8fhCMGjFwnmZ1b2oVNtWjlpH0S54gz9NzB2hKbIbZn/s
M+jc4UGHnjoR/Z1/g3wA5+zZ2n6+C/l33sGwnRFw/b59evoAvh0JKJyJl7SQrRpBFdNwg6Gz8vSn
V0NCgt3rdoLmOb2oqP2KUdTyzUQfLLSmDNPj8FUS3UP159bPt+J5ahVO9PTkLc4CVOqTN05DrGJA
77O/5KzxJh2mLOqc5yZl2KH3O6GE/bjk0OBbaWQ5ocNeGPTPT6fYPFiNbPKAoOsWL+8cyWqCvNtN
/l5LZiOd2oZn2JQw8yA2uhg+gMAsjyliS3DgSk3UARnQbk05xmvmg4Xd4e0+/dhQ0rZlnSR3+jKd
jk1Zi1MOhP0gB9yoMm6fIwymFUXx4WR2K9afBRZ24OEZhedPTaD8/mn3aDdJTqHiO4cxuOoyys2E
xNy2yP6eTmzhFWP9Toph0/2IvP19G0yM045yUIxGP5TwMroAz11IDGfXCwfgwQ2FjqfeC0GF6qwM
aYA7FpeSHtV2/E/nLJx0KSgjWLFSNt1zU8uXHDpPccXM6Wq4mTrXoNu2t3ZlX3rvd06pKzNKUYNB
32Jhp7YPxr7sypGPcqG1JGLKOA7Pg/eyngMZ1Vcpd3Y322eARVvN7GxDa0Ahfm97HQZwl037lXFR
u/QWPczKEP+ZiH9MvOmYMVZVyNlvRBM+cy0Q7Mb2pUEQW4XflmDIQ/0xo6O0qVDkj/teZViaHt7l
IeH6GqWVSsP4L64JYo0Dhk3MK1S/1D6+7P9hAy4qVOBhXS3876+TsPdHpBQshJ6/f4TUJQIebgE1
gmwzCJ0+RufFUZaWzFgiLvyG+pf8fi1vv0ZqCB2bKNcxuZmINRvXRUVACuNj6Neltk/9/1OXsbmQ
0WYOz3CGQJ9pGzlqDy4YOB4AOZ2xVWiO0vckcYW7VhUOwE4+Q8FaPpvrX46QEjpTsN1QEDdsod2P
5mT2nw3FUfqOV61jZhDag0q7qkFWUcY2cua0AXU8a9Xib6RriFZS2SFBMF4hD8CxTK0G26+wel8Q
Yv9vWuIv2nB31V8h8sxEEiRAvEEjKQ1Ow0iQX68nINrmKq1Cts/dzsvGsBxPRyQ4L9BTwDc9XUO3
jsavL0s4rTQUJleLp3P3YnhK1RFTvvfS8gigL9RdTSfSQvt78q3wRh74A2/wG0MAlpHYliBuE4lH
lfeXRwVSGgp7SJqwXqOuQ5fx75UawHBrHdgesIUrM5FnVxi0jEYOVFKN8o1VnS6Mgh29Eac7MJVA
wjaHIuazr5lJyKjFM+Vxt5AsbchVSoqe+wL0fHUZsasSS31hn2wwHODmq0i33tZVP2iafuAKfGIU
XfKiHWyGdVV7yZjkT51FYD173GSiGfhERJBwtlN72aFAeN1HDkA+NvGwKeCrmyFw9d/qUy6wfAsF
1PQFPswcqDiZ8lWSWG4c8q4ELnZAcyvqYnz19WeCl8vpNcJe+TlPiUz0GB9eF1TCMiz4ITKYLWUS
0FC42C9SNAr/pXnvsT+SbYNIM4oDB59Xx+QoOGPvAtJFDoZhxKRd4I0/FtWlWp6+hEYBcejbPpk+
RVH4Do+hwBxwqv5wG3jfwyqNFA4TXf8lGe+wczyEMj++X/ejITmxqNKmqndkAF4IsmqgUk0we1SN
Av9NgHqJ70xUHGFxjiURpYiZ0al0Ug8In/wvyra5N5HLcBVKhlx6ub2c9hsyTF2HpZ8jEhIcoIYr
z2y8Dv2fOU7+MD91q+NKxI+1ZaZhvL1wBwc3U7D7C0WihtS/WwJ2g63ecPyH4uPj05pDmK2XWprB
SREoqlvCkAn50dFEdMqsew6fMw5Uchg5ln+Yc8DoAQvhXJLaAWeA7bba0g8s4V2ayH3hrKwO7ehs
htNxXYUEFRhQXpj4M5O928YzqkLxznILWZn8ahx++QRR5xjn2gGN1iQZA8AeQcivxX6TaTLlqm1s
hzkdUMLhodAAd+/2egqPjPjvugOuWmuzbnaR0sORtpt4+kLEVLLX8Dn7WnEtSLT+HKrtqL2+tsgL
cjeg7BZJ/3hcnOuSSXJ0I+jUseGaSJQ34twiV9m5G2NDKgicUAcdt0X+DxukTNA7FwUpWbFgxpJt
IQCh1ZMhsQTBky25KvyopT4MvjQtotKazrURaPfaBogRPe5FV0wWnlPGOtHtmxKDaIJ4ePH8XS2C
sovWZ6t/vC6AZnz9TEblwW+STmQ6R4XXP4aTW7OcAq6y0HAaWOB4YWIHmKjyRniQ0MeZVKAUVVaw
nq49XhU4Urao8ovPhEg2GzYL7MlXGeWv2MPBetnuv+FK5hR8f4PIDb49tnXtvkxddm6EG68tHmwA
mGcDTpZublNikZE9k/+F5zVs6fn1+sLD6Oj3FTbl2LAwanc9W0/KYSDMYYyNE2jSJUYI1ERf1ncB
3NWLJCMWDDixaFWVIYU6nXDjZ0ASppRJWFNAKbaLH/5o5BWOZNFVbjDY1lfxgAWmGhdGHA92Ksb2
eq1YO2BwvNzyAU2pBXyfn+kqhnxG4cr6yH6HBoMIm41GDli48cc0t4KxjvT18ntse+MA7/Is+nBm
tGT/RTxHZNAIF3824marll2Yu5YL5MiX5skCIDiqNE069+DV18/pbwKbam59RUYP+i3hr3xXlqiW
S+bOknEaSVhHM8Ikjf/0EpOhvbs0FYKSS3LSKwCj8H4ocXcLeWEejf0hOOUlZXUrpWL2MVq4d+kY
0gW3jt88wUME/bBnVyDE7gbv6+DHPvz+QeZkRzZdb/yltt/bPdULnN1lfjm0e6wWm7SjSDj84VrC
0hw/glXeqVhLt7SMOU650On3h3MjBbWHXsnbuJ9eWX5la/QFWbakk1P/wjfoyB3aB1CEERDTSULK
dKkwT+7eO/3HGgcITbU1k7+U9mDnTQaJ5oFl02Yyx2laQKo76VyM30g5YB7MDhD1TtWi6kASGyvU
i1IYgQgDil83sGIpPV/iSxIO5zjk6o6aLfzM64NxgPwHCwTLaudVWiC1TgLMLZrzmWkdvmciM0gZ
Ol9c8yoCN7OZ9E9krJ4X5qQjV/vegi5T5q/mnZpGoa86vYAial4hFS8F6Hsq9Xf4Wyj3He6LQJck
1dUW0ywYeBkmrkmGcShRowb6LbwEXxV2G/PNXvteeAUt37ijvdRhBzc1PswJqIzSwvfVwXUIvwWk
0USwqGT+JWr7NDeI9tJoW9Jnur5+gJNC7oifkVef68Ked0lo/9bDFgHU2Js2mGCk1Cyuc15247Mk
Sc4AhiaR17tfYiTMMO2Ud2XDIP9rHPmbt3PIhTgetbEs7+r4SDoLPc0kw9sT9zLzqjWGhAILJLBz
S2VwkPmI9EUgd2oihCbP+RbBrm7Wa3gw9eRuEP5kH0Qn/XE8uAdg9tl25S1/XLCWtk0UhAvr8D4G
t28f6Nnr43fv/oYPIEn3ehFKgt/Boxkv6oLuALkIdVMuUBbZUlQzlhye1zlLxkqhVYlg/oabddZD
6ntvUbyvtXrm67pKmRZ6HiKBLyivE8BDMHcZciIJ9xvG6uIj6Y4GLRNUQQcfjECDRPrwweAg5nDJ
y82Jd3Qxw90B1Jq16S9cgC32R8rjVhYQCaBM7j0nZavibOFurd4Y9e5zyeibcKRL26DrHGRGWEmK
olPPm2saMrh3LlBm9z2ua1RRaFX5qVQCxVX7dXQp3Jn/+5a4N/ZDOm1Y7VVZ+lJMGiL6LyttiWDv
/XeaPxOaQK9G8lUN0b4FKAFh4N0hYCyUfkTxk61ufNMJZnOMcf4FJlyNbQpNBOfpiAXU4J4FCHDA
DokUOrh21Eajy+pFK2BrrSRAW90fxdiDi7BvdKuJ9Zco56LXdwVE0oQLhzbuD/6ZF+OeH540Zdyd
fJK+pSDKea9qd8IVBl5YsIBUcuZPM8EQcUtlKjBSgtzKUyrV9/tckk//ilUN/1EmMbUILoHf/BKy
718r6vY3e7g4VdSJodNbZtWpgBpEoQrQNUwVYDcyUkziszXouJwaX82CmKh4OdEDUYpmOV8+YNQj
CrC3qKof2CODODEr/9uEXUsr8rJlfPD4TAI3CzzBbJSMwT6Yb+E+I2XJ/OrxTIO/OErRZZaNJt1M
0TO3M7ncJomJbwrDLflpdBFr+RxpgjnJA1qnlD2UN3SRSoSkKeok1u1YEXiXn8mM8oXDriG0QhsA
OzpdDeq1UrE1FIs0Qxs5ckf2CCa0P3nK8i9jp/+9XXqa1ck851ZO6lcEwIkNiaaPt7wAjfQXSyzW
D9t/uj3K8Xf/CMmpDpaVDqOSpjB2jYlYfxTtiOrS1pgXpJ1HBajfMmHpwhsoAPDj/9Fk5GzTH35S
sGROJYkyMjOXY5Hh7VLxfbwaS3vFvEOmgOXMcarRfZ945hSfPa0NVPlSVrZXGrrFiqLcVUrbaon/
DWEflsakwDKIvUmwliscULFYgLqlhm9FSc3HOk3kWYpOnp/LqDYylY5vTI1QJ2DFEPcIDKI9fqw9
ruH+xz5iG9czBp1llCQIMvVMBVyk3eL3QrNMrOATnfJ47JHBUUVgPR3iqYwyr+JKkyCVB8g6bHFE
TPKjeVe5h34t+yfWtc0yCTYnzqKFWN1wF28+Ht+6/ZxrTruYewRF6ePpwgC7nUhhVwvGTWm7qSUO
K69IDuaBaU4kdPB8efcqcBcxMSznuXMD90Rrod2SdT8aUw1yMjTV1qsyIiiBf7OO4yH9uHvFsw9b
pxHURCAMMfGsYhXym4ONMW66vxfitIyJNOxDAUqm4HIYt+WlDvvjO5E3hxCq0ckBPDnV4UvwRjC3
wslDkzSKGrO2q/bDcqyCmIISz/MAqH29szHUlX16aueBoL2T43vQD1Pxsr3CVFu7M5EWAOqaepNz
p822Zln4f7tmBafsuxuAL7w3eTXDIEYHgeJL1Z/agMMdGuqa6TziGlS9fL0ZoH6aS6/9V1A53at1
tdNbb7pnCL0SO4K8vELJhFCNmln0did/oottdjSK0k2Q0BEF5/8il4c2Jests4lKk6a00gYXzVPV
x6qHz8Nqs8guyrgqOHOrKwlxnW4zuJ5vhCu1dt+N8An9Stiy0tm2vmiCymY9mWO7GnA/T2bZ644E
Y3N58VTusmLT380iFbYyOE8Ex9yy22X/OTISwO0eFUkGMjpRFPPGn45I6qhpWtng31y9kHgqk3X0
AANzSC/XkOEka+WV1MZcmVwS+89OF1os4ouGc05g3ygKRQ3a+20ZdLPv5T+OjqjE+vWowvBlU+1s
odqOVdwtLvZ7zCbsP2xdZDM6c2VcJ02rRoM/C/D35JWQZ+A3ofsebXSy5YsrJOMRW3nqNyX6sVwv
FjCPX/oVtNMVZyPREz8OjNqrYuvQHxwOEpZeGDY1X98DaTSXCtM59vBKKVMjR24VWbcHeZ6Z6RRz
Ya7zlTTHjkx3ocHRj5NHDCT4e66l+hIKwy/BQDKMRfUH1R290Gdz+NVN9uznjYmBX9/fGnL85VRO
ebW0yHvdobW9dSgGQcNfr42OYki104CUedM1lKt/NoqFEuyRUTY0JYWel4+ilTbifRIiTHiB8g5C
K3/TkfEqnCw3PRklo5GVd8ErzwNyjZYDmdR5Pq9DK5ZCyzSgSGi0qhwSJLxgRQ80KAZLdr1LZEJY
rzbQxYWN6eqElb2BuPeSDPg4CINEFX/wWqZ05lncFZ1mZNUNbmOJ97PRlEqGdFNjNxYVfvEmEzmQ
FK3krGW8lBVbORhD4zF3/nSctk17v3xK/6NnpO/8O8XYs4cVv3iTMApxLW6LQGd3M2OAXHoaji1g
/8OxXzOV+ux+/K1fqTITWI+WqnCLbv3qS+IzKVeNmjj7k+W3ata+tRmRATE4Lz3OTjSMUyhqiFNj
4W0cHsna3r5bbPVpT3KhOeMnB4ilZzJAmxRUCL1L7BJ3MoBrNt3lIo2D0NHPkFXNDln9S76MwM4w
wY33q8RI9joA4KkH5hkQXKRcXXguP2GZxIJXDJ/y+h8dOm21AxfEzZnvZAVTxpNGZDKkzW9cgs33
F46FslayjZ93Mazz7xtUsCVEG+de94O5lACc+HSJSDJI0XrWxntbrkxpcbPSquPr97LfOozEgUEA
6Lfa+1csIKYa50lzVVfpWAXEaGpz66RlgVmhhUIkibC3YfZcez7m7XdeW0QoDg1HLf4+kXWVpywK
2R6DevnRtZP0Ot80cQgqKVWvsEaUfXeiWJs1951qa4Qy/LkW4lRXxdMRCYi/rxfz9LkWnau+rN0a
WWCgqBVJutswPFYABpPBjadyLM2MN9fZn8kig0MHiK8E7EHI4mtC2Tx4Za07wze3t3NAUBwnf335
XRo3NIWujHJ0e8cAkCWYITGZ1c/A75eoyvXnjyleeevrCJVqMSnisKeMU7nz1SWhxP1swakxAN4J
yf2Dac/uO52qOPZUe6hHBrWndN+s2TNLonK7S3Rta+GJfwm9QQjCPw2Bj3e6dBMAD3Rdd8gf3ugt
DQL0WARNX0fNtD4d51E5/ju3g1wMjQ8Afzd7Gs0Ms9OlyLVlw9oADWqZZnF8qgF8EAPrOTdr+1MR
jJrneLekGTArp80kE7w1K3kaQsc/2vGqdmhS/Y2rqtl1lgz7DFzfWaJ1IcfiMOdrIt0R6r/WzSDX
JH+6wnzAUnNv/1r6LdDEpijGsAeIJIGnfDhbf42FuV2tokI37QrnZYeINY03XLkcpShzwr4Zg5NG
cgjY0+1IbHu8852DjE7ptBMTEm74A4SgkN5hoOf9LD26y21FkG8ImvJEKpNIeKSN8Aed3GwMVmjL
02627M3S0AKlhPD3x3cONpsHj2a6/nfhjpjPOrChpYH4tiqRr1HmZYM0iN/wadbvViTZXTIWDM4f
ixDPv3Xn1ykvIrYYA/ojcjRCdvGFZgg8EOhrst+KVJI0DUeXRZ5PkYQHrs7FIuxZsLqY090Yo7k0
Des6XgvZWTRzdincWC/I70pzaoQvB1rQHKMzmp5S6mJ8mXbo/IigsEB2a6UrfeJt8uC5M3k09QKl
EoJ/GoS7shuXQ5pmWjTyyKTVHEUM4UaeDER6629DqczwJLTEp+wJ6mm29jT2ify/8lylzM9GALw+
jPvmm5VKnrDf4QWfdm4bvplYO1JqrQSnytzvV/lbW/8pGTk38K4ld1k85dEQkrsh1sl93kS2ZOur
b0FmuoT2uoCTyfZjups7CJoeGQ9Qsqs3i5GFUQqqd+QGKLXPuh5aS2Uqpd8W72SRBJ9Y1t9c30nd
r9kCuABeKq9JNXCKnmLCleqib7j3TIGRTvrD9aKhnu9zly6sC7YBrV3n6RxWtE3lRsiCAXihUf3Y
EV8K7kGkg0AX/rLBiylm8LkbcN4oq947oG1mKS9IdjuJKAOOtd0wGSUv4otI5pDz4Tc77EE3pFJx
3ZBRbo+lI8m5lO1YXGzmBjVoNm/P1Q+uCSQJ5f3slWUt5RG6OhWkZekBJDt28wELGJryi28X+Byn
/Zyjv3bJ4gAigx9UzyzIaIwN9m7XgcKBJvvvtqOsp7pAz4wxeuXnDS+VdS/1HdMmwFJsTH4xpkm0
aB4l5uhsdiXGBLnLa0wa18LZX27WqLYcpWr4OslxvqbDKESAGiQEMZvxUIgiU3JoGepHRD/zVVKw
vS7n1TQ+XuFlXnz4pOBam1aSsWxrJFFNr9e1nlrM+d5bNDGPwtVd2QNUp2J5ntZm0nq3T/5+t1KT
+YGuiELnuBHCTH0RXriLEoQY3CJHo4L0uzRIC1/aEes72du3yhiCHLhmwBL3cd3SWK9ZvWlakOOV
l927wPBCjTRWKy5iaAFsElCzvlPGHyAAnqD47TcUJpQTmG+94u6AezpnPe5zUCyF23jh/FfJSOfN
UmEeHWSGVX9pfroLrWtVsrZZW1IABPDG3HkzR8Fe60IlyFYVLorgr9u+bGnXnq6VQvNW+eCQIdt2
bFbvH9Mko4qaJl4h8DqI+7ndqTmgmaoFJfk0wt/ViQCNsOLzXA5Wm59mlOLUGqWs2rn61h2/O4Fu
Z4jMNqGRQ+mFufCIvPUYSo31L/ZOkz8V4gsPkR4J4bQiVzmSZvYDyXqIeQfqsUi+7hwIKBS0IOEN
0flYybjIlrTuGivlqFXeBah3YDGUvprGj/AsgCtUlkLhhtIdRssNg7Ir1AvN8jN5+M39J+9nEB9U
JfNrJvMbBxgo9+x64rm79ELHC23s2pOiIep7YoL0n6+DxyDpuuEc+beA2/5Q5NY7CVw5XEqzhuLM
awFWGuMbkimoFWOkQTeRE2PJbSArZ1dpibZJqropZC7jlaSTNW6gB9FHnfDUQvfrYxJBfEq/Dt4B
vWqwgEZELUMzN1L8MZdcwa/gxNMgOjYBtD0uf6go9bmg6wue996qmH6F2ddF2bboIZAXKexmDZLs
j2kPqp7zCv5RlGayLnTXhFjz+ARrYHk8V7muBOlEdQ+F4xSzjHqQyDILY3L1B3PAy06WPfSZbwIB
HRB+7Z+vN5/tPAzXI6CZ+SBOTKEpemUuGn9yujAOY4ZZiDRe7q1px/U04upmYCm7+wDDIw4xSOLC
kj8ApunrSMrAizG9jDM0y6TgG8GF9J6YrLmIz1x7VaTqj6+epg4beLaTOBHORWJOyRZ8pSU2BOYX
xSaA+P71CIBYe+UhDG+jqykvRx737s14EoSicmLcqiIlHuWWkmY2qC3QMQWGaqIOsLbKRxD869LW
N16svpbcWE43MWCxXMEBhlPoTrMBgwock2IwKV9UqX4O65HyY+KD6jfGhyxxed5j035yw2mKtc3h
VlDJgWa1wTn4Aj6hQOvAvmqtJH0XkUDCssqsY0ID2YCbxiC48xqF9FztvXRNj6AtGzTDGuqpj70F
wDFWE4RU8oDLn2WxJPDZMYvRGFJu26Nv3o64or3CfNS6j/eI3rq1DyRG0iJabi1Jrsmt6rkHkoQx
dWMPIo6GTvcuyz8wWHLD3h/L47ghddiYvIgs6dv4CiocHb5M2guCD75yMJLRykiWsEj6oAm4DXKq
SH3rrc4gEEWm8icvsoPDQtgeHPoRLc4W+jSrF1ov9dI5eWqiO0FgIy5XBHRbjiofExN/TW3xfqsD
fYdRyt6lcQDqaBVXxguPjWkhKuNtMaI+qDMcCVKBibdqOcwK/p6OlnF+5j9so6LBbd8kJ5xUHrNX
De0gHEnUHFY3A4pq8E6V4GOP73OGhfbN37MorNhn+KNsdvBDkpf8HdFl9x2dr8Lk8kEC8tQVGdDn
RK3Z6RpWhEV+qu0M/p9+IafYlhTdNwfCAFfdl4NtZlUnYCGFHYtFMXJW0OvlsZZr/xTXFXtkv41D
ha9ootTEzy6ETtUK3duOXb+fjKLwo/J/gBLOsVLnqSnbbNC9UT2MxsypwX5Zk+p5SFiaFfrrXsBF
pV3VeTmNfwEzXEPqAfYSm2zMI3eDowFhobFNCoh7rYXhcSi7IcM9Js4PkRHM0ULGeWZWbmIKZdxA
+6ZeWKIAtn689D6mobLUiLlqdz8bZ8listXIwA4H9f/StT/gE/usLeUx5tZ/65SaYK9Icmo7Vl1N
amEU/22PZqO1FODGHp3LCMb+NIy9FXFAYtIEDgsmvM3g6jlpz1jONfUAepy9jtcunOMCfwicSIVy
tujlMaBhQJXz4yIWxCc1Zju45bBS/3Vdsu9eLkTqLFe/gx+b5UHHp3a3BTTPNnkp1XBmShTX0iTR
CFvMOQtrSAuai9SG0i6AcfHtmrSh7VKGtxXzOCxznCCCUEPhLWtNnln4pOTdl9s6rHNQFJlsoIGu
GAdSXFQRk9ATb70pA5hgmVFSSw7olwLDo3DbTv2jleh0qFX1XJiGPCwsDxXMLYyUP4ygGKG0f5gn
s5j9bqAlrrrmGshTNEf7eGUKjKXO5+L9CBHHilPvsfsOYtGih5Firdoev8OUv5CHXfFSA+8a1QQQ
tWqstTpbt4f6TfgWsDtMoPacoZB750IUE3ym38F4WD+6U5rIafQfz1sFso967lpSccDAWc0HCB2k
L3br4N6e4GmTUEyVVO+FCu9JInkr9IFMVYHWMwoq5clxy9Ed9xvAWrU2Gs4tzQMqvrdsfiUHQWPv
q0//GfNnhVOP/1DnsUuGLLyMtGLxZNW6oosYTM9Ts+ysImvtugQRUn0digyhWReOSbflr/7lFoKz
nITJpDVDY5mSuR1beXhTPsOzf6yMxtD2KmnE3ePvmpfecXX9lCbdBvI7jVJiGysxDWQ+iCaIBmF0
ysJU26sQfzhPjJAjw0f7uDEBYRSrR5LuqHiXvWTU0PQ+Ug9WvJSvp9viD59WP4p8DvsHrF2yjWT/
mo/iOCTj1T9gfTb+g06pXsrDuRF9JT19uQLEoLrpsIFAaUlKZzAiQS+r9qNxloT5i2y0/4IgFvZq
jri6HvanV8FOp6T7zrKV7Or3EoUmRKMv4T8T+pj8a79MI+6K2tpfS53rfiVNG00RkYyHzWnI3Uti
AqMBNqeMvWw+Bw9Leoq05itFoGJi/dojh5d2TnTLjpvZemynlP5IPyQcTmrhE0ws7TCDa63Ftowl
2qtoohHMdBzy+CZjPMKFLYoRs1rTSaeCaBOcJRYLanpQ6LD8smxUv4uz9MI6YIyLYPlmFhUF2a3a
/mryiwnGEVmfLc2isqrhb//ZmjwYYu5UoicPb+quwvyAVAh6hv2zFvjOczHg5Qzny+Jc1vdRqBoQ
MWbrjghplIDn0JEkfyBdhtTB8FX0kHLXDgRNeRf5mHunmzvi1ffzrfpI4ui6EXm+kborEQ2tWNKQ
xVFn7gqmS7Rd2q228t9dd4k5yRcdPTvjz1i9pLNJ2y1PDF5mPA00UfM3ZqmPDBINXLhMEuwoQY8A
G8adQhg0LSsmUuidgrp63Q+6OkLSL/3GkzSymGhbf2ROzI2E2z/y+YcM9o0tTLwgS4KdcrGxLQtK
mvBuKbws2EjXC6bVIV5+l6ngHe9kmPqo9u+UryrgdSlJAKdgEJC5Ab+aFsRLox4LhDc88i60ZnaT
TG51VXBLE1F/pUB4VupHL5pi+ZVcBhsG4cqyUn8F+HCuKodY+IrD7iyvArRInxmMdjzgaJ3pLGVi
mm6zUypYhixMp9Fmi3ikCl6JMDSPmXj1pko/OV+Q/2C+R5RsDrNyiflGgHMSTfFg9jF1vUrFzfQB
DQgxgDl7QXeO26n5XH1mPPGW+rkOOsLykCQWDKjmj96kg86sxnnV7EYqIVRcNalUrzlzn6OoPAq+
LLQSdoJHzUIZenZBoybJVbYQna92SkjgTXPRjex75yVo9zsM6akgAbjq7lKWGkJ08UgaXhw1iqRN
/xL9bw+eNds84ADMD/DlyKu/M3pUBiZVlHPndKyw54cmSESmq2Q12MQgyPtJ7w5RDQ7thTe0/4CF
oYizM4VlRvgv3SFbOxyZOuPBBNx+RPj4lNVGT35q02elc1HxQxC2Rf7yS021mjogXfO8lrFBA1s/
BQ4pqD0V1vbw33ursa880Wa3cCLcVY4tfyPLADvtjxsLnFc1QYMWR4mOF42JTkXO7KJWsAXAx9NO
Ee94MViN6a+H0ZuV29Uj9QujLkQJsj4PtK7bufqtqITMTSJYUnaN5MAxJ6TL5v4mJGfFzp+Vtqac
GGgAbwpQw5W0xHVJ4TTVKf8ZxhnHyfW5UdzMi/cSiuqVuLOrwyG57L1FbcEp1tlt2XbJtyv4Ynw/
QdJpG9tfCP0v0JOxMvtvwLBxOewZHzCM7HDYc5+YsLbrmuYoQ4HMocTaMBqjZ6EIW6HyYwgwHbAF
D7EvbFHBey8+drnnsYFM2wF4c9WaRhdktciRqyzd22rA02BttmTT5nbGATDbVRHOlG/B/gdKHQmB
nc5kG+cnDGzSRC0EmevLy9bxHUXKjkAzVMhRgx8f2NhxLAsxvs2R8wrGxNImyjLihzUPKHd+wClY
yZGmoPOG2gxboWLFOFzohePnL4HEW3zmWy97u27xV5m2H4vQyER5xlPUsctylM/nXhpuNc/5G1Zm
ZL1YLB09QkMqxXvZ5UCIsWFYXtsO3+mVEh8rNfCtyTQ6wHTww9WyfvJSMv3cnXJXJRF8SQA9EzQ8
iDiocB213zgbpKwXaHlFGznKueRxjcAUifI1fl8JvWkAvpxiBS12U10uHKelrXuXDSEA7LGhPCY7
HqyldDEgMSfJrZhjK1BC6JBEoEtOIRZQf+g0ou2NfVZjMhf+3tRzh7xFhrU2Mp9jA7U8GwBOj4YE
ldkBqnUWyLGq7S1DCF0hOHdkkJFhe3lV5VpgjNxPVUFa2muLfZkBubUctED3btOPHK9siZjvYwSY
C3pIPgBzRh58ERbEdpzMpOtvJulm6DK/RY0ZfkueGM7R1Vr1+xew8mwU+Gdcu7ubGCfGBH5BgI98
9CRmJ2+GLhF6YzPDjRrmb/USdz+oo0r7PylTjTU9o4ytyoE44ibMulnNax9MOgmpy5ykZRHv6fp9
FThJILd4TGiUSVVsRSM3neg4We5SSHmA2xVVUYT9lbbXoVrRNe7d6sHrdJr+t18ZCrfuRKdOn+Ja
CXEXKlaIy6ex3eYbvsVzc3gpZWCdz0EkDki4OPZQk7IG7eujU/nV2kwg+6M4eIavmBLTE25e41NA
k+M6ve2iEyPOOU4lnKaLLKskSa43z3LH7SYQ7MkuB81s0MI0o9OPrMqTZuTzKpwnaZZ58qmHSrbs
4oaX2vvIaRzACSmtVKMwmU8HjIitiFomboxE3J5E2P0zKyGsgVySH9dsA7e5Jem3kaB1PFjKnZIO
olPxWVyKtLCPxspQjikZRYwKV83hKivCX2HSj+jxjMTkUnpSBQbRDzdKVs1pB5DKWP5PPBpSqYPo
32YBFiKay/NhJclHRWxyebwOdFvEBh0EP/ZJ9jD+2W+9MfArumh2Rcjn571O74wHWghL1AkGPhsj
lhhI7rq0gGongTwA4WNX7ytgpx1sUxYZVgKox/WlsJmIRSwN7uJ28AuLP4a0+I4E5KkrkWTlFtUc
o5OR6yWsVki8GI1Byabyx3t6IdkrTJJD4zpigbkPrk29FL6Gpzzn2/0Ws5uKM5fIcJfmw4izNLpW
4WZmCDD+eHh/OpwUo66eaboS3SJWg3TUeBeQWxj+xHU0lmy7rKjaqM6+p44brj2pJ68HSys+PaP/
Y/7hVfSZNoVMjI2P8Yik/AidTAWRwmBSKr+QB6N98J143Up9jFjX47zHaNQyWLTejpzxfCHN00sd
6yhgvmeF9KSKvRvPCBlZNSPOjrxB6MvrSrt0VdQVNvPovkYuePmlHPpoN/RK1t4ih7lWltMlPa6c
ZY4W/lKCvy9hRyJ/F8cYNMgexJVl4kZxEsNlpdgM1Stro6qsPamWwKgiK9aRIoSTx0/Gq+GLwsCb
e5Ba0HkiM1u9QGXMyhCIPqSNh2z7fOw66jPwrSRQDw9sNoOHixwPj9u5GAqFIC9JLLLrkSGQwl7E
LBrbmL4JS27lrvaq4mER9yAVlWDyDKf7skowyusbranfMh7mXJ2nZmU0oB7ilg2Y0fdvPxeSrmIn
K7INvq0rTcZfZu8WxGQsCPWm1ZcYYo2VxaWO9BXYkrj45kskqj/+ygeLsci/DNoJmE+8t9SZ9b3s
6uBNdmwoSdR0FgjmWoqSjovghDKtWOAeNClIavoYrgazUYh5wMhmxwY1XKlknSlx0G/VrswaTP3X
6x+wBXxRmQxjhhULDYqZ5vqdWndXSFP8QjxZkyhUwgIuam8RAhIU/nExz/Bs205hBKji52bFOhle
b3gf+8FK/cHdsRwDxd2ggmpPnnp9dfcEkQLP175OrtMCh40UdlkyfIN1PGvGOg+sdtlytzvyU94U
5icedHflLtlNncIMNa/r0KahtMC7Rqped3zJ1fC90p12YXkJxwxoTYnHGekJ/jE9YvtwL8u7a6Zq
zXBfPJ0wkg2ToucWU6s+ciVz1K+5fZYcfvdEcwXC/5nQ3ix6p/FKruUP3j9LPHygDwDM5jmB2y1E
b9LGGBgka2TtDtTQwyTJSwJVgR5gPha1tfuthEpbQGedGNSn3j32DvthP2OAON2jbzUpdAPI8Pbq
Ygz1w1cHEZYa43KD37ZRyfWP00fGjXfHvx86hfBmNDWvaY4qcrgyasZhiDkXs1sfOHcSX8OeVqel
vjSFd/PZp2mOIG/1JV7zXLf7wyXEWwTDo5Hef8QrZJfqjBt77VeiTEbe3A8Ho2meJHGUHXYDRedc
zlwLZfqQASmqVdUic/wWTFlNr7WWpvoFALAvDsL0L/VfTYXjWc28D9xsGJ+VKlOwWCeSg96kk5gZ
O7jOBBrgcRRU3xQQognLwhv3yqqV3CM/d3/j9oc6jrjI4v+MlJr8iFDOexu0SzoMvX+OV871Y2K6
mdnqpYydnbvMcsKqVyyYJ52Ky2Z9E2QAe3rqRrAXZigY8NK1/bYGpGMO65tN9jj70MFlL6PEEv6k
1YsiwEy2UFEKrqj25aZz8Nh5ixYLvknaC4/UgLHIe9Fwdb6GbqtifztbEKegQAGCqGvOU/cnrfog
G0PC2EQ1DYvbcUSu5jYIK8VjLhFfY4Qu84tW3nTaTofyjZZUQFXTOCtomkL+LSbYmoJ6t7k63Y/F
rgOvegQKq8QGC7EwM+nix2GMT7BhmvEeKGMw7492Udv6FIn89kW90ColP9q/bIrMQzdf2fFSgJ5l
KqedKmssGwLjFWUr/KqOE9X6SWbxtu9/LMOG0WcA8ub7xSKRD4aqScCSRIMVTz4YX+loXs2Zq3zN
88RixXUN+5Vd9/ewswxSXs72FYU85nu39Q0GaWAbqiTQ5wbljhNkgczGFFSfjrZTCcv45ZdJnqiq
nUR+QfGMkdbdGcMmVlRLD3ad3xdFI0GL/IyMR7/HRw5uJxuSXdaMW2FtsK+UVf/ow6xJXnssKUKs
QSCBDpeaTpUVY1G1H3Xe5KOEZJtqgNjb9XWKHtgMmMya3XMfJMQD+e2O6YbBxCZiD8p0WA4T3Vna
dKJY96RxoiPXU/KY/Od5FpI/3c9/irWKbsvNZJQ9sI19lDemQx+wRntmjXCAg+csTnjWMacgbUlN
hB7yELz1BFWVX9iqYkqbPgHBoBATPvt4nVC7BH+Dc6/PiWXbhCvSRoOuIK+9tpIw+Kd6pvgQOGnA
WUZ3dkvwmeTMBWY9duY/SpZH4OSyMcU8hQe/+x1YoVhi825AG+Dvfy6ELaHJrlukbBUQZ30jyG7r
wjpHTRNSBVOlnih4BfCC/YxTK096ABOmcwalTUg60RwSe2ep+Dyhn1gAYoq37XP+7rijQ8V2YgTU
PLXjIvCTWoe3OqRJowLcP6fa7w/JdV5QtPiwN7kAuk13XRbytWjXjy2yK3iNy6P3SHfaPhyPI4oM
EDItJGqgWiqgfi1Egde9xsI9lLbz6jTs2aK7IES6VdpoDtfqDhCQTj1ggYbHUzf4Df0/WFyODbQ7
SrycIwIAo8ftz38H4zniFnU7SB0X9EnyzhHQkVZSzqKkKT4F/4rr/cFWyXB3J/yalU/xMIbMmcnY
z03RPD5Uj1rCC0jXs/AXE6nFWnupMfvyO/pOhhSDtc/sGUjubBeJ5Xdqbw7RPEkCCO7jX7DZwjrJ
RVvyy7N3EHRfHzVXbgZbD5eowZk70c17Zp2Vqdc6i/f6FGs1ISnHcumPtko38Vug5301VSd2iR2J
UmuExRaI4Tkp4hKZHfMMKbDT2H3VfNvfjAcyEp41YAruTE8faFWTRL3c509WL4YqGy0ygcAqcnZV
J6SrO9wBMMdd6/jvVFqxoTbBPjG7H8HlT+JbxcFRfg8bM1qvJo5YFzT5Uhy4qlC9UnxO7ZVCDzrU
V5xNfy3i+Zrf+JGIm8gXwh4UipAZQESyxUwnuBXjkla/k9qCUKXPGmLhJQVsN79Mh61gUkp1pzWV
FwAxIWnXeeycxjFjaagH15LGmWpLMBlgEk+j1t8zEaXA7Cm+MjKe4ZQefoW7oY7O445UcAUcSD2U
dhvRE8TD4M4Kp/Hw+AMfgX5vLmmFzUTEMw3Ws9QRqfAwpb4iiYfX9YZFJu5eI3KUD5hSapV9g7HC
z5bmCpKIoW895dYPqB7GvkpJ17yw0difEbF4P2mGWNbq8tlMOw6Gh1P6vzTnF4VBppc/PVLLKfrh
qUKybVx3fQcinLngVMmxBQVJsUiJt2WkiJkqfwhJ1t9JR0iOE1ln+Bie3SmD9+wumNgyB8R5jXig
SKOcVAnRxn7eqjetbpTiKR5xghf4pnemhnA5Ul761BjpRyQTlQI5mYJNdNRxKmOgUaOqicP/o+bs
LVzh2uJfHzgRhasDoOb/j3NzFQq3DdGvZVDkxGwV+A0hAxnYNRpdpsRuwL4bl7jpTzck4xyg4WrQ
O6vn/3qg/ZmYfGiXFIsxALsu9Xl3dYl9ip2lautVT08A4W1ULygFqHJ66xbVKfROC53d06131/zp
u37Yyk1n22uUGPNHvsuvnJaOKLVELiQAr8c5Lkp8qRkOuUy1j3s8PFguW6Ah4Dxyuy3gGjPUYKIh
jN/LVZynke8k2M8Xr5555qYbir3yUCgn8rwObGmgTBDkbNK9kxfgNElqm0xogosQyPuA66uB9SBM
TwTcyTuhUYjDqJFLoMsJveJYnVwidhECyY1cati8UYa6ZaO6yyNwpd7usvC8rN//SZ44BeqRnfq4
7KLh2eif6KowZASnalMpJ91tsNdqN2UB6OTHbELVkQwNst6HkP1lshQOJG+ohvSE1a16egNkIFZa
dTczDWCjGUcLVG1l+qzhTzW5dJMNBDMFZR5NBGkvpsH0yoDfvfY1bUddMmnln4yzAu0ajloEenxX
iu9EFgeEI/WYzda+amcnSEwwXcYJMox0V0nAp8UuVm4nQlQJQyKFzpxWKJUOQ+sKj6N/rbBRXQRn
/pL/QNf1HYyQGEWfeeSXsNlsyphjNdc4grIa9FhaYwGPM8g4gmPneDGT3+ldTwDK5dG0SLuaogpW
qf4MNE0CkFaEk/w2I4o/VBega4muWoD+/yyofIN9geJE79Ggof3GDvcgMIuPMLfHOxzGDeL6G7fs
jvVTOmuGqhtZDTOgz9jgSIDUnpBa9yVABr8hbhGErhzYuCVthBcg1V9Pff7xWjKTiMajJZucEklE
NI2dm2tVpT2wTEsElJSGxJqoJBscb0h4Lrk73ecqGr0zwSDaTW2KXIQQctUEe1hdGsnU7Qsg+mu1
G25KFAZ/QRsSSEywg62Cf97AF4T/ogSeAlRQJrCuZit/gMcG9vQ2F5amyDN3uDNdZVnjGSS2YlEK
+5DbXGinqFFejdnpozFmIr1vseIW4OZxnUDayAnZOco9v5/9J4w/HjYccKVlESj6TfXSkqNolFqZ
rd5NDdWd5a7SVCPMicGlCqBHLb9FixlfCy82Cm2ZUTBLK7zQCubVAmJI7ahO0OROZ26zIcs9p6K+
0oPUitPl3Nw8WFA1tzlkH2oiKYWk9s3HhjGJP0YBvA1xpy9BShL8jIjSSvN/B9leXc5jH7ti/haL
EAsj0xXyWBYhjla+jqbuzsY6lzRx9J3lOtpokGfku3fn9PCQp6JWKduoQCh7KIi5OA2tLiAZ/J2Y
6mpK3p6kVcuO5Pdv+PmB75iJzWdu9ugKy4eE+t0L7+vyB3a2NS1SAFR87yV6i5DSeBBj8AHKiWVX
WL/MOgeMYFG6mqlfD+cobqkEdrn40H+P9YiHi2vjK2r4OfkiiCNuSZxL8M32B5oUVKfwjnotB12Z
tzWV9eyapVmNmp9x8GhDZa8WLkk975OV4DYofZnbxK1LdAwveqqYS9/9Q+OweqiPhdxc/j829rGV
l//4L5NNgolQ3WSqXGhFccEaVdv4EvONEYlN174HTIEHBEKBIn7WcnDpzL6HC5NEZWRuJaZCrfVJ
wZEpQnUTO72u2k3chwlMaV2P3TQb4LW3H+LcJ8LmiYSJGTccS95ian7TH0bmO+lm0ANdh6He1tXq
fMEB7dZNEmtGE/C0vDqkzWWwYjavd/BC8KUIW3WbOw+L0vMINXVnZGJHYIIFOXHhxJYEHonhQIhi
oLgZgkjP4vtARU0Kl+q82oLQi9X5R7OfBO7POxGLRzPbem4OY8ozagULasu+b5sHSyEfC1uzF/s0
FUZE0yZGvNRqezUqhHBD9qqpch/SC35+GpVSA/zXK24wBQzXeFUzS6AwPKz552aM3jNCAkpgHapR
8Mg9RHyeqc4cKJnLNMpox0GE7oNgp+6pcQG2qaXtEmwcKW8HNYAm9wZbH+kCv6qd49mWVRHiAS8m
82VhQBWIq4sUxZByfBMSZloUEC4aHX693dTf03ChhGhLLr2v26v26dmcUTyFVH9kWzPltK9KyKCx
k7Ao+dPoSLZJlMEVtfHLXIg/NA8wKmBcpljwew5w1+2OeFXDieacIA/hlZtfhl5y+k3nA7H54bxm
I+P/sAkjA/8iMn7T3tNE4L3whZOUK0syXSVYWwc1UidlxRu3ifB/CQRozP6WExrDS288KWwgEn4r
mUp147muZrfxjnSuFbH1n4XhxSz3o67+VzZBsYRUrPXUEl2LcEc5nJodb7+8BHfYIeRycWfZ5Ckc
3ywQELMDx7XvQJqwlh38MeEfqJT4EVr3RY618OD7NiVVrCDbWjII2aAgMw1Ow6TlB6YkAzGx2ASr
PZFtoer6QsMTJGD7BQQsX3iC1tUjWRL4T79Cup2lh9XCpMiBd6uKWREeIIKlbMrGGlfiwhqmnDgB
gfdN60mJ0cT09U+xxcgaXXyKtRv2JW60GIoySJkoNkl+mYlt9mSO2mH2HbnPzALVeQjOCKI9OjXY
xZvEOCz6iJ6VBbXhqBGnMBuCowxhjWSZg97CiicY3/yIOZbdicq5MMPepNQlCbEma8fVxpnBrOJi
amlEEdh0fyJ21zVd/fWwlfE7BB15xq4/ud97WPnl7hOdzT74zp/sZp3EfCI677PPsPkOCx/SdYue
UDaAv10CIWJoANNgDlGkCJzplvY1TK0mKu+ojGNkvjTT7fBWi64pbQvvEFexo7Wosop2knInD6hj
6d+835lRZqNZZICPqll/HaYMULO32W3Gk/7mLFdf7bWVQrZRoI+fXjneyZ1Wwxo4k+FWZ5I6RIEK
7zlVv8vF9bry56eOHyt/IyE+Nc0oJs5GnMG+DTzoeFFtl8TUOYFXvYDe5vEwNQAuP5SJCI8HkhKk
jU17FM2vAZhiPkDtJVZemWbkdL6d1k6zpE6K+34chDJ6SabuzS/5tUcOvlnkzJVZEoiz529GPIcM
o7Pg9XCmFGvu1hNTGr5IjW++zMNAp3q91S58X/BioKu2wnPaFM/D3w4jeSbIjFxWBblZwKTZBclF
uvV+Csp2PPguzmu+hnbYQJbA9rHx0mTU3mNkgkl7RvX6fUqCOLyoKv8Q4Jscc27CPnni4LluCg7e
1mvNJtRVrOFaBIS6nfwSy/VoB7Oft95m0kp5tgaliBNWAEGhQ332zoRVdczAHLU/2/dODgv3A1H/
slN6nuNtr+9sgFj+XYLlsFlJuqjYm3/HGVGMHvvXZwQ9CdA/X3ZTXGbxhL+H84HJQ4iK2eQtLRcI
OpY11gOdXHoeGvG0+QlN1qy2ds7FIJReXVvPtO+GVQJAJgwYpYI5aAlZxtNckVrIYmXzb0BikCPk
HKqJyKfGe4K7NQDyLggux97dQbkbOzJkSmiubF+XQpujv07mZivT+gJzkgJCilNbEvWqN8ruaElv
JnvyWr4qitVhfwFmZiae+vJSzJAtCGg4ahPFxj8tJDsTP/hgCkSLvn1C/MldObv6479zHd5qstvF
OCnuBvx4xPsylzhv1df8bLD0sRV/ZOcVhXAO+S374rzh5efSo4iqB7GIdY9Pr6NGYTmK35XV4sjx
8KZ4IiJ4Kkn3QjMCHyRG6s0rEJPwG5LzTFzgiuNW6TlPpxY/EsxQwEQEhRS6LIIKBjXhrnR3634U
225tp3nfuSi78ryjd1HVIlPaOSD6oFhbGRh2Ov4Ek05o+56cZnotxU61GJsB+oNJOAka+m0z/oNm
QQ7wC62ys/mQzfzx2TgtbweltvS6HKFfOTiD2OVFRUi2+oj2GHMYztWd9r19a+CEw5+14nPpZs3u
EQNrPLNUXHHjXDG61/hkNjvO1/Cpx5yxw6glhWMVGdXYnGxfoVrCGKZtTgyU7f7RazaUa3Xopiqz
gLo9eQhBElZIwBiBFkYj06cd9M0lECUSqS3QAUk+GCHDBfO0dwx2a0uaBYm3cBxsgPf5GoLQq82Z
s1aukZVnzhsv/svmG1XrNgV9kqBu+ueaVsL2b40vvoVouuJSgfI1n4+icL6LUj1micrfoXAfIkN1
34sacQSJXAY3qpii3mMAYqLENo474fE/mXQW4CkisjiZMb06BHIsLqunazgscWntcnNl5mH9m1Ie
QEOOej+e9SH638TmXJ2KUojVWi3XE8qhB1eR1pWdiOQCb5t6Z9cDK9p3bOode2wjRaaOhFok1YrP
0XJJZZLkMRh/YGshEo0hSQjI7e5imcbljFVfHN36syZa+VjFUNvBc4nFfIQVAu1ualqWMwdcvJlK
GViYD1LFH1nz/b3b3s9gJDq0kI6Wb1RUoNFhgLXuXhk2rdU64FCa7Ng+TTwYJ8P4kwKHNfIbHCL3
tu3HP6aRtd6oYKSr9nglp9fSxBv/fvd+Q72fVtpq64nMWFetUc4/khZqE5PcLlfnn7CqXclclDum
yNIoWcOuWocWV8ZdeuD55Q2Eu2BHFdMwil0C32MpiIiwm/C8FzQvVqzvcgqgNsIIvz1c2291JeeJ
QxAJnELWJ9U418huZkIwHbEQ0O13iSZZ1Pp5KmCRjSxdEOYbFmR0lbNaASnYGGaIV4WAfUaHFcAa
6YJBEYzXT1p+OJw17BcH6uZvDWJNGpff5P4Ke0TeIhSbTq+9QeixUtTz4jmjKoeOTwNgeJPSiXUs
2RHWXj+bpi4J6bpi3C1dz9/kENLaAAXZLqvHA8NnalwO7v4fmhCzOOkOIa05ic1E4QVtQIX6zUBR
9OMldi6LPVVMcfx1oUOXeqUKPSCn50V4uBZQHg4855FheaU9Hm7sGupLkA43vVkIjth5GoddLcPi
BTYBESSmNyK7UfoVoNdu72yXgHN+vY2Fyksrd7EJ8LpvpprZtFTRDKN9q+TpSOOvpVGKfhy8M4G9
UCP435z8Lg72kR8m5+KrXAByeqA7ZqH/BiqEig1OnlWOHmLcKFZos1r1CkT6dnKd1Syl7RqvTAp6
0TAshqYMqiVkBVt4ZbrwPKwrBZS3mBarsZFP73e+S4g1QPH4dVkauCfXHhYCOLdQRyN4r0oFppRE
7eaifzziJnE5ZkNlZGp1O1tjwp+c+4vrM+k+3oajkvlhxA/jDLPZ1Ih2Hg8CrlkrgvPOCQoUU4Fc
ttcROcSebca5GQLjCfXhLcgvs1wIP5Rctf1A5og25sJfvsvzBOk4huqSjhQ/q1vHaTbS1UfTkaQm
M7czQCgk1z34FtVrgl7sG3n2M2FOiifJV81zownPd+aaQIHlDn1h4zz+2rpfNyRHxMmuquun1qY7
FHuVZosSJdMjUfshjs67taGTr0JzTs3yV8cIaALhTI7mGbeeY83VV+S2y/u4RcyZS98PkpgMVdrk
q6n79aBFnzLKr0197mRb+Iupfv4x7YVvRF6lAMpAshZsMsxTYYW4HXKRb2OzeRKq3AQQYZhAXU5n
eDEwAPPfYzdk5G7Q43NuuNnxXZPXR84cNTXR+9oKi07fgd9iWZ5c5KAUNUClhhpMk7E2KLZ8Bb+5
Ba724x5Yd1tuzT4kc2v2InRLUahLSqLcUh9dkuOtP3Qx99me0WuqQ7Ki9/NIbK+/4y32s2iM3R6d
Wg0No2MSDTKUA0FJdQivkwH1E9ZfXk/4U94BA4Eq4X0PRBqhsRdTq9FFFWHS0wJ6n7XksoLMB10o
ldBqZPPZhZnmACrAkirGCfE9K6VebtWuFXfwV2kQe04q69pqtTkt5MCXyrXvFtVSv4tpRw+1wvbR
Nb0oH9vso+TffiugGBrGR0dSYaf2pypgTfN7RBy4eGdDZp+c67+kl8lDxCXjOMyGRBOGKkbTTFXx
mXq1MvHDsma+SBenpcKgkODExjE8WsmeYYQmxXy6YIfHk7JfVKonWUlfQJFFfNnD47lpcbyhJJU5
GKsSuLmfjDqZdqXtke+cJqBQHFsabAIbV6j76YFhV68Sd+Adiesm6CNUCWXpVA3K4rbJDYSw/F7l
+8bst7K9sKbN3eEm88jmTNOQUdPAHZwQpTbamknmoc0F9ftIUUJjHZJtJym093S8OIx7CkHhUWTz
G6DrpUNRyAqJTWR1C28t9+TgfLp55WNHGwNe1a6wst/BBDttxpobCXJKIZcKpUUtqNWf1M8qlvci
fo3uGxM6HMHFmHSht9ApAH4PD8962u4YZ6c3e9np/yxjjD6OF5MBUrbA3g3K3tBV0s336T/8baWh
BDPwXOg/GF4pUKvQiQOyRFC8PNf+o35NKyjr8RFTp3hQ+JeBch+YN+3yN6SgZX1b3KV6VAHcuPlU
dgRf8H4ockVA7MhBcItAMnAZXamzTMPR9YgZcTnOeg2jdFCrtQUahs8Cf5N8baB9UH8AVFtXBIDU
Rkj5MrGKBErp+4pwgp8bO6ZSXqR4xkUqu+Ezt64q0AQ/EYXNRTK4NtGsD1Cst4XtjxRc7qmD39cn
IrdHthjf+MFQ3QJMO0m5f6BkiHaGYLpLYIPk/xxkH/QnezZVH4eHkx/BAIpudcIAEFjqadurbCG5
RnnTZVlX4FQ+QBNeoqXfT2qyAK3erlNBQMgGRpIo19xqBL/VP/VPVjkFhMBYMfODVoJphvzh6/N4
Brf1fxnvODTff9QentkIGI+binIG0zxK2w5sHzfahrA8k9GSCatUsLyfF/2eBejx4p09qpQX6zRP
19+Q3OxbFPszgKp3MyjpdMAQOqKqlBMqmKm+YFLorch0ulvfBwvUNx0aIoZRQueHFzZJW4Tj+jdR
qPJrddYSIbSi4bITo3Gxdd/nAlBuTLRKBtiCVY9gBCLjZt/fjzuFDbSzASIRUUEtpiIhmLP/b0JE
IGQZJSvUkEmPtL37fWNT0tXO0bI0Ch1O0TyxSsKbwUpR7mMsk8TEdIclYegZN0UHHDQ1zydmtCDp
4iTO0QCGefHdCsojHzFUWCu5f7sWQWk3EYWTYuX8X+abM5xzHVNOgwIp+kH9dEeMiyCjPIzGf3Wl
HPezTXKRRXf68w4bIVDloHzu438HnetYibnDIBNuM0ZTsz4J9mFjuF58g1e+1tMg0c7zes+l4XEW
5Mv4d4G3NV1rZdaJOLkeIcNUVDI3hKR33SVKT9cY54aoGjM6eM3VR0m93BV5eSG0DfMO6Vf26o5R
0AIROC9kA5c4lT38qzpguy+oUjyGqeAis6H5t8rWQMJyzWOPcmiosIb+1EDfLOSDAycRVHLjPdRU
+OEhndlkPmjF01ds5WqrZ2+zXadHVh0QjiA/IZb1dvP2Cqq8nUhkHEKqKnzZriighBxogclckG8q
EaxWf50LBAVxh4bBTTupS3NgdYSyAopVjW8eC2AhthrWNOlhUBaVWyPpipfsugHLjRtCJZDbaLzS
17yuAuTZcIp/nVbk7kdl8LlugwGnIA2k5VBiQC6jabUu3js866bmIozNuHEStjCVKOuDePtedinR
1Qnog51OZVCAlto84AqG2rlJOTLvchIem/gKmRMgtsI+D6JY3muZWpjQ/p3WmGMBgaPN5SxKh/QG
An6BKZa11Q3BriP+4A/dOLscEDkkKV7znV9OD9lFB2HDZ+6c5ekMfaHgENmjyac4jWthqsF0uZ9g
ojPusA2McWzrcKOWjR2i6/BjbSTJwsSgo8sfOqRlwkAtEdUEgQAAq88/XTUJjR59m55zwTVB1Hff
RrhyVkHJ8rU2AMpOeCHXtp82GEEqpdreNny4VT6oQiE+NLXiHEm6Nul6WwKev3vus+htPtYeP7iU
kYbhpmgxaqgm5NicAXf/7eYSPu0m9EPVoQtUi9ZoUqjmY6vnGe34eYmYhQlYARXNw+wuwQFGplyi
ow3x/WMJwakSqG26FAJJwUhaNJQ2FYkamQDisVHGvbU932eVUhyuU1F9splItFD5o43/iFqM5cGm
1kjoPR+dLmr/G6lt5L+nkZ5a0gccrOj7bCjtC6LIGv2B9RE7RCOSeu3XOhw6mnp5NP0l4c3OsbAx
FTONrWJb1wf7bmCRM+AgXqgjeVQRtrKcI5zzet2DaL8PaavRajXPLGmtmSi6FOeYhCEcpWX+TTHB
rfd/BTaumAbZpZawpcFMRbI+28IJ6dqwvLfixEhjwAgECxj0wVHjgSFOcq5TGs+GL0YR/qTbe3NJ
+qL9G6K7UXi3JO6+882UrxEupUqqAepUK+/IRzeXImlD0CVMmeVPpwv3GXC3E/4vpRz4XjtNTd50
KpxEX9kPQctQPjalECzKi672W6p5Tb9nbczWQLTO6HRm0pV9pB9iLTql+cMRllwGwsoR65awO9s+
hqVLd5DxAjehE1JItyQlkvBwCRw4DRVj3OnZ1bftYGLPO5LDxm3rraYIa9DZTaNBZdT9YgrRPDiO
md2hWHuJSw76OGZMEpl27ErP/sLus7pyP3jThy+la0zxtIWN5knAS7+ZJGdTKWadTSQHzNzfFkx5
j73oMLnG+Lsjggagwp84T3YNr8THn96sLp+Zof+TvEUeF5p5t0S51dx0AjwkQDzmwCBW4RySwnHR
NMaUYdsGTMoy6Jy+LLW0HBGtoxniczerEm0NJlNVdtT64kh8wOiywHynA3rsKDt55bBqsOgSwQBp
b+oWHB4GmfEn+5xtVJeq0/wSc9wU6KKeheKO1NepBFzryiWxXALdfQUB7YvBj1xzhBHpI+U9VKY4
5RWhORHF3kdM4jY6dkluXxOZrRqJfceOmN0YtK/zxwgrAQBH/0gUFamA313TjXDGwUjw2N89lFFc
sD6G7PWM611zKUxzdTqAKldkIZ3iB5QPQ7njstLZVSkulH7bVlngJRIskwFk7O/f6akDvTu0i1ib
6lJ4Ky1OQOsIThLu5olr7GxwoyT0fcCgNC4/80aD5KV5Ki4dAY1ZdMDOcr2xy926f49+ed0yX/iE
/8w9HP10jxh0tnwZkulhAbEvzCWCLkmd4or2GxqJmS/QeXTPm4Rf7KBTucpCY523I0kZGkQZw12e
Od7kL+TFmdT7cQqlLgOdjC9TIpT+zXsTNb3BC/6LMwLklZ0G8jlnSJ5sA4MJR8MBD7KEODngD1XK
duLCqxvW2sseWzHX+YPGHXJKscnVByI2hD8aMd/Mc11kpp7wWpEdcPMYpv9chDIYNC1otN4v3IMP
NXS+DlYExlkqBz8ZE9DyqyrzpsXXUEWf2DY0Eankmq5Fqjo6whO6iQZ9Q78iTk77bCzFFKSoLUpp
Yh8dJQgHbXGhnB6vI2M1LePmlD8O+SSE3Vfy4FnQPG53/ySXSM/3S0cA/DPpJDdrkMSulSiPeEVw
Y3qZ2x6ynmGkXHI+GAlEKc2+LNI9hjHuPEnehl7BlNcTqxrclcLx2rpXQJfYRHNblwsjEDV6DHTz
K0PlP65EBAN3YqualKhBZQAwz0/PLOEozwGGtOxxiNHysZf8vClBMJVVXqbk3nkGEtDmKeZrq/T8
bMrJ/aqpSE8UBo6R4StveYUfiqoqoLQ39WnpFq/6owAAXnaYwPfPsUAwQ9NhW7V/p/A3tdR8LxF1
xHTgPOnsLD792L3Dfbtpn/pWmwgXq7aCH6871eRP5QAtYKOfrZV00LUwvrMskio3kL+NU7DjmlAp
g0Tjj4jUzdnnxlb3E44tSgh15on0lrA0J3QpOGAPQeSmTKxnNIHueVWBcfwZdHbTDavMZvj5Smg1
gInoYt8f/47gXQtxl9WP3WI75Pbe2XyIs9AJ85Dz8BM7zLuFbBCITnjY4MdxuvWFXSmedgt/KIVj
GI+LAZZ2o5+k8wYvgdcKH5NslefbnToLtEHpkF+BmuNxgvRomov1+vSBNeTBHAq5lOmi3wRl3TP8
nP9rjIcxTZdkVUxY6QFy0HXqw6+mtqMh+d4eAcm1+nGU78E18KSvATshvXc1MmemxMi3sKbXsFzY
xSEc5YceqdFRkRSjwmqJlnxWK0wyLy0mTnHsXqLX1sa5XFfIsKkcrg8RPQM8SV+uN+0MX25VYG1/
0WdA0FfbDMAir//xdlAw6YWhwgspy8O+mDvd9jUKqxfJBYrq+Ku7lbUs4mQBb6OjI0VbZcIbnLDA
NLib6bi4UWpm2K+qcQ8vW4s7bF+l0FiWwOJLDxLCFmjEWMj9uXHBaQ9nrG8d1ZY46BMhJLYb51Cp
rvG315BN0zf8mF34yazHYO8IvTAzI+hf1SFx+q21Wa9ifEKpRM7RNIvIKxHsfHZWI/brEgxv5u0G
7XOMJHiRMJaGigFhFn5zcnbSwhD3vXokt6PEplUhsMvfF1mpsKobc6GzutDkeNWFk6AMZ1ZVl3MR
1PUHKTVNF63YxtbKQ93FP42JQjp3Rryr8TEYqXS1IZuSpb/bI6gVxwgTNiblzRsEQHj+QSBcuYdP
fOfCyytqEAGeo7lNEwhWcKH5HhM6pwKM+MaoBlA/2X0JUk1013Xas/vU9NsC4L7WQ1zNcnMopJmR
g660NDg2syGNXjkqg/zIzHElXrng3DipJdhi/8Br7uv0s5we8gF6UJNPH/hAVeJneijEgmpLS7gu
CKpPTwRNfaSK9+Fil/U/gHuFUbZI9UHl3Ro8WFixkeoR30IX4FKXqEXp3/SYuiDKz/hJqEAXQnQE
mhaOgB58lkl//egqsmo7N0EkQDUogZ4GkAOacPa6DCnfhIlcxigMQh+HL9J2jmWmgKORH3iFSFqz
XOuvmU4sTgqMhwhJ9FpieQpA3a3/BPh4qW/eJQR7cT7iKyMf5XblbFoHWwN+k78DXHOCfIT3tTak
9H9VlWuejutjgd+zGUBrJ3I9REDTm9jM80IvI1nfcEDRTGD4RkHLEjirf42INR8zRop1X4SxjMPf
qDQWZsrsI3nnoQWEZ9SIa1FWE3Qn/idqVDOgaRSlOCZEKmm1PYaWgP6/gV1Hn6zs6luxdtOdXERj
gfWQ/Er0c+2g3HJtJk4Bst/Z8SeZX86qXJkpgWY0ChemuyAoBQ7pmC56rUGTbg3+eGenxeciQSV1
ekoirukkvhz0R2K8mZkgCw+bWAUPrKpqrd1LQVPO4bX6M9/fNXjhfnvoTQ/ScrBmuyiGuxzy4ura
jkv8Cb39FsOpIQXdqYy9YX/JeniG9aTNaTqgjC4JOax04oWmzjst/da7pyBWloI2Wo32swF4ZAii
CuVOPNCJ6ba68xajD/0J7m5wjf1C3vWlbm/P38IpP0zxqFwnoJZSCq6WF5Bh756duJG3hdA5X5ph
medT+pO85fbeADDEHOjf0Jw3spF+w50CdW+LRRToulfYbmFeTYJrJDWUKxGltqEEDf8rXtaUFchD
ypSlCSAz8FjdZegKXUN/SOrwPzE7nwgLlz/mHIOkSbxt+IIBLmyg0u6dqslz3NuEXw4EnWVpMXKe
QBnePYuRb5zTJeZ/I9TcMJsSAGULl3yj8QORrDffSF2ZmAVYPHDDi6bS/wBKCtxwdUG24C44j7Da
dfWTFc2wpP90pthNQ5ZqhbK3oXEmkyXf8XNvxtnBqzMAX/uXXCQ1pohdyuB4RJkEULDeFBUT314l
IOSsjkUqeoC5keT+Mt72M8USyAY++aoT9cLdnygDLLhz9kPnJSIjJaIRQ5dmpQJBki5NPT9czUE1
3mpDFHOkK4SscqQTDeS59XO25BGxYcz0h0xujDkzi6CxNIldqOXjbwaQJPnh+wA2Cm+PGnvWKntx
OgCAHw2F95iYNQY4PsQ5XlPSxDby9HhEL5Rm/35HDRy7S2siTaSXG5fMKrsWL7BlAEHtUjYU75n7
/QKRFV/v46AQVzRgtDG+KDLNvl3ODgQ/bRkze6PDjs0TpKZu2JJD1d4zWLQ8XEZzNgClpaXSZ2BG
M3yuQaY0XTfxqlxmxkhbRaAXRyWBgq5H1EwvAaIu3byUl+dwjp8yMYpwzKFD8c3rQzuG/dkV4Lpy
0TAcrRz7Oet6LcEw2HOowhX3eRRsF9Mal/nh8AQSE2jrquo7hMZV+yVtGdiQ2FFaGe25UuR5eDyD
BjJvIH5ix3h/AC8mCuX3VaqSfYo/KsmeIhllx9KkofcmhPO8eHnW7j5fM513b9iTg8EvHVs7784L
H4SMNWx1YBOCABGSMSDMlUOVTxypXVOYk+0w6m9Aq2SEqb/LjtAULtYDRAPNuRhWGiFcS2NuKIe2
xzRplN/p6+I8WAPOV+djEWix7GHLVAFbrnJKLNHZXnw8r+Bx1vUZhlHoMmYE8vL6R5e18xrp2e92
ekHQ0/QKPbruzYwS3a8uiV8rhSCooikJ+wm0aLrGPHiR+ttIm6+1R0Bgp7hVDsXW6wGFIE5bcZ84
bzXr65Q3EKqmGJPH+DksVS3HW1WNnI37rGx0OtDHC57I6Rp1sRxQ/0KPHgENcSo+ZLhpz/exQjjP
AK8mp1Oo9CNjx3C5gwPMDZU+dJIi6jUS5bX6TORAalrwvrZFFREsByRKnt5RVcHowR/BzROlcRxx
5voNwJao8WPrrGi1qC7ifjZZItslfNxKCU6/eKlq8eVrV/xE4UFTdlrSRGrxhMu8emJr8ZiGIfZx
ZnZ5F0xqkjQr4UDopJjYkxCTu4Xl3r3HYXYB56Djx2fONFXgUdUryfW28iWHDuU6WdaEcdrepaH+
5HSkfjxuh5k+SKBH6Nvf3cp1ZKJR/QiSm7awVEzZLTDhSUBLdcXUXTHLLmFRuAcf5GYC1wcpyXJ6
InvPfB8eCyHYl85FTe+RbFEZB0cVkfswwu5bq3cRjtEUMsFbbzKHiBbZgUKuI4RFLOpalHZ2AnOO
dJB9JXl/IdRLlzOtjeoTrbtv6cQvPZkfKFZKnIa0YmjXqq2ZAtOGounun3KHh4OPYz40RBJ1o0xP
1MLYxuCft2Ckzp2XFb4JEiTvNK1XZ6toZtMRVTdOeUCQi6s0NUWdaRLQWHsxxODX85jhz1GhISHa
BPxRW/JOnI2oRFQceCn5rL1B1wyHpwwU+7DVjuCAv8dzMdSfL0EWzR7vZxmIPYzLtMbtjq+/LHZ3
nqrEtbcGK8Su0Yoj/ElrlbJOijwkfP5FFAk2r0Fkh9gA5aplOCvJpFShh3BfgEUzG7gx75qhO3pE
4I7Sy8V2fG/lqsmsCLUyLireKToBufpnDQZ3bMpu5MNQt1Msphx82T0R77HXSnQrztoXDTWQKUqm
ER6EAs5mZzNbLh47ybbRgihFWoV3zRT+zayVzlRs6J6snaH5v74Ua5wvS0lRJjot6QAq9OHso3yJ
D/bbjS6WKX0gOYk7g6s2OjlmpuRWfvs0CUaLNhtKGOAkHgF4XM9EVlYAfJWE1Kx1peDippD+nQEw
7ir27wqgdLntSMO7d5PwvtZt2B5QW3jgemkCGfLIVEKLIzJS5aOyepATg5BWCgnoQym0W9LB3xEc
V2vCpUssktCLoMmhBsbviu2zrABACaYyhI9in9eoKd7w9JgEfuHEz1iT9ZK+u1LKUszeonA89H0K
YmRXn+nN8J2CuixIH1M9Ms5t/B4c/wCVRWTKGY9FK7Lcmr9vHcqi6Q+Yz10zZaJAYZn52t7ZXqUf
BeX1p+08tI5hku1xezktkMmAtyUnwwEXKSZWqDyI0TJOOk/K5lioLySbltaNTpaQs6Ey+kZuj2hY
4r9jClJVQawbKGCuyfcoax3HluWRlGqMH1JcQeiGbJ+UybQl5xCh4qqAmezp6hVau/ccnL2ck4v+
/rxXWqOboiTj6q0xxM8waFFXxevjdVbYv0tFLEVWH5bFkpAOPHbqjCjiCdftBjYXceWxT9mI76L8
flvbqTKz8NiRt1WKDSR1h0kzqQLi0njwc+QFtuCoLDEerBm1PPsN6g3QspM7wgl+bf5EkFpq8+uP
TBG5cT6R54owtnNSlSnnNnGxbvCJM3sXbSuTob2NP47bKnKv5x9YVtf7/PMzTH7XaJjCLnC6BIPa
Umn/PHHv6x5AQ5+jcd6uomgrX3CICU87oAsG2TQZpy7WHk4A226pi+dm87HXZ2Pz1AS6zECru2ux
ApUnSNHPeOOi/kyxonrS6zjSPcJyWqWpEBrS2dQAwimph1xDFpyjQvWs1QdndeVI3NLQp8pvoChB
Z792nV+v5XXynN7Uk/3muo33IUgrdQ3Zied9rVa6Eid9Sgg0LLcQybNH8bZpelUc30BBZ58C9MJo
l9bV4kpYRcudRj8DPC1qRDC7Jmtxla+ytPEKattmvUKGOffZ5saRDHzmo6srmMFq22aE9PFXIM8A
5mFvpuQ/TdvIWL1zOVgQ//A9bDsNBm7JLYxGTW8kDiOiMjcvj8VcRnga7tl9xhap706ddYojPqXb
cR/rqIg5z4WdEkTeAlkgLHvZkJMNkmrNcXqQWC+Xv+FA5lm4nU5GkACTHrCtXhJriFtnxcCAHaIP
eJ/mvg4Lq/Y6P0SXBf/056oMMwx3vbrR22WWvSXeLVrsgTq1CU3LPEFr6uShjVhW1OlnppTXVWMq
09J1fNjy89vGeZRE69Bb3ODMwKcXFurfcuE4HhmKAJGDhIS6s7dIQm1wPQtsdDj55ZStx3Enq5Da
oXxnfOFi4jiLjZzEgJhi2Ai0jPb9JfbQHlp48d8BWGWX8HYxPviMXarthyjWyt4fEuC52cl2kIWl
q8OtXd3hA9geKR0IwezLPVvHiLsz0EiOKOjCigW5WS3INKUSS3HhIMjUtCEOYnLP5fJ+qHlBe4Oo
Mzu0m2134dtaeEsKu9ZIlFzmejUR8seEc2jDJ06Nf7DCHk76VYu02jimrTJUc+fuUPyrfGMb0K7R
ZU8ORZ8N+IRmheOW5Kf83v//cgufK3e8+qYEZZRc7EyJDt1UqPZnY2JMFrMWX6PdKRgUYHUkPMBd
E9jh4xN712HlcbKKegHBP+tmGAj4DQPK/oPWsYRtT5W8WmttfsyPNruKLd5tOMVZwC72jXlkO7qd
GJM1Ibc5kPE5zShaQHbYjqk519rsv7f+ly6MsApuTzRuwbmEKChGUUMRK8Qj/BkVaAeDtniAh75x
0ttiwJumKQ2SmF+aRDZqRkgniwHqL8d5BxeCTovCaOjKii4i2t3tB6+lAaZBWuiB9BlU5EBwKe0B
CrZrKuCBCBOBMnx0GziKMKSybUYUJOEYrKF28XM2iEkXgZ8uU9LFnW2v59a9jDv4Nbbr+ie7qXR0
JbrJ48n8EKHOofMxyLpLzpUw9ttxAjpGl+IT7/UTrWFv/wDF1D/dCtpH9JJCNH8/HeySnZqcFcLd
/X6im/YExNypobKrFjrmMmPEbOLPyEzQOCTfoRv2WvDkx02nH4732VZoky4c5fx62rsx+nauHSNd
Tn5aeQ8Mgn55bs0IstimHXlntpl8yKWMgUELAYeh9kxiVW9itdpF30EXy07QTiVCNizhmZKoDuBj
Mwq6sRzw0qfo+wCwDGk92jkjEKvcSyhDeoL43IWKL6Bm2lLshj+1T/GfSYLGFCDOPk+QimeYXIQq
0jdlqg/fHeQV90jLX27CNVGFUn1U9GqRyjzHHenjIsQGX5nzopa7T/ia3/Mo90YUA+5F4lmUdOTS
F9MjlJ9bxzRLohaO17X4ElErDTL/xZMDeZ73VtqSgpUB8ZQunGt2BcGVT9pabCnP8mlUjd1T4374
Vnkq/+DCUssk96NLcrYMxnM7p9f+m2AN0vrFMA2UpeqHdo2cscMUnhSijdeVA4NQamE5ASfk2rBO
KqDN2NOkEwUMjUTvHW1W8k8KTc8TsNrmvDekk0aAyjsr6j4T++f7YAGlG0RMDcjun2dP1U33OUZr
ULjBsz+CCoXmMm8Skr1LIee/LYc5TcGQJR8ZQ1Ub+T9RiukWmRIv3kH26ODheEfT4vg+jYnpkBTT
hM4iDfpR8xBO9/VBvhEWb4g5MbEs+KqfppdI0wKBLJhL/BkDu/KbtUQSWXH+T8gXUg7n92QZIqms
6zAKnxOwh61dzYY0ZsJ5nmCyBBJgksWitPj3fi+PipkTxJdRY8ndgymUhsfvfJOA2/yIQ5glLawc
NUbavoU90iUk3qPP+E999BmNbeky8+F0xbozVibXUNJ6M2Lxr7NwQL4hjUAmDAj9vb4JwaQtZpbO
CRcIWQ7OxB7mtVnnbNxAK0Tli1cRtURQ0MCUaDlqC+7Y/Nyfulxk+q7SGmMXPLVUbY2S1/1ujyHp
kN7T9WwMXOInVANTNhH/NwVhHUv7bKLVfOaW/nYgJKm+thfiEl66jOb1chMz6eS8gLMBEAKs0vk0
dnKV4DIZt3OerAlofGnz0rGydN7sOjW4cEozZNiONLC8Mz2jFRCapvFPTYXrYMffJSLDALH4YFpi
c+NGgqgTytR8Ny9vF2BGPu4EDajL82M9jm0TXWXTEkF574RLYo5Gf0eBP3rartViFjMOi6V5ROyY
PrsvUkMCi4zsJ5avptZK76FUkE+mk8x2/Isn3HqwvCV7pW9TqEJZkSNL/8yrdwSNFZzd93pwPaDx
BeyXN9+lUdAIuqSZTAG0s1FnTeB6Eu16omQvk80FLUHUQ3ELek6K38F3lrLGJO5BWueEODa3LBfJ
vRz9rHvDVDb8MoOrcE/Di93lUV/QN9LCVzxc3FvJcoTZQLpG2oq0XtyglaroAZhKSInVaYvlFKUx
V37DxbKyv8SJqh/6T8LNw6Jq7dizfDaK2oiEoZ0C0Oj1YbGuoFs5I2LigJDSFj2jEdlMCjeEX7AF
viB2wUrpuErwfCQo3SyEHuoWs2Siqz6lrGnJ2segGF74pJugeQK2rbvNGAE10k7DgCE4zixAb6ab
Sx7R8zsXoFsyVm9tZbTRAA9Zue5g46n0arKJtu/3qtEMSuGmQ/nz6sgYKyMjrIDTqp0jJzuhwFiN
pMlSHv+H4pk5ob1Bjg+Euj+UDjHllhF/KpUFJ4WCAwGXBrOXTbh0UnAgRsxPjQCnh3TYqZqEUqYH
MZJssTBNnt/oGoAwtp8QGY7FB1kANxR31IULpE4+CfGzXxqLLTg2UbmUW7UvLBY9VHxFG76BBW+C
fz1eEasSKULeP8CImzG4S+SeCFWns6gPEORN1t0VfybkePfta++3jkNzJqhYL5arbEOzJGx6fD/g
UsjFw9HGOZsihzIaOZhKEZnMEB6JV8RinL3HAuUzO2IdKDeaz1O1m1hLVweDh6y1BipZeA2nDbpV
ONQz83C3BOquh9RZStBelSjy0VoJp/GWLcPRT2jKs5JHyXGxQy3Y7MbfUmq7ksLeA1n9ePgO46bw
pbLooCWmdtgYdw2CB9tcpHCrWg69nzjynOUnyawG5u3l5KZrerGnO0G4fB8y4150qaIV4J1TsXC1
qhsAci3giom/Hv4AUFYfFIlKgCyKbk7+2zTV7SDRaYxez4YOFOkMup//exUZh7q44JWqCY9/WoQM
Wtxn6QKTgy0adHHIAsmRdsmVJTmZF1mh73gfWldwHISO2AgbMVNNAqDnYPeslXNXlkuVpNwX0vny
z3b6bwsw3rdPNLK9iOuytZaWE0XxoTjudbGcEZleHiUmvVXsZE0KqtZmWTaQ17D+kNKMQ0cIQnHg
TECI0vsgsZLBAmv+h+WfNSWsYm+N5b8XSh5mO73GFQbshfbimcp2d3kkb+hcKb2FElTrH9uwnVR+
Kf/KvAKjFHU4JcvKfsLbqG/0vNV964nX9NpFXIctZgyss2x+Xu5lSmj0Aj1pKyIU1PMyA98DWZTZ
QQ6toq/o+sGi/RD1sz5b4UJJn68+DG34FEStbPJ6J0G5IyqAzxpQ4jurVdpO9SIMRIgx6uDZTlw1
5tLKdeIKGooFFPYf29lF32pjAO8xvVLw050zP3WSgiFv48pc9LCmCkTYGkUia049OYAxXlCVLRd9
2vBk4LYQMP3y7N5/oDhiNW9A4PHXB206md6hYKNFXvk99vS4lZF8oA2tUVgY7IBM3EtfppxWL5QL
5wzVvZkP1dUIIm5HxWwDJy+ZgSqo+x+j1G+XjlBICGhm8x1/VV7qJK0270Anc0KQF0NJ5LaNxHe0
s1B3slsRpIDY6StfF855WSOF1x+fsKaOCwpgVlQZJVJPIGVJcoSUePmlqbPFR46Sy5DDb8qGvx17
Yfg9U1fkK1HqSioKMhNTbkkcTjFHI77VJw0VLXEku1fa89yvRJ6XRptgp22t5BtMlNQx4YNG1uxg
PvWm0NfSUB1drnfKQwBuU1tnv8g/ZMHrSC+wHHbEEFPkCFMqFo/HP4jDXwq+NvKMtiDZZVAzaf8V
xpKrIn1zNSlUr3WpOLtycb+c2cyUyf8RBSvvaz6Y56bGIGCJSdwDdKFYbAAPwJXKeLqDTjQvFG+1
TchlHvHFcA2cyIt/VeSXEfkICciPfbhWT0DDy97ve2vof/skOMZlCqNQJB2tEsPISjiplG+EQnZW
uQ53mEH/DdzVFIQQgBEQe5EIaXuaD5p5ETPYEbQMyPUTGzAR4X7X0UR3F7lSo0ts6vh5JhoKJPtr
nlEpgQfE+yrLlZ2ef5OBFWqfmDxJkn1zgDa0KeeVW2luOIMVJnnk05RUCmYrw35Zuhhbyq2ek6f8
qlQYT3c3nQ0d3b52jOcHy+QuxKjaFAgthV2SaYAODCxhR8yTqNMvu16GOZvsAItY+lvj0SXO5fDS
+g5bnjB1kRnE6DUthtDT0TLGKQwaHaG/AfIiuc3t/ADI2E1CRXTDYG4BauEJVeLTw4Gwbutu0tF2
hlY84pqS+2PM+1gn10TmhrE3okFCWo0pIPtcqeIz2cAEEF4kd6XoIEQhsd5pIBJ972yuxNCYjGq6
02pJrE0nZ9u4ub4G6zwO7jmcYJTUSgoyqM+jFsYz159vJofO9dOyuGcBc4i9mPxNkTzSyNLvmDGq
Xuc+87XHPlb7YdeleagPbhWzpPzhYFuwQKDZ55W2Qc4Mf7stQ02+SOOBbc3BUYZ8NY/5PfZTi5J4
uk54CZ8JWBw6bKoxGakBk6Kz70hddhrnp73hrmmHxWx2TwFHNJvFFC4EBFVh9MFw5ZzK79Xu52MV
pbC6kG6WP9jdVQ0EA8TNXU7dD2U23FMXcX//o5OKBvDLihBpzCocDW/YD/YAIfoWKL+Sw2lUbmVW
u+0NCZYsmDqECTsyWMWuQyhHqKkAGTq5upecr/GBvbJXJcrr39cnA5haRJpGTnedlz0UL+m5vxlV
vjrMqsgore2zPPIiGGdK6Y2jAciaWLFZPB9Bp/Rx4suRGf3lJ5/hDLnNSczZ3tWK0VwwMOXKnGgP
tdH+U2peoatvJsGwGmPP9SnoDrZaoc8ayj5ieB1ChGfIT46NORpNsTx2PEszdgtDX5Ym4RmO3wTv
Zv/csql7dFF9DTpEHveU9zbaStlB5reZrv0GrHiMGxHtsfopTDnvwzKHdA9qWmwlcQRziPtKb2DR
/SpTgebH4pzcWgkKM9Noz3nBFEWvM3Toef8//k6/AidByB2Qs2Dv6WuhNyRlQqDmhPK5iPGwVa0A
dUejNsuiGh4zfYkRDos9lzNQeNq1RJh47e1PMdn96MTOTiKkFMVzhomcy1eEp1l32CySSqEuZB2H
HFwGCyBzVz+j9R5pqpP7EP16532zV+bu5ZdmlqGll7WTvhPE5i/SUEVQcj5pqdfE6T+cgUObpL+w
L+jei9Hy+hgieSijtv/8KraUevrGGeHZJI98fkpsiu94n3LPnCVq8+Db07Tm0ed/jJEJ4l2KXrlo
mn3q2VmGnvHB6s5unD8cUu4OQcMItZSfP+W+djNWXPJjGhDhf13YwJil8yuvNxSXPM7Ri6aFZTkZ
efrddC4QlWavTdYoe4J7wstPIFxTkhA/yYvjxm5fioQ0FVroyw8jGqgVaFTEys/C9XBIGJSTmlGM
qjgBEvuf7qU0HJkOy+B8leeKM6DMWjTozdqYflu6+/EZgsFWCyenSyf2RdfkzEd9SNX39huyjLrx
r9Bs0fsLJ4pPAJwx5mSRhUraKo12uagLy/1RjXDdSkPQDQumnetumNslZTHxwlUWtterQtomnhh7
zxDbKi5VWo6ZAxTniRnJdzkfGFKAcPWV4xyKkGT4gsxIwAWBommDU+O+4JdVq9vhXIf+Bz24TvIO
JPzSdZiibBXspp0xkFgEptbaCPz0fTDvu6PRhv/jhCqnWfIgl+fZWCQDOnSALtbDWKGbbH9Eaefp
3QNZMqiWBY+YfQBfsF+5ggBAOXNRhYUI5cqFAu087JXU+9dkYG4r7BBwiTMz3+F94eJ1paTtpomO
E/emcacmPNwxs8JxHUvf8JPsMfNXlh0OtYYmJgf+IPIfJuHYmrkXTOad6a7drxkSx5+qaXwASgsP
/SKcmNp9e0vRiEyE8CBcJlJtDcbtGf9BKJGt9KfDyHSoC8O77GChfMIYjvwAd6aIPtO5bU+5+dyz
CLVYiJlY1QzRA0OXZVjv2ixyXetCLsLEFER3b/EFfupLxrI6qqLcN8wKK458v96SQWebDcKS+36a
kAJgWUZDADA5Srfw6zACnN3Maz9qW+qY7Qd4wWeesRX5eLMePfpIPbgf8fsSzTkMqzeX+1Jx6tiw
BIPHvMCKISRqLnOmnozp1FnVXyaZtLqVFcIctxfZCbouqg/Zz3yMx7OBiySW2NdXXV1B4GuuOcoV
SZ8l+pYeEtDIwFJk53afxfinJvzYvBN0o0Rek+7YK3X/ODqHhInhQ4STDglPX+T/frnz4S+MYkQ6
rFvy7lEvYFZY8ZrkH0M1T2yX9GIizacLAj7bb7p2gir9BKlFl8y6Cy05ovayJXvwBlrXY1SuAaW/
W5Jnvebta/7Yy+cEhTEsGL0PqJYp0MKfa5aFaf/V6IF0pGv3wZVjNGpanRMCDQqkA4CIbcz7Me0S
HFaR0bSy8OEOdcF7Ta+fGRBYeMeAesEdjvOsriTnvToLtq8+UnCOPmpWXGvkySpO+f7I4fKdMPWs
X2eKLEg9YI73dn+RoQWvao1sP2Iz5Zt+84AxDIBEJew2Sd7fe+N5qNSY0BjaIDb06KtoDrTRsdkn
GELGLhLLGwmMntYeyQyPGLjC4dPyc27WIwCbjKzLhVmkO5NaFZJovNK+MA4JZo00cXCjWFvIpBjR
p1GiNXaKogcWw4z1iiIeWPyWSn3JkD4IxACfasYhIbBAyGFSosRQ3g+M/S3ovHp6MtpIq7gFuHyY
ni++/yvW4ITeT4aCbENH9EuthwAK+ug04f3zjg/F3ZuvNEr2Yj41AQSsru6ImQxaHJeBc1iez8tR
xZddSUybbSl84PRzG4LAnK/QuT7aI7ycsVLj6FXCox/G+URkj7fn1UWhjUrfaKs8mSnGyKFVcbmv
uPsGzHKhfVhltpqkI5kCeKj+TGRhuUSGp3+9b/hzxmz78+HJm5Il1730i1cAArUssp4+sC/+fDTH
gyJaViUB40yFGF2dmIrYDMQ13+tTxHCjTnAVsRnin65qBJfWYakgWZav0vOTDf/fqQM3Y6gpEJBd
grxyHkDkg8sQzXl2GMqTpBGH4EtnUtDOyly1Qxper63F8PMOM8i2oLBUsOrlSJpaX0I+faTfL6Ke
LAkA8x2oEzvwPeIOJ517JTlgIZu2kaJ2XDWY4JZ/Gq8jqqVmqSw/LT7oKC6AVPxEG6psW65o4T/O
FNziIUxmyb2za+GeA7xvJbd75dFGjoNKoj1YdYjG2XNIP+5mLirDeiqydwweRY7YyIABGd26QbGG
QMnc/xCZzL4GrE3SE/BxB3g2uTWUTNef6IUo7VUEixFI7Tc7PUa8zmv0UxEG43Cg5WJExX0brZMc
hadeZu1hrEbom1LJxDTdWjduLfWZuakNsO7lp0k23fPTrv/MPydI+RUHgA/I7hR6AFwyJjDGdWI3
fmIhBiBEZGrGkVo/9iGS2MUI3bjbAmeOZ6Mf5/v7W85qkRlAikHrlqS2+2ojujc3FUVUG4CguJ7w
XVHY5jQc+h5XEopBD9MXudVTPUrUnCxsv0PXv378wQ4iRLG/5cakA9I6EWgFgUjEiVtvmqQjZ9bR
UCcBOvUBJQPKPF4wO00/u0g6cWMzlesC69XKEHkbnWJ3qFV8wU58f7tdEbFefHiwacFVVluIruc4
ntvtwfADSy7b/8A3wyPKZ1cDcawKOLxofmdNe8N/EscjLpHvtvos08gjV212Wfm6FNL3VFkpgbd3
G+Guzwd5m67MidWo6+IN8/iEKqYDXx7IJxGrxa1upUFXW1SPlbTCi1oW4S6t7nhgx2bFcHua0jxY
/WWeX0sMgA/4mbvq8tWciCtVhkgi6+rp9FNYUDkTC9cm7qsccn4//TZfHThDzfVOMOuMcW6c4Goi
YHoOaz7Go86o7GXGBUBOAH8xx27VaoeE8YGfZrPMggvPSaIJb3xrvMn6FmKfKhzVYNIqK6WBgOeN
Y3dnmEA1JsyO6dWE3F+7h2ynf4S0DElzN6rD830OQklpgfxloP5nlf36S1TLvwddglKZ49rCaDav
IQVkNaxwtwPIdz0mE0vrSzV/R1eh8VkqM9mhEa8TA18dGFTdcE5iUWiWltCT/lj6/kEsjfrw2sYi
TmOYCagiKJY/NLYyql6crvX/l8SiWscHRhVg2g4nInTFXNFesJoSriKf4J7UPQeBMIDyZBjnGRIK
A9/JYA8AeP2XSKnAEdIZi5ePStvqgnkXSTuq0QbKhZJ1hggCUY3nx0u8cZtFrFEnZPtHV88onXAV
pOri8uOrqnlV747/Ks8Du9FhA7uVb/M8UT3B2CWp8pooTKLcI4lugIHmOvx26ApXxdY0xgCzZWKR
Jj7vueNU9tZTKkI8LjGz3Nm+SHa9CgVFaWD9fNmG7rwQVR48cvU5E0gLpqI5xoAetwZ3oayTLoqv
scVP48Ad7mepg/mIlC1PfB9/5o5VUNxFO9vupOWSuFbEnp7/whZruk/ixMSUtdB0TB9OeRKryIuy
/pwCwQPWkklkHx0wfFj4Dpkrjtn74ZNlS+j7EgiJZs/GRBuuFn3F6NTy2YV79fMA+79GhrFB7/jm
GG9mp21pcFcGTbSoWnUjbtQp/teV7t7PAB0M1fUX7bQX8t46P5sch2DvJSCIpf44YE3etDjj7fZz
nle5/sLwtxR2iE3N+b3vmFDNsH7YMRuFb0dFeFUEQV+2x7iMGEMFN1DJBq29XqAElgyKF9hg3vnp
dLCpoaH86OZ/T0mAZ9UEo++kvpKjd6Iax8t2iNLCalnH9xirR/t52jqjYKHQLtDTmby0ITgi6Qvp
9VAPqOCitszpeoxU9AcDbHN8VDyg7Kb3HLqgiWCUU2aR+mQVp1PiCzvIou5F+KrtmqMTXmifOIsv
nsvaDeAshJr5kRFEfnSd+LHiBMZaxudBeZfsmXZC8ztAqKTLKLlLMKWAqLITQUq/aQnVODjmx3r/
uMr3TrzYvuFPISwwGi4M6Lrbz9IYC+c7cLGFWXXGWqc4ue9kAVpmjpunwuVH1s8VKpPaVywm4yBp
k49lbqpjhMV/eKg0aMnomPjccxnzhnMJCF6yXs3obObx4g/p+q9XlwX2sBy5O2M8ReIRxxTYCwfB
258FQfMlh+reCR0FxKKsp2MwdU8u6Ijb0FCDRoHUV2fZjdcGBW0LFJeEmup/Nv8pF3M6Z8i7FZMx
FVpbL2f46DSbgYZLXZeUYHSv1gysgfv6nWwCH+JaMX311qaHUKk6GlIWy7dekUhdIf2rmouLzBIZ
+qGpC/hREl+0lLHA0+p0eyxx2cE2CviBGmQkI6O91aeLUJG1tn3jU6x8Xk0si/8L1bBfjPSDkFkK
CHwOKagriln0uZ33Nu13ZeFAegNn9CmZGl49gcMXPhGKMYK2SXBsfWfU2CQdJu9xzUYsD8dF0iq6
fvis9t/JkHLJu2TSBIuvmEcvNYgbdmWh/WioBbvcYRNeoNWds/Uht7Ma0Q531jRNzWoh1E/87bye
RXHEknjFHa8BVHVnE/9YEVoDBLu+ja/QasE2BuUhjyFiPncnJgX2EgNBZdax5jiQ7c4tcWcygrOE
bTAX9Tiekt1Yt0rga0Ncd+GxhiGmfRxBWoZC7yl2cEu5qhNPjaS2T54MnWZJ+2uO/mKXiWyZ10hk
Te7oeBJqQcCCUIdboEIvfvP10el2q2EJa86hsWIw7LdYdGToPG/LkNZYnsIJtBZqjZHFtGxvDCEg
APIuoask8Xm3fUx9pE0896Z9wG0aKEwGj0u5Sls90/5Pzjq0KB7FCCN4z5+5J4w5McNbhPeXf/8V
Og5a3Ggu+ttsTKhTkZAQ7+1E15qD1ZlETdjFc5g4wvoL+ADUDG6LZYZTxyAKy2cyt5uwODjpKY38
Yvt2EoywQTUbqqpCpIrXM5TkiVHe5FkDpVELGQkLu/D1ZPkZEwIFekMoEOuZZHs8sKgbWIDcYR99
Jm7fbHutouuCF3zA4XoXkGr3bH0fg1twAY+HMnfRfCJKi1ND2T4y4fYoXeMaHXDJfWaYgnw6TtQp
Qvb6MukByNGZTUeT10w6pK+fpA8HdrN6Vn7CAxqxduuzQ31oYggUMoXp4WSI7bdbudcs57ldtuqF
Mq2ls2+ojfRrSo5IxS5E6tYlqEfNHl4GA9xxpNe+pDy1WNNRstO4vyYUscHBAGlwbetYZyx9Hajr
514xhUAbNGYrL7Rs5LXwTCn3kTYmgpF4McPlHncuE8jwxznKyxVsBnnWVnilE0S/JasX1woFexR2
hi5BSt/B4srdrrJMKWqkqRNOzMfKAFtzo23RyEKxnvUlpMZkB+STb2c2bodMQXCt3/vyqQnp0J3c
Q2dqaOKKRS+S5xRBhyJfhcaobXIJ6dsWjRFSgwMVk6YqDm5WarX14eNia0wxqtEVYKxbNevs0Gml
FyqJHw6T9DvIrSEngf98fSCCAI0pv0ZH2bLBeVdaI/yFuyRf8aiRiByqwvig12rMI+KjztbJI7Kw
s991XJ3/wRw+JlKo5OSbB/RgcqBwhuvHQ5Xu+73e6nY2i+nBu7tAEDvPLjQs9VT3BHbQqRblZ+IH
WsjmEC0qDd95iZQwdSATRrD50nsftaEj64PYUjb7nKWDX2T4CHWMA2irv/OVnjSUx8lzmJwLorlu
1jfdBFv17jn9+FM54RC6fpZmYY+0PCYP6KgliSeqjy30RqiVPfY6ZyqAwH5BfL34wR+D5/XCtHm2
2Yb6Exgd4wUV5jFv9TLNxzAQoGwaxkJyXe7rCJVTFZigWHfaTOCWlcOJwM9274HdhztNyJI/Z0MV
BpyVwRbsvj8u3ixaTEIBoBu06D0rCY7+5z2gBFwrqlWtHSCJhFYFyGoIo5AcsLEg78mpKe3iNUlY
mCzdZ20VoMU1vBVVkjGI3Uybc2+ySHC39duWHHsOiXzH13s2LoB6cemX9WOJ2JEC770kj2sAG/Ly
jNs5BWKqRDCbWbMAUKibX3Z71afY0VI6Sj6Y1NKJQsRtSvSYXekc3d+44G00Wr3qra2QlowbYqMh
Cb0AYx4wuUle7Y6h3LR72msn5sj9+AJT3GbSe/EsECawa8gP1YNJozg5Un9abDrl6mt4jbZZMK5s
rkNsKmr+4piOrISWyH6z/LhVIhcF+/h8YtiNTgtBddDsXtqAA+wpt3iZybnyhBSP23Rv1LWxcDwu
BYI4fvKtFuxexG1Sr0TvFsLPTMFO5dAdspAsmw1hS6s8dhJuS15lx+pr8FtbG16s+pJkYUYrfHhZ
gw0uVSCzCWe20RgyPkScBba9ZN/No69x0//LvQqNlnoxHjzbQv8TjRSo4qqjuygSCbGHaSlmuG9X
d1HSsdoHzjRJNEi//PtXkkJRr8QqfIsUq0mOQM9RAgZGcBueMfNdJJehWh8y9hdSZKC+A4i26D5m
ULZsa/mcN1ltLJ5CBk+ewV5o50NMPVMZrhhvFcRpSw/wO3/0uidT+gV58wmDnXlLQLdBCttnk+jw
akjEsi8/B52K4YC3yHzjWludcjKV4TdVY73SMxiL+LeSwnHUhAqFUl83j8Oyu2V6pQhIhZplsmjm
85NZI/Clz7fxtgbvHutePqTwoms8rXTd7nwVCeM9kND+k+Iwqm+XOBUI/1ikgRKN9D+fo7xwy6Ry
dqMMDIm9YmW8yi/24Zfvc8fv0pefaoQZ85w1V2Iv6zh3Xb+x9MCup3iOaOM55gercWhx7tZoewtl
HGZK40rb7kC4p29PuxI6NN/yunCSQsd/Ks10Z8zByfpZVgueYQlc2QVsud4nTMI+pTClghPWfLu0
jhWdwOT4Vd39M7HoQPL/N3/BJ0dGSx0IzowEmy7/oeUdJKiIR3flIJnznho88yPSqMak1KRRZnzd
H5g2dZQaBFYWQ0qv1dP2ut66q0rM6/lC/omBzJVem8sDsFCFOnowP9JihSt/ccmYhs0gtYH03I3d
k+87Y7PAZdIqE7ZJXu3WVxnBPytAiuONwLD89SUmlxiuK4lx+Z+PAuuL1q95pvwN49z6zOS6dNO/
CIJWmn6yIPPOt4WkZ6cLZzOlyhCuEJWA1iZer2vt0kfsV+LvAUSiWamADPPaDece8+V1BeTmRet/
CWgnSmxBcTgUDJajDEcvzzi8T086cGHQGwvvd7dZz0mR3fyrkoEj8Gql0CZP9GoH0LOaNqzrpv2S
GZlCT6/01nb1+ofoXcz5YSb72BkGooauQLGu1tS08W8QVZRF0nssFuX/kYIBHdaiMwWhXckE/9k/
mWeXWw/CMb7Woc4K69CGtYjXvbxH9Ehu6d2VCkN21O6ACbUCBytSKKdzjBBQpCbJKFX718x/9LQr
C1gWYPf52GQxZCmVCTTSOF+4XZkg9TVum5UBibJQngm/EPmHy7OaysObnBmE7fFbKkxQJ1Sjrh5p
KZQ2RitGvKUoGQfvj/Q9/aiG/tdyI4sB0UDjCM/PsMHe/7js7796rJ73aVaI9pdoy692PxAR+9Fe
marPgg+3hUlhHD/nDfy6f2O5Tr7eBrnvOM5/MB6aR4jttj0Xx1pxt/X6aWT605lqkCcM4sF54vU4
QYr65E+OIXgWUYdZvOGG3+IoMvnp1ZD68OmI1sQD0jqOtNqVvM32d/YGnPErwzyD3FVpxymI+Z5u
hy6QYDo5FO7KONvgU9YcpyaYmx519POecCH5JetsC90lbVikzsOqXxbXP4WbaT+q2k/sZu+81e/h
dgdoJJD6NBzBhGlngJ4R0ty62ZIJVzgQubxcXUza+1Nr3i3JKdyWEiGTyW/LS9Kn76cE4bj5O61n
uUHK5jIvPSYg1H5Ie1BL60HTg0rahicBBB2YjaRbgcvf98A0qoGyCDrEvFkM461ZWMiP0zhp5UD7
AfeGsYW1Ptqphmxj3Owqy8MwdBQzLTEzXql33CBqzylC8ayUtBv6S4Zvnybxzmav3xnvyctowqw4
QXcyfwTswJihrkoXtfSiO3OmJSf0hUXIELaDTcgQA2kEL4wDO6lDP1I0OXUITv7B2wZ8+pcO/MOj
bTTG0ypYSIrBkf8u+mkXJXgHJ2wjUXXxckZHqV4LjDodbIcQNIr5rAdY7NrRKZawZdj63hQ8NrPe
f7WK3UuIU32KVP31k6aGifn2pGPFOvvJznHxQFeRctWNryihYfPCS+ofg/M3jfLFw5YHF7D1plQq
nubYHVsISlNXwIR5px7m/UCneKys90TSdR9tN4hwnUcyFThVrdxrwLAcyz33R41mVKcTYsxU11MR
6xk2ulQwjOt+5iG/Ht4aTaK6Jrrs4P1jhm/1ZjsutxxSZiYqtfHVjwE46UVOfpmg8Mjr9zAPwqxq
dVdy4lHQu1ksSeyHZzGmuyR3zdvipOWnMJ8IbOve+tYi3VfMxtsBmwqha1D/8gEnCTA89GaoxggG
RQ44JM+U2SPa6aXfAQM5QNQPRJjZbYKfJGyNEggOpsZjj19kmoGWFSSsH7Pb2VDJUafMxsr543y1
HSDfrWa/O9FOgt0Y/UQhFIXTRa4jCFv0bu+a1T2TJ0/xEqjJHHyGtDjmYE6wmC5sABwKb1uuh791
SFWlzTC5ay5xsNItXB/l9XDQ0FJXzjiPE+UARxLWIrK5HBhilHGSQEaC7b8iu0pPMBpUlJzopPyk
hUKWvLGh+aYJ3x9f2JAD989QWYWIlcFKzNXB1RfuvwGcIG24PR/ewFROx+fIrgpok+idhDlmRQH6
x3Ml6r7aykkgNavf43GIxrQMs9Mpew9irfIfZRWzsMbrLZqZAg/3nAPFjNcx/TfAqulT2C/FgSdD
5oEQsovJdVOei0xGCd60yQKOeJb5hGWmeASq9ICQPKTsw/+l5YGYcmuUIqzGSzzUyJGMGxJ6wS1C
Rv4DVpxyRDztlKgPmOFIjyilIDi3Kc+Hbyoyq7cjB1OE0Gt91xlsM/ot14zetevlSqoWSR4UxLxB
vgus6xegtth7mZ+5MriPKAcW5mHNwGT0btJDq5/Qk9pRri9aRGk7IoJOt86DZYXXmojdJeLBVjvg
w6Mk0+xdRXa+O8tYBp9Z+jbJjwv7GDuD+Yvbl2Z0XM765P3m99jykiox9tZmOFBOkdnRlY0RKhkt
6WtP39TkYf5LjAatJ0GaktfsMXER/cQpU91Mrcd2ulOigUE+lvkkCqDdFi9tn7jkkb9zgjffajKt
mohkmK5AWUoqgxObV8KBFQy/jBqWmIk+E/mz0K55CszUXZHb5qi9kvmq2PXpjQIw4ZYlWIt2WDxL
HaljSgSHnTzPAK5LuXBWCOzcLAjphv4aJ3UCyfks3/bKJrFxqOg5uOIRh8D+DTEw+70yMymsw/NW
IXupzvC1snKDK4JS1cG+x88vx2gKBE+aZKonGKglr4Cle7zXGM94XSnL2Tz7L3ZtIusHM0IesD53
ielRLdZyt3uDJ09LxuI1pg1KV4W41aDJKg5MO1f4t+Ib2iDmiK3UNLWHryIOV0eCVKQYclB0RWcP
zsyXMiMUI8EvgS+QAhE3k5kq/qOkjj9P265WUuNEHuvmzyBnijK+t/ktCDSPh2hZieifKWtPSSxd
e5D9T/boqPWnmLQ6RWCbFZ46NAc7XNFr4gigh7OOthx7B6chfLSvnvwi/WEg4rqF281MeAKftlZQ
zgDgz7J3JL/IpJn6UjVThG2hLnzzxgsr72FYnmZJD9ZVYn3oBvoCa4QaaNukjiMSJK8WXvLG1A2v
D0sVIuZ7DEpoZa+IovsTuI4aiFgIuFJ5H7XbDehJG7DkDaGlhT+g8PXwKu7+zhf3AJ6z8AwpHnQ+
4TwpGMyG5pj12LEqsbVvYq+RGOMbugZM1D7vsKb1Qg/2vEd+5IiotX0h+kaDsKs1ydcqeHWc+n3x
cBlDmsoavXWQYe349ZPefY4jZzeKRmnP68h3jIT/QG6MLvMGCKrs45n5l31mVMpzX6lLiaFajXGw
QH1Ygq6qp9VnJuFMZ1BhHyGR13hBoN9DOiCsFWNKLQGnZpWWazxEr90UVj19XERYx2+bEEyCPHSI
/XKpnR/TpRDCTH7DlFEL30KihTcVK/rmR4qu3w4BIhgjSPGcc+zgoTtHPn1lyRW6xkvsggCaBwDH
TJ4sGzHNHzpu9suWMPmN5nJtHRxvmTY2/hbLAPdiTTOOW3MSIKGAKa2nI06C/yjdHjCRA0GwOOdf
p5Z6TrcoftT28idqhIMH0s4ASKTYK5tozFrKuAmxaZ9/GyibZ+jjObgXP6AssIxogd84hBzYnPpr
273kTSvX08Alh5kwTqZQc6CYGOIUfKowfOh17eZQPoTzp3PMX5m/OrGp9PuVuPUxPR3KnkA6lx/A
Y3K+zlN/EecY/onpmwoSTsnjGHkltVzbtZHSYW0x0Z5aUKEvQH8ac2Qh98HgeR3PrSAKiFGOWdgi
7Azp+RrTdhGLtIQfYmavHqTYIC25Sz6Zp7Vo7mmf/I504EqQP2I6tqRibSd/sM8aXmCt91dV+noT
Piq2Ajo2J3xElA+trCEOXb5zi4LaBPFB4//bsTOnQ48Xxv+/sKCj2Jsp3fLslPc5fA2CO2EDZvj4
6FFWCCfWe4ySzQrkX3W5gsx4/t0wDFQhbmedXXCkOjQ1FGAO41IrgYTrQ7Kpy0ET2PutEVxj/5yk
e6JXtvcZLaC3CFnnC7AmS+fsTNK0buSNkc3qwlj3AMuLurh7wvGh3igdyBekb+4mJLYPF7jpofTz
XDs/3hGSSGXWxRRhdiRIFyovE1yOYabWBwXwKEEyFXeUZ/LSo3LWE0PiHO+SbpYF/f++8c6wHelT
+TpH+32NekImjZuBOlfIxpHXfSB8Qu7tmOvdnIzszeh4ur2MDxDxReIR4HxZJURKnEFpMmOICCYD
G2YXqPm4EbxyepaAYiOcoPY5TinK09Cpu4sR1ACoYO9tqZFy9o+Gadkf08rCyYE4LfTstT5HPnN2
pvwCakFtbwrZEvHAeMJxHr13t2jYbULw/j5X9FdBfkRv1F6rC5oPPGA75UT44+zTy9M8TuT07cpY
QjZTGzk2r8YHG3rv5Op9naLHEHJ00MEf8DaZjk4yg9TlylipmYL2qS4cDQR7AQqbQwu45nsg8HMg
gMy6iezRfviEbUU3FVxSJJZR0mP1x72mY7pDq1ZhF7VyevV1a8QyfV7FdHG6S1wSAL89ozzCQ86W
LIhK3valhyD9hzUjFZRzJ60PD88yJhKdGzWRttDTJKib3BJvs4fc8x+KggNSPcd5U0ZESLCpPedh
HznoPBeqmZrq3sFs4Ald/H+Kfah9UlWjbOkga1MeABKh0ncWzRWkfJixHSZV0rnk6PUPaIFRoWPa
xMfHVuu6tS2iM17jwMbfUOoQs8dXHorDkkYDcv67ptepeL+Bkj8vdTa/kglGFXN9m9vjtpOpFLMl
8XQKwOIMIOTv+82kZUafEpQj12rpRbw2jvl/Oim3xN+Dwge2+R4h/qU62L4pvGgEUlwCMGVZgRc9
5RfYEP1vyRBUS4VTK50mevQiTzgb6VqqXJ49QIHxYKwarS9Et4IMyOyshKAJuluTBFLQorVs6HcP
dvZ/xJi9e9bAbVg8q2OpidIPtKKrjiy7fdu7pOb1MCVtUsTYVIKR2h/dglvicSIkYt9/EszorEff
dW6T8YDuSmC2tyfxKRZxFLGSEvgsAHv9sahzBb5ald9ks5mkpWh10TySEEzk94KvYvu2J3u0VKTn
832OLClN1/1J4+xwaFP/X1APEGZOwLgCaAYZn+5OYNV0VusfTYmN3bSuiY6NG2tHrm7CUX5MRwkI
L21aA/pI0uilJ+KUdQ043SegyiWYgf2BQAGbPBCnwlrLtxtFguw8mhhAtyVO/O8OABhH7p2D6Wkl
MmTP9RTJMVoga+CMx3JfRWIjwOQkMkoQ1BkQEjV7vxfXLCHr2e1dCPfP1i2JZcHo/FZPWyU/u4Yv
n134RRDYOTDV4EP2RBOo9/WrcwSOvKPQAedZd0pJgMTeqKHXpKbGsKIncZojizKbBp2A03fHtVT/
e6ER6bLbn77qywNP3hifPpoNzzjBlKlXn/1vhcxrrKfYnEbRjnQmAazpHwPGLN6GFYD2suEVNTsP
Odmmmk6xABeGm9XPPAVXWULztScfGVIGiXSTxl7hodIaC0+ocvRrqzlFlA8pNYQG3AB2/qK1P6Cj
M01XNDvPFH+gx+zzoVZhYM+908F8R98ylVEeTbi0L1c58nCKuZAn5LIl1r2+F42+PJoja5n6pz4d
qkVrF+CI4BkStGuttLURRQdiAinjysZsREgExcMBYzHcWY78mgoGcnIgImmO+FAMEszC+Oz25Khs
U9wV+2M090rQj2DUdsoCVMFLJrGOpPWo9wNJvwzAWHmZnloAFLICJM7O3jQ7huH2RmVczCUurwRS
CS8UIsB30tJbm7eCpTaMOOcSaLWi2s4OEw3syjUzOwkhLHb64n0gAmloveSYBPiR0BJHrsxRoqpO
mZjo8lw0Ajd5ij9bzvO+NuyOS4CVzL28oFqmWEqhWqR59r4b385jY+8bdABtaGZYkSF0Ta2rCSjc
Qh+QOWDxqc72VRxI+LU9CiJN84vkg35+JWdSFph+Yd2v4xVLBSaYhCrnSjfCwT+xyveTVvvhxCb6
B7WX2HnnLJYi4OmyjGT49pcueNsisadr8wkgBhsGltG8t28zCXVpHsQDf0Y6pFkhTVLIh7pz0BjM
KRZNHMwa/dNPHBMP581Q4YAbPLOVNP178usqDGXlalnyDPrv5FdnUTDcSuHFSGK7LH3x7iKruNrv
/5eWsFGTqIBjv1y+Jhy68Zv+hRornYbtJzBF0Kg0lDvWkmqU41lvoAY3zoiAPeSvE58RbQYIS7tv
UpLZ++GUd/W62LiQZiZ/sARuqR5mEseJTRkH/OE/DBWYfOONSKK0wi9gwhRUb+Uji2m23pBSQ+Qe
Mn66vNMg59mIa4XhOrFzlbsxLDI4EFxbLXE+e8K4n4j5tBM0359gftz7mtUDFTcHOEnOuzIPmfNx
q4zKxkTRBSr7NmNcj/9PI1xi8Y58qvkdTJYWVVcoQs+l+Sgo+fYyllhOUC2qCXmaidKk/ShwO9gd
lmeOFOHPR1DF4V5L7ScQmkstUVav31jsMe+dLXbFPbxCiEKMRwDHqhodjxWUkI69IL2Ke1re+lZY
0IDuA81RNrInZHH90i5FEuNfTVbcyp/p6feTFrQZbx3HDsGSKgdJfJ+PWm7715RmEMgFlzK7Zp+M
slSUPDwNKOY/3De5nEWKWOswxpH5KJHpEYUiXKc6x0rizfQZ6ckAaM2fqY53n/vvNiGWl4zCqUs3
QMnTvp3SNzBOoRI7G0DJaeCoaWpwb5rcRm1+6BPoYF+pjJwPkuQT6kD7oC/68UO1JpAquLCNLXpa
HLV4NrRT5jvlY0BPUEtOzqE5zsonFz7thBOZiD5X9lx0RxJBxPZYtM3t4y+CmabvitrH5e5mk4KQ
bVd0HdQgO4ZQHZrbYIhZg8ZoJduhUko8V8W5Dl2u6YfBINK3NgCe129kdj1L/CTycDwbLZJzusH2
396e2l5DbStrAdedFbn0ZFTYTY3Zl4FSMSAmKi4FGIVaY6ztZqcM0MqAVmj30NbAA24iYPuZfalZ
aqQBdDnWakVigXQhuFNruw2AqUuCyrF3LAl56JKp5AR9KWFBxvSlHrCU/NgLKAJe5GDmodGy5dQz
MCB+eyQASafXG+S1Lj9aR3YJ+p5Q1szzSTuJTMp8RVOMZVPUD2b/wZJxF3Tzjagg+iQdJZL/D8n2
mSd7LqQwfiK8/xCdDZOBZOEnkRNBp54BEsG0BWxp4I4GckiM11oYyeFNc7HLZZgBdj0uZHh6hO1D
Ns3xu4xMwOoOz696yLbLgV5u2ICgjZQCn1Dfm1hyzKEy8kGtEL27JH7GbhNK5WgI9GWoscJ2ZnxK
1wBIZnk8i22/1H9BEusZs917GFeOfyNgsBYtK1kox7cYfA9i2FUcc5+FpN9jnJsN4duWR/dV1mQa
q/JU399DnTXjRJtNqIFCAxoI9TL8FWthqhJfN2d8fKFDqWJPxRidi+Gh5oNd6dr1WdH4uQujwaaA
6vThBhhomrYJBAJMDDzHTjQyFfG7/4cQ+FwhBQp83mTQqUc8wCbLEEC0HbR5AdMEK1L955CfgS0h
MvKW63ixXQdIryk89Clxri/Zm1v/HtKKS17P+ioPJmN9DXwV9LZHLhlhFUAqRGndOqqlQD3AaLqM
aeDx4t3NLjFqgGVpKT7LjZodneKc5BeLnjWz99gzVe577doZwINwAyPanqtODc2YYYW47FMRwabl
W56S8xChGjO7Q9Hzao4ujNQ15JXL4psSQxazVYDLN+O7YOZgS3LPuRuDys/td66U5AmI16/+h56J
Xs+kBTVRFUKdqM/xdez06KzJatoWAH4H7s4oZSu9Aiey4I1shI/hapmo7x6mhjRK4cIAqEDvjblf
ZjdhuRCnL8lBpOMn7Zuz9rVWXm97CFrEuAREKqPEJ629x2FEvolxjzv43uJZ6IoAZth5C8JlMP9x
X/X5FPnVIMKZfGni/QCjrZk81E+05pnan74FyRE/yQjlCtkRs6ZCYrZnHfww7dMboNcW0qbtLnz3
A2lwRS+Qc0IMXJdGAqBrjW3AZSjKrj9l1hgIrjjNjtfJldmYYvb3OS25Ft7bNYQ36MnVfQcQ6Ur2
H28Ozi0ikIJwHSF/mHGAX9iAVPfEmSG3ytazenU4fI71V7eElHSdrFcnyXKAUoE/nS7QA3PYNxAi
pssFZjxaYRrWaUfnBKbfqXPAwmAclis9W2zxmbVLP1QI4utJfIG88vP/ttsSpAzynwrwGHs4OWNP
jJPeKbOQdEnipfY9H6jHoWSgToXYk52IBq6/RFGx0t4WmtiYmc3cLsvyEkCqU9L8cUS6C5JttZL6
DDejJCimJ0YGviHDcdWV30NHdNvaQPU9iZ9F9N/z3eRb7fnV0ZzODMJcYXeVNW1YSSv1iFsmQl4V
TGiuZpq65Tb63yRQuqQDvlOzbFE+n+26K2cT/+2ATxIUi5ngsIFua3A39hWsaWxuYMKR8g/Y8b+P
Xa059zTSl2qCQLe7sWSWrhx6KFvAr+82opuymC7ai8JenXbWOXBkqg1+gRKBHpxDsm22akhyQCHc
CiWf9ks881eg/V3E7//76OJyx+Tr+4N38wuN9k5RuD3rUJx1oDaOUxwYhJNt94jGbe+FJ2E33nlR
JTh6UskpYj8Lyejm/wJzY5EfCUJqlFWZM7ioawGzIhG4LEBDPcRIHVVMiPsNHllCnQhfm4xviaU+
qYWxdC6OWbipqhH4WVdHwiSyVfmIn/F+9ty7mvSYXRCk8AdUlul4SwJ7wpjkvih0blvZ7fQc0B1W
ixkDmyXrJySgqNmI2Pbq2P9sQukruQaOm8Q/wt4cszIqgyARxdrtSUDSzXLuEnluSBMi6rO0m2PJ
uHKcAiXCHgeIaO5Zb2eHzPwm9Yz94XyxiqXDx6vsJZQ0EeYpO7x+j2Nt+dTe5hZ4pMX7nXQzyslr
w3jct7x4AUlwbQRpiMu+qAs1amnErWckQqE+HF/Bme6v3RlMc3lTFyyYxGBT24crRjE+W1Be0xCd
YucSU3dc24f1PGcp/ezZne4bIDCZmL5SRaOTIYlhPfVBHbGtaOQcHfJxXYR7+9Q1wx1t4N/zBML0
fioYKOMq9GHv+5xo1xbaJ7c8nL2qQSUm2SPCj1d+wikKLXKwRzyrnoaL9JgagU05yrWi2ut0ReTF
TBvQIWsvWADdVXJyxnrfCeXNc3SwOT+82npDu2lMPyaAfV87o6yjJSEULwGgkQhZaTIlW4CO5Ffr
gGMVgrDjIcRqYzptqrHVqjqrU0DOTlLAFbgp3N1rJfsSa+hrr3GoHNbOgnLr9jgg5LQxP4/6tokD
ZZkkHM9QG2FXb+wbm27i6qLmaAw56qAd34tv7Kd7dJJmHTfb06spQMPuTuGTK0AM1ghPxEG2L+n5
6lyFeB1LWMnLgXCgQ+ky/01FpLrImPm9YcND5pkBRK1eqedQdvn0nJrsY/R+/RmoL/czMTbBMiaR
jWSic3zg8vmHvUAMFBjQqv7v5/TThcVDyg8BQb/AMqo+DSqouTs0GDnmtIopYVPqd9WWptyY8SVN
8kCvFEgvgzKFkkWSDoM+jilTrM0/2xqHY6qE2NcIJ/EylKq+V7rICEw4t+KuJi77coRX/JQRzYjR
54XEan/HvyVi5TrKVk6Z5+/cmAcb0NnxiQyUmDT0ELrfkvyG6EVbgaAXBNsFLa4e5H9sAnK8soN0
eDvgmQrRA2wZOpXQCbX+5Gay+JbMhzriEstSkE3G/wNgNNRqOdMZ34Po12WeGKfuyz1YGESgCzL0
RYnW4hjLdgHgXC/uk6fzl3UqhJBkA9ydvRZ3kIM3HAeJG9j1vcBX3lGz1PRVRbKNZ90cp+7LDETv
GW9T1wJOJKYeSrlMfyPv1PO6dAwXQvwo7oAk8DpECOPLxDUYNPlRLAYpU3Jf199oyL5ChJaDfe8P
OXhELxhofp0V3gyMSkjqJ+svR7252bBvmXo+T/wlxzMf9YCa283RfjpydW41FtiGsjb94NRw8MHr
eQWpvG7v3DvGtMubj+15F1PNJtlOS6LGnQG2PlZ89N1DnuAI/cgvG7u6Qebq+DqbH6ypY2whFr8A
EibbAqV2sv5YdBcug2BoY7at6gkgVMTznecy7s/GWA4sZE06Gxilo0mcwNI/mFP39bs9DteCwGH5
c4CcXmswVdznGQZeGPK6qkPAijZAHTvQc9pxEDJajiuKihq8DU85x7vbGjXshgerzZmBDj9Hv58W
7RgpWYsLKQW0Hedn9Wskr5TBVAGeC+BGwOXPvl8qOji9IlGsQPmnINwud6NIXihk7lG+5CMPQlCE
EsyBte1nNL96FoA1jeyWjq1RNUYDjhwXdy2M/PE129qzgw4ENoYJHjdpNba0T6Xr7jFwWuRbe07X
zvS0fHv1cT2Povh3m2DjDcYbswX1vHJIsOM3viYmPK86zIcXhPJyE56yg4jz+qPwsgXtmvnOLCgU
IqwRIrx0KmgOKEuxfI9q8Xiztq1F0o9pv0JuXpFcUlJ88xtjPqHtzg++Mw5sj6LP/H0PqbYMfuX4
TgsCgX6rGDNQXFZIBgDXmnQt5SQLm02J5SjmUJOZiFpbxLyub7nQdSS5PR1rwhH2nEx4T1+9Jpgu
UoPQCyjh9SxO360wWFZENYrRuGp717N06GivWJ6ZEMAhFHeJoZlugQT7NPbAaz8YDrxjKnmd5Jn4
8uDCKMWRZ6zCHsxl3tAzMa9lFA6y8zKgkKYjWNiBPwdwSkKcQSdCnmuunMNvJNcAb6U1/E4xOdH/
wjdzNmdHubDKDEFqwizXtdQlnDV7Fjydj77oxOFp+SCUlPN4tQgPUXKQP2fc7RTlaHueDBl5kquz
Q3DbkQSdMlALbdE2lGlmSThZ+bdpfgMlVkXJs15k5nQ5HS2ZzgnUt4WMbf6w9Gt4aPmXYq3x8ief
+UQX+32eA7z6sb+nghW6cpPsFF0Jr3wxzTnpDb+/2uSyZWEEOPmf24oHt43nI/PhMoCNmuBwRMiG
qDiP2s0ZnH51IQLE52tcFRnHhQ9C++J7iO6ZYEQSt3qYW9jhcp1l9FeZvLnLblV0jQ5C1T70mzl0
BmcygxD7NvJDbNxl2hOvdjFX3ZaJRL67Vjo6gyP3qX9Nllh/2Qz6jehfxeru3FcdcSPFTAGsutU2
88upWToyyPjc0qdvK4Tah0JA6UFQr/S1sBepDk4ckJbfyqyy/kduEqEb3S8hkziXm0TimF8W5IRe
7N54sfYzOA7U527uuD/DfWJiZJDh4/rSl0nkxR93e3vYjMpHRs5WyT0ow20ghYs5dZ9tq1qFyJFX
eF7kDkUn0nQLVCcYxGLxgIJIb7jcRh9zH5cCVnNrRw6D/3TLJpIGZtKimfJ5BB5kRQhQbh2g1Y/N
eDmUO6EwSW9apvgjalGljMHzUdik0Dgc+2TQ/79d3bRo89hPRvE6AxLPie8W69GXAq/q5XbvdXPf
lvReuu3QAb4qTC6RVgtEegfzJKt/R4TQmlN9V3CDUVh7BFpsfqckZyLw2KW3dIRQ++hyC4ug/ipL
ybNjObaRIdnGcbrqA8qjcDTKtMRY/hcoh0qPKiU3dazvTPkNo0nc03AKCzjkmC9VFYpvwCWoZm06
INwTrt2fToneYvRdz+mUJdSVYaebZ7gNX+jJ/mU+jvYVLPNdVjxFvbF57rcqSJ0S0deA2vWdxtpf
9ACkKJiwlN9S/j71M4d0+rL3GRtkd+IQtL9Mayxd/HWRlJnvNAf/c6VhsP3KQMR/5VlJ5lMHL277
rjK7FoMwHSqctXlugOHIVFazEjXzoHImQuQtrgFdwhtf9+09iwz4yi4JGdgSgm/Nb+il/UCpkTS+
jCbat2xiiS2x0wspzQ9vH6atUCCtGclo+FDXtc1CmvMh++cgGMOnU0LoPMD6oXxMAvhHNBiQuzgr
wu0Y75WgltFSvVL92a9Lcsl/XR+6sv9ooV4QJC94cWwK3X8Mn50Anur+aFoJ5v5Vp9mgFmt8Ymol
3A//+vsadKTxUYdzzDCoPULkmQLzK2ob5AY4wZptFfEYYkZpnmNf1TxavfjgZfhJRIphHboFI+SB
70/+MpKvQ+9tsZTUCWyaY+PqU8J58ZsEh+PoVjKMyxvANU2lXjfTl0dcq+J68nQO7GZBflvPEyNo
JennNnAVd3/10kVJAMPHHVLUDo1ZJ9A79Z42jnwgiNciPK1VpFH5O2SW9JreDR46pE7T4wmgngUG
rl2sWdJ/aZC2fJKc/t3uxENapDxq6lFVOAxx9ZOmv13ddvKIUQUQW9WpD89mObosK6vJ9uqR6R1h
23ky0HBwdDbI4XelQ3uDubJpRDaqe3Ys8S1wyAyQWtQ/GqI+cfa/KCP9UBaqjd+eg0oxgm1cOXNr
oR4XDgtesY28LwXyPzc/jMm2KOWJxDeQREcuObpvgei+y3CyNXlhjxU1cg4ZrwmlOUGDmHR+7n8m
d/LRQvs4TByuwJlowZhaPFnOyVYx2FUszwepq3Wl7rBxHVobuamfmtkkVMYr8NlJ2/msqoGHcj7D
r7t6vfEHKrIhGmq/u8yr6/B2Qk0KovH589YTkJsJSjGsUPitJV79irjQa1Yiv5Hp6HeyG/2r+Xni
exiYXONZyJtJ3KeEijV/3MpHTZBjeq2hiHNi6B340zW91CnTrFbflTDQoWkF2w+0TaPBq8pJ5EzM
iUTyIhMXfyweVBOWSHwFMjfZrNQe6ttUh1NXQ3bKoh5jYKLgoZm3LSsmTpVVt/y8qABsfbUgKoE5
jzjcYlGYvBFZchxzWTQ1uJ8OgnEfJJMZMuspjQjbPkrTmUwaXgyHj5HN9bHK5OZiSS03UdJMklaa
7ZVUAwPKhrwVMVytMFBhpe9J5m2a08hODPG9xXoSzIGjAMJI/8ygEJTuQqbklI3+rGwut0uAM7hD
/gg1C+kLKe5qVce3sruTK2V2mlOY5bMqXxp0d7lUEJietw0gyiEzufTFdMi9TFV1784bkigv/sae
j/b1OkpNxc8HJcf1YlEESYdqCOo7VrmdddMtffyrJBl/QpnDjchfxyj9Wu3j477Y4Oc+HD2RY7zG
N1SJm9mue168W04WR9+S5n7LE9H7qT2hAZzBS0pmYboox6TMn/ol42WTmxHjTfIknY5xvW/nIjvN
HPl1FYVw0qv8rhhVYWh2XIMelv9mru+nFIH67xJKFKtL0RXA6idUTv4NqZOSxzaLpdhia+csPCku
4yVrefBh2ZUbDieb9Z26+WjzDx1qdG3qqC4ZsfhND5d5/9LEQHkU88UOLaK3hjY5ROySrLccYkUn
pullW96Y4B/pMk/m2H/tSN0pd2zIvhmqYXJHeB5TWiWqvZdYne554X/P9lobNs4qOcvdIeitE/L5
F1tyhPHfs1sE728zLj+udRMSTV6L21EFJQ3GIeH9IO8XdUDb8rTKRYPKzshhsTMeLI/lZjQCqAxC
jUyoMhtZz/bMQNavYdU62Ok1oQ8OOFM0Rrtt6Ja2Fzi6dkfLvYHOgYN8sRhlagCo95vl55DRK6jf
uvvMuCbyWAs9STtz1AUESNUPpaiOiTFN2nq/A30NdCq9c2gMuSuiTBFVwAxXL6KFLqHGhES3GcEA
z6vBWJrcC9GBW4Xdneuo7vdW2c3u6nXzIONq7+wJu52mXJauwN0uQd6cDtN1cURtnnfJdUNsLYLA
bqLy4sFnMx5Dg71m6gsZea9k5bvQFqdOK0RxaBjfeLJAkXN2vuSkkfkzdLhltXY1pFj+vqCdziZV
vmxDwfZXkeWJuPTakaFhZO4q5Yg0BvO/WQPwoCdy+zXDtA0qWmTeqhDICIZBvQrKSJc2w2mUTMWf
H0DvtBHjHCl/4qeBlrCG19imf6zdujL/EP1vq7qZNf3VPVfsK4tDyZhVA8Rdzilc1QgRRMuhqN24
v3joEFfSF/oa0WK731ABXhuV/XBj/RFfm+7sNxyb1aw2UDVinwPNLW5bygf3R1Ub/MS0Z5r2bkJL
VhoQmdEc7g5cikbr6S3EaE9bEl4gy6l5wgL27ZDPC6DMF3zKKuTuwTBDLBx6kItpgp6DDzqJ9lVR
mT1CC2UqekaBY9EGndgJybRC4528SJpmHb+qB89bTYRKlhQVFz4fiBOBqOkxfHN1QK5brlGae0vi
xDlwXNmetEZBplL8pV91V2dK/p+cdIpE/N2fcdyvQlOPK6X/YqazY2N9CJ7kxnpGjaJOCVBEYv1J
HGyfkSll4zm3A53Ynacijyu4nSvA9vOv+ITyJmjege/G+gLhssooW5pfaz7DGXYdRmUmDkD53Sv4
oNnhFBVYtrdakAk9OiDj+nRvf1ooNdclce/lYAq1KmJ2KMbOa/NKaim0+0rPaFRe2FWaybYuQB1g
u71DwjoZ50wvsZwlrw4JVbskvzdRuVxY64CLl/V9BMMEQj6qVZG6iUaDD0EcZOIeGu5DoF9/sii3
wpKtUQ8OMAUKdyg8eEait4CJProQv9ipC314ZIhqTWHIl6K0Ml7vfAKAhGSWNEAvD+eAZSMTj+PG
4vM8TbADMzaxHHkcyuKsEgoissydjp/jlxSpwx0j3Jn3nxeTdici/9P0WMlV4IrdkEyrT3TlSrDJ
5tm2qLaqH6FkmJEAY7wwCIe4urmUSM64R7l+C1fnKmHpqAP1sfSU3TOUNvaJSvRNEUwYgawFpTnY
LqlYMOvn7xwzex8M+5awa1CCgdL6uJILfG0UpmZ3NreKu7kOYGoaE+dyuh5sI5EC676UGI0W5G1s
VAYwKQuJjP/fnV/fSpG6dzgvWQvCxoDvzHhOz4vwplAcDyNzKOgOVU7EaV6tctGzXy8eWZ+nlFug
vFzCeERX2M5J41vPYhLhm1H+2Q2JkFxbul6n1AmWE4XJKy2aLLlBPbNAklFqpb3uSuiTbudwI+yi
FgyXo6a8TwD2vVOV9+hYHjoJ3R8eRyt23M9os/N6Dtl9O3Trsls8gTYYHFbIlnz3/wocFnGRF36P
CELjE1sRZYH4RSSUVEFeUK54eoqevSJlI2R15LurIBA7YgUWGrloqapCrr+KikMbiGdxGHwevYbW
TNNRvdCIoGq+JTwsKVswHiXgvrDdvJcZLMNhAHceb+bO9T+PEzE9HFPWcKNRHtVUalLoXBjgMRi5
Wxu+vaG7PsDsSqMIr0hqKUHXE7JFrBrphzR3KS5oI5ikkTn28hEZgC0C2WVy4ptSEu4VjGynjnbU
hsUtcFKSsbJzyXSvahQ5qQsqMwv3NWSo8Y5ybHvJi6gb+G3zyOQIPGLJhYHdUg93ABGns3Tp7C3v
jbdBEBQketnszLXxmXG1quopjt9tSIc9mcQ7iF3VKMkGvzzCxvoZrR0EY1Pz0cX4jk7pd8iggWmS
RjddhBJG6ekJE54Ulfst8AOAQdl/JIbztNamNZ3ABq8D4oCEZaB2UlQgZ9VAIg1d8JIhCZLoqeYE
BzhoPFFqHMJG0dQmM+McKg/tdVCXvsr9Z38DTCOe65Wj6L515TgHHo7bfRcxnnX9RR13iKra0f3v
AZJkPb5l5FKLrhysJAzLs9nJFudVvFKGSlTTDjK46BIywXlJvW1l3+cjMvSWtz8dk1Lutq8y9ter
e2RGTpX4HeINn2sbBfaMqMqItNy8vA1OmbQHiKC862fYjvluLpIRzDH322WvQPuDiZ9mNrm4FsZM
D3kqKCdIBsS9Sow626memEVdocLwNIDDiuPYLT0KwnTnPKn4WLqkxAvFQEQ8VJRpIm1HLDA4CybT
u9Tu2sJKlGKeBm9App11EPazXs075zIPJqOEUVGXybPpoYBhOybXHhobaCPBq26L1xF9dFka81h7
sP14zze2ixw/8kjVzA2ttEweiNZ3JVxV7qwVJRf3ra4Oc+d6vA+BQED4mL0vWymwVj3wr3X9t7Rq
D3kpS/4rw+v0fh5jqrwLRCJiO4V5nFEnv/LokT9cipQ/MQGRZx0ZtYu7KHS+geg7r8tE8XNsoGbQ
sWvy59aFbZN9AwslwSG0ZHnUvQ1/0gAZEtr/nOo2fo0tmZT6x9sWb9eEN2JOcGy0F39zx/vXWNrb
Cup/p1zQp9kaslbx/YOvw0SFAIJYEgRYGctVsPS0e9c+044yoiKiscp4n6/UKHfjV7bGw6QiXMKL
qPsA9uG7q5yVVxMwco5UA9IHANmUbklaKyvuXB5aNJN2BH/TUPdmnPhHrcI+LGAZyIFse8AGlWuY
1mWQvhOjxYePRUOKsP044/t6/pgyAcHnZvGu4LWede+urDNn62j+kN+N/bKZEISeoRJopGmBFblb
huRotckQaK5Zj4Dt9L3i5JsUr23INJ8axkkjrzp8n84yE6VxVD5SG05CTMpSlPr4Q0XfLh3szNU6
OnzSne3B79AanbvwvZ7KrHPUft3dakpcwdY89+zNNIn8oG48pgGtiFnbRossUVQK6/FI+tfFJiMZ
zzAhRyYYFXvUaieQZ+qtWhHEkxskflunb67QExhAFLweQYsnlGDdeS2ayno2QDBBf0noUzzDdSES
cBpNh2RDVeAmFhlMZtBEwfi33hqw2AgnCvfIvSaDuvJe14K4siAe32uj/sAlT5TrYo4kODh6J9gm
TX0kI4K5K1ThuKnsoWfGfS3ccBMIoxssWXnpBOe5n7HspXr8j706jkdsfYWWjTuvbIss2ZllSQl/
4xNNqWldADh2cHRtW+kcSa1QphS94dC83JowgJ+RHjXGQAtVuI3WnCmuW9/qB8wOyc6C+F9Cfs7L
VcbLRvWqdsvxjPlCMF14jpWndW7BHabPQscADprmt0esLlajC6/nouSa493QkyfTpKP7l5o7go7U
fQ9zh6Y4w2xjkoPCU5mnFTP9VL0MYUWkBAysbQAIkyvE1cgbdtceU5hTUgcEIat6RlWLl25z8fBB
95o7qpAx5ZaVIANeXqsNOLLXGbblcf1kotz8BFt+/y3Zznir4Z0A6hnr7+git/UZadS+9zeDV95i
GynQskRSeWRBm52pWUExoqO2Zgfw3intJ/HS7mW2GEitb6UzbKFNN/5HdHJPYVgeDoO8TyJFMo9q
fJUzip5V9dLiwB/sazluVQa2cB5y1+bzxyXtI/Gi8HsSqSKvU8W1LhUo9q71w4fQ81HNB4TZ/I5i
h1nhAvaQXMOOHuu4McSBrvsukFYVeGqnjngRufAlw0aNncTbs8MCZviCerpqD4cPhaKfx2QkGc0h
/r5TFIJntKTrq4pn9RygidGC7h/a4i0AJIM+QHURRYCxPUvqVGsOiOxgIV0buJ8AhPyktA3tmWRK
3JQOfFZwvfjvpOlefr6pmyNUjTRDPKb2FdY9Fv7B1fVLdqgesD6fhPEGq2vP6VDLcyu++MgxJZP2
AY50dpKNA4A+SPQGjVB6AvBMiywOSylziQJ/PCwNPkO/vY8G1diBHTbFH1G6ex6p4bT11VTUr75H
ufO6eeBYnMXQdFBTw1D9pCHu8EuK6B5I9IXfAg35MvzsJEVyUYktXxoT5q3ECn4u6Mx9/IuCGBIk
LR0WH1EvQ+bjRH3CAxY1/ZUa7cxBCVFwp3+sDpjxB76Jek1LoBY8fvPBC3LE4NsLJalI7npKYlkl
+zOMxa7RwLNdP7VUDwNLtLvmZ+/4J2svIu/1pA+GxCRCOKDuUyzfAe0DKdKn7qEMfF8B9wzPsYPJ
b6foVDUC2wUHy+6EN7SFaawpiXhvmA7Ot9LbmjiXEnTSo/OBqdC39uBc5GMtGGIRSDZnvqai2U3/
LhcwifMzauM9fxoWeE2/EcKGEBFqZ7PhSIol6QBXFmr25r4VFbO6FhcPn2YlrKIO3jWjgwvCFCvP
mtNGMU/P6lgn+eDsBvf/t2B0154ITORrL/2ZkptmW1+mbegYQo4m5fdjds4ghNuiqhL0oJicjV58
8RvFnJe3Q4jT71+9Kj+KeMKLa+woOCvVXnYg3GOG7DB4XvohAKHX2NLA0HyX9+1Z518A2IPFTfWA
4kWpIYyMlHYOmP6EwHZpZq2qNpvTkAkiGWU/cUMHbGIACC9jRyK/Cm6g+B88oavG11s50THcRuPt
avYsJVlF+LZkNqScosdgealYAc83q+oyjZd7M0OUiw9wZhAy0lPpsdiL4bcS5FbrNbUDK0Cx0jql
Pknp3uNEY/tgVOenLm6iOvfsblwhWUMN6ULVFNB08BDGQ3G8prECqOZnTleIDUgi1WmEUauWzX7j
/6/rLsZDhmxRamF4891HBBTAyOUBdCs0q01pNbGMND2BZTzXMhqzN2by3y+2KG9cK2vp8ZUNd3OB
F9fjh0FCPKzRqNTRl0D+A0b0vr1WFjSLx7TBOeO2n/1W+3J66orD2Io2u+cufmYVEa31ijfaMjnN
ArBQqKk3wvBc0q9njK49ezCiqMJ97jaYOxCqhlrtMUxr1xjNFaWqouDyQG5ccw9A2OxYupC9D/AE
glUPGRiBthBdOeo3gxNgMlB8q6KXfrxBRFAe5KMm3b8XW15Dz/HaAjnX27rTqXQso00DFf6kb2tT
N2XC3KV8wtU054oW+OlMcvLS8W5Hw00Yv/Us/QBEiBfLzfK2FHaEHVYV3hbA+PaOtUogCqjh8wJf
byl1Rysv//TZe/oaTfPg9hx7WYIonwm3TlaszQO/YsIarBx5q78TPBVXA29QOq/pI2xD85CAMdnG
6PXHtWEfACTgx0+CNRhlmnWOSxCNwRqhTkNTpA9JjaKwZ3SayeqMK8FZJLa+Ij6/L70wfq/7QCFb
A/anMShlBMa1Jd1zRUJl1+lLkikUD2T9n597ZwQCeSZYUmUoiRxDQK9cqoQ/xx2UorRKCDc/dmuA
nMgsy19k0XvJBCxO+wwdSs8zT98qcml/AEALQ4lVnPWG2UayMXXX0iOsq3XVnJR1zFxEUM/S+5B/
JJOlFHHnhKUllvKzCOq/t8EsTKO2flA4BytdgAswPAottiJl71IJQTTIOg2BZacQXEi2DWVuJgs4
F/DbezyZ0ROPY53wQ08fA13RBRtxm0k05Rv0NbzXYUXviNJh8ko0nU8yvu715X43SHG/0VJgqqXb
maHg7FVxazE11Wa+Mz8/S4/6lTCa8LcmiLhatFrJSqLSdFJEm+1mALdTCdO79GIOuQNs+DgFHBq6
m2o9DtjVJBVBRbQdClQVz+ghp/MgKxJbl0R2i1I3MaG535OQYuEHLdBLjIzvPRdcceZ0o9TOyXQD
sEZJZ+o/cv0lWRrRnO0VPxOdXmcg6KyqZ04vayqctMuShQbjXpNSclS/mZNooN6z5qvOIId9JC4g
jIySVBSlgjQyE2C/0LEXCIvgBAWw0y8YpDB8PMvHGzEzwQj7uAfnrWjfOxhztZFv7JR1kyI/zDkx
LRmPOu05whBiLqrOg0Dwb54kmyNPVDniEGeC54UsuCWGZaXHa9GKG31OmeOqfzf1bPmtoB12s4tx
gpZmDuMkrr3baWV+SKWfr9NYoq2+mKrwoOjkFYjVKCZjdoxKNcR0Dbl3Vwr8OQCKWBvY+5Xbuzon
s3JARXt2GdQd5WrZlL2A7LqNGhSFjfTKjE29+WZQEgZ4xOjZPkZdk4soU4l33XbNNHHXsk3wVVcc
yZvzJLG9zCtPiLsEvxZUIR333qfhOzc6EoauUyM4mtNu5h+pbfhxljQSujZFwiaCXVXjupf14d6c
uuxwCv1klCYjctfnELRzdCua1GyduRcnCK6Dj23QFJ2ltaNYK+5Hr6Bfh26haj0yz53A8oTMFwra
q/G4pvYst4yXvUTK1r9bknra0Qi1x0/xYNc9CqR2jnz8X4xTByU6F4typsrrm9rqI+seBy8BHSUQ
zg91HDX9gXTqunAb9Xf77a0Z4C3oOh7Ax9EK0K1TfEh4kLgEY4EhOLop4fvYdmUrWDqsgbpdrrm5
EgwapV9z7zpC0hr2JJSZ+SiGpAGdfbhOvq9dTHHoQDF4urHj2S3CMMZsr6Pr88mcx+XRWI9Gcjgo
yRfZELwRW82Y/uvRa6PnY6FIUFN9t8Dl+fdze7ZAQ25thKRVCSae23dNlUBExhq53qOytIUSBKxh
AW/RSlOeVU8LfcQVA0vanCcj/QjstQuvtUDKVx9JAFYFl21bH8AjhiYACoOr0m6s2WxWtAbQPijK
VkYLtmIIiWqilTtoLoT3irK/6iA9ZdulJRd8f6UJZGV2/IqAnPcdgIKLpSNmwzM/l5Qrej6aP4CT
K3gLQGBSjqmCjj7QWqaokA5SS9FxHNlT1QBJtlo1tpi1f1H7FzP0JDIgHq7zBrD/9QTlkc9WYQvm
/a3dk/aVn/D7BxX8oK/ZcQweHUKIOV/oMVg1PnGVtpeBawcrpp943jdv4qO1ZYWve9Jhz4HwoxCP
JNlNePdie7Sv+4/9UrVB39jZOkn7hIkle8b4IIkbDhmFCcgRLXNEFQcnXUzmkfvi1q1a74AqDIJ2
1HFYNOARLz/L8GcdgiPBxMWOHqYnNDAVr0Qdll1p0ESwT6RyJPfKHXYQYB+1Um048TzDb9nHZxUj
hK6GRoYW30mLm3fOVER8+lPH+Ek8mFAq3H6j3Nn5vZH85nIKLQ4sivUSk1oXJgGGlY1mmoThO3om
1ap0yhNdg9CnVk0NATaO376c6YA+nWx6cReYrIryRdQGs1JXv8Qvtx+RneNZ4Pow/2J40OfyZZ0a
QHnUmDlrqhD4PtKh0QLBxFTXNtxAbsvbf5UOHf6eFoEUn5ntaakJxOwfPQKRk1luPx37vwMvaIPD
kuIcaXvY9yCJkLkjcIFJ6py/u0YPCqF8PFNdAjSFwXyTkkyGYnphWLtDUZj5FEsvUcu4qctx6VBV
SLF55C4mg+xnkMSbAiQyxihksdJ8NgNP2+tCgiyXSRQM/XmQ1ZJR4OCVorNE6eIgWZwliO5hhyee
fBJ+peWlO+FVsLTqlumq4uBugjHTcLuD9S0nQuLq36q0YbHQUGF+Z8nLulIwuuX5DYKB5T8NBvOi
/xOjHxMb42BHvWkN6BMUYT9ezi//XGdVEsFrAxp9pqUflCngZ9Q7nK2HcV9+xsnL4jDYv61tx0rY
fUlM8MB7BdBeJmr0iHqs9Cf7yqiUCsUbNW8F4Ry7qrhHCA0jbGmT/jwVCdRIc0877qn3QLY370bs
LwTB/Q4ztpt344+gf3/BLI7CJKD9GzxtgHT6VydEY9pYqskArSGDu8eS/u1eruANpAa5EHdcrUoM
hD6U39l6jWn/GM1lMXIxTdmObxRQhMshb01F1cieWCvI6yXHjz25HkdveCo2F6ZEsMxYOpZyeyA0
fEG4yG3ohgDYuFfJRz6NACQn59yfrI49GObmhT/SGu4RwD0NRB7gNnVIfr6oxOIdWi2Cmb3cT9na
onI1YhunefSkQOV2K6f+Pq9yncgVEwlUL89dKM/IJMT8Puxe9j1elZJp/jy5TG86zUFLNaE2UDK8
E+VNrigSTFlyvaK+VBraBz7aiT3ELesMMYvj93XjgIzHjF18KA/fqTiYr6805yaL2wFDacSEX1IE
MSWXvpfGhQNXRJC1IQn6QTrftZYoUTpEXu0VBEyilejcjenM4dndMHJ1E7OP21sNgVFLbwtRgI4t
Plt7NB3DpZNq+U5tX3aNu/LgNaPpwlj9nkDlkQD9JaPxPXWCDCOIodWUacVol33cO5jUzSWM/U9A
hx9JpZXa1RsPeScmjcSL7BHDsgMOsBac0bo0X1CEOhwPDEkveud3Hx6B6NT8v6uBnTvrbXfk/lVO
i9ss/DPYL+3ne/dLkosNugVzXX83QuiLCNrGFcw/3DERZ+1HCI3H0rH0wOe+PPZMRdCwDGzGK/hb
66qk4cMfFFQpTQnq54hPJy1Wyrtjr4PsFcNRLshQ/Lse5soziHY6mCw4lsyHrtAH8mxDq8qTwV6A
8fUNh8Uv4iP72pR+0NYHmn8XoZFw2OUKuNvYG1jczQ6QSw5ObmE0rcppK52YPqzqFb1K/mrwdGWn
N/+hIed5GK0utUbjScfGQOZZwxhiqFhcTOcGjPoOE3IC0Mvdj50fPYzPrZEe6nyzn5xwCkFq5rcE
uEenORafnRm8Piznc2tYXoNSl0VVicgm5u9v0ha+ugmUm08iV3VyDDTKRE63URkPFxkctYe8Bs50
XkNq5pRIx5sFZFdD9fdoGb1LbFKkYwoAiIf6yNrXHf6QSgmzS5EBvjxoJzCu2ih7RFjiqGUcVbLb
iSzu2hbsSve+KRyKcfPEoBkyOYUDy0aIyKW2kJMgpUsqypAvThvVRfLlmfJpDRaQ+ZN8brqNMPDk
wmT9GJmAeVBIR+XM3YfRrJEY68OyD3ReSaXbcMiVmFKrEM0MyPbO1am8oUclL7+NPd4W76mMKoBf
X5gpuWWcu2wTouRTMQXYXsv94aqbh5mrmPsbUnSsgUp0twjBHx9r6BOMdxy9y54l5dppUCulk3KH
yf3GDOiLY6C4Ta9QjVcxpTs0I7gqm0bjeqznXp8l8zzZefMfIgClW4TCCZdPrxtpuh9+ojLiSsrC
MmBjYQMumyN0ucd+qmLvLUJ8Qo1Pnp/IxlQe0y2xX5SrF33HKyYc/ON2F2Yh+hg3VIJsqK2lRO0E
z5RnSkCkmhL+WKIe3yt77MRDZYoazNpQcOTLo6LXBqenNDbWG0sxpvzCHX/olzPWwXGB9ifoSkYk
ygqyvlcnx/Rh65rLlWJuHt/yKXuK1gQ3Kl//3T7fvCgvKwpc/EyKe5ZFegiC7YYGeUTofB4qBxIr
0IG4LKn9E6p3nIxB+zpydeubLgwI7IP3pHLyhg1ylblOfQNgzdEkzu1qFC4VLBGcnmA5MHs6FEEN
RF1zhFaGjwnA5Q94krDGFCV2idJLjtZvLMt4JzIwricqfC/E1Rwiqm878Azi+0CzneOadKjf4bHr
brHwy+pKNJn4BIG0KRJCGBapyMedd+rg1jINjYXAriAuFhvcMlxu18z8m8aKKFWiYziDAa3gUhgs
tA8ZUwDq2D8HRdKx0Prp9vNf0UOOj+M+qBdipPVE/bDrxoO2os6qUuPEgzyiLdSCQXBSzEllpR84
tXI8qAuqGHd8nlZql6o2wNobFDk2vK4KNDdRkjjc/E1aNZvqbRIsKnYjYoAe3Y+IkaIPDWyNbI71
HTwlFhfmA6AVoH4ZwO0f2LfHoZttlosqYAjtjsbSs65P2N7cKhZ9XKhoq4Lw+P1xMwnstPYORBSo
jDQtmcs7Ten+L7HUusuM/zmREgPP203oCYBmw2lzAQYULKvr03ibOiCa87yb8HSIT+GFoxHR4+ZJ
CXk9tSNmUeRkseQf/0wBJaNxlSW8GJM8wd8Ij8ns5KzIrmpg2afris7qJPCSUiDea8SUaFx4RscG
zeDus8UFHAqQHbds2KZbpgu1Atg94iHMKUAppQ8l7glqteebvNHRa/O5wjxuw+33g2TNtzJEwvSH
qgqKcooAHDZGi1YZwpGiuvjBRoW/Nyn137wpmowrptm8xZlY4PC/HLDhSgIWU/tWL0nWGoggXB62
JmD+Yp4tVtWkbekOQ64BOvEy4lNNBD7XIvYQ+YhrAti/7sk8pWOwuqle2ksOfXdnhzp3IVr+7rix
HSfJpEuQzGlg1G8MQ0VSR3U/ZPqilZTkQqLpYqieJsZ3RtN8m9e5f0S1dRF9eSCoGQCmj2IVtnT+
RIEXdFg4COe4EqVt4TqjVTzM1fklnKtYrDQfLzBWfvx5Gf3A3A/akUWCSUq8n2BxMO+a3EAowcuR
Xgf4Y29u+y/yi5Np7MzBn3gl9rtYYSyujDgvVeG1NUnbvxpTNR4TBViqgoy9ZUqHJTUlfzRwprcV
1VTYY4k4CxPURZQ/n44lNET9CwXjYsv84HT5pYMTibP08EN0tNl47sezXvmc7TApBI7NVwGX8qKL
CaZ4pJXGHikzP7Ba0+DVkH5E8omTCW7bHgTFdgo1UhujsSmCGjg1sd39IKpq6Q7Wc5uFdeJzyVtw
YjBojbJ5Ee3iWst4EH3k6gpPD/vhwsmYdBFuJCpLNCWv1s4HhheMTLXasQe4lH/1iCPaR3uimfrk
MBW8T21wK7Wk8MZzb3OSBbvyJOgxHbbRgvuP3IWWpqTbY42pauadkSpMgSsn5/DZNpPRgh3ec+LI
SVm14dFz3wqmKWIPb8VdhPHdzEVcW7by40uThggpCVe2Ki75gty6OyQ0s5yMMcGHDSZ7BdKi7+U0
u9xkIOpdI1/yNvcpS8wUAJpZkguQWbkvqFgUPmXZkj8d2UQjGUOTcpW7O8jDBZu/Q1pdQdjFyXDs
YbP73YlBrZWLVk6J92wR/6lfJ1ZXXlr3d9MztA071H+EoMOW7gJa/xreHv2JtC9a2GDc8COK3S6I
mDc1XriUC5RygOBQhGtNVe11bCar7LwIJcYYXgILc8/jljfNQ84hr4DEGNscTWlC9aZShmh4zmkf
WD2a3s3uizPQTTNVYUdS4wVg96aBkts3RvUbcvh2WsQZNpzvCi5I+ktaN53HKc9OdBSdcbGK/m+N
vJvh7Kqd7QLCOo8TFrJkhv9x3TZhBZ2s6wsSk2K7rFNWtf62IcVccjcx9+lvhfyygv/szzjIuxvd
zBsL8sA2B3WvKoVJr8mCVmtViEQwDPIrC9QxcIHx6HxK0IMZK5HnDOGxr7Z4BYQiGmqJDa34tExx
ewhfNvGqR4yqNsFTvGmVsWyjhI9Rs8NgVhJjlYusFvSTBHHXPcQ8JWr8YdSirsFgcXvh2K4vyIbT
ydeq0QUo6O3R9rWW/WFJJp7fKiUnGaMBG3sg4deQx2PYT+1juz92hvuTxTzU14t8BZ52OMLgDaLl
MUsZlHeVXWPzIoLnWPd54D8/SrEKFwKeNQS3wT5/G5BKHRZh+JYLXj00y8VlQIpl7MFY6tSBJ3HZ
B4/oSjc6kMRiYKTP3Ak4R9Xu2Tq9SHHs6V5lDGelzZgWHOR3FxEV5apXeNXjR6rHpX+vtas1f+uS
vMlj2FsqSHUKJAHT4Z5t6ph4/i0LHjVb/daq8Cmy1YQbimeuh0lZtClt48bnftlhvJ8oFlSeu78u
zsjtqe1Jpo1+y9lgrPTJ0tGxzSfOKePLe6c70OyRTCS9EW+a4c8kD/tUS9cwYyVVi5OCVeGv+uEe
EKf2907h3B1cq8xXnjlNKq6p6e39Hz5d4P/j/d/TWp/UFg8dzloXazQNoJu1w6iiOIkitOmXLOx3
Ota3yb+EaKIoi2Ys7b1o3K34YbpyM2KLM2MI0rFQkgh4EExfCOt1MsDYQC2uvIMmqyY3ZNtrgUiQ
RV9mhq5HwMjuPdp+gMPABl5XeHTS0n9qfe/45cIkOVhCClao/ZQskpV7HXQvST4LmvQ5xTbZtzSa
Ereq92RddA09gFJuN1TEqU0of6mS2GkKLjCwdGUT5m6dcfWrgvbImVaPHrgfho75Lk+pF6Jl1qPk
99jnGGY8hNvoazTwPjIU6Qy3odiPlg/0g06gPsz9rTgtWf3TSA+rx/fwEnpOg32ahpc1fImtcaK/
vBO1+GzR5k4R6dPJGeg1/KxALXUl2yXDZl7KdUlDn/faczas45ms5ZA79zz4YziTqXA4mT2wkePV
glbH0DlpzXznrpXk5i7wG3eqkuN9kljUUOOM7e/vZ26N7ucxueP/fQ0vuHN6IDhEzUgzEM+Q7n2W
1HQawkmddpmlwILTbDHHqYWLAOMqbV3u4Tp94ZAguVsODVOBC8gwUGkJW27rAcs1iH75yfcVt4ih
vlfvcWwNpCMPp0mglRYSiBzfee/f7VmQcqilY5Mcanf8gV4R6jcZQmN49Aj7Izfa7PcKDfjf7yik
mCWc/ninplbaxRw3cRF64yPBU2MN1FljEHaF/qsQUH96LboOEsI5jv2vNn8Koic2lTHmFAqtkjsW
JISTmnWC/bn/5CcazqFL92sNZ+M+FX42+abUH9/C0BJhosTOan+LsS1ZmRGQjZNZwRz0WhwmNaFH
RRM6Qa0aW5kUpcsjZxd5GNzTsYkrHzkMogDOIP2MOD+wplcd0NddJCcysm8Kn35lWAlE2wMzGTyT
r4ZBOfgC3zHJXjf0ftqbO2HcE3AVX9GSZoPIi4DqOKXCLDTQedoXVnmKBqh3dpnGblKAxEqKaCuW
3uv5mGysmkjfcSxrA2QPPqhWhsZeW8OS5rBGxmqTm9VfP1nVouK2LuhJGkhVLXx2MK+JleMmabnG
aiEK3Q5lR8lsL3j4fSOsN1DLzU6rHpa4XWinIr+koxJVjQhnuJBsq4birhoPP7pAPyJIsdDlvoZy
uWRKBlivlaFMbh4JYnrmux/tq1YHMLsTOGQ2Ofm+rfaCqv2SQkb5q8+Zk71z1l1KwH1dujg0Jzy3
2D7lkF5uLopR6rYb8p7gmlWqJ8zWEOKCv9ZV/wiEWRb6USeWYwZIVrQKBX/tm4llmXE5YcsQMsxV
ChPyXPV8C60YTjtPXCrG+tLI7AZNT1Bdu3u9EkN4Aj/Lc2qwLmKGI9+1yKGdL6yRb7us1L+0fCX+
J81mkU+qBmmFmKQn8ALkjoxNwu+Na3hYHPEPuwJrHLXeHeBGsK/OXwIDUKWJCNcqAezuflTJ60Jx
Kb2pC4F8yAqEzOKZXOwe3HpAkKybC95VyHoV9txkpkdovKGulrQra8kO0HejwjyrBxXgLNvEMlIW
9KijRZP3k5FLuFtoWUj2zNtPZqZEvOWjKrsD3/B/7w6bMBMhptLCMyIU/S5gpBVlK08woL6stEjd
n855XC5gx2zUAG3GPghPkTOz0mMjCt9psPH7S9FENnT/oxoiOU6HnvQL7BRwoA+QTOyn91oPdRyI
+Px7IHvONajl8Jb6m0iiPOxhbz72FYaezm3myW0Yd/VJDcoFWPdoiJVDEjs8gLkVpzSS3qmEz8N8
zaIosfoMtTD5zg9/CMRySEz9svxf8KdiyYdVLoNI08nb0BaHXdnFetr0Vjnscu7N8towA4avCQs2
XRoC9HYADn0jYQEkHP6WGWqagWd+BQt2Sf4l3ZxzUV2wTdrjmdq2O/jIieL5IrOjTa7bA3GZ+zd0
62wQwMfr9AbqYzGikvSCOLRhINEo1J9O2O/eOfeU2fZv6l4nCEYCSMSb7kuEi7pVH47pnAQ3wvWu
aylqc/c304MXSZYb0IM5gXjZQC/4AzTlmthNnNVJLQj/BUpkX5ys7Dm9ARmBGeBsXgew5xBJSK/k
EyMuPyGNl58jkNH5zwdlbkjH0dpMyuHwJaNpEsDu3aZ5McDIYwscwDOBSqo2enHaO2lsdywNy1m7
vvY3DlQ354bfmUdAm4Lw8lECDxFldwyF4CA1Iafaip2oJjNfXJRv8R6WC5LMKATSe3BGWP1OjgkU
lzD9MC0H1v7ZHkW5v9xkloj6XGzAxAPNTsR3/4l9qdKXnMs1AQc3zCRZcurLE2SPxkP9Y0HY941s
IQbPasKnejHTjjzcCqqws3m5cOHbGtWxSoETUTZ6qizADFO05M90iZAMKhrYl5221RmvHC7RarBN
ljTnvMkij5JrW+2O8HmjDAP4wEsy/VdA0DiqL7nGkMrOpaT70exCCisH/Ma4r5rDkWUP3SNQp91A
d7YVTp8G44FIkXNswqcC4TiwQUVta7ABekJg4y/b6oBg2gTt2gPbNo6/UIU8Izypdt9zSKRU2QAq
nsuwLS0yEysm2x1v34/8PSCcz6Oy7/9jZ6p8UuRfpQhoRktkBvfGQLlKzVCVwPfQ982bM7TMsJhP
bpAtwYgUkJRCRqXhPbecF7a3q40r8sFgTOb0QqXijVnVOY9Qmp00UIBNr7SGnQkMsds+nUBD6CQ9
CVWsJLqCfSLtSGFF6QNm+g6jVptgbpRb/NlrgccApUBZuC63n0vxu2zk+Jk/wkHusBWBewtX0NOb
7LnOPUaTLK5DslmhNY90Ku81NiPuWES1zvCIFwM6C/tcx99pJFixZiBSx58uvnOmrxfkNZHZMwta
W5bjYvtw2rbnvmsO5A+bYqsU2PzhpxwZRWLHljvYojhXJsLM2wX5JsjdJyeioDOWy6QfihtEfHxp
7TWxIZSBa+GwZO4vYW4+8rqNAyENI/Nka4Jw3w8vUoknHPXqgaMZK+ZHQd4zDQHFZ57eNpqR+ILA
2kNA8+hpfQwXhBTymWuc8s9P2aP7jNZhHdGKj3gnDOpUB0iZkHQcCwGQuUA5IPk3wkb3Yv1Xcv7U
qWzbMWYKIkmfcCYB1gVzWQ0jsICSWK+dlZeByXCjvJPITj1xFGMArXmrhcimvmBQOD+fpACZ90Wj
sAtwekbs6IGB5LtoYdc06M26AU4ZDgjGEaC6HW60ISKwgAYCmJQydWmh0dOFCOxJ3Wmmgm40gAn7
l47KDbPIzC8OnRqFLbecaHu0uaS6GmdxrT+YDGcxm17r/LtGtZqskiF0LKsYjSk57GFb3RpxspdV
87PCZ1lKDP/Kc04ahD1IZdJfyyWc0MVlBAwn/zM9E0fBfb79AGoHJTE5Zq/STOgDgISnMYLM+n5Z
Ool7OPaS8A0J4WUutGKiPT4xC1azPsYXqCS7EFBxS4cNV8Z8F937+JtpYLs9C9eB401S2gEqnKZM
yMJP2Dltqrcw10ICuy0Ba8PD9n66iRc3rn3WYaky4kvjhbjYy9PM//N2x4pDn2e0JwG1BgWIErmc
RiQOW2uskBNEsY7S/qC58vUof69BA0jSgZWSrobyU+ajFntzYPjY3+KwAeo6m4ok8SWJYR4rPZgk
K4qz7bsn5ttCPj41zNX/e+92Kjf6tpFi5GoGRucmEnLalvOB1lnYTYjEC3R517Ql9zZ+tcR1W/U1
ChDygBI2llR8H3ohH0E3SQcUgJVBNGcp+y/jwuDpxePP5R5ttae7kV/renGhnZOLPjhiYLkZPErJ
l+cmv1d6Fm6pccH/LWNPceG/eqqe1aZZAEBRJcxVXUbPUQ6p8O73d9TcvY8nwn9J91DAdBvYDnaO
ndRV7T97z/WuGEn0pI8ZjaTdUP295Oi2kwqWt4dp5X6Bqms80xMGRhsiRHEA/FF0fYPibuvAT79u
gwIOfHBTRwaAF9nyiRUyAN8dquvUXd9N65OsIhQlQreRTpdVFRWXNBjoTMPNJV6Mdb4MPSxvgdkd
4uTheJO9pi+1Jq2QJ7n5FvmSqOMJl7S+Rb0RdR5NZqFNg/wF7eHJhDOIDIyq6nHnZiR325D9KQZ+
QAUyU9ZnAwVl2kFc8TqHQwMxcX9cgMOlnBRycfIA5inl2warGdZ/HI7cH1Xlajxu8+rw3k2C+WU5
ACSMIckytLItfX5UsBdlxdmCv8Umhhc9KBqmlXKBqlNbnOla5QkyvVLEjKvB3ES6dZALYo7wOkHW
+oA22veIONBW5oHNURyyAq0mgs7IbisF9+uY1Ddy3wlypkQfosEK4mVfF9BfKPfIGDLjVC3vrk4M
xqaYepPXNghVWDoxl73yaued631TrYesUpMkJRXXaXBzcBGI3jRWuRy+Sek00Eywph3HxDzS0+os
KcaFyIXMsnfwPXFHFC6oBSSlS83McLyBo9WUhUVTYCYt1Muj24Yv35yIL4lB7F/a61I4E79Ktjsd
AFryXtW9FjmhbUbH5AXx98mCSUd16ZgF3UPg9n52t3RRh2eDENUW38F6DkFHSi4DKO2lZa52W9z3
g2oA7286T0Ftbs6I2EKeLXhCu5WOdJZMyV8lCa+5HngftezYTP43sx6x9XBih4XCEE5lMiSt8EWT
2rz8O6mdAVXwNz0Du3P+6zbab1a3Mzo7pGlgLteabBTAXzv2YPO/+51Y9cCgNf7Ru5sz8EBSiUQO
irfOy4wce9ixy9VRb5pQP6xRuwq3saFdT1A4JJz2CiAhQj4evlEQdc4UZ3xmSqT2vXDfUbI6JoMB
/NVvNZA+VgJKs1/0n24kFI8xlWMLmBrFlssB7We0D97CRcKPLPyjeNQFZdaXXt9DsBjopqYK/MUz
hc36+AdKG5V4K/rMArboko2Hsy9R64Yc1H5D28J4Jnf7k2w4MsHWe51ccNOBf9hzgQfZ9bjAP6cs
kiHgxK4QylRvPsv+iUdDDtif+kIo4I1tuR0Q5lHxQwDGHRFw2ct7dA7gfaE/9DKvBSu0hibWBjCZ
8orcuWwCqb57D/mFgXa/jW9+fbI5D2olrbYNHrAh5XvV0pB4oEWcxAfkpQ/+pa5pDOJBy87s1T7D
IkH2STeVBDP2H8gMs3DFtRZViJzTTQ55nsEkl9xTbBt/yvbRkv4EbPB7ZdYBU9LkFQ21mMLGht2b
apq7Pr9L2wuHbmg/baL1f0BFaZHF2rz4TgB2CvySGXZeD+xKVf6B/ygYV9z6izkePIHqQxw9s4kc
tvVYgUBOKUJhYZOlrzqFBLKjuQXopgUV492bl/W0lKxibmLHCtFr5exPAqVaGhTtAn8guzSPzK8Z
tt1iDDrJGvzFKZUerIQnJiaE6BeQGfsgFD0LukmzpFu+jU10jzOIqkSajCjWFDyDTQVUJY+Kivei
hIIQ5T/Q/6SUQ1DojfC/bhQKx0hSr/f3rzKcS8OPnbnkwV1y7pBXkMufNrD1TzDZZaZKz7V+QWNK
+B3UUOTBdLhhCFVLzGZEkbn1FMQMsVJB2NbtVDKe6UqlJC8+GVTgnfYSLhZ4iIVGXKIjBL5FSBKK
exV+IUkno0j5+Mq2yR9ivqrIRqNdh+cRdVETWS2CEfMg2/HowfJcpUBbIZzGaMc3sKK21B7h6g4M
RlsKnXl/uFskwua7iWQ0JJVCyfkitt47eDjyOG7dinTEL4zWDq4H9FNHFX/RIimxMr9B4EBhrb61
Ye/vT4HFy+/QETEt5EsumzKKjFhAYGNd+xg55mpnbudNU8b5odbFLvjVo0wjxtMoJZLxE8HtcmYI
P5bfTJbhSJomRIZ/fHWpA7LpmplR4WgUBdf8rr9T63eJvIsO/GKpBTt8qmhKhXA4Ec1CHKPtg8Cp
1mN5XZnBYx9in8PCea1Zx3bnpDyo+9spxX5/jV2AcUiE3obLnpRCXGRTE+eghdzvTohkjkq55F7K
g0yDXmzk9hxPNz91SUrxe2UnvU+mlm1KXQakvryVjD8elriF2RbxoIf338j2j8DWhsQ1f/SRUsv4
XVkBopy9bgLDtq8/7sWoGQ0RjGP5sR6ekA88a6G8AUJv186odonJMFIZD/2V4gk48xzuvcasH+xY
ohCCeSDlC3NxHOh3Cdy/4Nq/Og0F7nJ5K3oYC1UONiIE1v+CBOxLTL7ogkrjbYgjwbofIynXUa95
//RUmuMMKI7kxuhI9Kh/zGobkEckihRgN/+iDeewSyVDbiyiHkx+MJx96HHcERx4UUX/DPaN0ZOH
2KKz7FkSw29XgVzmBhTeGveX3ZqLLOSacs4IxGV+BD/T6+GijqVPNkez5pTeA5ZpIrmABWuqSPaH
lqnsbY7NWkDxHJ884CZSMh6QU89496TA/6wxj70LnohjtMhcbemljCfCuKz3m7eSDrrrIZNNdiZp
MYZrLQNOI7l88O2VbpgZLRbKn94ZWap1FaAQwgmt8qHafWwxdA52JpiBf+R5o5cvqqX31fg+putv
P5VStxiAa+NwvnXCe13EvPnyx68rSiGmy6iCJlTtpKknrjGWAkEe7nDNt9RKXqnUA8Lws3Cq+eO/
mLEtxBhrjVWX57gz1VpbVVI6qR7Jea6g5q8fSr/dbl2htqZd3YWFhgQ8KucTUk0bY9K+s4+lJ2yg
UYVdcMf8DcZrzXgaraCOE+vOI5rd8UqHo7Ua3EwYIIT9YhLguUN2KW5nf/jHcXVT9DmqSdQeS0ZT
N7w425XT8eVJEwJTEEaOVB+thvxQqykfyuYx9wBSkHGH7mEbjABWYs+m5c9O7qBv0O4AOc1WtdvU
VSk8Z4D7FC+g6xHjEisGWvZtZJHyeguaFVsf96cPgvP2Z4gM+HPXOrAwRz3I96by/+QVTMhUA2Zt
4FdeP5rTXFqD3jgZHbmYXORrioDFq5aJoNjj4DK8mfLfvMAAtZB2Cn1nayvwy0HlcbYEkkh6V76y
1KHQayPhrQpJ7VqJKRc4A6GCdwEQhMYSYK5ctQ7+i8cYydsV67robLVt+W7mVqciHroz5podDpdc
e0F0O+06ZqW492sCZJnmivgQ4b9kl9NjcRmpv0MGnGQRRmnASPmZ3+fBEIiq5aX6k/hr8EOIzlQ+
XZeD/Las4BWuXQbO6LxosAR65qLjb12FumTtiHpnOLfX0WaZVin7b4EjAAZlKseOixDFbZSK1Bim
6eiS5aErsVqoXd5TqOlRSokgiJMWD2xWkTgLZJcKtfACKbJ8gxxNSRHKKErjMDQ9yj7dybYZPbWV
2tRmoVLnFHEsQe2D/f1NmElhjquRzhVR9JtwCX208RDica5hzs4Pw5z7cGPSdyw5BH84bFbGimrB
F29oXVGYP6Kp5LwXGOgNEZysP1chqKhVl4YaklSjl36IcWHPuqYBU++ZR4VvniFAvGHLsRkN2XY2
ofHk21qB3D1qUixdriSi1Jgsvtycg/dI6cmb2knkoUzp7c0d3cpckfMPIk2fwz8CWvQrY9RL3cat
3M92Me5edo5YJeOHGvyFTsTRzNt+FKX0i/+66qhkdALumMcp+km0CZp6eeIlFZxFkpHb3VSlgYQZ
e7BelOhDMfs5JIUFshG4CXOeBfZXJfLh2ScG5yHyMJ6Cq+SwdoVtJLuwwJsllyoZQI+LZ9sIu/Km
LbHOSLG0AzhuGFITOJgEaxe4728q3m0u7HGINpiAFK4Cp5lJ0t/sR3EEOs0JbsdgGgetBm+8K7ra
R8KtUATWZy/sHG5hIOZgo7AUP+gaI7mNevnqp1Us7fUR/0uT3gSNYhL5z9s93ROwX+YVJ9d/xNqm
XsC9l+kbvGW5RqxNgKq8MAiIt6Pl+rvLBENVnwn8WAijSwLu/ntYIHeW3xjOh6kNdpVctbet5UoQ
jorSdto1SDjtJZSLGH8SIqvWhdq5j5f0AI3zvz0s4jwKaNl+Yze6ewhC56RqtZvlqXq72DK4J5eP
l3oo4CGxvCmBrNC2d39m9sR7nHBHctF5K2YZ2OJQuiQwLdBbdlOU7N4zPLLYcBxC38b2uDvAxZyt
61Z2IRMJUuV+9i1BZLcd68VE/5N356i/rfAE24hQPQl11NOWKKjEv0DRf9Ojyt87Htu8t/0QAQHW
FUk9s/EHVsFAWHIGoPviD3cTx0CJQtuGMG/E9VAGbvOvkt2ifQ/lj7m2+5BTvakGm22OEefcOtZ5
bBZ1qjBF8KYpfC/65LzDvLQYMQSno1HUZhriykmSG/hu+M0nv3Lh78MeUyt06jHhe80yGx3MkGSu
/JGUfLS9V6bpgHuL1qASPvNCeRz4ym71BMYgBn/x+9Wom3cRfkAVEG42QiNyNWUPXcGBCE+/f4JP
f+I7Ni2dkcLqROGcStfo+jZt6dyvtLPZVKqi0ElbGKdWmy4S3679ILTWJE6NgDLBmfUUjoNABHCL
dJCF7oqMiDcAxERbNBfjiyc6A3loff/MT1Zqs3CuVMy42xO9z6k3As2031fewe9uuA9hUtZTjU4B
c+3iuiGhT5hn3b542GPP4zvoZffRGNvWVVOeA5aXsxtWSCJhk5r2/hsgBdqANVfg8NNiZw124Avm
4shGgr33UpSDIUJL5rysg2utMy+tDBjYxmNzgNrmHoXuCf46AqWdYd5UMTdpSBg0eftPpZEXM9E8
2kwA3StQD1n4ljO6SVMhZgQJUn5e6bkYA+B2rdBnubyjzFU7laPHGDInYkGTB40WJo8bKmsoqFzD
+aL/V4Bl4Oe8JJEWX5dMytemBzst5qcxBPCNWZvWrweQcRe0aEBCjOO1db47cUniJpmtR43PHN+l
V5OrGq3HSMg4uVi60hF0e9Kbo5cwO0/j+EZeNqnOI4hJRjOK18lvbXDceaFjhUYyI5Ab3TqKkGTk
fiBHAhlDT/6r6sEP87JQZVBo7kW1N5Iknrv79i6uLW7ZsQ9Ou5GbwPVuqGpF0nFDcUcS11dieFVm
kGW+SeaoCox07JNOwh1u/P3PInP7+mmdsllS+teDstn36eyixi0iu8D+nKCW0rPPX4IZIJGQOUik
Yketo+snlt2MuyUUDwnBj3SnkpC2df+BVJhc74rO1oV4y+lOpFAkfjNbgBaoNmLXdirnZ59YB5Z5
F27Bkg3M3ijiYzQJcwn2KyI7Z7+BGXdobItgLIPkfHFAvcxXc8Jpp6eAnQ7HIz9jLHeyrkZmVwH8
zKYmK/ZXBVoAXHQX0NGLiQuK6uDcIW3PmZFz5OKZcLsHWaoIs9A16wxHYAyiraqPfIfqj/bUCIOE
+jvCyy/f0OXU/DMesg8gM7O4yCjPp2h/fC1dP06DCv6sklWDPm2zfkHVLZv0UQ3fAerzQgFpkmQ6
OtilMugk6F1vYvJzEs8x+hif/Dpd8/m4lF9yD3kpRw7p3Xid5iGEizgTXeEUCs9XdPdY1LgZcfY/
YeyukhKirQzghnmm522TuBzwQ4qt3cRR8HcrORv8jJ1PknzZfp2luqfTY67fb6flSod8IFM1rMnT
YpZp00v0tgaTiIia6SUXgGFen4mc3LCPbFjxwOM/PDHzci01YrHDNw/Afoq2QKj0K90nNSwEVSWJ
di/mF/zX4BqafvlYMbIll12n9ILNYebA2yvVON8ynvDZmvVuf2TEYOnmocKLLxeZQpnkgxOTZirj
KZXnUDe2bTL09QUclmnLI9uTx9Lm103Y/E68SDlMJRS6sSbr4eNhhZlYG+fWdgjEjWt+P0y6FUVh
/+P0HEZcPqyT6sw1oQkDVQKNBFFkbwAZeYJM/uamHYwhJOHY15qxtx1F1R7smBScGYUGl2SBXqOT
5QEPVuL8A9pifI8CZGeBBxFTtXukLtuq0vufEQmtvYJe/S0LnM/xSE2fZhlWMm/jI4mAviDZepNR
Id9g5lbHXmEv3z3Fy6VTGTnhy4zfbr5ylrcaWTR8le9N22urvVRJV0b0kg6bOfm0me7ht8M6LQ40
oCdTZYY1kpKpoCscWE2hM+BqJ36w6Hiw7gwXnrDZGkhyalSWyMk/9yNRI/ewXXdVLkMTyCkfxMnh
Sr8xS3Br5K5EYDCkV8nRjkAM9DZ05FcdJK5mZ4w6zUjqpduQrefaxXvZ4me+gkoFTTRLv6q8JG5B
EeaHrc/VPY0t8ZuAF1F6hrS3K9ShEOUNuRN/4RRc1EVtb8d6haBLbydziEO5kB0nppf6D95ZBnTV
W3wr1wAnbjunMefhAdI5nu7+SUSVX6SjsG27LIYn4rZJFuwCLy/Q/jHpljWv7BxgDSFJDXpHNn3Y
/OT4fcviPkXvQQXzrcs/SS0Bie57bXiEpeCGnoUOlzgPu4It/qrR6Mf81nBgTS1EDGBuKeQg0PAF
qSBKTPkHBA7QRw5rJYljTFrk3T15oxTeOg2eYwfJqXsvNHdEp8LiB0v2mssM1h49TsWmlivVV32m
/cJ1x8ZupZeXJA8Ex9NCkOI1W7l6TntfEBACIF/iHVloIXoPN0GkhaStm4JwXiNTYXfajjyU95Lx
qZfDeXzCj5rKoK6SzcWKe3RU0LezOO2r+muEuY9mUroHIFQrnID+gvQhpwerA9F6Jo/aj6RI9I29
UuJpsMO5m2OhD/qUKyAsWZ4CatacCgN/XO4idE1YnBZ4VmykIZ1650TBS8UQLB5rpLSDVdUCtAwv
s8kYWwdYPaqU6GHzj8nonBH+7KF0qMI9HsgwaOc7RQ/0Z2MG94dSqqiP6BE+rGYXK4CNyJneMyfv
YFa5ZovVY5iCjLWFiVSymhRZJ9LlIMSUUMegclnNppiYnWy8KN265J3sWPKliUw3Q6zYohKyfMAa
qq0AmxxA8gOJzdM4V012vo9MFDxyGIx1iZeH2LiDxn2/wcgjZp6NKSblm2tcG86pxz/yEm49gdMo
CiUOq0RadZceSYtmBLpbrOZU6UJfjrS8bSQT0rws4YK121TevQqbN2JqDGTyvKcKHbsj3EmBwnZs
ve3ERipYt3ZcYMcBMIwXRVLKgBWo+V6CFwJXLWUyBaRDsJw01CEd5+EQwkbc6LJwtyH4qD7KC47r
SJjPbpOS0Yk8V2wICYy5IE+zlHz6YVA+4c5kP68F+7dquS1C1K56v+N2KPgEmyaiA9Gaf2fa6jz3
UywBffbiBT+ZTxuMZgBSQvNUIXayMnOdpkkSj0tP5iw/bXTyG+rh/EaNo+PNE/kvcFcdvPZkcx6V
oWoUtIODr+5TWDJyarfLNM1vJbzHo5dBj2vVtMGwrNBRGOL2FpeF6XaIU9qDDxJpouls9fUOJrZB
+tbdHkDP2dTcOzYL4sEz5PY3vDQuXOkHmoM0YazLKF0FAViBsEpFSoqrGCgswXJqw54m9EX/acom
oCCjYs6KWBPQHcSVvtDmgramgwnfSb8uvqNhHfZfYcGQrhHQ2lBBfKcnrDW26fHMyjReke9tGCE3
9VbgCvVDia+bVNnQuXOietYIBLk44U7VJwr4NnjM8d+97+KHHeDCIFUDFyu+ZNd97OF4jED05fwX
yEwyRpeJY+ViOj0sHSDbQQLQWe3hWauZsyQRYVGqsBTP6XuNlvJ5aiMvaYLd27Utfp+W1LzLxFKc
elWteGIm4SnoeiN+C6fLGlO3K9RW29hFpBep8/5gpu6hjaMrLYWRxTWpP52oQioJV//YN39U5XJ2
wK78uwFCHg9YJjjR66fXqlNtPSerDETmEvvmMHZ89k7CNxd/ISxmS7vmMUjUlPHIIw1Zvcd+cuxV
tCJVuZorQDE7LaqaX38nvOz+6l0cO7s0cjrjkT2hllJ02Qo1ut2BtribFCEIJoo2vfOQPWQv2gwX
XKM9CKEy0ehNdm6cFwkmOqn+eCQM09cq+m8bm8++VZESkAvyG3fVqt5StlLHAbi0l97Ko2LUWQwT
o9LoCV1g0MrRswiUl4oQ/qpA5mOAnZwTa9UHrj8Aw9gr2VA9ORFPVkPniBHP7E4yevnMB5ZDFCHu
egHlRRYb42w/4xqJh4/EFcrtatvzcujQO9fbRoMIVE6pFIM7OGkOx3ZACDLcbjyR044GRrpIybHK
/SGf9zn23jQ6HoVRmEqT7lUAX1K7194zvgOqgehoPpr6Pw479PoTT1MDlqNFTARY5+rK2Oib5bDj
98iRgePZ4TMOPLMdDV+CJFUKWGDhpk6VjxaehfgwllC0Hx0Wi9k3bpiV3pxLguOHIFBFRDAolWZy
kPXIkMu7rM5ByWXsRItJ1EPGSPcK7MDhZQL0LhuOLr/Awa/QMp1YUbuasUIzCmNBWfCLAV6kUIaG
VtzOjHpOc8KuFy2ir9vYuQcqlY+d0lWJAIdJ+2UA2j1xxDw1suTU7oFixwB2LdtKZ8BnldCTTJTF
QApoOeWaS40iMoV+sS0ARIfenN+FcbsPfd7dQNId5UFwnFbGd/2oJSGyHycTd63tK7aY5OPG7tw0
o3kEWgTcSfTa5qY8jqZ96Fpf1sCKWWecj+sndrrEQ3bzTpXX3eT8Apegm53CjngzlOE6suDWb9Os
nTWWeIQykiTXcWWdIvzuM01eXr+HyWfX+qbBqYRAtGi4xdsjggKu6NI7gCcseEa/wRa77SYI97Pw
XL/VRghpqmzwRp5X91QzrPEwgcMQFJTHvvTW3izpFJdQrxjB4PseA/hU3b0sNg2NLJoUynftFXZI
Ef5s+xsbinb1hhiCxFd61vhq29BFEyqheE0/KF09nnXSa3u5cFJ4a4n7g97aXWhObUnzBqlVy/eW
HwrDwkA8CCZIXgON3nftCCZGyKdZB7ap7d7FprQAfqepuRrIArZ1vGPsdgOg1EZYNq9A2/+hGTYP
0AWYO99aYbbjYbtr3z6o9MNHEkLCHPZxenYMxhhOZymm+/16xJGlt0edf376MsNTy+CHi4uK+BOf
+neQXsZ0T9gQJ+VVfkmNTnGn1UzYY2GNtP9EGnjoNN58YH8jB+AqcMj/RCdeVKTeH1V8pvRotptY
SKIOt2JOeq78s4YK7y8Lc3b+zN62+0HK4s0RW9x7lTb7pwQhiuy8IDE7aZ7elVP3Z5oIASi95Lzn
UFW8aUSqN/tZYicn/HITX3h0CzszYUNnrQCGWMlMtnT4mmwZ0OwnFzEAMhFc0cVASipAXoXzR6C2
LtT+COlSskX9KRsh/s9o+m3z6gkhEJHC+ubLSD3IyvW6l+pWaM5BibHPOGnhsgp/hPUar77VWTHr
nearzYRo5LGTZpUPxJgNBgpeiOb23+KXs9b3Pq5H/Dh8r5Mk0cBe3NQFLE3flNrlhPytFP1ZPSdQ
LSgSOGSUJoULf8XUmBQC2uE0DqcbRKc5eVAMD5fwpV3th0ZZSPebUNa4jHPpTdMKlCBnbI/+Kwz5
A+JIifVxfwH8bMuf9uMrNuKiX4BQS+1C7UNCdIL3JXE1UOfbymrq5+8rGLhq2I0mJLeJiRNLk/Cq
EdzmeccfDKpB4qTPptxfrV3iabFp5tZ6+gC3326PoWh/LwIUwvtqmdy2wYUVfeD8FDQT5sycPSv8
DsSguh6AlYcE6NLQnR2au1MrScAUEl+8b5yMmxDw1/0p6OGLDb3R1CBxXtG4pdAaEsjqUUYN23Cc
RIsi/W/0thqEfoyge7xl6NALkSPSbjFX91W+dhXNScnaXISyy07GS6ZG8flhFmJsCeHXTX/lUZWx
n+On5r/6Cx/yvIZTSXPe6tKGAjAIkAQUdExBJ55xWO1qHiCTVWRcKl2nVQicPhh7Iyx3Id183sHp
aFf5/0C/y+osPGhvv0OX1r+Mbl27UXOIhlxla+BmQocnXDyvpxbvdIFCUYBVDQTwaIQ0xJkIi49L
4RAm8qHkBqWx5qovBF1jYaVHYA/+sjHiD2n9i96SO2AU2EQ+hZi8Y7kwDANQwS1PFPDe0Ow9pWnU
N4XgiOKsD/Cl/PIBX+Ngz4sRIA3OEeQVeuIqGubzyy8zR7+z66TmRm/YHv0aBBAcwGpvpTGNOkxe
OCFwLgskim0aH+83Vi/iS97WlebtwtgYD9EfA54Sn2ZCWZlNKNKlkt74PxQbTt24cP0lq5QJax0E
O1bO0kgFf4WuP9R3RcdgZN6Wrq/dYI0ro4T9GD2PBsZmRdeGqOI0SZy3zSgH1CDIsFrLIlqvqtky
aF9pUoEOehEjb6H75pSXfAdffcig9pgeU0fSQ8U7QxCzI9mTeOX+Ci2dKj/WlyXrGFxygjx3G0IO
iemF+shgwgspi20D3YdJBBM4lgT7JwOP5jyElG/cgEO82kLWgdbzhH5fASjYCILf/IliOkGYjwTV
KC/MhB9eXkxeMgXYcw9NCitQXciIRFDLaLLMOMCkxlXVUu49y5SSqM92wIJ9haDwCKf49l1pcgvH
wld2GWN6fPbA7pogvHBL+Husnkb67ZKDOJHNyfavM1UN9dZMF5nhR/OCh975DeqwvMPRaM20Sw0F
TcPeq6Uwr4Wqd71IRekgcYSuJwLX8vGIsDhlED2dNmjOI02j5cpLcsNIpvJX1OQCV6uEJKhvoVQA
jDUN6r1CGYJrfDZNio6V8VBBvS3y/wjbdtqIMMoYvxcW6OuLlKAJwkhUtq4xKNgPDzJygLEHAAXW
B+lMo9JC1AhLHsKVQ5ATxLpzbUEYBK6nJT/PmAS1FH+WrsHmJJmqtFoY41xc7EtcmQHdbrDAw24o
lo0VfgQht2AtKdPmc2I5P7XVgfWhbD8oH8jumeeYeVAMF7a40zbzfwJA0tUa1wkeVzWRTvFN7wLq
dv7XZoLrDvDje9F7Px4p2irioxATJnuTYIx2YJVBE6OPYmgvKK6hLt3wjEWOlTfbovtnlYst2Vjy
GpMxDn6UvR/+ls8+bfKdwVv9Y47QoPcA12JJ8s4pcvxkoNeDAGe+KwBluw31G8Chmmu5IRwV0jYG
2vt4ieLvTEUnb6hdhfVRA5ZBsBRwr0g40cwcPxEmYy9BHOVOc3C7u+brkhfpEVgpVMYw4rM/VCLU
1sEu+L7QdfvbPKohWZ+ngd7rBoxuJLZ9FzIlbjiCWmSdkIilEY6fybNmLUufpCobLuv52Urm56kJ
6hihjbFo3/2KcPs32PlVUKEpKe88Zn5BmH43+cnxtT48IIRULQDq8sv+ewMu6Ln75kEATpH5rx78
vo8Izk0mX/wmBk7QZhYLDQZ5nbikN9ahm3vnWuxaKJEZNfl7G8KUCbRu7AdHoA1u1t9QSPL+9/DV
KrnBe0/aABnKnGka8J0ROHcVLEr1j/ZNgCV9ZHn1lWppNygsGakmRBpgegijS7Oxxw4Qke+1my3e
3SS5BMmfmOAMrPWY/RebunavpKKjcCar11L64EOGRo+u2koyCBrxHKGynSnyKTD0x+B684wjTb9Q
xi/hFLAbyRybN0HxPT5S81jDvndhdZIX2vqM5Rvx1Ef5l9pB9fB02HLsr2som1pSNv4MEbgkRDs1
i7sjMzTpu0FALB7134zdm75mokz7EPUvBCg32LJr9cUa+9fSB9due5E97f9gaxtPin4EJgUDzucl
ZpRriX3xuxjEoM5NZs0/sLq0wezuaW5hOq0mmFRHRbpmdU8j09T2vNhVhh5fVQOENJPm5RiYNtWA
vk6X7PIDKyNW/oHfHOmEGAakWD/P3HbXo9huTwLLLI7l3QlQBpxdPn+YCmcaw4luu4ECx/4J7syr
pYiXygZEweJ6MFhLpaqAWFQGtWY3lToqDlf5EpHRzd/U+rJHpO3vswxnjoOT/8et3mIvg79CUPtn
2UfdwqUCzy1EHDHzyhBiWSzA6IEe5cAcsXj/eL2GOK0nQ6xSAUwGiafoHfqUcjU7k9d1tLV9+cmA
UfNl4VmRih927Sv+/2oufAeLNuNRNgbT/PE4g9VHEWQPJyDoz+zP8qS6oAMdWTphmfCxTiTKS62S
zJdiP58giMs+71pPYnwmGNG6WgLXDVY+qb2DN7hW1FEaLxtfaqErGNw8DWvxU37dR8bCOEO8vWHH
hAiOGfLKppqt3lt1Io79453DIGb8k1nvopJrcdpTeN9oOfUN9FC/QaGgdYZ7LwheSGfOIvrCtphX
WeO9D1F7kwM3a2lOvu7Xtfvl/qv7og6yiVhtaaJ6h/lcmh3jG0VdXPftYVlbC0RNpsWtUqNm62zf
PR9rgSugnmFGJ5pz2GRvjMWS+Ds2o3cQ0EkaC23u8NgXf7DAHwFI0ZKC2CSAifZDwpBEwBs94OTT
3Y24A1JaVTDDZIIdVSluzYaSp6zkWbRyFbCZhZgEXIJgETG1pE9FZc51qC7IEmjG3dUU9kPMjPDA
jRINyvVJ0bo2izDRqxPPKETiqx3SfWs7wLvlQhCWngEI4eZSgRzBVi/mHKcq3vAu7EKdxIoAjxmc
BYelRk5jwvK6ELWlOkZd5/gjtqQbDGrZrgHTZtzwjMAD8jQuoq4TDFVy1YPD1lE78kn9seQscNZp
0TXF9vcz3VlwTKs55/8dQqpY+eK/rrgLiWnvFVZeSEIeLPbJvF3e+3KwNtVAI7DxaH7A2skx74sj
wlnrtOLCH+CKeHYfbaMaTupIvuPmpU/meso26bB+fugGlNsb1mEVd/b0NS++YEH+seeayzxk/FAh
EeKlgtET/qpBMGmzOoS7NmuhenO4bFHicWDdpj9sJz/Eq9LE381efvSeWKfhQ0vxBkoTHrUFV7ew
ya28j1GMJxVuZYEl2hF7PXs+hqnheGyA6zQRJ2OzndD/Uhyds+hifXFMyPNpF6MVEuLSTDG+z29L
U2eH0kX2eZx9HRPr7mUIeJVS8SVnbDVY4LVLr+S7FCWiSzkZqwh0cVyktPckva53PP8LYgFMzO5h
rMvDvKxputAR9q3HPFSr1Ucm0sN1J945WNZcVhqE5M5oxouevSyChvLiKB4KVzg7Y2NwWqlQxd+U
sTjFOHwbUV/P8bOBPkjudF8BEMHvx0+4NjC2tArIAdbwnAbWnJeAlhEV5EcUaxxQV2e+WwTP5yzz
XsCq/EepaZDaArrU6PoFO6BAayK/OSdlKaJ5AZTyIkPTkqcsJzeUxwhK8ezD2eEGT4DeyDDzQG7b
owC6+E8netI/V/9Z120CzJjaaAhpE3Dar4fFUvE0xfdCUAPEVS4aorAb+DFVv4tohs4YPGyQJEBS
jcHLB/WvtTkrH1vVcVvb6rSNDVUu0aOoA5sq0vETfsP2hu8iDk0FKM8zLb+A7uOFUuMeKfyBRXSd
evC7UndypUCXy508RsujB3Ytb3RbzTFzZGbOlEreaEzJYemIMl2lFzJYaWiwzOHFdlSVnFlrxi3s
QIb2rAzVDUYrA+ZKlF1MO5NVq4TTEUeLzwhD16SkxDrHhBIGp0QTwmbfZfx+pAPdcqefGgBn14zn
9xTpZpsWg6aUCqRFn34EAto/ruZDB36bRHJeylwSLWOQVbPcOktflyc0bXCKkolPnsgNTDDgcyD8
J/kWa3r2yAnHXxlW5M6V/l68myahJ++twZMRXF+hhQJd8MPXG06oUVlmRlWxnBsY/20SL9+KJSHL
G7E1/IR7xQ+I3IFIGlQpTQ4WiSEurv+lj8KOygy0+Lv2YMOijkWUVQj3g5r+d9d5EPx2cB/SIpR1
yu3/Cz6EEx8JIEdw8IJFrBcrtovIwt/GZkCeKxp70UxMzHZUPj7XlqPzaWx6yraumHSEfMpDW0zt
fuHwlmsFWai6tR3ZlswiiBAsjDW2rh4mTS2PQxl4MlJn/wdU12GDhvJoYJk//rwVHV9QMCFSlvwQ
s6DKntrFUJwobIDJ1mH+g9O4Q+cjcKWRGdNR6OtlJpMGDEoD8k43XpLLhoW4iMhr349J4Jt1QZLN
vzpxWvCiN/b+a2hemIZOwI/nsY+/SbTN0Qh/Q08khTICvpywRWZOF9hukgU6EFXtz+mP41vZVsXa
gCtPdtLmFGjYjIUqywB5x8KJV10DhTWqkrAAE3TTrstKGdm7xW756OqypQJjfedLS9kdLpXHcDZv
xNdBd+pgqoNf8txN/u41+sfQqBrpAJgvqb8Cz9hzgyllaJGDqPF6IAegyS7YXCITIGS+g2lUhfm/
YnCVI6LeQ/4W7+Nca78A80+LVwFJehu6rPPgaipSqLtkbXSouEDC4M9mYA9z7iABQoF65BsbzX1V
BApcScDeKWCkQNwpNbBceEmZIvc7ZtC81yy1+6eSCt/1E7sjn+4gOH66MvCK6/+9UPF8krE5i8cu
55i8YtSf9kNPPvWDXv7KmmBZQA7ktvyeqmgiYNvEouYfbEXS3kRiLQHZjqzcSOKQq6eT19sQdZ0Z
34gf0R33/MPQ6b2SZqROkgkxStYZZGMuxqIr6wJ7Hl903JJhubs6QqoJvNJOEncOxxyU/HHN7P/w
fpNgc45zkphQH7rH/p6GT1ik9aw8C5tOknxv9lYwzkMIH2BlenM+P5CDPS8pb+vcCp8igBDh7t5l
XIzCeCHIQHgwv4u1xaL7YiHamWD2oRkwSFqm0bc0SnE5a12rFoKOW3COJx+PpI9MEDtSyYKkoQAD
zwO4AlY+5vFiovVBPc2C2G8IxQcRUQxMoB2xbzVNCC2LSBAQILD5Nf5lzChOzU19ef2AHCqg3pux
mLQVzgK4q61Z5LhQPiGvpUTFPbtRQeME69zA5qlhG61y8ZzzoYx/XQ+WZkYVwQTm1NNWHDPiWI+J
IIVWUAFIVDgihze5zjIm1gDGSugi+oHMmrLiIEO/jY1inQd+6/1fb+amwAzessfDkyl+NrmEYV1R
/Ttt3ihHpnjdtPw0+9siF6g1WyzqudoSFTjJrjEdGVZwmiUTbmd87+qX6PYQbiFZqigioLI8/xNf
nPmuKdbplHWoFCnvapelDj+l81ylztz5es0XrLD/AKlttO345QO5bslQKeetwYtFFvcgXBVxSF3S
rvP2k8CUd5uP9R+hEijWT7PxSm5SnHz0V4taRRhb64xtZF9Hb4Mc+oF61d0pXCviDVlgSPr8pRYQ
CrgWe9iHPygpEZ8hG10MfN0Ujsg5ednFnA7roDdFvNgNKvnzDwCvaFrpxfNc84byz5cmdoZjvIvx
wTIQRB6QadghPzUyHnD/AIZpIrjg3lLkZQUsfE4dNxIPVYNjNZEPOHc73/aVTCIzQ5/MOBrOqzg0
L9SoX4w+gAqqLuklt4TR+i8k1CM8b6T4F6Nfc/EASD7Qj8jtp1J6Dt7exHedDcincshoi3s2N0VB
kOkEaDdiKFf+hrQG/r7suvWEfE6Gf1pcImJiyfJ6j2sx4HNPaXbbnV3SoKSzrwkm2s4jT9WOm84B
wsm+ZwQxqp5pLRdOh92HuwrfQUKCwlEa5cfC5NVom7JiMfFF32CavRJWWR7/I+kq3iY+WKJ9udU+
qFZ15YsuPUh/adzTw6IylpX1WEkB0VOL1lgFP0SV1AAtJbBt7ZUTZJsTZKroTpki4meMPymNGvOZ
sScy/8LoK+W4Plw8UpNdWn2k4WzGmcLvctfKZ8K0dYearZwuPLwLBLHIQoyMQAJrkPd+L23b0aOS
OVbuaDHd+W1QmP1GVTNpZZW8lj9qXZTZGAi4eOLsmtDyMqShNrfg+raRVi7eRqCPFmhqUkGzDmVp
vNr8Xa0IJO62hxPyR0cr42sznfze2ncgYunASZHBHUZMIvZRkkLV5xX7hdoRDUseiOBWAeYRDI2l
Cs1/UlExei3aRiUto6GJKDLqashuFI9q5yZnirpuiqIKFPrWEw1QWo407Hqb77pS3sb/rq4oli8B
fMxD0D9F6AuotF4WgpSxI+c1af9uMFHZsimBMyoUDi08nd84hoiDm9JvvJm7kEELUAITtb3xvfBc
OQcHF+4v3axueWNRa9/QUlUp0mu7eYnb4I+fvNnL4QEHJT9ZJU/iiHJyJKF2TK4OGCk2qZdY2shW
5+y5ei0fXbYjny7LU8DONy5AAjHHOGewwwd8P+OdnOK52/0ZJ/1TlLFkht0s/x9okxzWUFSvQEqj
TIchEIAkvwjiu3ZN7+uBdlsFJafj0mNY6CRMroe/BEnTh5V4XG+I10JfaW+dERg7YCbLKdomSYo+
gzL+mRJu3eHn49C3HduzzN9JBI/Blpr6KEhb6zv9zNsJwZrf+HT/FurPASvcA+ASNwIFpxRfF6d8
wMRTvwhQ9MI2mJ2g8FHJ1rFXHyTAqoyPWBWSGv5uduUZrvbN+jJCC5g85bLtD97zuC0WXCMyhIxn
cQ/JSvwgLeWkBiWg14Y3f3Y7r0XYMDkCffOdATl5G4SeXFcrajj8JTgV1mRn+pLFQT8mul2ovQSj
G+PVgAFxkKfbQ4eprKveLtxvQRVuNjECIqwCkyrDsWvWT2Hqali74UoqPErLyAXoPtgKO59P1412
lo8XMSA86EYQpdkvJE+Und5xkcRm1pWtkZrlZB+3Clx3r/wDhjLmlq5xArPNNaSqiOq5rgQhx2i5
fToveEoKqsPxCJhZMG4qvTZQA5VU8SP5K+M+k9b9bt/1fChYrhf3dUXyiReXfeXMZL10P77615QY
LM9wwC8/QT2h+RSXNVr3iaX57+kFhf3egdFzpPjX6l4JTR2TF3uyvVNNY4UTlCM/uv8GO/M6EQAo
kb7BU1szKOLqQbre6e7N5Zuix6QV9ibxC2twujJxSlHTyIvQK85erzG6rt901uIHRZc03cpXnG7o
jOlHM9rzX53zTii4PqYA3sO9Mr8lvysG4c5/Y8mkJb1XtWz+H4eT+xIdMBtBB/slC6+aAMKbfRp2
nzIg88SFvHmNmFZwon9tIlUsKmMjx960rc0JNzVoPNyRGjaFqEJjbqxtigOlMdFBYW9sifia97i/
2nAxXHTrmCZu+NTYnQaGIMoxZu1QnCOJNzSJdhY+yIan2tWB9t5J7z4YLb2Gdvduwu4HoMcIaxRD
HSLScox1VNxYOfuCT/INvHr0lKVNMpMq/qW87AcCNKOQ/WEIBE+nL4gPX7URTGFouuhRG23st8PS
SnIUpXyzwMurl1HQsqEZJWXp2NUYzQDj2uIi+XHg2dBUqTQ4z6H33j+se/2lK/bpFFIirBTrM0c+
LJhFTvNdLb1IPLSRCVYarKyC9sy8yLPW1A5vmopEWhk1bAXDN+lLMnyxGF/68zlehUVFUVZV/KEz
eMDD+4pk7D5Q8h2V1fLaB9yR2YYF9q1RBEFD6X0N2GyL95B+F9Q9aCt9Aa9NMvYEyvZrXBKp6sfa
GoSqsN2Qld8DB+/+uth27hORIaaaHVjZ1osdtrq/jchV9FJ/T1eeKW4MsiJc7pQamyRJElWh2csX
SrOJ48Qi2cZEgFp3DaRSnbo2Tlc3AOZmDi87v/6XJnXQFs+pRMfGSjgOLlno3qspPJFpYj5qb2xp
gQ322MYcOgyZuxU1ngW1B7oVq9fcx1qHCHVhvrbwMlS0/IExzpQkD0SfiiAqZC2VWuEYbylbNYXP
vWY5IVn6zvh2/NnA54d63zzqHv4gCYi3O8FwkyIHlBtHH8TivwcDNGYdAI+6CywyN/DjJBNom6aJ
7aVVsvObWIUeGatXkx2dtsUN+xOxz4OPctyo5dAFOeDEWSm9AIRJowxq7lKCv/JL9YOMF+LVYYRN
JmuJQA41Wkxd1JqdzXt7FRW6JKKQFFbWgsyta9MxRgsjJQf45DdTcQdaW/fYhUJZIzjpVH+SH38k
wV7Sk6CZoSLO8lg5o1UkTk44Nzvk0YArT0eivYrIh0u80DDO0dHwBH9FtnTuuPaf5F5FiHZrLHVZ
ivHlrjG0QB5f/VsOUaIt6oTwlVz8NU/pSk0tGdn5zApE0Om5VOIYdzarsEov8rwgqJQublAJp8e+
PU+hbXNvbwiQmsGGY4d5mbhzCQKFcp8fMc0CKW4ClwmnxF5yPsrq8PTYeGdhoZLoZwuQodkRTJXu
u8AOpmz6CU4HAkIs8wChBtDnP58lK7rvwrmKFTWz//5oZOl4NP4XoMd+YqeyRStWkEl8XCHCu6L5
atf0gLwI3wRfmKamMUO09oUapl/fTalewG5IGPzHiRO4P3wiv+yy2putDdDV+yx3ed5ZrdhAiQKv
uTnnZIXdgQvrD6ESI4O5v0AI70VWoRDVPC+0PltVOx+NE1aFLkFh3Ysh/383gJsM+6rLOsYeznuY
H6j+xnj8XSFO5XK7+/IUYWBX5rvgUpIskrVg7iPFQm8NphpnwnYHuYhRyYdnv4Yp6n1gyZbD6YqP
YLOZvVder9b3PMk2/RJPZwfcMWn++ERZY8oN3ZNICE0nEwq5vZPoJDE2WJqRv+laY6ZmSqzI3xKn
FqrOX8161HnrN9KpX1D1KXadlYEv7lZEJvIgf54L/E6FrI2WmHWm2x6eQ2LKWjL9tGnGJIouYe1e
iE9RAURHexeIyVsEFxP3Lva612Wg3b4ORL1BthwjKyG5PlcXTZdSPpQbgf9L6ZyBWS2RDGTk9smJ
Vee/BOo86V593/j01wVRKsmFrI8xVQNeajRboHEUtAL4T4SjzgbTsAgzjz1QDnf4cc6h0Tvxkl/F
vO27owFCs2tgISMKiWlnk14QVR9auIKWU8jh/El5lA7P9P1S6msoc9PlprU2wJbDtPXoYWoqRaoF
ZdYSB/IqJK2CKZHbdJEP7QcaJfayIWxdA8bob0tEyBo9LRnF9ElqP2rz/1qst3+GksegEAGlhuzY
q5B4HNRz6ICBQ0TaHN3Oxiwu6GLNV7jCxtwOM7TIYC5O1vtigAnmMvW1yJ6fodfWLYo98kRoF0lg
35i3BY9G/9fbcfxZSqDrwnOxZOf6vCVOAjvp8t6Y6hs0slWhqASDDCZi8cJrhaODJMBr0z2GSdGI
/hPmIbeOQXGlurCnT7qu246Z8IiqsZF9dylaTAzpmHqJjN7SmftvuWMRWPsuz5YHO8tbLgGjpnoJ
y94W4AJcWgnpaIl1/hzB1ACwSoBpd6e6TmMVQo01Mz6k1JVm89sBU96L1+lXdNU1nw7gU5wrKHNz
6HHq/ANnpHEXCYaKbQQeig78oVEQB36LPDvm16K5qGCefXtB5TerL4nALXhwwC9TaiboI3KsC4lh
US71NDxsLI4ayVGc+AEzFXhgJesXOSmxNK4QXYvGhTr5WFZjQRwqV1VattyhKiYo5hPiy8zykzE7
IJ3aSnKXZgdGu0D3Mi/+fnVODqEmaq/bI4EDNosbSI9rxdKz9vEYaeC+ogivNjroSlwEhNxdRjr5
R6Ma4T6NL0qQgDMi8DefiDJ3GPGSgXUkJ5DHZ7Bwj/6YUeo9j0uwUfGma6QD0PRFO7PIu+TyxXA7
3ndXlYYzI/3/p+eam/NXpjSyMzOVxxzSsYCGNa6rRSXwMKkevHkVS9MztsmGQm7iZv1ozjQXkQz+
aEG09cVgZyXWChjVYIeGVcjBj0dfPtoFIwtYrtc/j16CSPGsbiRa0twxD71oSiWlfwDBJeTThWb4
adkuga/0zRiS7j7XcChg83BTAgxLSp08qlKKouGcGv54jRiaOMwgE14Cimp7jkcbpMbxzDEAdX/1
eZueHb5QlKS+m8KG0Ps0I6mX41b9FbKl3lMb8FCr7tDgedX0DxpzNk3Qky1+1grb2GAXhi3f/X6L
er47N7yvgHzHx8oTVnsCuZkwfcFdNieOo4v8C1h+ykj6arb3JaS2HoFG0oz2+MOPS4qsRUNwltBZ
5WxMDe+8KHbSO9eHpNEuubQXoY7aM+OLO9Sy8+8GiIMgB61+eMOOkM+cUUuSM+59QpqsyUhyPtDG
lk6Uq+6PipKsgY8BhT8Drd/2FffgQ6Aci6zDP6OJ2VhNK5zkKwoUK+gLB0l5eS9a4nukmKdHOf4X
o3yAvqSHvy3Ivjk7QBXyUm+iek5mHLGOILYECAS51GRUFWA5URxrctobnZymvTyaeEedFS9Q2NC+
sRysTvWU3QQ0+UeA26sL+gmB+5jhu9f8rWB4/eg/VOTnqZFMqs1cP/xL2hnHLGPmOynqYqpk0X3C
VhLpJkYR9ky8bC77XmM+T4C1lEcjyjQAE8gerv4fV7MACvrOTzn7FqtJsRQJAByIDeyuU4IKG65P
2NclSkV3kOnEs5zOtpLmw66Cq1o3uqww0p9JkF0qz6ovgR9vJvh34Wl/E9zWcmI3Fd0HKjZG6409
OYM4VMpl4oI6CbBZKyXPQhKI6CgzKAhfeIjm9MXrb5debqo2QfVDPFwJUiraKTMvssALENLS1OMd
QvwiOsA68+4zR5lWAXcZP/t8tuXDtOUjCdoy+ZrXFuF/yh9/g40/ieYVUc6A8Yfe0vS4taSFvA+h
ggYS8OzfoHEoo8m2Y5riqCZ3MIBNU+L4FFBvMx+7cTpSbIOyO0fByaymgZynqsM4Sp/jhvO429JK
9SPL5xNbkTjSjhvBvvsf5qw7vrm4SGPCIqacWID1M4yhASAJnu9LVxXL10UuACw/aPM7RaLb2Z8k
F0oQD2zOFzHQ4ao0nTe3OSLKz5kvmnAntGOLaLDZp5oLhdAelhVPQQ2E3kz+uxNmFdzFR5j6SmwV
tackn16zsyGbC7Mxkeqs2bVpNkWRWZNjucY8jmSmforE3mg4ZWBpAqAbw7buzr047ePoq7Z/PuZy
KI6F7nZukU/0FX7FS4om6Km6J1n1tWzSl6vKZXti4buxO2bgRM3rhNtS9ydOntgMDF4+IGBYkgdR
I47go4+r3sdqmQGs0BhB7fgI3JwJThl81Ft/iTgznt/5w2LFn9m7qOqpH4gFkhjZWpcIeTVF1vWi
EIy4Gdyc2W7CGyhAtgAxrJoq1CrnXfhJZ22XDJqiv6Yl6JnkhWUeDRfvvGaf+9PhtyMOxnB8xmOl
5ea9Uc9+htTj7f6Oc0Z2CapUwPepeearN9w4jNrr0rWZD3K3otrn1vBWooLhU9M+vy9T4Z5FG/5w
sYIp5tzS+pzh4+WMrjYRqPrM8IiZ1OgfGITN5Vy/9vwOW9928ANrDbJXIJqeEsafGqtawni8o267
JKkKA4rN9rtZgOdoQM2bHqVJT6YPKllNYD1Z/oAzDM2vA6Q2gw2ZPVynO9t67OKa3g5i9MgMUyzO
u9WvTxrrg0+ocPirbkrEL/3bdWLZwSeQ/wbHAYcKSm8HgBW5fmKxiqq9/MzrtNtN1wo6nZLIANf2
G7Cpsstra+u/dIkAFp8ii1LclJCK2mREiwXMybiQZCNqPeX5siMGZUuWYdnF3MdgniTk77Nf9WFu
XEa+PzgohoLKFDYcOSGoA6GYkHaRiJQx0eHEjllU1yh153GR9JZyNsf+Iy3F/ATDEIQzzVqnihH3
eUtLa0W2LuB5no+QkyyFW3Wtu53RCTwZR7pdBl7eEusAUCtQLqdUuA31gb9qljr8CoQhQscuZ24O
ZQJ2yAVZjCUjTReaZMFpBdxZpdvUaw5F+3ts/3i1vGdNSDyg/dHWO+uBz86zNirbCkuOg9KuxU0Q
xXCosM2iF7RPZyiOtArzSCqdDyJBKQYNBbDXLT7K58bsHmprjhe8JAXpZWyLbU/QlEI/hiVFVcaj
byy7+3qQ0yOK85mSVoFc98nFOGWL2apWcnbOvs1/+x4RrYb80n/Bh8VePJknedUWSsahBYO+XT8y
HrwgxkeyBQkB5yi4NRaKbl4eHcQruonJLtpsYRZgn1Elxyp0tf91DPAYPM7+A70QlwPUJkzQQr2m
TsOOuvtkPAabrMt1gMhgYuzWUBKZ2K5EO2bb6HfJc3f82IxC36nZoUoEZH1erHHwPbFuQo+ul821
nSf8GHuvdzq+2rbhShHZx5X3IXzAogw2e9KC4gcIyHa8acplIEC9uRJwwuA4u9raoUXLg5fjjY3n
6UJfcE4ZpOSEm0Yzjgb5hc45SJya+ZJgOtk/XbW9ksHkdwxi0NC9B5G+gK5voFCMbWl8gJSz/lTb
mWaT5ru9+C3SN0FaGMm8yb8sdxIJNp3+EJUQapMkbK/DHCzwSynE1S1ewDG+qilZ1M6lpxChfNZ1
/1tYXMZp4UfeTMNj5olfjch4O4g+E7c0VEFg36IUfUjbTTD4KKFhLi+Q9NSFwRV9HtgU505husuB
clQ/iYgQeMqM31rVoYTUwqbmmwcApqeyjV3jiz3nFDbfnjOL0IXql1VU5pvzPSNvSXrzg6VLZAIU
UqvP0vwDq6SuEYbx7hFhP40GnsAr54rl84MAArA9TjXByunXdsCad8bOpp0NAtsLd+r+sxBQxLrj
aoo/bchggf+tGVEKbsSbUXHy7LZM/OGL5bdZfzbzeZzhphpxz7P30bTucnTaxkK00co83VS5Jzxb
Nn5t3W642En0aA4rWSEPA9JxSBzUJ/zasuf0kZGNqss6FoEGbH5/u2ufIfzmA9JEVWA27XjWj8BH
1JM58w7reqIOm8Cn4mt45m4HLsNzz4ek7iy+YLvI6c37gtt89udl67sY01GqCUX3uSgP8XeXgJgX
sKqHCvchiAX1uaBf3iFE+nbCsTKNu0pE138KWOy01OyNEqILDzxsYrYKm68epJT3AqM+JCikihsh
M+Bl4KaCrewsbxH89aUqNZ/TNxw1f3749YZiyS1XJFnmkjo0LgMQ+55a88qkOpbgoVbO/4j/EVVN
qCdxCDdTJkTJk3rgZlwzPh2cNOlK9PNsxV0TMzpD+C/kPFB+ejYtrplG+7tOOZoIsS9EiDmZUCjs
GUw/NldQnhxqlw/WGyJTEEPZ5BQVR2lnjzPV6KGDOMJDrVaH4F8s7F65GHv9hgr0q4qMPmXrVabJ
/FEvEUqCHklwb+gsWRBe9Oj//LtnhsF4oGapQATERu/c7YLvmWfNTWhEf/S59YEVFU64ztyF3r1B
yjgHU+zxrneBVEckviKGpOwFgPC7LqqSTx/ZmCWk7U4xi3kYORiiXlmxOeP8aRTI4UEomUiYJ6j6
V2RBgg2HpES5SXdv9wVIZ2x2L9K+thgrgLtavXVhDW8Fn8bBpyADjSTmWDrX0lUUM5n4TYt2pHd0
1NKJWdk/TE4lGLm7ecUcWG7PBfoYzeVR1LLXWH2Bke6v7MYHfOgo4T6z7gh9DU7zJB4l4PcTD5xu
ZIDwPekdeeggJDZgeUHq4voTlAPe6mPKe0ZfAKMlhWkMMlBYvBHCcVK4TU3DhUdWR0KJ/hLmzDDr
Zex6KOGLSh1R9zU0IuhAonOxk8kr8oAEfRf9ch6Fr6uJLmxEXuOcQPIpFc3v/z9BK7S/F/IqrwqE
gcSMcQlheh6TQ4B/IcBudiHvR4XNwpenA7aKk2we57sninOVMKp8Lm0yqneMbEqDVXcqCeOfsjFe
+Z8Cce+yJOMt3oLPVpM6ZCCxWxMxT4O+eVRIObgZmIXZdDFw3m3j0W8K+PtXllSDyVgmNoLNz92V
/RTGxjF2B4OcWgazfbaxmZBhnAP741Ylm5qTSjDud5wzKpZeGR4TF4Lu7hAYNUopljfeMxZTCXcT
U++bzROWIFYP68wHMR65jpHX50qN8SN2K+6owGMZBtVpv3tVDM7GJlYPwWJbZ5SJcUbFQX8J3IRT
zQZQLZxM9dG5cLCRmFkOwR6xgpAJ0nVE4UaVUL1BiDO6uxKPrPeyIIY9uIfebYaFybd+X8E+2Sp7
R7SDKWJrDDjtCeS7ZmYSdnER0gXD9flJEuOJKYvUfHOqfAJoIdOgXeJ5vB+30SHshiY/rGlFKrJE
Fee8V7F4/NaucAKK5cJvRJMg1ya+AAHm1aUU37v3479rgzPs95/Xw4dsEXGOCLuvTxIJBgWwjR5O
gZPxW+1FF/LkNEBhcqQl0Vhtz/FCN1oAgSkmx6aQd6y8H3pAYSoVGxFiBiguIrD0d2iU2rqow9XN
VjtCDKT2h9bAzzwG58KKf1+qxMi9g5JaUuAtXHKnijKayDUXyL2Wkpt4jm+RSuBlnzjMNxbS3Gjx
h8PXBhJt0FnOZqgq0x1RHr4MIn3C7kjHAGXhjSKJNH/XoaKObZFciamcZMvmrupOjNIEg1iQaVDe
8oqagmSG7ktyYjPmzJZ+nJiv6eVnkw0Am3cup6RbCe5BNyfGYjpPO3uAgATaH9ZK2UcOYk6aJX6m
xRkhBFd2XvDDxvaJ1hL340vQmrIRwpHAhQnIy8hzyVLUlHwL6ilBaJuwk57FxXNEyCRnvn5Bj0x8
7tZtxRdCF+s6ICN3JVqs8LgxnQPUBq2GQ0ni1CPfniIX8i6nlUvxHDZIeMjIzadbNdojWbbF/Jvl
d5+Tvtkww8krw2S77eGm1QkThkhClU7wyKP3tYenxdCmmaKYE21/ZjeKw4Ac7ugNcnYoIA3+QAk9
ENwT+Yl3hRbIBsdW1eZd9N4jcdbw8mALNjnKot/1HedLz5+VDSuyqMc85qIdx0gyuNc3PyRtkkFG
qKSjl283NSBloL2s4RB0M2vJRKoFIGSk3feNWagR6LRHJ1tD69TwQjHZckfL4kh3DF3tXf2YPHiX
gtkNjJFeGTSO1DPRUZ+0FGvL9oz+hzKe3GUPk+hpWYcui/Vg1ykQqbsiRyPZt1SXGEx1GeJDnJ0E
aQA9lmxInL4FZtMGeZDCvy/KEQxkk9yZuFCGhTzOWAL7n/zynXreKh/DebR8iQYOnYuVEL0g+n+a
d2fg+teSTQQsYjsUawKIj+3kZXk57PvTcFiHamY9wBrR9gfpVb++J+j6AOryCA2lMEmG0TXhUePv
/Atua7+A8tJzXp/ZbACD9aA3rwCzMJBm0NFXaE/HjB5YCfkNAJyEh4IkBAenCzuXRyR67jFGluvl
x0ANBIy9FOYgBhyj26gbLdGAVNARxsG/p/p7JEZyuATEhsSZ3Zk5hlehu5MGIPVsVVK7wYBnJ6KW
oyBsqM3jM623oQONDLQ6VyQsT1CRMZtvGRYuJX8bKi8KdqXp7N0xCMU1Y8JbEchH4gJIIjJdQ8eA
NaCfx2aBhEGUtLZRhTDk5P7f2phNgSmigdv65FRmcNXldAz3pREONAfUBuSi6VyYlyr6VCTgWW7r
eU67GKalemQb3tebEAdCxMkRzACLM9o3KUMoCnRNidU9EF/xmb5k76zEerOS3G3mNP93Tf/xg0Ra
cTdAM8a5zk37kMdJsN1SKEh/xbBBkqOI2Q1eyHy55GJ62BsZ6NclPmqxPqL1jwt/DMRPh4xNIt2y
EUaXWZ8JUM5RRV7dutoVN61PmfLi5eInOaY+MAVc2yabNyo+ecNlfBfE+qG9h708z5pq7hKo0n4w
xw9cbpTOAMJV6FMdbheqy8RikjYQEFoASlKLYfBK2EKmWaUB3g9MdgTqndDK+7LoWyPtLvKA2sey
8aV6oQm40PEsPk7m0yXJDwCUbuGKaoDi03kBY/3fvTzDxH5mvtr7LkQMh3U89G/7fSxC+lC3blxR
ES4xyVPPQNd0SspT6EyALB0Hpg4/5rSaNPz/y3CXWtqXDKD2Q0HYzFj1EscWvQrvOAFHPX/HEPXd
vX1pK/Nfqj/ZPgL2IvDNavOoz+0o/OHu1MfHuKm9UWqdU84HYOFn7fX7WHW8X/+zzKPXvPI6aJyL
vc5L/SzxJ95HXBJUo0zjBqTYx9y8f8IlMRpwFcpSID2lrqdtLIJnGN0EQ1GupdbjrqiwT7qL2ymv
bjS6CAiFgJTd/DIylVLfs5J5nR93ZIadhjU3SPedwQwTFXSlkHbkY0chEPkcb8OdXkckU2WiHW6l
WjJNfo78CcOOOxrSbtWHSVytAOTi4SvmeXWjdkNdgRGSuCEe/b5u0RS9aCH7VvL/BAnOvpJFMq6T
lrkKlROck8pFVm7TX+RAKxWCR9XD38Et0LBf2sUhdLQbj3kpfAIr4isW1tCxCL47ntLKIieQc6or
TTmGOtnTxh0+ZxNzYijRyfg8j85DE+Phe5OMKmtNZlpQDLaOI4B7v6kQeIBdRJRAdgzjMO1zxLvn
a+UVlcW7Y2lJ7w0aObX1ZTUCgKov534hooZNRcCfjPutBdOPIfNy/Bw5KfhBIiD3vF7+j7d5P8BF
sZudpyqppko1M3oTdK379h1txYkjgfQSYrnDNeKyWmGEVzIGEN03lQzkOWT3iIA4O5Q7aQ6xb1if
J3Dcykg7E4Gg4wB2n1H5HROe37JZUfUiYWthI3w9NuDPLJWPV1YpuH6lFfMhihHqzzf4EBQMLWB2
t7vUyNWhzrRt2yiEUyhFO1zl1JS06qUWkd/BFeNQWl+Naf0EvM2zJcWWKQjJwCPZkuI0RALutOoq
NiqSrUTQBeaWdHodhh+PwJa1TpqWpxG0lBIPlgpT4fSf6H9BMolwxTThRVNGBPFp4h2X0pOHYYL/
khpTPAR2uFRdeVP6loHCUvLbz8e8Sh2Q/Uv7/3VIN0aPy0pTvmCxpqMZq7Jg7MMi6/jWsfuRbphB
gNRVdM9F6RWN2J2YsHd1LucPGSnRN/PA/NkRgxxzvxu28IOwkXKFCyxqFHkfq7ijPUMAyYBBUcBP
xNt2iCNThwWjIQx+4ePqmJUdTajEgthyaVpaR5C1v+q3zA/LCTzUZae888Lirn47YAwfCEoZChzB
VY5t0bL7kZ5VqWGKi3MUzJqFQVt7mGS4XwqE50GSuK79FxQa8EUU5Zh7dzD+VCdEE1QXG7ofbXfw
hG3MxctK7L7cEVGz7sYWmcEdmbDssvbOxZkHAZnX54xkKcZgdlIbpDbZCEeh5HDY1cv84spaluN1
+cWERYzNH3MzSQrqrG+UV0zaq4Qk861Pr/jycK+7NIjupW9Jt45ThoNzjxlhwoGqr1BAF1Lbf+Jf
8cJKIH2L+cqzbVBVPUfBEZLFyhAaBTqPimUo+ahVAV8IMpvVTLsptcRTC2LiQVXNzVCjKOTLiPbI
IhoSajCjsIY7PaMwIz3GmCGCH8usa1KHkmukKAkVNQouw3CrSxs+hQPi8IC+XzjjK9deSPzXAs/H
tpefvAqA/yV156ZBvoLLVS4EH5SlKo+v5f6I2CslNFWwu13Ftxy7qJtZJwkHqmOpLD4LjF/Fdu4U
/UyIGtY/uBNukE9JYXw+n/nkh6WTnVAxyiUriWtWY5n7oMWgMjlzUWaV6uVN+CIM3rtWIK/fZbTt
btOTESmNMiD00CE7IuJd+542hNuJMBMMfdSB1aXsBkwmaAJ7d9cb1RfPle2i2lptCOJA/yrol7E8
BYHusNy5O5Jw/oYlG1RPtu3T+aYZTSVkoo9ZQapKW/DXiGPdjaUVYNaiWllpuNvhRj/U8LXcJYDw
PDHPtGBcj3Iwm4jc3DgEZJCl+cPPVncy+Z+d1bfAgLyawGqwv3mtTT9VD9L2L5sHtxQ16fojLJre
gdsSpHrb4l92ZvZQ+XR8y9JSRWbhmo1kC48M9D1sglLiAqAtDPGfUwGSmHTdlxZKD5VFwlN7fJSd
9/eLT97VZ5VLk4vWx4u5IJPO576dl0/2QvNoDm1sOaJGZVYWvsIV3zgnSK+8w4BRBmc/LXO+MwPx
HSH0ZMvaU7rQ49QEE0YN38CP5Z5NNdJJ019sn2SyYxbywrxjqr6szIMJkzkYPic/LPQJwynzVHwY
M1Mw/f4BHxP1f2C0IPYI12tKp3jVqj/rkvEKsiDrY+kzqL2nwvD2FJfCAzEIA8zf3XguEU2R2zwQ
072SahD8F6g6Xk/2s8LNkwtGsyrfDP5zjcuiBHXl1Byhv7x7TUR0T7hPFA2UHFr1dUEGzsuC0ifX
rRDXMbWCApf5MKpnzu3hFyjKMQSRo7Gw4dMaIf+EwxCDbL8fQyZESFFZAg9SNPv/UO0jBw5UOcSv
LWLMWix3Q4cJKS+Zsvbwu1TGi55+rFMrzy/RcMVYTf7CX+aZ0Gml3mRFRHKpJJtTPPXIxNQhpn/U
LqAGwLsvpMX+a8p5Sc4a+B1FQty9rWoJAFSskldAkyPVvmVfSfGyf2sjpw59W8U4RDtpGT6O809i
KzkMC6DPtT3SGdkXahtx7rTjDpAG9zeKUzhvQYwnvJ/F3d7iMT6/i0Mcgk98D4euZefuV4bJW0Hh
hyuUpI+/xJplVko3qAQjVdnLU9T1Ckuzr3h88z3V5eIWsPVvBaqkkf+BMRDoZvtELdtUkk2mxS9G
OgLUM3p17HZO9DBlGagWCh4rnYxHh6hx6llZp5eeNdFFGcgXGL/ps3oqeJipLSGca+vj/C1rIUqh
qVFmzKxPdZLd0LiWBsrC58UluQFHjbB9wbecDyfuCqK2YOTLCQSW4ytGA7bpVE4gGGCPg2J1A/oY
14i+gqJPnTCXszqxnF7yZQeasmqAW59U8+zC2yuav9QEq+DPaWsbX1Ocu1FnynwvsY8MYiMmjnID
xbPuutz/rCMVVLUQWcgKKpTHtmru9YPBkXhlOTHvRLzLXYRvvotrP2g7dIv74n8IerH1YfhlcoV1
XI97vU/L2m3iycrT+8bZS72ghC3dF4zHkrHCKKd1SlBjfnMiQw01DMC219Q9DMNrxrZ44uZdNxed
N5m9ZfQUNgK26WqP5B8KZjjWGjBoOZIHXayNOdF7kB1vTOSpDyg6MoeP5L5Gk8g3V9Mv2Rn0fhuE
7TcMUZ9GzaH263mB4VovVGhVfUdQZJaEEfa6D/T/ppuGCsml7rATIzvJ0t1OC4BnxiujBIfkpwnN
jcAsJs21q5x4QDimQ82xFTVepuG0bqTveZR7AZB/4KSiaRzyxjwQafqwQOCLnS1/PLSbI+OuxADX
wcwE349i/A5Eb8t63kbMjWOrqAJiiZH1N9wuTBe+9QW+mF6ZlgbhiDXrldEsPxdIaP7Ts19j9Rvl
8tSirlX4ex4M44RDZ3vxm2kJ3ZPEtDDEYN6DY/GIVyIUQBV4W8jQldRm2ekmVmrOMRucBcSEIAVg
oEC5LW+6aT80NaRkM1PGf558d8plwFbTHIpM/R0Ij6gJl2UgJw8pLyThluTRQh8fUOXCrCIQilfJ
Ch59A/y7txz8ycXUMfnTj6tsTnuVYAX8uUBEAL9MkotQiOP5FirMizPKMsJGS4aApYJI4cG+opcu
mVJFJ9ZYJ8FximTiZzxkQOGgOWNDRboE7iWgUkr5p8xyERcgpxuadLxQKnuPilnwbTLLLV/4FuNE
UukKRFFQfFw8udcNWQKtcPIKAg4koxQZVRqsp/T4xLwLXy3fUFWsR27zA6iueY+B1m+FZFxOalRi
ib+DQWppH8aVo4H9zldEU5fRbK/+yRUsWFrRyGjWezeDZhHeLMMWtBehP7dY5IUJIZzRUEH/Uj3G
Z/ibE92dc2O1bBG7O0b7YQbqTgAqdJDp3DtTBPFCuL505jtgspBLcaKyT7+03bS1BdH+JToPAtCH
w/tSWEC+/Zq98Bp7h8YukCehehZ/si4QiWajmyuJQzXnV8eeXKHmr8H7us+rKLzQsnPJvKHB+qmK
fepANDPYbAWadNbZO9LeewocnMT/2Ng738SlG/ozpn1oS0Mi3lwNjc1s0GsYOTadXb+ed7nctUM5
U/JaMDL12XAxV41wUSrjVC5Czj2JqZGXV1LHUCyaLt5aAjbonsw54Cr+pumUqpHScjPmq2Vg43K5
eueQEWZahlgbu1DB5jidn1utnX/5XeNImXXYCCDDR97r2bbvWdBHh5ZdYsakhpq/kKeJraEHsGXF
9RRzhEOUkzXuILTk0mYb+42/0nH91xvrORQrQCX6DRVJs2WptfejTKelSku+xmVNQ3hcrxyvqKE2
EcLu0hCVg6zvzGX5ZiMP0ae/B9Ew1cpWufz+Y9c+UUgowZ9TrHXbAonIzeIw9Axy+8+D8Yl2qHUe
vxq0V4o0y2yhy5PFJEn1bNrmGPsMDXOqzSPbanOwzOFBGFaGMIDHqENqAiyE8ES4cRgyD57oAk2Y
atCHzXmCH+Aq+Qun6CgZObHeQJeX8vS+9E5Cdra2ziVMYU3R1TtRKjiZBzGC+sb/upJffMXugmnj
48jKlLhdINoUWU5qLeTcRSYXWCdqImuah104teFhZWpBO6IzlsnXiJ1QBy7lfS3xXc3jQQ7nC+IH
zq7yiwX1KfnrxHbRdES/F+7LtVEnY/FgRa9J42QGHvHL2hgUdjDdZyC5s8UjaOAJJx5TQ9QAR0Tv
NNF8Y/VZzH0Ol7t4+Bhcz5WX2Xfwi9KXsfWY7vni/zbWvd0oJ9cnU2DNPd1M5hh/gwJdvWETBmVb
ZRA4NVyrandK9GeFDY8HEbI3KL+3G8m190KmXG8pMJL1xPu0An9eSMHXjGkboY5Om79KSUNbnSBw
NgrWEBXB7ikASHcGN4LVs+A251CntbSUqaZgpodDFbwQqx9vuHwpLROGX1V/ttsphpqCtD+YqqvS
rbf96vaNTMjev5gWjetHRovzlTXZnkdGiG562qfTM593diKtTbRJHHrPi9IcnjceB1cUHVm0JM2S
TlHkRegvZu810BWT6MZ+cNcgRZIZbdVvkp9eYgBbF4D+JrAUhSifL0Trk0OoMM0g5s5hL1Dtz7mA
/49GGCfd6KGE3zgF3DUum1HsiHGT68GKLWlZqrsAJRKVhbiraaczi8gbQ7C3fNzwfRc88uIzeVpS
HiQLaiHZTp3FjtCNzFeDranMDiqle3+MG2k8EAAQ4QRiFwbhzvxAITKjiaCJemy22mDOdDGsE9jE
MhPka+OOez+41/jhDvTzzFvbYZWqRq6Ol4PdwRTu8Nb8YEWWIW79cShO/tbj4Sr41U6E3jHTToqT
OwKo6DVU9emadoCpzmDIAXdsMsC+POGg0aqx4pocJC3L80veJbq0SNvyNLSElQE9r1mM8JWBPQDT
pzy/wGBlIYd4unuwEzWZ4AiTn0wOrSwhvOBEaxf4BbvSVDW+p7kLY5g5xg0ERmJR0Dg2BUsVCBLr
HQE+lmQQC9UTGg10cW5sZVE1zbcFtYZspUCwgcahhile6myQZrFKnXLA/xyA3ruKHdu3W9NIQ2h/
Yt1XsXYZ6PTPlDF0Xbc+SVP5mO16oe8ryDkxwAWgl5P7tiDjBLEMDSQpYRRYR4rBDjqeQry8eTJs
p00PbIV+6HyVT16x/63qZ2Zhf850V+AQJbAfs6Qqsd1f18vSpsEQM8Q/mprjNRFKQnm+RPMQqUPs
tfi80CkD7gAFFrmc4MZNu1qYWto+zTSpyg/BkDyj97fLOKQL5f410TFgOFJDaTihdlARc5x2CUsS
1UGqpd8otfAZP94ngLQ1LFJ94O0Ub3h4yj5CrfABP8mDOie6GDWEwiV6l16WMtuilQjEjfIe7OT8
v8pVvztqk0BdXF4NPlbCstZ+lZKsyHAQKHYHhP7vi4jV5cW1ldFWBUxO7VLppApdqQAp1+mzNq1Y
4Xk9ICGoWlJ8IP+WXfHhwOl5C58EUbNzbGNdU4nSCt5IHfUkiG/T7Hm0PqgFUBdhH0HLD3csna/+
3TejX5R2F2uBnTT1VbTD/8WKbiM2toO/MBF8UZekOjcDo8xsPDmghjRhm8GndLVs/j2hkjHL5Sg2
2XjhdeJeUgpcae5mdS3N9mHickPwt8trOiHQudxIrLoWbyq0gYDlfXyiXINSHTj2NClxQ0NVVTgi
9QChUCwHSec4Jl1k+bpXz++panIJWLaq+kiiIQL26E2gP0q5P8tFB6SenbnWbGitD+x7ktR9neho
9L3+QZyYIFzN5J+6xCMfwQKd5tIWtP3ghFrfZWIvNxULJ7vvmxRqN+48s5/4ZUX8y2Qb9feZn/6S
6+3mZf25TlCoghvDtI3snIrd/MhRYcIkV/LafsFL57BuYLvRKAxpHQ7KP/38EqxNZt90Q+H5jNuK
0WHvcoMOBaZi7VJJNaT0+PiWlsoYZsmaqE141OsecrzUO0GIctD9wU7YKD1CFAhVe5ACHyvh4dX7
NqUJMnv794tgZlGuxKDvNBJq+09UxBMPiBpr14GVt4XtqyY5YNB4my/JmJ9t+thWDLRduI6cLRDG
mdUVFsEXZX2wRSFGBoILLiE+3843eDc/i3CL4GOR3XZA8hvpr0D8nyXoMmAj5tWDmZ5KCYqfYQUW
IY2mTOWs0NzVR/m8JAeTQ6JWIZfTYkP6LLCya+t6BT1NXK9sW8UW8nd13Zu9okzQU01YqOEm9ems
CNcO8zIGe/tT/eBy4e4BB9ZoCQzGtk97FPJvzjhtds70ciMFAF2tJM1CUhM23AD+acgvJVY88fJV
yb+08UK9owfL0Ubp5T1LxL8ro9W2cX4YPxN3GnbZ4nzFGOfT6HOVM7su6IC2mRrJEUSIvo+mwNI5
me+WYSivDxEingNPY0F1OgWHd8NOlR2r67vxzVLgzRxTt9ewb+YXYhRrOjW47sqf6A2JFc20ncuT
72AcvR8IwCru7dbAyIlBOXfjEMxr+8nrkB28BlEH3Ip70+NP7X9AJKhB8eqD0AvG59XOPQDVu8XZ
IEa4VlCYIkq0PsEcr9pOIsXsl0MxoSsFGtbbZRlFx8jm3SO2xPsVhvjU0b0sTsrLDPjKc2y91+Lm
q1uiZMEaIt1y26iFFSOy6piGb92RaOJ8kKOgGyneNF1zUPT9nlAzIjJCM97jbuhC1+lnoklC7jR0
2DjRCYVDwKCP3niJggVMOpf7r6dDYbhDZqwznZPae3wtb6SK/3oxOAx2356XvA9cHm1VKt+Y+37i
cVUUzusk66Tnm8IClhTCOz8omrTuUC2WPTSlmMgDogEfsnUkwoQDMjks1xwRwYnz5SyM+FLP59h8
Cfv7boqprFFUlp92S3MjZFgzfaY/Q6+SgCwN4QBIHankKZ0V84j3I/SUIkNgg3pn4lGu7qEc36Co
bKuAM9c1ddEJfIaw3v7mK9jx/D85mPexzLTJS87/p490cFn80J0A28QzwXeNzq8TUeUjp1oKtPUL
bbeyUWFrnyrrbyzJeZDyv6lyG9m7vNzeVcJvePbJ3AuY5r6LxuE5rMruBMKphOFGH1xIpgNBLZYp
cUQPPyuKfIv7z9myIHy1bUWSlDUIiE2baT3p17a502aDw86btpcVZEKDGScdVmDXg1U/CTn6ggCT
wk9X+VqnsetJys9B4GBkRKmAsjZu7Dl6X2Uxvgev5aKJIGN5qTSR6iqek3SbJpUXVUbbRXjKmlRv
yQXTgF1ZiN7PhT89yTOdYaBTWwj3WXHhyINYDKYI2Ds2OI/MrhHiRutsCp/9i+BCKSC+PCLdFPmk
YdBsuc9XJddb47RrzWa95zWA24njSWlMupr9Qj2pOe974kf9J3sH8of91JiE6ScUNHRDdHL3mwS2
nO/of6dIFNOYW5xp4X5tJd/QBcnZC/wDmWz0RLj7ZdSQo6Ne6LRNHB0UO8Ny62PteuRg8XOvTSXL
XguioRPpr+TR6dh9uwrVkoQ4ugGM4cmoLc5xk5kp/vzCSwkX91GXA1aXozsKW+kud1hGFda34HMT
XyqMqvu2gv4FYv7b+ODiLrmXy2Id1W+xNzxjE7Rh4/yiHLrH/PpxOZ6xS8GGJxsiecoxg90ksJO8
RzvG0pZ5UWer37FfvwBBLD8zU8Q90tAPiA9sTYtJoDEFkc4N1SB4fQ4rXCb0r+lKHU8idzv0lEGw
gD6ctKKYzfpGSmghBzNGO8I9QVvPWD2mhPh1W3tRQp/CxtegQWC4PCid4exj9H+TzBvzJ4bjJUcg
xz8D5PkjnD8Q2tQPJI6r02Wx1hojyxL+j8wG7+Rak3skb9Wl+51bJuceWmuJtu9r9zLVYgRa7rEV
Cl0jLz+JOZVsvv+BbaTGaqNoMJvHsRDiIlftAqwwX85KXlAEwTm6KtoBFp2eMeFsQIseOKVEauj6
KuhFJ59H37VMg2GsYTYAWW3bBCdqKVCfDcswQa4PLQs1neh0U/NLniE029/MKWhc2IptM2v3jC91
P+UTlPAI+qfiXMMFfFH3dNUHn7qgbqJ487QLWT6HTHyb6c1tBpCSXf8TrvDGqnLLk+vY+ZQR90p7
MieD2z3zkpPvcdvk7h43kpBA47unbgYXUCTMa0JfcMdsvKpgWJEYFyFdE96fb11IEBi1JOQnH+P/
YjCl2fbSIUzDw3Gq7EKE/aBCb0nljDdofvrx8sVtfO0AE+akLqR0tOgKoVqh+htEO8Kt96kiMaG6
3VJSX+GONg2JlkKx4B648eMSjxCJ7GNF74ppMjl9VLnxfU1u0DvGiCRWYknJVC87N29hI2tWGXDX
8PnIv/kpj39ZnVY/IIEQbJsxwA1hIaJjCjZYTLu3PCucR3SP05SpUAKN+X/micHjCWG5ILdVdsM3
p/LFPO2ML5/3jFT3nXJa9ORc7r8jZlrU6MR87ydxXbstkw9EY++9n/ide07hz27CEL1KcAUYFnDc
wZM9MV6Er7v+NGwrU+hB2JqaLdqrsx+U8evWoNg4oXW2k+Io5sVjwRKhuziIbkxnnmrRpYV0ZLhl
Pr0dv6T2krzRcL6o/ea/AV+CsWCy9YI4JI4Zdx6B3Rpq6yaGoghQHfS7+mVKpdoq6UzKPHBNsdYv
CSAcjURRGSIfyD3to14fMZq3TnQTVMTOZHv6ejCoGU4ORPO/l/5v5/kZUjclX9BvxQU6p3gwExhB
DyJaciXlmPSoLqRtlW8I0tIGh9iJ0m9tEyelZfYyFW15xVaAYFXg6DmYR5EzZF107hHF6sWs5x6a
uTV4wwGUZdw0luqboBrC5MHlAiK9bs1u9pyuF3aBdLrKBXA4KaQZVz7SsL/OnJopvqHo612hM4DT
cGOSbsSOmUnSK4plbmEEf59CQy+7ehU7fAor3q3m7NOSxNtC8rdxx8rhkvjCoLBEf22DZwBQ0KXp
yFEfxb3mbfDp9wCWCu4H5Oeh/86bizRtQEE7W2qlUtXpeUZdey3sRdIT96XjonpYj9JQrWBUPRWw
rINzgLkQEltTKiBUH1jhINkrnkhcq5gvGdu5dDJgOAU/hUMprxJR7en/fyn6DTTQ1fPmtlDU4xDC
L6GpC3cn+j7i6mkhLCEvHpF0H6K0owK+5RjpZt0SRW3N5wgCszl+31pyqTB4JatyjOttKPNFrRNR
z01va3T7w9TpGvfw6sN9dywdYHosBL9jtToCIhdBT8upq+KtpkPYxoWYtAetSCsZsEIK+bnU8d5/
O4BomJwZGFjlHY0XyuXmbm9GmJVxMvzX4LC1XKTok745BvEpJK8X2O3bYKkHLUBBg6isep2mu/W1
k+Gf/WQQV2Dod2S0ZVkYq9+FOTFoIG9udZmfLOJ2ZWM/94VSfrz5iG43UR1qTET1kzIaLvgNYiMm
JP7M7UQLhYnwIjkKZfa9MQuHNG/B+fKXFTge1u0VGRNacrBuqjVvCMg6qct7sGQoGUmNQkUi7m0k
mkf+9jaivC+X7KI3LrlmC787TjIKwttOt61EllWc/MquQPQZLWvg4UYpyOm+1zoSda2s3LLS80Nx
eSnLHw9BGGngOU5VJDcsJ9QsqPsBBPQgcbS6eqD9arOJ10x7u0mMJ71UgbgmYPSEcWWcVyOoxzgZ
5LiCZcL3D7nbVrHpEMvP/a8S75ChzxltZSvNsW9JwuMDoypSYRdL+i6OHiE3jqRAyIvXK2wRXLrI
624KthFnZ94RUYT87PscbpFLN9NaoWsO6u54DvYKHfvfPgjwOktaN9ZDN4jR26cocnRAMYkI06Gt
nuHL2s852B7TGV01X1dRiX6N+D2G6hbPew9AgzZDsWMhfRGaOZK7X5HxuhZjZmFt+86eoaC9hqxQ
KdxN12wgUEScUHqDCwIga39uPZdNrEzQgNbc6AeNb4ZCrA6dcBub0mwnaeteULax4HOl+GZPIOJF
2R5SeUWJVnh/etUYICdnrm+Vd2smOhoLk3X1ePH2H+ykzI33WBSOt/K24G67hp2lOIbstA0gmQVM
5XBFJmfQ2eLZ1nG29sxNWFh0R1UZ48LNmevOwoZPxwmosO6keBQWyn2oMfwijwbfq+u4CMZoNHsQ
NXZwm2XE0nJ7fLmRALH7Cu0Cpa3q5jfsqBU9VaLXwwlCfnn2geffbr3UnedfWkW2M5/90w5FXm5q
tBqj4mhN3jlMN0D8R0rTHXN6G+wWXAzoekRwBID5ZQHomyPYnRllRcV2Klbiu+nZVGA3dxjK3ztA
3oZiGg0o7q0UayWTY57am47CARsRoUxywYGeY2vHEzBOeTF6CAhBGjJ6yX1HllZbbTvJiTlblX6g
KWnhlAqNH7CGw1aJ6Kh5fjX4opbJ2y/95hxB5pJ9Fbj+m+a5+4IRCHd/OYrrX26DZ4Yr5bi8uFCZ
NVpImSgDGApxQVkf8/y3H2nEv5DIL28Dk0B0ymasdqKijJXVg7NyX96mUq2v17XpgD/iMJXfJidl
pkSSEKjZHIOy3QlGZoEn/Nmo7Tj4KO7z9k/h3YcUem1sLTBRwWjaVDlmeibZTS4yacr5bfYcrDo2
6vTLg+6l6Y7YNSRjodfdIm5MP4Fzm7/PoxeurbVMSY/uB5Y4fmLrnk4wknKdtbNdQ3HQN1lp23wm
gLV3QuGYSHkNwVeQkCmfLeGoVB5sTGnixEbcKecQc0fawAHUcwBfR0puGa/FZ/Zh9DDkoQ6m65Rk
cfJgy3QOk6qZVtfp8iFGOhJ1zYuMlA5j8HXacdLk0Xx0apVggcoHqAl/nXfe5eMkIzZSe37j/1q/
0oOJKGpN7DnFBTSObXpvIbhuM9z92FuLR7U9kVpjY3L5PtQPQd/0LPbWUIuVram9sbsfHNdZCZpQ
e3mFrGa9Z5V77xrIf35nrly33ZueGiqVCc2kf1VqTn0fGwSwHCpqGs/YyKrAUf5TifkaKlTeSyUs
Bk2JLNvklryJ1I5+g4x78TgeMRhGa5QISPsvckMYPYNm56VOstX6YUj6Wa5gH6L7VPRUdcFxD8Uz
C8+Ohee8asfRSO5jNkxlZEkCJyOL+Gq/0WvaXy1j5A9zrS1WADM5iERDH5LdUlWlGTxa2z6o4+eH
sovBWEs+bezffrUcsDa1CgRwGnEUBQ9fyqCikByGGXdpTv2rfFBhaJIlPtGDrNZ0GgjmrlMlD784
4NOjhTw4sFO1cifDz+rNWL5m6L0frue0ufjbELuKaFCb+7meGPGlCL6FjdxVzn10ySc7c1rWLWSQ
qEnSX/k3Q4k2/RS/RMB8JDp7eIju1MwRSMcwQymRk2Vy3kKBY117aZewbhCZQiE1tzBqt5hLvqLN
eYMHV/nJqi38OVCguj+3udZL4IgTR8QwJdlLGYGWJ7dEkuuW3ZNEEohKTBrQs/oIvMZJFM6A+Zy5
a4Il1gnAds+xKU3ujTga8n9NAQfAOrp2VJ+iCI7rjKf0jccw9eLfRXv+F6FfD4FIHz6y14YKVZp+
MAimPIPCCByxM5ITLvpMeBHgpSuRlhDGtJ+kfnyTY5ROP+k4QqUq1BM63cbSOG4OBhDz4TkaniQ7
oM8BMD5qoR7s5mzWraz4RrJWuLRT7eWjC+XWMfs0HMJ6bpXkDpyNhC5aIpQuPYdOng3GEabuEcuB
pbM8TQd46Qv6vsDaiLDJVyw57TF2gPN/B4Wgf61a5trQY/UrDZ63OTX32berMnPdDXD6EApwXNeE
YYXlcsGckcnAA6x9DAKwNAP+073Mt3q+l5RZZD0qBIykhd0yoA2LsK8zkGKcr0pQEZioHU13s2oZ
KlMLKQs7gQ5YItovVUHR5eF/JwUmWQYgB2grr7qKK8YbndBbfELiN9TlefSFzFVkYllAKP8fDap+
biht7WNlX/gquJpwJ+RU/p+62F7/t4ShuFI9U64mgdBTZksY1thkGjenjtDeDiGEf65OYJZcsBsh
8PE/J9xn6qlbvHTyndQPts34E+Qw83Bfh8qJ8/DQ6mTI7ZyqZGE7FYPsuXSQi+MDDE2dfYy5mnbf
QKEM7eZGaf3nOYHq+rW44aoNiP/TJXtRi8M59yWjQ+lMs+QrLnT2DqFpDodvAJtjXGHtECSyK+hT
TZ/aphP3ApCvunij4zl/9Gyl3UlT3OY2La6eIE2aIp0ZBfDzAwDBozdp87ZOg8TeQAxDeY0wMKWz
DICiR50dkd/LFovLpEBv5xUaYl0hBnuvhP8BWBcOagmCIqDJj43/OamZXNVvjxPEqOiyKUcV9e+j
TCWvIUDdRCiiNDOxJR9BkspvjKouMFulyqqpKUnJxKXXQFa2PYAtVg1nuEBq02z9R88lH/17OjBs
GOr//S1SumND0/qDhGPg+S+6J86hyC6iAqpykhelvUw3UdPDsm/gpRLlhU62KOBFmEhRjNl7aW68
xpQf3iQvApXKw5vAg/pXkdQHWJea0/3JlyGj16IulclxfISNBx96wrCKUNFODAtFEn5ugOFC6VTW
MjNrj4ADcwx5goWjj9nT6G2jZT8R8qyOEXoCgqcgQ2pIpCQUj4ZHhCj5mWvZ2SbcB5xblt67klFZ
+8Siaoui0jZbimmKyRLXnqEmOfv2AdvVUWqEutVz+idrxcHDkS7cIMUGUeMuvdq6s0c8pNcWvN4n
yOpzslRkdeKbnROTm6Gm4HpD28Ov62lKJ5blDPWk2VjGO4bso7GpmL3vPo/YdpbaZMfqpa6EFdS9
TOoh0rMxIotfQnxbsEr2RofSyH/0+aUWou8QFziqnvN0HYz+UmN3JXz6z2wRt7ObaC+bgAphece+
NDey5T5f1KZYw5mXsjMO0Zb4lEqfra20H8CsU78rNKhXvXDN3Kon3pGtIVL/yIV49n6Z+4c1E5rS
fl/bF21OcXknpVQx0aQMvB9LGraIXi7vLrtsJ0+Al5t2J1n4EgH/99PE+BkDUfmDtQc/weR9dlyJ
a4FkFPAUPaiY/iGwGB1z7JKPswL6d5ePH7LBShZxDjuUBMo1J8/0ozXLq0sdWpkZvJ6YspBqiFlz
gzZC9qScvlJwRoSsV73ckZM7bWZYUzdgtN/TmXQh8jxOq1fkGmjqWR4VrZyxgNkcBMCgbjzVZukb
Mnu2FIfLpHML3RZXtO3mQsbV+uA+Jp4305uYIi/Hi224IOqY3X6j5r03+xRO60bCKSiJMhyFl5R4
7UN94MM6U9zlb6evva1AFYxIVlXvXZ0XnNt5p7SXwthoJCwvZFZUN5JI5oVEslmA8ETp5dauTjFK
b4xhms9RM4AQNOirtb+d4E1N8S/h+CAijInIoADPFan9Ru8XFX0YM6Ue/PVhBLIU7+ckSvt6mfdS
RCZmV7qoDJkglI11LoY9LRzTFt8awbb3Wmo/ky2Z0YlzL+1pJTbORSYznfpex2bS8a8xAgRRkLzQ
zHUwIZXvF3ItBLQnGRARNug7YCZGJoudwsVT4OIh/Mq1fJWQ2v1xr+HwAq3+QFKS0SduKmkH1/ha
EnqtKWr7vAAREOhaOD+iiiOdMDwaq2izKnN/FfQyXW+Lkh2ut8mb9Ca4CywLqpX49xl/OWFD9q8C
XXIM8zfp3HXA6Xskuh9sddVPCWJpTEyEQrlQQnjumrHlYfrxGr1VUEsbq7wehfSy1vAxtUhhipbm
pQUHXPTsgw764L6kbeyEHv3FK1lMm0JRAeLTyEHP6ZcSyJ8Jpa+6iShCe+tPZJCYvCz01lTcZ1aQ
LxztC6rL3u7IQOayqxnrlCut8KEctlzyIvZq54Vt2Dib2PN0rv5mEAPaFui7rR6b083Eu3OHNghD
JukCdR1jNMSFT2wR/olWFPJFHcjC8fYYF3PpZscsvMEqakZMUMItpRa0omx80NwuUrWIu3mW1pso
z2pUevdewGsxrlyOtDWCGwXcRyMuOZWFd1D0Vt3759v5fu5+472MW6F5V42UNjLB52IHvy2DgLb2
S6pSdM4EQ0m+L4mhQae7MRCgYkkOU1B5e6r9SWl+j3udZt1CsHWiiJk1S1IA8a8DVD06rftJIg1w
tHLsmJzs5CGdCd0QzOtjX/IaEO9a9k9ife9OOns+zKC2dlCFN14/lojOu9Pcaizpx3uMcqengDGs
U7wVAYPmhlynXEFVQdyu05rtqDtVbBtdWbikZacgVKQ7F85WouQ9WWm9+Wjk4MK7XT3X7Ny000Vo
cQZoA4pDlnus9UEKM5ylO28mFpsQ9DkOh9XsgNzFFIq140iTcvROe27D7mkKe/NMUNJ+LhbmcEmv
8nYFWA3wQ7gKLdbYu2GXMNL3GtSSTPzs/z2KTSAYR9lnXiQ6qCmum8H1LN+fHVGYXxiZyWGENdWw
DZ4FhMTFebDMq8KBc101jpw/WLUlmcPnspH4I3WOZoSBpW4FEl58f90azq6pFrFOv3t2cO+1o8nt
c8s1etjlQROIz2jpSKpPH621khZvAXQXBaUOccxixVGwsLA2hB0+iEQ29o+5ELH3bQE7avQxrqym
0RBNcpyexYkrTVeQ3GiR05ErtHYR8ZbJyufdUwia0UZU6KqbQw+5EcxcUJlGzK0tDt72qocMHJLS
pjqIuI6hCyk8hk6xysXxLaEcj3b+nggORhek1BdEwKeZ01DqtRrEWP3RBWgt2sEFIhTRw+ghQrLI
QTBi6DelUq0nolPiXnh5Yve8LFL4fZLCYpAvblrzeTqKHif6+adbd0pgW/HmfTxbOBEWinhpQm8a
mv8Y/WYoH9wKMrXZhCdrVGV2J3LpWD2WMhJn46IEfbJdLqXjDDPC7xgJXxNtf12hQS7U++Cb1CpB
WmRs82i9JanOxahIxayuR4SNFjej4hYy20A5W3bpg1Y5UCFsEqe6nIHK2HdpU4u3nvamE690fUl0
+qNoYNkfnm263nSc+PVIP9u5zfsxzlu07rL6rCalEzHS3HNmuPBd1fkkhssD01/L48m+toujt4za
Qbo5DabsyY7Kl7fJAVQ0Nv+2xjINdL4lawsQ6H+GNHV9bkHP4wNsbOqdX+SdmUcdK2mjp/fJoZAo
ac5t+3GajuDmIRia929ozeQcWERMVoIypiZCvVZdyK5Q1t+s7VVKe8c5x2yayAwXnbeIYtENTirr
K8BdFoOIWlksj1L845uJwP9ZL8AX/6Qbg3kmNCdW0W8SLqlEwmdg2OR+DfpmICF2Ln/CK93bzNrG
Vt6sJdSCxbF3GncUKE9ESt3a0Uu9l5hfK2C2tHDaiPF/kRuWh6P+tZWj3O3VESO4C+KMkRPPXwxO
PfImnIW01P8NIP4szcr6S8JEzIxwsVzgYadhmUZeeaibTNqw7x+X6LFdZiKN8Fx729Oh7KjzWR77
Cw1DSb3Gv+Dcqjju5yNPirf0PJuw5/6FoKP9CbbKYlhDyvDenb1Rjup+CoDeOrWwMYzINu0aYuvi
CVJfiubOf0KyY6IYqj6zr/2JYqW14w0x//e14vkp+ksqgp1tUoNxscYhJq+Sh5FUoooeWQ+il7Y8
JLvlgq+szbV8OYUaPu/J9MOm+PPxxRMULkj3uq6L5wy8/tzc0uywz2tNBSCzaFzVwF1mt0Dk9vez
t8Lm7cFkYqs4UC8seKnebBRwELNSTW4QCOHd52eGovcyTpDg0mbqu+EPjy60B+q81eJz9NRgAx3a
3tvL5ElGB5Zec7h9I0bnFPVs32NUd/p2Jc1JJtuWpd1AnPYcMWQP4aljC87HYRygwwkLwYAB9gWJ
7s2x/9MW6/tZCwhKFTFpSrw+cOPUDQENfcGEB07m6z0LPWhkZ1ffo54QFVbGH/lM96NikclugNpd
0WFCGfVjSAp6UTSr8hJI4slz99aUzqRuBo7W+349M+YIwGq9/Q0zp4IEhdq/QOun9m/jrGpGjLkg
/m1YIH/KXAU35NWM4H1gIVFszV2mUJcMz6+65+ejUXVqkOCVsVvsJTA21GQ2gb4aXxRRvcj/A1Ks
7T/YDS6QiEqblusAn7Ym3VWlIGPLe0LbMgV4i4Ajvyrmu9Uqu7FpJlUwlLE82dcL5XFnok+Z/IEo
GiGuDWPuTzhEiEWXJ7fHqbqyhwz6OafkmhsYqCkP8pr6BhPzqCLA81sIl0Br1w4l9DFQD6heGfgs
0oBGs4d4dySH0QJskAp5G1E6srmtDM4rcTIM78VneJjvbcfOHfyK5un1Ad6x7QBO900sQenpnbdf
KAMZ8YLUaE1Rf/ewvhSNbgFpmIGGPcmUe96gduLAwIAMw1FvuI6z6AqgKs+fOv2RuZ+nu4MPcXIx
uk591Jb8mzYVLGggbZaTb+BkjFMAuxfCHk84n9cgtA94cQRhT9wtFlSZG5NafPaPmDz8rEvHu3PH
jYQzdjLgaacbI7WBzQTV3YQcKyQyOrL0wNy3BBNXelS0czZpmjpUptz+x44pZ+VekNtc2ZFM3txC
kWk/WWlALPQijCOnIbP873wguc12UlRzR1yxfDbg/QZi6kgiOeqGTarlX2nz6q66W+a2Hw6ruxA/
/ZdHNAfjdKPs8hiyhk4PpAhRf1G37hN5u0paL4+bJdgv4eql4Uz/C+71zIZPO3DGdD/jTmI64dgw
ZG+Um274xaglOr8tuVj9G1xaMj9ASuLdFsn1hSxYoJaRKmLtjCnNp4hi7sv72b71immdFCkzRTid
XfTiTXNWNnaWYLGPkX8SP9tZb38GQ7GPSsWarx6aWmPBGDVMxXE5ngdTUD75JAwj6TNhwWFcFbhS
3EiaVmkNz0jseB/JNV5sC2z/Nd+G4k5jSvQ2jXNvc3TPUd8xEFk9ggNY5beBiFGgyk91xb5c5dBX
OaqpnjyiqOghoZVze6nVILs/tsJVyd6hLBUKTtfDcfIMV+NW3bXvn8Nd62oLW9doGaem5KQATOmX
WeXceDhzew0v6IVb+M97o2zuOGg1a3Ncx+BuM4n9RltJRQyStaKm3r7NSRU1gLP8S8mmVbuJ4Nsv
ZjhwzZPBnM/PVRVcQFQQWNKOnsfFo527mKRt8KaNf+F6eiFrJ59lc0nlV6XfkwKWU/zRpE5v7Q8e
UkCnJFyz3ZvUFWRgpXXXDERMcApsMRXDH3LP71b3D678dRkRTdJgyAMlOCAICK46RgJL7maua/B4
EihSVuHV4FJC0cRoVykWoLTswpOiVZHp/IUAGIoo1Oxg12JQr5+LrmmOTXIE+3s93soyvydiflqR
v+N6p8t7m78kfX2PREi6AlGa07ubamthFqQ1D9iDQzcihDYzXLLaY90XadiHmAzvMZfS8o/O1bmq
wPgmb4Eq1pDkNNzLid7I+Vf/KylwtCA8UbdkXyfx9TR9Aj7jie8jhQwGvbB4ncbbDQI3p8m74qGT
0/ocmxMNRiutDZPkavoe5lnX4Z63DVubKh0QOhaQcugeH/642SBNKMf7rsOaJrad8Vb1ZEoMZ+H/
DVHSRpDw2UqfY6ebjufCXgSISD3L7FvNPhm2OfHSDtd6t9cTXJ44QMeg9BvSUTjKDQlXHLTzmD4y
XHjhKE6nonrrf1im3CCve7SwwOfretvtOmXGqKEv0uRlyWZ384gURyY43UtwFh04jRecViek3ep3
luEwmGQ5AttmQXwjdmRIVxKutZV9kX1Tl37YWGMgDRrNzY/3uQdRlYEiwXW/hop6lVkXChUUYXrJ
e/+KBOmLwPUokr31omvVuc4NHj8ZZoSqxe1J4bhNmJMtVmbMp2F8+yO9SjxNRFd8N/4DFSObWo+n
9rTcXWv8n2DY5HuN00LZprMKCtETL+9WPjeO68/xAQmZAyp7ceR5B4ZRQKOphwoQAekrsQ3h1TyX
/GH8lJGdPtNtzwTcMTdGqP5giGMxLnWo2/kq3FGFF5Iwl44LQjspZc6F5yqJyUwtwy17xIcOZwTl
nhUAEla1Lv3IUwoLx48ivhFPyniWFWKyfMTk6d3fbom0E7TZGfwv1bUCG6YGU3Y96d7UJkojpd69
+2uogBQyGYJdKiAUUIswkPtXjpR2qWZVUrP8fzuE7bDrzmcGE0ZM5Re368tf7zTD+vv2AApi+l/I
qyn+/FrpZAvHF5sE6uu5l4XaoxkhhOKfBPTIWp7dSHZUo4226xIeZXWmOmj8oVt92eGcRz3iIBs/
OWO7em4INqtE3tBfkMp4c4jsAc/GZSauTEveC4KPQwCr21HOazZi64pLwMRS+8QPzlTz2xhbD+U4
I1/Srae4nf/kY36bGWXA3gFnFMCSR+7Gtd/znenBmrfIXIKwpsOxUBFORIUTGXz7h8PuJFuNJpeu
YBEN67ShPpF7ryNeyxZRII9pjMM73zHykfNprnPPaZ2KfWiSjOV+IR4b6v2+k4isEiR93Cu2UE4M
sy5gjYnRW531U0y5mHiiV1hfV/t66qvTLEX3lT6DSiqNkxgAIbhPq4kP3EVipgyJb2xYzFHeyYUI
oDr0JNE1VWjQ+v+4iW7wq8xkbtdoxD/OH0l/ihTyld9zvxieliU9DmLFfXblB7aW0javmAn6u68K
jEoyjLzbdsg80ll56RhSb7+4TqmMa6k2FUbALrj4k24VTod6Uvmnx5tHEX8TnsaKfoAJ6Hfh/NQA
IztFzYvmMnxXuDY4XJ/6WBb1lLGmNKOmTmRU762m5OCUtYxfcAy9S6FvCQEpXz0Sx6g/BiZZ0JUk
QOeOeYIKa6nU4hYGFCc+r9glAlT33NmiGSAtcc8ZzWlQ4WeVbl8DGlFhXw5aeF3WnsJKZ5yD5Q6g
n7gxEv74HY0Z+LdZ8TmEe6g65DuBoj4hpRfq30KWWp22ECBDqk+n8eWhnXCqbj5HUEwuy7tDvE23
GavllBL34P4VbKCELF5AlVQmoL1CSXeENN9/qB7MndcHxhTZuXv2uZ+RTCo/DLSuaO9u/ZcdCvA1
fiPb8jF2ZalDCs+xTRPELTACMRz3/Zv7atNvfVonAob2pBi98lHLdIy2o5Odr75w/JUMCkZVa6F/
Dvl+oNWhPndyp5CuKE1AYiOJdGm1YJyLDyDAqdDYhZswWqTQQ6aR7RTPgRnkaRfxKJogj8RPuDzk
kCPYu5LBcbEkMAHD5qlMSwxgcDlFYJtixtK/uNYbhTPjND2pSVY8o3Z8IjYx+n4eSAxxOnQ5bg21
HMoJJqJ89sSk2EH2/fe4rvADIA2mGQD49+w3MWTbjq044OMQjo2r5ULCeIrsA+08r6507x8pkIgr
D+tfNNmNiIBuLB1gwRZMMVxtU5iYkvRyd2pcINB2RcwJ/RGeqJ3Wzpy/gc4YopA8iqCYzZmPmUUO
EnzByx4BQQHZxIpv3YRWJQ+wdKqczeqP0dC8dRTst5r44dwAPDRmCHiiD5GRQIRBNiKqRZQuPLfP
gdEbzU7dhQVdI8DU0DRpGsdgBCdTnrj1bMPC8W48gPb5mD/Vh/5CDpL32tWS2dGGgNtPI31rCEZk
VBAYyx4gifJLf952ZvmYVG/trRWFU8T+HQdBmfbCTuvSGRKVaT2pdLte10T84VL5DAn53v/P7k+m
QucAZejwajDJYCMOsgnoQn5E9+D3UxOPtTpRNh3a/XJz00Y/Cd+RJiwJKlx3PwnfVPxpk2M6Ajfo
JFpgda2tDVAOuyJY6SDxMs9rh6TurUIq3Efnt1BQUqd5GE6GC9fF3riuWrymGVY/PVcRR+csaHhK
38rQ0Ay1594YiEZCmFtI2/YHiNwXOEPjrXjc+e+SEEy3peG6d4sH3o2bmeFMxdXJKObRaNllOfEk
ZY9rQhAVRb4ybTNX1KyEDJyeo/4NB4dsobHhwfsUnAB6PWpe1TSOmZl7zA1CwvQkKqEevOa0eL+9
RLQCnLOYc2BJf+IAjbp0TganR47CrR9Lc004URGmmK4yxzoTUHBbrG/KP2aU+ALMeO7koQKuc1J8
BARHCqa0eMoOXOJ+M2FB9xITXg0X+I2NCcCGU0Rhl482UXeSuOqOUdOEzGLtoY4gUxFHs1m62oEf
nVYG/Xce92MD3JZx/zwNxJRPnuRYy1ym0K5asWHDNZoiPxe2tRh84tT+SmlK55P+Z7VuyNDQ1lvB
eglhY/6LEndtwuPxXqy8M3/M/Gs5yXJjPk86LgIxwEjF/oW4l+9aJWcvao/zpN2N/vwysP8WPicz
SSVnEnDEpbbjsQYY65nSdJP8ql07ydwJRCVWFh2X/9Ug6Sosxh+nHfgmWUkeIv9PDU0hxg5nIKce
0BLsPWdvC3rX+26QLd6OL7AcGtX6pQcwBc7noLC86YJiW+tQI3IKPTz1bn069qElkz6lZX9TCbSm
Ej2LrZK/D5vAH5v7dne2oRIyQgS20ZIsa86U1ttN+E74LgrpD61NawYiyw5sveBgFGA8Eg3mtAJE
I6rbKiI8TntrJN5ime69fQ7LaVOS8qlUQyjqVV3JyD1lQvuV6ffcUoPywXa/0L9QAXEf8ynQuBLM
3E2GzxM/dcJqAWRPPs5JvVqeGTUHfqYE0TJ//pjlu/jAAOTzedoih/MN3sWqNU1xXu0wypMdBV0q
+u5N0hScOHDvU0p7VD7g27D7PcjZTfnywcWcnDnFvuMd7UFxP6RE0tIlWsZC4CU007zaVMXvDWMU
gxfSdWeLlguT4/Bi/4c4DNumkaFuBazVrCTg5S18mT4H49peL9OyBcJq6oMtv66r6q8jZeGwaiG8
Gs7yt5XIXHv+b8UFzXMoeU1Pz81PqN5FQmIrlVvujlQ0LB+T5WB5tLkLfTXgNjHEKyMkQlRBG/cY
1xHCyJNow6AoeS5oUNKFQNM4v2Mw92RIMlpBknhOQpfa6eZtGygHrkjfTHGaJxoMoUxBdXS6E72M
WKpU4pmekJc+5J6CcAI+yXK8iCdbPJJ1ywACq6/OnSZd2Khv4Xtz/EdhdlgfTPp1vHCfhgetdKCj
lwVIf75eHoCLlclwly2iRjkKdIKg7MWMZ/7VdpZBO2XzbiWu4ACNiCEfszF4hO2PMSrB0EN18nw/
cDX9rjPNzO8ROkeX76ocfvsvbIMe28M0bXA7MjxWjKYZ11Sdm06WXS7hG4MHMEmOCLM8TgfJHApL
HdF9HcG5A76H26mac2RJySs5RePdmSx5aJWRdvyScMWkmIHf23EXkYJJJvrOjcg1IChhK4vrjiz8
Iq+/YAw0MbXmFYkShy+lw4x0qseO3AXdiTJcufzO8CTylcRLo9HMcD3627umMSkg7rvfgjONi2gt
JW1VZcf3786u2g9e+xoemeoGbJyazubVmcwNsRyURKuXpVI3EKjL4THseSFd26o9zrjFWLBV8bFS
IH+eCey7RNgYdoRz0ne3d6a/obNtpuDkAkc5lAj5tKEuWnwrpZVRmcx9hM5620qSqTh/MTVlD/ST
PZO3erqSgvFnkdIMsABzmYlom5777OGRvVB5DUf7uoN5g4IeO9wuyL8UDMCZwEnYdYWSmLCRr8Ej
B5dXEPZQAU192U8q0pvH6CCvnRC8U82PHTcAjEkzWhmtfUtd+o2f1S4fYi6rIv3LW/AtR9RoEtFE
v8MeyeY0jWDgOeHcP7GtUqyqYKN2XaLl0JZse3F3d3kYSrrbwp0qoB4GmrkILYOvlro39K8+BWqG
rm48nzSUtI1Is3Utgeff9mETdfd3y/oy44ZpsfaNtjloc0ifU31AUkFQ1n+sa1jOEL5E+EVB5XGH
LOUZmjzJhuRAL1eS9tfNg2vsw+WAWDAR6ZfkbqxvFONk5g6BEor2q/f9ZmGNKxmn462jjOwxVJQE
fO5QiEvTQQN9ovcAFd6/IvjmipRGCeL0qYuVfhbuDOrV0FviBhrnwEyUWtV6LwG9wQgepddxI3Qk
zuxCNH/w2cOI7zbaT3Dc4IHUDRGcG2OZ1lfavYQ1fJSjGzn29DUGauqBzhbYlju1uYWjmIhsKz3W
1Yul0HOL+wQPBdsLxpIKXhm+R1wnKZsozYSBwNrI6HnPwIM61S9/tGJk/cC1JTedWFMjrpvWO9OR
NYV4lYrYLrck93ZZsoBF633Kg24DuLJ3s3KQs8tvGo/QPgGcSsXPTmwqkJFAP1YhSLOYhCMFR7Va
lOqVjpB3ezJ6UkaHLTNItZjSmjcVmwkZ2rTrvN65Llx0gPKKpWT2p1k358BqkIEWX3Fu6bhbdE+B
K7eTYiZ6qaMyIWubD7b9Z7hTtBijmGxX4Lcxcpmsgk/9jkX0dVrdrLrzYYMYnbelmfrjAj2rMl6i
HowScNccqwYIjOhft177jc9mHWz1s0vxJiucSVQFl1riJmxZODDX+aZsM2m8OGImbqcy6mdtUgwG
oqwHxI0GAitAxKVSoMffwAtm4lbDDzSiy9ABSIL0blgRR8J8V8KvVBCtCdNrDFxb4JNECQm8lECl
EmRnMIk3TVkw8owtnkv+fx6OA7pvYK+6KkZyrP1WF2ZrJpDkbjNEOPnWCuDIya5/eywDLyjst3bK
JTvsUBQ5YvtDKOzsNqwORagRjaaNWqcqTYKd89T2kD22D1Blux0hVx/cPRG+ByzI5G9s+9urGJYr
iJaibLLyZfTcG1/n8jwVu3fTjWroACR/W3ImHVdoOP3m0F3fHW3CyQThg/TrZFAqnNDyz/cdSf1s
jXPzXYhpXwH4bHKwXvsfYqzgAdgTRIwG6RXLjxgO3s1urI5MSPLHs7WfBHwJ/30uiH1EaWgaAPFl
8tcRoUlb6z/A9bYbyVs6POYlzG04Fu8b4rjODsH3Eq//SZzMzhN4bDM1r143pRbgUlpMWZmzINSV
Gd/lUcZGLuTCCiJC7f4+1T05UyaO47DdD+N0cd9SLyNrGMJ4aS+9inDstjCKBGsCRrTGe5iFFqGb
uHR2HEE3m56jVP5sJWQhpM22J5MCNS2WxrSYbJc4dgURxsHNn3mkZR+8xTvijuvBpA1dlxO2C5/+
+OHsLME5Oame7k6TCFJ/OUQwwgOvxrCw5FAWMhV2QFoLxOMqB59F5GQJ+JRieRjio3gy4hW1wN06
zDYEf+0nqJj0qWYbSnFjYx7oR7Nkfv+QSPXZ41nLqq5rOstxcs3Lc2teQ5OMX0auIYI+4ByDDSjS
PQVWeIEIsw7yEjYgn7E9X4EM9MwErUHgNdfzwFCF0oZLn7EXOAIvFaR5ge9W7ziK1LNRAW2mHr2s
/0k8KWIbFcZt6o4JskI49i19QAg+w5op4LfPkYR9ezV8oieJUH5PPQEIlayHahwqiCWnOoDRLxRC
9Lqis1JxNbFNchrstBZ28EqKLLDhAE7Y4e1H38KvUzKKeUkDxPm3peknY+IFm8JxI362H6IT67bz
6DzLNMVT/HMja9baQ9PVlqPL6+uknCbTHXuqS7jTAKBVHuTCsfmwtuZ7TrIh5SlxDtOQoX/NFTdA
5ehU6GOdeNfo2x05pqMz9ctWH6wOkNozSz1E+11TbCUcfgrLwQBg0hb5FjcZCSpBuAoSnibP9WvI
Y3gImBwXbZkC1L+WCqb/9Z32AG2r/mMY1p5ztY7a3kFNX4Dc1D93WjxjRDu/pGEYy8MPPT091gSF
cYRyR2OX4z+vxpAVBlz6HhjryEYJ8O/+VuUAg8Zv9V0Or6bG4MLBDFJ2RjIXiAmuHfX5LI8VzAG+
urEINq3KjxR355msng68vbmUAFV+JffQVLTrMYtusOH9U2k2D2UXqkk/s1zLG54P9aH+nk9i2y8s
GPiTDMJBYDbxFZC5QYwnSpfweNc2aBXl4viu7PY2Ue78k0IdX30kkl3a8OoZAaNZec6KU5NE7NN2
UmqOBton6jaaY1oIXhxfKA5U3PVPnanfI5hOaU1fPzEInKapB+edyCdeqcUrv4xguXhwOdXJZFcx
HMIktbaz2IUMZ2MzCpQfSZgE8R41vY1o1SGYuyMspn+FJpb1Lmb5l6jiBKUYt1qTdSslMq6GRS1f
dzGDPocJ5DfM3odDDuB/rP3Pfz5epFzgRalhbf6n3Bpp8R+Bre0hCHdU9ACspxuVc0XgqS/KogHZ
0h/dwYTnwB/jRe/qVQfYA8m0/ykEGDqx1Uoom2HpCJSCtV54YM6hFRKAP9sCREUvTFNmYbSFbe6X
rQJfJjS35pPbbLH4cH7qixWAwwmTJ0S3HZhLEQlhNTDRmX7evJAqrl2zCigqD2Nym+yBRRcsWyej
Pl/7kRfwzlxyJS8HxQSIQup6DelFc55WjTzZnJI0Y1qoP0ztpfEIaIqT69A/dQwKAgRphet0xwDz
rTxRCIzTfmGlSrUuL98SzEqEPbik75k6UD5mJyjKZm+iGguoW6aqnSBULfurlvMOCk24yMvMZQkN
macXJTLNP4S8jKutkaGUVeLPk5waYz3i6/Gs0lDY6lvCj3WOhC7XlogGzCQOvYatIS4ncJC/inJR
sEwQDaXz0v/rSgFcdj7/c/s2+TsOQFVNt1uKhaPkNoVTZ6mZ4erQ0d3sLSKEtG9iCwiF9HviMc/b
rFviOS8H9B4HvslEKSi9JU1+8PKVInxgN9GmKnPvfiyG+BlCIFfT7GvLReHaVIBO0rLqHauIUzb/
F0lkGNtdrZvx45JH7Q4VbDhHV8vkNzBbEQALiGU8uF3KwILQb8J/N/tHd9SN8LQMZ8BZaYSmmYP8
g1ANeoTvnHfe8ItsYcyeSQZby4oU+hmJ0qnlbcG1HEcUiaNEDN19BedBYcUu+aXGWifuoOdA//mk
sjFuDKh+paMvrJc6joG4AaTFPIS/gVJgkrwP1YoJvdCYCx5mjOXiimXKGrH3HupIWt+pbPiFl2Qu
B3gYG/suBEHgUDlbcYffXsVmcvU3z5zQgx4W++kWDrgProgFM6hOwndlBuDBR52Fp4eFcxROJ28j
kK+cSV4PcFPpOsLPfZHbLIwDSzMaVZZPPZHBtvu22bYh3shUKKDQaZVkTjTKauQ7m1f0xl/4xGra
qO5PA4Xo9iwkCir6U5eg+L2GUHcDPHPe06fJ9CE89SXbVGYnQfRvff89drhMYv6xHE4hr4LzNike
dDyoETq49eVO52y63FuwRp2bEXjKvthyEXi5Mesit2KF78fyPkd/D9a7FJ50gkiTnq8DFNqLvB48
QxFxrSJ4ZfeVt54pVtGlOzbIe6YKqN/nmLL6tAKZ4pawX3LRt4HTumoxCbB4Q+fKGpYnQsA/UJ5x
9MkzlKNMctc6jLDyjyywlJ3hjUhLxvqfTYVLP89Km7hEFphZzwBvAYwGmBWRA+qdikIw21BfkzdW
sSMad6kx9xM9Z5HmNAVN20WR3kNJI59Cjl9D3Wk+8akKZTikomqXt8N97k+XxGdM7sRXbS6YfNVG
fCt16kKwxA9Oektbb3qnOqQrPxU0HVdvJT5r07RX972VpJ9Z/mU3YD9svnJ692VWNF2tauU9C6ws
cBCONTo9i7tCohUrSAaeB8wH8g5uDqmjrSabriEgPT8a0kTe4hjQlI3QYRAUfd8dsufGTzCd3YIP
InbwfA4pepPN7vd6HJFRcLySCMoZeDsMTc+FpHm3OpT0GAPudkSO5v44YMUP0tmU98U0wPLg84/p
vIST7OrHu5UibKWH0Cz6rUEdPxfyd9k1B4mZV3yxy8TR2flr5qX4ky/2XNWW4S+Cyrm/FHyLl4y6
3ANgz3JwcVDQLGA2ju1HdYQvt03xA158gKLCCQ0BWrnPKIWi8xQzXX29yWtGFE8qWLHaS8t9r7wC
Wi+NHvhRYU05oVyADqDae0vvP+JFXkonstGL2fA77AB+iOgskGp9SI9fgzCgR0+6fHuGOX+mzbNJ
J2MFFiVQFuk8L/6mvU4ICmGLAqSBhz+Aq8iDEoZSR54ClODbLUC67DZxlzKN6BDs0ZzFATFr2kbn
PSo3ZvejyEerLm0C7hEgF68wUM1u8uawbND8Q4YuGkobIPzO1VYIW73/MfSAi396X5QAhuWb6n6G
UGfn6oqrUVI6o/gnN/fQ3rUCQbMeXKA77rIxbjo7XOKrpxtqf67kFskN7FCgPLMJ6BWtb35qyhvo
JU7laV3z6i6CZKLZMJ5jvTwVZi1Z9b3mUTIXtKP2T1m1tMQN4zutH4zL+jUVoscVy2tEK5VPra13
R7hJLms77b8COWoeDtZhh9w6qX9qM6DIgkdB6P+bbUSh6NotGh/J7ihVJnINtqmLzJSYF6oRUXjA
pLd3jrzc9WZ6bFtFxLjLvLYSG+VaqKONxDBmULVsX+UrKbUrj5k8tsw4PR00Z5mVfwSfHDaoYhSg
tt4GJpCLpJ+YffN11DOYV38GhaSU7SLJWIpd8HcLy6XL184sJ7uMz5hhN/Ku4rsi2Nnqb+MFazRr
jwDReE2nuEvExdIwGSEncfOa0p9w8PassgYKDB5tLaxJfj96L1LIsiAw6I9DeEtFqOLroLOrIPfm
hPTnStmigQLeQF3TQm32LTMzyqgk+Ytp1LGZr1go2knlnVcRm/ZmMGB82WqUnE1jtjmkF+z9oPU7
kvwbZdjJFU2/wpRlxOdmkTlCSPu0RQbX3J0y+PLQPEo6NPVLdYspCpX5ie3AkrhlFGCx6gS4emCU
QBEZevwj/KSlQb7EX1v3xii/9nvpvAGHf/vQW5lerG44fGdI3Bgu8AEoQv0f5GSkVX+n/8pP0qey
eKbS+Tq8Vr0KuRnVvk2k2/Rq9m1dtPb0lS3k0BSPkSMnAwOMAhX4NKmV54HCBdkvu+BU/UJCy51X
3VNt8PECQoSiUr3yVPXZSYjVBRtbuMwUClTHvai552/tOeemH9d6vCpPaCfWnJjIap2Bb0UlZPtg
uQBdusZM9jneigKjk5YA0StB3HA+enr6ad69czERxI3wV0+WS2EIIyhO/Vqqyip9G9vsayfzTL2o
7PwatoT3tHPfh2y3Vq6M/GfjXXTPN9uy0LMdfm34foWpa5HQgb/0nF1F9ugeafMnoHR+HkFPZSoP
jvDowaBC2yFk5fU/Cg2xVvxgxmsleOthH++4sTmpHZXsuvlV8bD5KlXhB+BZcFauQjEAqC3lru4e
nFmw7hAOkpquoqZ1bN//8RErkGFxoSxdzGilOCKEbl+7Y0HwrjGmKEQD/BevyDUKJGmDqMnzPQhI
RZBKT4fUZ1oe3P8lwqMBWkJtB3ZS6eRQcJNaLV6XM2Mdrv2LMvvUApxS2xs4jrvS7fK2LcgbDrZW
j3AjAR6PIVcB6mlzsfp8wOuP87ar+ZR6IC5drdEk/p/z+rXKlxtvrDZ2DuN7hVt16uHHykTRoBmJ
JoWOD2j3SFM6YHfZxPbtceWymVX7oNQx7y7drgHzipcXGds8g3joTiE6uwvYpi7y7DP3uAMVZuQq
Fus5WLQdDQfKr2/Vn9L0/pK3p/txxvIs3HWexESPQdmxKi9dcbUGVN18hk68vCdEBnnBor/2AIkK
Y2KgIqLFHphQQ8bE3OeOJzGC/ttBNiy+kbdwXrkPjq0glGRIYo/iCPGOvhtj3fmZ+X0WhTZfe8cK
4C4ilgupnIwmf5R6X0O9BP57pVt5lFb/DB6dyBlg7U0XpjAlIw2nU6p/mG7qbFVxbUPtc9L9jViP
kEs5szwsus8cDFVfBqVm1Sk2/XhAaaQWr0oYzlLbP6Y9uTvRNy4o+RX9hyX5MHO0oyey5swZ9NyY
aDWD7olUPvjRpzS03POtLV0/IPoLE5Ip/afhpl1uVCUYEaOLPmT3hBrWN5Auq0vFuRI1IkrVeEIG
fgdQo4CJjvnSO/nLOAq5kKau23HZXmU3guFlWzjvUTdMBj4O9nq3Mm800h7W19gPe7V0dMCFnD+g
cE4PsY7IZLbZTPYNjlvsyjcxNWbIjGkSpbY/7rpmjFiUpRDWChDfEKbCMkPcayReSfLDrGZsOHqN
XccjwOYp3m9e2LEhUvlOpiKfx3BvnACgT1RAA/V+5LccTccjpT/qL3fzwqAnw66E+x1aiK9JlgpS
mrtyz+FgcBRKYhcZPNvFGt9MzpfksE8OrcOAFI7Ej8WwElF2v9DDrh1jZ6gwO8hGi5/h2f4fhBBp
A+hvskcCJat9h/l+iD3cU6H4auLC9Hks8EcJI5UZpIylCdpFaEB0oNn6NmBqs6pDrjIQGEMg54EP
9RYroymQVJDbPO7o7D2YagtR0Zddud/+X1gOFSdSIsFfd10FMcC5Ye9Nh5I665/W5yhfNYQ3c9X/
dTHpQ8LtR481tBMdvWZoe0FTG8gcv28NyK1lhRXnuca4p2D3u1C8zK3oG3mUs0icieKFvtV4YbdO
mFJN2gyIXyn8vumsHM6/WPr8KPyZTSsyDbL5/6Qq8QgauSSKHIzf+oy3BS59875rZ0faoPEpzWsq
avuBRz38NIvVoDaiimWgipNGqu9U3X74npJgmk7dqfebSWYLJXHs6wzeEmHpevdh2Z9uBaxCPOfl
xWofxyLvuGqafefIinCnCmCgE07CyRHfTNiREh/CBPq5DjVvs2rLKEgVLUMuTojVmjLNb3BJ4ZOY
LNzr45Y21posSVU9B6v4C+mhqIKpQT5/V/otv2i5DHkLyMV8Ma1q7ACoLiJgU4NrttAJBNdYasW6
Fdidx5N2ltYpk1/Rx4ZZem0j7aYxfwbjBi4odBrZb7aa/T1uib0mqzKFMY515UToCwBNXRZaxbQA
MB62NwPDoV5XnmDvMUavJRC5nX0qjln0x4LUnOkwwI4++DnYx6LvXE/Hrt0EmjgPTgM6YibIfYzU
bt5Rd1xJhUFKboQwPVDkwedb8QR4BzyNYdKVVhYW2L3EIPSGK4PEmofkkbxOI7mnrv4jfUHvupb9
yxHDrdyUhHh0+mgiYhmUJkhUF3El40SQVt135//S1aCS9yQCbD0ntnx2hSGpyFtGf1MY7BNXuoCq
TOnMXgiOV6HMgBDpHpZy5VjLxV3cYYGUZ1ZuEjB43+uEDC01Ljr4A0Ne1mMNKm8rSssdjLdkLUvv
+9MjwIe+nSFAeay15Ulvq8OpSJpX29pJkLZ6NK8wbOBFEmT0U3/d53lVmiyHq03P22Q8X7NvbpLV
35d2t3fDQy0R06ZwtZpPlpPGqWM4yFKcFOGEgpKEyHg1LBlKsH58T/5uI+2eDMMzxDoNV6Dz07hp
OSPkN42UyK+AXEBbzc3g1Ub8Id4Yw+KOKkIXk9/J5nkgZ+KlbDjZBF9VAX3d8DJUJIqf2hWvPpYP
Y4IBHARG+Z0yzTCcq3qVQ9LcQZmVnsotajIGEW6XtV/9YxiJtHhUHwGekmRP0+lNmH+b1ugiVKtK
twmS8q45A4I+rYXS/ENvpXJtoFTp1H4XdVFPIht6LbqqwU7Zd8b+ZcBpnE6q7uvQbqTGvDrU+Ogp
itxU6mY8Mss/hETBsLI5UAAub/nZOjjfBu481q4Dp42JERwyE2zHGx5KX89gngN+Wl9FShD7jKGw
uQEh8lov4Vg0XK23j9NeZxr6NsR5+3e4H2GmSnP0xyvBmLfVl58vLYIzHiDJZ7O066G+DuUxsIWZ
GDnYYTzKundVtwxX9lN0obwu2OWzKIQGYOqUBoZUPlnHsgVpK0VU4lkUqK2R5rcVKYlf+wiI121m
1xcKN20ZodBAfuad7l6ERliTfTC89KBFsFKjtSmp4k0h0sQsv+Nb2eOSxri0UEwz+7THAl9MRg1C
E64q/F0pV3Gc4PGPA+QYQV84kH7Dask2MIctBuamnYiIeP0KSsbZcHlSWX5AOdVJWKaZ5iwpEVIV
dfTDj5O+WbwBEoBbIcIPAtshA7gVTR3f76JaiEQOavOD+CayFJy62IALuFhDm1CK+LFpd5Adb1Q/
gLCqTjF3dBA6LpXXlVA5DBZWbxFcLyCFZzAQtxnCNSQfT/SLYAXPSqztxX49eEiLgvisLS6sVbMh
RbT/5xj5E6uA7iCx97VfpALKhj2nDG8y27jxXxIOAPGkWqdGIrIx2GAMu+ArUQO0ALMgmHr8+7Rz
B9kpegS4h7DIhEltsKaA4rAf7Sfvd6VPooVTw0izqqgzF0gYgP0+l3haHyWKWXwFD2+hWS0S0WmT
zTrp6Lkf45Zbb7RQvGAanHtHZRkQNL4KOb0uAQrQheMF4NBh4Lbvx0eBR2K3a+hy8Wds2YR+RTUN
/GiMXv+Uv3zR2UR75AzBQT/owPvwA8mqCQ+hxnuwqqad/PO9d/gbLHTq9BDUX0/ok04Vb0bS4hV+
kC2o8CfFvM+P1+Bbn+XqrRv9cDJela2xm2dHES78slllqaNB6o22cezdeBKc0hGA7/qU1S9qywOl
W54ppwr2F2bCGo/b5ckZXS/Xa0zFVwKHEvK4/WBftwSJIp8Uft0ZbmaRwIsYfir7a4ttgwPpdRPW
2WMeIA1DmZeeVBB0ITEfLmvgPvjAfzokLejK9/9fCoJ2PBQlcUfoy/IP2u26QnlPaZxgNdhNrLDD
EtvaUTpt36XCY9No0ImobLtgl0KpbhsUlHTCSmKC/4NJjyuWIm1fKYpb1xj/y4nP8srNDWEB3E2v
nffRKkC4ZSP2cSNQodlO0RWZUjYBLsR2CeaaphWuXT1fFEBmJmlSWl3/ZoIbvRLQeRzyv4SOoAOq
NUTCO+akbCigDjhDokZ8mXDPGg22nkrycnq0Hia+2Xj+mQAR/wW4XlBnSdwS9Bff6g7NBYnx/Bdz
k8BptRsMRO5m1LeHgzJsd9bX29Hmcg07cJHOcpdZXVxD9VVty+V+9M27HFDpEdpT20l+xbI1ue4Y
kqBufMf+TYtwpYup8gkSyk12qibeKmmj2dkqwc4FV/PcsottCTVCnCQN8MvrXqPp0x5xKGr37m3i
DknnFaMHHxanoIGdDbutIr4YOXxPMs0v5y6Jkmff+g0ofLhysUx8KHNfI+Strp1ksDgnOd6bdfLD
b+3xIRt4jzQlt482Q4FeXAyFA1ee04hbb8+N6oOHh9eBcJjONWDf9AQHqTNeV8qK7BoSZR3iFiUs
QPWrQNSbg4dUWwCGSmL6Ptq48kQv5TqxeSexlTs/A+nJ0czHU+cvHVUw/lGmK2gLd9M+RVQG/Uhc
IxnEIs3FR5pdq9lDA8Rvp2DiajAvF7Z6mHMToYuPvvNRRiSyinknfS5vQoplPqrtQgdR17bRY10u
x0vlnFxF/TUnB4h+ASpyHRHTY4jbvIty+FJxUxAF9jk7rG3m8HwN08SDXm1D0N82X3FOoHiGqLaQ
Nb/Ee8PjO9TxoUPUbSzyDbVkKlqOxAh0myArkhOD8xVyLS/wFqskxdh+EZelfoHjMTxc1UPb666r
Eb9NukzgBT6/3tqXtxyQ3g2frQJh5fFcW38jC8/T14byvMJzHcF/yyhzHPcET6Uxu09jqpgmXuAt
/twQFtisvVquYVF/pHmupHAYNP41k+se+YTRK4v7qof3A5v+FSM65k3pDKz3UHWR6BGVEHWJgsWJ
w/VqHuz3Xe98DfqymdJSvDKJCBqTYaFW4/c3hQ/UyVaTNHVJ75nedgh/r59r8OjWcro3jyyrZaQ2
JU1mlK4Uj0EtFcDXykyofaR2lC39+hiAcVFO3MgQTcX5lQ/cQxMLvKICUUJI55KU1PSuqFQ/tjlW
h1gS6UEvzD1t3r2XnHkOMtlPSfBDZIL0mVvI6MYk23E0SvUwZ6PMKNw4S7RAE5lYmEacVQ0Kp4aA
lgSPin2/Sdri8p9uDLksmsXmxxAHfMbDICUeWOQeuPe9jwLDtdjIlfcYxOSz/rN4a4WuRH83doEL
p5ch0LyjwmYMAYEw971Ja0wfBsTklu/KTV7RFQC9lBAOO2lJ3OEhbG2tRT44O/nBLNQ3O+L63upc
Ze/I5952fdX9zmMv1lAYK+7b83Gzc9dmT1eZ8DNl5h89fVjH/OXWxx7zyHm4NXMnlIR0lf5peYcw
SYS+s2nZP2dGbZ7KXqmEY93fC/BD7dPdkfUgUax24Ifm1AIH6UahXD4/4yY1gtnZvyQEecL+rWIJ
vnNSN0HJwpn15DP016JIgF1mLT/tscLru8451N9zbKWv4JHAgFJVy5ucnhDGIkRONK4e/6cAoN4O
pzNuyJJNfVdGeLAZLa+5JqXh6zhywS97lDt+BCidy/3PMqqjgaieTQLfpRF/5oRiR4q+1jjNpmCm
g0j4ylJ2uk6aLJwelkRoAGAR/lFJXjPBtDs1k8eEP4O+BuVR5fPdBL/Wky+uK8e9l40sTUq+zOPB
Uw1JjB6mCIdmKWV4E6bLA3KSHB4Bv3SnAxtmlOHqsKEkBPXj0Q2jidy574qa8s0tVDJpmjyySWUF
UDHq11egDEpEOLtvFp9DtZ/ADl4r3eTdMhKdBUoJtlIOfYxSpNpWG5fSge1Nj1dYLTZWP9otHUp0
yqtGbMkucRQ0IsYyBCGFpExt9s5BfnrGiOVeKxLVO2ia9EgM+nevsuu00VstIWljLu9sef731Vnf
y6fQn8nF7VUaejPZF7lBkaZN40xs0evRkZcNexZW4L4j4ijd6jX4XlON4kV1rXQLHYEY+G3lPT4j
Wk6pL0Df22gCPeP7Ta4nROGINXbISi+MVDLPuFMAm3rGBhjfQenTSVujoq2MkNYmc/PYHyZ5rpJN
9aSFVN6ZwX8VK+OJeid0NZMha5BgNjQvwG0glIyLEhijpaLfuoyeyAN252CKYfneaHnCaOQmgJVH
0rHgbIJ7/H+cX1xtdHRIAIKRn9WEtD2PrjSQB4Asw1nsQ97//MauBjc7oxyYRh/MYTI9nHD2j9LV
/nC5jfQx5ojYkzQN4QnxuwN+mf8z5anpxIx5P4kLdgmoqZVbGjZjziu8F/369YohD/VucZnIxgqp
lfONq/QEfcm9W00el2zXsHeWQGYE/b+ATroXAmk14qQe/puG23Lt3b5295NHjC2+SmGHdO9Bs7gW
S710+S7YAXy7ap776H1/MqIPO1vcMKKV6hBNKyudUIdIYk9cIRyKMkU1BDkMLVqgWlQJ8QeFkCTl
MeijaQubECDCOJ3dlJB+iFfyHgqtsP01ErUC4Z0h/OIj/0dOGxBg4SwzTlJkrWTmZ6IWGgsgJBPv
NqRrfcLVBYSJv0bEfbt+DH9ufiNCmWbyD8nLdqsyoMoInHwE0Fewsw/iCNSzPwQxJKJb+ordzjvt
bRMi2dfg9PQl5dnWg3CEALXzU9wpghqlpThQxqqAF+KTTl4YGMRf1hdI6zyJ/fsGROG1eFzr2mrp
seXKDAIpjNSruLLf7FiL04f5q6aycbSRk+avn5qrunuSe5uVBkZIDsCFr6C5e2o3ztq1j2/Hi1eo
/Z4o49MrvOMTxfLPAoVLarTMlr4Z9Tu5KItCM+Y+7/Ag4V8caiwjhwIv8Hfdd0vLWyTWkXXFsXTS
5r7W+tJ7ZY5OtZdxukssUiy/uGtQmSb/baNyRJuNN4DbmRmY54HVqX5SGcXZu9asCFOA+iELoGvj
BrbogFOrQ7V2FIgjjNeLJnUitVniUsdzqMU33l1WGJyx4x7hVMLJxrdDpzB5Dx63v8Vf7FUEDjoG
usjwZ4DpRl8+W8I+B8FPRmR1duyJEeSORH0ZodYNJ9stV9AVEsZcX7o6UMwi3z2nT4b3VnAM4t2u
BdYsiGu4a0lAUpgUYIgBulK0dNrsqcrkiHCKBdGoG4F5EwqyRzfdvhfR/QrmXdgomz3tlPdKY1z8
uq371Gbo0cy3UOYL8ilmtx8ISn+whEX8KOcXalQFeDs5xFmytljOsyKeKdOtXSwGcqfhBpxesgiF
BwiOC4vuFCjYb6z0JZMfmBLPtL20/njc0kjBV6/zY62Z8fHl5HIjMcZAr+YXUla/kosfoQ4/h3sH
FYhFlMEDXaD5XyCx2Q7X3umW0ymNOpelbh37AhnJ2sjo6uZ3zBEgSwka8YX8cA80xfwksHxnB1u8
Gq9y3hIB72xcXNKSYdEp2IMct+XmXXUsowCGNTbvJ58nT2qbKqmRtwC+g3jYbXPKSd+pu5bv6Tz5
dBKQv5rsZjvBhqk5xFt4FsN+sCmod8ASqR5l9mxcVzHHTXiytxt72CRrkgX2N0NLtF7+ePOzJRB6
Yy+5rtVO0eTct7F9m98F3KxPW+eSXzG4r/3hmcSV9uPZ6NOiqO82XjNbpGZOaqRalQwcvwzS2gdp
ODGYKPEvNnjB0WgXowQy7Fhzor+A38lQ9sS7t6mFA0YOnhY/3KoPzGQab7kjOtydua/HMqwu6KMw
UJaeec2dCqsRgHoCJAQEiWMncTyvU9s0+U/zt87xTrTSG/6BjZ9i1CjIjTcmpDWxt8yCvAKEQq7F
7eYApF+6+kGl98CXsks0VElaPOr+yDzjlTbnI1DKkzQDq2JUchuUOj0lDuRjGn1UH4vKUfxXAqsy
yNqIp1aime5aQ6uvOWZO+rttCNuBU/rKqLgtJggN1BeiSXKDIaRUpCHrc3UY2uauS5JcHwvPm5Wv
igXOuULInp96zcgtM/6M/qa6HmATfwGeb47E6TGTCEVRzGoJlbKoLlUIWahH00O8bsxIp0ytJi82
oUZXPx0FoMzq02AGWHBGzQfkhU6pxEzmgWBdvQKOgjMr2+3zyalDak+MK08M2FEKm0pp35oK9A7r
xKYUYJhnJZHax99Xtz7gxaaWWDMutHlvIVMxWoXBT7YJvQhpfrvR8LQ/dJoAxzqiiasF8BlRu+2+
OdZ01sUGs72pAEWUl2jrkgyYPlOsx9W66hOIvNudhDnEmzQ2hhCQOOXbIYGCM6rRO5bjeIVf7Ua8
TTnEssqzieCxGH6v7LEQg59shBvnXnUJdwlkWAZgrXYDElFc14VDMrIyU62NndQQBJ/L7qPX0zN8
apwI2gU+aRBGTOXZyBqi6tuGh36q4OkdHZPLzvU/ruROhul/jbEc8+oCRF1wJjZ320RtZSI+pdFC
Gb9onMseH4f1YFVdsw6m6/Bc8A7UZqCJCSkRcaCaOVyrNQiirHJ6iKcVokbyh3tyH2DotE+q6uio
AL7LfByYQ8WzslwrdpGkyyz4MX2mqlPhAVpzGxG/5TstrE9xiJyE9c62DGpmGGTQhIhWzc9jMPNU
T8qRaLPm8jqK07NcB9tBvlv1GUeCLzwAyDbH0BPV+f63o0cokCmtoyNwCYkAsspJkrT8JjBVfSwz
uR0s9g/ZH8+gaJX1DH/wM7U26RD3pIBpt4/xojKZT4mJ9p4XN5kq+9/mgpcmxK+bCEAejJcuLGSt
4dXf9vRBKUmXTWdhTZAmy7CpUTCTfJPpGE8ACtvh74aCts8VQvWysb6NplSmOS5Ibg9LchIVBgDA
8gPSoJhTmTvCcwgPtT7wW8/g37128IgCPIrh3HIaaRewOuIeM30e5w+QPmZPPINffU0ExYIZaf56
h7/K4GMSVE3vwIrtDT4o1AkrosIbkYJoc1L82dS9nzULG+b/sWTwhkXkOq1kqEOY+7tWCKxW+ZUZ
HfX6fGNKLMhz9reaZv2L7La8iXLkJqbaHttMaQe1DcKbvVcc1QfIkzMHxQw1lSseLycHtB2gxgZC
qG2Phh1gDu8UXU45WJbeZLBunbcZdNbBkXoQ8dKc0R2OVzy/HLP+AiCaWHQM62xLPXVPjH47Yp7E
X1RKJOB0VLiEt67fP1nM4uK2vmv62MFqfUTpGSrqNyMhvUlQ/IBtn5xB6BIH8wmRohLIu7jygwcj
eS72T94x/FM5AHkOT4N4HWhPI5ZJiODqwMY4lM/oOw8wyM2txzF25BuVkS/X+O2mXNhtqkyR0Vre
Y4yyCNB/IcOsJUX8WBapqgHm4k1aK8ClOUQHMsTyTaOeqI5YSkW7LbrBkxTiW3jJ8h77MW7laCCf
vPuYXpnhn8MufhpnaAJ5iHrBBSqfqRci0qlG+ETNdtCVZIAp6E2J76GsBVY8d07aMWz/C0/6QQcX
ToppUTjt2A5NE2kGrG/yOx7Fva6s9dZA5DktzgIvKmDf5EjxcbjBYqIxY9lr1rqkUUb1jJjH0TrR
Q6CKONp5X9P8/jxOB9F+CsU4CFK6fsocSsnVQ3EBNzlOeraX9Gq1Dnypi2ae7oQPsNI0tSSVfPAK
necY14QMaujtI5+Ua7/YHpkZ4+39NT9nJXL/Up2YKjS8sVzP6WP9W+1YmoC9Tm+YfvTLgP+9+2iS
SxrcXY8EyzvoB+hxSZHDRr/VxLt5scLJYOZI6xrjrUy6a+wv340RIKhy09i4THqMwgnPmV8TjVEB
pT3mSiAs/JftRhiNmqMPrZTpzJjYO1kA55F3N23IJ8ptxNBBUZbIord2H0ko+WrHBQKxcfY57c36
yUKy7hti92yTpkWYG3k3IHEr0LThCgn9CaCpVa/IzXKVoxSlnR/Y/ifHxR7pZsdPiX3RZdJm3Lph
eiYD6MB8S4Z9CGXYi/mq2QgO3GU9Kn/2jX/g0MZ7KnLNzqpC4VuAhfeTjZXBc+SJJpw2Kh8bHKwt
cd03C1TjH5ISB1alQGHFfYnAivHthkaCCVjWIK9mCHzFmuXWKBGqr+CVNGcrUtxyevZ7WiYKnZdl
XHrUtzsIxtZwPbuC0xTIQTs7I0hOfoFJwHaTT9ePrchMm2WUbfwLtEyPD73YCzJfhkIjBO10uY2B
DpkTrbZRGT1mnPKDHAjTiGQPzD/90HbZyUYmURCjIYTZl/LEsUupg2YD91vVTQK3aR6WheSZcEjW
VMCzaSRwzt4ktRySgqOMn5N9W8e4KuH1omlNCIdT2qOdgy21mmct2khY5OwdPCKzzcdroaEwmbFa
qYzbEpcP2myJN4soBw16UEWfwCyluJO31DyptcfC4fzDXagXflpqFFIEff6UnIdHvUUKk8Ak+jCd
u4Qpum8sGX1c3/v3JQZaBUI3wUljUTOcQ9PTm8arI7mdayJsc1OG1zkVuC+Rpy+9TLIIXBBDr+u2
6g/t/RbdQyHnISizrdosVPbRNoeb+aN7efax8MvGCO2cUa56Us51gQGCIfnHhEvD0DziZ+Ctwd2w
3qGxBaQoPM5OVOE9HIDx5aUGB9AM5ZgscYBOuhTUUPGWWUb849JyCPXgh5PWlETUGExpGz/z2qhs
etI67oElNB+MmIprgpLQEPffvEyP0EJ931vtmlZlcnJr6UfCCuFiZ+EFvSbkpNwhnVP1XAhEoEq8
6jZ9+bs/6KmvePeytT1INaUNSndWIepYDvtQaiZNsjIkP9/8GGTNMhAt1CevfU22dBtCiuYE1SdU
I4eHc39M3FLziuhkYpQEPga028cTPKxDXC12Wi9H/cJUMG2o94cptUfeoMoVCz9p1dPT1hewa3fy
ahOsyHeZT1EbSDbgwH0q6jsySqQ0LQ9rQInSxS0gEk/IWaEeKjHcxVqDhUTqBmOhnT/8O6j01sbo
nDd8ogmBCYs4p+aX0ii4nKtfmIDRyfQJMJlVALF79pXQUTigEHO7GanWnPTefe328LyvOclTnfOI
+iLZQ68tVwtjposWBsGXCDuXPxKbzq5bvL4ty1f5MCMDNwS6VvOXb4a1tN9U3wUqwNFp+j4E+6d5
iAGk3iCfCDmeQXegkAvRlELk9HH0fvQm6U1hIF2JLJPFPRBY85WjIgpJ7PnquBLxh7I7USEA8Qbd
hw/Hy+DufKM31QW9L0Gy6PvQ+R8yheWVmxTF074G7ZRFX28zmPnWD4beDPtNaTbn5xEhr3cCsNko
HAU7Uw59GRybvaX6cdv8K1gXFzXACC5y/2fIgmo17rL06aKUJ3x2jA1vqfqhpLWK2dskrK+RAMfD
jSNp/BJoGY/N8PC9YnrUwf9Cipy7iFvyjvBu4QHexhfgazmEgQQayn83hAAnI00mUXOsreT7r+Ca
VteNkNxl27LqUfRCeXhOQouCRsI42DU6v2vq8ZwtQ1cz14ec6EmJV107inTdufGdTZneGkwG075a
Nppt8kOU+2r1AJKHJNhPoPccgbOevhxSyMyMxPHFP1pRVgH3rrqYC3CiG+x5dqs1XXLHj5AQF/7e
CkhpK3pGrMrNBuV9YkCj7wA6DhAKpUMDlH63iriagODVJ0NBqmRTzu+od32N++F10pMMLVLJTmiB
NZjOazzVj9ydQsfZ9jSFIbFRh2PSy1YSoBa7syN7itNH3/e4GquaBuVGWpM+SUXHCkdtbo7OxhCK
5IIMgFyqIhMATinGaN2MuIDTcDEq2tNfYvAWMveoAQpX4sUEUE3mJyD1O0Sw1Buna3ZNX/zgHWdF
Dac6bSCcdysZH7WIqC2dGyzceBlafIz7KzwJxGd5kTXdkg+RnVfSXEfrLVsOHK4pvesl+DdSAnT+
ol/IgaN+PhO9Tdd5Sby8orvLTWm4u/WsQzx1dMCOHTXeAi8hSEYNh1sVMawcuJzyJO2eR+SaKq+s
B+e3n2TxClXUZ03IKLjiTd28tz8wx2f0oQ/5VrNoX4oVxDDyY5kWhJqNBVSpFdlXbuSMl949UVIk
vY35I8uHdohD7AKvBJ6AaDWalnjMtS6O5BBHO9mlrW836wWLxdPdHyfJMXf9nuHSQhPgDlkOJIy0
DfjUx7FVDmb/Trh/mv2UKwkPETW5dgXHFjo9sygMCA/DU6L42qaKb0h2gGXZFkrx/yn6Rm0EuX/n
tOhp1+wSrpF/bgzQimGq8z3HnieJyyY4nWS/is5rAh04TFITJGQt/v0qF8tEE4XhEhGnS04tP8KD
079gFjh8vSGQyTY44KPXp4cYVHMGXhzns3W/ULbRMlWZ6PVl9FnVW/eHRXjVpX10oUJiqTgpKsOs
zZ7SvxFAGHZgrMH/PB1jpagxONrdWG7j2oY/DumDqQPfXyuCUu0zc8uxZgjix8XEgQ77Eoc8F6G+
9OWnpImKjp9psL/I99aAXj3pzcSuH8tNdFSI3TFUdFr/5Mk/YbQRYd8WChdivHXP0g94147qgo3l
klqPUloeZGso5i0j9W5/J595Lh05jWlQ71y+ieesWPV2dXyH1ApsLo6ILzCEys6gbSGB5kqieHNr
exKQDKPPcBVBA8oBc6t1hYmtdknpNhYXbpCDxxO+XKMQHEQY59tJgZ5R+EYqxKB1L53ZoE0tbWqz
jsXoJg1eDetvtl8aVqOXQ/phoRtFlda7ZYPvwCSWBC/FqEJWByPHJ7M7FdZiQPpmCKHqu6MU2w/X
SFooL80iL7Mhn1Q+jeBhRPUSZuLwgXJJbQ//mX8P3Xxmu0/pUo2UjLJm1shmlsHXimUFS6XHykUv
dx0QORhpYRboA/AM1ZUs8zumy+9ZBD3dlhDFRl+7mY5tYcvyKLR9oHEyX6iyE8YavjwRws2Rod3n
YWRzMsrYqdb23P7Q8S7ob22sF5pIwlhd6VX+iGcXdbfG/eVGOJjweUxLxtjkRSEhfOkRVjMvzyQC
APfsDIyNq09c21jZTP7O6CqipPkMqfTc2yiGgUzKcTZLiBsFYF2w/KCEBfq/ZBYVpCd2tkY7ow8H
59JW0G5Le+3g30pTAIhZiQWC+VKUX+2E4e7DvQAbe7zUJsiF/gGqHyLrfpGfh4tdfAomIs3nGH6q
JkXQm8ofPpSuFXfVvGfzvMdz+H3P7OblDArU4ToDPmR/7UK6ByQfPvwpDe6MYQxc38+k9lFmHaIn
wcZIvxBC7iP+8Z7Gk0MIIiZkqM7L2VLjaOM+YjnU/dHqgCyBYqPLuum0tTWPVsemdecRzBMo1t14
vcEJ3RUZGYrkYqwF/RTIE5q6mPWwcNxGf+kI86ivZ61pg9vBDDfAr7KNwTsK71RfKixsQfAICDJx
Bt3GcoFWTk/SBhWQjZrapmEnxbejdGgwHutlhlzLxvfHk4MyqQpvaE+mzSNXPTdnX4c9Bw0gpBR5
vWc3NpPPhcgqADjbLo+qZJSZS3MYS6X1qqPHjx1OKzDW+j7TjcRec4OiFF2TvY2vEJShjAw39grJ
BHdSzVY88+zvtZ3qz0i4E1NOJk7OsJbUwEmZBBo2rDuQtjGv2AAwnqnOB4N0geG3L9amw+ZYnSnm
vdWuMg6/4A15Sb8Pb2JsP/USJOs57iainIcXWrGj2jwkjVBCLQqmNYYB1zs1OzzqYsDUnwTLaMBa
4ZumGgl+RY5hCP2UXkFjTyRWAlTSzU4kOulTjrBjviQcuVAfhsvreRjhPMjOGKNcJOQKNO8LmDOi
CjO77O43ZRX/LoTRFZwlr8nrMj6E1hHA/8KBmdoGR/EpPl2aRq2LD245ejpki85CDsz+3Onrwo4K
c9Rhd43VIZ4KHqI5EmwPue2jyXW6VEbC+2NPQIbEneA3LA/Dv+ZaPKr9FxDMJPuQEr9FGFOrfveS
Umm9bvKXL6SwikymOQ21JFEcbp5/atOdBXAPkwYTFWQ8QdeC7dg+yE+xcV2TfPPl7lNxahww4g4p
Dg9C+lzbVW6I4nsfwys3ioInTZfr4UBVn/Ob6pNU1xVG35DdIRHPuPK0j+3RjbpFQg4EXF+rxrdT
CmkiSEY7G2hm7/wTUH68aoXAsW6yDhHqq8+RtGFIYCI9KiZYONIRzmg3WMhHbOh0JfIARAR0JL3f
+KG0bSXFUG4vkTgiOkXr/5eiUZ2N/jw2giw3ZcuPUVz5rI+cZ6qjgGeppjN1TyUA9VrUXq89CpDy
E5Nug2RMJj6qrD7D888p2VGpkJFJHZV6ilWiZ0JCkAsER2pqGF7ssYN2k7ZqJBE1mlO8lFa/sKba
qA8ILcb6SRkC8OMot0hChulHF//BLmPLPgOt7eQvW8uy8pQMcnTjI42wH9B6gBjbOfjALTS3nPgt
ZbfZ3xYb5VylodBHOIjVDnCN7ekejnIfv1kHEOyY852oXaVA2wVO4dv3sZXi3ivW0A57bSDz+31i
PjZsAZjjY1pSIMmka4+W+ZGg8lhh5m3ltmQDt8IEPAE1PZrVshHjvsj3G7KU4UnEWcf7/SlIqz4V
/UhWIX/s2IsEzC90nVZLq9HfJaSxUn5FMO5YwXfZSeRKupGO6q563zP0bI7Gh1NKrrAzZ4kH2RtW
2imNCUa747JThKT67klzgbqFzuQgLbONUdtuj0jUkOTJKhD7ek6UnzkGl1VI/2ACbSDITY6mWTYo
ZUF21AvLp1kY9gXyX5ObuQTAKxodjs/fV+u8x8zxi12HCIXvPpNfPWnpZC7J0mURmOovPhMz7Qof
PxtgBBlHFsOUVi4gng+XhDCXpyGSIdqjxfslqL/cUdVVY1nCeMBqXeX05wUDN3Lh53KhPGI7Nq5J
v+UDN/Aqb5vY06YwLteDoZ0rDtUYse3nO2WW21JtQCcnclIDqf8z7gkprmvO5VDKPhh80boQsYaj
W26ubumCUziNkfT84toc6OItxl7jil366HrzlJi/aflw5tXHWfXkD3FzPZkUlYlBoShC3JYgLTVd
s2ulJHhFIvQrhPDJs6s2p4palzG2FUikNI9yRlO5WLfIqkIBq7i25lamlSFuK72KPdxZyKhUpyvy
tE1nqO1HCnnUVNlxugDdDtbMrZxxihuD9FrcAZ6NyoJSHDdeDj1rUhbx4X4CphtEqLeJvqHqlq0m
EG0hM8LMz9Z2Dn3rOvLyOGcdZxgOIt0ndo7JVAaSSaa8kBNfmAAwrVyEZ9St6yEpc8Jzxs7RfJ69
dRkjW2G2ZkNkuZPGqw079rRAp9NpS7cH0RlLmKtrX/mlXQ10+svmHeZLFrEoLDIE7sUnSMNtWSJl
4zyXa+MkKGdmsSsspPqDAEjGd10FE8SwgYjDfNP1qB19aCWyp6q9n0jl26z1rJrV+CCM/pLREJZF
LbZhduotZ/nm8kNnKizabrzMgOH6b81sNB2VfuV2W4IEMGTN1bddHDWfa07OVOXRiYCS1Ep76bUW
j6iZJ2AtaMLrzhNRSZ0eRu2YFRx93NEexRRZUQ/cHDs1sP7UHXkIWESSZhJrSOO8QPR4Bmzc6bFq
wmWPiycBjMYoC9XqJDaNE3wDzLtrgfAg10uWtYG9QbUDPNb9u7fNhcrmPJymna3Z3K92saoxZc68
8uhaf4bi7r+rE83NQtTekcz7Qu5vwbAlIVXbZjROVe0Dql+0RLRur6v9S3Vla8UiNofW1UKZxs98
CxMPdigTqPWTJ9kK/y1lC/cXhgqpHhpMU8/3cqgky6WVvYm+fw0IQjrsvASCfYZtyCT2xYskLm1T
XyI0c09pBROQsB4Tx2RExBfCgA5sdxIquxq6BJmIQN5kAWYLgsnbSFV+9uUHdP5s6G1P6h23Hi2h
1MqqSPIBSAXTOnOPyMgLMLmDaNch2Ou2pfyjV8eVhrzuH4GuiC3wRIPELTx3/gUEHQ4vmYDzMn+p
e3UJULv9FvkXrVcTuN2MCP8Sa9Q0ItOSZZxQJjU5PyeUC/CPVMnTpgbCL9pz3/5izb3/otV/2UsZ
YWJ3qTSQNhM5CovL4LQaMpX2+TNsgpIKb4DjiixvAS/6ee2yPo3Ogjt+MjupXa0rAZAIIQ4AsvlB
QU4VC4Roac3odoUFUnnlj45LEimQyID7hB7x5mgZB0W7mP9EwFN4RCKtqOF2qUDHz+qzhsVjdTW2
HCEGuA/n0TGT1n6YCwyPyDACyCfAaghQE+E9/XF+JKNYjGzXfsf7qfFivZLhA63HxEsb6G8uBAQT
cP3XUoykybE0o0i6K4v+tLjPtZRDWsSMDM5dCgWr9/kLxJh5+7j1qUAjl96UVFLPl/z+rZ5OipE1
9Kw6NPnmsO/osK5x3hrS5Vrx8boZMPlq9qhfIQQPXlzmE0aLv8tIKTdaCiblY9K7dIWmpCWz1fKB
3CxcDZLIvdWlIve/ji2/OgateLg2SpA4H9AhyekVLfDvBbKi68V56+NIxeqsXnOifd80YgV8kNAE
NzaKcXtLzdtHdmCt8XbXqnT8VK9wLFBUqAZMk3WW+/RfYVdE2w8RrdImgqdhWZcCQeIz87OSeDhf
CyHpNEqwhvrx1Ajvvx4yrxuobYilUsD2qtQbJzqngmVBM/6NBJsE5uxug2Du/Nsp9/StDLb0I1Hg
y1REqnvFmWVHwbBn//zZ9DbbOU/yeS11/s6DHZUEydHeRgbN05lcEJBB7bICnLs8+gynxIInZJ5p
Hq8dRU0QFZLonXiifsJoEcHqCZcsKCJicY+cDKhbfYorp0p454+Gw1iP0BremAgPe9olXSUAtUtd
nBDrrM0/HBFU+gvnMVJ676kgTU94oFJy084WQhub6zAcKT3s8JKdXzYc/wXsdvBvGluHCeXOJMFY
wQ5y9AaVOLsm0HHuhianqcGWMfhE0MLhGk18yC5R4zeTlho8g7R0d+Ezdl28p/vYdIc/zwEqAMqv
QfBGYMXWaNYgcXPsq72DCg+fZwUBR/BZvTULtLhGMrAYEHgBtlPWVHSI52U+crvuLwo+u+HRHPa+
TNiYwQ3d/y/ICpWZMJpDJW1BeSAOzqDA6HhSfpOVZo7udrI7OVHvaOcKqC91PlVN7V5xhqCwJW6z
KKlb9J06g6yUf9RfUi4A6xSawozEsNKyYdCiSm19AXw+5ktlmdLjlAc0umla5he0twEYNR2Vgrh0
IIRT2poClZhELYaQgNWLMdSXkHqtmI9+3h/s5OxyjPEM5h0kpftuadmgvSMAxtkHCDem1jv1AQ5k
iN3IT/TF6y9Ojf+zcejUgdeT3TKnwEfQp4hXCHoZA3K+JPg8w+TWGx7uNcgQhoxzX9qZoNj/htwi
prrzZ3EbASrOShJGhovpjxIWNb4D1SlT3PX7umMw+YoVAOfUYNBUSdRu0iUYeEkxlLaQPbi2trYe
WsMd8K5gw75Z853DlncI/rnb/wIKcKpMG3aphHJeuseFXu+HDVJfmVNtbsI/XtGjh6cNvFulk9Sj
BbNLwqDi7aIAp580A5qG0xLGJapa/zO3iAnZN3Loq9c08kYke1I0MhtE1WGa/w+UYLQ5Y5O+jXkH
DalIuhYvJDIodsEQSnlxMUp8GhcHiN5z0l7/Cnl6U2nIS61+3AEBKg64e5oLxX27D1R/7N26fAm7
7gKT73pBoUA5H6jGYKUhM+XH3kstf2p02OnHo5VB5nYeCpbSljSZp3Zd74F0bnlk9oGc3JdSNCJD
x7HOt6UxWCdADWC7DhbO4Ah2IBNfspdQhPlobMzL9aVDM3L3y4wPD80kRwYkpmA5AmFxktwn0T+Q
CAh3P0otIDIoJ0fIRD6z7wEtv+9kxlaT7ZoWAgDZKCpX27BZQuqrvWGQOPmgBQZ6DsScBPWHZ355
fwGiOGhv7uc7tU5RyfzEXEEv5W0ttFIImXwjP0Z+X2UYLyD+6Injm+at+cd6k50ciIJA6e+1iVJi
kyOlNfVnkbcRx7j6mvFOiK5UxRcGQpgjtw9kvZTWTZ3izNzmlLHmyWXzjhzRCkF9PfFYcLyMtk9m
dURGBcoftUMcV4jgsXPwxmnqL+PdohZOZ18/dZwEkvDbW0BCv39er0SzEErNC7xi4LyNoaj073hR
x9cXbHXJdjKKp3p6YY6K9VGFCMSsrZ8y2PMlQAJ9GSs5+VsIiI0bRVPUvpFGl+hQsZ3kWNBd0Zpt
GaVQmsDE1StcoTHAoRqrDhnXEAnw77iT7dYYWSQASunf7vvU7QPT0CbSUwieCu+2ICi6GXHU5jbx
09Qtr/AVbsuwA6EkxnJ/vB/Wfo75SeS4SwDOj08A3UaVV1DB4nffilZ+ZQLjX6DLjxJ9ZPW8sP0S
U8RFQzoi0e4rb+46Ai7cEOhRvF3JFYOaKhHJl4w81rp1NVr7c8D1szkeWbMOFD5pVO3flLukSmr6
8rf4gHlsPfZHosXmUpWYXUTMuRdpiiq5cZaqiHBx04dI3XMIzAcsR7/fyHgw4LBTvkW92MZx0AlL
6zocXJU0DbaITi6MYA5RSPnaZfP6e4RLHXC7I3m8maeej5XhNCM1iSThd/hkfd6mVNgXJYnPVXrH
SxNIr7h1FjRf5uneWCXqPIb+EXzKVkwkWUgdapyScYEaAruDiGxO6pkJYc4Ozj0PxDpdQ1l8VlRW
QiaIuJCXMCBXHPrAUHup3W7lW0LD6Mn6HyKtQFkpwd+ViB7nh0lv0JP8eVcWfLUifGAY4DbsZ+or
BaDBVA6Yupk5Ch37zEqy0G+Z+DqSeCWQAqsYQPzDAXNEzPuTxV875pDa9A31NT/YxFVlOouN3hzJ
f3Bpe8CPL5c3Qzp/Z/spnAJAz6RMPZYrzVLipxB2qHn47rq9lyo3hQy+RC2pLpjOZuaU8ZaNhbko
NKR4DWBCYaBWGA95tN/v3DPr5HQ2DLf9bzihsCYkDDqnAeiwpFKjhi1vSIs2FtNYBwdxwsLGofVI
5FYRjQ7D5XfbEjuS+7uCTTxcvBbeA2fZ8wjvQCv8PsXVuvYKyfB9mZd7zcqPgouyefm+cYjenCMB
F0EcB82aR9V0/xjv1sN93fKxgF3H0kJou81LrLp36OddFs7GEactKaha3qhl0NmWZrVCZi5aI/iO
hB+g1LnQlrC8FZdHSQKxfiuEU37JxxzIxfOIagSmrAWMDwALuvQkk8SrOK94DaXGIVIy6j9rD1Xq
HhX7hBNGvGZRFD4HtFucKON4BGxUM9O6rmD1qG0sCNji3ATWernkY/AhGB5/a+LMKD4uwsA2uPoe
JsWA2+HlTrd/EyVXsIGSbaO53fyqYVuIN3fmD84eputq/TdsuGjI2zKwQPK0RgDfrv5dvqQEv+mW
slwjb9258ao2Sa9EG5+XWXbSuvSHYujzeLLAI+vK30iIvaPO74by9VVrbc6nKtxqIxnrJ3POmn5I
5CscFHbYciJZq9+tQOfgO9Uy42zmyEtvRqywVz9oTGIn8dWhA3Hgs27WsJRDzLS+3HMKlbZpnVbF
eghv9s4V8RxNbsySjUAO229VVJwCPtYp6Gy7dbhF7aJJMFHNFE8U9rQmILyZueprnCOGX2/8TR4f
SnSUQDGnDd/nIKN+yUAF0u6Xz0eENcakbSsZ+SL0Fw6eImwNA5M9YT+WLAhoBF9IXEZeaZGfvnw2
wGPn7OaixoYGUAs+rWm6+oqhsW35qZvyJIfxp4UTLAvaLy+9YynjujqGlPjb2Pm6hKaIPRE8c5dj
Ohq2EMOvSUMrIn1A/xPh7nzEKHY8UHpFfuDMuAg9QQQG0I2WjuSvkBdmA4I1PXQsS7XeMLmqVpdy
/xWm4plIfAmBIsHq5zAwCxtgW6AadHGLZI4+u582p7QOC5xcThLyASy26KesX4v5kHJhYRQevg2i
uUosFQSOxajSKdFcezLxZIUWwvT859YMji9oLmPWaGugLHv9i9ZpSzIHgJgUGgKzwq3G+DUVZ3fX
PwiTIjMCvgQO+mA0dP/SZlVvh7GChbnqMhuHYzfeU9xD1AtdnlsukSJPEiQQ3R274AsBZXR6Zy/8
6j90qEUDIi90nsZBGp8wjkmyLtpNzNh7Ob2CR/MI3PX5BwCh0cGB9usyDXqiSM/er6rvSEyYxxuO
xPuNLz6q1n44ZjRll23qyXBVQKnCdN1ZRQRGMVROGCBzvk+ruJMVhP+Issg5pLbH/x5JN6+LOXSz
mWihhYKKURtEU/tdqjmxQMtis8WGFqLbDx8ZeySuPaiHcMs6iUeM/NwWkx9l/Ph9Uac9ZhtBKQ4X
CM23SiIOiaXQzWUJ0dn5dczz/aNcmLwdfotZmoSuLxei21/L6Pe8EOwAEev6qA+ronDi5CQWUxSx
5U0b8BqcwMgGXTN7wvesh0aXQkHML+WoF1x12BejrUdpDXgbRpXsdSUWUlbl9apFFl8Nyd0HeL72
1z1G7gkMOGF5MH/ymL8hER1YCkgF8YK06lWto84vKLvLnkhNhl8vv/N89UQftfcVwJGokl9ATZc7
/0O/6r4eJGrW0rESoyq1tHhFY4knMzwrniBDSmT9TjptPnoIKOyeJT8TI/74FOGiwJ5f7xGS081J
naAWyD+BsrL15B5zjpCP/GAYVR/XsHVdcUcp0M7nIWD00adQ9TkV+X92qSi3tnIbziTxjNtuM8Lq
JcFncPiygzyt4ZqsIv79hUv17cOY97du8GxfsmrmbFPVrfnsfwKEzWdlRU53XFJwwo0xwqjpa0E5
2+79OZstDacpcFpwxKDn1pKHYbQApPkPOhChkP2OOaRqY3+vq1QTXH7qJkrSl30a3G4w+NqPiwi4
fJDd8xsSYEC8Nte3i63qiPweP+2Hb+aoPK/wAa2chzpV5BP+FIx8Bgab/wbvodZaKxN/raCoH4mJ
ESldgCnR7BA6xAbn0VGFbb55EW1pzmJ27dVt0ezxYUMhlSgyn/2tZgauazwQ7IzIvpnC1UBFADS1
TXsX050VxPHYMBRlylnJncmgHplltjWwTOziCXnhYYEV4LQBjqbllBCZF6gy3ogO0gwC1AJIjhpv
XpYg9oJMBPXt+fSlybT+SjXUtWnLfLBhE7uFZBZ01X5q26911sAYWwgRs9tiZd4Uph7w6rzD1t5q
Bkb/cdCeyLoJw0/zn0zQYioTO/+vbIkl0Z7x0YMvMJGn0qLlyJ2rgElHbCOmYu8suD5cGoayR4EE
x/V79y9SUxd2Gsc1RuHXhCeC9KhRhVNwuKVmu6RBQCqYznVcgssAMusAwMr95SjKaa26OQnNCdfn
mHnfuRsvdie9PHBzLWlvfWRHn0lnpGHV9yOj2BXla9wRRJ4VfuIW8RC3y7EPLB6XzPrzYLTL25D4
idTrRfm0rzEKKbsUIs7oaQvD9wfhuFioW782CI9y/PK/yxJBBgHczixo05vMSlvEn9lSK4imG2/R
uMQRnpARv3JhZBd8m/2l7YMA63y2H6Bh9yRTUTHIr1FEuVXU/LMnatSltJMREOPcnJ6Kum9ntxas
fKSt7mg2Sbalqbesx8+ANas8QgD4HhZ0+6ZK+pg99yhKNrGHdbbI8iAVrMGXA1AZIHxFVRVB6MWq
YzBlkRjak6c7T+C/EKXNEJRNqaJyJTxcxkmFQiJHgNYE9cb1iQFWHTRrU0VNsED3wkO22/BV5PIE
af3zz2jvj6L+4nfMaQ0bo1RfVdgvK6Ni5uBVYQ5XkNs/qMxaxNBOb38OHJq45zrKDHPngldNNe7L
N483hFrkOYFkOmSitPxgj7RcZRimdxePimSDxGoCAahmu4tu2RDevpnWA1rL5CVK/MxwHmiBX2BL
C76F6o94mnuqiuAc6Dlwige2FF0ErqafAb0MAe6nxecUb+YVyQ4w9e9O+65SH6wNR6syIiVA3NTy
JtBwZEkF+yRHdPXFbx7eaVpHCaBG44lrjGAbwnlKrnESih6MgAdLXphNGldCDNFvROoZUPvN2feP
S3FxjsmDDYO+uuhrLWkwiTbsbyUTV6QGA53aeDKOzTfEOerbxa3i4oU2XrIa96PHURnKmP2QfZoG
zXnp2wO+6c4PzMT/UUTLQVSPb4KZL/p50vydaD4e5vsjVkh3W6bgFcSTRhcJKN/PJ/Q6Pkrc6FF4
x3TaS9bwG7dowK4uq71MnYwTEKX3gViNARcFQg5FQp5ZirAenK/2TB+XGd4wNMVcnnJl+j8bRsM8
cDcme0CW7iuzH+Jx+JCE1D7vYR2IdxmOr+pfVJAiGUCsPrztr79GyCvjkzu78cDjLPFl3AhQstWx
WQm1qbAgwH/+BiZ7Vy+K1jcsU4EhCb0bRSTI4kVi7Ob/VnbgIiy0344KW7OqlDQ6bMC85KZqvLHg
EIIUCM4jxZrya7ETTr1KUST/9GK+s6/zFmYSjV/0AOS7Nr0UdKxrsmRPsZcL/l+vvXCWc6vEmORD
wrEjJu0TjWiqgl5OWOz7/ZlP7CALgkGnGjJHhvx4W5MRzFJVt7ntduTpWvsQEhA5xHzCsCIc02WJ
lbA4y4wdDtTufi8XFwPUUgoRGUQe0HEq8/tOHDUwma16DYzBNiGffgiuLWUDiIjchTc2+9vhET7Z
WrdjGf7uFT+0o6xCMhVTeyk0aOmIDCaT5lrIUhPgNLe9A3UWtlNF1Y98ucgzVn5QeIIb1uyphhWE
YPmTNpXGRGZdTuY96SSP9hTIBczODSwfNjw5YOeema9H4NmtlwvEeGdIrq9gv8Dn8qM8m1OOw2Iq
FXmDt1ZpbhkNxPxQZ5Nhr5dP7G8VtCk0TelUFffEQF4Q4S/UeIdagMQ/LXmmYO2cm5CyiJzVgP/S
43tpZs85QHyAzYlVqOni9pxABC7mR1JlkyPLNDa/93Yg0DkD5ewtjZWU0Zsw+Qnu6Jwf/PBBeDCk
jSWdGhjxVbV48Vu2G93VGpiEW9kmLTn29SEmybJoqfgcCXJ3BROz9BLc+sta3F79aifA5cdEkpaq
jsWSqKHZSBqOWYWR4LxdPaYE9sp2LNOlGwugqRzjoLkitCEEQAfaWCOqiqPfkGbD9CdWjThTdw14
F2kjksG+XTrC6C4iTB9oj8qgoXssFuGJaEE1UeQZXXmHAwEPTZWtnCmFy43wSGvfoPWlPknuMPrW
UBVxFKaPu/nOeE6rXAT1bxZcSOmGfw9w1x0ucwIBn02vGviurJcxS9uC1kZxATrMk9PjtxR+Jb9S
Bv1hyw2KxlZ8xTYWwL44M7lUd7rnWQ/jxm2a0mczzN0hgSPxd4R+Uzh0JAJQBWTetfB8qQcfB+fd
1LAm7MJdTHHj1ECkEt73fnDZ8ItmAOJoosg8mhG+w/PKYd+yIpJk5w9udtQZsNW8ZgULPeR0uVHb
hyNbCqlTkcbwjMcy8RUJVNyBJ7r6TcLl+IoX5wCVOF1QM+5IZ9t4wZWueChDndeORgKHtS/dBsds
36O4zFFFyEi7RVpDTyKOMvXIfmtpUUkPujVayp/nHVafEpBQFZvF4/+xG/JQqJfMCSKRw5IXVE+i
uKJPrftXAJMhCOD00OGcVxLzxkvehGWZ5nz6Uj44P99zj5yfO5vKt/EP+duxDkMUb3D6+gkkXweK
RQ1KsLKa4Cf/W2nt0Cggtt09pzny7zZhyGatBU6i42Lyk4bir7C4jszzMlP/HIj0uKyCinMWDqPh
+2G5nLbdDzB8uXSdpKVGmeetPl/IoY0jDF0wKz3qP+NU4sukA7fdEDoHKG/asfbTqMepXOvTo84z
zQQhme9Ab+IE9LMbtUBbyi4SHv90w4c3dESOrrnR+vncSEE/mBevAyyPSyyR5YoGdY7eJseC0X8R
Hb9qNoka6EaOPR9f0KE3NiLt48xiH5ADl3+uRteaeV2sjoOzV+2KoFKvwaY/I4nQJRDefftRUcg+
IIivqftRQ6fLG+s3v0cvXE3G8IPFl5WJo0+e7WFRFPmoVnYKWIKfEEZlh8RWhSyKNLuC9b4/GVnG
+gVceTWFlT8Se0z75iLbtkPkenfyVnzn3UWSV3OZD6MVdawdzKDVC0P6Zsv5j3s+XQ5UbnDYJWBW
4U5TAgTQGIk8t2PJeGfJc3JMdg6jmp0gHQwqEND5M7EYoLddPde916MCECiHj0xcmRmH03IgE9BP
xTMmnIfrh9U7WTxh7cE0o6tnFLgaXVFZyH+VnH8wsd6GMv9p66+1TuG+E6HlMqfpZKFF7YJeFxjW
e7EHUk0CuVMzf7xELGbzMVXuWvwxs9UAYAXG1/piVfcFtWQ2CEIqK4lNkr2Q8eTU5R3z7JTPvEGI
k0owmPHCkja9G4AsCqSs5G4w3GFuncd4BtPdQW7OHUKRWXDIYlj/RYlU9utWUONW1F9qE2noUBn/
RCh9WNfEK3y1An/hop3KbFREYNHpJDvh2i8TlpEeYFa2JIib+sD6si5YcpVeVWiqAHfaKoHQph4f
eMvMcQ2fuyVICh/1npnBh520OjWNjA/eCXYGt6o+X7EHFWB3eDMupkLfm1LXB5DDMRUdVQwpryQa
SPrV8wMRZmYvLwz5jfNczGGxMA50o09RDCYmzV7SHm3tOmHf3rowQpURN9plLsXZjHcJ5Yyohabd
lTln/M6Y8sgw0NHT4nmCcDnSoLXAgEM+4dDkY5Ano4bj+dmXlDvCizhm9iMdjUMVgyDVDXnNLHGS
qL+2I6o/8+5XkR2y5QtoOkh/Qq8H/WXFX8yDhhSR65MvXMUaRpbwA/OOCOw4+CJdAiCedot3K5oo
vtJ10oGz7EaZJdnPJbJn8HhEd1wwuXL5EKycou//t0Qxmm2JizbVoWeYzlKShPnduHud/t/iXGfK
daFP278xCQaG1g6tchVPa6VD5silO2BwFUulJq5DW/tBn+F7O+/MkEDQyW9qBCEvQqcxCvSW9CQt
4TkJtgje8G67SPJoAb9E0A6AOnWjUVwuW2fECe/vOJpoXBs935J4fCI56lssI0EQAmj5Y1XX8Dtr
ye9EftaboHN6YzCt4iMtmcjRqZWklL1GWJpyE7F68qQDb3ffavOJo32fDQYAOOU7GjMEmG+4pucD
1OnR+yuGO4hr2DrO3gslHIBF2Nc7VhUGTRKL0Ui9aU/fxKzbp8Usex/2ttRWc67MGPoClGuOIqOW
L+Qw4zwgPzL8kO0QjJJITDpnuFyfYS41Q/w/I+aPrghokzGBtdmo7sRz5Tj1i5eh/7Ag01hHkAy6
Pu5wloi3qJpCw1e/vGMeiwJM3btt6BUTEQ/vqbA2UfDCZIcl3Pc4/LAPJbRW8XQu7gt9IbuZ8rNk
UPfBXnwO5l11b2cYVuRSnQ5qkDeg9gNgwjtKtOKjHTpCWK1z9HMWYCdpVg3NkcEejhiW+WyzELeA
BCbvip6TGNqoFVIjVUM7OI9c5pvX1NatbVHUv4keHuu0FLR3N71JbT4CbO7KDvYQ2xu4vCs4Myux
QpWGUavyZrJSNF/E5J65IflZL9S1EF57hc+FIkmCHsNrrBlgiPpyH0sm58kG5II9Nxn4WIM+HKp2
S8Oi5GLoVPfeoqXDF1NOrWfI/zfxvlKFAGuR/OxQznJRVqV8/30vdaurRwDFS39nv9/ZZ4oE7dfV
xs7n3RDZ7VsEXkHPJcjh1jTLTGUqSu5m/L7sOr/dcmG1U1QnVHPmRyVL3YYvkqc1SvpM6G4agLZk
GLqZk2QsKTUMlrRcGDZBSRdZeJLKh+n75kFjVWtHHDefYOxZZvhQqh0xLIUMSVWWbd71m1IGC7w/
6CUFRz9JItMW5R40GYP7C9DLr00gXJsRDdUzjNErLbxk4DOVpkTCyN16wHqATdRroLZbOEoQm2sv
YOmIrf87ebd3kB57W8lvrjIvOaQc5G63yYToDpO0o0rnviLQrfTlIKGd0B7HyI7TdxJvg0+fi3xl
NLQ6ypMxF6SgpZnUd6p80qTYpMTncgot6fmziTfGG/ffSzLqSP18JjmX18qSpGzzqtjQZ8AP4qb8
Vj0xm4QhvCuHGBfkMpeUVdrg2ZiIHKKM5fbHxHoLt0+zexc28NmWH0eaGqBj3JtLQyLk8Cst94dD
0/pJjehkvWClL0vJCpjzwsBhwhCJhzyx8hkd8MyVxuEsKdVqkgTse16mqIJZsogK/vo75nvNBanr
8FXKdM/TJTkjZIkxp3F2HJ7YOMmHbCrQVmmDhA4Eb+PNF/NkyrDd1+loUrtd5aMfNI5tomSzOkO7
9a8+YhwugYHv1v0untBn8lwxAOuno+gAzbCm+9ndMRAeWlmdwPAxHd/4ksYAfr4/5eQShRu+wAHd
wYOdWNgBGQynsj06GkmBLI8e8buXXFUYs7FPpozvDiaVBCmIPxqwLnI9E42gRksqZ5VBoJZMFtg3
84qqoYi20c183r2Rh24UuG3WTyM/qM/h/ExUKkPLYFUZmgon6FA5mQyr6JEtW2azuAK+hVdyNA/r
hSUkoH3UdwndT8dJUlpLI+CZ7BSzAZsh6wN/STY62PJK6GiLTnPNS6ISXJ/RnZzMDBk9vboNZrp+
KXApJVwmocAdnm+7ePL7f58DMujgRnOgaon6xU6nU+0cEUDroPz1mN0tQLhzf67edDIiIdfa1IVQ
TJxtupczG1dEQ9s2XSmWnpftHyTxooktdAR7mVOmCj6ioLqT3BYanXrNcncuWAH6U75UkMCI1Xjr
gL2jnrY0Zf4Lb01Lia6quakzmECXy+YOqLkCEenZ4CEptDPWOuOOvP3bZqILTvnIzAjCjWQZ2BLy
ni+bBfCCxkRmbVBAOKh0GCj5hrEpTXaUkkL0n4iD0xHWslpypE+4pf5ntlkmLXTu/b6P6e1JHdOL
PpD1hxYau6yu6OmEqDmpmYGnewRoy1pBV3nNDBsTqwgPIOFdcP508OQoZdZ+/K/VKG/kKzLZcb1Y
ISbqjLHHyWdWoxV9eb9SF0VKxorNbxu4ylyLR7UO/vTMnMCfKZKhfi8iUNMKH4UQ1cXFefBOSwrI
Xb5iCX/7aYggr1orgD4zcHCQnBBZTfZKsYmhFA13vb++lP9mgjuFepFZXmDZpVR4u9tH2Hz5ZWJQ
rqJ8OgI10x7z/nkhcej1/1yeGthQsN1V+xlr3hy2PDJoIeCqljdmUD9hmynRnM1PnXOAFlZUWmlJ
Xg8FAoc4zOoMHhgMWVbcOpqwEqu6srFCg/HHYdwdMu6tmDryW2tkOVp0JEAoEkzVCVUGc/V5GxfQ
Ak/68+2PdNA7IsNirNANZTHDukE1mS66FaiRpc/k687o19mMojxSbICRQcxICttmCy2gUIDoMY/k
UL01yig5EQdbeYvWrtJYuAY1biw7NuzGI//cTIwsgg6CVdsVXhcTJ3PNgR2LsRbRMw46x0ufw/os
KTi3tNLPRgP0VqEJWDRpLEEAiaW7Lrvi/yi5zMljyvK8zxyZ/nsfkFYY3FVBDTO0jqacurw/ztGo
SqHlE4sYvCrWC7WApw/NolebgnGmmbDoODirTBvoJfABxZ9MJQMxp8TJ73YqeoVpk+PSkbAujzIA
qPjMGSVrz9epZom+MboGTHIntRNCULvi/A4FKekK8fSU1gfV29sg5pRM4ALKCYcipA3Gy6uzPnTF
2LTSAPIY0bHyQK13SlKIZSC1/RepKulcM0E6JkAIVwTrX8X47k/98zlEvdSx2BFweXUCbIV6jCSs
JYxK5kMxhyhoCQmNFrWNwBVmWU1qu9nkh8zb9dwPMpPoNlcKpjZOR6t1hjs1hR6u4cKl8GkTMKzo
Y5Ekql+gbHcd3WopDn5rbJOoyFpnZGbUFeDRz59li/GvZy8MYJcogL7hNF84U1r7P3K2pJaKi4QR
u8Mw4B28LKSZ45q3ZMXFwK+ahe0mbQerHUyX4vFYkRA21huusqSW3kJKhC8iJxd2PFXbbf+jgO1O
S7TyY+H94ao27CgfDA8AN0U3JZsGfEqASpfO0kdT0x+VdEkh00mwKK3aT9+2TcmjUUlAAe+GEj1g
+DsiJuKGQnRW1jL+ogFx8z4Nt19JIfG6kyCHT+E0HRujLOa7o31zGVwEZEhGyge5IojyKaCH9G1x
rVEqo4vaKTZbswCJVEUxPO7fEcx8duoprxBYvtxgxJYtTuq1ovXnwVPlBh2PuBH7ACkjTfNHnabr
zF7zQkhlIQ0bc3a5Q3JoXH6aIYatXIN/bNN0cZNQEOTUyStzGvn2EHcVqdQBoMS4JutJH4RZNGaU
JWihznRjUccrKct5+Y8eqbvPWt7wmDgmjXN7YL3ATMhbZfLpIjZWGabxxpgulBesxpO0u5jKTB+T
Lv0zMXOVgZ3Ave/4oydCTT/xsfmBV2qdmewFV4kITFAjFIHBnFUE13FtcDV5kyHzTmknp2QquJrZ
HkeojQGwE9bBHsXZKKyRBXt1S+jCgshQ88B51jgotjmOHlvWlCAq7RmHNn8g5Hr8Jv6GhzeZsVHj
g5xtfw9aHniKzRcKBwWF/3DMiVVnLFQ300jwhD0H2a0lBhiVLMP/CA5h31KjBI6hNnIYc5r+20mI
KPA56bwivhFhOdBWRwaICgfQ0IrHwdyxsdYvPm6TObLe+Cl/YoZkAHzMU2L7fR4O0+pTPKjToO1A
95zHaBAQG6dedw6IAPhbuyEb8VjYwtOVVPc6N7pEZ2wKCQXMR+t1+J5xwzNF8bk4sx9J7be6/fpJ
i4vZ7rdqVC7hSMScS7CvyWYaphzeoT8oJO/JXweR1kURrD6hIuxOdSo3bE83YUXdxrKMJ+yItUPi
rczEBsLMfZC5mP+Lr0dMLIeqHVPdW4wjPrCVP2hCckeIHFPPpnXghRwg6TTORob2k4uWDhGGyV99
XH5gaQztAkLbohn3FK+GrzG4hl2eRp6qByWZUWqrNS5XdDXABFOPBL2/0OasSXfT1/iU3awmVM67
Beu0BZeCaEXb4HiWBGvOJE+qxtDdxUoYtEEySPGI4yI2f49YwigiRLalTYFzt06noNySymTPXD8r
wCvOWvs8YxwehycGtMKPb7ZWTTqalhxo0gAkJhdImm1SaGilNj2A2ScKNNISxR01jcwB5UL9fChE
KWHOjikQnwklcbU93GSpG65uAyf2+R5jiw2Wytg4guU+HNtaT+9/jMvz0NQaSTJq9K1P2HEsTmPb
5pUzit2VA8B4TdzkjazPzuK1o4DfqnESeSPKZGYo3nfDxOSA7URRZTjh9sDg8rBIZmIy56Aawq4f
GNWun53Rv0mOHWUQRFld5x99y+ZqYsKvDa6zq4rh1vu73es4JyUZBdIICeemdv4PPRR48buv82iD
xYc2JrzXEzFWQ+egJm+GNEphHMDub1RYW03aRloeZWve5xe/TU6eUfxQFRybhiXbb62+WM/6nanm
vei44VqPa11P0MAk7wrEDcgQOwd90RIlAZ+l+ltCBbdvxjZXnnLS7bbSGsY12yeBygqgJoWkZYn7
WgnxrGpsm3Z6GHTouDdkx3vT3tGzVGIEp3QensRsC8PO98YERdn39mr/TR3eUbnvje+d6HXUr8qH
Qf7AS4qqIwFt2Gkepx0DhBTV/Hc/N5XJ4mZdclQSujnHGu3rzYlHUGgBWc/VFGOPBU+xYdsVp6j3
zmJgsfHsFbUicpaLh9w+EzUQyrhoJvr5QOm2VB+znlL44IMuvAe5TR778dJH25BdXP35MK9F9DAJ
aQ2B+TOIAAk1JxpXTVErNL8u8oerWpx7js6HUJQ9/rn/sZP0XBsdaW2+0QPfnJa9//G5kufsZzhT
xO/qiGliRng9AhrDWhEQ7iJ+uRx349Ivx1uPBskEsxLe9LVbR3iHEopTM6cqWM1ZVIx7d7uZ5Xh1
RMZbl46WS5BngVThW6imW8bFAePj3fU6eB3R57QoUAn3PSHaH52yZUrpNPKBRjiH13kCKu8OISiE
aDVMUJg47Kx9ozRRlfFfEEaBuPtXb/w6WRcsagOhqFjT0UxkO+C3LhH1kjYxp5XYwhDAvcGI0o1A
gVZqXaMEi6Rgh3DlnywhO3uD/7SLo1sdwuTWaHJT7SnrinjH1lD31Rp0eie03d0yXtFZ1FxUt8EQ
LyugoIIIvsT7xETEXQpXi92ReW2pqTkZDio+03DicTNhz/d7LYAlsBRoNNMoOIA+lZi+Fv0mXuXF
iEuBUPsrHe5dMo3H5MHb5drLbtWiwcwUhHCMRzKwlZUe6d+cE/Y2d5XF0vCngeV+mLRkNP38PyxB
DmdWE5zE2+SAMJjvKr9lSU2iufVZS/QdNVj9cg3UM0gMt83fUtQXAqBL3x1qNEfnwzMYlz4BAUBJ
XY6wVhv3VPzW2FYp2bYyeGtjNH86BzieYpH1N4LYKROHO9zJu1Lrt2oWDbBWm/wcuY9D5ypR5798
DoWkUslhIPDNI4xCYaAAZE8gLBNhJHGvbHVxSjwEUJpow3IMgiK/iq1impvcubsumheENG4RZ9N1
2veyHYkQVKePC/e4ZvDjZHwavqXkfNpUFRi2hkR1XXZtnpDj3D7iC/baPA255aQAZhlNErsQwks1
r1TcZpOiqbHkN3hrzTZz9PUMkhldtTfSTkwsx7He939Hd+KVPz9Bxl7yaOPPiaz+5rM8Okqn2+jr
YVcpPhDn2ODovUD8HE2mx9D7tV3ZcovfAkhNpf8ldAf3s6V6n2wCkh1SIXxkLDJderiBxw+V7Kvr
52E6nBy6/fYIPDtzrHv5WmeCyhjxWS0hVTGhR11sImjmdQEx8M73Z3slEqzfln1xqDuSfwnlxogc
VQzm3lr+gtTTuDNhUFasdslkMyBwh2NI5Ju/jAZOLmMJJu62MWX/5Oz+bGzRVDMZvb407EYwKwfG
XFP118bNcysJPMw6Sh0SkXwm4RLgO6AVuFvNLNVomRE95Y2i03cNCCBFi2HgCjxuqUrVmESyGzV1
osHKTub4nNYbJ9YaqVOzRLoWcuhfbj46CRcL/0qHzLtYjy8D3qmRmKxIX71YOg1oJAdL707LJmlV
9e8ucQd5gFd3ACmbbVol/c4kpauWSWm+4lPtbYX24to/PsdE3kcM0c9qxOLX7oD0huJVvfMdFwDr
xHIe+rBG2PaSSnWGcoznwKkR4sZH6JY7tWlQ+P9Kx84bzFmJ7yJl6HqEb3+LSY52JM36wyOz1f6y
0X85/H5yPZinrRORW38jmFznTs8rJ/4EaVUu0OR91KclP/QiwSS95pbJIItDwPwGJ8DDNXnk5Oat
zVTaDnPagqN2pDxtC6FN+odGu4ocLZSeONWZS4IEcXrjbQDoJ9CtLuV1Z3xd+Y31hlPGqWLNne84
ZxIDDsSttaZDMgXQ9N5QN96uX6PU10Zly60pV1++RmdoMmhmrv8PfRQSgsgSCCRBSDdCncvGpTl9
U0d4/X1pBlTY1Aw24PYjljdOZjhlG69NOiQ96xcuxGTVd+/tnM6NFC+iko4cSF8OkF78ttf8lY+p
cbeipZfjNxbiYT64qUwFLTgB7L364kUhAVXROfByFHxXoqbLDpphaDKMez7JLPd+lQ7GlnAQ5QGn
7NaTnmOUKbldB7VCeinVC67S6EO/IYyutujIhIucT8nwYZxZ+Vc9V+jILTH4Jm1Ps3gVWrJKcsj9
9vWAIj9A3xLCTkRjC1YHKdOCWm+paQVdW412NcFx+GDs51TsKp2iRjmP9vj4PkISr7xX5jXF+MIk
kH5lgXGj8ty14zuVZ35l0f40VO9eTDACDsLo1HtgyhK1F6839uuRj2h2EpmS5ZrnbSsGdgHbDUv3
+T1LiU7Mi2QD5jI9ccViaPRW/o9QLYSCO8bzrx0Llp9CuT16ut3fh88QTK/d9u0oolg0Ir/6iYW1
vwi9+A34nZ3Qv+DH44Tg8/I+a76gU7msoMTc9BtFKUKuvfs2MrJFBaHm216e9QuYchaEVVTqRiFz
bdksgXtnLpLXqhMZ84ig6TXfMT27aLH0xMYffKnIBzYocQmX+MTWEOsmSxTODrFY34D14za/bCsE
6J/Z/fN9vS7PUg0JozORLnQajCAlj6OILZgLoz6Ckz1anzr72GMyQIJZSiL55zKEnIuItqTcUJny
Go4vDScZ4uBfLa2P/tVOFjhbGoeq8csdkbczudpcIz4FfGlG6heken/PRMRcVMjesAwIUg3x5YoF
sUtpmTwAGnLNAHnMuxFMQ+p1oyLusQA95FFokCySBzG7p7fPrxNSuWJVSIJWzSoSYh51k5fMb1HQ
eC8u8NoladXF6mPZd1DLZAUpRoGYt8V1stqpezKbWg8kSGnLAIzy+m5cGjKTrrkydRbE3VW20e0O
YB3TcaU6XqlQBomvZkRqCyGwfRtz6F04eVk8xHfxQpRqxf+UFiOtQAZEWb9iEeGYjJJv+G2MJ3nk
SK03nMwsA4mk4alE3IHkg3WtnpWsSaJD1zVCXJQjmZLnJwFWU/YldwTttCrYWqABB0SmzJfbArvn
5u1R4H4hkQ8pZA2QWQt78QNCQLPEaZg4ANqpfBUlgPEaUH5DGVZyX2uvlGj/7g1rJm/M53UnoZbK
TFft9w9aR2TM0/wwK+aZsCAbBfOcJnmJoLQ1khaVYQ5O6XJnZPWUFgbCqEwRvl0IFVHAuMDRYt6T
5sKMX4+a8M+KyRmTmVc43XW9SK+1diaepu/OmYcwXmjnq3zmB0PG9cOqKEK/zSSjTmheEHWmaNJE
bkDOFRBV6tng4kRqpa21ddopV66b016LAV/YOcORRvG62RyOfG6d3ji6eyVNZyX/MfVnx+Mm2e19
xRCovnTrhN78AV5pArQu3sTWdfJ1pALZCAGimIqlB+kPXHEqeH8B9Tixy9TK9Y4xhYjKeNAdfiqJ
WPTsWbSsZ+1YkaV7jn4yMiADQdlTBx4f2WSVC1mNXyYBxYcHUGJps3BcZovPC4O/88Wbb5JjAk56
aNNCybmHTuoJTQQZocz3bU4Wf8OjiXKaK2/RLcKPWE/ldnZKZeYMKSbSOFuw7zVWq3fjaY4ndaK7
W+VVclTzANn4DebF5XFkcFpqhTHJzXmHW6EqxFv/l9CfJ7gmJATJCWNeXpNHBtWC7YMVbxCczxIj
2QM/d69zSKV7yooSSmjqm0rYu25oVjE3VZT/nmk++q552D7rSADen+CmNWlLdeU3MGLx7AhGc0UV
8hJFCyHLuqiwsz/g4KZyVugJ1mQEO0QpWOBlW2zjS/E8LCxh3OPvqUHT7PSTxey0iIqkOVTxiVA+
nID5aU+zjRY2Q4TqTBhdAKYH0YO3YqwGZz2z9CPXfbJ/hwh1shUHV/55TNczGAszyIAa7NMNG2/H
vIBJTZ+dieGoovEq9qX468JkOM98ZrkdQoy2ZZbIyDeCRUIsI6+WPHnN5ddIycGTwvBjSyLBXHE+
YSKk55Ap8e3kHvVG608afUq3ihGApJL1LG8tEq3+EVGjcLRJv0ioSpC99ZWCOoXQsj2uaIkLayTD
YpSx/2zECMfIh2QUbhSfDMIU0EaLV1g9qrw3iy/0wedqtkGdj2gqgJ2e5z5MYi2ztYegxtVYSkLb
jc1IGqtx4+0bu1dnMIQxq6kQMexkZKXD0ckBkDDN2xajPtIiKJinJgfm3kf/4vEXHdYxzPeH0Arl
CShVtGHzHbN1EdMsJYiq/G9cPXnIOilR+UICxwAv5Ip0HDMK7nqZ0UPMH12E+G65+1Jq3r3wd6Cc
zlCBg6RPaG9UzW9SLBx1qDHI7pcnLXXfyq0RpqK6FfJD0LUUFjvG/2zSrMLginacUReViFpHLh2n
+sK2yDwYusdutI30+aTldqTZbpjf8oQCOWKUKHB7GIod4UX48MUjzd+2n0qosbVd1/yoIiBB9FZT
o2xbg0buGlGZ+HeW4kaHrw16ARskDJ2P9NYDoQjtIXQDJUO6q3Iv1T+e3tBe0hGhWZEDGGsX5XzI
ELE6doTg0bB7GzVixBh/zJSZWej0asaIVmHMJ8reDSiunCTVcaWpVqB22UKl4Hghnz7vtOmOcYeH
cK4PVSc5kt2yfZC+pAuV3/kN/XSaHwAwgBWrBuxRCjWQJOW3we0kSdsYMco5LbaqRjjpyeKXS1dz
YOmBlctQaIqAMY/iyBF+6wRTugsDKuPKkOzdl0k7B2kfLfHFD/GIg5MDvC3P9myoBb+wsEn94Y7C
i9d1oI6yiGm/0fpS9k+vySMJf0BVmQE08R3pmD1vzu4iIXFCYAxpIrx+CtJnjABPinbWobt/iKrD
JFDMwP0n991hCP2DoxBxeOiUtM8va729gRk+Hkf0j3MBvJXTf8QH/JZk5GJqSVZPQAULTq1XyahP
pAbve38kSSjWsBavobMIUSEvlUTFN6dO33C8sAzBCiXjgKS+E2WTb/3F7gGaSCC/ORt54thw1RH1
oF30ekRQKzesiURD0zNMNDe1Uwb8Tjn1I2LYHwEPfWv6rpzJS6jAsLYdta0cTT7JRWX5tTQTfJEH
GELwX/euYTObz+gMbZlZIx2aAXbGJQQfw8rrt3SO5ypaZxJxR5rfRuaJu7cX9CuuDHdnHMipTF8X
fiAa01KRWf9cCgIlWn8C7Bextg3WSanWN24u2AVpu7B7ukThh3V7XSlyr4mE/3by2lUP54IXidM5
+GX5cowyDCVbyVhRr4wMHBAlUsFx0gNrPaJwts7z4m2Locsku+k5ty4/AccpXNY1God7CPSjfSQj
mXK9/daN4d3vbAEBbAOfGStIqwQwRcdBDmGn2Y/xnijtzIvOVotPFXMEGmL89nqIcOwCr0HejYm2
ytX9MqhtjHY9ZWg1JHKvcDLxZZmQ6ylBBWOrGan+WtNjhjMTD7y3yxL0SmM9JD/JO/P87mtl97Ud
vPyjPgJZAMjrFNfdqFDJfYhZ4mQIPj9mAta1LzPKWSOo+8MSjnTWfAstFgWgcjei9B2saCR6DXgB
j/w4Q2slj5QZKfJvTPQ8mTzbGFYJJRYb/BaCpPvR9lFUnTEQGZWVGR0PcBm9Fvtjwf8S+HZ4/TyL
Dtoxh2zjNaEZsBQGYch9wB9rFMd7NiIV2XurQ8J0clNwVIJo22EcueqMLJF7HzquIHkMO1m/DktO
Tnrp5IzL0ji9hWqUyXXJmpXBnVSSXibobdLsD7+4q0LWoXONSjJjqyeLpYG/Xn5bq5uyBUlG0Wxh
H7hcTa+2+gM9W08rsaSF+8IXwGfXIlRm5BSXrs4dVnVD6W2ZnKi8I6xcSxAVHPrZATqpKPTHpkGS
2oqJPDZOOvGtJa4r4gq7sf3mLY3k7nWajhgSp9r6TIjxOhQB6SWzhKXao3xQSTVSGovBug3ZyFhf
Ra/JrXxaQH3fZ105mBS3qMaGMUdnxpxc15xeOa0MVvzvZjMoa5z+XGcASPq4RkgowYul8J7HYSZU
N0az0jCkI0D/fqaoUtBALBmhxb2QuOia0B/7C7ctgH/pqg5pULix48qJhqfNHQzmgCc1sgg0ZdXv
pcG7ddhRXFEFvI63x+uUrX3U9ev1tOtXuKd6yR7xiCL1HSyd+wEfrRin1+38x+X13VB0NPGNFz0a
eZ0TBzsXJM4LTCGGmTTlDARlubsevyCqArMpoDQhtSjzGJvYioLtU/R3j9gankOW2TmmmelBIDfM
RJejmoDkylP2t+KyuK80RUalMKF9bW/JTNc06c5ZLIfGuLAQDhr5H+VsmKOE/WKgUbYinRBmp0Pc
kI8o8NtzbX1I+JE1az06GbWAO++1jwKwbegyIWSVBIRCXB8yEaCAbdyCPoSRqdt3VtNc6t8tn8Hv
z/qmpfcqIYpUMMrO5jqywGXWEpTJ47ZVUIDcEOeTzSjVaAuA6rVw72hiArd1xXPJhrcBuXTcRETt
EWNQi+WtISmM8krT1Og9nSBEG5kzXEHwrVSDodvyr7UIEy5miMLOb3mshNRh0ObkwQweSxd3NnjF
8sAwcygjqpDCpP4C5fc6S00+wMb2BNQ1Diq1KeofiqGsp2n7W+eGn/j+vj1721D5kzAumO9kcM4y
vzE58XOrErb0twdOLhV8X0u67ZrJtCX4B7rSXhGfHfrr58iiShBOA8GYFkFEddWP69sj4qR7ILLF
qm21Qp1n8VAIjTAQGmBBYcAQFh/0NbP4LV0FuY19rlX6e8FDIhkyC28K6ev9MYbfoGmvhiNGb6y/
sY5dyyHnxIPJi7bYfG3YyezfmYWX7ZQk9cVg1WIFnGXyh+KZdSONLR9/eRG2gS3Me4q38JOu9wen
gizyNy6qOBXLzlQ93O0uNgnwHQ6RvqvHPyJ5E8L42hdp1ePBPA5ML6lhbRwdRGQNXk1556/Uj4rO
4vN3psqdZCUaHLcTnFMSfLS2m4ewjvimmZWZEIQH1JX58LvEvUvg0BQ8j1NWPGQxfDGnThuy3dMi
D3mSe1kkNhb3UCY/DrdDkjldpbaG7vLCQNw6FJMBKMNP/n19TnO4lT6QAOoScU/AYX9/6Cn1Fezv
IVMz2wlMR5iOLwjG2zWEsrVFIdC/8oD8RmeGsG57adXAdETfqLCib9io4QDXg3dK5vc7MYSVmU3i
RkZmiOqFYxUSnBhG+O4LG0tQ02SlYMF+EvNDSqXJtOD+eJAnSgCVIvsMRq+/Muj/dnMf7Fvg4lrx
ktgzrfqHazvMT9TCzOTtqJzvsRIKREFCRJLo0Skwu0wAUVYjL40GIK1OYmKZOegMkIe6D1CqLzXf
Yb7J5niRJtAJHY8WtidYAmSzUGInwXFi/W8ZgmkDJ095Vy46PuDqV08uOi3+blUyo+ops+jOgp65
oCETl1fIbcpAn+AbBRuOCSnjEDwMclqytVqZJ45RLlWcDHjtxRe2k5jZ1e3F43d5o2yCXpEEZ/tB
Ug7u8b+0PjXdFD9OnaT92WQ541NPxgnxaCb00RY7DMZJqrakgoHbUFXUtqZfv3NZgBbwiolP5fOT
yu9xPWcAHIhAsVx6gt2fMs69SsoA1T1LrU5k5dfTqozThQ2mFnmsI7MZWXnEcuMnckjaNDDs3e5U
VNt45AV5jOQg5NZJupGrgYaG4Zffgw9YVgEWcduRCjLu9tS/0Nr7uVtbLPAEQWSGQv6R6xLaBbnl
8Qy31CO3+H+t7Q/okNOngOsouCvsZtFjCWrKHcAiDG9LhQKOX8b8RHpDNPQK5X5Vc/5Js1yAMHCo
3QfzF4qNC5799JJlFkraiRYMkpwDTj6fsPGJAZuBfIwOV2/p2DvjOAByxdgbpVSJqPPOXzWnJ9BB
Jk0KemICIiCe9f9W9rVfWFEPUSTp/tBksPgnRwbUHneNKP8Q217JomBjzqHHjUmVgpyES/hZjpCC
DfkHAAv+6/Rs5xeY1ZLzi0kbUq9AuVURNxoPvJziIkSzDwEYwu9Pjte0GLEL6NTv6ZEfAbI6InQg
Y4TO1PcnGkgJCs6xlB93plwXVxeAzKUkdp4BaaOXa6EzmqKOWsbjM+zqujKKg1AG3jS4Xqs+ypuA
FvIjjmnpOJuVQ0M+tY6fEoWXMQ3oWRu2ifq9TmBOj/GKFAE1qPQ+4SQ+LDAByM/W2luBPReO2jKM
adomD31OjA/U/0khLlSvUF+2l+AiF9rlRkc1R5/+Y6Kb+Rpm2cCBeD2BCnY1HEG/IVc9fAeGB1HC
Y/nci7vYxYwGOjr5nco9g3UITCReZY4xeqwXK8P4tvtX+7ckA2STPwwLU71FA78N3bKJMlmfx0GZ
GZRONZ3mOuGhRvm3CBNyChxGW7sbF9dpuGSwTVka35zjVKMvbSUvGlcDTy6Ra0EM/v02XwAS177o
CGiHa6Hi9iA/axSqgx2GN286VFBISGpDwUK0xsnQd7xfe0qBexgJpMSjDlqQOcrHEkzo2LdYJeVn
0QIxVsH3mtoah/x1/eT6zM5bfIHbrpVUo10FciYsGdwrFGpSFNXNDFf7spHvZ0cfeSJvxlPTjrDt
HT6FQSyrbVdaXv8w8LuJ+gIYLjIixGkPH5kpSBYIYSKldUUkDtgE2hDC3HRZvVYN3ujw0dzj/Z6o
lwpahegBDKo2+iiy3/FmttxCXiVb8PmgX7TJmql4Q7sXTy1nV0r5DXetQ/1m0JxUjsoU3BpBk9uM
lOb5ZogT0kwREKRfwY3ec8dStzaSdqtjf80iUt5k5tta0ErYPAvMUeId3A3oFoUPomlVvwt/sphu
qy9JOWby1IgHIgHPxPYN0lLI2FXOxiLfd+45f74GJnbp8w++JxPFvGQZL2+b/koZ98C7UZM+R8nB
R6TSZk8Ypv2JerqmmBugXtxT/zte92ehdnWqb+RxQiY4QXjfWioSuA7ynleSXmDFXMOUpCk4/sIh
lLLID49Q/8y/9YTY0/683WImQKrJIHwMl/X6oa2jfLoDx9AQtz9PxmiP60DZUNJw6VpANSTC6/S/
lVqZay2msK2svzQkkqiIQwCb4mNZ0UEaK7Vl/kgpHngNtTFu2uFj/+dN8SeS/Tj/5Z13hXe61n2A
o7WvrL0am8mzIik206OrMEjbJoJ/zQrpu9nEmlC51QDEnPIvuTxbWznUXTHO6ez7h9l1IKoTJ+ka
RN3ctXFq5GXSl1l1TSWXnvig7Eg123OJoHNVCOh+Abte0+BmUmyuoZ5RsRgWBmU4rO6H1s6AyXGN
Q2DaVcbj3JRXfM9M7vrE1t8xGUMS/BcIHHEhUkO+kr4OMx12n8pnS6p/fObjSUHL3Z7ht32+mOuC
NDRO44IQpm7JNjYg4QtTpWIdtN3tgkmKu+tnguLrnHmXVuN34ktBXm5aX31H6fwU++Rb6qdwOqxN
JnneayjLIQmmYEq9zNXLyhUKqhnWCTHzvAa4NBc9iIrZFswR0JmGq2YhawfgO4UAfix6u8P1Rt3r
tnmA6MV1SN9P4fsU92Qty7PRtEj9Fh8TMG8SgziBfPdcZrEUIc0AKDDjqF+YCJ7uZN3ab2AFkeVr
/5tLDDd6zr13hZJFh//2u6i17QElXaQNEU9Pw0KVjj1+MCw5Fs/yC46ga2B6pNu3KAkOqKT0ZhgJ
Nlosy5SSmXuIjFtEQJsvdPwxlbgvU5aM2iwFOycnF+te0gm+uH1L6xzpJivqFTAbmTibDWLFEh0w
8ElmIkWucIJIauZ1HKmewq15UNxKEwRimAxErar6DsM1rqEOmDcc1CKhl5OHwYzhpGSWoxJh1cUA
C9Zj/FxWdTUcP/TigjyLO+393Sk6vq5ypL8rvpG3b8Wa+VoY0X/M5saAWGqXnGFo2D7xRgwa0f4U
8lbb/jQ0quYhT+Gwpx3ikzOk9VBOJMtLeszC0BN+q5c8V5s2mFBVd7Wq4tBG3oY3ItBsHmgNOUiW
POAwwMbowgugHiirRlQJ5iekH/Ua7waj+tJQZSDhOBDEUi0SO1MpoK4Gxu2ll2DtNi4Z93U/T2vh
/5B46bCyKQrHMMn6oAXXEHSZnZXAO2/HfEqzzfU0vileljE2aDrt1+2tOkw1NcGd2DdaMYzAyAkj
dyIjThFRy0knDUDvd/n0aLg5mqFjZAEER2HBmGE6QqpGOiLQn5VimijQfanjoieYXO8vHCnYxMrZ
3TWLadWLXm75mn8zVLQPoazJ3Cl94jM5iDwiezWjM2EviMwgaXt6RtFbWqmd/95i9Qydme8rcZS7
eiaQTUwyrL1GD+hiDSaLW5hz40hdsj+F0DWaE/eRWPwS9gtg4LqnhntI252F1ri1Z+Zu19aqE3mB
CZsXposfrMBPLI5jE/wjwO7sU0YNS+r2jdBp5QhpOZQj3FyM4i4ckJMuNPMVQw2tA/LwDu2EZ8H0
AuZx9DjpBHiwGX6ED8zTvdNP16HV7HQZIRYtHvQ7u5cIW8Cp8lFGaecO+hp+/jWFFyNnDx6UgFhD
ewVyJYj2FqHA6GdcZEodgS6bYRj/tiwfQTkWqwNbCqCIzNaylD3vYoWNN1ujp+8U89Dv2Nvd9ydT
l4Wmho+5qHcxeySV3UrUPXKpxTDxrD7Mf2jdpW3ksMdBA3nW4Mj6Nw1EC7xYovu+J8stXpzWcy0q
UrKwnH+9wTRLpZuqDtZl7Q6JKCGRTm0DiTm6IvjF29DdEH2HBUY8zUUAN2HDdhuJ8UAwiswdwv38
0Ue0x6VRj2EMM2pzOtR3Sage/XppftKWol6Ea9NgY9liivI23a2MXiZ4YFgB304V/8Y40Ke1DWcW
7dTwVgpAj2f58qIkEMLu3b20b1EaAgYgInd9qMm6w4ydfar9sqsyRItthgZwg9dbHhIU02+WsOiH
FhYbWpdjDahfZx6PVn+MdbUxrHt/oel57Yx1LhBPeHgwnL/J1SDCh3YTfpVb35VxyeQKPesYWwwO
JcxklHvdyv9fA9yFV2edm0Hmpfbr51NdCsvvivq70yzpvmU0/jXw90XmevX+FVNA8ECjINrQ8dHz
phvrx+AJ9GzMIuOS8wPx8760+L78df8WlHQaA7XZk4+HMCoT5+uzXS+Fr4dgHnDy3m99RZgyHk27
pL9FSMj+fZwcjbu453VfRwLQiFqJcQvnBowCpFyyyBSWraPYqn45WFlQvNQiEegzhUAXF+AWV3YZ
MQaW1rPKOG6c2tf8qmzbUwcN7qoVDjEUBmxzWBDVuwC/yAv52n4P7yh2EIjkALS9ZlQZF8WLliN/
qmXrtLIwAgSIe8b2ox9QD+rxeydXbgE5C4JS4Ood8SRcOueZjAHwkmC1AEM2YoaQzYekrMCp5nH5
HlAKQMkPFjGvh1otESwndJZMZNpfSeL0JnvmqhtP4/OPxg0yfhc79jQkTufWS9c02oUx8b/+/KMa
CDmD3w3kbl7JCZ3SU4jDd8MUkuf8XBuh+eFMoz3wkmsW4kX6BrHz4XZ9UPQwJjdp9Rfzm0YI2UjR
ABwXqOFyePgySZFZNMYFmxiTD5As5E0nQrct+nKgE7l1eOvxL3gS3y+dqTnXF0wPd9NvO9PaMwnl
5/IGZuyZDmrsZbJqfawinkEyJ1xdGF9D5ZQ3cIZnNkq0wzpeIrNT/gjKtMU0dHJuiJJxg8Z8GVMA
6vdF0KMf7eGgjBx0wjrVrFAFdYDPWrUR906qQ97bJ3GaHAa5vTN5w9yIO4d8T5fGxnURkqyLF8u9
KdSY2mwjJr7TlyYAiDMLSotnBM61cyEnV/VZH2jxGvL8uXnLBjUNw0YiffvlvgJBFZXCojfyzU5r
YicpP6t7L7g9HCHtakIy/H5UUZ1ml7cGbqFYh0aIXMiACFCU3YlD9EmeDcWaJPabdNVCy18oc85x
X4SLrypauNyeCvU0rTO5GJ+HipqqgvxqU15B0839z2T4hvnN7synssQ4frsolB1moHwfekbi0G16
u51xQL2AuSH8zwya10kt5+DkBxVVWAiS+0Rf0PLRBSXeAuj7RqvxiwVvZAagkfUfcEXRTD1vhqBF
XMtX9Lqy86ZWcs9zcHPiZL2oFRWhT6s9mIbqYuKR1J9+K3lmN3f1mdTCObeNqyLglwVZI4Y9Ys6V
BKZfawR4SbidSLltfpjnJWW+WnBkiUI8te4fXEAcXxOdxeZxD8AZUstYslveCSlCODSUTO5/0EJv
LhAspq/nfodAFAmU80LQ+1SU5rqrYG5yoa6tCAxGlMscLwAjE6918i5692PBrt+PxDZqwPGtnOZu
8dzHQjDYTMzVgtFBMjBxN4fHU2DRqqxnE4AnQ9a25e/o3nb1lQLkGAjDqWgRJgrl9GjRWhpM+FWL
ZJPnLdPOINNGN1+WS4PYlsxyWE0n5YmcPGR3sgbf3dpYOy85n0pZiGMuOiHkjDgo1VvSXyt/kIAB
ak1SFZ8kcEkbHdYwu2V+FQ5htfiLdZ2ZOFLmCCMnnSIpO5u+juMZlgFDlQYYUNMKGpr96SaAf7CR
v6KO64hZeqkxb9UD6ECv+PjC+olXCd37fRpQPjOmD+727ktJyHC4wYQLyeevVTwGeuAUZHEvp0oQ
RFg7sKO7fMHtoY+1Tw5/gd4LQ5VjJXqeKkKzIHjYNkpvtEakNzSVTJ6V9VX88JEv8KLOcqOStoj8
YttBzGhlFw3KrSjxQtqlc7u0gg/kNQ9vaz1NkGpdhuoRz5yM66HhiSaZMONaDNqC5wJXwrFTboKw
xzKLDQODuYNWNZmCg6l3dLFJt/leWezkjgdtZUOdE2w5BnAlmLogtjPi7h9xyvlFw8Z8fJFvgY48
vCrCzO2T3IHWdkADKkehIVja54XoyP5VNr5toW7vi4qxxVX6doYkJWgJgvfamX9Pu3rOuUJhymwb
HL0inIhFKpYeDhbnwjQervCYN19g3CscmXC+Mzye9SfUoChxPRQrTagm1Eod5TD46C80rJIxDcnx
IW5hsgnkXg4jXPbksfT4YC3yTtoa2ltR7sfdBOZ740i6vMV7l4D9At6A2cEJX43H0nXm6ZQWAJ+g
yotmcwVaU48IcgKNSbm/2BERLu3eIX2jSoGGR/nNtRj74Dw5MEVA3W9aVQ6bT5LDlw4Ewqd50VFC
g7W9TRn6F2nCkZiTsnBu7PiWwMSxWYRYLERN9YVChCsqLhg2gF41ExJsIYb9/2KWI53U8GXhKQxm
yH9zwaGRy2rXNW6iLqA+vYFK1b4i/LLjKb+5pY4IWpKBfrvthS+ZLrbEOt9KzA902Bpqm0ZpQ1k+
us2Wltgqnbx2cZ0ubHUVOoHbnR49W7+MMsa6Dql2OqnE6SGVIvA4RVlzjRi4XvkBKJDbMa2M1/JC
Zu9uysZmQKYGB7sSh1lXVBPPpYVPvhjHSgpx3bhfrEXmDRAYl2+6IeEnIEZlbja7ESNWu8ebOX8m
R4K9BhAlFXJ4sxFIlMJPZNaux6e/J0WUfUmNKzKlsz9hHKzpEwyVuJsrN4T/VzEXA7zdFFZx0cr4
anLKPujRBLCp0IxfJJU0j287TeDi5LotQE1XgAKn2Xe+vGF5RWDNnLxubo4WAhrbfewMhbhC2FqW
2o+JIEo+zRmL88GGwJafhmCaF//nkr/fREyFQ5hIe3X4VUaWLUnEXNtuaip0G3qUpVjWnYgOUoVY
cwwZ5arXQdlgMMMck/6sCjgcR9SVogmsdK0lMkoHwlTwcG1GgndbSjmQ2L4AzIonOUgNOXu019Ek
jwweNq1TDFK7NBbLMxXjouc4jbK2Xe8Sr9LvXQ91SG9BwHoJ3JvS8rmPKCzBMT9p/YnF1GJSRaKd
tamrl99PD4165adQCnMFC0jc/a5seSZONGMCVfLcGEYldCXFHqJpcJsdBJMSh5vMhYvZBcW6dnbV
2NyTEmfQtfaDPSVaod0RS/naOwvGFGgOShYyTn3mpkUzACpvx4opwJX3QShXuSXmW+VCUxdGhWlO
2Ncd7aboaD6sUsP5AVBulEwJmlSUq+fPX3lzEvwxd5sokr44IEhQZsbJYXwTbLEPPrgiuHuU8QaX
LHLBFH+p9NWXqjRpdLZT9ohGpMtjeB1quITn2z3YEJRYnZ8TTD7GtjtJLgXVCC73LeCc7YYrZIhP
AFbtyXLyHa/zbkV7PZFi/Caz1OzsT2XxXrSr3U+hjJoXICAmHKgZQ3dqNAcGiT7n1Qwo3L0c/6Vu
MBPsnLVZElID27Sjqj3XKr+WCZJtFBY3paIdos8tMHxtDLTJyjR5mOiOk2NmcRsM9B7ig+ASiRm8
ZsVEJhCcaqLpqPSsfsi2jKTig3ETmHmrG/yb9Bk7LRGVpp14HFPRvqL7IWlG0TnHSyQrOBMSf4sV
JbZFiIrHrTXqvXNCxCnD+61rzJUkqhMGpty+pGtsBEsy0R5UtfRXWAfqZ4iFlyaT4ro84fszdtn6
EiVhti3vmu/v8RzXAlVhFo2421CDFrBSMIaWtCvYYSEvO0Ay+2AqTbaVQzDoWztb67B1xYl9+9gx
vn03mtLBXFs0r/ewSPWiMSvJHtS42T/A87QZat1srAEmhMWvlEFpOVFd2uRw8Gs9AppLe75v0/ns
3mG69dIGOsnWP3Dt30/Z20KDe61i3zNdlEYboWeLrO07+ePGNRRS3BuJ0auiUO9TMjPF9jfES/MC
5ifI2gohrkZX0qB+v/4Pva+BldBanVzIX6Ptej475msbwK8FAWWLkBgiYk5NF8yEepNkfR++7r6r
TVXOGibzpOP4ZBAy/uWk5fPzcuIMGfKAh+iwIBXqW9XXvbPMVh2mm+DzA371EW+RPHjxwFlSP0mr
FriIluroyOClZlfvwpKX1THJ2F9vWgg+CjxrWlLs2HXJYaTpDN/exkccMDQrPIiERoYvEs+ScVw7
CJYIcGbYN4nxgp5hcwnArYQHhGyWfE15NwC3PrtiCNVqSn+8+bGSf8mjiKd39mPgEZX4duLDXuMw
s6Z8UecBipK+npSRJSTFUIV+1DbwQPfaH/WkfrEuJu+RkR+tMRAzvHY9y4Zb0ytJ58NOdVA/kg8t
3c6xENGrVvqj0nnAc4W3HwwAGIOIxGc9VvbknxhL5VF8aEW7bYOBiwDWE8/UvyBEGKGGJsjnq2Gk
BkCCa7rWF6ri8xdME7di4Idl/iqssDQdAIjbvPbrpbPX4pWzGapy0D6x+4xRxvZDVJjgVPCWB+sQ
PEUkhlqpdFgKkFw5GpikNc88x3qLlN4mdSVy3KjmAqDy4GzE/1CH8WK0fctxogX/KPjgVR2x5Ivy
NDxdc4pmB99/A1iRPWw42sMBupW46hpZN2CUDmpaX8YGHmOzPNUk3mNvRxp21Be/lsa6JkXhoPV4
x8YE0VQx5go0qmkwjk0mchaxzr7H28fPjP88ueiCJbK16fGIPSpPPFMAwzeQrsRfF1jZbORvm4PX
ugayV7JGGTq6owqRfzkWlCulP+pXf+QNa8Nxg7rfZG31SAODz/csfAAUdoQ57erzJ5E8cdhmVDfc
FX3X50ZUxyQZaW3lainnvnr1aBy23itmmcR2amcvLY6f8hjxuOC+/bMtlXIE/hKwr/UPazWQWuDI
62/pDoB/5hnXURqvJcymxqCpjT75MmQEXTP/2ZnmMXgjTlINSd0iGeXQNPQSp8gCLzstFLNi4FyO
ohRF9A9FM5ZMAk7J8NWNGvNrr1pPTjKvNM0k3lIUeclygfYggxajQ8GKaNcJAeVYCLsV2kWpIsKj
xcdfWYffyl/FMSFj/IBucG4pcGMQvx+9w+o2Z/8jJskXnEjTK4EclnTLMZCHQEt5Extj/9pYzTK5
8DhictmBzqHjQgTY7O3QJHVcwYtOqncxVK7YO+fzJgjxhZ6+JsaTtKciDOSYzcuCgmOJgqys998S
rBpY+qx+9SsoBm+cacahl6BnlwoqvwBvIxMNa5B8S3QLgOVlktK2bV2o+YrvdrNLGKp3Z/NEnSmj
CDkU2eLb1Zun8Vc3FuyM54Ju7NOhc4AB5Lzopr69w+hswyy8LEIKet7WmUl72U4XjXbRqE8W4WIl
KzPwh4NIa3QF1eOAPm3jVRkXsJ3BOYyk3NE3U1yl7684jaf5XfJ7dJrjwddaLkFPLCV5kY7HHrJF
oK1FK/ITDcyPXy2xNKyksejraYK0ofA/gSFS/F1ggvU1ikWjh35VUI0iN+k0hPP9XNIueY6YW8un
Z9ipkbViM+cGpR4w9G40PUZwJ2f5hW2qETOvGi9t4Ik5l8nmS1YyWbpVTKB77pccrh8vavhn1m/X
yUmsXlRnnZgAM5Xq4fdVxlUQl3L4njWl6Yt8Cj9JgLuI3hjatFBLhFSp4foD4D30u76gJUKdkbik
9SnAkJZJpTGQ0OSSy5AxI8dWaLJarBkyEr8Sy/9U+TaOnK2dnTHCKdkFXcHd5EODxnsy6yR9KHdm
B4uXD8IPpKsx4jfuKqY/x3I+iM3CcD/zlxDt6NFKQGI0UiHZ7BnTX32+2HclirPGSIfWuLxM97jE
81iYOn3NlAmesz3QuVHamBdfEkS1R73wZrpf2a1V8oKfq8zcSs85YWZSmQ//04toCLteRxleX439
aa+f6AZ+vF4WfRdu+aC0nz+AaXXRZUOj7IzFcUIuYo1ozKN9nMFTduTzwrYx3KNCsl1V1rgHr5zG
yE6Q6GjiOD9pIlk7cQf1sj2nUGEdiPvYrdFoZXXAFUGK/LgvLr3WA7dC0PWI9BMfpcmYqs0vXki0
4Q3lH+P81uzxDyCK7JBlsXddlZRyapjqVJurJE9h+LCZRodRZAIw7Z928lH20L25fbkyH6lknMkg
2Se6/uZsOdznDCWq/pKRw5X+lcYIrAquQBeXbKMofdeu6m9EuX1HI5yYAUJK5btk3lSE7rGr0Dpy
wk1bedyFu4DcViiJZ+zBxtkZ1shxTG/YiUfJIZVxI3fNq5RIe4MoX8ZkuXmXYnhaL6zjU1hRlRlF
XhStFm3fYg6tDTfvAQcMbLci6VmXrzTJ0VqFqGyQcVwbIITA1nSv7Zajgj3C754MKQjUWUdZR/TC
6FBzDHk4kpJAjDmwcBSd5kUttUdIUfXujaxkOSnkQeR/ZHy/C3LumnCb6Qtv9OkCYJXiCTbdhxSJ
4SR1YaO8HYFf+0mqDhHg9RrEuuK0+Kl/NpVqCbQciEb4GDjy3uOEh4bDyzovVVkkZ5tGx9Nku3oD
PeVSqwiTAz/BRlHYvwSxu+ksQxD8DW+AGfr3IqXI7NNl0XNgJavz4cR6yLO/yWWFpjDFRF4eyi4K
0d1DpZYudDFF3Oryai19RI52G/V7rwS6lBgPHnpCqcaKPlXqWTqBWJcly8EbYJvZb51jdgmtpupT
PlMpbt+pbs33OFsro6Ihlx1f4QEgJMK5q/tPAbXadGLFtaWwK73JUnm82vW7uPNAhZbPcbIbgH0H
e+K16Iteoqb566lbZwEPw2yLR8Y+K3NcTc5pWp4zl2tPVcBHCecKHPpu7cYSNORjapBockbUJbAz
VNtKFSXCXUUm8ksac2DXEaKvJAHBv8mhodILK4sNsu1co8UGsbJXtgJTzrxdISk6wuYm8buVV1KF
dmgacJ47921cBYwQYzRW/Y20W144gsOvC1ByGRVQwZyppxGafSHbclSDg5kncouN062htmMKwSLZ
e7zHbsQC3paehx/EF9cJdGaEm6e8s+3xQSk4pNIvHAtDktDZghyTmsasBijwAcxWAfNplbrJGSmW
3DdEx6IUNP1IoJNAJV6yuC/1ykcJo+PVTzhNy/DlH18ujMCbPqYD6WlvD00l57inAw/mrps6ev8U
4UE4oV74ZbJ+BA9RNJkUmy2SSj4/a6LZecJ8D929s04imVDxcQ6DY3MzGkGhhmpcoW1FzQseMJDS
x+lKIqPqapp46x27EyerABJPKtC2hX8i1TKr6U3WhXrI9xAHpnp8rVzjbvHbdeK2NUF4iKbNGL/x
x4CQtjb+/n49EBftE1A3rUpPQ5UKtigYT0icXiSiHjlridL0+xrcj3EajZXN7rDHevzjMfCJUgAQ
tZ+RMp2lRW3IL4B3bJO9HJFTNkJLoSS+UzeSdsmlwygIa+a/3XZVPKvRNuQaFrBU35BR2J3qOM+l
uRVRw/OSo8Eh4hguEL0+HlUJw+givdhhCkn/g+ffeWgOcfYN3Pu4UPeO/lp9k8tmuEzdM+3NWCnA
m3S41qyiAcsZJaOe4P+7bFGBnJ8T9UBLg8ef1NfwDbZtznNVq0jam6Rl5fyjOsA7Wh7rz2waoTlc
1Lg8+dWDRWO+jMzG5aGhyIq31e+nUoZ6UvO0Cic6j/t4PVhOGgUUTqGVhZ0NJ1+GI7ckDyaXYmSD
MRThX75OtHc9wHoOJZE59k0xiPPz7IYcs8xyx4nIkoU+i8xbkxjNzTFSfwKyXMinscK3SelrvdjL
Tl1INMqSPWwoCU1x12wPsxtv7fLMO7upB7RSen2ggUWZtvAo7xoo//DjJ61yRtm+bWdGhzVvLbW+
2IpoAvUq0OlE5fouyqrkuxNYABMX9NXn0KQN0aPNyL+wsVoX8af8FX0zuCHkr3FkSK33S+TpL+Kb
xaTk5mnq6mv45Nja/jpK8WQoLiNKb6lr4wsm8Z9EkOsrcvOylyDjMRPEYRlcEKSCRANKcdRiKvVL
jdydUEYiepaeBvvQDtRN5VUzl3L4P+3Z6qLqDhRORTXiq26foM/EVnqo3h/9etUURp7cvilLP+Sh
rxdjcWyMI4YhX9WLeAUgcqPevMQKunUVM3TP48lv9QTPN4wnJGVBTbh9tRGiAh109FxRvMLFHKDU
dP73SOamJm6I+PeDsv74BlMEhhN8njdxuM1ItArorUbrjALxzpELFdANR2Jpxr7KR11/9N/ufynA
r0RM7GQd6q98Q3XNmzI/8X+U/UniMarA6aJI3Y7sR1qYqBXguZQICS+BCznug5HybcESCD+12iOv
XEwQidZoCMy0DeCXatbJvCrQcWI9e1V3HoX2OHaDuNq2fnPuQ+FfFvC3lSQt/f+qOxO3nSPw8VJK
clikL6WSOaBkgNpcqA10G2yQPh6AI3n9bFzFFkQV2Whvbo7Ff1e1hKEgdiDmHOvUhgZTlw3aZQ4R
XAW3Z8GMzPD9r6oCCEzvGrozHXAcqOxkTyKEhPbm8GEXYOujOPkd5D/Ieg6hzDre9qZfMHZNGzyN
9iWFAVIdX1H3lp3OdWglkQjtyzwfZTgTzBqOtMzM0Vi/YdnxSMdE1APK3U7kMDLRSnTD56K16xoq
O1CJEMAUW3gYC7FZrC9CmNnCnu/OSQdw1XjeNFUJ9Q3op5MzTvoNwmexB/UHe7qVIDaziP9EhO5R
S3MfsUGBM5puH8MHqQByH4YkX4S3yhCZviCIDVh5CG4dG48DeS6v1Qqez870G4/PKnqD1M6KYKwZ
jaOnmdhJUw0KVdFnw5hDfa+ErIYdQ+zlPoLJEnfz0lyL3eQJSzwgKOQm+q888Z8ug0A339UIfgG0
pm9rXPrxW8qrE8lEPQlfL/cG6jMo5a6oJRegwxcwWWeslf5OFlFTqHz5l3RDQju9maqSN6QOWH1w
qMbvM5eD75+tc/UOAje+9eNsizrcNzmx0VBLhLd5wyfUy1KtEfIcO8Q74/vGJ2PMY7sgR/KefSNG
NhYj99mB8a3+pLvIp4ZhjDeab2loBQsyDmGziJ4/AxeLs/cD8N+0CCPGAH4BpTXfrtQzHcZNxdxv
1xnwX2pJUwOO3Yi0uqf3D5RtOMumAgAoawWNer/hrG3iCZ6qJHFA2uxjprAzsLpW6AUEfcz6Hi9q
GyRTVGbH9fOuSdQqhWkWhJjBziilaqDmjCAECQPP/ZslwtTEyJLQaUx+C3gXZ4GGRfBxx5cXnfMi
DZ8vNHXE0ot1Yk+GPaXmZAp3lB1TmxXzHGAj6O2G+bIEKTX9JNeCyrYdVGosSAbJGeNUesHsPVId
BC7ny8J5wi4rr82lDP0nQkZ39LnD4WNdq+q72odj8MO9OhCT7LJ2MeFBV6WzRAZtR/h9sjb7do+A
DGlzeyMyWA7PtrAvjYwPuVxR+UXzjG2fWUL+r9OM9mk/iEKJu2BO8wQtqMSXOyh7zcIvyrfmqu3Y
JKF/ZDg+elrB8+uf9TEQMCBLvpWzj7nLo9CC7qaBGlUtbzxlYKjE3jQegf/MuPDGRUpXlI7yefvV
RayKP2HN62/VKq79bA93ljaoMMGc9oEcxzBY4+ZefiJlXFAMRqylINYfUCr1AMz4uEZPrpvffKoO
AIDLUGc6e+SS2XkKvHna02BdTqOam40rlsuclnrI2Inm4M1eiTfxM9p6zKX4zW1L+JFi8HeeDV6b
0nMXbSGVp46efoB3cPeuRcnrgcbUIzw2yoYPUj/gYHfregRAbDl90oi8eFSbPwo1gPodp/rJ/VsI
8DKgJ1H456fHFPGwhFrHyIATlc/tkN9SyoySbak4XbHStsn40mUvwJhPVRqBPkHDUZtbI3n+/ZdG
haBzdljA8kdPwI8duk3SBO/IN2Xhb+L5Wvluf+ZuMjGgMtxtgHYKVzVMA1gK3mmUUGwlT1eXDGnp
vRpGqyYlNHqbZbXcXta+rKOqFPsOmlCirVbKad8vct0D02HU00fsL52qjWOqqqAVH+gCXaAi0jaU
WkeRGzgLuR8CQe5izsnohFs545l7ezycw/0j56oFkiGcUb8iQOTd/qlxa7QLUqTR0wkVmihfVp8b
CyVTpgIk0EN9LgnkemLEeN3+9dlxpw3wYow1QwHnqmBjz3wGlJs9COqZwkSF+RskY7zxV2ZuKPyS
cbNgPePABIMbrt0T/f5otFFX0jEjOjpkdUdirZAKdeQnp33MNq4UwvixPkN6UJWBXv5co8XZmVu0
vOCw8t9zlTD3csdW97ILSoBZ8fPVt3561ZasNa1nQWBV17NP57/Jsr4vs23H8SEr1ezRLa1DWXb4
wjQYzv0mizyFWdShtWI/6ol354fIN2IuYVfRhFDIdA2Zd45YY8E5PMKiZ4TNm6IbStmLv2NZVqOW
OQofgJlaemFdqehhYmpRnG7k5ggeWw3OWH6I9X1vfD5AaL5q5yhMFVsWtIaurpGrz47E/i0P37k1
T5IKUceTJkTAO7kNXydUesXCcDBuM1KQpUbPZjJapl+rPbBa7UGaPFaV7B+AusoVqjlNLsqIHKFz
pEjC2ci7v2FcwmT98r19x8Gs6ZWmNJYNHpYI+v4TZeY0cQxu+hcGejRu1Kf2ck/8wXbUQ+dTDeOa
E5lPKxenVvxz+ttiCoPNl1Up2EWYlwnVgsGl2Yaqi8WJCD677kaIXR7xBHVRldYzGY84mzWdSmng
1FgHtAKRx3uAX6jY5KrfJ4+FiPL7Z7dfLA3qDQdwj4O06c6iTdfcuzXUtzgYnBSuzrZxnwgBLj4e
wzrJbhhYs9CcQuq68ryruPiAF/pqkuX5JvpDmVNTnMPFwkW6OuqUp9GmWZ3oUabIRP4cHvi1gZU+
DokCB09qn+P48Sv3nXYpm2/lW7KbdnXOkRWbgKOHF11EIS5vma/3a+rpSjRmHuBabLq1UvSVmdT9
vrfibxhnOncqT/tHIM3YRtrU0kj8LT691KKdDF3MpOilPj9aZlSZczp1wOKCc0HZ3tqaG+hAo9MQ
QLd7iFCJCclPhfYIf8o6wyg9Y8G2BOpcD9y07Ztoa+n9jW7DlwG+/Ek3CUQMqwVdZCDyqAENxPT/
WbH76/M1jlYNxkoHFcm/67kS0zp1JQo6KiyaXJrL08sAQtkHL5C3cmBxK5OzVQLiiUGKGm9PW2mn
NrmkynxJA/QqaqTTUruKJanSQfaIWtT9gemBOehBQWICZS3hlsPvWjiHCvXx+42ah7E5P3sopobp
LNx1TZ1xhYqNapvMTPEebDAojY58bGWRvUollxTuEiBa/qIZX3atwg+yDOPhVg0rvNCq4+RhX13X
eeTIxKP+xmL/g4rFKtl1/g8iSapSIsmvlt9cyG2068i8MdbRBWO9GNOMWhK3XV6fhWB4w/3dUHZJ
YUAV174OU2ioxdQGq0xljCXxiJa6WOLzkjcqyChMRTldkEvkHQ75XwQLumr7e70Mx/sAkZpyFoZT
gwUgpgBFHJS5YhkT9KsrKP5ByTKd6zWAQL04q//Frxx1i41kbYtvnDQczGH2kaWPB04rBjvl0idN
bIEwS3bv0UOMqbGzYXKDAMuxUzriK3159BN2kd5Q4sZZorio376Mr8QO0nVoITDnGrD3drLAc85S
pS/vW9jiFH7Gm/M0E5AeHQw4DLp6CsO58H/Lwir8pfRUNO5Qex62BkrF3FbqkJI3ilsrprCt01HU
tumHmBqbrW+aIhNpdnFyt/AZH7Gn8Bh+0SWtwlhuy0ifsFPJt7ACeEJTP4vUWgmVEbG22eHH4XO+
I8nqDlHPZLcW6gGLwzEhSxI4Pxh+BREuMBEKJOz6RDZa9D/iLL9YvaZLljrN2nXlbxFuMSOwnGFB
lprbyOogrjJ+X1bGrPKktVOCrEEti3ahyUiiiCIAjS8gsQjC2n2spPjp/KiZRMlMqsqeIHqkHhw9
jWKdj86aqKtHotMgkKQh5kXSi0opYTLJF5+5D9338kQYoBpg4BGCKzNbkOr6FRcHKTrpPyPYRfYx
E+vL1DgFVy6eZeVi2k0xLeY9uSLYu8UKWKl7rol6fHCtQeGFfuVC0yG2YjkQRvmGHiW+mjzE095S
yiWDPEGB7y768yTbIHRdw3/aGy87eOC0uT3TSYE5Jme8e32P27rcVMRrBVJL3Iywg79QazfgaSdn
qZNd5EAty6PM4jEA45OTdzEguXlo/+aB/RhRIDmrvd0sc2GKhbis4fvvj0sa1U0VWsxvanBd3ZGA
mIwAdfX8WICn3Bm60cvXGFz96cspVdvUOHfgo6r94P1xoCZ0aadXquAZKF56hylhNCN0pq0bbeQd
CjR0ST3jQsMETcMLoVNhzpaK8NGh8SWZxk2xMeXfzpHFl9Y3nbJ3LG2Fnj/vsHvzayYejgtrBYdY
kF4RSOjTWSZM0sdWyMNc23h+X6TL8PA2EpfopU7Di0cda+vyHRgPqR2ynVrrvIfD4rqiZzZZu2hJ
7DRncthdwpjKu9wHvoxwjRnIap1GgvMePNqY8klxGQTlNOeztCiP7gSO2oH+43XDCdIQSxUxfNxb
9Jav6ApeAIpWHy4cdrtwYA50eDRQhROrseh91FwTK3f/qXFqO9yEuQaBML/oZG4wg8EBO+/E680+
IYtgmMpwFIy7UqnJ++nIYUii1q2ctLan+dkBv4l25osgCANPbJtYIyvHJ1Ag4xSBXRYinaTNd0fm
xGNw2WJmDllNImAKDv64yGRhtvYpO4mriCQK+pGydlcPNeqAhCI0OdaJOM7FdAWH6Z6iHwDcU75I
nY7Ix+ixQH1v3E324FUtbNHKuVkzsScDsAg2WurOoQtmoPnA2vr/5Lj9HKHqG8ZrGnDK5IOdJVF0
oJvysR6/IFsbZkGFFdoXdpzzUWKlnfPhg3cqZ7/4rtY2akh/C+RM7zUnlD7FZJ7UxBQBLzWabNsT
AjytqBmTr/y2yHnjfSG77irdhJxG+v3MQfUU3q59KX1Uk/HfR6qlIaos9TqEHBUv4spsBv4dnOLt
lnVtINeJeoOSpUEpQINsIsdpfhwzN3pp3uHI+tuEFKCy1/zl2g7bMoS3zP575rzA3I1p9pPZIF0j
FUyOP0lrV4tY0GtICGIg57bclhidYWYF7ehFRGWVHsJO5RCqSnLYnRRzmxC5eAth+X/YHujU4stU
n5Qq08LqevYeiaq7F9XQKavBTFILiXGDM8t5riF5uDO4haDumAaOWbfLTWYg9zhDHFUD60yGS9jD
unml5wpGYhnwLPMqzZryN3/KN2yURE/1TVolR6nqG9DxMkfPKzTIyiHmk9r+VYNWjqKEVfmw20W/
FpG9XLkdulb6NKWG1AB6PuYAjWUq1wIwGlaKA1ow1n6wVYTvVmVUNyM6631ESCAZSREnz76O9cnu
pD1m1ScOhNKYeilBo+lUQqzT8EwM0wbjOrciqAk9aUSihWRuv76qs91OT4EJTXCVcJ2/KI2yomJb
tlNh2AoKlzsfYR9Abs1HWFiDUtqudBhL6Jh8ph2VElOEJqDSxakvubvO8D8CipPGTOyAZyfesgTH
cOpkl7uWf3VvFS813q9D0QweWkWwJ/iTuhoxI68nrSwknk61oW+7bz9iG9R5AhIhA+O3t6EHX4E/
iU/Qy0HiJ0F3nWrDQfXe12jCLNbjvb3+/s5atPPGe/enYmxEmpMaVvGzCo53XR3zPQnhBgUAf4dQ
AjtRR2iLouQsCZYl6L5UtuwVakZ9ufwcYO8dp0MHGocRunchcgxgdzpdc/bkC8D9cqCLQd5bomNy
XMqHmqW8dBu5AkjPpAkkaOBaPBrPGl5ihvRStoRkCvxXgGm5nVVysxCdclBEnOnbzfACjojNoqGt
iVtAF4YBDTw5Cx0JWj/Zrwfos8mclbkX7pFvnvbpPZh+X05qaeJC3t2iJkbZKieX2oPzWep5vTUF
4uqfCwRwaCh/J0je0GQux9EwzlSbRnv8Srd38pMGj2XfJcZVkbjFSaPZburipEklU2RNQuHkyctD
6+OsWojLljISar62kVapeChZaRk6rQ56DZzymZBmkgwy1t8R4TgSqhJfqyWLVLNPBNSzAKcEtitM
P4epyqTHg3XOYDsVMXA6zeUavNH38mYxEbC1SqC1jRbp++C5Zjrj2mUKyRDxbttMO18V+LIHaBQ0
dgXi0dg5br8Ap+bvSm0TmcrgZQ4q00tdxF4mttpm9pZriO7EA7lsFvB/x+31qVEOCW7QlF5mHzVJ
vEbaodEnCfYqu1cWaU7DEHXNDlXRAWAgLoqATSEUzFE54f9DCDKLm/B/fwykwpoergmsV45zuhNB
OPGre1WZ95TLTVLNhQHNnry+0qpDe3eo9xFPc5gAfBC3kJWl4FUyze0EMz2q2XlyrBLwAyqBCVQ9
YE2PPYu1rbG5ptMQVi3MP02LUU7kXrmPlCM6SW5+VjCKvLiHTAlB7YHyDImHFXPoWgS9OVqVdvb2
UOaVA4XgReHjt0t2S/vNn+G3I9adD9FtITehzpqN4xPZ0rDQEqGvsE56Pkj2aRZf6zOwdBpQVY90
/28WxIuCunl0IAtPbwlLE6QEqBEopNxWjN4UKYB3ealJPJhqtPFfdeGrYEY9BOLQhaM0Y0QNglZC
DxH/qUmjQk/Nrf+ERzDagUBeB0J5d85AFzCSTTMmXvIkSbPgcI5eMmYUBfPpaONSWSYvX4u2HYVu
DUtT1h1ZVuSR89G3li9iMl8AXNec9UtvYi4rHy4lFokeApGw7hE4oghsePgdbI/syQ/nEoArvSb0
3DomIauUfboWIu5xlGNZaOzO2mETRSpR4PvQcOQ2qTqwyX0iWochlNE/gbBVcXuE3Hfr8O9ThISh
oLxoaen7Rrb+fU0kKZchlRA2kwUhKHi6yI7toksv1NRvldG4WGepy1emv+8fQidutIe4HbHXNhkb
pwWRHNAJ2L3rhDmlKaySIK/uFECZkNPZcJ7+cz2cja9Ard2RnWjGhUB+os5oiJrX/bGCBPYQNnO1
G9dqsAtU9SeiCAlTxpPrruQIvzUQfbHTZ59pT+SSgtQ72lbO0K2pUz3RR5VJI4decn8S/4EPHRlQ
z+125Um4TOi6bhNRqtlNELiec/6RL1Ery3QHX3FfnN2JnEJuQHJ0eutKKZvEBJoie0DCRCIzfd+u
yQZkC/vcKF8xYgXAkHXYYL4/gYyji95J+bxGuzVDvw2iWXUYKwnb2WnBbNp6sg/Os1EiBKomQOHC
cNEuWkpwkBuDvAkWSdfdoRBna+FR1OsZHuXq28h9Uqer8D+Y63AzfW87K0rRXG55pNoU7zMt96vH
W1/+ObIYM0GsyEFf1liYSqPIDD5t4xU4ZZy9l3NpbkIC7fyQZQry1KOkB1eVoIuiO6n2kS87oCdk
ItjQN9MDlSthGPVCJpf1Lw/bCcwM7So9FA7BLNUFJcIhqIqdfIb43l+IJrtpEj6oSM2miMu7PhJJ
boFzzPmH2/kupW3o6Om+Pj6MFg9AfvlyXVFJ+UGcDUZqxP6EGY0/9iCacNV5Y2HsfYAtjEn6bhQV
Gdt+NK8ZwxrJoNv8JA64p+oZxhug705FuKQWYUZkokVqDGKBcA0DnyYpOiozY9kP3lIPDnarqb3j
rUp/mvJApnXQUcJzEIHkcEJqyG5Uo6h6IjXEIf1ccM0VxqVmpaE+GVlYM9CntaG4jqgHzIeuocJQ
b0su5iWOZA2nVwkLiq/pOBey15CqGg+GKbQIwlopvF8LixRH0ULCv92B67aNk8DLZS+kPhACdfjj
w9Wz2v+HMNZvVlMZQtUOOZ0o3HTQtcQs1KpnilnwRUMAHm2bm4M9YxJZMr9JZqHgSrW12uaGdsBu
56dD5Fml8EmPr1EtqSJO5ArbDvKa7bZftj4+BUVakP4UlnqMeHgpAXNF9QtbrZ1eJtiWZ0ycRczi
dJ8vRKNNHgzinXjWVf87+gj6o/20BqUOF5mT6MajqbzJDXyNPQfxAWdE1Mcirbd52Gm9b9nr1Qnf
eiOW1OsltX8KyqbGCVFNsmR0jv//ayB63rqbvH4thX0TgQwrWpVL8SRGDxqTXiVM4YS1A8zKgemp
cOSYMTDobPcCv7T3QfLd6mYc/nJN2u2c7WkcKaR/8zCviDJCG5qjGv5GL12zh8yeo3+2G8jVCoSu
l/q/T7gOv7qpZ0lBY1SNpAsowXwlijHEmPySWemwZek6pyJJzBLx1ufuGN9XE50UEK+o7EYWss1f
kJa7CtRLdSMJEZ0i/Q273+h91KIqAnHYHz/R3qb3J0Q0NpFhcklaMEBgo5RTrHv6cg/smh9biTTE
WtWfp8YZM9BL5JyJbB+sNan0fmFcB+o114p+O0mvOAPpQ4xezIUHLf73DHF/CZvIvCdK1z2T8qAr
mVH4gZ+UYYGO5K/xnJmk7OXpgoHrOn8YhOz+bEFqt9xkwHUWyGSsCX9ZVQrBV0gK3ewODq8pbr4s
zGEgO1DNeKbz/jJFfvOxjJjFXcL3ydoLVfzfK+VNDpbsxEEl7olsV3F3dtelu1myrpoPio1WiUoY
B7X5t9VrnITvEMEK8k93SHknpPxDy7yuUX6Rt63oKx7LHebq14b8uyIa/QjpC+GM4VejlKjg/hxr
hGUtGNNpdptGjvxEkgTYCOmLFlbvBbktgsxIWbEYSh5oopSfelpJN8fah1m7cY/sSQmxznocfXB4
gA7HwQ1EN06J8KpYr9rGAJzNJP6399C9oMvEpyD2hdFEGuWdTlOqeVzB1Fz0gPIfgGPrnJp1a0E4
bLCqW4OWgS48SQLRupdCtCVTAh1ptCRpCGKINHaHTR9YmBq067++IlmJa0ve2FV9NTOut18B09hK
zgUe2ROW4k4qgGY62XeLTZ4mUvFME5ew8947TJfxD6FeSmbZdsPLeiH9dokvkdO2e7h9fAwLPb/E
uZY9WRmsxc5H3ly8HnSdkQpF9tWn0dIgYqkj+XfnDhAKLO+hhrSUgEliR8xLQDjYhbYcnhrR5oPR
bq4zN1/qF1d/+nmOJlcRYHxiHjkXpMOo4Rnmb6zd+XDJMkhE5Kii/zRrWUEC0pZlVpD6LazVzNkl
GSfFBGhnF9/hu1mwHDtD0DNQh5jjmLbPfj6CCxMZE33uKuUyUn6HrCZUXOpyYaw3dD8mMF4tZ+Eg
5YcJHa6vlXz60p5E6bBW22OkSfCvr43AO/SRXGYZgRxgSM10cT27wGWTWF6/p7kCxFudpHD4w/9c
RbWyjwN9aYi9sp/NlWMsueoEWJq4pDaBE9QB1PAAsoVs8D+rlu112MOzu/ptxL09AG1GyhUgbm35
c+8lP83YU01SxuTvBk4Z2hYoqq6JR2cgXLM5HBTronYotWpVo2uh2qBIJr1xKJkJhfZNpJm5Bd8y
UayzX5s6dgrZy28ZEjijgUF4jzW7ti/SknlfjPysAusufUx5eCekENFUZWzky457LpgvNEoR8IiK
ED0m+7QO083jRUxhp5LBjSXN2d9pKhGZ1U+CrDNKoJgLgYmxl6QWY8Xc1hQctDUvehmp+AvPnSYc
4GMYURWGOP+cQaRIt6r/DaJLpeYN7Pv07dAfgR9N9QJZdBmriBY2XS/endTcs2Qf3GH6hLylMa9t
fTTvC1t9yTQ1Cz5V5fwe0qVydSp+PKlPyTLBZckSHvgiK2kz+tXtRo2tC1SuhAv+APH/sKEFMbyb
8JCmWWYIkQgVP6r+gup1jB+GkQBuJtRz8QtGambzsZJZlj1FfrqcaqyDSH5x5opFt4ZQbEZrv1Qh
4K2ycq1ZxRvYSUwWxVKRbjn7u8qqjx55YgK5DuZRPJWknQww0mdbIQcjdlD0l5qbeUwxEh3M563e
t88pu7KN2wrPNpelq6KU8GzmtNAgZkBHccOablOtS6gMzIRPpcjXUJfP9/aViiIUuvwFZ8PS1rJk
fIY9+LxoTQzvc/T1XDfG/9Gazfd2F515YXeQjtfxOG23oSniMRC+go7UyK56tWzPj7QMtIDI8Cgd
bMLnn/AzK2Kvnk8Y6G0z/x4HX0FnVaxsCOSh1yB/BkSkFVMPqumg4+DFpkChkIVYDqclbpXi3wTU
3m70P7+C1PeZ5DzNzg260lFKbCMO56iaEqIY3yTc+SQFUGhuhsYr96ASNol0uFcpPw682hh86Ut8
LfKmh6JUUEOVBsuez3qH9Fmy1kzvK5kBZcqfr+wuAjczShU3WNRr/TL1mNwQjYE1JjoDbMCT5yTS
nR9BP9/Fop4BXuGYOrdgiwFqsVrYrdwamI63VCa+DOjIILgvK1ZyyXI3fWfSFtVaD+jV+O629w7q
GJHYrU142YC1UsO6MOaNm1C/uO6VH2pAqxs3A9WXijxgxY1SiyzcS2UqymIyU9p3X7P3ff1njE6R
s/OD+4iEIHbTxE/n5PbrfVz1PdaCry14kAuJNNWCMwkB7T/exH3BSC0PNpOaTS4U68Vw7GZucjAp
4ylAz8p2mBSW0XdMdzoJ+Be2H3u6QLUuNVFW2H5IZMm20trHx6Wadh3WyYdNfyR4jmtUOaxY4hp2
Snree5/kB8wKk4C6jmQORcTK6M+6pHY+qTHEeXgZv7p5fBjDUBTAY4zyuZAeb7KGoeJl9p6zT+W6
f+/oHSIthKAqsUpxOKHVSfIzgbfYV3JvQwWPFcfCfHWtlz1vqDub/mUNfyP5QfSyinTjLTePKEUQ
rJ70eAxgsiAKg/prqmw7MJkOQN09t0prJIStFmMgevoLcUloSp7MPc5voowkTXea7WzHqIrQu+0g
kedu0Dx0qRcm5noSJspHSmOTzX09Oz031zf7pf74PBMGIVNz7IC8fJgnMekgudsIcu9wSXokHWIl
+odR0OXT9L3ad6E7ekZLuFOWLYjMx91a4MKAuwM6hfuQX+GX85D+JM9N5TgOjNuwLcwW7RXZ0/T7
5u9OCx9cvphpIuRUg47TVrWFhjIMw0I46kSUbDOLJ0lMkEzu+APKVNN8OzN3TZhy6iDicNlQhWBv
FLWguAisjz4v1E5X6Lhd2+jcm9JXPLOJB1Qdt8fa/GJqtmh/fG6LeJazzw82ipuQudBkZMPQssLV
w8fvHJif0xM2pl8OTjhySsjGxGUPeMFQ2K8voBaUnnzrd8FEgWIlg4gbGo6CndlAE8Iqnbs6igwK
EbUsioAGnmiTasmGBAbsIOv0QdjYQ5rQhX1ZfJ2sv5cthcFmuIpIQAvmK24hWC7xT5P2MxhrnUjb
qGID49Ntzlb27e50IVsP66QbI0OorLQhWfPBi5UQOkA1EjqVC4hSUeAhkVEvRGwwEVeMfsrGDnyP
ey2q2FO4Uu4tR97zTh2GYVVAbPwOsa5QDA8dZblzZ+8JWYzr7BtTFnkP5Wu2KDcVDRW9JEdak+ir
+N6HMx2b/mfBWIMaES6y9Mk734eyRa5Myf3SDqs431u/hLjQDP3VscZiROBOjiJmk/aD4gwu0Klt
8HJ2mcZMArZpr8nac65BdsaKsLM6wv4LySlUwjPw3MD4DE41iin9Cf+1SrHeXTgfx5sKy4dHv4/k
gY9GTe76Bv7cz6TyYImeBJ9kaiZ0PxrcVeULnMqTMtz0ANdpHRF5Jlpaod/6AAVpULRn5KZp2zSn
BbVp4MK/hDJb0Q8K9zcqX7FiDThPl7snnYQiM6Db+FoavzxiI2+AaGRrEetQDg+7No+ZINXgJH1O
1/A57nxbamWb8Tp1M0nGnalW9OJJhEBMR+5c+eFgrwzzaY+bb9rbOloM4rcM/nI97cyWBZiv4En6
eC3hollC3jqNRPEgyNc4x+GmLD45oHleK0HRKkkq9d17X7k8+YjnScdgox4vNEtzw25toT140Ugc
df/Bg2OKwt61Rsht3fyIdFNDQrAiR1Lt0yOJDvRt/aYOJobs4Y1w1qZkWYxmz+NdixpQsiqeWuAe
8qUtmnnxgHCLX8uC0nwb2+uT6kC2SPWlgm8eXcpAX2dMoGHTffbyqc0VJxleF29CzcmSeqQl/6ON
Mws1nPB9ST+hWCUmD+jWG8XUE4IeWJSm8EVM3buJBwO1XJnaHiUiPWlNQS3CWlvINrDjxZRKyxyh
LWVLk1x16fN+HUuArE//Lc9b/VKrx/nR3b9sN97lAjIyKZKKdHIAC6rMKlAOs5CPUdLZOm3w5/oj
ZKGpAfM4TUNPCrswRFkFNPyWIx3+4QrAzqxJOwejPn8rTPe8xI+HMG8dyy917th/pxAB8nitDs25
SB3PRi/euP+0snmU2pcnd4WebJatwFZZmITbBWH5U5L+K1rEnc8YnhdUy2+yS1p/USskvKv3xEJO
4kFvrYVhtOBmNLXW61NGWvTStMTAgfTEC5/AA8Fh/bgvXCQStT1PY133TU5OOo5NoPPp34eU+bwO
rLQqd9RAU4WvKvvaBj3Yelu02LLnIrHZblSH8lDmbF1vlxsqwlbmQKEGBfZEarvJT4k7xb0ZTUXv
DqcId58pNsyXsnRM+nhP45aGLTL7hFU8quYRGAqiAh1+/FmAXjhwx+SmWNvFr1Qoon6SkganQn/Y
L4jPFWMfKAffl7eK9cQS7i/K4uFh3Qyu/Kpu4OVniom1Q4Iz3NkqYnZ9SUiMqUqC+tzLcuDalZWt
8EOtXycIhyBmW8fl6pMYfapnyeRoCU8eHNh/gXBGY4Ze1RKjqBCTvL9s6lDGCP8UPpJLS+2vpry4
Qqo46R11i9wrCWv/NHMry9O2GnrwBSmuwB0BMIPK0G1AU6LH0kFgkoOuEgxoAniUSP4WrUvStIM2
Mt04Dulb0i1skHNUz4VMBK/bMtdHBd0fhHLNpy+5TOQ3PB39MQo8E1PcduGU7mRnAFwbacNltFOV
J1v8TOFzrJwwntWc8VNR0jVoi74+WzB0a/X+qrq8rZhCjvuRbVGWfp8mJwAFNERfb6U3+ZfzXFP3
WYQWhuDQpBa+sE48XLiDU34fJB5l3KBgq8y8MW8Zqlkjcsf/sD6qB1TfTWYxBbsPpbwZpb2qRMdt
YSueZMkAIn5jlJ9h4tSfiFO02ZkBOpu2Ha6+1lJ1bu/4OXvg+uQlIVdLCNBxSrg4/+3ueYLy00Kr
X5DJfQveziMwsr43GX3ULnIXuv0LBjF6f7fXChk6gDtUQ4wOxkOnhNTMcslyqKg1PEnow3tl7FDZ
aKR9UgDXs+0hGjYKOQlTgXFu8LH0onR4qlv5FngpomInS5x/PvHaFYjOaclQjIHTcGVFt+NyBmun
QaMuPX5OZYeSSxz9Xi4Jzc/FbqHA+oKozz3xk9NRRRiqrJzbFtKlwiNpC+UZLX14JUNy/uN1pTVE
vngBEQ/3I+uqS8dU0dKWkX2rhxH8GCjxfLZEqWKiaEBVkxXWMG05GhqSmtKuYw7TDkc3n+8vP1vG
J0FFtFtSsBgfmbp7q4v6agZWZ74zrhxkk3gSjG3teUFs/SaZ3ynHdTEBpUjbYorFQBjWm2WAWsqZ
zxmgOkGArBuKeAixkL3CohxFU3jTz2YRpFnTRcm9ixsLi8nXUIUITF61ah9iFOj6oQPCd+4I2f+u
cJNH/ann1wLVaZyZ3Yca9G86QCsstYXs+yNBhkmjCZ4XEBGvC6qdYfvpD24O1M0nYMY0ndDsLZas
GsP7+2WbOfu1mAexCBKFDmbYNEzTKUSYYIbnEm/cw5veDhBNBa2MO8cKhoiZKb0knG1ebpNJfdX7
mUjS5hNyVHkOvlIrOtZlCws9qkbPUYMJU2YAyYS/Ib2yUwGArbH323mVWuZ9NHzMS5zop5vnSBZN
KccifrCbmokWUrq0DnfBsBNW9yfV5Sgt/2vGyT3ppWbqYmkpyi/2bziS8ig8jI/GdkLWVGx49iZa
+AE4IE+9vAW/lc9kjpi00XvEhYz2iBovYTb28Rtp9nNz53B0UPqknzHpzSobez2+BJVt2nCalQSH
eLfnlUMqMd4uklTDvIDPOuEVS7ljSoBDhlOAD7KTu+INzc9DXbR8SjHVG7+YizJLr9oqdGGWcJtW
BceLWSfjqDttI/qGGaWV+5Vj+2kGJFwBIuVzI0f9uHBPqAYNQTuoB1k+XV9Dcc2LFDNqh5FcxThk
NxmVW/Bv1C++ayOFVgFcwybKp4PM2G4vPwcLGyfFbhUty9SUGWStGVeQRh26G1Y3kuO/VYl4Glw0
fyb3fYq41SKvw9zFpM0cPqEkf2+aUzP0KYM054lNa0lU/0RGYXsP9lH45S9yrb8u38ujye0DalnR
jfc5u/JFPzO7SEx2NDPrDYCbkqwuvI5UQ2kCuZI6Qmeg76boubFKojniDS6Zl52hpzhuRyjHEUKN
0tk0kQ5m103Xx6iNA4ciQZQ+7I1ud9HmpGzSeAwQq50WlrGMc4liDez0McLeDb8rFra7L99ODeZ0
kwwkyCowg30pya9UYiq9i21SSzB/R8CoJIVa4uqmgk5xLhgVcwB+k2K1Cv7hT+uNVIeW+wvJFyw3
bT5Wxlp1cl3Rp3bazHyO0QX0nPybXzHjCRLrOK5Eh9DfUS4hdOAiHcvEI0yNIWfgM/vLXBpUIq2j
vMv8DdtL0QD7rZIwit3yYOF0Mgor2IEh4tDDGvyxqKv9aKaSe4xxz5XCPi/1Chs56Su8gOl9ReXz
YsrExKsi7VhDkv1iNcGC+KK13ufp3t2Tu9vZZhFUCF27SY+qsTDwnO5Q0svlcJpMEAoBaq4qtMfm
ptcIqoRelvOtZAt4nKpNfyYPmSfhPmt4uaMTx4zPuTyvxA2hO7JHEBTq+ZjS2e9Qjc39+ujCvqAK
3VjiY6fBzKyojZxISAivZxMH/tCbYaFIBoeShtEn/rWZlpgmACssSYV0V9Mf5fbaECpSXJ0a+rqH
A5bRygZk7bvO02NuC5ZQUOVBTj9ON86V5xzX2/6NX/JAp0gERo1VaPyhtaAHqsMlAuflrnRMCLBx
PifiDVYfgPCRjrmO0AmhzGI/ljVukNUUTF9CNk4iSlKdty8tbw9HOvKppKCwD1x8c5Xhs25L5B2v
7AK9w14fuK1u7ckNhq1osKl6wwHxik8AR4ALskb0JwSWoOmusyshbUqN7jPLeiuIcisRnvJ0bVKV
yMI1/FylGV172DaZnmyJaiNThtKBkDuAzeh2CeGznoIMpKTfCr5woSvAJBc8C04D0GsLibtzuGzL
vSggibIZp+PSOcAoiOpQuLAFkJpyiiX4bGnkKLsEiewLFZvtAFqHXatrmMT256B+MrnUS7+t1qCa
9ar+bVx7gZxPO4xAxXalz449Iemh5EwMg5tbuKeFXKk7NAyYJ3cKQWfIEeFneko2a1EkIKGi624l
yxlaR0sAQnSA4qSEtcQHnPmmReq4adPgx5G7RsscmFUbSBSWt0WYebEFMtAb6DMWekqHURfzlV3k
t/TU2TOQmYYGhIIn0DRhbZjm1AyxyXqHhB+LCmijuiZmcUUyNQtXBDmn6aTMWIrfYmSmrFEX0dF3
74DCkp0h1nsWApQnIAC6FVHdJmDgXb9Gu1iE2W7kPPTIW+9OMcob23Bo/rBjdI34fPDccrFuKdv0
HLCt0pdNBxQaSydfqWzeMkj69mcGzcQ3vqlydIVht56Zy/VgnP/+91eGpnuU3BaXpfC+nkaYrvcV
dPz0bJk+t/f5Bu+cMMWt8sUduwY8IM2rAPqaq93WIZsHRupokVIu64JkHHrUD//y4lzoXJUbT0ok
xa5uLGEfPZ+JjeQ4a6MmFaZrRen/pbKtu8FI2TOWmOgjSUyOUUpm3rvjMb9I700HsZi2Ha3wc7n+
3LVE77MOPCiXuTQ9bELgxTOyjPcyMX5bjmxy4omKuvKctTAssoKBWEuLV3lr+gZyyWNiex0GHlRm
THe98wD/prh6U4BnUCfvPaqp2yfqY92GM/x1DSSJdMFik2z39w2W3L086pPQK3ap2oPFoK820feh
I4baNNCQyhEfwrbZyX2xS8YS8UANn204lvhdeh/U2AbLD8QvElBQKiDltXlZhUQyizpENISyOiGu
IespICr8O3STFQxi4A9IfO233vK12l4ZUViQ3S/b7Mt86nB/PeOjrZ1/lkKXbA3+BXii46YLmsWq
xXzP+hdKvQ4C1LDywXa+FYiE/iYVuCOm8p90Ofhr833BlppXfSLcAUPG7cbPIwD8yedFGnf5QVSs
VJfXosQAind4vSHREzX+Le5tejfbAuaK5dwHHuHXB+pNpPEcRfZj0a1MJsdphtun56rWFkvcCp5i
e3vfx426TRKoo5qVToSb2aGP3KNgO6TTIRcT7Lv+Soi+IfSfsP/tzq6zg6rwofBMan/bR8nvCgg7
gdY4saNCXbH1F9hlZ7lhVBz0ysvxdzB/pOQafxQdnnK7yOX9iXF9HrAEl+pTwAQg2xiuteHMNdJY
eTqEoruB5KHtlBmTejdKhwukLJwwuDEk0Acw8G9Dq/EY3lQw+esrpSvGOJn9rgZUCIFSocH5MfGx
pTLursTL1jd5ZTh6r5lcbWj1xG4v3QnGwiGF7X/D9eueaGX3sHR/OZPVeGJUcmY2N8sAlcm4AbZT
dpgPQXfJRW0AJ9LimeXMthu1bNrd3/BLttETomExUYg0OhmwVZuiIoWavmp08vo1XpijicO+TKV9
j4fOXkuy4yAtD+0U/Oa2o2+kE3GmgvPvWPZluQEuUHRsUqnLSeDds6AlTcYVIo7ldgB9rUFKhY9G
iXi+4p+MYWkzdMWtjwcqmMTiQkK+uU4XZvAsLPSJHX9AiU7aidWwDd+I64GuLjGZMNCCjZ816+s/
uujJpxqihAebd1c0fnEvk4FdmeppGcQnqdmdWDGNThN5cAZyHiNaHL/hoKD2Dnn9RpWgMzDBVpnj
bimJeb8jtjSmAFxntnospSXlLfjheywP91ZsFvKO0y9gHysssJK1CD+DKHW6BvBMR+KqFaSH1Xo7
93tlIhmLY7lgt829tTLpqLECneRTs2ghrDXIiNav9Ya6DqwTsVz1t3E4UxD4tckJ/SiOE9qvbcSW
KnKHXWqYiEksYSfn0RdjiRaI94POOtBnHpuamYbD3y/TjcVwwFZKTgazwRDFEynTwyzDSeBFRU2D
mohQyc+qjKNTTqQ8ur/PiWzkAUrIDfQQr93IzzxYHCA2t6MX4BWSqgsTdDvHhXWU+t/jQuE1LdDe
gsMpYQNovHSw9FjYAwiMW2KqRMB+zujxjJLsN0/Iv5aTUonu+qR0moiP3/CYVrBWK3ggbekS/Mol
toO5HwHxVHgfhPqUQtO1FxwACDdtnaqb4POQCMms0hmz5O7spzm15zic0uiH2G9LO7HXBNeU4vjr
d9w0A2DCG0lfj5FLsHo5OXlwivGBVdVVH96y5y76lRcw6Od4m9GQFnxIuLYLOg2uxnhTiseT112I
71Xu8prDS7RI8Yg9Tu8Cjhfk9RfyIl+s1IrEoYaS9M7I2jzI3utgKfdb8d4yPuXrnjATtB0TunkZ
xSOol3DkrSMl4Gktmzy0n8b1oRwI2AIL3ChlORaTFgKwOsSMMJDTstn1WMaHXxhAlFb24kw/K/71
+QsVEKtifrL7NdDacM4CF/FCEOEA7cK5E6RFnhWYA0OVaqIEa8KsWbKNHFiHtziSkHxBEHrN/jy2
Vr+67FieSMpOHmnxZgWuPrNLz1gJQ3HrZD92xWCmyV7vRzJB0BCG10MYJcKDsL8ouGf0n1pkWsTQ
w+P/Uq4RRnKP5gZL6b/tiMEu7/38s3uKkW23vsW3OKf0cwq3sNV2eSAOXtGr1bfxNQ/Wi2tyzxvH
sv0DQYusnucuPi/O4Uu5Fde2KwIwT66RN0BX+rdIL6pQIrnAIHuPvtpvLQgG3meUuCqzt0FSjlXM
yy/92FZEb9Wie88fwWflfXtTHwUb+a+rfjMQmumrRr80Pu4aNMuyk1NWbAprFpqt5xx2fTxa+jjz
/uTlRHeE2BtSSKFi2PctZKJURBCKThDZ/lD+HGfUIiu9D01u8UQRs98wBZttl27jOEVJhnQf1VDC
WBlG+vCO5Cpb9XA6MYtL7o7KwEPS54IsEIv+05FkcsBnxbDeiLTKTW/2Myigrui2wgYoi3moEMMd
w8QtDp9CIZV7QrGU86RmLZ3wgNxkgO3Qvrp7FWY6buLgKzAMS9HczDOpwYVYIOVmiDXOFDBt5gHO
rSIqco7YHFUL+Ot9CtZftsIgnxEFf/8g+4DF7UfqNJVmXIHgtitDYcYh9hzy0tIuUbBdjt4Z1kd+
3M7zsVtdQosocpXW2tcwz0VySrJ1SXGikABWBeWjSWxgkd0FFOMnJPl51H1J9FiGP3jvoYIe/RW0
lV404ahRtHvEH8UBHcJt/WxRuTiakvv85PdU8iV8xgvG7NnFacfz7MQEV10tEWUmjaT7KT5X6EPr
9IDbnN4Yr8azfzZcAF5WAq4MOm97GzS0HdKLfCyhXzTRhEnX7MTpXYpzynwnZynLbJ9v2ZA0fuL3
/feRNa4MRr17wa4ozBgOmYY+U4Iu1811wJmy1ad1syyWsbfaw1rTE7PnnxmAqfHdv5vGlwdq1IJ0
BUQVygxyKkelwApg41Iz709SEfuNNpvqT2eiqRjn5LRnVawwiq9rUqSyGczL/3bGT42oD8rkGVIS
Qy1ZQRxXiiH94Q+iPOi2Th9mS7fyp+Pha5qfSb33uzJohlrWjeIIu06eoG8iHDYgS35KYY+/SpBA
t8CreZiSWXN9NPjSdTyAdXFPg/6M5uUtYOTwX7eVvwZ9w9szPaxRIbcfiyt/cqCp5XCJVnnIZTsL
yJcAKHbJY7WIDPQmJ6+VOLEzX8hnZ1EPUKcfnM9Exhx9mJBhXbs5A0DN+WuuKM/A6Au60sCeQ3sr
rDLLZCwPQ2TRstnxqKk44KmV5xLdFqdj4BtYC1adj3NaSAqZTgn04eCD7Q/+skfhPSKFNHUErJS4
+WcJyL0WvAnmYqAcV5ncCt7TtAwg1xc8uOiGp2PLObK70BaGGYmsXq1PhyhBNfjzNt30HDRncWMT
xMGRtq7fsvU/0WiVpsWIpOczYQkA0bhPhi/dWIo24VdzXVVunI+IFD2GLnzxNVu7CzJ0e0IYPqfc
03/6vQIJW2sWk6i+hHiTpSU0ND6oZw7ToWx1V7fAsxD+CgS50r2y/Sj8XVBm6rr+pjrllYorvQbB
7zNERtT8nOq+V/H2brxZbJofhJVbTQ61yn5ESqdATNPaB6Th/8VWuJXSJ5WrOYbLRQHWeoxNys/j
EvnrxLOwwHa454XBiWTza1iEuIysMK7wprA/4XhoelDCeWhBWpxksER/KTwnzqGoy38UMtXvjLXE
keZLy8h1r3SLXhuV/IvuXFuh/CgNpl48C56wB97nrE+yZ240Pqi37pC4NS7BjB4udBxb7P8+1EVg
bCyhaafAy0viqSP59rYH4wl3jbNY+IE8Lq82JmaJA65o2qFp8CJ16g9cEqZHOjqIcP1dDc3kuI6t
XFsgDnEZw0W6kWkNUle9UvUPkpp5CP0l9nFCFkeYhA+bqpnCKQUu25BODIaPM7Z3eb2t9Jc2gaPx
3rvlWnSB9a7Q/bJE4/c/B0wZt7/vg6k48bU16jiLL54sE+f7wjPhiU4TMclwaanb+jbH2Xr6QToR
aCCvNEeOvO5cQP/Mvw+Gszg1+gjB1dP0wCJ8Fkz/f3fQnwwi4Wd1PdlxvHgSuwsPujL2bJwQ+kpb
PVmmTUI4ZkAFeckYRHDBerjLhAOwarGEvYxRzmudtsq1v8FqURrXn5Iaf27LhvD7BpKdjaR+WSPD
mjGUz3F6hNQ8sgk2JMfCZos8fe9NuuRTjoENJoHCJZ8xRpQj3tfF2yxMB0w8j7QZBq5DHRxac+ez
sSGbsxLYFZScrQlO6AWyrHDr6eyd/aWeQ1juciU7ohppfgmSFNbcuDvTtbtCUlDbfH5y/2ufGha+
aYcnuwEOeFNiUmJUIGixMk1GbqPOrHy5RiCdkMbzh3Y9iX91vEYr0NLRhopxrAk7FahvZj5lgHR3
QqiZMGlQRdljhufPJmQKoLjrelMYDUsF6frmRdZ3P1uxyV23rIJs/KgYbibV6aRVoU1CuzOyH7Ux
O3pp5+xZXDwqtyHYXwjbH0gw6DNh1tnPKBe4p4oX4i0l3KjY3vGO4+OcrJLBxCxILF0vSqwvOszV
Ef+6HsMPDtPF96nbiI1eGpvw03pvZWLj2PjsyUK7KNTJ2ws/HncetWDxVVTCHhReA2+OOR+ldNYL
Z03JBPIyzZdymBQv9X/dc90qL80VlbAtoL+nyFHwZLei4MZo9g4uLJqkT0/+oSz/3UffMneghN/2
5BGpHGAjTVy6buHAaoLHIL+JnXhmpGHfdm2FC3p0ZQtJaKD1NAjSS8YqmKkJHv2usfpmAD9dwW6x
xARQcJsYognb8AqJ38nMOtP4s/tYL6zgO0Fwn3P41s58snFv4rWqrFnsv3trULDk0l+qjraxzXCk
zYZdzJmq5HbniyBALhS68lzfn193KeXBVqWWSU3oCgzRkd6COcQSinXeP2pHR8mqF4F/wnSUhEw/
aC5NTkUGAvba2LWG0Hcz3bhq36Y94zpe4zDjueJyGYG48A+iCtRyRz6s6tBFFGs2Icr8spJt4a4V
NanLGnRIA0od8WUCLCwZYhAi2CdCNGTSuSVxr2CMT/fo6TgxtMOL7udLXuXSWyaq47JzO5jMN2+O
WtVLX1bH/JMh6Bxqy2JShfgrKwN68hDCpkJJn/tOmg1Q9cu4l1N7nQiOQuHB8r9jIYN9/aRE3Ioa
WgpXRsOIqIKH5wU2vC9khUytjqOyFlGUB835Dy+4B6/h59j0L8INvDV2H6nUDThzewkiWnoOd+Uo
awKvr6anRow9yFJlyONN7Nl0DOS2/kCJk8vEx6qdjolPsTg/DJs3Jpb5VzOvPRetDxPNu7k6ahh9
MVui59aWKgJKcoxaeu+l/QwAgewUkdAbT8uxizWorsVe1+smmw6AiwuYjqP/LL5ehZoCHsE0JJkI
3/BSjI9n97gF/Xgb+ykWRyZaYzK3Gc0Q0A6hY20lqh+dpyhvgvMBDZSEPM2lLYtxzOJwK5hH3lMk
H1XjxWSGPgoA9ZUh19mCAd2lNZXLowtxasefFaIu/hiZ19WonG9iQlIB6FYShdVuLZ3wpbUi4EE6
sk8lLWoLIxMZeI6OP+XExMO2V6DQPJbB2TQrntrY0RiZ+1S8LPZpWMQ+aWzc5sBSWdOt0B4BjZ0e
19c7oDM3fb7NXMohAAe2M2dbCQDrhXK4zPENkC1X8KrAcz893PoHHgMj26EcX+vlGvjEXlaJrm9U
TyTeZYtPh3TTfI6NTTrgn4VIybZqQRaePx9Y30meVNYGZ1lbmlrp83SxcZMbgSOUuIiXvp2KIQ12
boWSnRXrU7kqj8o/mX936hqUnR/ZSAtfHt5Dy/RmyJyn03Nmp6fLqbrVE9iuFK0z57TLgEqMsA0o
9YNMyT3Gn+EL9yCbk+jYQqse10MtI/C+EB0br+4ONonJkfLeeS2aIgQPtipMlgzGQ7D8kJdEkkZQ
Ffu91Zee1dX+jDQToqKToov+/IY6Ul7mUZAnDHJRnMKtQ9dhFmbkRJ7izMgfBwyIaJamKWbE04IW
eYjZkUc9t4uPZQGm/XOvBVw9ddvEfTKfpt0b229bTfo03l7NaqLU7ZzTWMCuutvSSX87TbkMIN82
MuilD99KT/fyyYHqhaTF69I6AA/dPRxP5hHbcmsIL8LGkbIi0ifNOWwJuAn+WcXMFEe2+1zCDr10
c+U6ZoW0T7HsmuNuQH6OQQRzQLyhMLvNUpiv12w3TUhjEROmtNdCZkejnM+Itz9MBc/8IFOBhs9I
jxGOLEcvI31+BfX1W4Gp56aqw45eiEiiXLzzgAa2YRXT2A2apwDKK8MuriXQUCAP849DqoYDxi6X
XAn4WEv9VkCfTGT5Jyb0JHoU3GXZ4JPtYbwTMn7f3IhO14T1RsJrf6KF5W2bVYqcohDVTFW3AIHq
6A1dM8jN9Thcv84P+3U0EDh1JPGVtcDKV7vKAEuVmO5j5jQn/ot6by0dv9CC74+nTyMSVaN+K6Pk
+cF/pJKcXvvSOz1aIj7W+++3vjK6meSKs2WMtSziR3fDzEFisLeVM2lFO26A+QkGRRAZp6OWH1Wi
SzPpQKQJIgcCbnyVSSIUkkHpAXlLUWnRhVJbzVwK1UW/sDUBF2XqjKZQWHGHVN3uaQLU3ZLpURPf
ijpHbp1RHrVO9WB3XTkBBi7pXN95eyRTM6ZD9SMJmjdAMIqKPYyUUhxwj86SjaLMrY6lQ2eTj736
YpFtwwMdghNHVmVKL6Bs3iBx92cNv/cuFiy92vZnPglg6RJTbum6804oytY2wbHs77KRI3xXcPvw
ES33Ax3x8jg6uWPeorRNEKfC7oud8CLkRVzMD1s0maT2kbwtrUvwsJOvgBo9PO389epYVhkNrbxJ
JxClMLa6FsBu0QQfl7gAySOpe0Gdqsma5sLF9ViywBp4ZceMdyS7J6vyLK+kfMsZ5CL83Wda7tY/
+u2AHzFHu4MpkABGl8jYcvnqI+4bGK8RNg/1TvOMCotrjnuvK2V7tCFN9jJsZswjAaXZQ64Ll3cR
aUCxYVPHy3SoEoXBhPkpW621aBo9FyxDRQS/9JUFnI2a3ev4EBg+gmNj24Co1RZPAX0IeJmG1FP7
dgQUAPmN7upIhIhuCiITk0uvtfLbYw2p3GrhJyd74/6xC0x2oRXhX+zi5kwJpAH9Nn3QMmUvd4Qe
UtgSnKE/vn8QUmbjlDZ9Vk/quspOT3Aq3jQt89qWwXsPzt1WGMIo2C889HkYrVHAYlhInxeoXtCD
KL8u5JcdRQ5WJAoE+XyCeZJ7Yts0iyQs+/SkBdm/fUEgkPR6M1pRnCTJwD74fHcEaybB24N6AhhK
bWR5hHCXfyC69bBGgPXZgEmcsUi3lP9Jd/JmtEo93gpCoFzBtsrqxz/p0sJPchBugIqAue+lhpZ6
wQYhyclppSXO3x/kV7xGxf3+Wl4YvItC386xbfviFP97x73goDTmRqBBr+M7xv0iR7u7BdSAT5DF
Ij0l46vmE665dBZgGcyZeDmNM+UQJrP7Jp0HyxEsTLQxX5Egd1b+FWfdXx+7u+n3I6E7pOMeMQZ2
KoWfIpdEJI+KCTwtjJzifwVKgwxmQAcx00jYTWN6I7DGu+lLLgEW7drd4qwdOmaOZUErekumixT4
4tyAh/OmpUTM9OBL+vQal3Is6YuK95kQn9/pMDDIAMymO+GopSbRf8ON1YVD2VqF7+C5EZWaIadZ
AfcUSGdkDTJNQu2ZTpRPlOw6HOYvwfM1iUt49mlcCQZMxgOKih35ooicCBbc1yzYDeqOyDDkI6SF
/z5YfcWdLz6WlrTq7V1m8z2wYZRq+wTiKGV1trqpCEJrQbED0BmBb3TWVn7SRpH9bps6QJBG3kvD
dTctHpPfJGL4fch6tMNiJCQLRJEjiJKqKtSw/xOQMBeAvhAOuarmfs0NlK/+vovd3VNMrTZ510oP
+wO/85Y/+eG+hWodU5nS4d1EXkohzhMqdM6t1ztKRCmHrAAck+dNa8T2AP1NEDbKwXXZCxTenAt9
HD07unlOP9cs/ZCM/Lf2rRU1LtxiatjEAyV9P4vT8431RwNXo0SUpZptf8QYj9RTywhFLoa+y8EK
HaoKfDW1/hGJO1Frv+P2vFUT2vBR6GDLScLURzSFn1nglOzYxr64SIEqczVvFjbwNelsyi4H+uum
8J8gJId42AltGijOmDEH8uqya809ryo7+EeXfgefyLPlr5zH4PHTyyUdnp2rEYM4dcKyxpNC0fku
xKh+/CS6XjIRZDX4yKDPITLXQJ3JAizBnR1hZbleUQc1SG0MsirYklhop19L6acPdsw8QHNUH4gk
u7Eza7KPCOKmLZrsgJq9nPCgMD/XwwGj0JK1pTFR859CxYtWeKygxNvEXk5uYTjeSmHEDTedssLC
iOMGtt8xUjSB3IkURxGFENK8k1FpXrFu7fpe9j5n6vLZWzMZ8ridYKSOVjX5aFEMupzg812e/w6d
n+4DLHsXwOa2cUv7XJEM2S4IHtNVnT4/S6LMXUQSLRQGEzg8eSPQd3BQN8jARz3UPpBHevk7Rzv8
4hGTuZwmRgOGg5tqzqd+uFC9D2r059CeEf+LdOQQ84Nvrmsip2FJoXPhsm/wSEuPFw6FtHJwGaQ2
593o2fCJBXbRsb2ewdyPQhzclvwhiSm0PZRsmugJEz7cW3xGqW1iHy9zaK5DkEnZSRdPTBD2SR4a
T/mOTQWnJ+lncnsts28U1u63ekzcXhQmiX0YmayTQeJh/zeZiqKE7EP1d8Ib7/3NmdIvWPRYJJ3f
cBGSf9FAziF+SyOYpailGYejG+qtxVM2hs9alDVY6maYTchXoXsZavZo3utW9aVAAjPCoAJzGQRy
LUla3zE2n5NiHhGiXyDtx5NWfEgmmZKLHVBc712Vv8hi8FuFa8Vm4WdNljwobOMuStUjIp2uHq9M
y64WHDHGlR45vySSsQAM8WARBaXLuUjBRXgUWubE/Qbf67JdwpZf0pLv+aMw94Sh5gWz0CtzNvGk
MbPYtIWxzLMiBGR3qDbp3obayC1jiFHUldyH4VCdIaIh7M8xIq70IzHCerMBQ1mhtDvQIohx4Fve
fo8A58PhLZOwQRbA+GNVyo7JaECwK4hrlzT2rwQ9sK6EfEHsc6MHXP4tjZS8Lmk2q3eVlZ4bNAjl
wy7pf+8m9RsrCrZ/cbAEtfI2WZZROYefHhltZz+mBS6659lyrxvGo7AlVInoL3v1tqiWgqpOTEZ1
LLkBdg133slJk+2U+dlO0bz7VWwUolnAFrDsfqA8mtVPLTbXtR983rHj15JVujZqI55E29g03wV5
Mr4TYsILHqEJ0i147n0WMUrievoKUm9X8Q24nyctuSKLA9YEEEAWPywkO71ZoXG6O8txNBYne9Qr
sXvYGuXJXR1s4pl+RwS2OJWMpjUQuqONJfccPT3Y1hLTL9jtHN+lbsPkGz/BybRLasdlKMe+n2vo
yGOmJ+S3B7XQ8DH+Yyg/potpelqRwouaabbZcaFJxAHDOfdyVXvFk57GCtxe5nNVpLYWH/fVE+jW
mrpDM/oXHHNJrVzch2m6JSYkb7OwTKywxg4NCrNumY8gjB+egauHcoi55REMNeSa6OaPh6Baeafl
Ivbp6FGZzHAXvD0IkA+VYmuAEaT2cFhiznzGMnv7NFm9gPe5Qp/+6wM1rY7Tpg/eGMGYw4aUdrJ7
uIV2Wjekk3Gnz0Jv9uS18t1mOFUspD+emP6zPm1hBl2JH0Byx+SWqATfyE6lmmYBSFpkHNBKbEBM
2kR8XO4o5CZbH2SrhVAbIpH0dtumAFIzX3eBLPSrdpi3hd7X2B4Hy29gIDG6VyZ2kkwhKLU28IG1
iljTrMjCeBYBVikGYcUK4adNeYoD6H2maci4UkVg6YFz/qBYIurX1f81LuGFZcTrM8nXUt/DzrRb
fkzc68/xwd316SE1/ihd4El+soUvDpESfUtFu8CC+FBjCvJLO+3FQYgv2afreUhxjn0i05e9sQBf
jvvHbdaqFEIBjsKgL+6H6BcsPAhbnegIL5+efLd5WjbzQcwd6ANg6CpkIZzrS3ILPTpzstT+nBJ+
DQr4c+6d10HPz75UddkT8dWbXbBywZXR++TpM6yL3QUwtsxztAGrzXqPnH/a8whYXDtvX3auLFMW
nnaQoYBuebwelPHLkNebykKdvmP2tur+ASB9c8hIBh0jNFfN8XzeGTDx4kotRtWxZjPkz1vChipA
bqAkCG3W2frrSQPO9Dt8T+8nfXKLgIhYecC4lL6S/LNZBRvJBNQSBm05S0mli6++0Mbg5WjkHzGd
FgroMN+6Ra1zhHBqSFiDrzkS7X+yNSaMmZ0lm+SaJnBhSSW1Sf8utraap4JLpR1/xCIUiixoTkds
s2U512Mplja7MwNdTUSVIIBjh7Uzh3y6sNhOfcsTIhoZHY+exaX4DXpRKgTClxY/jxor1buanlEB
zWzv0oVUbG3vVko9mlCwx7OcK3ESyR3hRgfcmN+iA2AARt7jXzha3PttrjgZgrvDJn6e9LHPKeVj
CjpOIO3jlxsFqzWWlwzxoka2U35EbIqjK7EQYYQSkDTnby/v1QUox4X7Frb6zJPrq9eqWoS2pHWa
C9KfSWalzIQFIVcW67lWVUvjlYWX3RBCIkBsgHqQnhy7r/MdkQq3VK94dc/4rXdxDc/3g4GQzTGG
lh8+GRLiYa5iwR1hFErOIlMsZCEQENPHck2b4oczq1HVrTX7zfwsc/PrKZvtv8+gC9n6sPY/a12L
vez25IUhyTZQ8bMJGGH3YhvDDjXGRNaGhFuNd2PIhDsZG/e9hAySNR2mJq0ko6109Jm4vTQu5S3/
Ls2ZxJUmD+Lemb5qsqeni5f2GhnHw98irpAfDBezejb+cmpAa//Yl+TFX1OhnZPxRv4ORSTrSgI6
ap3XpnK0VAjVkGS8BvVc43lXZGYAEQ7xB3gpWwy+fPyIntfv1iPglGPt6zW3CjSYytCKZwSl3LVM
IY5K62P9NerOGG330DLA8N+NrhTfc3vpDGWkfBiz+n1H55arpL9K6e0qTudIcvXkGnvGbVjbklej
4ptdzK875Vyu7R7Un+2LGFIqCTC/GNDY0Y0taI79Gc7imcWH75AMrX9Z9Qkuni0P5qpIJiDzLttu
RHeJIw4hSxgn0B+9tIkjB/q4FpHo2+C3j254DqYTtWLf6XLfSGM/rMH8HlKzyLlC6s7zxTBTqrvJ
2lSkqS0f2lnCnxW5TmvLFMbd5AdX2fUyamq7lHgdGzRsH1gCubQsU0RHdtVcxgRjWVDCcvguh7Zb
FrHVjZzN50t/x7dexG8IN0S02Yq9pxmsK23yIiz94FSfvwmzD0x4Z29QRZYqkEQJEzluyRbUyNPu
5s+a0qrSKy4L7kjuPQiLOcr0rzXpQwL3Z41B/r9zB7YeyEYN4aBzjtEpEPM5GKl1EJoGM/RL/nhl
wYMusUnPTXbiaKVzNhuYG17YuKDMIVDX/kCqvJ7oO6pFwORqWXJxGAMlfKmARShpfYUyW+sBqqEC
yhX0QBu+HkgZbPgW3/9bMwtI0cteanuo+Ttxx+ni7LiR/5nKGgyEzwyR0ZgDnQLRfV2MZEUVKWji
ipJgegE/2LrATaV6vVbxodJE2nJ0Xac9NfPVQTEnwq0wfWHWSJWf3GnXxc6JkpViv2kLqFRfjVOp
XmXZnF+oXPbZZ0jFXLREYBvjMREmwbeZngJ+tnK/6ZJ++Tsxj2stvRWBuPodJMaJNWeUfI0OivX9
Q3vKWb0ABzCvv2MYZ9bGEZ/K5c64u8QRLIbrQneBzp+jC0yk7DCuPFWSTYKVWl4CVPe4nmEN+tde
VmodPQgrk2cjXowl4wS9rK8NTnGLEno8RJfbXKd5YLZQFyneNtUjwUx6ygcts/WRFk6rQVsFTa2F
Gmh/0PFgnqUCdJTr/M3xC327bHhe6eDj2QtZZkOGfYaav33Q6MhqbxvnC0QKOF+v68UfByA1bCIW
7lamyVzmNNbihtSP0aRUU18rgOgAlre8LWscMyoeJVQv/XWqSl9wjTh7Rm1u+23P74zZL5zOmJxm
2XXSd09gN8525U4B07X6+K0/301ji/mdVFiHpps9gxClSSvJMJbQWXb6Sc27IbdrYj810owUl27n
67G6MaH3F5o/u5DvC3biWwlaQpBy+BJi5DBsHit75Gl8YSY9SsoHorNDV3Bvb3JealpWemb0W73K
9n/QIFZhU1sBJWMUFWbypim584SfQyOIT2okib4TDctUjp33vwi4MFCiEE28aAhKLSNG9HRXvIbI
NLMjdQfaezxkSM7ITijBrQrUhyCBVtmlEvuYuhsSwXwSnhqwTAFhnVMCWf/rJz/1PGKhoW4YpDL8
QXQdQmfy4wRI29yEfgOaNZRalpAibP2pnG7IA4bDzrIZupy4EL2XKEgFK7Zb9zO510V4jxWqCi5k
gIeKjBjy3muklU4t85L+0CVa2D6mr6g7c95ID6/60dRSiOBHBjiq5tdNniRjC+9Z7oN8NwQkKC5l
aWbS9W/49DjUnIDLZ7Gu4luonntotC/4Ap1WphjFcyK/9/0JQ3JPCJ7DjNcyCw/f3QnUYnh2K2yx
rLzR1g36cjQ6fWsN/f87Gugzo10g31hPCDbncgwzNrcsljm2vdMCQL3t+VCooDR+hMRwom2eiX29
+o7hZ4Dvj7ebJw+s41kEP1ocYJkYkmiYDNYyvz8VH5SIprV7iKSwPldhYaZ65WFHS7xWe3ILFwLe
uN+Q3q1eWI3awyK6liGpm4HO9Uf0ehlifG5nGTXZJZ/B+++OSRnxFFZHMazahB+t+uqRv7wxsoYR
62PZuIgug/OpXx22Sk9f7XvsOPZq1c8LRBnRAF3I9VyB1DAQYMxbdacWTIU30x8toxCLYsMFJ/C/
FpZ52s00+Vt+N6YUCtE2ukZCTN5SXLZiiLrNr8jE5G/VTi3+5oHBedzcmCWpUkALOWFaHz2F3T2Y
gHb4/RZFbmumwPVAvXiel2D9D56EhvrArbRcueykxD/DSvpzG66BKDOFYbnIG26wKC7/Kq2ESYjv
jVAVbLMhdxiSDZkE8I9hJDybibyZ+j1OQjWPoFnQieOqUj+6bC3U+j+vuCAGvRLAMS4Dz8LjU7Fc
F/0qxbdZv8Vsr+i/4kl0PPVpoQfLkjc37NStjOzSVIcbdr7mJqntZKpdU9Xw/DiqqWL15AGbh35e
8qGCJcaULrA7Mgk+OLeEb8j5g+Alw+HwTW/4LiJB1en2k58QbaFARLMcSbUM3gnxsAoGMjk4vNPj
wuNjYYdc8YCX5bVOa0fr/4kz+7+7bzuVDQ/lRoKJlK7xo3BHgMtlfxjwsfMiUDqttYcVVhOWqt+J
Se6y9DYRyaq9mBFRka184+xgIRoLktx6Qtiuq01jrUVYhGRvPpr3ivqxlP2Ed1KiDRDZBCymKrm1
Izbyd2NTBuypPtXn2VExjV6U8doCqnDJ966JTGvaMPgBgTzBA138h9LkYV9O2h8gUDtUPYkfXgXO
JYU46kr/ebHP9d+9VkRaf8e7Zx3XLz1f0ymuG7+ibbivOMPnGVBppvJqYlLdjzSygsMnHFiPBmfi
pe2lEZaVyKNeTxamnE2iZAqzkyTcn81LpLTKzJuQzroVNK1zSgfEfkKZaV1ZGcE28I7sHuzB1YNy
r4oSAWD2aJRGJ8Y7IzIWJKr8AHwZj0FDXve0u07+zRM8LwtUlbcmAMQfAYHhC6A3TvgGlQXx7pef
sV93UfFR1tGem3SlY4p2l518t81mH5rGD+QrQhemluCphSH7z3SLtPeXUrVf8Pox3bgDMztXn7sv
CCU1XpA6Vplr/hBoNGJK+oiCBSWND3IbQVbGUjEGqD75IFt3aHTbKDCF18Gwe0i6hobEvngT1VP6
BCAG8zJH4WSPDGYOXmEl5+VuhaPpIesQqFjvNjXhE3CsEArSFsu0UG8lRmLq49LVoiEo2AY/a+Ra
IWCftW+KAzbCigAJMJJRBeFHWd3TJ59Cq8JWL7ZW18c5vDM/tpBFj5A10a1xjIyDbyCgG7mENINF
szCCkKF0uXd5SX5RyyK2Jpg+Vu21xBuNiisUZumIxI7PP0JQEKfn+ajJFUPEFJ23TM7aHBgHiVaC
s+zTkkOizqrW1Ufy0o1OLK79vZETVN5gre4mJKBy1P4fJdknNmyU9ZMPVbotf3H4evkg+RZXfJxX
QuXrrEc/RslSEgExZex66/5LWRzg5LnmICaWY5Q384DQUCdjxPc6Opx77yRVqBFxrQWNXBo1BObC
CeTqeF26TgjVTCkKw/eRLPUjzCheI+1FjPA1gbbVQuxOYQxMPE5WJ3r2dWLb6T1Xjj9MAtMl0T/l
yZHCyLFEFXOKzJtMlw/NZPwxWgrBWA0csHgrtUSmtdHSJyuTKQ/PMS/yVBtgNfZ7xH9zRoNvbXy9
HPKoHZxBLI3MGy9JQlErbFZkUYzXWfIva0xYLPDMV1yb1RDO6cX7jq/a23PFntXkqZfPOChvEucu
Fmzk6bP3kQYfH+6GSJ3HY39Gbuk6xTqJkZKXGonTHnB59FcdhBkqSKJ5s4FbRrCd+DbVkC3gzv3h
ldY2YRUFnwCZkpR3FRDt5P8RoMjthNkqtHTPftnwRZSejLlr4LaJ0W08mjhx+jLsuNquXyY0DGEC
v5Af1z6R/mR8Rzfgp+VTCL/iIkOkQd8VBti+sOoI4IYd21DoTTwaO+ohtlGdiuGJ1+yhIe+sPcmX
YogoS3W/ch7DAFMSCu6TrsYQ91smtER6tKcyr39fOVDtFplHdqVmKuNvMOV0dtcNXuJ5mTVbdgB4
473Jal0ohE+dxpcQSJq3UqnXcs9sxYJP8Gq8KZpIVQREux2t9wdShF/2Zn3VAsv+DHTr7bQbvYNt
V80NNnvR7BBciWtZz0gwqk3h6kiX9DlhZsTP9MHWV3YrbGHvbd5EyqdimRZ20U+vO6EdhNp95G/x
8k36Vw47DyTV4pg2iqry9rrqT+S6dnGwprj2vz8SO77Pssp+4jRMlt/OTBjNht9ufiM0KeTYKSdO
YifmELNpWw2YNm0X8su8Ak87chpv4JVRnwMA3iGKt4tpUjhL8IIXmB+2a75Llg+pErZrJiIkM+0x
S82aqOCjE7PCEHAwqlLyVKhcAW8ua9E3jrfE2nGGfL4dBLUerCqciH9nNyIrTh4uBqjwNPsxl9gf
tUW9bgLH4AcfzwRf34s84yEvcXqtEaLr5oEgwyFTJBcJQUwS0MeiRWbeo2dA/7HUmXqUOsYHCB2W
ZLkzLCpkRB9D8i0+Q+JELZXuih4IP1z3cuHR+ZvxQNkmMkjUe/PFJWDtMlR8eDwdtpNRfxT09PuI
lbt0aVtXalSV3ex+6hlovBnBjrJKzlA5QJK+gdwkP0WJso1mqu38SrtjHTzDCFEiDBlIwQiBRq9k
j7uyHVqFQL9hi1X63CT6pyIT3pjg9VkD0TpLUElbAzlFa1Egw2L9fXVkGxmW++8oMUl4LpQW0U+3
1ex2jgUlJmPjbG6Q/D0fD/HI+j/JazyCBVbYhRRiCK6MzOGKDXOn7Jtq8VIT6Uc2DoepKE8cS2bp
Yz3f3KeOW++Qg4MO15G27g3VdG3IVYDi2H/Axk0t3L61nRjpKZDMGRHcqAhqsLrRjvrhddnXTnGr
w6vt5X8TwiRBjUwfzSuWAibg+T+We6eKl3bBJI1xj892d8e7OetQDq2SZbDoKsppUGVtTgbJR0ap
69oa7yGjlDyN7QhBcFasLJCfV6LO9k+4xAq17wtun2gVHvcv7oX6+MlZ70+B7jttRtVyDWjttD4R
uHP4Oxw62plUdykplpy+UnXnCrKdtK6X0BhfHl+Nnz4NxsInKDRo3A7BRcjsXf4vn/UOHI5KRrao
sXVJ2qksZIF0/pGukqHmaENN1Gbbe9wLumK5UOWbRQmmKcwFNMBRxdJ6tAN7QcVW2inhAz/FF6dn
+kt03FcNKWEKHdnU1PmmW3YgdJs58kBOLzGM/MsMxJVaE1xTADPYFBRe/Ad+JXIuq+9S/IxPJxc+
24ejHc1IAW9EHPiSU+K7Rrnk8z5moXjkVRcvgMXdhw7lvkcg1YKM8/hGRRI4dMO+7sZQY/bsbwrl
Fc6mpBYpeidUvVDsPzhcwH0+1cz20610MFXFY9ZGg5V18YklYmDTzNtfgGTc8KbLs0Yg9WWbtE0r
xZIB/MxjjIdkqUddiQIRxUVeM8jn1i9vnglCeKxGkqiXFYh1SwEZg/AOJbWEFMvIvhNLjNJtZsnU
EXsbgIR2km3f57MWJuiQ02XIYHUKu2flzFmQIRwEnuHwnbfQJqzToCT+0u+Ixs3FxkjeLpa5HiVD
4D2VgirAyimSUrJEu9Ye5FD+M7M6Zfs6OXBSnecNO/TsOI2YDBVmC/CiBUB3kLzyq7M4rmX9vcse
Km1Cm98lf1pG13lU28vN1HY3uqglaR3ChTt/ytAakNkOEOHhVxva2jk0SBkademVliGmQYn2kret
eKv74XICf+wrY/24ts4Ge0OwXf1UUIyGqnAnERGYhvjRACWp7Cy9yub3AWoSmhTs5dIFr5v/QyZ3
zLQV6nR5lCFiCs3g6+vRSZEpIPd2SkSzR9oLW37VWPiEjvu50jFx5F3sQyezOfKcpQNVn8iom9Gr
2D+WldzfUlXWeRS6oDCFNu1FYlNwfh9bHEveyQyocooc2uS4dFPictuDSy2v5PamafQKGmLv7Vip
nDGTPLbVQ0z6XjZy8e4UW7jIsAxd5mfspQx3vXh4He1U7ZG43l2Ly4A4V+vhzH7LGrcVSv35f8Xx
wIWdq5zv31EHmDb42FP9N3OIv/4ipTt1vN4PoMPNkwAndLmq5oK1ze38BqlatI1KX3YhtR6VBBRh
pjfehyWIWrprlKNv/zIbQ6Fkym9wHO+YIax4YBDGAfVYDLhetNknQL5tHMqCJ4gvYivZKJbeccTA
fzD8LjcqHKBgx3FeKKn9OdSJQ8MXrCbAUYY+Ap/WRP2Pm84HOud6lqV6sCWENgT+eNPZ7+Ueq9yA
9TsnZjO9V8aKMJiLqRx8QsikTjgyfAx4XygmXcwtCQ3l3OP/yrtLXkerMb7gdS29Tspl/wAN7Zyg
M8WGACVxT0r33qVE3Pyd/EiupUrDYhr5m06wzxI0DNJ3VNZVDLyuQxha6jeK5jtFETBpebgn6UB1
WLRal+9i+QHOdb8krLPzy4MFc3jSeXza2Qb/S24nfU42h41cmDvGUks2ynPF9IFmbY70x5NJvX6w
p0818TXTGv0fNPDfNS86MpZSo2h3wrMBq3awCsZ8s1xHsSu7Y6ZyHuh4Zl8iZeChx0R820xuaalX
QXX7LNMYBD23t64Wegviw8lwbJRInz4Ia0Vv6jjHdhIxrW5u8YLB9VY39bpmCPGxuxCckF6kEa8O
YSD9yxKuvAunTt+mqvXU52y+bvb15oUyCr4vHYKlRyTV+b5szxWsu91HNPIW1laGiaIK+FV97tg6
HEJVrgFBS7gpCRI9XCrtraagn3NrVEFltzB2Y4tTMgvtp/vw7CJqcpj1QnQVspU7edNj7E9EUjSn
LNHD97cjZ1w48Xt4riqResv2HNCxivdwMLOJVbKZAnZjPtxJT10nl4owHsxhaqYJqpFYbGdxQcnK
uOG9OzYALs9v0Lj8owQk9mXvy+5F/0zokUvkMlCrd0RumwODdho8iXgcj7tr737kz2/kI6WQaM4H
xh008RMOiH+pnzDZHaeCHvPCUEjIeu/H4oZFc3IraFyQBXH9kSZ9NkDAj7fP4gcQyedvFF89cVPk
y/MNP5fDeZnpgd06yn7cQHLu2uY8L7qyOreL+fGy16dBZk2bd+fkYYoMQdpqEOYtBCFO1iTpnpBD
F3GWbpZ7an9WlbB1rQF+umCjLgENYN2Vwmw0PSTOhNlSGi2ohrPMCJcRe4kdwoEQS8bbPPBVrq2W
Yfzgp/VzW7uGEeZVbjcenVTmOzt5f9XMauPaTD2hLpBA71uN5unkuvHYr2abfL7rOpslaJDHEq7o
pXehw3hZAD+o/sFDDrF/ZSNy85Plqsonyd4Bgz/tmrlfsrP+7eaOxNnBrXuw1xk+D0fT5CkrkaCF
bb4FRF0cjWdM6QKf7/2yJHaV/VjTWjU+aCjV0T2GImKU//rYoZxCKN1sgfnkRHMB5dxW1XTlDTLF
nBFp+XKXFf8wzwaUHJ7F+jkDmRuDRVWqYVqq41GohULbGvGAcmjdonYSzdH7DOMeanUadfwF7DYf
GqGdOK5Y7iRICaqqX9TKHoLrl61TSJ6dH6riwyvx1H4SQNKeev1BGyFLf4hI70Vzi135AFHxnaqM
7KQGyyEdcRBq4lVa5bGc9HEjL3/3SXfIKgUENUcYouGLwomq2qlJlM+S5cA9iHQjvd2E2t/L7SlI
Us+1Ff2P9QoSPTLrWX6siGB2ZMolXifddsDQ1ljpc1Bu4UikLdPfQQlPrwUCFfDh3V2AT1DexAyv
/DEq5jrUzYo08DhDmCn9i284pMuEeHfckpcPvbjWfy0Cqx2jOzm9knOA6z40Mi6DJ0/AqdNyftOh
8fm6LCoBbNev7zEZYOZHglG0rD3mjLJtbzxUVailj5p8Oi5ZTZNDJlgtHX5m2k/32E1aZOrFIRa3
YmsYPXehKW35sNYq/U1LuHucTeZpmA9C3rexMlORVEIwRoBBbVGVPEF1cIi3SoesZsadAC94qob6
hXKFAmfK1WZXeMXOwMMtmVn1z79Qv7oWGRfIEWegHqolfwlgOQdAlK7FO+IW+1P3zGuPV5jGrdoO
tcXqE2gQcw7QodV182kGPD+8diMCMssWDLNsJ0Tyi3B9UrfRrL9FHaghHnGXnC5oocQKvILtI0YH
bW8AYYqlpHXRzOuy5uW3L6A+u804PtiGlmHGISuB8rHxgti1nhRHXr2scZ6tSUjYkjaF/oInoJOn
7+o8cM25h6dywddusdsTbJVJVjKnjX/xhslYB7SUsR2X9YvgxIqnYggOdGKaZs2k4SlECM3+2D98
aXP7bPoTdBFIqFzMJmdItlNELA+T/RlX+V5WXk8oCLMj5PtV3rv/DTYfx2EIwikZ55Q6VkVw/mAT
Eg/8EsntEEV+iknImSk+2jNwVfDED63XxVRonvL1zrD+P1PGAsKidprQo2yXS0Gf9MQiHkuWrYQj
leRQ9+Td2RiGBtlrJOQkNaTFa2iCOWv9bjPP5xysHwZqKW4WiI5uDZBoIoRsAF0cXyrBq38q2YsB
RWQTGOFD1vQInOXFf2vxqyRIRVx6OzWM/5iaHr2gU+rQs2B4DQJF0Nx25AH/8LAQFXgC5qE3NRUo
BydF9mz7PiBRlaXp43gFyqTGagzDXGwUkI6cUhDkovHoWXUIeuZQMgOekhPzcZj5S2gB7kM5iWpD
Qh//45+WIjI8U7a/ILzKQWQ9gMJCsV76XKSZEX5Vymut3liCinI8H95l5W6qi6OkuGB91Hxc+HZF
KVAlvQUEHgaRD0z0pE3uaUPioC0uEH95eCAtkWvNFHBqwaPcUjHNQdPcfLaxVJBQvuHpdN08y6sH
boPFo8Pkqp4yGxjvjjziyC1Cb8bmwMXP1KR/3LaqBQ4Od5W8wGw9IvEgjvfrxmr+LMM4puecCwv4
xc4oeUBdaprJMIfG8aM+qxkdOLdOwHmrH/fCzwVoMLF3UU6rGqNEz4WNgzxgMsvel/hRvJf7P6P5
vf4mo9D+goMasF/YGNLzMdvuLsOeE5vxhRXHQCEhHfRxcdoTkckR1RZecA1Ousb+nHeUUFLamCoo
u3vbFvTJe6OMvVwasGoJbCobUVBU08HlMyySp1J9qssH+KllcRXTSOkN+c/ZZPX7jatO5eVWnAZE
KBnjtW+7yuOKe371Ms0BtW8h/oKgzIQXCrR8pSXRPMzsTi1R4a5FQVvaHxLooVpLmCzIVin0ytEb
lU5O7HP3SqcpfvGblNfsJRUVcxVOYZdRBlFcuspy2z+ox38PZLlMujJUb9vHvxx9CV4NS/Ryk8Pz
GwvzBXXezTbJ4R8TprzCOU7mbn1Ss5YqCMdJhAnb0+Fdf1deSNIWEdRszoYGrjsqXXh/gpbfHzNA
swploYjSJEabIjqzhZMIsbb6RRGwweyEbsDjeJ/8dybMW3EV0QrX8epZgZr+QXvB5WtEiXysf67y
aKETMkifD16gEEIa6kz22t9nGbXwwQy5rRmypkQkY1l7u0OBBK09sOOQA9IaFLFiXp5PAmHvI3yE
0hlVtZeSKMQozABmK2ryw0+QQai3UES3Mq/gq/hMGHVqoDnHD9RP7wddIF7483Onaemo7K+YL7Cw
oCnRfWzSeN6RbUvm6CGReJaEn18kffiGrwCIDHmvroZS/MfQlglDjlwqHuPxHna4MFM75lSBRMJG
xTU/9sdb+L4Vog/2/h+74XqGQV4Adj+9hy6FqGzn8xouWf32rVph418cOWauGtuJOhPbXvpT7/O4
YU1OhIbnXzl+32JA/5omyensbPqqQjBQTk/R2OuS1x4vPzSAN8kQ3ed9ubWNMUsG5pYYMq42yyNH
iQX30yzKgUQrugBeTjRmS86ZxPtiijtJsv86dZNuimWMrCTgqveEf2JIP4+sYau8pPPvQLOV4w+B
ZDMSyEasFkCBOMUqo8QTyymLvJ5aRTjhOyGviGZlOCCar+yC9eqw3krRCvxq0RHDLB3mzygzNC81
VMwCyRJqr88N1ZLrGDh9QKjuRFYkqXUptQib9ojG+Rmg1vvvhmq3OlGZjOK5TNkdzcZ0d4gh/ha8
5YYzhw2E9l2wt5eDb3xwIzJyQjFVuONIELiW2hxbjWFIX+0mSEwFuHKVQOZ68Ea8DuVa4Ma8oJ6C
13nM6zDyQbpXLg53yGxXQ0cIyWCTirNpK6JscPYrrS7ZOtEAqSnXwDg7Q+BSUhORgbMjTp1hthIY
XgcwP+GB7N+7b5kZY+SUuBv8NENFpUygt50jBcRirLMkWYPI6id/7dKZPXPCRlv3l+ZjNKeoimpW
xonEn7VlXBMEOg+1rJWxb4SFD2GIcKI+E+W0TaPaB6z1yfrxnqo1YRnqgB/Kr0Kc5dZV9dGkv8n0
oW2+GzaTlJKMjVJyLqWO1EovI9JH/YsuR5yjHFy25ek/KBMTPUZ2eoW/id5768fKOPkp04HF1PLI
ssoMJE7T76NZh1ycXne/j/DZs7tihSxwweObQ2loGJ+H9l8+vjja4ldQfrUQMXl3tBdd3PdQI05B
RLAeXkplC/XGcqMrI4sqLnQAC1XqbMJBPb9qwOa6hqPNUAf0k2MC+AogbY6utAE9Ln9A0GYkskXG
dzErSeHu7tgAfgjaPDyQrXu5c/0OAAtTnIskFxStA6KL0Tmh8QZ3sd0v2ojosgXj5gxliIFOdDEP
pF9tAOiUf9P/JosKjrGBcXpyp4I3hvkG+qgqoAfvTZK0wTcP36JbT835vC0sWo+c4BnUTfdnCOPi
+iOfl00c7PuBzNK+sP8xj/O5RBOAHuNbIgc0KgP2lQhOTydcD8zRitzEvNYaEi5xa1X6rp0JUgYs
NmDWAEhJQcXuJ+8doGwrfBjPRPCJQpWOozDgyUjYTcpz4uufxF9+LFJLDbRLH2Xa/L2WzATvFT7I
1nHtevDoucLu0hPqlUFpa+dNUS8/7zd2myuxaUKQfUk93ot3+S571ctdXBMHryEO9UgSmVI/HmOi
iJOS/zVZ+P85nrMbQbWfzpYs+KDgjdgK8wqZN9DhhL4WKcQyaadKSQrfggufTuY3yp+86Zf6ttmf
pzdT+GNjBWVl+fWWKN0NqI+YLIfU2cm8l5icrrdh6zhuPCbMuZ9uh4zBNVVyPYF8pRNpdzYRNza5
1rc3Ole+3MuTfT8U7/+vIx7ggOC4AU1zwySt42+x6R9oVn/LEehbZlNxUZTMDHyx76TTWzjKVoEu
RA+FCIgTIUSgS3aIvwffb8u5F40pRMD8sRrJZZpYhAcTSLcUl3ds+DC7GT6zs+oQ7oec8ZRaHNkd
WKdGm5nnFNKS/rZJbWomjx+bHofwRJO0SrO1EUWuYo6r+l1/6AYBqnCZ0jvbzRxi9Z6YpeG35IAj
BL84be7vkAaVN7w+51brp/mAZmG9qDpQYgToBZjmL0xJUolpa/u5+sz+RpFw8vTuFOEpj+hm/wHP
R6BOjwCQlReswVZ7ZDjr6mp+IYoiGnHtVD+t0acS41zY/g2QC5Y0b6PEwZTqXt1Eaqj7gA6MEpbC
kuR3BEaXEdktJ/12dekPm9z29oxCo4jWrvoWm4Y5L59RSW8gP5UUyBP7Cs97dC7c1MHs2ELKv8SN
9M/vDFgjxP1QU6foGIIcfHcive4S0VL+d3QWm1NaqWKKy9RPyuWh3NKUMJj/AfHK1nXdrg8BXHYE
CyWO6gebRrnqqeYH3ZOfQyK2F62kZWnklwuNJCyVP8SoMihJyGa7p7qPrlALgk8yncPolu5GkSis
PEZ/z18QmIHg8pdR7Doiwa6Q0LPGVFosFanL7+TQ+8sVSAdH0Wa1zCpyVsCVVuN72b54Xyl+XxMS
sk7Mkgtfjp5dEgzBpIINS3uUiMQsHdxTRxf/K8Ar/B8qyxveAypBMUT6Pp5DETa/VPo8vayyYn2l
aH86smG8qpxkZ6zdfwZFC+bZZI68bDUOxjnf1rya4iqJZyGJxYR4tFg/rcvwheV8To9ZJSXnjHps
6MT7cRl/rzFjMTIo1bf57/It9WRBAJ3d8SG75zUXZWpAIg9pLhRJSyaqhPbvRnkjJp8gDjTPNzFq
KBG3IGcHAl7+jDjXhd7MbiawfBk8pINFotNGhAnrYyJDyzq5S8ODu7LjPEvKYkOXtnMEbhCYDkki
sptPqLHN/P6+TJTC5XLB09Tw5Xm7jrlrf5BVcSB3oNRDuoobtsKraMxCAjKObbKbXhom7mpqzklI
tX3lQ3IKfs4SUSXkakBIhQdpPfvLSYmo38jr5j25jTqR75Ljv9+MnleNGMl+GIvaTQdNDI64D1A3
hwK12WeBzrLZtdO4WYqpt4M/EZhxohC00/e5WXsa9KROFxTuGPyFV0+6GGoINOcNYzze8EnVIPwT
rCWDvlU7BYFq/GJwd5CHeQC+wHv2BOkiToGkINFgt0LhSHPupW8LYnC/+JsEgDd3zK6hp9vBWx+2
JKQuN9+ddFqoFooE1wckimuP1uukbsXruh0vHuo17hdMfEhRK08gnIh19hPZa9m3Q4cZ7oXKSoLx
e+TCaVV/njUjL9R4o18mj/tJZAj0bMVEWtfXPq9vzzeDVg2zo6/m41qUAvYDB3GEOs1/HcmqcYRL
aLEZozJarO+q8Xslp51i4c5NLrIyXB0V5l8TN9LOKzBcNeDFUfHeqvJ9SUxe4tFBqZQDURdhRWCB
6jmyRkjqGTf17CUzlsjeQWk5DQbLhmC0VVn2ZEH/6Y5926QlYRJS1+HWDHBdpkcHuz3jYNXrRUHx
JvD8E2jmNPl20ZwrIVaIchmLRhfrxDfl6gAAVzx1XtoQnr1jhQNQOcHXy4Dekqwl0paPgQlG3Cz7
CD/tNDlWeqANyPqLm6rVYBDuSGqeyrj4GvPImBVI5Qf5R5UORXRKQYChQzEinjWoVkxQ2fnbkL8O
ASG4KLV1msMGJWWk1MgBdOwlrOYPg15xKlLvYLUkRcAUKQRqaSNrQK4EuS0xnJzISiAIfxafm1+N
kCBxL86xqpVmpm9jchFafzRRNiicQtLZRckMogx55A88aSwzfeMZo9S48SUgJT+OCUIIiNlxyyWd
VjyjDb+4VimVvcKqwKPFnQ+YQx/XSkt1RVu92OcdDCs1o/M3zuxW7RxxkSW2+fA9m0y6tXnBqgka
xrIq8GOL3jNMuof7HWXhxUw47UIQJrzyApgBrUZqNfFWwYoQ7hm75i9cnVLrUplZwYVJs6lqlJH1
3PUyH36v+gm88yXInQyyuIZHBBTTFS/l0JW3RsHRW5BKVeSgr/QkkDeqdhLrvJDtjnWQQQC1/gXr
Ce6QahCzGEKPwQYut0hTU58Zog05S1zb9eHod0hLIDHVhFaSJJYaVvDk3gvAoNy++ktwvSHlylYW
urgrtTuq4Obi+OJPAkMgV85IKiNP0ndLReBXG/H7u0sEawGn2OlpZfiulVnprIRsF2sGp2UMURr2
bWAfgdWQhEav/wCtTIFctbbqbl8/GQK4ZeSiJEbbzeoleiK8dQ6fqHAMrs50TcqIscNDhpHnvEw6
g0l5VZKJccMuyzH/JzCeRPxcNKYiqaRJpqcSHYbbEl0zgfq+SLlKnaJ4B0/b8UM/9edBQwhwwnuj
ktxAftWTQDKzuR4VShfITTakaMEVwyZ2qUYyNVRBLRDl19fILu84C9KydV3LK51ZrTTcZRg6Bkzw
DSzxVdjafk9xoj71uo4NhkbB/8Pk0X8Nz723FhVXS5diAauRh3wEe85BHjhpNKs4Lg5ru4LnOt1X
5OmnxWwltmusn9GZinjJFIPXkZ1ybiSAWWkHMc2QsnSaj3pLAXcLXBsITDFhFwPbk6KulqTVfOX7
KRre0IXsur9CX6nEHf72URYDbFCTcN5caEx6z9yvTNTpdXYUaBXZvT37tqrrUsrdpj49LDXG7TSv
bN+BpL5rVunDd7RyJTC0hi2ePvwgLLOGxu3IIv/TFW+hcJmLfwcRmy6H2eGEx614XDWmRSQoTtjC
0VdCbXTbYTTwsOnJCv6LfPdfHfgL+VWX8s5g+7J0RwXxQpxTXVAatYmieb6IAJglguOFj5O3moSv
+3HeErfnC/9uKluun54mJyZyKslo9zu3Hxt8C2Qtsd8gKhp78g0LrTHxh8WzXFC1VAfLSfq3yz/N
nYd74qqsvW4BCWblc7RF0N9f66JWqdBsLN9Dn2i2fiDCY+YtZ4CvleRBWlK22BIsH2hCOVouTDD2
2YUn+3fBvQg6Er79SQJZeAGzvc4rFHWdEleuIS1fsR/iq5/DuuNyvBXT/nbp0r2V7nvaNYwi4+K/
RI2wGO6dIHo9EdPl1z/UoTOwJ52Darg9pGN8eGRKMn1K5hVNq/QcPYMumekbxORA4BRVAdy7PFb0
RdDmDhKQFnPIQ2stuJHPhf+es6PEguQulgzb8RodW75CmgPVCeTdFeeBp7Yp0qSqiUzFF7R5vAUa
UevQdEUeA8pANvtadtVf1PDZQKIbkzjGIubD6v6t3ZC4dWKcT10ayY1N/1FWAECkUVV6VG6zlFWZ
XwPgnQAnVWVT8Uh5ltFvC0UBVo7i5v8eq0U+SnirjXlhoOp0laS6fPHUeUm/pgnXmOMscYc1i7uw
Q7DL1k84E3kfAS9XA0gURLnXfbIPqm1M87xzCI1c9Q0YYQLf3bHH8crCrgUktbnzBeLAfl4F9bz1
yrLjvpNkTPLR4QI5FxJ8YReBbWwwvHw79rbt6n87hvdq1/JJOmgWnOTTLkGP707hi42iegP35y/B
PxBjroETvYdqT2fDWWn1lWLTPV98sgDP+Bt2uL16CMdXAE9VKbpYNk94dhv16U5gYtRx5m6h6GvR
ngczRyHN+C5h/uiigGoPF91q+0nGwbc+ama8gLzX+cnVRhExITU17YDXL1fp3wMP3VV/HOEJGxZP
SP27HlsQ1Lg5mdgLNMA/EqmjolK1FvXQm9plhtP4x3K1YOn4jPnjDFAOyceNbyWuznXPySPfu0CU
1fplcbgDyhyGyxJ1vgVI5pe0yaJtLfy3micfuMTztNOIKmHKkHvu8Ki1dbKyPWyq28W32uDW7fBO
A0qSBaXMzlHLL6YMkuRrKMdueCDwRF164Z3oih5mkX57e3E/bn7/EHyP55e2Pfbl2E9396IHy3vt
ti3HuXVxFcpnMFzxGLop49bQOzU1dmHuJkCqfusrmJwuTD23CeFEfFIv4FraSe9mnpp0C8Bf52Kl
HfMo5DZuIDyUIntZPoDbM6ARdx8Na1gaz4Ox4YNnOiWed2Sizx2lIMXp6yvcr/1x7CfuoQU1+Io2
ip1qtCm9oC9lxsLYG6/0RVrktEti6oZcSIvlNbu1szbx7VvKOA2+xj7PNz2y4m3dPDMhwBkNYY5u
PnKPUGo93vdP3i/s4uZ4N5Ay0s6KzrI+3lSuGhXTorNeNhTaAsDNp/mNnZEAljzP1ta+2AdNQoGL
Lp1eBANsk5ATaV/q8/yUk/fPclNvtCkYVE85I8NdwQmdTCL24UVWjxJc2raVgnxC1HeuLVe8NE5A
MqS29UtiehhOuxdyVoJ3ZD9D2Hj8grT3Jw9qH2AChQgA43bpd4MO8pJWTsqiO228tR2a8fYWzMW1
IAQOk5TZ1fJxx1WJVIIzoI0XKnIyQVqEB7P/Q6wAqqBz9Io82qTBYWxV1TzXS6vzm1PXdMQx+HHW
7WQNLB8KtzGREytpKw8z2ilUofCdtR5LLfu8h7o5DR2b+9zb0wK0sheSi0wvorGC4x4UfzQIg2bJ
fG0/oQY+/7THE0ceCsRgy5YcIADUwaIXRFfjHy8b2A1jLV29wvxxJBKaW1+O4CHN/bK8As8VDLkD
bylFmOlpnC/7FZa8FrDLwxfxmqyWYFpEbvzpO0BI4SsFswDzUrCn8VbUw+xn9miSK4XC3dtPdfE+
ov7+EOf9YafPty4lQH35Nl/MIWDvcNYdU4lofiJVryNIAa0APcppOTHVc21hjt+J7nvG7hHEZyj8
4MKclaYwDZcnl0crpw1trWpYOwk+4LepCJnDyusd2c7zitekymSGkM+sXqiVkO8sHWsl3vVZM7HD
wd8CB799AQ8d6zT2SmB4eVFvwj/llNtjwfM1fNFmvTOvEzzA1yJEN4cu47X2J3tBa8GSVTJb5rgx
e4ms53y/fUQDop34Zb+DVyJPE6UuMLY0rMYJe7Q9ZMyuwuLpA0oRwzCvFJLYWPZep5jlobvJUi8z
5lkgy01vMZEkl7ZdDnmJ/8hKDudSiLDmhBhoXQEr+gt4bGTSvv9AY6MnQKTTwXhdcvE1+yLDdxwj
wv7Aud1kAHgOj/YHI+nKjxHCga0Eoy60EL16gwlrLT+BCpHTFCEeseYI3NyMYQk5g2vwBWQRiyid
G/9B+CxnIwx4mfHio3ZksJZiQ2eaQN8LCd+wZvQmiQO+4P7HtSayEDdhmQ+t/OKgjlXWkphYa6Dx
PuoxVPMQwaSCqLfk+b5biaD2SPt9WLhAqbTHXTmSMjZA6kW7K7LDC+D6vHIV0mylknZC4FqcAEvi
WrWXv5fxiSR2egG7ReAPHJlTLuzy2DRdoUtci3yMz0eDF8mpIIgCsiRF3dIlL5QpWeopNzzcPz1+
4gu+agQWDmd0JDo7d0deO/3MyxKRDDT5O/apzipZqS0ycjLv4Ore1fw9ifrTmyfsq9Ro7kKg32TT
5tmW93dXZ9Z+T/w6oWosBhtd7yXGQQ/cG+raHi8Z2x2vznki0PopKnXoFUEht60UgDzM43PrxgOM
W+4KyWDk03VCcQsrTt7urCWa5077CtBxrlECTDC81qEZL3PVwJPUJSymKQzARVu+7UDYREwhl0pC
uFVw9j41h/kPd6gXwC7jx7OggJjgcIVRj3FWD+p/CKLdiyNCySsMplNaGx2Yzw0mRj2IBfBwp4UG
DYWfYLatvi78MlZoptkFYqiYMm3eiow2RNtW9SJhNHdv0rMn39qrdGYmUBQlL6sUvJhvFXwDYNYU
cTPef3yzmIkL6XqVpAI7h6eNcAafR1NC0Fsb1iFkBUldNinGSwFyS68LzD7mDcB2TkAp+HJA8DHc
aCkWQVAQtmW4W49lthP4mGubUyGyhC5i23jYUXn2Npoa920a+kQBB23J1fEO/4uS30935tZvAEXm
qz8RRGjrE6wrGFYYlX9fSw2sv4zRwIMVYFO2dyYGk56dkbVhPJ7D5/S4Ph/YeZsenEvv3t99eXJU
ogYcazNEzamsiGVdyGcDruIKJ4AfqI/K10JVh3zbp5ZQos98oNK4kiDoRQkGKFii+xREQlKfhqMt
EZge5eKri/5jCa1ZrAfboUHy4PozR6if5f3yKgFY9k+z/8G4udegpsXL+29esSGi69XDE2rMQvjo
2vM9tbTeeXyurkz8nrlUhHzicqQ4kuO3oHLohhoyYWrpSJ2Xej/wP6Kn5e1AKbHJDI+rOWv7KgNX
wH3bboHWR/4ufX24QbmyMrfUtt5Rz2g2EaTt1g66Uo11tVdRpJztHIJLBzLUYAOfjwpYfeaNPRhi
0yDm+ugz0M9mSROQvo8PhpTzGVhXxSr1GMzn+TmJ3swtFY+RvGMKDvre9pPWsxZpSb2sLeAoG12W
sRe8DPJwVLnprmmH8qgnwLjI2lw/M6PM4nW/M61R60q9Kavp1H/a3D6VkUCjv0Jp5bVo6bPlbLTQ
ukDdSuYzT+vidluT0Z5P/seJ0Z2nRzbrKnVNeHvLzCmPg56ombSMmXPFCAXxdoOfERHBRUqR5NKK
3e15UzlGGrXjISYQwXV8FIdJQllX6yHW/rgC0q3q3kScpwr0VABlDs4r1Vjo8mGDWmPJBn4poK01
rfI9ZbOdElp61dDXNLtu3XYLejL9Leq3DWj6nCVIFuvWQyfr2AG+Pa83TrRTfIkBPa/kcOsHlOTI
Lqm2GtmYKGknJShkiEkd0BE2Nf8mFsew7CIY+XBtNlf+ekClV8kW8wAFIUGVYo/t76Y2vD+sJmhH
2Y0Cpt1nroshcjAQvBDsDfQaevCUNSq4zcRmyP6VE8FnOkaMmjpV+pHNwTEo3Y1L8Uy1qhxg9VIG
X2a+KZhebEBz8WpwvkPcAagF2GPM0hOCwvrhc5HjoXnqs9No76WmSXgErtjmTTGy3xQl8X4t0jLt
/LzNGmei85y2WBBf0lVToKHPyc8UwXvWGDhMJYmI4c5WDJmR+6JyAULEwe+UI375jOJE1Kc99a82
ereltFgNODtkCoEoN6fi8YuZ8EwXojrkqcPR1354R9Jm4/XTCNt6SRKFmzZ+kfl62Oo8KtkDSgSP
4OHfNxOSpUMCHf6x8Wa8J2hOzDeqG0PD+zdzQSdW2uGcLHpX3+waf5GzS7rogp+DU50dbJ6qgHQa
ZYUdD5u9SEUrxUVd3tpTCSlueuW5sicp5guTHLSrdoOMbHa6omVdT7hZ8MRijgMAJOR8jAQ9gMHO
W/0pi504lQ1TKKd4p4QhI9zDCooVkIPIXrRJXbzxpzlludgUt4H9M5ljyUdi50uLgPixXXlvNCKb
LghNBIW3Cv8s5o7ymPfJaMNc4W6yBMZyHicsfE2xumcEzvC1SroDPMhz2nL2x0K6Lt4qJ4mRGWT8
R1XTmsqw2mLoNKIlZI2P//LqhCjSw4mm9Oz5I+i9z1Qkloz87+8H4876mb61tA5WHORh+9pAbnVH
fF19hm095NmyYyo/g2UEsb8AG4CLTEl8TUZF8l5xGgfZOCOEjB9EJWyzJjlB6ALiC6ZL4vt7cmym
ixEZ2aQM8veOlnDARcm+77SaHB/5teYOKutauFMeCaUs/9UssmFM/i4KUaBkTBcjWsECDVDNltdC
SQYCe5HQ40WJhZ+sGVxys0L+PwG46ALsHmRXCAizoLVVvAUdHwW8xLIvMC3lisuz0ZNJKPhfPAyQ
A00/7MZTlW0YD2aJ46nD6AEGQXGjTllMJS4sCyO4nW0PeTxCRwngV0GUlER04MoOhEffutYPp2x8
a0/WiA2bAwsBPNEYt9E8YojdweqrvICTPMTo8lbC7n6rms2wnPA/9XFQc1ZUgjVSksZqM2f6Z+YA
kRp6llruQ85Ynrhl43UuNUs6DywlzmuQaSm+cdoNJ46Nmxv8nQPGb2HQ0fMHISMjf0ybB0yId8Rf
QHf+Lq7hLsw2sq4+llnZ5ucfjHfIhUa0FqD1V6Wsn0h/HIrsrhfdwYQSTHPPQBrNaO8IpIgQj8z5
meCfDKnYgnB6wESG+scEVKRWTdDbgpVFd92zb/lUD/C6L6LWkhRkyJNzdVRp5gYS6dyuJ/1m7r6q
aMvK2ZdlQs1+jUlk70Ux8wZKtWpmS1j9BxlGvb4oA7kpzQqSHKiskktpBdjvX34Ivh+YfaZM2NpD
/gAwwYoJN3JhMIRBBpViYiT7Nbq4hiwumN7CTHO3L0o4zUKmv+jALi+uCRPnWaaVY0mkPEakke6m
tmnZ/q0LzAjc5eP7S/XDNLOzg8RvlGPBriYKeiNzdnr507FmKFCgWjsmOZeOmeajLvlkjw+yNjqe
fFUcOi9LZYRuFh4/KUcszdaXGpk/rEutOPu64gTFfS3vpCdKhlNls2joL0gScA4VuDsTNuE8ttJq
rsRI40NuiuRm9NXVMVEbo3KPJalufu8xXIzUXhTuEnLNFelsVEKrQAc/xiZdJPwtb5aVY9Wy89M8
l8Q18mCc3MB2/+b98zqKC2Acd7YLoI9JOW3cX6TIcAUYutt4/yQTd5B9ZtPCGXt+/doNFP+Ahz+u
d6/KRU4+bvVwNN5cIDh7V3saRs6qUZY7oywSBwja0SIe2G44JGY56ILHbPacuR9MkGE7g2DMTiJZ
mwAkOc2NbPasnBB8Yu3JUONjSh3TpudbiPHXBvG+rs0wj1Rdmw+Al931miVTqWbcvwsXXUubt2Zt
cnW+u0/nz6LSSdKLVo8/ZNJEyE2Ef5hOHlUghgvTCwC1jqHVVekV+g0M5CTrpNj6fsR5AGfCeYHJ
ubKRXHPm29gKv2ceCiW373FAWBrvhMWc53VVgXTQVkqiZvZkleM7KoU/AdKGSTsH41dSM81R/9N6
pWm1IcVZ/5nQku6fyuo86h/ORzxQMTudC5efzswDCAuk7KXb3BWIiQiJwcIJboRgZV2AdejdV1G7
Uq9MMKh0audWbiZobztXALCjMvNvIYbuxkqeuxVZNWqtbSwU/UWugbgkmN9jj0FbXotjVyEKz9Yn
mEjyEYt9kBk/DgVg3JNZSmeStmLj3zHBHOgxKWEjNwPUcY270KCTHsqaranAB56CklBgBsxgaPCC
0koMsrgddLwm+AQ5EmO6P8+zewHbnb4JRK/fz59d22Bj7GcCitT387EyQim1Ud6HBwg6Cnaf1tW9
dn2UrhDBusJqIdJRHbIeUbwUfTDOBUaFGIvdwVamKf8sllHheLFL7oWgLphuzH8TJHDvNS3IILYM
z7P7h97uo+AMBRqVsCPbQvubUnW3PG6aI2tUic4Xh3PgywbkX7jlTOlR1Sq7bi2Phgo3pUubtAD4
ijyQhlhQCaBDAj/E5P1Yox0NVMSXXKC82EVn+GiCT20J5D/x+GNFxWw64ZW3WLypbf09L5h5LUcR
PfhURcPof9r0TfehTkdqzPHbA1GMYkM9NTLLy+jQK/HkjrXJ0vdYnD7E/PiuuSAoIV2wPM0nwB08
t7femT6dWlJIXBT/kg8BF+oQnEJ2UoYU6XGDxB59Hwoq74QXFse9ShYloNCYoGtEmL2OukC4XzU5
ECSjQBK8clDZ0HsCv/U9Ihf/oqTrNj7u16q5lUfWL6SGC1yZb1FMFD64yMh5qMUoyhIZLD14Xlc/
3H6fE5bvmwnQUqUZ/Nt19FsKTUa/U+Vd7VJOUB14oekqVlnhIbvTqGEzWOEv0S/ao/yyGMk1ZyBa
WizDebDoYq/EdhUueRLNqJl5E9XJd+vougoG/Nl8i7qBvmm4WrRCwLUV/QmqwwO2DVN9pJ73cxNN
OKq/T9p8pza4NnhLczxBOUOWOoMjP1xEO15fVuoz7H3mjohCno2me6rCp8fWNt6R8BwgYg7T+w4x
J4S7/iQr5ymtj3u2B0vml8JK3GZkidnv4mnYgd/gfrNngDNsgzCj1kzpAPma9Rrqm7Z9VawBmtWI
FVBpLje3t9cpy8QSEj822fwccphIqkywfcu5UGhwYQ7hYu17F4Qs2jv1jMfRYitbhdUMD2SIZ4Cr
RAuS/Va60tgGZHgnmyTJufqop1l6gk780vvgtd12IgEK6+4C+OjCKNpKcjfNtC2j5PxCBitoXPN1
UEiBKKROJTwDtoR+KXazpZdr+KvktsHo5/iyTXEhcdyB32U9sFA3wbgOewiYfvlkPvcLcVwLeHHN
FhJluTx61y8Pt7+yH6KmYJRynHi+xAWNwKU387fnOtik/OFgIvwNEVYbK89DeCzOjuXvG4IzlOv5
O055yaIioqDj/hO3WpKksjkMg6HEBea1SbkQApVcdAirpsDq85Wn4/waQjXfvGMg+toY2qL21S6c
OpK1iEXQ15OfH4MurLxDceZcERxCzv58EEiGeVWyWozmGELIUonj0s53QbCJ2nMAN7g4q9H07EP+
l+lduetvBBU76xffyJOdI4AVX7XK8aYvQlFXKpvMMfF0IomLnUBZhRD41ceaXLkT2JzuYnzOBM06
G286usKj48GKgU/egYr0nrmKXE80o5Xsa97aU7Ua0I+Pd2ebpg1ciA31bLKTAdwc9o/Z91QhiHdK
SQPt/vbFWDen7L7NEsDJEWMkeC8xGmmxdc8lJD+yDomg2vr4RnGdyFnB+28NrUSRA+Xo5DzT/t6W
tTHtoswnviAYOFSfUs0Cso09td4WKLP47vYNGXoGjGdhxAvmADikxwSckIBouJSjkoBI8Imnabgv
36RMNM8B3++Rl8VDLTtYFCzq/HLC3CYfRALZF/CNzoKQu0BAJP4bpASE7eLLQ7y6ZGCkSlX9egVd
54jH3bTsfuusqRZtTTGUjX8W/w+Q9/07EBwOZZDnEg/OTkrIck7YqAY/EeN7H1dZwL3s9pAvLnme
1jwzi74MWnj9Qh54husbXqWzZwr3qMX71Z5SoadsHAUdbFVTKWaLL+fVwNSoSa6IgxkGjA1Bo/gM
YFsrqUV8XvAQXqy4x7kT8KOtZvNZlHwTqvln5gJYTeyWTy90dsK0T4SqaDut7MPBxXac3YhwIHhj
cWFIVKX9c2OaONqf0UNKb49zJlt8NwsMlIMwcQ3qyKDZiLGeXirOgxMKQbVO+RCsvtXRgNNHexZu
DVOV9E5HyqlK/8Ss7j4d5hAPp2ZDVLb03LXI/JXvDEGMlgAYD6S9bd+l7pINVwXJetm/VyW7qbam
wJemdE8zBxpkOUcvEWjJF66BsnAYV7opcylIa9MZ30v0DBmdNPR81VVcbEaeiiuzqWL3Ag0Ex+/Y
94Dq9XV3ww3mK5Jm8E5tlzhHF+ZlOWh0gYUiqg+AQ24Qic7EuTWpc6bdAptJCrrl7Az/1YnrtFFT
wd9Le7iuhaivRn75Exz19JiBe4ac/vshhvhyQ3Ove6MvYVGSfYY5+BWtZdVGc6XdPqmaye198Er0
21jvOWXwnpe0Eb9vAMLMcP5Qtc5GWR8dwpsQCQh8S/6fcWCbBAjex/AH4Q3jd/TrBQhWIJwiWPYZ
A8uI5m8asNAS86lEK7xxqgs0dCTx4ZX0Um+x386xNRoN2tw1sg356sZe4ceG1wd+JLB/y0h/IBOx
/U4SxiqQ3TJL5GO3HSwSH7DKKJwo8K20VJYByKzCwKkXbNstkGmmLkG3i28khoX+h2XB/TQMF/3l
4M1l9ftmRm2iT2WyGLd2G00fzQPh8P4emZ1kcBF57dgKtAPsMQ8kJdocqR4m4zE8Ge06GMUItZGK
cuRxXCjpzxj+70WKJ4IRgcwfI7NjU4JxSateWAT/mqVxOMulZfUv7xaTo2VTXya2MvXBcbD+BIE2
10a3bhChAgXl9lReKrPnG9kSR7qaH8ZkE4BKDONoBUz07hKkoldSipOpXaNKs3CCOO+u2on5+aMn
D/Ey30PdKHDSCbxrQzQMHQZo2R5U/zbArlzF6y5kfkcTSc2uZ+0iOSOmLWa7XrbxSWLklNHs0490
Z4A9OKOCedfzAzm9yZbVis6sVW65IRoQ8GEJMqD57HHmApa4dYr07eFwjpki5HN+tVJPqCB9Hv2Q
qlL03fZ1lP9f415B1vuEXpmp2EHhyOppQzcjBTNzIQh1jphYLbq2T8A0f6Mwb8cP4Na3i5qU/ugn
Seakv4jd1/J/05RVzbe6/A7Dap1Hxo1HLpNQub5uei/n0d00Ll3fjy6fxSirmAQ0+5ZFEtjEBSyr
d47d+fV3BKLQjw7ffO100owWtFON6BVQf/QaFs2Jk/8GupfkTznXCmUuM9kfhat6m/MLyOAKru/b
UKpdOyhrZ69glgd/dEpOVIHGd8AColJV/Z7Emgnm6D5JIxuOjRxdgmGwSyrdOrt+/aqfM1t+3NF5
1gV+bUKBzI2ywnjRQZDx321sI4AMUtlR1a1ME4ndrf1odNAsfUlwqAGQVp+PPxJDAsyUx9Mqt2MT
cf1BoP5vmrpcb8CtSwnl0fMQ9//0FYmTfahDPZu86KEkKlrLyGm5utODk390RlpFZfTAGA3Oc2c9
HZG/QcumbKNs14Hh+T0Yu+CroV06RCd2hmU4LfwOTqA9ou0AuZy66LJLEvEB3PUlOFADgepWZvu+
iQows0tJTemGTBNLUqE6sCrMSZ1Ic6veWYtmQZRMX7XqEkztP7tPJe6JqoPT1ECxYluHB2a/XVB8
QsUXShGgrq0It4J5cDYGw2tmjyk1fPggIHxlRywqGQQ1mEd7BurJTEGe5u6POgMqohfrpzmYuPZ/
qz3USwmO8KQqfbi2Jp8K6wYc3RjC1I3QxTW2LP+LkhUOCcdoDfGv/qm988dm7LIkGaK3pU/WViWr
66R4LwZeCrQFxbXfXM8Wnfy+40mtJ9WaHIKHVAN5Bf1X/LEEsCezDMJ/nDWwmhsldFuZP18jP0OG
WMkgflEWnetLM9BCE4dA8IWMW54M9n+4/laLuuLSmiVUSpKoc9mgwTCL9gIFr7lCSWfrFMY/zeHr
gcJqcAcrG/FwtknkTSgCA8GMgbneQAVFm2RP9ckuyFOVYXqv+CpY6tRREq7EFMNgOpLHh1C5QIa4
BG8x11vi1TaLakvwwbFdwIa/x6kCePh8bpQjXymlzcKrP6i1+PsH5lD/ozswKvK5lVakQsWa1SrF
SniOI8XOi/lDPfQtNsGcYb/jqphIFdbyJQ4fM0LQR3l02H51M6m1sEvOToqGlogSLnZx/oykedV0
HWDu+PxcwBBAw0S4TBXFs6QGBwnfU4PdZg0NkAwJxJOZrnVaB9FhVn0IrdozDxC7L7lvN/lOF2vs
KMpTgVPAcfESbZ4XiRetKwAiP5LjdUTE5pookxahy+P177S0pTqF/KZEQlpzSYOBaLKxkSIz4gEI
CsclgpuH2p4XkOCUFiukZXn7J67XRkGA/KYgrJzEJ8o/GPFBNmlAxhTytoFI2widcAh+KdkNCknH
J4ONh0zUMbUAKaikyn305DS0FNSkS0kTcejAtCsx2m2+Qia/9h125OWhNlrfqe5ViyEq0XqK0xOq
QiZV8hmIXTtLEVAvNtmDPOqFAzdXBECQa9ySfg0YnAfzW0ZT7IsrSkcoTEsxgMYdnWw8BhnxSbQc
rtrUCfd14vPeYiUIakg17MJcVdcShZAq0apvjZ4IXAiboTdkDP3aw77trSf/RFXsL80l1b5S7O33
UMqOkr6PXir3k1+K7Cpf1wk12sSYt6WH6LKbJk/IIwZWz388bRV7N0X7D7JGl/EFcUPrcvXWR0VS
Q7bLr/qsPE5lkHBKRT7kRyDOORn65ZybQYPBbOC2C2Fd9N43rwTVghlhpCpAAEdeUwRtSnKwpiMD
h+12j6rOrDFT3eyFSuIxngAZfJ3zXry3EoKA7HAdVC72qTNC5Y59FHd/1m8ebvd0HniC1lPn+x/C
//Kcw1S7blfyg6l4zqZHx035o7a86ZPjxUNCAFCnMWYFg6MJP5QBbESznrv3KHIKXuZKB1ICBPWW
nIXtDW78QhW52ts/P+hdRmUJ1ktpFtQq5mxeaLSlFPXNyPrQcgTyh+aDwXg0pXqxxFVUvHIGS79J
nim2qam9BfLqfAcigP/EFktd1kELdhqkz5p9Dz3m2gZXb2tSCfMAs/+2C/GrTnB3xkhkRbxCNw64
F53AnFttoA6jx2nYeJMVAlsGb2x58nnUa9wVvTtMQJAXQyht9fexztOsY9FqwK4fYcgmFFZqYQLk
C0QM2Mn8N3/ZLfRWNgQiULhHuOaYYBIb4peIRO9iBHZag6oxLzZK4IVT7Zyj7UjpINXe0H/vur95
q5hJMC7KG0tPaGjmFyA4n8fdPAhRXzf+45C8loul7hnOrEdmXphkh3oBIZM1QsrrSuGB8/4BkY97
3f15X7bGuZxFQwjFA59DfFC067CwExpaF9WU0vHmklNW+AMZk1aJzQ8Bd367b1QOMApzwq93RWGs
2RpBtBuvBduFwEK1RzMs+w7deafZ6VQo/UTIpn4DVYYNiL7/X7JJwdBNlY8mkAsd84qokAxoJ9WS
ZPhKz8b8yc34zcvIzMeTEPTSYFX8+QacSL4OvNEk04Z+/LVKZ/daMV4hzDqn/WyIKE/g9Wfe2S2f
NTVnW6YrJNymIC0WMf0A3i0s24TwK/+i7I3dwFh4vSJKeMeQhoRk0zb4/aQ4TuSCWE4T3zHGn+BG
cYxdF57sk29LrjCzVJIAIYMMOZ3ehi4X478vRg40i/r+Vd7TvI1thMLdls9V3qcanA86DvHgix4i
j1FBu1rdQApf29NePZpRy4HO53+dxFTggJraCKjzOa36JGvxY5i6phHygEuEx/K3qE2xqxFUsEMM
LIUI9GCBVHDx7iS6MBdkXWb/aCedobahmRZVSGvL8EIBD1VRs+Ew5T11kh7JDy4JU6Cw8xXvgCRk
9jHuZDccliMo3+fWdIDG36RIWBfzmKFXSXxr03GJXxwuA+qpl/lLOI4reXM8QkVybE7DrnSwoGYW
IzQ+JnilKvMMSSmDmwKCSPQyNg6OOUrFa0LQnNgrdQCjEQu+nh7YIKnFqZMP6g6SCV5kwp8biJ+r
Dv4ZwPNIxoWEE6TSqlm6fH74I5xQLwo/ZQwYHuLyyhTfCi907aoKOJUSh89Wq0ILv5tcHySVuBgL
mbPB4XrLQSdU7A/TQfW/FBmua4oVGxFobl2WCuXw0061h028sHDSsB0+PpvcDOpeJBaAdRMogEKO
Qm32Vvh7fwZ+jRtmVepxPXQ9mjFQdVPTQe7LuUfn+nmcsHfpNSe0Pu7g0hmCYVjfUWdB4GwbcDMM
PAceW6Ym1NKTpkuBLtW6ifpP0tWPy3ITgpU0s8Yu5xYUuR4v7ZvAY0vC2Ne4NSr7tMJ+DnXXlpQN
qWSFiGey1pjGtRo1sTh6XdDq90dyyP+HiUg60PT643iq8KgUlPR0AL98ee1tRPaHtGgX+l4H5hMd
IoS3rUnVW4UPkpT5zHKX0XKuMpMGymprkn6DhhntnWZrbxL48RLRdizin5pwavcapPi/OX7Y8Cpa
75I3cOojoy4TDCM6creTcmDdlyfidkNg9aG7MAwOND+K1raj2X7ouwvaDGzpf8TPxIlnAv/qzO/w
6cEsN4DNImyieueWr1JJ0/LvXZil6irREcZJTWD1RFWWfeGaNzluEaJr16J/ZBWzu3MO566GD4RW
OSaw/hurbkYEup+U7sFrew5Gim8dc91vAfyCgF34t2YSkOnzKsgP0BIAJ77zQVGpP417z6Ba4XXQ
MWjZ5pduOdkyvP3tZouLuNqN7kgJi0U1IuGuD1CZnEzaZRSd5Ka6yeEUeWF2KvDQQmRHfJsP5TRN
SQ1bWSXyGcSw5Y3BJe0z3+pvBqRqaVoTtzeiE0jlRx5g0azQBv3mTPXZHhAodBtE1C2Tdv+iOH9l
eKla2kYjmtbH8htIsIDWIY0ZUX0Tii2HMys4SWyto9f/cBg59Ic7EW0pd9WrQbDdy6Tc64ke0ccR
q9D73SMQF6Cvg5PBnHBnE5UbR9aJ1bDA6eE1O/zx1cVi4lHNo1JEcUAom/NiWPziXeyO991NGnQa
ibmTXJAyQgmReCkN/0HSCC1sKAKwWtavRF0+lQaqj7BcYbR3y/avQSYFG10sL5YSZ6aqNPcN0p8Q
Y5SQe+GtRrD+GY1An7Li1WQbcdOWbJGdaSDCqgNONx0KWd2/4mWawJrZmxDXqI37u79CjqNr4ON+
Ik8/04migv0es4PTowdIQHbdUpYE+qjq1RygAm6IpV09E7xvQ3TG1Dnw7DYsZ+Yrdu2zDvfT+0Y4
uYA+Oz3ibl+BanmOeWB8sb7oSZmN0VGoYgVSf5c8BHJjZfYBUMRdJjLAQJaULuv8ck/XNZktkLxK
9X04DPAV+RY3n7OEEw5Jnzg7MIENJsSolYXDJfiwsFmI0gbvkszrvMMYk/5Q4M85kJlj3a7iBW+9
f+QnGLyKHjQlZfmTiwPhbEth58tEL2aObGd2FCrn4Cz87YvU3jrjVQC7nqr9DyUGcaK1TdPNmgRA
pBLSPM8P7asQabxA9JOyJJaDWiMUYzxNMBJoH38Ia8hneJ30uQsUZrOh2brRfdLJE0OhXipe8zfB
Y+NQOxPTOQOMi6Q2MXr+b2TgKinaLGQl8jMFRJMp8ATZUW0meGBPDeYq4Y6vRxrVpemvg2ZqyNIy
wqUZ68XA5vnvzFAE4bUidpLQhPtjIOAmFJfxoSa10H2nPYTuVISIsBiVtJ0+L1kuavuguyt3tgmC
ved3YzaT8Ke7058jfo6sxzDLFqC9+Etc+hxhBlMJnA960XotDFdsFH6fsuzuUo8JrQzCDaWqZ9Ro
RorHCap1mGeq9/V1DVj5QgdBQ2UwjUYdY1blEkzGwkWVPOg90KT0XKKuvFGea3UpZ/X7VlQojgVa
yBmejEHjh9gNGSjkh+FAwhFEHqlog/czlPqNUMfnVHC1GP1SRj8SmIouPK9fUPU5teyGTltoTwVN
R/Iqa4w/czk8Y5wNpQpSM0vzpuTw9+WAt7oyEo+FieoTcgt0j62jgcBOANYpC/oDiKMae6BaJWw4
wOM3f+cdrgBiR3xv9suvjljjthlaKhFKtGadhWGbfKdexvrUTisaxKUjp8iercOGBgg0fGFi+dHo
PwVF9X6ZXGXZkQzY0T5poa3ZD0APnnaH6inZ/8iKh3i4SlTPvN915JV7bd6x+3oidhZyYBajlIIG
sCI/EWZiFFs3/U1EUZFsPDTKW84Wnf6l3QvBxr6weiPPt3/hNzC6TC4l+07pw9tHADHuZc04S3pJ
6vOUn6NZvILhy1JWDb57y3MrPkaQOKahzhmgpKmMQWAcXxMvStURQDYdF2Rv8CgeQp9Gs+dmQVF1
oaWYGPf2Mj40/mwX4KqH05NIICS4uThw/RPKq1Tn2k4gGuU0Hggf1yRq/aa5vUF02rd0ypNdPdSD
8miMAWMjfnb+fk/+xTJa9/8gHjLi+1Fe7VCwE0qMbUjSOVmHtIP+8yhTfvBXls/Ff6MPyamN3eSi
S2PmcVNs2t0a4nHyDsG/U9m/h4rmuere0ZAAZeQyMge3aGdbmxseVXiPa2TLTNWJb+0JmhLNPdRp
2jS5KEg13AbghEG0jxO8emgQVGtDRfIoSNPRh4nm9yNrY8PYOOOoNcXZByzj3FR6TedEh5pwHeBm
D/IA3ZPHhIRFnu2b25+u48bzNZk5gCtAZuPoJYTn7zAKx0AGfkmPlZ/wZjybcz001fvn1C8K5Hru
AY+jMLVMH4Rd0OAkqx2z6LxZ5vf2nBBZt3//9E6Tj/UhVWT9kf5lUNHbgnDuQlNU9QcZbrr1LQgU
k93KVoSFRii/tQmNxXB8RPLDdAmzymlJNAxAVAPVa+nG8M+v3AbPWRFA0oOkeP4yyflkFldIt7jA
HGp2yNKanBpulj61p/B7ldJRvxZni1j0yH35kzNuBm0fce557ch764Ub4NJj/imjfw1fKTTilgJG
jkiGb1momCIgp+q5gbzq1pkKQ++B2airRjJi5ltp5YuFTnQj880fZkoJTcj87lUrfoQJNCBH+sCR
rbsLwwtHuZJp3+QPo+Bi7yW4N3EWYVmnpCuvDd+hhp+whn4LeeWbJ3LoF2ukikpttMo8DHQwMHa6
B3wiPPtIcflhdeT/9z6DnBVO4ZJ4DvkeE3I3cJLY45epSFqs8w5Su3SMBPk6uYijP/m6HHH2E9/X
f+uAaEsvmwXtTua4VGuwAODvTNGFnMNDIs+5Wx2H785/3RhRYVw7ItuEwbE4+Cthr26CnwbMnRFF
yHmDMsLAFi1+Ft3xLl1B4N6TW0n7P7NrGbV0N9jcS3ksf6i5RjjLqigByY64CtgXj9HHw7aK4SQd
ezaqZql07zt8cZ7xqKXE6sEkaz9mkQ0FortBvFxIC808gXhajVqlz/HSRpOSxOJbDugY0h6to6o+
xzy1XZa6r8TC4inPjeU+YLkdL4DsnIIYqIE99xKtWtNVEp2h/N1IJUFaef+EStPlyb89mGy0IWno
MLzQSnm9/VeeYdxPbJxH693Hs/61V2+ro0gcxwSXZsLETxpUX7a+AKy07Q8d1Zn68qo7eSNNI7p+
24dp2soAxGbl5pqPaqc5epx1r3OA2yxBA4MVd3m8/c0zQZCWNxmq+AaAsWg/XYFGxgVwA6bBXE9u
0yZMnkDOl0KP8gGXQULV7heD3PdPXoDUSrpokW5XkWAfIE3pwEl9/ahzbwq0Nf4wggHRpLzr+Sec
01SHHQCznG3tA586hOHV7ZZT5XZO2bgI5rk6RYauNiDJCuY61SoUlgYkiF2tJKXPHlFVudq0NvR5
PYtcRaI+ToZ/jE6IYqb4bCD+F88ehykqHOMG5200LU/rcqtGC1nN5KHgw/ptggWho9vR5uOHoVi+
GI98yQACCTHaoUQsZ4fkP3iJyy8kk4nCX2nWR3D/jQb1uVcL+ejeInY8RkBCxXzeSU73ZBAtZsdL
XIUaGT4LrE99cRI3EG1IbRNOLzMzJXhSAX/zmdBNgJrHJvmki8DZsw5fIeo9mf+Hu1n+dPYJoS6K
6vhI8qKiEqRVyNchYHs+W5Agr872S/gWAw7pp6xgsqVEkXr2HfTd8XHtiLkc60UxONXoZVXeFedG
O//sCNzi/I1TZBMSRa++0RrOYTPvfbfUwcqASO7zyjXRq6tRv2jGh8iMWkz0TWUUy7EaEJbP/eTE
mvBFAurf8xOWYafYvFyKuvO++Q00CEzNCanSPnglkfNBGmohj1T1fx09kXtGr1qgIHtHCiWv+yfZ
JmNJhhKsu/LAmM2lvGQlqB3terrviktv96K2yQEuueVOWKfSAmJCSjZKrJENFu5a8pJ/VWwWJ9Ar
7pKIkg5cbbGbMv+1ZoCjHJMKwz37/ggWC5DvnFyQgZkOUW1G8flvFF3rYl6ShNjOg4fGdtWNk1nt
Lu/+zPwt905L5T4pJLQxmnzSi5LVuiWI/XsWMNoAHuWyay4F1XgQipu9SHL7tLEROdWppj19GRC+
Bgsm3jBLl6pZS/bKEBRAcpl/sEwVgtA8wM1rORYTAjFfk6dvpdTyh7PdUyBuAmEh+7jgQ52VYAdT
cl0qlL5DxeF/n4UcGeFY9WElaDdkfrdnEB2/GGEj1Ao29pz/IME3M+dhMkQNawVTtIvspOASgAOo
RP98fORJ5XMQqswt4Is1PecaKr61mcz5Qs/yvyau68V2SdW/MAU0kCikHG0vMUfvEgyZAQLe+kFm
eHBQx/gsH4uI+D0HJKBzDVgUZzGorWxiAGPTRLbckVuV+L6qUsA3RFSrqDiX4aNjVaPTlZjkrA21
+ONz1lDD/rEJoSXu5ZBCVl4f+s4eyWu8piFeEcdxXyIZHSip/YGRFySVnj/F+RrnnyLN87Vv5bog
wUJIUFBhTk/Wb3keKRgJ/ZeqwfSctWwixBnfeVF1RYTRX08v79noliORlg+Fc7u6OyE1VWPVHxMR
0eH34xDnjSboylQFma16WT68mne0xlqz0d8rjICPSOrKnr9osK5LIx0TTEgO+H++iimNdiOLjFU4
a5+cvtZ1/UzfzAPB8elg7gfN9nkrQnxVd30atc7iJCGSgelQgOF3vvICbhRWGVv9RrwI8YF9HA03
isZsPKb2OpkIBfa8TV/4BgCIfoU604fRtsZBLuWs3zRHbOQ15sVB5cy14JJANwT93CWDzOhzh6Rq
IkOJIV790d6YexZVx6AhpDc1Clm4qiEYpgcD7QiDIaClKH4eLBCtp0g4bIqAV8fQmGSv7YEhIHE2
SERD9+f04dgvpfZoTu8KgHAdFWFqxQbn0M+BQNp3TRoT5fVj44V1WPlraCEQ7oKyPhuMyYeRQmo8
VqYRLDHP7IDWNvVi50eKk5WBX3XXs3QkRgdIEGDV/fFezu9BDtx+v3Sa+vVg4S6BXTROnukzm4CO
8AhVVeMIey230m1gKu4V/jCbw16/oBuHT6qe9hXvVz+b1JmCTvxqHLKgyyC6UQfpnMjEFisRheK2
bTJvNEry0jATAX/ndFeWebkVMZpTyg3HVs5Gwdr41CDqGcQczwvieTUOMb8nG/6u8+eRRnkjJWCR
cYWICcSr2B10SlUBxMVc/B/NDiWb1VZmsa8Ek3yPeTOLV0h40OSi73NhrIu3JOF60buMMW8WSNNV
7xaea07f1sg04+l0bGZqTgCbX29/XXzGOWy7AZsOQnEQWF5RBWlhF4HLDaTorJGU1roDHCd//U1p
v/h3/Nwe0ojdauHce8/vivrzUZH2h0WqGwNOcBC7z83GgPRPT5811rSMuP2s4S5RTGgK7dSSU8uM
m96A3mEmVIkqNVi4tFu0llbOScvDXqKVTyhcAIzf3EINAcrJ1Yucm7aHCFP/1tkc5v0STp3AZXjj
zvsj1eTDF1LVJ/VrZzLmFs/uCn0ivUjhyjHyZ8d8/FjsNGPj9Fx5LWAZgdUkPa03xsEZsepCfcqo
o2QTZERKVDdQ3UvRNxL1f1V/0ipd7bxc/mIO8ACxwS79f+UlHZQfphtZ2gFlW4eOiMshsvLxhrl0
W9MnUngv5kzEAvT6eFJmo7mKTsiRaYw/EoCiDGUqarSsdEy35qDBijTRFmvqJiYfIQ2cBg0Rphxu
e4Rf+uHaklxGShPZ/oSyL3r3WRFluPIGVdoVtefgir7yVmlt5EOJVNaueqypyUKwkW0NO+LjMDng
0WZcnU00dpcJBLLS9PW4wgkjzvG06jPbUJltEYDQ5Dm1z372IlKDddCaDJgAccLrCzwaDyNvXu5s
mEBLFGZHQHGm/m7JjXDf5IcU9tinPElUSEM3XjDYm7vH5UWoZRt4nLqY4wbPtVoju95XRopV/rLD
rM968+5Pe03kXPzZy0ll15nppjXjG+xlYwev4mjIOWDJ+AiOUJKlDByKHgBSjrPas2wQMSEikHkh
+GsQpUoIrN1L9SL7Cho05P7ChZKxTA6p09BtFBlkxyIsfO8tpQKUr8KW3H59V8qZRIPkIsGQS5RM
3+O0rWb2PMthcI934NJQRw9tmHqVli9avnLq3bn+yOS+f41RyXJ2spgwDMtaAEhokixoHIC84VEs
1uu89C0gu6C2RnEzsmLuhjv1olVF+s7z7c8ccSlRM74aI7mOdUZmAwQhYdYVy2/f1RuIFpybmUzP
N5rDxj5sQ1vSWA4O3mYgaxZ7s6xAC8+yb71huGiyH4hyCB/1EO3U+m+/7qIUVnFE5BwcOEOKj3M7
bqPsPUXK1WUol/SACPrbqcvSSRIkGD+XIHvTeXKDmLXzkD5nU2n0b7+lH+4NpeNRLz/GBwCF6f2n
xBC0PgLEufKPxqj4Rz0Agxx+jdXFiU+OScl9tI6ZmHClO3vG3+Q1LSLjw5M/sjSQ281WZpCPVex4
ThGrxCjc5J4k9NtIQCsVIk5RdgsS+XjVs2mr7b3cLIbzQF32VU3vzqZpOxd+PXSJUIJ4aZzGFS6b
vBhaeBvZNnM6sUMwMn9tBviQwPwuzPJ6tUJbirY8B7A3O1X9njuXAj7C7gohk0rJWP9Xir5qktAF
cLpzhe67ji/OiPlm6yXso46XL6zDu5frxFQ7j9nT/d9XF1ajcfIp+70RrkG3x7PhHcjQfILqa6qc
NiQbHaJWkMBCNLIGmReqMie1IWmddfIs+cSL8Wb7kcP8RiyukhhGC4Mk8SKq4hpJfRySB6nT4Zqw
/goQ6lKiic1D2nLrWzqd9X58FZBYmT4wl2ntch/nreJSStFG4WAwwqCWQHEkW5Kr625gMfsgPHJh
4W1ptIZzE93p8EOMr0crX0LKzh/4v3AZIszDbrZHbgCXBt/vW6EQG8MTI8iB+Q4UxteHS5Gxxlug
vdZyj72uDsa1oey+yt37QAKg3D0MJ3NiTLZo8Gyc8KdRJw73WFcsS3Tm1LPYkXjVlCFY9W+Mgt1r
d+XAu12BSsNi5r7pwY9+6vPx5MOY3UMqT3kK8SvsbwEYYi145K+LYORGuiF5isrUYSksFr6VaCGc
5Rrg0uoRmduH/nZMGJdBFQZtxXT3FaB6RC4G5QClFrN2HaN0Kbb1jwYQ/qAVbnOUQnvq58nMTHlx
yTJXMOVqxdR945HJD8cQocjbCnvluftQpH+EDAJhDSL5BfTGfbgXv1qCmI8g7rVql6IEnlLxQ8wV
zhULAdaUAT6IsQXD3m97NfaH45h5yXj0mfRgDMNmyrt7wRDN2eQoW7b3kULvgt9QIkKgkumwTT4d
aZOlfUwBJ50T1Q/O/4dWgrcMizNJJiHS2ZYZEQolgc7E9a+Bgrf8vlNDKPG9y66RhXrwSqFNTJVk
Fnz6lJvRCIwDxDix6qcmJDPxTRC75VIQ79Lit2Myn4f3P/Ms6zjJFeAV2jqvEGNkTSiyzxVqxMKX
D+WVfXPUQ2J2C1GoKVIazd4+W8PmFy/GPZjl4T7+ft4mlFIEu7fM/6sE4Y6rDHKcQisZrR8WTtF5
ewCf/5OqqcZF+Ot7aPHLkykoKAHFU2G7CpJYVQXler2+/3XFrt7ZZaDD5tlPw6pBmzOfUSeRSaiy
AshwMhpexqB6mx5UYweWEykA7AOwYwvIWJCO3KkjqN26YUmfgdBSs3aqC9+NwBIMqhgy5wuPjJOX
hi5ncHxWIzAGMOheXBijxKPUPx5laLW68qUoTKX+Lf1dnnR75852d9dmfJzERYSFUrXD664Tb7gQ
0czdXYO1PyFhMyF1YB4SSY05TjIEonBpbif76vtQ38bwuQV6xkX7jmrG8anpQTV/i89PqHA2N4ge
OXOKgWUAKhrgPPUCQWm0JUIddD85KBTyy94DFEW8XfcShjVUu8qR+TRwCSlVgB1sccEOO2MBS0x7
LpHFZQp654ay7IwX0KRIyFi6NqOOA9Rf7sfrxM5y67c8R96Aqexk0G0Db6QC/IVI7a/hofZV8JfR
qVCjrWhIvy+Oc7y1qph0FsjgXlALvqMe1NZ6cQcjmKUap0HPBdndgcf44lKzLeNU65qogm3PgX7J
JpJSMSnDZxy3TEy0YHREBd2iLAf91BK21XtmELvxfpC3U6i+LG2nbzKH9wwxt7JgCblGl+uRlbGD
I8RjKJLpvnRj++/m4q4OBmc1bsWRrTyZf0IUKKW0Qpxo033QzphAds/aE5HSSS/QU16j76Jhea2W
xP0JspKWSytekSnStNv+iJDfE3BOfm7W36XrkWf/oyUQcS8JEmkEMFtMHoVyLFRNY1Er6Ns3bQdh
0zLS2/sYkq5jq6VhVNDlV4oKY0rWJz/6Uy2vyRCwc3E5RD2sDfIynLK2mwIJxofHgtDWdeTHLg9d
bJtqvhqCEx5tV/RntlhtDfKFdGH+f384MwowweNMdBHGvE3MwdGcAodb2q+Wphw0mtRp3QeqGXjA
4kInjzCV24qM2NBPmvD5r5I/wbD/GK9iyJLJ2F7PM2P902YK2FXyu2UGIMP/NcJi2LueSLIVZrXx
62+6Q01p8wBdm2kWYDhieRb8i8Gw32qo17c/aUKGBXGXkCxW+9jMZboo0fjezTvLfj9y3DYSibP4
ySI5u6QxkSAt8JHSrwfZo4EVI09psApNxR3fjTsqqntuZmj4iNixbHEKfQ/KVmJLtVw/gP8lERC9
RmpwifqTlw7ZRW8P98NNL0/HLnIpv/06xngH885r5ksm1v6uHswQXybmMzKDKyiNA6yKAVlHDzrv
dx99/QrFf2cYfmLAvlHEJhKLzBI1Gmp4Z98b22MnGjKEoqVYcUp+Q5Dmp4sWUbIm07ZIN8XhP2gW
TvalsoXDE4+5yi/CV/4CGcqZuGQrQAfBf+J6hoApl253H39+GeAQb4XN5TrfaSeAnpQr+ApnvMll
z03/NNg3pUpAv6LUz1GtB0eMp5qaijd802bkpu31d4IADDMO8WENURn8CNs4DQP1cyhOPezj4kbx
vJH63NVHZ/Ffc9WMOakUV0MknwyJuoYsVI1ImMT+NRNiYf3/F79/mLpn0vxivJQK8V7lw7PpFteA
NQYB9jkqg9R2Zhptb6kY9NO1KvrU6v339saNZqHmfRpItR2aNKbwv8/oHt9cOZANx+w7UpYVEyaU
5CylfI5YRIm7Q06cwX5HwWya5wbIvbLGRh0+oG87pd2NxNY92Jg+v3ySFXamhFC+3IKAcm+Ch7rA
beMRJ8EZXwUY9N5Q7+mguVz9AjgIkK1f6MWfYWQYMxWDsk0hCKuJkqmz3awgfMz7HmMXcSEDxngs
Oz+T8IswJMlSoVZxEI6WoftxSHFO+kGAhg+lTkjTBDCsyPl/sA/k7OJUaOoPdL3PSJ7Zhu2xVCMS
aUBJXu3bL8nNK0MtuYQ2O5NSnebdfTRfFwwYtgcFNiwjMTSJIQSvm3/HXs3hPLsKQuDN1GM0B8Au
xa6+6vhOFvQbvKzs/nqH/AciquAHHu7olODFdGnWI56JMRQN7VhAciUqFs9rymgaSd7lDw/qlTOG
T7jWFrAd43lA6HccUqDlCmriCwEn5JcSEOWw1Mz7RvaZ6hg/+MoI7KePx2d4y6mAVwGtKm9nXEU8
eUUyTGOBP33QdCbd2a85U7iIXNj27KP0KyRbHcJ//Ui5OvDThxsxAYZvqyFSe5MJkbIXIQp3+sty
CARCWdLRrd7IP7XrOFoMlTC+Z5awxy/Hmpp1M1Y3vIO4WkntBdGbq/rpRhM4yjb+1c/2kZL+8uiM
bWJm/A5Z1xQ8eAI/bCGAbHYGv70tcDF0PlPkv767dJPXSH1N8xgjWBlTaXYCpNNCrC80vnv92fTi
X/YcNH7NvZsHXnjhlBNKaqfUSt7iPIh9Y199AZjl6ELgkMBUsgqGSWB7mTFUpU3t0AP0zyWmvAss
1QnYNsi3XrFcvTpz/53MVMW1PmuLkcArXh2aqtMNGADkomk2iDtR947luxVeghOyJIneKM9wkDwp
spLF4jc98lvwf6Kr1IO5go0lOxw5W2ge4uNmtPrExH6TxxwQSx504x1o02vKBYMftbf/hGhIWUbi
69xBGTbsCPBJBz88udZMCFwG0rWSO6KDPmG4x1nlE9iLd8Fk5Ihh7/ma/RWrIw/aWQCafT59GnTJ
cUbxsAeQ29ISWqjv4QlPR+f0BpCzad6EtpXyOiyXsM6Dwx9B4ph/bWv1ydngz56dw4IfAxx+c/Be
jHeFeh3fbEYFjVCyw63vjf7NC2l6y013GqNvW8C6L3NXcWCyDXMQ+N9aYq/HYLPsOy1AiIWEIum3
oI0BUNbXyZuIIrN/cf6nZRp5MbQThCs7AkLEyvW5G76EVrfY6r2iudSOmVOfNpElu8HG9YzgVEbm
KjEQoHZKNpYlnBVDpiudFx+pvi53LlZZl0V2TiVwDKPhuojNHe2BgMD7cpQpgffcyX0viA+SYSqG
1jIUK6tAhIu/FfSXPTZlhUuvWvn7E+nOOvyqeOAl2h71WWWfaq2rw5mganEezV9TCUPWpcWEQ7Zo
ZC3+D4Wg6jyavFOLR94pDRSodd4ntyepLMDqR/7y6LXRKseGEL/xql+QgeRPsodhXLT23ooeCO7J
HqHqwHyIVoG54QxTip+e6aAta7KNT9Qv+zzY12wRnniwvzAuKJ8wVUhTJ5xuSjWZssGVzkozigMr
TbC70UgCpdiZKMavBRl53UUAuYBVywm9XEaBK8sAKVhiabraUJJfzdxq6ReTXqLHtRGPJGJ2Hp5/
jOYKHFX1CcrG3sFGP6XOxWWqQ5r067/lrZlvscJcboqSqT4de8Ziqc9cqt4hyqHuYTvYeAZn5Kgr
qDEuchYBa72udDCj1QjPCkGy88vxV42DwsKWIXAWZNwrZVfUgSWAZFYnHkAX+N62gbLmM+43E+ut
PIc/tmIUwlWH/76/SnVj4ZwgRaoGXANMZrtlAM9WluVYs4/lQ/WpTNuShxG1ppByX8mcaOwyA1X6
/8U+MUdBxgMYS26Vtwu6HTe2NYEJdAeaf3BIBW103NU8+MT7HBXk/0GBfEsSxJxVZaQjKtwMk7db
kfr3d64/xX9HHsKcQ/0MDreDXM88F0WMhgorxiW9ZPZ6gOXjYZf+DFzFbpYiVbYyWEuB8IMmfu9b
ROorWcZvzkrDy1bTk2f/jUvU67zgvEgAW+OwWmtbmRRIpbo4g8KuPRV+oggCTlQdghtAEfdraXwA
FoapFwecjdEypyGpPS2s8iXwPy6VTXjr6/LXVPHlRNxjFcuL5TirjQe/FugsBCY3zmR2wFsAJfTm
+F7HvAYrZzHi61c/JcILWCVyWZAqUXAlclofIY69G2ZQjQwI7HvxYtnhPfNDGFPqM25QA3XzvUgB
PvCuX1A/+jwerpU6x7UqVWfAodIGglHvxbg7Mk/BZzQGOM22iOBMZLXAo+v/8Mkc7w7aJJ6j++vH
TjdL4V+E1NsbNoUk4atUodbbZgXC0cBHQcLCfqHEWjxSdl5Q8RaNmZr7r8bpjFijSLAIR7J17SLo
0c+V0Z3+U5XeZE5Fx/mMFBohrMr5oQ2pmqFgIu9UGBX6J/e+/e2YTS/LGzprpvTo/yYCbAnfYF4k
YN3SVQ8EZW/RvcyeEXtUPpfUI5DSBcg4a+mY2O3/x4tzwtKV0x6RkcifjHaHwm836UoI5Z6VcBc1
2KptrWZ5IZ/Mo4wkWD6csAffeQrrE2xmoGXBKQ1x+xkRSXPaCAGMtjUafmHhm9KV/reVGparkt9a
2uxcn0W/Z7l2Hrd9460o+N6XErds3xx4qtRHnqB6vBcKMbqIFL3gLPcH5uhetJAaAttyhLdFUKAZ
OR8W+N8rtMcjawxMuMzlEF9Z3KyUNLOd4NIARkdNtXOGgzp9daKvsclTIY9bydEVp/c/cVR8Voo7
lY4VEqk74MF4fIv73AmmctS8rpqDD3E/ApEyubsITgdpM234K1uyTBLZDD+CMAARAuefy6KaxXrr
XN2bpOHZk+VLKsy226RfVPRE47+D06sk50fjq9GAHemumsAIr6ai9X7xhY2jgVXVnQwnnet9C7Rp
q6wFTR9TEI5Vn42/wbpz45H4zBruzHne4kO3gz0GEYdUNnCbyvs5rWDQQ+97ipRWZR+Vfbnn3aNN
4fXCKYlwJJgLATAfUMnIctCRLo3hrgSB8SGmKGlpvj82t4Yf1X7f8lCQie1MCeeL+HFXanDMlTzA
MyB87THS9xPxaKciOdZa/aEzQDlUSRwT2warLY73WYxh948KljtWeCpMv55djJelIwuxeLdgS+59
qstmJ/NZCjVRiXhTIUld9+LP/lR7DO9GH4yz7odOwN9iE6fQ+zRUv6LEGzfDBQoyMEkFwM1xyg32
wa/blCJYkqSG0FrTHV/GO0ivpCGo2ksUBY3reEFxwKdK2V5Zf2KgNLuFDBpDchf3vE+Ct5dlnvj9
toaGResWStRavt24PjG/a5jrL2TmAFGGrdeH8X8NCVDTIZi0tf5qu6EoCVpTrVkm/mdqIAa0Ulsp
KYJ8NCxI6+kyO4e3NkiMJiQ/T38vaPi/OROCXVskHNKeFSY7cULb+QFSXjjsd+sVaKwmHtxex0yT
A2VXITzmkyNllJAfZxs5x3zrBbvEOp0fcLhb6a9w3I31VkEai1MbsNJN6HKXL7wO5NRfvI4M2vjQ
JWCZFwldbSYjcJKeFqNvMcXS0ahjajbf1x13eFMOJKCi6igdirFOtvPEMaczLlykBANKxe+aMRJO
2wYz5OMdY394XQ6J6FSlCeJlZn5AD7u+UYpviX4xTNv9KWlUgr8pNRHZnQ49lYdFCYtAFIiMbfji
UbEmCMDeCDDYgXt9kxYLgE/zrFAOp9XUz1tRSPHD+9w7ixwaqVL89xMAk2rZeewjiJ0fSKQkszFz
v1PNkC05wPNaY6UcxzLDf1Vm5OpPkQwo9XDON4PXwXoinJNvtWJldRnbVtUCQ5DJU3aFhQD60nUX
b2FiP7/Y18LzyYT3GpCIc2UkzDakEeGBVK4k7WO69mf/IjUANOZPb9pnOPe0YVkMa6sox7RUzGBF
s6mqgFFs8/MS/cGaRcWV/ORhREpFfQ5eISxi0DeL264XRkU2TE6/zZ9OTItY/HzZTuwIV6jedbDI
29BjDyADmJ8oXDeFYXq+JP0c2KrkO+9Xuknbi/IOng+FOY1D3sSIw2bSVRyXwRvkXLCjkAal5J1O
ixO06uGO0KSwokbzI++pdrLGQRA7zM7nlvjQzv2k2HvtzHDhm64PN8jHD5u7x3cBq+t8DlIf6HBi
weTLu3U8asF0l+F9jMriOQNAybzWzEZ81GyGzIqhjVcA5O6DcB/lDn2vjeOBiS2Dtmt22JSqRUxo
K4L6cYF8v+OLiGjlZ6rUrPzhMrDm0QkIQ/bGdcwEcyQfgmbPKVGLtjYl9QOFHcvKb8eqaEGBhykj
UeXJdFcJMx/j7SBODlQR769hHWwt2Ebrw+KN/j0phjqupsiryAxCPco21XAPNDywxKYGgNS+FMwL
c2NR0SV+Awq+doB2/zEZm/0GcOuWX2bCctJv8ix54avj0dnSxPzteyC7Bk0xVwGnCvQlOu2iCpD2
5uTyqRSusROpC66yfan+DWmPCi/fittCaZ87f/0rd5t/qtyftAqWR0tNfqTklOrmS5mSvg6/RLt0
bpW6oCLhE6b+UlJP1EDJVw0xkBpEzu69ACdxoJHCkVefqL/jdGEz9lFJ/U6gYKl9J8fiUjg9Cmrw
TyFtazrNRPYufT8LlFXZ71QIUdZETyPB3oGO76SDekXKzaoX4OxcWYKLBwdT4oJxt2EOdZUCGCSU
QTrNmv3e6xh1O19pWz9QN37woTlbtuITRf0jaRFbplbtppaK2TzMzqIoF06qqsLfKah81Fe1v7Ia
Zs71P0XXRGS28qjDE5k3iu294/79W4c6U3EBdoglLdw/qi7iKV7MUflOOzjn9AyHgGdJunOVPfZX
TjGtEbGJBnwqG0YMLSoI0qT9hySdFOLakt/+7HeXhFzJT5AfK4qGVCX9bRK7fZVy5Dpar+W7AbfD
5CUHniqttH/rz29qeQUJaYi//A4WwumwFPWi3jajq37aUC/gOi63NJor6K/0es4fDQW9OVhmdJE1
zgAaJSQe/EgW4QjhpC7bQZPS7aZ/SF4NR4pr20H44qUos7QFWS3c8vFA8R2m2cxkUS6BEc1oyLSl
xhzu0PWdWVncQ1MgK4IVbYELxNGS2mV/PaL2+0a/EC7r35l4ZM6BqeAiO51JxwcAbK0dPwMeJ7IM
A/QFeAJUTA2MjGeX7CRoWdtm1yTwIsZ63/THhqim2qx3Y4nh0uOLCIluDXNByIkOQtAPy2nlc5LR
EVRYUbH2ZTq4XQLEaemHUFEofhnqC9YZeI2QIXt1ZQT7DPqIVX3QHVybaGsRsG1vvrpXri/6ezEl
c1nTZTP1javJ1K4owiMJ+np6TcPG8UrG04ydjnlMEUIwNY4yKjP63iWebbCFoUIF5aZrilCdboTt
gt+ihs0/kbGNvYUkl3v+M1wsluMY3XL7Mb6P3mzCoY7utbWppNgsuC8I3qel4cDRpJ4ezHcjG/9Q
JGM0rPuYWmLKSjF31pwe67ezcjvpyhTAVxnkFEGHqJjrI07K3Jw0nT7amFMEZKRm1xY1NhKRvkq0
j38MnIZ3Nt6+ofMBGupXgI8BPfSGr0z6syVK9iKbOw43tZ/S6NDJzYp/BHiZZ/H2+dH8CHMT7Poj
Idlak/ISmtBSgc/IqQntcVoGo/c9w/FCRArhyJVRgLy8YNozPlUKmX4nm4z2qM/54HZEfr/mjELj
UALQjmUhT3B9Pz0ZxinNXwfCVW8fyi0Q8lCUKUlKWq9P5LGaj8FU+73YoYSA1nDoU5u2JXgODTJi
PNJ5xCF+xo0pgE+GpzlOqWQ228qMh3qU+l6YOGxz2jO9VBK3R4ZrPE1fjccUqzQ4NUJnz+Y19R7J
DPR9HqJvH1EtoS44vN2KaUTn4w/PN2xDnsj2iBqxzvuJbbjtAWRwrzYf/O3CpUV0CfzdxcsXGISC
FXV/xRX+NmY8GVsFZ06OYaQcsmegbWpQQImRxiAoeho+hWN10/9FauPUn7fXQl/YdW/HMm+hCNlz
Gdc6C2wQh4lGYj8ofNodss/sKonpa1cyc5deFAGTgXK5bh1W9RuSHFKk0ibEZkr9llgWV6YSxYE8
v9SqhssUZ5O5eRY/vQW6eauHcEyVHLNx2xJlCH+nJto1/ZMp/BhglTU9BS8/g4A7qOHylPgN4NzC
a4C5iWY0yNJsqShIy+Hgzdl5vd/sAFfLe3H9JFo10Afmhr+qloXvlOSbh5kiAz+n4ryzVi46yZsc
cmlosJ3YzLgZ0hMa9Jn4JuyWdLqJyOrmLsd3HR6PafRSnTFLnTeca7Bd+uRpIO0K37vIx7PQLbg7
Xad8M7m9L97X/tTEhy7SXXeFqGf4N/QKJdMGhbhSRtkYgcgt2PHTLKfraY5LpcqFgQ/eUUDV1bvd
a5Y4VTBR0Befsbfvk0b8J3Bgv4x53wSXT7SKxP/K2xQfTK2ZEqkeVl9/zEIJobcqS0ngA6T+oMID
Qo8RC2rNrvE0WHkXpTQOmgZVX1hH1CfVjrRU8qM1typatTfXAS8BgU9zkPUEOLOOdjDAQgcPYAwI
ThHW6VYab9VqR8Pa4kzCrGN2w4HGBollAeG4RHhq0V3bWaE1e9KJz0jZBD+CXZ74llXYrbG1zy8G
QwJffAZ5hFfqfyQQEGhkjSyY5wutgqyoSZQrN721sQZug5qvwhYnsb6e3cN81s9X9N1ZfchAWZAh
lgkqG0sBD/XMNi0KCAT/OhVJWhbZonh4mpu3Z+UyhK9o3f8rtXXEWUIqcNVqVgJFqkJLJKRw35Po
zeM5GRhpd1QSC7gpDaivlBm7Wj1GBW6RlUUkoQxGUPegnDNTo84BAfnixN2OdBhhLiS2B3i5aK2G
rGrnSEC7Qh6uyrRWHzdozKfqwMYI67R/Hz6snLjwcSIiPZeVK8SYRI2rc0LEILiqbbO7SEZ/VEf3
O8w1jLhVanSB6E+Fi7PvqVko8rz9EwYYYegYyOx/pHTY7gZW1cvehemODmz2PwlbnouDl/5iDXaC
8oH6BP9JGT33aN++xP6eTUzCguMQjQCGi/lVf7qdG7qEhj+kq2AdpCUMlkBaVybGSN7gtPXo8+fZ
t2j2BE1/DddO4kFNaVWVtE8+/MTsXfHe0MvHShwVSvnfnhaBM3n+W7hiAEQIFdM4ugGqc/1U4GIP
ktyD873Cv3y7l6CRT5ISTI6wkLAnETwk8wOXuVs0mYL/2eUWjiH97yov5Er+61rj6ea2tKAKICxO
KZZrcHYwfVhr5NETkZ9KOUYCnoAmgsR+wWRrXepdo4euBAxgZ8fq8zz+qP9ytN1TL4DcKc+4VJXo
lmFyEqFuBIFHZhQct1h6HJ7hYvhMKxNLMKQ/yp3Pv3EL01alRNoX25kvioZ9yX8KpdH1RTbva4AD
BCdSGtxTE+TaJLB2bf7u3JkT3jSPVcEXBdRRyGd313epB60dwWZM5xg5HiFLLvOLyjGLPfs1YcLj
yO1VDRK7PtyVyzY2GA8kezUNMlUxeUG6jGAvRofQASV9mG9UFAuB04dwFTPfMkMnKyXS11oYt4NV
7FQOpVKmlBcuGoQMjhKEf4SoJAZhThbDuTUvGN0Xh2LD7y0x1+JonM3rFBHj9e7CFRfu2VmGg2Fo
9PAN7bgCppNacm6Dhz/lsuOvD6xRgIriP1M5DpqjeMb4G1CGRDEOImc7PQm0O+pg3XASE/laRKQt
uvgwb24236W0Ja/ZizuzAKH3T3quqpiGZ/nE/Xt8QRr/nsQgmLVn/4/246QBR1lz+gWD2uaKXwL7
2bCwLWoPPQ8CdoUUNT3ELsSHkSGt3mGwGb3Mz4RnMsa29FH9sjQmuhjqiRmnyUIOG/vDj17J+UKP
56cFFmsvRRR7lGkD3JLSOhlb1aV7DeACw/Pp34QUHFwMuuz+0R0ciPujnvrZSphAVFfbyhPzaYkf
T5Ghh9wOsi3REgEWKZcslAC50O/a9VnQVuHFF+DbGIzAuJS3Wrjhkc6R/zsadn/+9cMbFQbt+FgU
Ywab9IiyHKfkGyuN3ATnhDE9TCWr/m2RgOxFcFBwcgWUxBiw5beboAnA4gqI+lh/yc4VDsjjHBue
Bp7ixYBD30o6IpKv2+8CkgmPvJOhjrh4XD/GYD5KL19v4Avmp7GlrzE/02ita89JmZwIxIg/+dpP
jXRLQg2nDFnSzfpVlJnYbw7y4f3G+a8+TQG3DKLCOnwG+csaNqNEFPwtlRnYliHAYbaRx8yWpCRA
qEBy/nFR08lYE+mKDAi292o8ehSiToEPX5gB6HrDHitMiR5KB8GPyC3uhxVMHiIwmmG/OcutLGXZ
RMN4Qpx9u+ZMzQMLTTe6VboVuiWiC3gHP9ndArnvNGGj9d8pXY6DUfVMXBH/Tj98FH7lMUmQrx2u
xvJxExkCHKO2n2IB7vrFnioNhzchoKqtGEyx+iVFGufvP/jlyyjAvRDsxxmkpQqTFiX7CCwgtd7x
luNZ3HjZCp9KYEeaupHMJAJa8LdSFQfY6mE6hg5frM0OSPB4WKPND2HXM8OIVkDAHm81MpTcytrA
NzOg8vmt37/8RM7J5qnn3dTx/p0uPAMR3K9WKzcj1SnxNSw+qMHjAZozNHhKMaFD3RHoJDfevPx2
+82CCzMhqU07xnko7K9OVT9xg8M+PcP600138oV5XtrXgw8nYKn7kGaYJhok9ya1Gde02DvjYUOK
OTCBC6p8pieTuZ2i1VTuX+T682AcOv1WQcQDuEuYAPXjqNLwrA1aB+fBB+Rr1OXMUtXICjmtnJzU
R6982r2s9WhhJj5nKBwp/La62RnlQE+HLJEmPMdHfkyFf2awwtPN5axtcYulva79SZp/YkVHitaF
EmXqbWU1rXrrfDFIOMc45Z3qT9HmXzzcTmbeQWtPTsRDP7HiFmh5HDz0M4RGlIvt7gBrG4qLTr68
qEXDPBfWVqa4+BcEmldPXRdfj0F/Xym3k/5VriluxONeGLyo8LyKXDVrIzJVhwlyDU6jdnwY7Eun
x8o/o+CQAoaRDArH/3x/IOqAKLd3MOvLTdFEP0ZMb95b+pUwQ9SCTu2ZZZgdZYdVX6mgZGnKMiOd
srhZFV6YcpyR+tDDHq5VLeoi0MOxyN+SMd/JWbeWTd5AvNUFtBZPvfL7+8DqAL8CU82niM0S3p7d
PIvilBr2UkmlZ78GKdqBPCD7N7+EorGZWwWG+0/leTNyxFA0yFId9q5FtqrgNBZdcfMYnLQbMT47
4V9vIdvd68FYrdK+OjPDyiVrEeLyu3j7FOQNHMeyaC5K+pXXuqCoMWCcbg9TmAL9xi6QnbyzKE3M
IKgjnj7hYPrVsHj/suHLvfCqoRZXGNIfd0PJXxiUWYIH6XPC1h4PMtQ+BykwROWJxDidzLAvwsXj
dSc8odE4d9McHt+d1AP/Mo1OTyJfzZ3F2P9z9O07R/CgB409Fd/cGASY7+McEXVxlCoMi7yO/L/I
+Vdrf9U4+0kDjjiGNalsRTl2vNpuUcjTygh1oQu9jjQopjA1Pf8x/nTaSQ0i4Jp0rIs+AfDMgTaH
gDZlF2553Y4cBrS5u+3AZ8KGQX6VGCI13NrZSsTKtOaVsCumOlD9hkGoXSk5OtuP7issJSH9euWN
/D+U/0pSu7lDiN1u2wwib8e4ft9y761VqIl/1bleRBF4UTEmKaED+9HF20fw2kL2+4SnBGMPw8os
bx7ClcDrk0l45neYzhtKLwl6txZxmYfLvIEY+g58G5mFIyK7XGIgTpQ/ieESC/XMTrYsECxMLnut
pwhpXvziONv72p1GPYD5ojSX3IO+CKPtaK2bpIdHgM7U08p2OGazo3+TvMDN3PN2M7ufRuBCI8EW
bp2dZ3GI1jmkcq1Tc2J8tbSNHeTexSWJT2ssI+wz3iXksysLM2Nj87tmFT1l3UWAoHVSKQmvK/0E
xIADfNWuZfvt+x3vXswvkh0XOa7vgnr0erdoE2RuSbh7uYYzBMgfCc/aKq5IjKD7uPyMzSTkkwAU
hNQHUb9hYXXERyBZe48xyo4+gEk5JdltAssXLUXIhWqEO/cSv2EzVPnRthjCyoDzSExvSXgh5LiL
bNOYkRDH6NFboQDkCMDUaEQSf3YGiDLtGvUuKFogTWGHrA6ZaoLTt0DCIr7j3PBla78NzN8LbsRd
uaZmDllmYLllLaAMB3hDc0kShLxysgQIcQJPBR5s1Hn+lJOKMPbrqRskn/3h0hMiUIL80YSuEXNi
1WCOnONkHjz7HEjf9bbCDAuZvhd/QvbJUad4DZc477X3WxvIyIjyPHfWAOBLz/mbk0VsPxV2mmtK
Uoe1r5X30Q0wI6hD3Rjb4G3xnnM5EvZ4ZmZVand6VNTVygSOPfBl1HuHwjIJt+a4D4el5rOpL4Dh
KgT4hVQxc4e0x4piNzVz+7PtHllSxasExdRDo0yprxAcwonv1nAD4Dg96b4RFrsc1baIbbCRhiwe
JG7P+qevsvkFKMeiyJ4tuihBn50b8gwlEMrtnf2MtsMsMNuZJG1rAmTZbDWefAF2V+mouvLqHbAj
INU1mIGumxW/eTSFA9Q2gzPAGSlg9RQZGiDtPbg0B4eVQkVcJjl0K3ocTK4Sbhq70bzTMWlo4Qve
Jwov048IssUcJsKE0lN0/0ODEZ87Rfb6y299tIefamR6EpKHF0YUu9mtjcGwA0b3ohb1WJzyg/a5
mLcLB9Gj22dMPxm6aQSuBCA/IEZnZjogWeoI2VGMBOqgHV6cntNg5U7tHuuQH2Fe9hs6gSEKF06D
BTHezHBrkiO4WPx3InjB+jjJD9CTgduNlAuZCTzHXKcm33dVhWz1F9r4zyuQJH2765F2higsfJOl
7rf4Q2Y18av6rLdo1U7E52reeX6XSx9ksnQR8kdVp+zENQT5kQIeIQCGMIgBGGd/v4nF4xBIuSXH
j2kXlkyx+zd2LOUiE+hoqtqzQShwD0XjhXJoJdl/fAgOtgQ/L0opgihVcTL80nTOnTPssldFZYJs
PYPu/d8LuxpceaamcIh5dw2aOMpfgyfJofA+cknNm4q2t2A9Wpy+H2zOskgwGBBwlDn7NmbyYjrl
+8VWGFm09KxC9+bZByH4L6CsoK1Bc1C0M4g7qIAO7VuDlQQPBj7Js02HoECOfQYUi9C1c+zsVt1i
GgWoi5QuXELKRDhKfQsCWiEH0NRrygFjuTKX1ckVRnDEoKhqpkdNUF6J8hoJLYzkX02wG3h2vf+Q
HR3lkX2HQIw5+5QrgjQzNm7Nm72r9XnY+cFE/KlWtcawNoXtTsvAGWphPmOdY+pHr6JjUZZN8DxY
wRfbXLh8UAazk3RfE90bv+g4QsIG8YAHhGaTxubG7cijcNTFX189NmlOJaVoSpIIr8WKfnhnIkqf
fwrCr56ZmvAMhzKSVIh3ax4CqHOtqgVxQB7GTlYj+uADaSRMnfC4gHnY6sNGQGxJAIPOeYNUZNQj
r4N/8/RV7vGyGJWma3yHJNjPljoQIL+YbhLUMyMHQlAhOo4ulhE+pLaGkmlBfsT56VzOxKPxV/Mw
fFWa0fMTpOBBP+B5ScikdFOsOMI2stdSAu/B3Us/d7eptzoaS7l0KiJWpDBk1m6fpgmWtS6PrA6Y
N5G04kGssujHyROh8Z6qNReIWBOdHlszMyAzsdj8U9i0S4M8u3js9T/Xzn4tE3FPPY3EmBvN2vtT
unhRds7KtJQla5IPmNMj8jpOm1aV4vXRVRy0wxhumjbIaxIPac+pxRIoQ0ZuAI2Trwl7Pg+4fTjB
imzHJhV0EUVQy+MEfuBa6kQfWUzX43ku9njOFdIXDw5JAEQ7TMPVthrgM8flQIkK1G18isVb/t/x
L8Pc98zL6ipEBBNwyTPpNViGw39qXCfnVvTiEC+Gy8nUP2DAPMKkrf0J0os+MQihhsevIsWqptJb
MTZxsACVDEvKm65XDe55tGIPx6OOfuwNPTk5Ik8qyu4zGfAUjBqIKHVZM5uPUVYydZKUwQb16k3o
XDVohZoucwm/Ga6EiCawU9usMmtO67Aob8YemenPN2BAWXQkSMKRbGZXqlZU9FShfnMnJsmvw/WJ
1qSRVOM7aZsma4vOEFFE6rwimnZvJD4gATGfWGxT2RRMovLKzj4hZTRKuY99TDTojSx7SEEwlhp+
UTpIoGOsR75BntCEOcrORixSB3xnMuu1JCkETJhEsZd1UgH12NwldyOyuwTQIpFfVx+gyWsRU6o8
RXpBzaOAauquz/JWXODbweVRScRXod+Jd62gu8lvSLF4HxllEOuwoAed+PTGKg+9vvCq7chFHd/l
fD7a01fwHsJhaHHLGAMoxzipSpu4qfNhdBhKwngMWtuXHP9fbn4Qc83v8KvIv9f0Mv6p/4I6q0h8
7o980mfW1ct4yYLjiIfnaDON2Aa4qMUJ+a+Re0bsFPxRoudxpjoqBTBV+6tmcDJ1cqkl58neaj2A
PnV6TyCMcu26KSiUaDUwW/8jLXKHv+Js4nVFSTPbKfYkGTq9A+yDP453OM5cWbyko/zLfbYXF54Z
ZMGU3WJQvpCIKiTq+bwlE1VZ9UYvUZrxFzYQdN+o16+Es5iPmbpq8pPXP2lvuvGaxIDkK/xECiz1
94nLo+x7ktihGVYGd4pheQEkVi1mzXDiBBdMaX6BRgzy5IyZcUU60gJ/uV8A/0Qd7PmThGp5cd+b
jxCTyvHdGKBwkyNJRIJcA7iHsl7jIpucZ5aIT3OO8dKkoARPmC7lC6HwnBkqfrzMUMLbkpN4YBw2
xjDSJpw20vrPLB7Qk+pDhlWMmpSLrVqHmeLc8W082PYXml84U0Kd3O2KzhReziQMveLmTku9QrJQ
T56KWidGOGtTcGds130D8PPQG5y4JQ299xyJovYXl04HkXdeKa1pAsIcLhWsCYspaUFe8lFQkVnY
jHmEkmu0k+NbnGw1Zv2/pxThBG/lFKvOyubvAf8v7i6bV8iPd0xrmXJd0dn7yS5vHJUrbIej/QZZ
R2URDYhuxqFPwxvOtzBHod+Hr4Qu3gNP/kbXrO6e/1XJMB46d3uSY0JV3HftWH4ToZGCmi3ceCnR
J2H5wk82UuZtXChSIfD4H0ceq+ZIlazDU7mTj5xttgwAKcDkVf4ZrWqMiX00mxDStYx5NKhAtJ22
uDz4g3+VwO4mWM9yBqQ0XXFDJ6+vyXLoJ+f5TZhWRCVJCAbTo0Og9Zrx9xpA7Z+vlVkTUWBXVU+9
9BsAcklK1Gacu1jHOE9v8YZNaMAoxPfI1ne3wY8m1xuS3nN/coOXQwEHtmkrUdnyFtXTEjOXsGyy
FaCQIvdLOD6Ho3FNEVjQh8jg6FRIbKNVLJBtxp/fpM53Bc2n5E0QuV35rGUEp4qmrDMpdsGOXRMK
U6bAodQxMRhoxUmZF9KIbxJsgaHerzhe2ivG9irBpCJB7OBj4Xi5sPmt9y82Neg/0riEoBL6P0mJ
gv14ZOa6rKPIUlXIsJ+s7ODXe5zk0EfVSM3fcLbEO2TrOT42xrXMVtGr9PCy93OD0vlDY0Dk1utY
m3o+XCcLiS4KNmCLMHYXzR6ZjPdgDBZI1SyvMGRosNrZ8yBZT3Kafb7lekEZfrqcbkz+kLqnCtGQ
A21cNLy4FoNfkhHl0Jl2te/N60GGYfVrMkBRQse6mJ15Z5bcgdHQ95BhemKKDObDeQNupJCxfLhD
969bJp0bjV5pUnbPzhN2qp64xhC10u4t0q8Vdnq3wFIFSx3Y/ZUzLvyh384reppfTazzNfmAYaF1
BKN82cCtSA6ocAJR3/1Q+5uFYLCxxClzWbfBlcjhCbjabbyyKd99fzXsKEfO/iHiNnbBFP04ym2V
3WXzQtwCNYbQufOf+7SE+/ZzzUuyUoYMiTyyb6xTXas65sdzw3vjv7u2X91r+FOFTfgJFFIwNSX2
rE5se/U9qgxjppBIr/t3xJCZMxZFFOZ0Y2rgDC+pig5mCD6OeHsRUlxaMe+nK7dON3rRs5Dp4Tc+
ovpeBGAEkkX6iu9KYe9MoKUl5tljptcmK8OHrntAFXiGRWsaRasxzm/l9xex+QkcrCnF8HMP/h3m
rbp4S9F0B3BBw5u3YYbXdBfeRkQPRzmgA+QGkeDUQVPlq5E8Jx/omHa5j62IkJuPRkvoFCE9H+qt
oIALBDdzFWuE5tXIxtq0HUvgnsMGmIebyfPdu576VPjlcyTL5mzVZVgPWMY+EAOuRVG2nuR0opek
YaP2H/MOfFCYbFQ+VEKAJsQX9cXOECeQe0v1tPMXe4mwBVniFExwHi6ixK4J/MDlEyk4IB+rzJ9o
9ZRH1/Vpq6H7zshvv8XYnsVZd/jTAq1yVxD4Lou2Gn2UOlh+5gabYKGaPE+JF9IJI3mlOPCbX5rE
DthJTa842vMJ8kXBdyCtnKZccOl5vpzuVI7CqcdA9BCWGG7way8IWx1OSdRjts1l2YpGhEALwwPp
IQ2V1ydGP47Fr18MDxPy1EPBKUm4OVLp1i1QNh2HXW4D3DoW0Hkp3ZonBwrdfCcoQ/1osTjYcbp7
lhcFV+QhQ5+mKOMAsyiAioCimg57kP5gK46xRCFzxQq8mBWbxnKH62M9irxtYwpYoF5krzu52s/7
VjwY8fqzX5jAVv0hLi/ZHqJCaTYBmQ37VN0IpIxDR+DdlWI+KVWouPCaBBFKaZNlinKSHTMbfvx0
2ObfQdw4IIMMyiKNMQtbmg4uoRZK7trW0zkPbpcuMNPqhErMWiVMJatAduZeBLXZ9sUzEX1XDTnU
ckZCDyOnzuGmWMVTJegil0ducCyOCwjGJEuMChPMOdcuWG8xO42GpZJAj8YOyWM5n1t6qb/FdS2s
cXU7DDWlI18yGupaJvyGNJlwhbYgMr7k8OtXOQ8J/4GCliSomHezdrTiiOFaG8D88ZkBpKXL+D7n
rFthknWTJBQyWbbvtKU7uetsqGpmGXCtugXcK7H6rjAox9nF/VlqdAda7f5erDWd5DpTizAmqv9N
ME3XMA4DsXQ4xN2TgCvq6lrlgzIUbUuqsbx5bMvH9azqGC2vxqS8YMIg0mYobuRf2JQb06eVK4Yy
ZVc4k7Hv9AN6cDV4m3XXJLXgI4HNrNW8pMr5I6x9JI4mTztznunLVCPBRFZBQDOaly45z1EQPm9N
DI6XqH3TQ6PkKIqX+J8+MEkh/D/3slQ4AoMB4GMu73Mw8OBYOW7Q32yM69MsRUuMOxfQVXpz/QXx
Wzg9SpjLZS9FbG5yW/2bIniluCIwD8O1XVRs7iHQShnMjWLynUZPNxzPco1+zBCUtFl4BA0dJlkS
7YB3E5hYPg3cIaWV9VNmjjzmeZkmZzb65B9NavkpaznZPmJoU8u6zM+oH7TNJTOnyUiIvC993h5S
sQjygpxkCco6dg7ztw7wBcsHBvjwAD3wYN6NmW3ZnJjsu2Qd8nj0/CLTH7rNWnXKdrgwhjCm7KQs
57kHcjZDXF3VmRl59T/M/kRPS73nh/WpMXptKjfc6jCUbzkxbeMhg+WmN15FCumiPVfM9FNfcn8m
FYUiOp2w8cJL4EVEg6tH0Q4wWKAh3BQM2/unQGJmt5AWilzkGYKt3xwgrM/HHWDwuUwkp6Keffes
U15wMlsSINy1e8T6lBDlsl3Jv/p8bTHYceHgHu+nyaEcg0YNBdU8NK/odRUnVvH0evS2w2ykkSRa
cqS5xkZsYfqVUeMpX6ig4KI4RGPQIF7IwSkrTJfO9T1cbsZ+oFuLPyaHOMschcTG0ePoY/+X52Xv
KNyOk3YjMXLJVXGik/KqD3ZFRdUu5IS/nFA3x2P/Y8p35k7UMB2102AGdRxVsYShY78qh3MzKN23
j/EQfc99u3sxjTvSr13tf0aImY4iExNVQP5Vk/Ss/Tb1/1yLqqsfw2XrPVUShG10Bgb3I7mc+hQj
yjifxm85941IuyjsfAT1e0NxLDlmBN2W3mT5Bqnx1/BmFtvs8CJqy6UG4VO9ks7vr31tqR0BW0D+
3cDZzcN4jFucyrceWVmTeOZ5UolSwYI+eGnbl7cWpNy3nGzzxdN4YAGwus5ZEwK1CtGPw4IwJd7k
2D6nE1NjSmRje2P6WKvoeohiudPcHnRoVJPwSkODY0OR/59dQzVVrmPtO62WZHKQRTq+K2AMU6Zw
zI+hYv5lPcj8jAveauxWbqjP3rw3H9kifu5mCKwrqHICYmxrBUBMmpwoTQd7SRa795cbzWWCAe4k
XtQAPoUj3MGiguioRzG4RNR/aw0WzVJyxrnMvQND1M1n3alCbHY6EZt1gtl+VtlQD3DN2xYd/I5n
MdMQfqSQZuN51yeaMy7/QUtx7y1cTzxRwvon9s5MwsF0FjBEqXfY3ruHYkY/AtG3sY3GgBLkiIu4
JzaCzhinkSgk4DQu87bjAlHETiad5XM7aYzGM+VKWzHqUlEDzy19qa5K6ha+/cQj6ZnQkYYmevCg
swk7rVBG9oePG9Watg2ccfNldr/Dsln4TOhY5JaKn4jW82iUP1bqFUIk6sND/wt+rOmtmjWtc2Zu
jifHJcLAwALI5qk6Xc5T5MqVq00R/YepQeMJPLLlEgnfp2vbq/aOyxFK00DEFN1m2GHaIQUouGM2
pZRyQPMVIbNwj0DNh95CxHf153X9lso0HtIo/dFCndzPYTXPTBZsPSvpklvXwUC70Tu7/69Zwe+p
1a9Cy1Bzr4LhyxdhIPWp59cfsi3UHCZnw7LDC8OgoCIMMFAr2cPIjExxwvi/Au85taRkr6m2lFRJ
SLHJIL+TaVdPjUyu5L3N3jgQO/iCjcll3UJfGEuImHqiBLP02N7scJoDc4VqeuioI7e/SvebhBFK
pPJJ7woKa2T9WJLQ/azCsBTB63kuDlQnBWYL8Nv0DjpW88F62BqOgm+91ZbFg+7WWpOYOsuWAWsv
LCjKxFdsNn9mwQJz7MtPRYEvOWTIPLhrejvkNb1nF5irJDWEWB2ZywWrTuFaHsGHG9quaeSD/k2n
aahlcPuj0DKGc0M9BafRKxZNcMjB/MP8kxMc0rRaN3+IDgwcoMiI/3LFJ+wVsvog20EPhp3WGmZV
dQu8325nueRs0ESh6gky1CP2BqOlQOotV6wTR+tw5c5Li8Gmx1Ds13cyJ0tLhrQvvgwspDdnu4zh
gL4HpHMQ6gJ97Rgu9jFDychMltshRREgriPr5aZSO7LR0ojApgASlL/duZkAo4sFG91Z6R00OGWL
Xy6oM2N9VA9LfBVfqyCDL/wInCpod4jQgKTQ8I6NpN4nlG+WFvoItfJ/LP9MVyvPO7h5M8uSZcJ2
cFr1ZBaGttiUEW3ltYuXKzDckLDpN3WSN/cPflj+9ekrbAfAbkz/he5I8/Hwaet6RWthRiLb+Hxt
bEGFqsG8YGj6qMsc8UDeI1OpCyvkBFWWPT1APKYwWGnQetFqbVUSc7s1fsdSMY9cfSFfSic8ngts
6kSla1nUBNTVNwlNKcSzga5ioc78bRlaVAOQxNEbduPoJYdfZAsvGJSCL9tK1dg2vvxOjJjX+Frc
ichKPPawt72KOGtR6bDY6fAjMP6FJHYq4+Gb6h+jR+2XvZBzzJb13PtgtleMG+RcBO+3Uq3uqkKr
Zaz4pkGLgWGc5UfNZtrdjLr7CsZpDNJAMv1zepOqXOKJQHcEdJXmKqmyyN2N/H0DiSX9XAH9ShK2
ytrXCKwZyaj8oetayVDkp1qFVjlQ5SFRCHy873Y/Jix7NLJtagiFv/K8aK+ZbOHApMvH57h9RVrQ
yHwdN99bBBG4Vwu6ZpLk5hlR+yPeVYwD7JiglSf4EY37aS6DEY7RGB5Qfex67TALmmB4XMHt+rVp
IEFwCg/WPaQirvRN1G5f1J7otqG0NU4OrSrnztErRL84+YCYyeJFmxE3lecjU4U/jViNJcLWHZga
PzPRF7TU0Aslm3XzRFUFrneoJm9tZU9qgFmaZ5jXMY5KJKrBD/+Az3vmM2xyzHP/J4JlxbZDHRTk
UlXKtzCxvHVWdogH3dZm8QUHCc/+9e36UE5q9jElYFxdDXH1neQQUmn9r7GXfU3tkNxYN9ceC5+K
5EJvY+0dw/2ek+dyQZ8BGj+SUph5s2lhRJ/gBDBR4Kb3goKK7UiNbRC7YsbzDD1N8+4+DPrCHpAV
IOsFe+LPJk1c4pW6zOc/5S58PHRy/W/HDRowh4k8mpqBmZwg4cHUbFOBwxdbjMf9eNQRsptgBtom
6C0JRITIOEKYr+8Zp4Lko7z1jPMODa9bXvERIfT3Y6NdxCxV3oFy1EqtDpUqlYXMYa2/E8m5evj2
30I8wuzFQWgNEXp4TNjSS6dpXu9Fc9141iYxfYqisisCD41L8mEKLLlkLWUo4k9sPEMF/AfQ+soV
N0/0h18wkZbW8UIS59kevKNUkpv47agH0cxDzPt2oF5WZjSyvy7KakKD+5vssxIRc13c6WWpUOaI
t4Rp2LQ+c2Dyp8MN/hZuFGa1dWmA31e84oDcF3AfYbG71F8OlBq8Lh4377Ako4jVTXqZa8LTM5uI
ql4ZrXn3bJlSfoARqaEuDz5efQahzMK2cww7cfAnsvCUqHbvU5w0tia6iUZXT0tVLluJtqDYK8Mb
VA/SJia70yVJ0nFZ9mTonVVLQak1uaMTcS7GUyu/FzvgscdVsUtP59YrLAN+cbnvVMp9V6wHiiEX
aokKSr3QUnQiLN2r2jhg05c0sFYTo9UgGJv58OThlrytxXXVdSnIVxuNBfzjoFUZkbSZvqlImow4
APv4msbG/PZBSaLcBzzuVxhEzOlW7RmuA6219lge5L25kZHiUTSizziR/gJ+yrkgQYSuc2PiDrwp
oBmRyNVFU0xraB9QTeyUX1VTTyoTbik6tQs4nblTBnpXNLWLr0s/hgAoN3X3YPjNUmQYLZ+y6dhW
EDq/e82zSv9gPROis3mUAH4F8N6rpZMQFt4PlqCCfwDnxEM9+7ZzZwdB68cK8HPQfEWS8uoUUIyh
Ns9Y/JAkVEnzxXSBABwvnTQhZuoQBhudiaX10dWd4cF3U1y6z8IYvc+7UnAMab5B1XK1TMSwi4R2
B34THxnE6tI28tkpvdfCBPGoivUqmxTmdO95AlxJl4Iza4tw9F9ChJ3BxJpuFVBSC/f4jk8Rpe4X
xxPDsqsaVnDHTOAVfoJxoz8YZvIhwruyFchmz3TUYEjXxw/i5zoPiTvquOz1czAJ1lbs8IjfR3wu
eJzKH+yowvHbbI4VocGQQJ+Xfc01IwEv8lCYiVldh+UQ3ZGm6DLBFJ5Y2956W1McxkpY47bvU1pA
tYHqRbZtQEhpaq6zfPklDmXBJiPBdPy5jA1aNHFH8pcs75SYPTNPbi3YpWlXCoUccfxlr95RQQ5K
5v4NQ3bHoY6YzSSyrmPHPP9Pu32R/AjAdIn6p5tbN7/l/dNl5x8B/BlEIqR3Lyh1A86b2eARJCA9
PgdXU1k97DhR97Mp5SLhIwn/B+VVqz0pDazVWNuBBRzcS3Wfdr3mhCE6591at5eUiozPBdyR1iMg
buTZ7Rih6jbUFhJ/QacsP4yITaRoa/D/JI0N5+ZPUXvQ+DPL7VNTuJZI1z6Iudwd7ojZ9bM1S2/A
M3t2T/r2dsfQHPy+rS/IAAz+F2Mq7lsIZnFS7unfVpLYFKjppFq1Qw+ZJ6DaFQIvv3StuWQmM36h
va91M65NP744D8JPAAIvAMB63eRgDtuL0XHbOHaDd80y0LdDc+3ArBninTbpiQKbp9OILZ/FiTgY
uN+1nPKUcLJITgHXQVkjx41goa8Gh/f+L9iNL00n8sz9LgEmLqGpOJbu4ezlCIly3D7P1GI1HjjA
dhnlvaOB9slUZ+TDeXMaTfuqEs3rtGhcemgQHjzF8V7ebipsm61fAw5V46y0m8oBWnIRGdpuyy+J
xSJuNLCh6I+jWgzU5U0RGMfKo+mm9cEbsTNLaK973O4VC3kLegKrpvYWvbVfzfno6phGSbOhxqxm
VEHrI81cyVCRoTJker3cz0vH7mUsbTYYYQohZJPcKp+0tcYWSiQ/iMg2noi5XDx0NGQPhgPfl7Yh
dXrqm07NOvgOFKTfGmd3ne2AEoEGoE3oRZ5M6wy91z/JUR93AI6YsiHdTsWZkciYxFBBnvMcgFi6
VY/K24tZAxq7pXveLrixKz0hpXcsy9FOTHrA7g5xQE1QZpfiV/CxBxkcBt0iS7CPWyHTsTkVYpVJ
78trQxIpFAytpTheUX9NImEB/5MdSaZm6gARFz/Cf/ThFVwbgc3StI4WxGGv42XmbBrNm4VGVW7u
MSZDcZrefB6QU9/84aqPiL5deF8ZteysCFKjYG2EGaCnBvmLSvwv9pk0hkHBGvyJCIVCC8zWmzmh
YHG+s4BR6FNk4X9CQeYYSXl5IPkDQsmRKlo+4Ttv16MRwRxjoxQ/g5I4x5demScrF6MYpQZ9SJct
SqpWO3hJHVYo04IA0OBUxKU+lui5cmxm+DOY+SDg9m5A6uvnnluQ2tn4I2Rz0Z1u2YEfKPDqhw8q
e0oOPGnbsTBIQIh1Ni7/UfJatIHfejSszAGxmpNht0i+nXX0YFAvuU826ykW7nJckGd2mNysKR+p
NGFtsshXQYBYC7CIdNMXf30W5JHHoOmM26HJu0NPgga9s5kvxI6Spp8G4h1QbbBK6UMPFtleBBwq
Xs5hGtE7Pvf1ARFz1jEi1zrXA20LC6Knbk1nFShE7mEB+YRyuYu2WbTac/vLw9/uieAdNf8Egc2b
SezVWx2zDQvDDT0mUDI6Ulycd+s0BFVaEmBh0r1vFZdNJGcID25/92v/qcKo2/ukDkprte1rqHsd
URjxYftpCrh+a+CgCtTzD2UrbPjJpgIjPGbYoTnGR9VBY3hN97hOxpcldEcIh5lewWxAPs9m63kx
WtLTHvBrwEwk6mInYDPTOlqddydeJ4RurWVAUyzhzUHtNkwt11tPtfkscGPHyLxwwhM6kWYqjfT0
jZ96TGNssaBvxgFBjG9D+7bFrhWCcrSLzeut7Yf3tOC3VjEW1kqEIPkTKwido31Fpw82xaaXxF8m
bkq0ICSsTjbAhMIMaKic4qeQcezoNRmC3xztt16tlkN4InK4wKvIIfu/OeFKpF+P96vRsyCGQIxX
WbDDIE5NRmR5sJMce+5pMtYCVCHTZmNZFI6EQ22J6oLh9togRhb6z3/DcfqiGJR5HNrBY5Y5l7ki
DHUQP87lJZw3gX2NAkapZaZtkpcTF/EMXyeFlNy/XuMLMrTbwlu93uuSetlCTIKixPNOmoiLusZF
pjXMNq/qhpYiZOKc6EcWCbjotc8GZPrwKGTXZ2o+9K3esWwbY0fwONNs+vTrxAvnPD0PkGb+EQa8
mRkkH7oRsQNidTtn2q2MqbjlYg8/c3Aw3f9jsBx+ehviFKI+D7oqaxoUNaPIafpZwmwl7VOOLIf4
Y+m2ZZq+UCQc8aE864kOVsz8tJlbIinNZQVSHvxykoqqeZFz+N22ri5b86ki63txcZvEU1Tqq8JZ
ydtu2cqehnvxs5PTN2y1Oz2Q506O1BQpCoqSYrp6Ziizava/hT511YhQaJxVZDMd5IroZ0OCW4+g
VLaCD9nZs5hjCIRglBBEKUkd80Ek/KXNczqA6SKQBKHI1M9UnLkE5fCjQZ67WHQNYm24hdVl4peJ
F0wHioZt0QVC1+28v3KtKx7IapRY13OUslt+cU4vYKohin/0twsRmjzaVFiqUG3BH8HKz/b9le7Q
7V/PKTi/RhvuHz9tSoH7G2HWxCCGIjnqT/4XABQd53BMbLapzO1Cd5hH3ZFVqdTEXaBLkultcMLq
BoMmnvWKCzJvBC3OognbqheK3rr/dloQuL1gfNDnjjhWT8UQrw53ISmMvZSHB3c4afWKU7H8Svg6
GSIflwcQcs6S6LUctUf81a7CUfqivxn28nIdahJrpbZonBf/9qTMG5W0f4K/oYaCByJJI68xCcpC
0LOeg/3/RZJqMYXUAPhltVISupEnJRnKMSnJtOm7leiwHIGYZbo3Zm3xt7Br/1q3BjHqW9A4AO+s
fVLxoiBQsCg+ogbriqb6v/hM5AYnQ1rcel+6leFxlmmvJgsXIV9cjnFpZ2RxeLcy01TCPhOoTSkt
79b9NLNW/4jefAVcT4sAUBCue2HAcY6q3rQnyHsOocRXy8FfGAQjKZ4BBz057x6fYUJ9Fv5KVWs8
a3Rc7YBj2W9+F8aewK7HHRr7PJ6SvSPuS2bmSsTqLVPl4lBJqVGLuMcFoE/YfFSAsesq77kmgaJN
l1oUR9/W5BU7V/3aS0r8Nwuhh3bTQDGQIU4O2vNAdWo2ft4GANCXR/lD5Qc+TOW7LndZyh9yIFNe
GWdETcvALCWftJelIzEiV3BVWzfi34y96QO1eKOtAZ2TSdAXAq5XQSQ1iRr4wHVgrIoYXnEeHWHv
5qjr5jwKHyG+TvbJQqusmLnRB2kuumCsgefx8bWgSJ9uszIk2XHPZZ1AJKhd9bcYFavYJSJnh/5J
0f0rnaexLS5hWoEhXUl7oi3jlgmZCQ+1e6zAlJY6RxDfUoM3veqePVYtnnEaNnIOeXz8cG3RkmFU
TJOY+GAY7BmzjwHOo6P/RGVw9pPZl7MVTA20pYm683PsvsiJhhkjNZ36kaj4COCvjjmUZ/lb/ruX
z4e1gXMgwKkBulZpRmA/g0m6CxCHQoRYajd4iMFESHcjGbUdHyt3gdP4JMZlvCbsS/JzwDLYtTCp
g9H/nPEwt1yKCeZ5aORzYzI+M+G90qjhp9DDQbpJMXSXdaGFvKm5ewbuXvBTO0JXNCJ+MVjkotvX
y7S6R6Q3m4KlImC0zZY+SFT/K4ASRsbzlNtDd9cGvEuFGiucV3B9RUe4Atwxt4z5QZN8FCgRgeQX
2kRhMRrK9JADdPIY6FFEp2SB4aul0DxaSRK8kII5iBCu3cdOrurEOHHHan3vIa1bP4Fk8kLo70Th
AGJgP5ddYkq9dHCCNubygvixStWVDtxoDu1mg9cN0Q3U1PQ6o/bz5y9v5u0cErkUGCUvra1OwvZN
P+jcAPyMHy6BHJbzaWW+mAUv5OFBMQZz8szrTtHpuRzoCaK1+6RXq6JxeeHtk+Lwif1lvm1OZkZ3
YFRysCxC+bS9Ki2CQCvYk7SkvM6pkq2PQivEN32mzVmfXzkZWLtFNu7hHGTHPr1mKGMTHBKy47SD
U5pTZQIRFdaL/eQZRTZr5eIRcNsgKVPNrY3a9DT2D44Ot5BgX8GOKok8Cn2MxvVrNvVEE7fuwnBq
3hm9yWckScxc2hkK5bkvoxGcPNLHf1JoGrOPozW7Vkp49Wozuey4lC4b7R1jixmEC0i38wjnGl0d
PhCud2gLucE7VaRlPFb3njzqfag/VwOk/Ah6vBd5kk1xHw+MRSiokB/KoEVZDf4dDNhaDU/y3OOn
OawwrO0khrpRAjn1gJZh41fHDOKAgy+kmNYUxr2tuQiOaR7i4z6MpZixqKeYBLK719ynjE3zlPLw
r2Ng7UM2BWmvqNRbOwku8Gc7dg8DD9pxfkdiHcrkLdtHOc0eJxiklgkiVQT8vYH1S6Z4KtYLM2m2
uwee7DVK2EIYjZz0K/GXPsMhJ9v/ts0Wf7/BXgfUqfsouqQ1Z4WP0Y5RqCWyhRBtvzlRYpcNobHv
V9ZFqAQx+atxy4Sp7xrgHVNrdN3PaulyfHrGHlh9qjH3yQLYlmWZPJk+V7Dg5rfmnc0zxVPOwML/
A0JkTK4e7Nc9MaLCPaM7EM+/EiktieC+qlrnf/+46nLKDYDJ8BcTCdU5Okev5rlQj/IgfyUf1rbR
2zhEBw+e5LZxOvDopnVWog/E+atFqM/FpfFpSSV5JpYCsWmJwvMdGicAWuG5l7kd80PGQ8dUlZLJ
7YS5MLR58XWMD3ZNQjSxCAAk18apvN4fyGZo/TPMz3d8asMmtjsxO+WXXiC59PM7OrzHzvnis3Up
KTrXaKEZEVX/5KIuVGj6bl8mLvaDXZ1IRDmeZv/+X7i5Uu0EgkN2QNjx3AucwNa7WhOEYKRdd1sf
InJyvgLP+2+A4LTWms7xWjKPfyWPP4/7xU2GSwwkZvzBMtYVqCwd8iHoZoLQbrPkniaVgrLk45O3
IMNUrdEMjH32espD/wIaKFsLi6vXogvz1/v2KW1ZC3SPEVXgHabjfJSnfhjswO3k+NJYDo/bdIZR
tGMEzLelbgmWD59ojrb+K3nq6nH2kB9H8bB3/nD7/+oPDFlrDp2rFke0N3nVAYouX4cmGjlUhtCv
smYrQuXb5bfVlmx76ZTuTzf7OFCNFWkWcPsYNT/gSAl/QdmU+nyo6wVrZ9plRBOqFEIWGNkadhfl
BHeUHQZLrsg6geyE+jVJnlkliKTxgJXXXU5xQzHFHoR/JkUCVkW5JD3XmvffhgFgo7gdO1CeMGno
41+81Zq4Pb8UvCyRWDOIsP9LPAXO1sDIXYPDPsrITru/MoKHYNMxKzaAVySdai4+KmCWAsY8etuC
7NRcTUuIAv57BK/Wc4u8ZyCXNMeKSp6ZA7qkPOQe5kLdXy6VhjG25YADoafTPvclDCf1+mKvFUEX
BEphsqKw+z9zNvrgflHqMAthSGmkL6RIssbW3ouYkOMnBKOhfVPQmWQMG4EewFbG30eyfLOnCJSI
QMopUolPkCnRlpTxiy1pV02HJYXY6qzBtLglkFWU0fD080bobknkIt9ptz9eehCjYWdUMiiWehwr
gYWvpUu1Bh58fQ5nPUfVQ1kSAylHQ2gwUMW3UVQtW/PIbIhvedMnIm64lMePbHg2XLn1+0Yjv8se
3W58leWOc1lGknnqBbOVT8sFn1TcSjqN0+oppTsrGhCTc8LJIu1mYDLk+3nmpt9XMC3VKbGtv9JM
UvBeP2CSeo2sPchsj6gCWSW5HjUw4neCogiyMWxar00Mv4/O83O4ORrAoYoLXfwMr6FVDji6oW30
29x3T7thVlcGs5bzGgs3wrgOtyEQJZq7xm0qd74PC6MDWUWz6Qp9wVQ9qGTJD2FFLreYiAmo36qw
hzEmr2x98FTs5RvVwTCbGpemZmvakm5DWn1hIWQApALjA2WuCT5R6Db+MWpP2ftbDXNk9kCEWhzG
SiOFKJJ5sDiQRdoxsSUHi+Zm2z5nyzSrUgU2WsoYU+rQKHOL0RaEam4ogcUCgsptwZrkdVWxGmQ7
3EDaEpnFHB+FhHUi6sctWmkkwzctIXzQfOJwEXq3NeMLurd4cGNwoSfZRA8QZhwPxmCMEHkjxnGD
4xZfMMyOvwHP6ZY+aFST9osInLKDnHEON3hMHMIg3mDVomHn9jensB5QYrXH9pBfVV8XZ8Ro7nub
R6XCq4g1UPjz/9FkMkQQppIgNUQy9/m8DbRe+6CGNBUgDBaVFB3Z9cxK+K6EJnGxbcquXBCiIS8s
nNcC8rewSCfv1R2qmdsC0vK39wMvAinzL1qR7uG1TYBeGbb+euJ1WdrBMYij0TezL/M3tCk725jU
Nft4D8QyOxFj5A6onmJ1nnVDRiG8zZfs28xGHHQJyyJOODJ3aO0eZvWB46xIbzFQwcpTV5smJqQk
Oawz7jbpBL6piS+9mmyR2Bax/UgJoLzcZZY3Ztz+1KXi0TaY9yu/Osx66LC5hyWrOb25bpM/49S/
gjr3xoYwNNcxk/lfmjHxSvYgF0LCvnRij6OlQ5CCZ60EoWE7wq9wgcWSn3J7JSyXKeNaQdYHHgPe
3X+P+iSvkhpihN3UDXQFx1SteIbk7hqSH7lHgMUxk3E9vtjQEdk65ZugGxgIJkiCFZs9XSZUWGOu
QrmrFoWWqLY8kK4e3iaxKbf6HR0Vi+GNtQOUD0QMB4oTWqNsCvpgqt3He6wAWV6aBIET1I5odmTf
/M532szx4nr8o5c7Rs+f5XmUpv6GipQN04/9Wjtsq2hzCtIAAyhkGPFEsQ2yFoEln5v+ZzxU1bCg
175aYi4xOrxednYQTzW1F7ueLigDVkdugjUsm6dYT8BtLFKeO6AkJa1JhAve8VcKDLYKOfvAwe77
+sQzpK6thUADC3Cm46MvqhPKfceCfDEqVvPXPnhRY0TKiw4vtD7r09XsCad0yblwYju+qEtn5TCd
x6owOsC4q9r3HzrKMlSlFWTVCiPwkNfDLodgH4gETxpYzrirfnp+BQjnK4WMUewaDDUeLAK/NiM+
OPAKjvKwcH8J40ePbhVfY1Cg3YN8Vv1x6Ob60eaRnc4TG8Ec6AzvmH7phCNKsqk70pB1TNBBjWcF
Yp4OUvqsgwzZdAzur5VD6ULKhXo4kXbbzhch9v5SM3WUljN8V7DTq6O/hduzucnluNWpCB5rjYbl
/XJGBWPNrGrkaBwKdjxp9gyq4wuh8CqWiB5zXsSByzVBbm4zQzNsljXNe3lTXbGwGufAvsQEIZB/
UNmj8Vp54Fue8a5bhvTBc5a6dEkr0kP9qdFGtRtXt5MWcDMz6kAT+VVibCZ7LOTVJcNTXcYZShe6
p1iCp4513sN6F5o30X77rd+NTzUYk0d42FRpzxi/GY/in33+srx2K7yvPHp+bOcf5Z71SIjjPaLt
48Vxvh1s0K1/6+SRdfqs1liipQFXfJZ9vVmBoj9W/S9aBqRRknEs1YY9hWCtJUrB4krU7RLLWqWW
uPhFpeDsKeSI6tCRPNPRzMGi2g2XLcY+SnCMZoM6kodjv0DikiMJ5qgn+89rBz++kEc5J4YG03VE
U88EHV4Vll3Lk1RQzTEq8Nqz50rHUXbEqeAtalSWa/guXpopY1tRsnfqjl12/r5tBSzWthMRm/0a
6ozkvhDif0CCjk1koh4kTWYxCYrXzKb9fD6QGdCUgzGDDztMGiA4mzCNQqGSSjl88A4wfG6y3/jE
y+c1Ae8q1lYfd5okAPYa5DRsovK1aEQCQoKahv11BIM82kW4EaAWeudJxqnkWMS2jI4DRhiAvtF/
sESkY0aGX39DpdqT4hUcFF/es36RxRsbvScF8ypw28PhULoMgk91V9RWZIgMjL7AwgXgFAmECV+R
UOcAPSQkty6DY5gUTeoCsY8kYjFHC8tjNNEUV3eiJkEPV52Zc/Zdxvc4wOCrY8MzUIDNVbq60ywB
afLakPicsyanf0fy7S+aY8gQIXDWt1fUo9IDcy3vJTp2d+NgDnHQp9m/8BkbXlhmp7eEPqKsGqRe
0V/UVDiM05o/52WPpWa9WO4mn84Gec1ysWO4687S0A/Z6zbQZYUDmw6zZTVBHbHE8rzMzs5rz1aH
UkNcGq7ys8GThgoAZTQYKvWaL2eA3nL0PJJT30fNrkEcZBEEg9OyHieW4eaDasw/0Qlx/hEWR0Ai
oHmuOj1+UNoGsy9POQ9uYH4s7iO5/QpC8ejYWYud9ulcpty7Nc1clZPPpck60Q8zopgbrdd9aNjA
rBMeC0qDoHhqHbYFzE52/yvxb70XkWJI5j9n3P/1X4Q1ObqpHTfCQEJkRlEcvpRGiBzgjoTv6/Xm
kxcKKzowdpiSqqH2NGBtZ1XfED53arITDQShxF1uEmhYHr1+ciDViZuo5SiT1e07L+JIe9dkYNcV
Z3J9vWYppSD4SPjA+gLVSLsRCyJFiSv5hD8A5RAIUpq7D/VPiFxNzlFThxy49XnXndSK+TmgeqjH
ii8WaWWEw0EFmJdKa8ypVkuyKeA2FY/mW0A2/aFMOqaVg3iRJgvxqk+2RoaYwrJYYHoFd4VnZGB3
dDbUuTweaQZUObvVxQQGpK5PQ1Pf8W3HQo+Cu6FC1Pue2ObFZZwDNYiiH1yjYQLkLoFMyte1+buK
TFUPdC1tQq2675fcQQJnbbwBkuKlvPDEdAkH2rIEPdd7scpvDLVGwsHYGfxQ54L7hPtUBqN8KOv9
wXmbvme14YdAV+IPtMpKF4DlxwsEQvn/dhsnGYbb11KU1fHKzVwb7fMRlS+7ophALOtKGFltdPU8
ZPRmI4tApJ9xOA/v55tjg8dUCEYlrYOti5vz8V1ph6fHeqY27ZKgpvRcKK2w5zOTVbZFytD2tWq7
8p4raxStr76NndESX7Azrz2n6lf/w/+b1y2GWrVbHWads20qXKkrxbEiWSmFBbJ8AqY7tKNiiAG5
dy1+Nfb2UWglFuCpVTpYyBBZ46i9nV5LNcbXS+n/+1PLNKRCKUlMGVJHgeRq7niswgIwL22xyOA3
cDll28G25pT7jESWvi0SnFe3Vc/CGRTjhLrUGdOOS9g1PkJXARf768fKxfmtj4HE80NiC/woDHA/
Zwa7bTX5HWxMp3LF8KkxIBgs7/xJFbpgR7dwB+1e4TNNoysY/tQrMMlt4U34pzeLD5xJqZisrvTJ
L3Pt7EDTfRqifIKnoodPcjWHFidyLFEXg/fbWWRiSU5LI2z1kiWWTe5L1RnrEwtVeswF+8VAswO/
b+ckh+F3HNHJajIsiU2zaRy4LEebFKcvDukXxUuix+wpfnucEv1+wd8oB3Jq8D3qpyRqTmsycIPs
7vpqrtBr0AmCJBbQdOlCXBbqpTbzIvFHuHDznvLw0LpKCA3GNM2q8gHsLm/L/eRnwvmDPmrMR+ai
sM7v2Kucnjp9JJz0U094xdnrPcC32w5nzrnF9SiXx8kJhzb+i/4x78dFgjPfAPmkvwPpPaMtbpNV
U5yuYlUfKXUk/4h5Uwpubqm4K/eef57eiNGEXgLr64rNo2AYwENmIn3lyo8e00heO8mhXMmiuRZs
sBzqZEUbGr1nHyiBavoeLpUhZW6/lS411tdrmTivcC2ITLYjlhxpycrX81+tzXN44GTNekIRGPix
hvPAmcCgsudYoquJRpHRsSWLO7mgXeg2GasNQ7JhranwtZsiy2jcBnBGvtTr4VzICzZpIIRln6wC
t9WkNeLNhsnMGHl8v9EaiYpCTN1gmhAYA4eb/kyhICDSfz7FlJAKEC/S7MZxecI3cGxLB2sRj0MZ
NmMJGmj6Deq88hWMkbXKymOlnp4A2MIkJc7qgjb0bznSxocSjfL+tHMYF4CAlIhQNXWFhF2m4pmJ
OKtkEjaGNMDAWWpu9Y0ReQSJV6S9FB2SB8lcV750sjzmrU49bKL2Dr4o4sj54fIzSQAZ9K9x68Aa
6Nawab9XdyMOxIwZV1XM//h9GrV19XG7o/ALjzv3udkDsuf/lKmvqa/m0KBpTffS3vnx3Qdj6PGz
FnpyMjN5t2yHLfDI3V9E27rZAY9QtFIFVRU7/FoInouBK56au/krcNhW8uFNEdzO0RiIdKqcBB05
6erW8ocPRZElIa/QIu9iXUGSiIassaIFy5SDGSCm/GQj+QZvWdLKFWb4PH1zGI+PCexYX/YNTG02
alBVhrCTgwoC0lwCjaJ1wnye5qpq9yyG2Jet09KszsuJ5z+PwB0EKDDif9T5PSEwKwBh6pR7BwDv
hQZZ42eAI+zzoVT8Sli31298rDcER9l6fWhAmtnVFYugvY6BkmK7gkdbNJThut7Pp8pUZt5aXmPv
9wldp3BUFXJDvGNdvVlTHxGhhfLjPZl3RdgvrPQYgnFbUbOuDhoIQdjmnYynL1O+bShhNFuanunR
oBcEfStnP7OT5UEI+pzl9SZ5Jx4JJ/O5eIEGfPmi81UCe2g9BIfqki1ZPsTUtxyYwD4AaG4BWuWz
5nJ/EMFTi2rWg3hK370wQ9I6dTQLXiNP6ik1oH5+Sg1gy6/wiklnFfTEeOkK2d0ukUWSzYTvHYbO
eK7VGEWgLzIpcpTZslqKTorKl7bYnfEupu/OGIkYuHSbnYnFSch/tNoY1pTvbPkkMmA69T/MP8Pn
Bm9DPkoo1y/5iJ/uZJJDltAGbAErcuMntSrFUYb92UDc4xUYyhUvg1f4dLMHysxbZicssCN9GDVe
5V4dRWCCazKcrsI1PT06T59VIa5PRD0zokJ7jc31Bj4QC6vr8b3SjKYe/f0kdFQq9k0YtKFrwT1W
4/GuGojA25aJUhgqH3f1Q/bBscPa2UICDRxwpsjRKGsOFlo4ogNKo/wMd3cgm5ABmvdWoC9xD4zG
n7fYLDJX8d1UUo/Psy6OV47A4k59vsOLI62l8kh4m5K2HECR1ncvziyjaLJRsi13mJSHL09sq1M2
BrOlqVoPBu12rBqL0FMDHcok21X5iZwiElAhfZR6OGSTtLZ/r8v3vI+A85xNDaUYgwKTqHj349ci
Q6RwtMdKTaa2TDJlLnH0+XSeHznA0QSJKXADw1nMqlXgwAXibKQHQRVA3c1iPXbfVONMJ+CYNjbB
ixDLIui3HRhjRt7QV83RlSaOPdcU3ydXQ/pYwt7SLzlzoRt8Pnj528akPoKFRMPWjVYwKofS0wA7
wI5/jlR11a0MwdtU0SlX+4BZYeoYoQlC4NvZnEaKDm2eRhG2BdB0TLdDZ7esUNJZXIHMBXDGo+cl
ULEUQvocVTnIU1jrt/CsB7fWU80lPL93WrK7ola8eGbcHdqsBXOsmgIWKt6mJ1Xj/m9vQo1mIy3b
RK/TYzXypiMkn2+fVYKHQvwdt5IMI5eC+s1yHL8loT/wSe71fkPsUoZSKR/qe2fQVwqpwUFvWqyT
v6/hjes7g2ulF+sLP1UVXLziw1AuOSrRnX12KvrBc6EXQW3GYt8gvMb/6i114bh95l8Dk+//dJdW
Bpt8pYFUX3PekPy+VKPsFlsbrKDGD+y6cO0aRe5KnD+QFY2LQnj3J0zwPzlUdMjM8mCq6iiqkG54
S8lvOvDnoFcb3rMFhQxL8fDw+4dPOY/H4yf//tFkRmDWYMs3d0GQJvf5Saru1Ldx4VPIXjWt+lfj
qDPkxLCEbrbGfRpuQ3g6iEwRa/zFHSBItKoWaUwt4j3S7urm7ljb5YoP9NTR99yiN3+qeX2nCR46
PhPOUR+gpmA+5rBZusocf658QMiXvx5INq2IJrappCW3PWyS9479MSlYX70XHH/4HZAWPWPe4WAS
EkdDyzUWzOnfR6zC1CqKQhhJ0KU2dq2CUTldWoxqp+gNkf0t1gaOpAyaN5rTKcZg7BFZphVjNjOA
oxv2NJLTUjMyrmJYV+Gq1FNQrsYRgfMIZH3fZASXmGS+CmSSC4UtoVAxMvb2GmPFuAgyhhw+1ujt
rQjqhYeTuVygav92MjmqsEd7+4QeRPZXxw0yMfamqgW/8h34/88LOVtGILgKNHOgAKboyli/IQGz
Ig8JR4WZrs5RYxZpk+7/dakIYJmfdjzhPaVe/reWvYQVm6x8pm/JfKqGFOZ5Dj9ZiMtA4bJMqms0
kGwQ776efSG34evzbiJKtAwdbAf4m5glXpC+WNuAF01qgYzZrNWmgoRTG0c02xPI8m+g/cXqRpaE
8fNodyBHX0XHv6/1aAlvyPX9zkhna8Tln0hY5Y4U3bznmfMssZgPRxmwhk6mZJ5IaavHjKYit3LY
MRlwIQdgVpCVFWrCj/7aLrvrb6c4KnqEhV+TNwhx/G/YaODES4fCZzi90atg4zIXHwBcUGgqcEQS
dYQRan7O3n9MjJZH+XCcRzFq0BdGoCuH0wg8CHxnbS0bw0Kh1C6R9JNMa8Q8hepadTKgGVqR7NcY
1TSzaXWYpxZCcb7qale728P5mHtKeO0AV6wtlBe+vj5AOxmUwG5sGPaX2rdBFP/FadHNTqbvClvv
UNJOWo3H42FDSTqzt9YyujXAlfC/wDzFWWwLrazpmAerYGe/QziSshMAVOz73xwpqJ+MqbGWYeil
ciHlgvbcj4xlPti12UGQ/G018paEMqAZ5qcjZKTD2bfbN51Mz88JkrcGwSyIYRm2I5Qq+TZFRRxv
emgBG2ttHfYU9Ah00cAC+6et10ToYyuzJAasqf1x/Lb51e144H6OHX3sjJfDY7akEyHl4Z4ZlqY+
n3Q2+5UnTYFRdAMEemnHx2Llzbn7ZAkt8u36F3b6eKqMxXh8ub5/1ToAGR9acUbVKZpfIYcaYiHU
uU2ffteALiE1Yd7RyszzDOUE8oNOj721geluxj6WfZZpPFgQmrYJxZSsPtTPwpaBh9dd5WTTNp3h
DOhyrDDTLN6FVG8yhmApC2b6+GxedLmOXunVuJHbxNrBxqjgT/9ayVgDhU4c0SfA2qIzN+8qQxGN
u8EpIB8rTDIWihBouSOoc7eLXY3eVPI49RITCoWG8RV/S72fwuNZCxBI6Muv80bRxcRnsFWHmG/q
oC8MHxGE9hmjTpmbEIW2GFK3e/Z+59V94wOYqn+pUMX/6Cyc1gDP8l4HjjowUrOq27PTIDtruW0t
iaY+maH/mcfKI7fsZlx3DUJD7NfdksIm0ScTU8lgX0SVawFG0eiB2B5ImHacNrdABKSyrubY+OGm
IA3rCdGXjh+fVdDYWMvne5D3HYlJEpl8hojT+gSDw+9iVCzfNqT2PtL/C/KJ1b6kORBhZGcCb0oV
uZC/VXHrmSdaaFBOQUzo9iYxYCZgPeQ7P7wwEi0xb6+cVazONuts4yB2gfOwCffro1YxkDRLj+D6
+3AkE9xG+F/kMIoYByduCPz0c0fwfHLYIRLApy64jaSEUre9oQfqe55Om47aw8t4LFb9S1Y5fetv
dkD/Nf7Yvv89yVVl2px8GWNpGKduM5AcwWQRPFE/hd+oKyIUNMOeMgod6OJf1Og74/PcvsWZ99fo
FAbddVb73UY0OkaIMzVe468VTPMfYSZ8Pyov4y3moLLa6pGWo7K6/QUT8EEn+RpU4iOODg1iy4lP
tzcpWmh2iRQTTu7YP5hBMo5eJ0T0cLNvn5XUtysAWaCEKr1X5fdJdWMc/DrFmMhQZlRmjRRgYAXP
JxZYmiZADI3c6KF0HnwzLBv4yfd6Uiztak/WAmw7mQYo+iF1W7I0fN8KGyW+fP0BiAIWpB90Wd4t
USSuWyR5RxvgT9WqVtL4gCE39rBSiV8WAZefnXBMrCkmEfM9PrpBhVtVYixXGXTo4x+Hr4uHXtq6
NjSTUz1hJEV0TZj6GCK57HVX4ZYPhUGtG8dSi9D/5lCxoUTibfd1UM+RpuKkx7tHD8MbvP1rhgfX
4oiILeJPUSV9h1T9mJivblEoL+ZzV6P4NmMKS7ZvszMrCUSJgKx40j6xtpBUfQRoc/nYpc5OQQ81
wyzXcFApiiUBUZ9kMaAhhBsg8aHzQKRpwJx+yBgR73RKPZ7YT9iJOBRVIEkpF/nnSDgb+9OcFdgf
tJ/2ndmpxS1UVv3OtM2pX0HGT+wC4deFio0SOKSIdFtVqOqencII7TLtGra8J8MxFZ9AMIedxmq1
E4VaVjmptRJ+7aTMrQ7eayuqEbUmvWiCVKGRFACFD/HJl70L1WutgbQ7fgIlGVIXOdOSntnBQrgc
P7pm7ahlh84Ly2IX5n+A6QwlYFSSHxLgXgiJ3w/ntEpwTBarAWuK5XdTqYNspV9gH++RRbXrMsG1
VD5bMFNXTE8erzKPng+XqbzgMH+1pqCwOsDDd6uXSEl9vlaASQ/v1gGvnYy0+sSpatFSzKDD9Man
3wi2lxlNFXvoooGHjhtJJToN0kbDXAjaGH1uXqk2tR7AVrJ5x6R5suA3lKfkWjaUCD5XFVYwCSRr
BZlMfHuPvBLv3At2LDDEB8ZRdMCMoX7KPG41VkzJmlq54mJsDqjfWPca07HvF9GLzdjTFys+aWcW
89+bGQ8iNKbvJkH3rrHrxEA/pARYCxdqdutRkG+lwraI/jjT/e7dWdu6uXRcDFt6qZhazeMvYTiT
0aHxBjA4AQh9JGIbMrH2Moj/jg5bHUFJ9pkiS/CywHHXqiSabBLTiMNba5sG3Y5DLe6G1UxaoaXp
jn+24EIUKT5INYrayAr92JmhUDmZWN25Z5i2AgTe63dmvMeZvmNi9mqbJQ0kHxaaR3ecYrtIniZb
9Gr9WX3HfJRyaYsZ+PW3Hn3mFlRBMt9QpLvkDCwArmgUC00h00fpEcLr+Dz526zVUtAAXyPygBq7
u0oQKGi+DnK+sfKqQqHAdHDKo19L7WEepRoBp0kOVVO/kFfrkJUGWm5L6XjVSAhuRyGjEYQYJQri
67H8l/Sy4gaYb+Hy24H8SZyezQJ6xO3aDg8jubqI5pWupYH5FB9OykIOvnl3KQZal3MhWEOCB5p7
Kmt37Fd17M2KPf6767ClSk1fG7xYFyDuIOkbTwUGU/wsWYbBo2PM9ENwN2bnJJ91/oqi0oSuyjZN
9xRD8q+l7BchT2uSRM1WOYJnFDfU0DRwwVgQU0ap8RTU1tjEqpOekp9nGQ8NCgevZksSiCSXa7R3
g1PJu+RVgEweFq4klESj6QeQryH3y9FTMfXDet3k1Pju4j3NLCaF+cYc8PBGTZgak1iyBevoYG8l
/OcpT46+r0yKGIliqO92t8HLBWrrEOhQAnyg1OGu9veIF0Z5WvdOEvkHhYskjn68Mr5WgJSZbEQa
irX7htCr6OE4dp62SP8Uc7lKIG27w5aRQyOSLUJbOvba97z2bXFTRRm7c+Ej1Hh0i1ehJmx8atFK
Dvqxw3nFGQ3JSn38FOYxEcuBLdGRrVMDHWr1ziiYEx/jUbSI8KWXSDTAuJG7x8mZEKuO0QSoT2dc
pBnZu0Eq1iYq/E9nJ4LGq0ihYb4zrIvdR4XWpYWIZ3LvzmPkTKFOfhDUgyFd7E+7YilXAYYMBngY
Y4uyRuc6aNJwMFQU58ipJmJM3ZkV5Fb76VWZmGJI9F3aIZBRgcKFaDwJM2QoguFW6RGPq0jdLtya
rEcwHiwLZVaggaJynqsFjclaA3nObWw1EE8U+fbSCko4hulDUHZ2FFyChpHxZsHKAVvsHwyNgTtN
5GZH2zzxn5Kq/HzOgbnm61BwUOBBwIcd2dbW87MKDtkXglkah1HDj7xt5HTpe53eQPQ2IXA4PU3O
n1kLXpkQbl3NiPnpbF0fXNPjzf5I3dGzoVz1iJw8TuFl3UvpPVoPywMwtbzEIwWRMBIvdWSp62JW
nhlCJUuDsRZJAqAmhRVoSOVh6IF3LBds6HKFgFMKQ3/zQIEHp/syjYztD18n5j/QeRFHfVrbbP/p
jtKNQSBohIpOQPL//2ih/DFLsg/lfqZh4+rrZcta+EvqxXJwQ474Ukd+kTmBUkEe/DVJND/OkanY
qdgJHIJJ7s6O1mOGcnTTk641+FWAnIDMug0v3l0Ew3sVaRfgDMfLSf2aEEoEdJ4S7p+FkGa60b4p
OOYyEBk00TelFDkmSpCk0q8kUzq+W6dHSaIsHpIY78IBR86leZKrIZT2fgu7FoWToAaZ0RXvZts2
ekDM2SHONsvNhxJvTGLGEHP9X47qDPmnvOl5QoNRRkPx+vdmVwUnXFBdL0+9LpjG+3rV/05Nzrpi
NEuivlBSD/nrR5qulLcPutmMaJAd1sA/wYSO3FmiMFkPV9cuWhQsAWLQR/kNQvinxABaJlXVvzOW
FzF/MVM76RCRN3RjlXY7gjBzclUccoMJ38sx3S8VOOI0z5Xl5koM4Gj9PHpU9dopCfPtb8e3ek/J
UeUN8gdefZu98PT0Vm5vPo3BE0FgqyOZ/eN0kbW9mkEatprxWJDQg4RuK6zp5jCo0PurO+MgZQM2
8AB4bTxinv93dX14VyYbqEtCkA3ZhWxcLNBiIRyg5AeW179NtHu9bFKbLrchjOoG6PG1JWMFvYey
iwNCwhB4a9A7PS1eHGIX6xZSkuJ1QWwUud6WN/lWVrPe2NG3PimhPgVRN5gA8J1pS2VvNqP810l5
2cQB5u60TVhvsXoPVT5JHk8W6B7lPu1cPcT9pTdXaJj//qdFGlhgil16stphpdk4+TCK9ZXMen39
hBCa3sjEf0wDc2jb04Q2n1hjErJmGV766zHE48IXTWX+EZWd/oRLRscnL87qkzKfn464ocUrwyzf
x8vn8TCOj4fJfwtPaK0lKPrn3GJSPymtIxdCo+XHfPH+Wjjcwu0dzn7CclVYuSkShx2tCYplx/ZZ
e7oDRCEw0QFihtoYUOiomDjCq7srNipZIicJLktGR4mJVWwkL2lFHweFjyhZ2FmHMUEngfviWFDQ
wPhBgyCZDlrSd8KbqROvf9QUUbg55FZPndVWBm3uTwJ1rjdwn3fj4ilieXi7nprFprw+H4wpjfmk
MjHECn1nH4mUWQvsPYnpgLaUmEdtN+MFlzJXCViOr4TnKsDlfVoTXjkyBTFH0+I1tEDQQmazG4oA
4MAVf+QGmO5Ec29JjArB2jg3SxBAIiVim4QxyrASOnOMl2gFW8QRx9s7oBF+48shEg4oeV/NtrxS
wRrsB0RyLwKOD4k5V094A3f5tgVXyeDoGzJizIsqXy2w2h08wvxVQ/T3MfYWvYk+7w/N5i0S8p5K
jr4l9/uSg9GYjrhXY1OJDVVSJiLD2pcGv4KdjV3guQrI7QZ9ljpTSjmnial2FAP+RD3M4R3n976s
qRlv9oZ9l5FU0rcTfHXDlUi1Tf1OR1Us89HEZO5kbAD21SNilfs3XK/5lu7ZfHra257t74Kdtxrz
sC9hTQAgqMZF74hHIzTphpPZpeagu7l2F16VK1m3/tf7soZbwt4o8bqDFG6TIaGmHskXXsG6PzyR
lKt0D5Qu4BpkKSP1VGoUVPjb35iZtrbx24h2kFtf9xOzODzqmKuuZVhAd4LkZTpzDICKmGd1rOqr
gUpcUPTPk/Z4epRbty6fKEVB+DAWwNHkW/adWoBaIDQfHBOiNoQNM4pUMqdYM+I51YJap7/zVCwK
o794xm+y/0+55TUM9PRX3HuzkAiY+o8iQ0f4vf+jSZWwCBt2vxlI3N4KwTD4Ijbn5Volb6mbsSd2
8XgIZuujRjT4WcBRxtilXsITu5ttESkA6rGYBHU1Fu5zv4b4+3jZGgSZSR1d+2fLXpB9sz2ruNmb
yQsMrMZGSqb7XO92FtIRWD67PMUvKopaXcCat4CQ1QUDmh3Rygw/Wn92rnjTr7T12VDfjbafXcug
YI1l3t8ufWtJXJo4kWKPgGMh24ariKxW17Rybi8VGmVlECQEWl54h+de1kYP83TTZn8pZlephDA9
C596um5oGOg5vDg2q750jQ2TuVe3K50I19PGi3w/g+YR6moysjkAtl647+P63fewDJlPO7tALgnd
gAgK1uRsxkOI35uDxtQ8xtQtfw5iA0tXn8FT8aa1R+567WNwUVNFHsZBa1BDHwFx41PYbjpoIHPt
hWjmNhTz6tj7mGZ8O47j5rh2JXZZiRnFjUNF9GKrk7OqcxUEyD6Z3V2Hrs3pLV8RGgdO3oABep2/
Tt43gzuLfM4FzvIAMv3o1Vio0O5H60Xww0feYCwikCNKcA35Maaw/77FeCootTtz2mkFBOeOnrx/
Tilj+jTAXV7E17jQUn9HaXzLVydPDmSxSOf7nVTajgVqcNvtxPUrI1jkI5HYvbT9JRDycWpqtpYs
E2PpXM/IgaYSfjaJQpx+yHLJKNDvbat2Y4O8sa+a18RhtEsSQ+9UF3hGPoy4RonDyd/qDVYX+Ft2
cNF6CjriaNPoTCGwiE9hn0ysv4RvCv+XoUc9e+tfsdz8ORBc/F6qX0ShMXVe7sHXPu+C5HIDlYV9
7jxGJvsCOYcKIxG/s/YUsL4paSNZGAE54UIc3jMlqvwQQckl2PA+K9d3krmPO3l3+VU+cZF8UNUz
+ObyP43s+bDSxDUbYFwYQMZAzXkYYVPogSzBxC3LW4COQSHvF7AI/UMK6fe4uJ3dC/GassTRHZV4
7126+Pq30zPSOTZy4LAEMOMQ7mD+rdeIRSHPCEKKywFPjiT94hAz8kQBBj2WSBrkqQYzVxpWo+sP
K2t9pcU4ZCuuUi3W2GggywqLHixiRMqGR9cN8xURlWTMUQNbE/Zz31XSQyDTydMctZ3b6ZSsQeOK
ozrlz6rQ908iUPpPHIjQUtVrktydeJh95mJp6rLR7itS8rYJZv0+tkN/rJDvV+5ZUsBeQ/SCsV1t
cKyXw7cKY+gn3PoFolaTLGPu55VVDZh4AbSPovStTJgLMSszI46FT0sma2DCH9pSQT30eXEAaqNs
jLzqGF8Alc0dkgk50IPFHCgU5d976/NJpweMyLtRZ1Y2pz6jUNnnIrj95yNMQhzlnSclLdrXvgSJ
0DLVBQeEG00l7VkBc4CdnXxla5wWwfdz6neDmeY+IvIertTaTX4tWbHQM0SwH+fsj9Zx3xvmm0pL
jDRpHvGwFhC9gvky9wWLr1OmzFNr6vuh/TyS/b8m10Z8Kly9TQDIzwpJ9desQWdDXT/EhnmotYHC
FnL55IdqE+j2tY/hGtUvLdX/5qb1mXGEpAMH0hadatdZWoNQwTGgSXOEo0b0P4JvXlgY6FGP4AzL
qI/kcl3KsuVNGnTGNKfuLkVHfWfS4JTa+SzCZdymrQa+RrGLhaDpnKB0jGxGjntAB7goLwSM6rDJ
o1VZFY9Epf2U/LN/AZ8iW377e+dmboqFKN5yToPqC+JvBEjX6/dkYVdLjx8I/1hgmZdx6BsBnJqO
xe0fRKlRemXBCWLnIMBSmDXBTxKtgbVI59jBJTA6oLJHh5RuVD17sMhaev6s6QaohRoszyTwcIg6
bqKaUoQjeDgMzloGtd4FCqB1B4qxaSgTlfwtqb2SQze72+lo2nqDnD1aiEgAddSbRSr/BBjElRz4
L2VH/BblK/Wr0yZjUIJ3EaEp/Pc/DBM0NwbjmMErgrrrmpHcRAtu7C4Ew5v2LPcIEZ7YBEhV1YZy
9gCEFj8J1cHFQF2FD56gGI+iZ5j380/Xze968Ku7EYZEbUmbSnmtPDwu0YZo6ogHYlQVdn9fyRUN
s+0PKHKe03E05bxua3UCWLmXobF5ivasxshvKjHbYA1DsVyNptyFvhtJQ5Zcfly0snABuQ3Bvp6N
NpNWE3DCMKKMk0Fyor3yYuHQ/mTreXutKW8f8lMKf3PZ+n8JIcN9ExY/4f/YJzvkLy5Mkmko+gix
w4dzG8CPSNEd3nzl6TZwk2RKnVg53YRnhl70oNFzdGySQGiVAry71ieS25Vq1SVgUqivHc9fkcP5
VHOk8/PFFIvSTUk7w1Dw8vj6XHoHLD1d2SXxs4MXIuVKhnjqMEa3hAl7rS7uq4RfYRbMSf8LNs/f
bnu3YCuqO7cSxRyTP/lNZSZErBQf0/GZQRri/maQ8GSinY482eSg9rm7CubAsLggN0RsGBH2YbEa
em4/t4HWVwiClM9n+f8/7fohFvKwHGWDiWhRLrgPT1bwvCjeIFXaheZK2UvrPu44JVOMzYkSkIE5
TYGpk4mDEIybbzu49KCnmo8Xy7CAT9CSsz3PnwgnYtyZQ0BOtMzZ21FwB9LYtzJ6h2QmQ7ad39bO
jIPPpL0pkTyRLtqmCzKFrbLJxvHYw4L5mR9lr5AjDARsgK4yVRwQEw+1YgcTfC30lEfZS9WDbTck
yQ9RjLywsrko1LvUYxcToiHoCuaV9/t0Rxjmlej4PWPGqP2A7EDWp+7gTjP6TJfFnXly3rKKQo+W
j6gjvZElS7SzXJNQF/F/hIv6Oxuepe+upkh/o0WagZ7u9fhybRPI1Jk0yALjQEJ/SnZmW+yD9405
N3Shav8DLXuoPDhL108VhOhZK/iLPW+HhT0qUP8QH0b6v3dfZenCCHGfOM1ORNzk0/zipbUuqUdc
gSE9Hu63hO0JGCvHNQvJOTzVEgUfDWigRgs9w73+DV0NsJOcXK5bw7+Je/QZ/IRu3ICTtGRkaIYn
amN/xK9/8VCuH3K6WmdOUZEqM9y4q+Mfs7aYfRNZmspITOkO0y0wmABBiLhxBlXHi6rySNK3gIIE
trCM9E3shSUxba3rak3R158tEF5puluswNmlHcfXpr1Xsg81HIlayA/Rs1x9C7B9aO6utSagza/X
qPDGIC7oFRRQ0pdgSD0caBOJ2doNh/6S+30M1idQnG6ZeRnW7Krmbc5byOskHYa9ZIiUd8agsrt2
bwRWpt9Yiebex5YiRTsJJTGLY4uEVCNgCCKzEUp3lQy2p1e8N5BXUu2LGrF2LyfL7mulRygsWZUm
C3URZhC8S9zVTBatoB6zrvefiUbKTG78Yg4iLXAlphVDw61WHAb+jxtvT1Di6KEa1YKY9+jnEOLa
c9cgPkF9R3s2X/ErHQPPLJl6nNEaWVL5ejDtWab4toLO4C5llFnJwNBIobnANQ8C/sFQ26cOVEgl
4EnbJIL7iMfMsirtrLEw3BXVQaWwvUQwefduPQwH3vuTD6oAiWedcXBoPjTB21srjFpq+OZO/nue
T2zzjKoOlbAs2oX7PHCSo0qn7Q2hUGzyL9qSlzHySag3TCvG+Wd0TuPo9Fm87s3hHWzRmDVFJUI4
Hv0Z6Xmru6nJd5bACosl3pjH1WodwUwU3cUDmIy9P0muYsvDxdBOAzfGEkJBnWABfQCLIErXAOlc
fafph7B41Ve1U7coFHM3j/NZMN8O00WJJk5olKoYGeR6IgcQsuPaQ+W8yWMhoVhyhYYglOUVSlO+
60jhtTv+Cnct5Xw4bquxcHyB0oGXnl5UXopt67R9YVCNK4PNd+Anaitrsu2mXJyROb7QT6cooZjb
GvvHXqW0fcei2srvLEok3F5372SzjnxTbqs8mrPHRIDETc9fsiR1n1NNBUil3QcblB5t+bmkqv0E
3BQCl8Tem6qydLA5pjEzLmpxQCrSBoYF/RmR5xt0aT0EKJuq109J0p4enQ7SUX48mWE+MEUl710m
k/vHu4XOCr1TRdpYOLZtXb4VHiHbudtV50yeFtk0LeBMwhaRZ6gEipb6P2ojBv/CllNtnBtSJoFM
mOIvz9mqiWMQrGKKpdydp25fRCt/Oo5RaBrp/Z+3uKPFNp8CZC4zrHZ9txgXB+YjG+JcfiByYzDH
WATDfag3G6h1QEuUT9joBGt7mMQ5Sz6VolMcRUdc2B9gE5a4jRxMiv4lMMwfqssks15bxUswNRI3
TgkFTxLn1TDYPT1FDMaw0597U2XyMbedIJQHSeoaCtZg9CO1k2VvwaFJWoUWb4GCUPk+UsTTEsDC
MQ7/N35Xk0BL+A5hPUZOhcMIZtSAUvDzAo6t90jtmw5WWbZuXUZiZGgTGs5Hfs9zJlHn0Q7NIvOL
II+LaW69Jkm2O5V93uab6KGaEvo7d4IrnabPjBGYT6u1pSwz2tvhHx9jvdJ09eF+kwEC2CcLCT9d
VzpHp6A33PL5KSd91GqKvDsyp0AUwZZw6NA5hXDu0DTkPFT6/PMY0E56+ZrmD8DWnuBw7lRdIZyF
lFJSZlAFfoC4wrZfDWyQQ1lC6exRDgVSunvSJbroxRkRlAD63PNGvj724ww1QvyBOIFAPvUJVC8Q
zAq+1RGdtA3pN+Lt2bOYKmrltGZtFDMZOfYZLWP9V/BC7KDrEyD4MTUe9u9Wym91f4PJNLk0boWc
aKhfQFA0e5WSiXKIIVzPcsnEtWw8eb5tKb3X8NfVReB4ipM6OH2yfL6kqGdS2xjT4F6/QTrS9vCL
F0/eG91vcwfb/Khfupcu1DyTRVmXbbu2IMqwBHfZaJZm+yfu1pRHSeCVqGkM5qJzxiIwUFTSYF7t
+t7B6hrYqDhpjER7S6hE39Fbgz43B7zBhuzS1DmmKOo/zJ4ELI9A7+1QnZga1wbPvdPYB/39qYae
mcEexgzrZLdaveMBMf8J2tZmgRJqqMLbYdYshXhQZikWP2l0miRH5EM7nuMisD+mbydXOb0tTp3G
koEmkLM7SB1zFUnEn0bdllA4ZhDDuliIwGqV74W85lZrN3aEGpO499LzUAHi8O9lKBKwH+saMWym
ON4D/oRpRoznbu7NfUuCCSt3xKLOLFJe6yLtHhkVb0i9UGHtInyWNtr/Sg7kwMtNSunSUBxxHkIg
nbtjUnrjaSCBk7Hln3sFkwTsZb0bEJmdTnY+S5jufbJ3D6Q+WpDPekd+9Fl/i8nJBmn0EBnTBkwk
/xNTixJkzNX8u1QQF1p0/pAIGnc1q9ZO7esTXiIBg/pJJZeAICa4FnUFJxO9g0hbp2MB9L58mgJI
QLv8zYGfGmpJ81qp7eGEn9K6j0dA4PvWfEHgNr593MfAmmb1ouVHLF3xu1cb7faai4rHXu2hOrNe
4Q0Jawmz0XUVl4SvgfrKkY1IdYUv5Y3/JdAqalkT7Fi1abDAs8V2jW58mlvZTkdt5ufZIpkrAIHm
r1Rwfz2AX5c7NSuJxYyr07qWMcoUDPG5T9izYbpD8P6tBhTCiw1PuTwKLkKMXJCbC3irjLFYKMAr
nGUV1MYydU+4bAUstL4oOmF93C0XV3kulucf89jr1cixk+PjFfZisXqj7aK1akThEUmbHkD454Q+
PTquWv1R1t2m9eWUj0O3LBjhFXD/r3ictHNErXi3gUGOGMOYkdgKUu6+jwpIoCeUEA7fdJz7noFx
zqO7uZ15kmOuGdO2athLFpE8HZJCF+OrASiQ1EmU4X++W+B9IketCIbkZtoThLUmk66iMnD55QxO
LuVblm054IQSWDsQZNxh1dc6aC3TDd96vbz6hNlAHVU/l3gu2Fnv5P5QTswepZY5LIktmZ/swO+9
8lxgGziQ7RWFXR1FevDN1gomn+jrrhVmwwe6cNOthMM9LY7sMCA/5+WDj2Va9Y2quYKE6X6be63q
oQaa1xfu7YibRcVrKoRw5uJ6uebKc478DZhkJ5NgIT4X46w4UgOKy+zkkog4v1WnuHbzAc5fDdAg
dao5QsC5wDaoV2sKrRjF9jAZSHXo8YyJT6heCoX1V0ywLBwtM6sqH14gQfl967i3UjWdtCEf2nGD
yNsxHLKf1ksy7qTBf9JAMTWrNY7zfpJA2RlKYTfOG6L0y8SxxdrBR1G/mdvkSf8uqYy2Hyh4Qx9+
+vIk9rZn8t5ymL+VPsS50COWE7mI8gCwu8mZE2CfHBwJijX5tERn4rSROJQuAR9xMgy+yoibYUBX
r+Byq7OJD1v+u6T+cAHQ+26J/0LyzraL6P7ZTyZR4F3SZTKUM9JTsXY81Yk9u4Gl+klTijOfFaiF
mvhd1AXvS81NHBVqon1zkE8n2NiobaDGXRYu8hSeQ10AADgfOSPVyF9BzztdYHGvniS2fEJFkz2N
D0fX5LVAJR54707fFmCsLg73Amz4ZmCsmEotwkzaqGcYn4TGAs7IIE71ROhb1f5QFHbl5RbJSAd4
JM4415UV2c3VglSMTceTWqivTziLfxpfIieK+LfD/o/ac+8zq+kUZDP0DGaLsC45Di8nJ/6nnWtX
VOXV+nCXAxzUUJa0P+4TsdSk/oLPpiinOMuzDEk68dua2loCjMub6u35yIEDC/W2wWlGYr9/Itc/
2/Fim9ENuJRHhhyOcR34ehW56piEpcw+lJFBD+aSSl7kQmYKmmtIRYBMNYBSIIJ+Dl4kmcPdp3M6
BPxhzl1LmHGzdQAVDAyIRDkgzK50jCo+OtEnnvt/o/HV8gQzSCH2LETGM5Cq2NxQ1cC6z6O/n6bG
Ftr11s6gJRxrrzytJ0D7zJCqJ0ln9x/rKJ5uLuw0ku5Nl7SxUfkhY1CE7zqkFqPgBU0oPFoxflOM
o46DohZLNha0a09rm/OUKyOUGoEWzNTaQs78NNsz4PoKAOk2tFr6SJOF1+U8+o/tALYpIxkSDmed
GqJgUzCbLyRNtziwrtfgNtZhdd9rWIPoIAPFrYh006P6jm3WH6+WdCLaMoETpsSPYk0dMHblQXaV
OCCVwX30asiFfcVadVVI4HxPmCnMM5zsPVtPhyYNa25vyu50w7k+sAwUplj0myryCnVFLU6/QNR3
ULEydlo7hR7kVKYhne8bOLPzlb3h5XbqI/t7Yr0MJe2Gg6PMSyMYix/JuURzoLsi++DuQdJ/ke8c
oWTaKjzUA0Bbe6glTkUBFEFJXsU8b3g42FWT3bYThLTMQcGi+MhFNd3uOA8sz4FWpaZS72RLDDrC
tBLfPFizRQKMsIWyd0kGPi9iMVc12KqrTzhfYAXMbbj+a9GPDKEnQjh4efkUzMJOYBmlPX4Y57P/
XwbFs+CXWtzXxNJfIqeCvJj4xm0m6qWt6Gf/LJGqzsjzhEjjdozm/16FNofplJhqAk5+g+3EeHcl
J+jhZqx6FmPvaw6TUtQ4Wj1fUZrSxt72RNq2Ncl/J5AaJDcjNTItetAB9Jd9HZbGM+iwVta5QWOz
aIz/wcuyOqANDxGJjsX6/Ld1NKH97w2nHe7fsEsBDeavKlgbx1qaFIVYRUwQJJ9PjXqJ/3Lao1uN
m5dE04L1uqEwr/3P+2FDj0HwdhyjnyuoPGgRdXND8jIes8p89Ar6zwmf+6rSdqoj4B6qMhWiu80t
QSxGMESOtMjE/6OXti2NsHNO6CaW1Xh+JvspC3d2gt+Qil3LM6l7T/Jb72hYDsHCnBbNaP/P5J7y
CR/wU+oG6JNuZce2hOc40aFSauyapJ179dp20Hq3VCrpZ3UT9yDJDH2soTTqQ9t7P1wEBon2uHee
K9qp7m/uHLNlHuwvoVtWFdXvEfaRMKCOG75FDggWSke1om60ENBzEZbdvvZ0GBgOitwtbByCgr2K
VHI0XUw62lhluspO/LI3VZjOf/US+jNg6RzAiUSQGGaeAnXz1tc7puwn1EM2F2OplVPhnvzX4PIF
v5VYEHyjf1271vZDR8EbGJQVhvdU0eDaDA7Tf18PVKyJB/cbotwCiFh9e31gc69eynj0bhtPxWmq
jGJS6KRrJfQBFNAEvFeb/ELMyWH7F166ExL7D8XrbbUQMU4ldGRXL5lNlQpnxWYMpn+cJ9AHylR8
85WcDdyHV/ilRAcDzJ0man+vIQ4TwZueb23AqH0SnOenUX2dhVOfqRkLFLyISgxVcqi2eskE0/wS
MVbtCwnkfoGThsxPNRYilkR2H/feWNDnu3xOU9vp3QtvzFSHThIgH9mPxZrnRFY3ve3onx1hLz7l
G02haxuRkqhz4qsXCdgV275XeorLLJagT3tdZB0AMh4jEDrk8i307GqO9Chglvk6Jk5aWckvfBKB
bzLciYsrhslc5XxZzsY6f+jUqKgsixfbOOY4mGJ+8y1ty8QfgiFhVHi8bk15UdQ6WYSfosIv9nlx
v7kgqWSe3bkCmXTRO14sxE5P71HpRZN7JOjCRatm/R2zO1TEUnDioBEXgR4+aTrhKAQQWqKH8qxK
zpSZ7HlXRj5Xmyx1ehH81kwtHBh/9d+EYlDWL5fONVwcgz3knYo6GYgu+jg61THTODf6guf+E512
8WRuV3ya/skhsOWTlGSMfh4TMuLc4Le0OYLGq4O5XoMeVIMvyC0mvB7xYgZrd0vyzVMEadxUbtQv
/0dhHKQBJtPX1IslXj7XNbpQKwLO+ATA0n6XG28mW4ZkXSUMYOb2CszhOm8Rxn8fqG9NWEq7j2cF
pberKixZmCUE7CtGY43aOlXfbN09gmgai676rT4w2AvZHScTku7q3xeidFEK3BKZGOxR6hb8jgDx
GdT1YKJKKxwHVLJ5je3lEcwtcSo9xX4jW2hDqBkw/ysmPl1YWQ4dz/R5z7guRKR7Iu7VzcgpsdlC
mQ8twQ08/eaAKrfVMdlEscSxv1MqgobTj3mrDtP4t+FnuC4X5qhWQwiwzWPZs8yXYltLP1wY2ztP
TBapS7OGaiG2KctZYjsLTZiA5fFw9KUgMqxGYN62AVHefh/53UuHCMap3gk7woM3TXe28uGf503L
tTo3PhxpshAAEqs5K8/JhTMEel02QYVflweGKRGasM99irBCWczvdUqFbIrYw7Sr1z9qE2MqOuig
jedW4XoUmpxMDUgFIB6y3HHg+PSYjqykm5kDiTpgEgsBGKCNKc22N1irE0T+RcGwwPy4g/OmO7rv
AboA9M0JRK9Kfjl4HZYHvOXt9H7PPD+i0TR/avpXw8whRDcH2Bgt9x6zeUbVhsEMgYWRTDm6IrKD
/RvcVymP5lL9dJ+wP0ZGJOkxDF5ma/3+hwy4bT2MeYLvb+uSVx/s2ENamp0Yl2fTUewYcKpx2LZJ
6SQL/AvgRqCuBXoBaukL5Asw6omdQs1s/jf4QfPNYVLa/yEnaKvhD4lpVNOObo97wA8Ya24mUfYv
8GKP01NPXArO9QxkSSML3C3UgA6h1Ro4GBQCCUpOMtZxP6E+OFuZpsz0HRM+Y+rz359YNnHuX2PS
70ERfg6tuYYpPxczM0Ei6Z7Pi1i6DbmL7XfTmYNH9hlk56Jkf7+UkvXipeRsaujMcBVltCYTz10E
3J+dx7G4V0Ty1KHXAzG1vK4V5V4+i6uoGda27mUSBGrSTzryqEzkjhK1mh8ra4723eJq4ujha9wF
CZnAcSXnHNLQh0U6gDWThncZjNAOG/8aYr1x+mNyN2mw0FXoq7gSY0bKK3p9jidipV95OSBFnDHO
chOz5JgttjiXvpXPNYG6Npy5mQ/DFOuYulXrCU7Qrmew81AZGvgsSa6n/ur75AYeUGI6ypqFsh+R
8o1z10BTGMaqB/HKNdY/vvOhf8fViYHf1u1pHJzqJTiDBkFHRIhxa5a3r/DtYZTM4hNEAav70v8K
koZIAG9eH1T4MhiVvPuXxjFeQqR0xlD0HLk1jn7enR/0kyDf+MYqRKZmzKzCioFABnGRT4tVckH/
AjpcIw+VdET26LzyURDiyfzztPfNa7TS3390piV5OCb4QylwQtsUKARB781Kd/BFnaeLmbDXd+ph
yjfm1O3Dz2/+/+CX9HN93Fq5WSXIW6J1pobrme7k3SIao5i+dtUYvFqiHe+s+DAQfbpJQl+a+iBk
h9fS++6Qwwguk30wGpSTjwrDYGnq2nT5xsV0REkg3yhPVPbUFH1rRERWU9wKUPaj3iNNWInaoKHJ
mvFU2yTTIGFPwIYi7a97G69IOsiFDshs3dYWNPvIJOtEQYLwf6wtGszv59zj+fjmLOb/HShRIrs4
M57rioGe02wKj609sFGLM/if6d7spMq4WQFAdotodGepPfv1HyzdP/FylLxjqjS3Huf52uGBN+zj
3rz9/6+w7O6x6pbK9vQ9amlypzCCJNPlfI6/y2n944tey+UGqlX06tZ1Chkn9jAWJTEW55IBXYgB
PLt8H7IU2wN8yX3hiusbYlK7jM9IxoFdC24hMN4+AIB/J3kHwOi9GHeZRsNLR1Ifz02TdEuck/uW
ojfydLe6Gpw4uLwkpqbxgbhmaVzPWPs/6g0wX4oX58hgB1SUbaVKFN0UJ5CMp323IYtb5QQcDoqT
6oW2m4xJC1WCCVsuX1mbqzo5b8LjvpXi8F6KS86w8BMureiYqk+nBXsfaD6VWJYjtLTLXVJkhZVj
dxU3Roat0k2HU1H5qN6pjyTC5sCAPsWX4fyGTAfpW7opA+tdeR+BGv3R5oyIRDpaUxyQWqE/WiRT
4pe8q9p4kCi62r3ifSX93LKUfedkKa8tTIEyB8iKhwXhp02y5s4V2sboQMY9ksXyURymwYyvsYLx
TifJmoQqDU6Bg3iZ8N6L4VJY8bmA2qwMLk+UoRvH/nmGRiLS9wEyJl76CqVheRR3St0JZh4qRFVc
bzM1Vcdk6ba4hpE78hunK7s+PZgHAml5t+Gorthl/11si2S/dTwWlNsdu5DUY6fHxKT143dXGm7t
msRz0Cz3+Fntt8DXaxTxHHJo3Sr3+YR6WnpRFi4XOvAgIjYJxqXbThpNK+CeUHBqLHJ37ExdrON4
Kadpbb5o7FNZkixsv+bTuBliKT7efvW64lIT2p4f1z/yMvPGGPb6Gv8Z0XcS47oW4UgTylRfzDWz
T5VrQAB3db0fTyi48MIy6sMAP5NVpkFlxzEGLfodgisdoY8TeTE+fdAepX8VFB5Eu9p3kNwMBGE0
fbcN9eChvPfecud8RsI340klq0R0q1DenqzhJMmVo6OL4gXxgYHwvYg4L4xlC0Gy9i0tacSccvbo
SaI790FXi1rjVMb+tP4UuoenfhRY/DBvJngWnRXumPvR5zMWVtLr31RPnEsfausU4NSEEdAMqube
MhGn048G7h1Aw7NXyQLDslQVLWnaCo6sJd2r08XGaxqOoBtNNK/KZR7mgMeEb2xTSZZdvobSajmk
kuGWYDX1kFtLvVckFUgrYjVBR9OHWIiE5nuWUG2B5kNvrRp0W/gsACUXVc26zhJ/Ub8eijL5pOah
2zIgzYes9LgQh09ZXuFuHoUKbq8230EeIJ8XWYPX3qc1mAaksd7n9fSB1FdhYpURs0+R0t25aQlC
W+vb2WFKpmxq+tPn6L5YXOWO8iCYaQgyc/B///8ffFhGfA1pCYAimy5SKODf0A1QnCzxiUHEqFl3
iuZnustPP6uxnEylTHIUJlELSVjWeo4n6mbPDSVZIHnfBAVe0KN2IScLcBUOv8A1BeXBJAM8o/dE
GaE+my7pVlFf0vGeRAt0mCW5tFlkRnXx2nX/wLg1Jjf/wAzIU24GG3QC1t3aAC3wtgnoVFwk5Sx7
1vesB/Ty4yPGAtD7oX7OZtZhA/QgvvmpuTR6D1tdCa4K+L8uXCjvmYiVjPHU20+p42wR7cKvX0RB
yie6xNVabf8RFhYJlnOqxPlw1+5tKuPtog9x/Va3+iyGxnY4ckcJDNYf7Iy91NI7zcqRIINH520i
/x5X0RvgUXkyJ1xITa25IZ8riNHqtg7IHmozXgIRhG8vfuQni6eXkepTT8Ws3fzDCV4cq6ppKYvz
Ze5LlcKxOXviLfyeIBwvH3aNb8BViU9rf/yluOaOGcybkjaM4e0A+RuxWskXLrASku0k96aXCnsm
Qvw3DkmSrAL8flTvHidEl94VAQ8B+ABe5xi8r6dFeeo8K5qwyDtaRpNFRa4yparqiqmy/B2gQOkR
UM9jQEgHWGRovTut1gG15qs28e0f0FBnwvRFHjPm8fKgXkwzd1Fx7+MuScFV8Q6mAoqVIIANrdz0
pxsutNpPTVSwiOI2paugHuZfDCzHA1Av103DsOqQJjfNU6hK7aKWrAArR83N2gUt295jSPXwdMHN
461mqENxQoW9hGbsXZ2RtzhLGbMvyqw6LaMV61d9R7QVp0jIyC+42NQcGtRFYN1oibBVkHKwWbzJ
qaPunfijRgP3alB9NFqzswEaUHSf73CB7xQgr5UH1AlyIyI9RyPR3OQJKE9QkOEGk4zwnXuDdjxK
loV1+K3jiN2j+6x4mreGedV7wRD65+WWrUKqvhUQJf2hgqJsmILW5BPxL1Jjl87l0HFkI4DMMCmz
9tliVi3Z8V5v/QDxhmnZxZV4+XdxnLtZtcyyiqs6GaQAYMILRQn/G4gQif1wyMVUca6lP8CIqa1D
kT1l7PeHmYkmI0k4x4ZRfDqDdheuX+68oW0hPk9X42gztEyqHqSmZ24XqapFdnoVCcLVFwA33xuc
LjdTKdqP0bT2L0sLmTqu6H9OO8BrP3vKKKRzn+2+zSPivB25n+lm7XkRdXrOXAWNcL59Sg7vxKAE
PG1qgAE7EmJX0Kd+zqyRMRO+9s0LQbZSJdGHNwDhI4XxO0Txs2DK8ZfrsVkx/DS8uBHKHWQ9zQlZ
N3YWjK8pyhmVTPsjdsk4Cdbs7gY6PfKe2p8oTS64s8+NMMgNcVQAm4VX4/yi9IsEeCUF7Z2Zec/+
eUCdHQjO0xab26mZFlkuHkxubIuL08cfJ2kgGQ9CHZku+UlSlJNrlYGhKel4qZhSEVKkw0MAWACT
MtVezH+umQaCguCz7eUdAiLUCodAf5RjvhzxottkKkdGKiWgxG0xiYjNME0JXjuuSXkrw7ea6fmW
ej71NCUqphXObguw3EcCFrj8SA1wlEsJgNkzMXVgxCi8HWY+GQzE3QPFgxuXVcaFI8GFpo86Kxdw
+0Q2s6WcMf8zCyi+f3wZf+6yQW6jVBQRKJz+SVWIflLF30ihhTFwIwquUcAJ0cWm/5r+S8rfBWox
yg7XxYma5mb2V9oFxj1AC/f6ZNOSCteBasDl2Gf2Z5Z5nrXHV+lUUmVl3QO22OIFHYTita9hzjbW
0pGgLzzH+1kbOA0/tNqwvvJ6b+zRmHvYiLzFqPIhIE3rjXva2uODX9SYRvpzT+5JI7+XxIrA76xe
xnUflS3maUam2mslOlyjlB2lFD/mxc+0m8AIioxReJ2jnX0vbUbb5rJelk860QD/gueX4tKLtBec
8J6Mf/So51+FGflm16DUTzfY77/Ky2E8gnAkpA0INxuTMGGid9M9p03YPmVmkGPXnwZbeCu0wXuA
VofdUm0ttbq/SH45DPpE7jb+mxptp0QnBNkr6YIu+CmO3EZzUS/lAFpZUYvw02WwIKTlOJ+T2xCC
G2wuOWUpZ842b4VDikyTQ6PHvMKm026nVdHfdZb2BUnht9xjMdxk9j9EfWuqIohNUDJFNff/8otI
AOZJRIspj4AV3d8sDOtP3q4lpHzGL2QPVINE/MhWOm3G4uyCXkIkdYQhZnZ4vbeUWa9+58WCESMD
RjCUpjHPhMis8F3haT0jzklYuhCFJeGslvWrfYWPxGMbtvitaxTCxD5hUr5QMtVlUEmBNlxdBYAC
YjCawXPeYRmdR/TL6xJlIg23YdtcwRmKiK1idwTcE/+qkj26avib0NbB4lvPJMvVfI5T9cjXIkGj
zu0PvXlpmdedI12B5Oy6Z2+HHDTBQNgUzNr3B7iHl/WVM9WgUhSfMj/2a5iv95jXq/QRY44NEJZf
L/D89ihTBDa3FO42sH+qa4zml4FZioi0/pHyBCzyOErix6iuX1UgoAy0ciaWmS1msjs9F45TKdEB
hGf6pd0u5de9UAdJZf19KcvkiMu7Pgqe4pSNb5X8Sd38Zb3t57JuUmH+TYKlS+uQbpffsgOeSATU
g895JZ2TN5e0bJgAnH20YywcSrmPGDtHyNp2RNiUCmKfqLdpta2j2zmTA0TuAJzboyicEVs82C/j
vIWDW8EcN0mnewyXpM6kYT7KMOwq0rjHceuOQw/B8XApYNO1gtdO7gDguAFPeGGHP2Cbc039qPTl
orrrWP7Tyq7kAu5Gf1JV60ngun+4LAg6hiC6+vXX9xUOFNtFRe6ZT50pqpR7iiqRbp5Ja8ExZoqh
D0GqNfugaF/OCkc3dIK77Xy0u2OsW6/yU3Ysh5fUrxUvnHNW207xLuyxzVO+hptRt85PXgvIG48W
HekV7oan0rvP5zfFSjY6rq8hNiytcMH9/BIVPyNf0VhoNi42MSTXS5wVPVzx2dYvVe7zHegUVhGr
4Q+C3oS16eEyHcjbNj2P/aaPRoSCN0P3xjyZ845nQG9w2utzytF0JRR5vP43TuJ6k7uGcHfsvZ/3
555Wk9r53o2Aqz4R5OlO0iqcpxSVzpWHdBzSydaRe612LkedNsradaP1LGO2PhdAUn+4bhkUrf/x
fVwWcEPq/rREyEB67m7KhPFOosJdhFIeO+p5fQpeCKQ3IGXC7WxbUuKZD6TISAEogSsrNyfNlPuC
qPda9IG2R7ZYQJGYVneV2TeJr9jnbXFxcadndd3bkoxdcgVezGqHvJEPc+SxBs0lXTdrsPvhApHe
S0YWqZxcAENe5P67SkKmlzDqvf1Qj6jXo2J9OCYDTIBxz2VTHbeMjBSIVurzu2FvwoQOXjunU5au
F+cey3U3B6v8fh2knDw7CBg6aCNJNqSzyGyT3Uj6coXyIrP8QfHrtthvsXOK05UPkdCk3qRqLGxi
3my4gCPaUl8NWHgVFU60KIGmc99U3n13e7CjzfHsIMNpdE7c+dthIWbR7xYsozRip+qg5QaADDVV
JAd17wNbslvyfK0FN3pERcuFthGfM/y/f4ijdfZTDsrFDmUQx0er/EqHu7cejUfOsTcRomAxxX/c
jImu2eHoNL2ksR1mwlKZl+9RX8+zBUmaemxkxVWziSijIopSyQtJwTJIeMyJVI864SK2HkLSdQ1s
VW/jyUdVpnmxz65mSDPd9iXHjMAYwiqgfotx/ppXaM9DjCzKkD06LZt/I4RqxCAgzJHEXi43dgue
NYklEkOu652Qo70E8O3FWK0NWZS8/koAT0EIlWyID8trx+LO9ZktXk3P5UV1Mlljm1zBYWrzv0qS
/+xhtRUeC7AHPPq9/K9+d8CAdTufBwAdd+lS9sEQ5zwWB9oEHW/Mu83qmrVVi7UXPhUC5bnYVK5m
CuDJalqdwvepUG2HycbNrx+GFdz165is7EPMZc9vlIXSD5b3Zj/jmPlQOlHmoPnvl3fUQ7RuP6oe
1XrvcK+zwAN246g9Fpnq+mLm6cbQTpTkfeP4E5qY2xmxSBvU6Hi4V8ICyM9UhkaD6xNuZvshtuND
Yhl9XkJs0pYzhCwHwRgjCkSBt92/PrNajnY7OOTP7O03t+xbbF9KgXr3MajOwGbnwd4Ln8VTi13m
A/Zk8MiG4190g082Qk5ATm5eb8jgNugxqRWBCnb61T1lyYWyM+4AhVeHXJeyu0+tviMBEecmtRR4
wrWd0IRjsegVcr+DnbyMcf6YuIPp/HacLXi8EpixL0iMj1LCWN1o1Cn+3Wp0kqc5xopE5K/Wxege
mZvaRsLKNt20CQNDaQnWFf2WwMz1J4E9hlcvVUx1IrESlUePVvg21+x4LW9kZ3ueZDbw6sabtp7z
NAi9C89uYKyzLIIlgNz5DW3rTj8EJBJcEm3nRt7mXpX+y1bVhwLDUkUbh50lL5rmPlrVRfNz51Oa
KyYgFNeEmn7ypWP6fGHSozvOsb1IkDV0DQdBtxpka51jOK3p1QnAHvfoOv6NmDAtK061DFxCNFdE
UxMjjAPogIie7GvszhGiqrNBZ6LfR5ggFo6sEn62baA8Aax/9/wRMAHTXZmZVqWl/l+ukT2exXoI
CxAaW3X8j5/x41y8hW6Ktci+XnJ0i7++hAogwEOToG6G4dLNz0thyNKA98+rQtqi9ffkie5xYadU
hRhTehjKi9SXnHwbtDgZgDncj6CAYFtvkyhlueo/awtZMJ4pXlCjPDH2tHT9VripQQIMAgVup2wq
/QDpcwdBWV44z7b2c3XPNg5lfe2lBxYI7v85oTwsc82JoCNCX6fEgpMVlQzo5XNti6yxfCjzjfVV
zmwlPTfucRCjJEwuiaOv1AVB0j+dTrie+8WgytMK0ar64WAU0RcHgPTcShE0yO1TBA43u69LswyV
lpmVlr3uch7hmKEzsZOaLWd96hfNugafqRW5yo4bO6c4PRrTAdpdU5sk0D60VgDxuD2dZh3bl+ji
x05sIe10LEcASQp1zk25E1pwSRccnSqPpGoZGUA5hzd6ioFF+SYJdaeXychDwhQQwTXENT4iuoSv
o0WFB9TUOAx07F8MWpb9A/TBKa95h/k7AHpO3chBjpQbK2qHxh6wfIBa48TRgzGuVCyBXBfo4aEZ
y5mJbcIOvqwgszMAWc3Ol9RnwSOgke+IURS3a+YXUP/TgCf6WaiW6ALZTX7bFuEXTX7PUKE+yGtk
bf0DDI3RO+i1Pb+69gI/lw+K9Ls+ts6ZHfTgRkMILECvaMZT/y3DvD8vowtPZ9pPM5TWXDmiV7aa
5ZVNPow5nat5Hte60+r1ZUYeDIfKbup1gWZaN5Qp+th4eR6IsdtRmxTnwvQvXkXLI85d8slTUeZq
/vS6BwLXCZMctHdo8f5jivb/rAbFRxlU7ofHvili5eJ94hjOqfG241gNaKcwtyrgXsR2RpydxhX/
R17y6WmbqVOLblW6+UbUmVI3RcTerY8DjDSD6h8FrPQskNa7bOIgHAJbSx9BZp40ghxLyp/tauv/
rbSkGnYssKxHmPyy9A836r9bat06D0TWYVSpi944F8ZKSJc7kb4yR9lt5wBnmcMqotR9rXQNY2Xp
iwKUZEKJOzF1QfD3d6nZ7JJ2JMgTlUbGHOkNefOBHlA3FEaiKJL2C+HiW8TvvXR9pvJy0b+KhjL6
jv8P66W/TK7Nit7BqeW36nHllLMtVxjz1AS4DHnxr6zbpLL5cKms/Xkv9bAsAEUlQCCLzOR50KCv
fBocUBue0C8xQ9PFyX3TJCEkhEeM2JJ+QxEerKa+S0VDjydJVtZlAzBWm2XIok0LCHIZvkVGNwmn
CzFccIJBYCSbdVfqw9p5DChGHtgKYZndjin0BhhABI4pmmoFpy1hIvkWmkttzD0AuyQs3TrBOeLi
DcsK4rsSLeAo0Kjz9Md3TuzaWvZ7WdfApigDjm77CLPLdob04VzMWwBsBe7nCEnHI0mrzh7ABNqh
pcGjzgfv4MSYnNjgeT+e9zfdXj3i8ERVsUaQYPTTYqdjQLAgoE+aJDPlvx5gQ+GrZ3fj/66XA+xe
4qWkGNieIzq9YCUqlbCDABoOstF3DIPenuf0Z5n0dxj1rGYPfZ47INr6jo5dl03xJzT91XUFYeqr
1C93ybx23JIUgOPj88yQ+enda2K297PpQaRryazyjUvITakWbqUTMzFJ3zG9tvMzyuAtYyQbu438
GRTv2MQyEDoxlcwszYeEtrH6MBn9R7P0BHEDEzQIapqyMjQaa7yB5C6dixNRI1OBHn+f4B6a4qA1
dIJwS6nm7vYVVjw39XpM5FKpIME8MgOxy6WbqzmE5zrl/qc5i07bML63aELOIP2r1m2JxnHlqnYm
iEZRYVdIFmp/F83rQTrNZ48v4fm2MnRqUa/nk+dQBQ9vfLE0SpAvjzprsjYRxJlOnkQPHMtcOUiK
AWwxNwnITLKnEABJH8MelVKDky6AB/9i4UvYkzVTHVngoKi2T+UH5M4J4t6owDDBbbFo1jMSqexi
IjUGJzinpRwGgCm6kS5y9AinjWGWyQ/w38qyeYjoNzuLDDhUCmXAYVlJjifyVXdYs0b5rI8lZEzi
k3XWfxXodUfzoWVfoAJWPALxxlcKOS1mb83ZBuVHmqV6Ik23FLf0fPiWr+RKtAcdZCbdQEz+zIYO
XfR1Eo3Mpzsu/9Nq8jBbdSdgmQw66OUdurMEKt9O0l35YQQ1FkvCfFktpC9EfDcwOWo40dUDJmqi
hgAiVvXL1TpDOIKs1nHscN2vhADaSkblM+TH/hgZSfEph35s6s8w6bGKHNzXLLhqZoWT//vSLzNi
mb/yrlVrbMAwkXyT/kWYoeji80Nj7lx8QVsJjjNifWUN/+5mYYpmCVK3Ngr0Rv0W7O9i9gvVH5Yq
g/1PyRZ7liglmZnRgWWDg7WMT0iptbJAg0rRR3NSv47RirOd/EpAQBIL9/+4h03jJ88OLVhj+3x1
U2smfuwWu7tckcwcqOVzG5ay8GHYvsiUE7PWllkLU0USDEqAWKf5Psx/fSVN975moTz7tZxpmpeH
aXWRGR5wsQS8ND17//4pNV0GnyZSyRntFXVyOXaMV57f9wIEfPjzKM19IoJjCpCSRkiaV4qecweQ
1VsUXRhwBcZ+yt3Xk1s1efwg5+BkqKTdIe6rR4dutBXLWpJBdsN5UZfney0ljX51MnGn1chf8IOa
xJR8D/KH9EDWNLNxdT6SjlhkfYcCJsG01m5WmSKN5jiNl73v3wXR8saJlhDMWWzrEQj57WLYPgW6
AMICsN9iRCO4e/CovUKlpLaX3lfRXHgd2Xouu0/4qxxkuc3e5tng1NNvYSzImB5QDWafsYZR3Ik5
SOaAXs7hsZDfK4YmMz6t4q4KeSTonkDO5m/c3JrpFHJpnr6knEvTv7bT4hGDvNfX5yvYHJz18Q7k
jZU9GOAkAkKAt9n5SmO7q+c1c2NogcYZ81SQpNbEu9D0H8rBmL+jnpZsHpQ8LCXVzXL5iuUcJz7s
6b9XH1JOYgq+TL5tTBgT4tJ2KzInkkAY5VtlQgXUrYQiLfh9m0D3QiDO/8oX00wuejj+kZGGJkI6
YqqduzJrrUnSf5j2lbVlZ4/rLetVuTNHMYfGfwFw4UT9timgy3MJDYhCmQYAI0XgwU/DnI5hT3kG
BOzTr10U9JjAhemBuoHiabWLCiLRT9VD8wv9TG3dlM1Ez0qAZ/HO2PADFifTjMldDRqaYihH+crA
HGqKV2hvIepnRnfVwlLiZVazkpeubiqhC6qxdc8BfFIZd9qXGVovTaqRcWnlem/0aQpnyf52r1wK
Wxjv55L5ifuU5t+z85c+BM4+q25VCwUdoKfz7W7OXMQKrUNRGQ4lP6/T0i+yFNOGQugcSd1qU5nR
NTC0QVe4WKLUdnAu7bzhCMF8s8QDFaWCYdCazt4IKMl+bOo+fGOXsf3m6hpEgg2WrWRCFwXx+tFI
oaasHx5pgi3GU/oV2LklqKPmkJr2+6zlBw6s90ecPjvHwh7yRTZhlJEtzFMUfWSyZ6hjcvcubfFb
0C3aKRqH3j3h+hqqIO9dUPYoGU/gSXYDdpqCdPmpBsrIBQ7E+yim5Q8y3dLLVaxfmSD0Ny4DbWG3
+6OKRw3/t9ME4d4jtMKBjPeuyfRN9628js1v+RcA1BJ5OoEw6drZgzEzEBIehMSe9VeeApkvqV5Z
mq3H7KUVJKBL2vMcMojRq36D1mZNoZvDNpLhx7FodJH7Eiz1L2n3aZdmSShLY0dD1cgNg/SDqKVr
lmv5v84esieHI8X5Pclz0rLju5EmiFY8uie7mshV4DDZPNpbhwEaGvp9d18B0hsqQ5JP6VcMHv0V
RD+gc0BMjQH/9xzICgUBMG12P7f5EbISRdRIO/VyJbIll3fAnMjXn9zCne9rblgT+wTh/VogPmX2
dsC6/Q0F1vVcmFDb51P7X6XiFwgeMqN42qPChaSQRke9zSdA6eV9WfkfX2DIiv2xDe3Pqw4wyC5r
8sJ/GpiB9Ka0N+rxGH0hPqhp0xlCkYlHTuOt6lJwk0caOnH1kDciJiBTtEU+rUOVkkMwzEj8I0Nj
XUOLZBM5jTS0FuTY5iqMg1a5bE2GRwjOL6z4ilun9FPOSidU0ZadlrXVrEPe6W1hlL6uPu6xBw5P
sKTeRmHfUNaNrP0uBIkjDQHAZ8mZgtqJ2g2cn2Rc0If225Xf5q+QSmvUByWhDefU0+SMYKTNVwyo
gPwGQE637tT/GVkkYFJSdwQpV6uKKs3jjrJJbglBPZ7FTU84RjBbe+Z+sDqmNRL3LftLweXmaWXc
bkD6+EZWYIPuSDCHr5mGhBVZk7y1NgtEcTaLeEbFz2ut7KZKnkqkcmTT5HVlhqhokbkDsySOtbUf
0UNsjdf9TD7ivBTDc/+FgvjEnEOy4GR2gG5i8/Zc0rlIye2VnHQVd8dRXcL7bgAEDho568XkYVDn
9Q42MjInjXAw1Hzy0PZHK/RD+/JX8Ka9+mjabPcl3G+l3Qju7EmkFyvLXzOvc3lxFQ/GiZK/sXXy
2EREmuSZDJYJgQv1sHu/BRiq6aCCd5guge5Ob5wREpaboyKbkWRIzCif16m9/KMfxO7dsE5ktsFn
canIRdcChkuIHzI3YyqiOTCOymiwjQ9lhxWeQCjPA9BevPhBSEPgdgz4KVB0mZ678rx6X6dD6ocR
jiOOnebMr+BkkAI8Jb1CA2XTHfVvcJQtDMj+hUwQKcLK1BqULZYM03lhFHzpfo0rIDBxAarMdK9c
tPbWkBgFpzEHhdfCMNbh1v8k3lkNz8ELwY87kj1SlLtbpLZBzhSTt/Xl54eSMqGe/OiVS+CTI0ze
uMHWIUkJwcaVrthGq15Ww02mpB5O32yV0WIAdI8+k8yMBtM4cBL0px+VE7OqDL0gf8gWszWd1Fas
yZrGGQjYQSRB/dM5j4MiiPoi8DjI4DKwSqxJUA4lUMKWCoq0eQD6pXlniwbcJBZyohACAudaKaEE
v/HEJD1+6Ryu6lwCH4EcBjqTzoEXCF1cGGQ/yETmoLdnjtqsJ2FIKzsXNvPMxouuM7FV/XCJnDQz
NRgK8tBBVm7VpBnrt8SrZDvSq6lmr5IZwGm3D7Ex4U81UpVooECyWCb2tcL7Y1i0WZRSe9JIpM6O
5yByVsIT4B0782Ajkw5ySP1yX58BJyVx6mttmTLcrXgSsJylKsfxTYvXr/R+oYQrONHM/AhCv59s
VnKMqZ+FgvmOXEhhUiXVot2KW4IiUOUlRzBb1PIsTcsYPXo6JSBvgiRErqk3igoxT2oemT4CtFmQ
7s0KHsr/pf/w+SRZwY93kzKHn3yBwNwn19nKuo0v71EYtGU6T78rifZLU4pl2j/Dk+feZvi1DdEN
lasbdIfRYk84o191ztvec2TPZEmwbHEYDZ7rCgytnA6nA6qZeJphxvnPoGL+RPAIsSi2U1yc8lwf
i6HQFNrT+0dEMzntf+3tiQ91T3RCCwk/9WN4FxfqdDKMeI5712yJtVnlpV/0Dbj+e5a8y8s71fOj
+vro7o1ddfRsU3m2aQd9FZWodzDX9b2Hh4igqEd/zCrlP7q7MMQvTeeOTimxALQj8pA49ZWas0Fa
L6Q3hUSxnxUIy/U0p8eHIlvAG5lLqcNCzOr/JvnxSCRZWNtRcU19goavNxmIvszdm2J9ZWt7S0BO
8vDXzjpglaAjWSUa2PYpA3FyRRc213wDuEUvPwR6JbY12hUYVvDtN1hsu8siRqoXmRGLZp+4Qwu3
Mh//KRZmfW3xCRa88MejVCuWXYl/z1c34yrzMQnB8GDm16zAGkhBapMKQUvzI1PTdlqYYubJwYag
faYGKqeZamIYJi9+2r+XD+AqAaEmtMpjm+CivO2SbC3TtQLGVpYbdiJmpFxwGNO4q1yVYJlEHwov
g10XWjfU9DA5Yf4cYAVbvXT8IYaYDEc98YM24HFzpJZ3gAys1Ljfsudy2YgYVdQYO1nkq6hVOrlC
xqoaAyPXAj+WyDsxer6EMjQqtfPRHil1G90v/a3SGMDV72/wZsGi0IKTujp19+gDqC0JfAXfPBQM
OilEvXAvPyJVeFCRioh5Dvms6rbf5lM6mB6zxUNccZUZtj4ANMWL7B0JvbeM4OYLizASmtmzd6Gv
oQTFl3L4If4vcrdVpULqSd4gxDzuCUNSuYZxAxnzMM1VMZtpdpSoPEMQKobS1H2NU9keakvwtTbI
8vJ64K1ZkicFTyK0L63//GtPrHS/lfqq5GnyMcjGYC+kz3ZcDRBb1rqMcRjC9FWF0akILA4qIhhA
BJS84ZPUDaFgNykGpediiV4cMp8YUFon/ua3zk1ltz+NwsSFyPgmeOzBAfAllQN6i4MqRRtuBhXO
VdN2LLp1AXH3EFf8IDHB0cp+lpYNU6o0m+9RhD2/ZZMHF0xagW8eQM8ZtKd5w4E132qDfUXLj4gk
lRMRArDfV7rUX9PbYt5ecCXLWGeRdtq9nOjY8GFGiujNNBGLQ+NTy2yUcsyOvWnPU6AAapp9MIrp
idYVVq6YLRPE7CBnH9Lf32MuwzDlBVWPMlRr5nu0SL7HnG+deCzEuF6cjLSKiYBeFnc4U+0UfNkb
si1okdaD8LDuEb/Q8Rqy1Aa5LUarkBy8rgQZwQq+cGWjdWjlw5pidhpXchwnsF00X7yL4ivPCg0E
1Gri1jNqlPCKdkpGogv3fbC/uCoqrRtBM3F2wb40LmcnQ3nkbXjFH8w1dpf2iJ7OxdmDWGBY6bc/
Rl46fVWlYnqEvrZWkp8jIeGLW1HVO9BaCCsn0Yctf1nGvqF8Bcz4c59t1UbUUNq5PHbkAMCMENLX
vt3XNHPiEQFUXd2MOU6R1dL3fgWZ75jJarvTq2U1O1Af9zjtMQntLd3VCo5WPZfP4CIwyBhnYGQ6
2BMJdB1XuPoWj0wQpRQPU6Y+GvT90mylNdkGPxW1+yBKL2sEdVe7bBmR98sG2cbhibLxarLOzP+h
IgPtP10zXn+7Hq7phFt8KLe409Uv/V6LaVNsEQuauTSyJNkrdwbnuNL6HrhMHOFyey11dG2VsOfk
+32zYlYkcEZBeCv5hah06YVe4TRb7sq+h3Vpbia2+6SAxkqEXykdmdFLoVwJGiWT4qgPZPxjm13E
nZdiDypylJ3IF46a3gPAfbRSLj5Lg2635sauRWl5XWXPZLtNwUuD9iAoiTaiuTGAMcgE46mV9XmD
UFpbZYRtJJfmWZ+1ex8+yr0YewpfQgZoglrlUbHrb9jDTyVJ7iFYJ+xJCrHImtkQ0UnJUc73IrBM
ncXCm389jKSXIN/wOgklmyT2OSRchpdY6EfZk11XU7X6nqPxLm5ySJLOGWatgGxOXI4abSlhF0Et
29tTKMrfIrKyJJShkgMo/ZXFJ77IPH9lqSiruwTj8QjOSPjrT14Phb+7A6HUV7rJ4L38Ak1OA3vP
T/Fy9ICuLo95g9cVaUmXiDe9lqCWQGvTOj7h2YWcjfxqYc5KsYMnMWMyy5E+1QTGgel9W8rleLhP
qT9bWJ+tx/XmvlslfWvvM3ijT6+gY+fTXUGcqlhoMgw8HisB4++4hBqCwnjCYJ4ZmpIcS3j3KHsm
gUdAVCD7XnHOxQjqDdvtKmZPzQnXJYjHmZYqEDTSFWMlDq3i0+zaLn4q/DgRzDgkxFwDHpDUPvtx
Pi1coRVpRAgTr5Dfk7UXtAGqfGgWyjmgyhknUWTTlcT8uEBR6u9G3oQtknO0rw2HAz4jJZ6MJ7EZ
ooXd5XzhemLYmsMQTqyiavzN7ok9wkf4O6Fhph0rkN4nGY6TuUVFUfkuOp6PjXPRrA9I7uPOdUmD
g0Lq5fW1+F8hTmRNXdoJnW/v7CSXvfX9x30IBU1QaC1OBJDS9xMm3+otPzpEC6jyFuBO+nmzf1Bu
UThcPIWXcVW4kIuo9RQT1Y0THrG6RVdUQXHtjhC8tPbbEjhYfulx+h/lF0hk6uG2S7f5JkjU9MNq
n9LEBVgTtpFX4MrUuZIFfmseifrM4L3EjMTyIpQ2Pa4zXFNrQMe28G+fDw+3IN1Mj73XxUtyB+L2
M/Q/QQ5stkeSTIHOQKKM/rwtMwQh9RkXzwA4r5fz/EqoWNtIatQ/oe9bnZFRG2Yo+A8hpZM003S/
b0krieQED5bgj8GlRqr/ehDqYKMi0IlbzQ9OdNZF4eouOSUzx3HWFVyu8uc6ZbMse3gL3ax+VLqt
UoOdQYU8XT4pSATFtB3Ky2xM1E82GGvAFNT4pERRq02y8z656ZwW7vj+0zlfIB2HmNsy7Qm67OGw
KAH5Icmzs6UxkTQHmBKq7LeMRoI0SB8bSJm87ZW6K2IdGBqQc/DUQy1FckgDD+Ra4J5uYPw+pWtP
qNMijLyn9NgdgdzzpNp5bO6VNo07d3I49xp9/ndNhXfUQ8c9RSLDCvVcSSDVpI5BYXDsBmwuJlDd
64Y9RWByTnxg41r/FziqyqAyJvUMgDA2+FfRSkaMn/6a070a2p0wl+PS9gHCnMRAJCih/cAKYNXV
oHmH+LRJctuKk3hnFf55HpBhszs6mwLHIB8SolSc907euUSc4HBED+TfVkFXPfSb4P56NC4ly2gK
A2Pg9yqfMcazMk7JprSiJFmOJPRwS7yk+nSnKyGnWN8J2jn6FY96bDKkySnjLzJ26PMq6KpsdhLL
eiYU0VqeaPK+jScc1WB8LO2pOGMuJ1kVTHUqI35K4yVY3E+Ts7SYUP76utAYev+WlFSj0lKmKjX7
jvMsLEYndvRmu6yFJrNrR9+miTEiFxYGHAEgSMgaj0GzTsyZLlymL+wdzDW+ZmWxXAL5R53y6BQm
IG1RXRHc6wG5vJO4yiC3s2hxDr4P6ynCK1sefISzvIa764UPEVe/NmbieaFo2TNE3LgvecQLmBA1
AT20vpcrPyuuRww/9+iamdEUYGeWG1eQmIYO8wTLYx6fukokd89hRSw7f7+LxmPwH99utn0HlPoO
8a5neRxBWilxH2a00zAnAFM+8gEv6VyWzCdmOxe54fI17E5/J8Q5b7jzmLXPEdPZ+4MvY7FMlAZi
69dX2l14chLuE1kNavUBZJPlWShOC7Q4uYOasXcYSR7ITjIQLhlwQzhRj82JInq4qLVGJfAqxeqU
PoA0xE6fIIPVzrkFWit9m1T8K2sPdaj5AeFOV4yJMkwMEQVifKMi008TEpL/l+Z+i3cAikzDKxY5
s8SGAlv87vZKG+5/LzhNtbI8iwH4LrXm8XMNzZo46ZArXHByLXtQmI7oOYfsbRzGwGznm2qQ4d9I
wwxnVcJbaBZFTZOuC2F8Wak0B4khAnicWqzYYVKKGnuZgHtM1aPHy9Nb9oJcohcGVtrA++6r2+kb
WHyn87+iiHog+zVr2+aq02x0b9vKQTJ2NMX72uTaCL1vdRmZ+DKXK/MbkJkjq1yPr8EmUcKqmMf/
n6s8+8OdAhZYvwWombTIwgPav5GfyzI73QI07LrHNPbwVTCiycevI5DVphTFuU32nefUCkJgOCv8
lJMltee4FhkZRF+0K5jZiueFIsVmgqx6m3aWpd/gqSs8d6KBaIXG5MxRPUKco9s+NzYBjwtHghrV
GvvxQpjL67uLFd12Sc41hXP4mtkZgVRPmoY6OG2kQmmYEmyu8b3qTXqExMjSpAX3QuleDrRfMMTy
iMJ5/aK6EjtgRPnRZha5qeDc6H1E76VL7Z3w18Txn/qRHWlNAbPRPhbXa1Uq9dKAdeTxQKX50o9G
vc/TD7DSkZkIIlFzSCLsfjLX1bUWJ3aX1Z0w9HXFf0XC1sZDTcbi1nV/JhYsqNmBD99ND0yPAD02
iIPT6UQugIDjhnV8WijBfnmaCZeCPEfjaX5HrgriY41hawJm8KbSef4nW/MgcJHIPbZ7lq/esOxz
fzHnYsNH2tf+0vucpTb+4zfiRNzJ9yAksIHTGE6BFalir+C7dNs8hySUlaxFj9J3k1htOngD7g0m
AI181h2IpLtiTNroumf+TeO+xiNweiazXD85kfUrY8HQBen1F8hkvyo2IwVhCbUnPv/yn2QxQ3xJ
Du5iYwiyQ7yE0UucBZSXvenb6FKoL27Pvc12msxCLPqE3NZBbdF4ZGHJccguMIypDnnKiE132/1B
HgUzhkWkBW5uDswUIY5+A9G4hg23KwVQOnPP01NoSCTIiuVTHX9ZMegkQ3Ks6hokimghR6vcnpSj
io/cVRCausaMwsUv64e+TFhuuNsI2y9oTDZW0Ck3cgSLRfAtZhjQ8KQ3ThvnccR0YPF6PYM2izyK
Gz5WK3QvfxJ+A3CxUyXYmJHmq6MZtQS9VrkeWw3Aptw8r6dCwhXVWs5PcBAjeG835GGXimEYhXF1
cRj6KmdcdFawaq0zDTCiPn1C4mbEhQvnlAdbtdv1yt4bo04szp3/enGbzpZFlFOEtgRoEI3iQYdD
sYUOcpK73iT4VDswdgCX+F7n8v2VPsWWJJaI53Z7fBGgzw6v47hM/jjL75c5kl+honib8Q3C3aXX
aUrM0vF5f0i6kjpIxDd1AtFo901RCoKvRsgjdaBLiCizKkvUJRWDOrBlBtcaUzhGSYHPsOflSLv5
WwKBvWjpwq98YTCKc+nPHjb8jClxBmwqa2J0/Q4iJfQNbnC/0Iwp1MHa6TI+xreZHgfCUVAfcE7E
KmjE33+HwVFB0MO3xFah57Q/MoghWVwHIKw8S7gvZGmTmE9izH8eJrqjseE+WjZyzThNfdg0J+e+
J5PydVKl4o1KVoH14xt//GUO4EJzUzPmcQkjSRyko0EyS89nYUdRcpE/NhZABrnALNIXV8sbYFcb
0Z10s6cgu54/EI4u3FI16ME15LfPQOc5h4PoWUxhlzb+nGvqkIwEMgUvF/XXvBcxCqOe2C4PtXg5
G+Ad8vSUpwwvH9i4ONm2RZyXNKQteavhe4A1eDKmleqw+9Y0Qvjs15GwHrIFztlRdDaTcyvhT7En
iCau8EQ5YWy12T7B8Pm68Y7MjFkbPXa1ld5P+pU8z9aBzdHNVzF84bTHI6uKuipi7+PgCBkJPZgV
AzmgJ/fG2V8gVrXDPmbWjWx9HTlnwHw3WhQerIz+VaIBtCpgb5IcevzYs9unVfXSXEddALzCSTZo
AWdOWc12QPnMmRem1U3c8kuMk4o0mIrjgxFKiGyuXgYlUuFHNJqz2qv2BnZLw7vINzkhOBgw9Orr
f9ZrC5mqVhgrHVi4l5Buqb3DaFZBlv0BMi60R3ZVCG7AWDNffm46UWPIXgjMeloRWftMRyYMGbCe
P8rCfvMsHPyWYAeWT5BWuqVzGarAvNV2yEFfQ3FZAx1mWsaA14w6T1iP+aPEhlBBiNuubTEajwLD
xVps490OWf5whfdZRjWBzDX1Hyv64YLfUWiVSmuX/I+vQbDLuaITSKQUIPD4FcQ5V4MX/DfujWIR
z5anEMnxO4CiKzeS9G8ea1Zzo/pY1yMX1nEDhq1Rchl+NNuNVpiT7BJRQqbcXWfrk00h7S8dE2bZ
pEwm2a8DRcBMXXv9qMlJCj6EFcQqjShIiZITiMP9GfR5fIgU4uC82kDOIGBx5Ib7zxYkLX5yLnJ5
UGn4A3ACs5YjOu9hB/dXy5W8JBk8X0DVYLL51rA6w3yWy5kyzpg5z5nv9vutCzGpwR9HxR4bLI7c
bpoRKjLT0KP0ghhumVrWS3Y2tCZKM8Gm8yD+mqfMEtAuxMAxObtGQ8y+wxBz3TNRRFxgwk42S+Uo
AqryQdXayUrDvi75FVgvSeGvbZ8kX5++njILFpkDzapYbD107qd3HiGaQx5wPl5V+oufoWZQcmTj
bpB2N7M4+6nbTfaoQYUqKEog6CVGZNYCJRr55u0Dk6llB0vFRaS5TlT2Cya14Gu9zjErTntVyG/J
9LONvlCG2629uURcKtx0/43kWYZkrCc+5F4ybUv7mYMnl3deqcuTGxdg29f4mTPkng2hpFUrE1EG
9MitAle9jXieGhhfUSOCFauy4WYoGuh4OiaUDFgIuPbR+dxOFo7d62VAdMvBuR65q00tR4+9Zbpj
8Dhg7YNuXPA6fAk1AxOzy3M0LmmA7YCKtSvgn6gyQU5/iV7nn7kJNEQvgGSufWMXajbSsgidqTXy
wW7HJwVBGx7NGcp0ADn0Txl+oWLa8b1XEFkftsb9SSmCKRClHiPUewtwpAfjHc2U7nzuxW3RkeQh
lMK78J1OZ1AxPotG9KBz278iEOVlbewE1dwurtHJW2zqMJt9VqFvoTYZs+/VeHwldMMhTBjkJQ5E
k+uSqmzLHV7kPuEn7kzI8Ny9KLZFvRo1BOR5Ode//qO769TBY88DOlQ6byEznW3qMBTRbuOcTeZc
4fu/rUUu//8TP4gX0DSP00JVBiY5gZUAC+pfFXM0/fXlHmT4GtlWDUcQLOCX5nTOCGNjj/y/dadX
mBJ03qIm2DgZUkIfSQtWpWQmr1qW1jG3Oe2LesqUHLtYxWJZyNJ475F+lwOoIe+B9tETiXY95YDO
8tRlwUUxsrMWItyx5wzC3iu+vw4HO51BoNZr6uTQfb3kMisxgmgYrvlKl44hnDY3NafumqcGSFxI
CxT5cR4dhooTrbHImA8ugR7224ZgQVdT6sDLHIscMag2xs09EyRtfu1UepSwSd8FwPtZjj2C3V5k
9/3KPfljIyLKF37fWSeeIJnmHz+0rad56NsBT+e+gnmQqeY6/Xl47EI0psV96XrlR9v8U38eZo+7
BqKhKlaVeZwzEmq6+dOThlTVtpuYG0RALQZPb2TobbCB1RaOcPOMoYyWB8c0d0m86zyJ1HrUptER
5fscQlRfJix1kK4ILBWwk+zwV9+oWWBv35FA5EgdbhuvlIXfDJVOJe2Q+S1lxg8VsTt60Dp3EVjG
PpzCB6JmYXT9Sxd3pTeT8y/9V2x7flw3YN8neqla+KrVOepzkKe8EGsPs3CKGVVvwM5Dq3aQsb0r
Bisw7U2Xi5e2qd/lhPZAqmGfPe4wzzi0fTJDtNn4z62CdvwuMbhm3coZCpyR2A5XF6BWr9AK/8Um
DVm5eyfxMpPuTmYz60GQt34Rt8pTxaTLvRIMmr+lc8L/PZd3UmlUf8S3XiO+7Ke8b3YraYrkHTLC
7E5KT9nPxEnU9EBHWs17H7d7MF83nQb2VDS/ZoXJstFjNx+7WkZg3F+WK+h48U9LQzG9DVz1SLqa
hVmNzxuCZI1t5GuS3lUzPTtWqOq6uxU2hDXO7PwY4Ia2wtcduqaSBqHpalDlFlYbX7NXiaa8Wwpt
mWre3yNg7WXjYYZ5QECrCq1Qx563vG6Pt5FoMTkwHvZCHKt/A/9EoAdfDsMT+vA8l+0SO8b9sq8j
U2UoAVfwHSAk9nQb66Y+8XizAQfLtdNeqFpjm4uoh+U/SbYdM8Af9M3TTJvIdda/geSC5a9VIXAR
uY3v6vpxEkKTyVcbHsICP5MGCmq6i64hvt1sCpoCJ11JMYYMfoidP97bb3F2Pf+yxkBW0+1mMmuJ
/qhIileLtg+GHBf/2JTTXL6/iW94J/xmQv8XdQPL62LMI1XiW/CsP0Utj1nM+Ingj0q49TftjQ+p
zy3uobg/eNf1eiyrfjs0bqe5Rwx616yDrCd9F/yimcKCQY7l13i4HUJU2LPnTu2CckKKhQBRQnV0
6OQSgk1vBrByWrOA6J4a+I7lPzWYQqoQGZaaDGDh8m+wf2Q+WgBghkL6m8XaLHIm4x9dsFvbzlyq
+p8BFCDzOBJY8J12CgpNHiblqWtpHyQgzm9obvuhm45Bswv1Kmol4O70sjqHUNGHjFVrHRYRhhrF
Pr84DXIV1jf+NAm/S0UaNJKXHDEIBRugmQntUpaXvCDJ6hBu9XfdgUjMEFgYYejaTPxHNvMPNMvv
k92Jn4Wn+boZoRZYUc3xMwpoL4mKazcIK8cgvzPRbemF0Os/ZUrmAIIg82MZxEd19J4O4Qkp1Yug
Z6rVRgUGUb7XqVIJGRxpxvXmfWfrH3aOoGCuB/weHnoxYKxGUM04xx/75lyf73UrNq8ijml0KN5+
gOh1D39zRM9mviKPP3EenlyZQogHQj8XdhGi+E0ko80cPm7fNq/WmK0S0zru0h8dUQKKvHceuA0Y
pD+4uUdMElqPRiVeY66pe+/cUCw1azd5jS8iaUeOUcK00M6QOLIGJYuICPR06DFRDCdVi9ZqRmb3
nacy15N1PKHXqjwa8BwYbrG8/1oatFvSxNh8bU2oDCmu6VcbL/dUvYlr7OV6kecazcHmaTuqiVmE
K03rpCRZJgtmQqzt4jTNxSYJ5OwwLjhsbIFuyaxN400ZNIdoKbjDviIY/3ughYaH5/QKuXU+/M23
G9volIjyaOTSAZYazyurDJbZapJ7iivprA2NtP6CQjZlSKtQkuOCpZBseP1lphK+8LzDMWqiXP1X
ecUT8Bnff7pigAcb0Kn7hrPgIbnVXUSo4EIsCaR8CgZNxgMsE+5MTGu6maPCkdrqS3HjtDLIQ2ig
m9aMjLWozwZvRBlRwaoxB/vh2RpyPSpPj4RKsJu+m4IeHeN5F6C1bgT36VxrtcrQIt5Q/7p2hf5p
Aek0bRnuTrHk/+bd19U/6MRr5XaUJbgrzN9v0sC2UEvd+IiaDbDkYVtY8Li6CQak+pgOMQnZTFLT
1ehFAHYbsWRBJxu9ZLJ6idMzGihDOt0oZsxYHnzp5tadSrUbHW8nqreYMdPN1SyfGmQDXAFbUaLO
EyGVHV+GpHm0t1uJ60USBNLHLWzNxO4f0wIZigjge8OxegQrwOda7VuH0IN31lB30Uhc0uXo0GWu
maMH5LPekKCcBiVfRaSFW/VVTUKxDrJFKyySBNVMFEW9dKnfV+QHKpzQEEMZ9+stWibf/z+L5w8l
Stc1bAgP6XiZfSz4DmjFk9C5vRtUSynfFUUqEDDzN2PA7sYlMu3Hw0EBoDLw8gcYpM72uRzMurfN
tJ/7UcD/zZ1YcZ0athJsmfZrm5iCPfHJKb1+TL3wgeAnxSZAEamXONJKGxgK5HN+T2V9o1K0UYk+
4JnIJjj9EIsNOqpA65gvLCuXVszsdujpHAGhqFX6zMOfxmmvhI4rPwzP5KobfGPYucIcHOX963/t
Za9FDUEoFPrAxuZxjpxR1Z9Lqmd3WgGby0QaE/s+AlXWXhbq96l0M0MJy04x7ZBqAEJUFdZK68dP
deh+BPPz4SMtkEu8amY8ftUPkknNqVCgRbuyXX+1BWYIL/UK8O7hro2dF7SeKpDhdHddTvKh1hsK
k4EFDW79YJioSvxAjxgIUPbRAZQYKZTMnX6HsnMePlkYadi3Jg65BtWA9kP+9US1a+f03/Q9osK5
EOfr8hZVSqQD/324UnIFwUdPYJc3JI9wtmSgoKiz3dn8PuZYRsEIICoHn3X91WSmoqF4NH0ZxSRq
mTO37BgCuncyO67zx4TeZeTAVMc+ROsmv11jdH15nu93DTl9pQgVrZurvhcQcaUY/rZUqmwltX90
pNB/LQ8ARxQQdR4VMK9JeU94IiE9AnlcQ2LO9iqn/Vj+r2YX4wvHdt2L+e1H3QxVjWH6E4Dh+OL/
wOC4ffaUlxhObZGo9wNohS0zQVVGvX0xmlrU85Lyg1OEm+X1J/4EdXpyoiDZhmnQZitj2obc+QiM
KaRNF2CN0DjvJ7tt6X2FBmmZknUwZXmd/lXCpee4MuhUMAgatTRB97KQKotA98x6znd02/ykeFtQ
061mDj/Qss680sYjWDUgjf9nUEFkoRivB5Om2PN3UE00HIzpj3eeTtb3wqpaqHpn9BENhbmI98QW
XB8IYcQG3RhiTNkUB2p34BAKGAAlPmdJ/NYzeUfP8eVSFzDmL9TqOXCs5pYzCcqkEoZN7PZYidh7
FzsUP2i7NajbNqUXnAYDpTz+DlItp6JMIlKo2uShiRHq3LCEDBX0qshZDs6KKV3F137sc8hDObTC
7PvsNFXpk4Idyl+w0O94R9SaBdiEqonb1Y9lrpG1Imn08odtmCsrZdY2ft2qvd/kVd3m0Tk/uWff
M5fJzymfhebPFbqa2s74zmE6zUylg9v2T6XWIHuqb8wBkX9cRoIJGAbGUXZzw5knTajvwTNkNEzV
LZ0g6dY4XNUu77/ha8foYt5G+ZELWSK+whpA3OeqZheh1BVviUp/GWy2Bzp4P6DC5c1gEMRXH3KX
iBbVDISWpL2/jpxxyLEe5sVSukBNWnTaSbHAjWUc/ghbKrscq/DvIyhEwUFKnII9R5FEKFKscf9t
laWcmbrbIewq5wbz8Zn/kZ5AhNjEEhPkzPFa96DnFStXtCb+YdVfRLQRBDdNa63aV0eUzUFum7Be
XRncFP36yhoD0KEnZ8rZeKZfAx+5sGMQDwejIlkjPtWePWL90GjmERRiwgSPBK6ISvOUvz/Liljg
zEyUNEZMspHuGb8/Gdt0Gj/dHC+MYiuu30pEzZVuCrWGItklt6ZAMLnBdHW+wVt9uxvCxIJa/VZi
xc5sxsymgQGThdmFYVd+OR0Z3gvZ7X/PPas7OHeXbtzd9MnejetfTIZgN2WgcWoNF+YAuZENe6Uh
PN2mVA3dURmfBLH7gYe1qO8UgY466djN1uziGAZ5hZHtoUC/rpfM7897jjwvFa/SJ5mv0NhfbKsC
UgNZYi/AfovjlBa7RL1aMBZWqNVcApNf81z4P7s6X32oslpWe5Z5fKYS7Xi/+ChymU6/AouFzYNM
MdqTvecqoLuLiydv67KLU4+2MARuAjnVahtucZmEAUvUESZqSBGr2H01u3Z/ZDz0Ls73Ie6XBgul
BuPP88jchMMGC0bVTPVfHzyPCseYc+quT5HrD1duunuNPFbUaSN5JHuA2xRsK982bk2Hg/wKg6rJ
FKvRhZpRucWweOpqW+H5nEdOr8MKNWyZrgyToAMTr206r4hdtjI+SuUxLxacOD01c6pwZVF2wdG9
kGMUJXgwZNyGF8c40SgZGD7xCtA5sYtno7i2ciWIBukDFqVggzuheNurkU/G6KkU8cleM7ARg82P
OdUB4R2h0OYmuep46XacMgeP5Dqu+CnTxawecVab1jUu7+ftDr4ZKWtEtuoa0P2uwFXOIVm5cTsk
NmIHYi767NDrKnmu7/zJqqa3qcLYTMkfdUmxovQO8CcjWgp4TNDICFsxHBDxkm+tgALXALCiM+78
Q5/dQwcNI/Sn6e//IV0hMISeMDBAYOZ99dpfB0kZKT7JNOO64MyZMmKvm6slxeEcuU8dRMUWrxui
TAVtjFzKs20dc8DBdXbWadkqAU14eKRbNGI8YV+HUFlblcHj8OANZCfMXWmWvWVZMPFQAQtwHnXm
pMeBG9vf/5AteKkj99vAU0ydCZUDxMPR5ApwNWOMfkk9O4LVZ4RzBE8cJsPPTsUHNWrhHmuuZ1/J
rpNW6Knmgok7IfeKlDCRmN9T8YGts+0nVmlw2EcwRdk2B6VC31BLTHqhnV8xu/dMLveqGPrb1o6W
ZjuOe0X4Ld0kXbh6jDgKwKk8DkWcCJ4MiBEpPdALB6cD2AWRTxU2cog0BP2u74caddckuYlbE5+9
WOs7KJKt/8dBj28VjPOLiT5uGqp+PNNuEttG9lCiecUosGKqAFDZQFjl1MziAQ4iAM3TWw7Su/Vu
FvvXoKCLwobnBUCGvamWA2d+v+XWZmcGoWvgVcJb+77Yj2caekkzFY8hj/UwvCnT/7eZNIFaIEj4
4/BhH2HDd/vHiSFIuKVBzrBbIk0Pp0kbxNdupbvCVZRXQYa6v6v9UBdFtDZWbFHxXEgSHXnCnJtm
W8lebCmmmYS6pAJ57ERernJU1WcSgFNwLdZXqvPPhwgjEXT6YUPACjT1W7HiTJZzcCzJm/tz9ZE3
kk9B/1SpuTwU/2qeu+Y06PAGe9Mf5plNUHeLlyIDMavsdbfaIwMPaUnv5ITFhdZzWX7IphrQly/t
iBV2LOkapxlATCgISOJkybMpBq7kGGEAAFXmW5e/CcFebdklJE/Z9YTHPDudbuxaPQZk/+F1UEjb
Xkf6a/6ZeeLgXer8qh64Jbtt+DshxDu1NO/XFijj9fsjCHW0R5zOpI3fV10aPYnaQZLBKqRbLnrC
+DMpqTWyESO2VfNBX5cW+PpOEZgNA16nAzOn/E9mv4rmktTzXW+Kon0oJlTmoJbhrZhhNRtD/ab4
mrOb5KSEu18NHLNMDk9kFoqt9hG5KwzWbkhy1vJUKSyJrRiVWr901JrgDvzOM77YFxC5znnxNCwa
LtPRBjV5hto45KxwSKKHP9mEfWbEQHpUmkHqKym16qyIdwI81LbE2xYi9CqdsqsGUD0BCFdMXEGw
EaSUzchwR/Zpf2Mesb7nqJXzDpVBESaRSocO0hObCvFwCknWPkUqSLo7tBCwi/dorVPCWeM0QmYF
8QaB2TMhsP+Ah8tYvlmgCmM2gBKmwJuyg+zDT7H35orn2gOkxCelAXwX2V7YExDlYT4dZAocIGyD
LIpzBKVcs6pajyHXzmJz35Zn3sm/Rd/X6/eCX5wG6WMe8c0CJDOJIv8jNuJ+D+h08tEOiYVDf+TQ
FboXQm/TN5HByuIEssKlx2ZVxGMNmb4N8MZpNOUNJDOliNh2mFNandA91NzLRNE46pvkQWJJbVF1
lOQcUpwrO6NaSZRzkPv/JHG8AHwTaxOTF4HWiQHmIU9Z08eNIE7VIzf2vjlfgxlr50cbhpGHxA0G
3mSt3e3c0DY5V2HAU3ODtwa2RUwYFGBNN51Pp1Y7AghHuU/YEhnrxzLLNwUXdkQkAQKXpwQBg/3d
gia21ni3cvsSE7dpFAwZ2Z+H7Twmntg9tPyBzZey2lyy5oVByKKMymA5JDyJfioRiw2edueDVIeY
L2P5IMFT03BS/RbyZpC0RMGbuBe1XP8qynwAFQDZ6AV6ANDUb92zjAsQKPx3ufC2qJiMIu9/BfA7
la06yOmAwaZpwf3ag5nFjt4zAJPIWJquhQkyXuLFwMuTX7jC/wmaOhxZ8Xy+vxu8/Mib48gBY0so
0rCHa/k3dk6VvuY7EaEPJCyajbkcOO1AFDZHMfGZWQeBmikCsymv69M4RRxqPjgBbEBLyJQ94TE+
T5/TH0sPeCoJ0tdLDN9snjeKwmIqsqHHmq5j688KAPa1uLJHzPd6OjPqS7hQwqSxhxRyQtdJXgXL
rUR6ZVsNfjx+umkFyzdqzRtXbP8xEAbl0Fy9W2F9BM2KHsRqIxUEI5aySVEfLWnaxmwZfnOAC/ik
yxe0gpg0uyMxkMqrPX4DaM24RH7rQ2/+kNOs1NKFXE3RNM6+aNhFQWrPds1dzi4M39mRnFVZPyv3
GBWfqE1HtAFyGkecEM1QY1TD5M3q5EwuP6q1AnVRWfeO/l87OHsNls+k7MZ4meP01XNlH9I43v89
B7UmEMR7shl1JHFzH+LjgLYimpXcT3V0TIF8FTk0IFLULL8x6hEfWlbj3Y9YUN0LgtqAFluAZzNG
rHQlc/wrVRaR+04zYrmOOAf7uCDr2OCloPBUdrq0lESXZr9Bykxz3RE2N77FcmWmP1RGCM6mv50e
anS7G7fW3jrw72m7ilwvSay5njt+HeDulOXaHqRMoLHtrSauXRNIVCa4c/Gk8SLtu+HhmXapQUwS
GfudbHktRTP9Tn0s3x5pPtHCUOBWn9g7XBu1tTdQHeXorYmxKO2FJvyRm330odFDbgsAyiLqqZ4W
s2zzsPXnxuZOCS6/SJpur2FCBcsKk5FKkmK6RqxisRcxZMBa8J7cwHyOBmDcdEwFn1Fl1crWg4kx
elQgPOBkkTnfd9Jb8npu9dnDyQ3sqCSDiiu6F7lLacbwo2/uZWngZf7U3RUhfyDrMCOTUDKuXucl
yKVmdVk2Vh51PeVGJv4yJFoL+SkaUYz1PPq/EBzkBj9DHSdQe67nNkDNijbt62wCA+zz3loCdQL7
ury93uUpEnorwbCi+ejR3y6ZYiopQa/8RvHD21mbLO8khWsGmtTKixP9WyXq/ROYpcQkPQk2vcWE
04atYlhYm7QTfBDwjSVFi5eGSfrEcl64XT0Xz2M8HZsUIRTK+CzFPpjZ7YUFc3/UqPq5G+RG9Y7a
fd7ayn9aYpkcvLmh4tQgF87WmnVq7pVgjiIM622zi+5CtSGqL6BVCYndZVq56PGpQA+2zcN838NY
RH5K07+zisvWs6fhyjG35fzOq/EeIEGQ4ItbV8+oWJl4TL0wQP8N4erdKyLHNSTSoY/qX6iRHUJ1
CHFUt2V4kIJ80C4NAFm8xryZBB4NGrrwol2G4BaTdcHU17J6C29It/2M7RI/ot8yX5PaOMWtXtIs
WmcRtXmJqbDwp3VP1RBn2J6Xe6Cg3g7RWnd+jpEB3Rr4JYc6Q79CLZKMhoc8gXKBpdYZzISA23ou
thDHLag9031gfBzGti7Fg633ZDPrGoap8TAF8NV1rodtqu3T7h0+1wEc1pwfSx4SWIc9FjQK4hPP
hS9/od5p9/twY2DBWtHdjZt4SUYQcv5H1SP27/9fxGTVF6H1lT+nPOSyr0ZxA9s5AUaN6QpKYFR7
LjtXQ61S1SU7JhOy6S/9xZYsJpyWW7Mn22E/rt1z5eWCROm0PDeZ3QG04/7R1EAMQbf9ow+GEAKP
qKQjgIXvzZ+W9bftuQv5jgTOnWnSSEmUu0ho+C/ihwBLEcSGcS4OiEwDgQKmt3fPzNon2gdZAIE8
2Fu7AmfMzl5SqAvKJl2PSkPdpDOHMULcnJ9vac+CnD7JeKUIpCpahduT7M7aUKbcn78w7+N7jo0W
HTN/S/v0ZiWSeTe/GS3wQedx00hGFvQKLo9H92bXvmfMvMuepIiPVpjDeKJxow4HQMAPMRk94aOJ
ffMBYD5IkuO8Dgxw73ywLjKQa1Xhksfh+B0uMGsI45snwV8EXgvwLMGMDQpsi/wdiu/kPzb7CggI
XOVATdyWoVkpxvaC7Rdj1M7atTOI7ByXsytsg+JKisodjt0t1muFo62/yYPBxNlIvSCu2wQ+mThv
A4rwfsve8vho+GqMx1LyJtgx+LiPve7xdEHQa8wP0Epgnz2MEPJkt44QcqBci42Y67wfQe/fW60r
0qL8AuRWZk2c9VZ6HJbIIagCjEaU8gvdSDUXy9juJcbOcF8cUlNBjeIdYqywmu5LpYsGmjtTjp0E
94ArQJGpMBSfa6Xz47Wivc+aVr7uhBYmfB2De+o2xViqxhSYk0Dq9weK62Tr8rBSLnHH/ZUzoizQ
O17Inp3jn3dGipcgT2epj54VC1EMVQBgL9WKogwAnejQDolQE698zUVx1f4+mH3sLDJEmw50RR41
FqYb0u/1jfvLmufBZAfxAfbiXwDjZIp4DSJcHwIYr2bwJuR2WgCoKNQWd6esazeM6Bcu+18mdk6R
Xsgnfu5lQUKWet48qEGm5o8fvAV8sNIUTQ1nhREcbloqQGAgsbP4A7OCJVBnmKPYr8FI8QhzEwsn
OBqbNx4A9TwxAPznAv2Vgh3R6QGA0VeWhASu90VippZ6cqhnfT2j3aGJLU+oLtXjAIbsyU77+A51
XC+64IZlST7Lj3wYM/pbMsC7LK0JxU69R6fqZB2EVvC2+mTl9i0zSy8+x7Nb9wttiTr7acx7Xel7
bodKI1HYhClymEhdgEY04WL+TTp/E6N7erp+e/iZofNBqA4rYM/ix1c1pQQzivK6XG/HZxKkUMFx
nmoVo801Si1BIJc08jsb8g3rPrNPfSeC9R6mbz649+Zlv5vjrvLdzBtBTzeL3QraFD68C8noiGI4
zk6UC/My6UR5b7+1pn5ObTFIO4GEYgEA/YXLMjb+THRY55wAWb/mkQugNVUWKtjvXtbtadLI8b7G
Iwagvf7jQysm54F3I1oap0xdzXHt/yIZw8xteJ1Vntnmml+isgPmP36vf8IZ5rg8Ihmpdom9QVyY
iTHQ618FAQ+bpSh9QNeS0aO6L9F3RkCrhROSvR6LN6Sr3eg+AS8VwTtyyU2esoTGiTRbBQ6213zz
fHNyNZ9W+gGMZ83xLTbNM4CcnWfi+FyTnT3pz21XYhpXPIeD34XX7lS23WaeXvATSU6znBhofQn+
wzEAegneR20uLVV+8W5ah0Fa6OgwEQGxKNaj/haWKK5oozE4roMeaE9ClHY2JDPQ9gOpJnAOWfxI
LJdP4IWmyTYdSv1FwBGo+5OCfrF+XDXuLtpmY3IHxJ1+/+0pG4sZYt4DhMO5KZVaGrTqxjSy4+9p
Orm/S8mB2JFotaHh46MaUCdiVHSlZn29b4l4tPtb463E8gEVjsSGQ6ZPM2NtjRQADDxs7cCFmXdH
tuniP/I3eFYuO46PYWsNg8KErcalqxdfBp9tjAVcynBqBHimgw6EAZVMI1dJD0LN26N5Imkdej5W
voUtK5761JWGO4ODXmq0R9Llf6ltflMUZ492mhe68SThCwnSlzkGJPx3Y+ShvupKLd7k/B0EArvq
wpE7BWT1MlZ4vZpYWwG2OvzVuTI00PHxNC7c0SJPmD5N9j6Pe0ErI8gArb1Pcs9Pox4fK1bp/Zeb
tIOnBQzRSxLYQf6lUheH3jSQGIvKSufiyAo1mqyC5sssOtdCHcMGl8LVLCx8CiY7Sw63c6wRnU70
kEildMYG5Wt8v6Yld0BB5fTmG3cSK2okVcqKbRJWbcaEBqzDZgIoC6el6qHvOl4v/APVbf0oPfrp
h0PkOvD9nNnKZ3uqi139sdYwfh4JZKcOqqRWE+5W1VyLXzJKQlhBiqKD8B2iOy/tovYWBySwRYhb
HIYAQF12p60VEhti0eZex0UjR/cUpPdaWIi+qOGihgfYACNYWj91uH+9t2+h1nfsla+1KEZ5mXuw
7u6fGnPBpG3pQ4deGAYHsHkhNaWIp/P22nDVf6oCgBV1Z2LuLnwvl2wWFl/gIwA5VQef8KCyDqP/
iSxkhYNNckE5qK10nUFg/FJwln7lUnf1pRZvQqie7BypmRD99TAguKNmfxCJ8MaEs+KRgp5ozpKF
MEMNmT+4fbzIHOlRfV94TsiGqb1Nn9G9/nBQv7ZjnoMC76imXSpE/bLJtjDphAY8RwrkcJ6UIpif
NMh+W4koc/PzosAFB3OC5bFbTiktDY4QDAODfMstFQQ0I7qmX8h3sC7P6xunu1jJM9xOTMkir9M4
08oeCGeezwA2V8RJq1eQlIiYVv0jaZDZNL+Vzw/0o1tXFnm99BnH9oeS/PMrxdNEU9L7FwqK6OP4
4gg58Gjdz325NM/kYKXHJEKphJwUYVwS44xJUUZX79cxFpShmWkQdtzvRb3fmHE6u6yjSYxwGsZF
GZJbfaGaiTrrJ7sWIcoZxRd6C0d9m5MsN9c8X+DNqAbt3MXxpLhkYwFpsd5t96I04Y7vEoWqbLTV
i37ZZuvQpLnm9dGgkNwg2uBevXFn5+z7EyuVlob5pvZMzY5gXo3Zgo+/mTe7cHPS3b2rqruuWt0G
IfaDdjP1/yfbcq2dVbt3emRAXN8sV6bLd6Xpu8Rb+2edZPk6Fav0oqbsTKaZyiRCu3miHJ1P4oD0
6lSpCIhuTWRywPD4j5xcefe62S3c+s+S3LBPph/dM8oLfzZpjBsfA3MyEN2M3UUwDHOmREEptpG7
dQlT2daYDTFe7s1fE79bsDSK6n6h9U4sK6WcRzxb3ULO1MZLLtdj2amifAFJ46QQMzuwN3eQoVT/
H+4hHMYTH+45eH4P4CFprLiruA6OqPYpPQn4wUJ6NHjjvl3XnaB4xiuPMYtmtBr+ZihSe4vhJrU0
PGBx2kCaFIiQbU6Pe8CBb2/TKyHtVMd/NpC/X3mNt3jW5L2yMLBc6QBcEteWtP50skic7mnwxs0Y
VtqhS1YsE9mQ5WnT5U1XYaOyjGZ4d3Az1aqGXB/JGf1xI0fPrMZ5jw7a+Y5swr2urK6lSuVAH+HI
AFUpC5T6E6r6fAIyRIJ4Jo7qGFW1H/BTVTZ9lcUPF6qlmDvlWb0OT3B5cIQkQORV9zi8sc+XqZs6
slqeZYYmyHDiiWAu0M+AJGhpfSbhXWZa7Z6KXdnrny4dyOHeeOzF/ZUkD+bOA1W6ZGj7HMzOsDAc
FBENeZKRHOJLm4/E2MdhD7XCcTZ/pPFN/Rf+tY8IzZ8TjXqFSyYaK4qBqoL53r7SSbG+3WQ1llhv
CUCE/o6gDzsKL71jzh6FJYYf6raDZoLz2Gureiq3lHC7VewgUPBti2Es3FmtHwUGEjMiGLxlvdhd
IlDVslRAK0ok6PsgioaSPIC345VRKPZS9OBshtSLrLaEf8iuNc+XAt3mFFEqRPJjE4JpLVCU0f5v
ElO9ig1NhkqqQYrcLM4xN3ENHd8zEIqftA4Ti09+3NVpDhaKxsz0Z4cwgASguGGXGx+Oymc9Esou
pb2LAp1MgxonB6UnscXUUoZi7b7tImrBfKHfsE3WUbnvensJHrpXdw6wviosxrieQNGWn+nbZX+v
yPJHoG5oop/PyxvVza5orH5GNO/3S0dX0TawLvyDAp7Aa7sBSakruRyrgFOA2/dJD9DAzKPjiPcH
HU4M7A4N3XrZ6XAKw3ZoRBCfFIeH9mIWUn2SkXW22ruedF6NRxMVF5JxYPS4SCtFDE5fpOVL7k1r
WbUSbCtGbrKcgjPA//cMaSRHj3Y9g2XjjB0PfPx3Ni/4iY+fI+xVirCKMKfxIXu9H43OXC44LzA4
x7wmlkKeogZ41KyiqET07ScEu2OeBj63zmeguvrz3QSvUSECwCKZHM1FMx055lzlpanK3nP4b/zm
k0yjhVJCogYanPllwxMYeFq6vqGMOqwM/hjtNhhrUImFG1Zax/CkOoroRIq94/Vg6Aew1d6ihPfr
cT5cljnDIUFBCdylU/MB6qqpn06sQIERIpCYribokFeta1xVD+0JgHREDK8WEkf/90UPeYiv/Hwo
c/+Sn/+GIWG+YAYca2Q6Ga4clmDrzebKSrm4JqWK+1cHQeoyC7QRmASutsgMJMounksJ12at0QJZ
llivzRRlEYZVQknpuvuZhniSnFqvgtMWuUXxW2/J7om8oIyJLo7VzGPlmuzwsgwbB4A0jPARAQXl
+l+eFnpVK5UcYuSBkkAPdV9bKDx9Jfa4UQxRSlIIGBN91OPv4AmLXIORtU+61YGvzP6VhIdpBCbm
QsgCek8q9QqMMIplNaklAUK+OCeH7NrsePFtgAhWCjN33BTjpIxwVxiqsect9yp1Scr8BFsHg7pi
R6NDex8enmOiRoQW1Oca6hn4qThFi5pyjxg8RjPEoaGmUmpW6pgLnGM1L4BRhBVdNiLINbiSam9k
MvlrZn9zpLbYXK66TRTNze2EKXv48P5bxzk2VloeI1iCsdzTMSBYmN2/qXAuq1YwFSqF2G+LwEEE
EVrrOdMAEuC0MAtmzAZ5owu2OqBy0XWbtzi8NqH8tiOQGfak1O/79B90l8YQdFl0glYZ3/4I3/t2
oTATXR2+pkndLyez0wAxzRe0Lmq55q0MKjH1rMd2SJeScA1J/Ze7esgdISvhG9gOL4ST4rCOVkDE
YmE+jQ/1ixYBFRPBKTpC/kEXsoKt2WZULQUetyLWTNz9VuZPq9nSXA3gJaO8/7WPlMT4qsR6e6SR
uQDIkAkYD1ZneIGYXTapoUrrZhOuvNK0CaYuI2ZaYmYJ70A2uUBuzxZQlI7HnGQ9LDLsAriMNzyG
NMIF7AFToB+GQ0i0FbSITvvWZu3d+bMv8PwDJ3CPFoKdT7wSBItZc72oQK3sq6ck0OUQu72ok4nW
XDb2k2+Xovwrc1khUso2dKvEH1I2GgI5mwmFjQAJg760krcN/dzUPPWQCek+ciuBc1uaf9TsClr/
ReahAVc7/cGAQuHzXlABZp/P0TJ4ow4l3Lrn6yeZMt1mkEtIr7x7NFyhpeEwP/8dTH9llRvJCBuo
W1gpuD7QFh0lPTicc5amir7kMitNQqYCp/ncYRiDd9FPyzs1WLsEHZ63QCai9kJ5WrcDDayssuTT
OzIBo+SMgr+ptqmC1hPG1twnr1f82r2sofd0yL1L6KxBwbULhRUQz+GKZ5mXczMtFP3fkNVSfxZ9
KYNKIQ3x5IoTia+fuVqoxhnvXWjrXYtmX4CoGqFS+Z46vNETqE6jRaXAIZ6woD3ik68/tBLGYFiO
wC1IB7BYmh7QtxV3wv67bSBVDvySSXUwaPV1gbmHzD3wgXRVHZz0Z+1NGJzAN7Li6R41b91XDPZQ
AlX8/CxDnj+jyonErSY9jkYIX+JkiLEmJGBmu1FAgaEbcYuB2dU2pHbMdGiTOveyXtMcQo+J8SHy
/xRl/yf5UuP8lCOtW5Wd5diC5KmK6dv7hMyIwCKf6JJIrwq5793lK6i407d/zXwIPk3up/oV9AH8
3M21we36tHO+A9UPrZDWhEjh7pCeLSm2KMp9lC4TaFrMQyhJKGbpY5+/24su19CjwbzxEI2nZtGE
xz/Pi5z/RPB1bUN4k5mV1zqev/eBBPO9FTR8/y1ePYGGyhDuufFkfWygcT9Q/vIqLFvwMjPqOvxj
Y336HhzVSwNhbR3uNZNaV+FXNHNobbSs/8Qon2F5YYGbP0nDuOR9rPRrC2cl0qN5A21CUxO5cGeN
YQ8Iyic4A5AEFR/FT6LWqxeomUgEgoHSRNhOf6LxSifA7TNjW+5Jfbqo7tjF6GIrTUKfbF3noY36
cwGKqVz+LAFAJWk+EkANDhueYk4pokv/2tpkg/3IP9ZIz3Dx4+10+POuOXLMs6amIdppty50taev
BcfMInwVvvZL7gBgYPuD+uvmqk/6qB1OduqdRgAgI5O9UpDkd8HHr/zrgehT/xRqaGLwJp5wTpxj
Rlwr/JbaZVbRByPyGr7sEKKejYyMCpfGuL8UV80eq5YQDEfqYbRFQRGjHY/+90RQTEaC8xL+zShv
mqAacWeAKpxMNgWDgZ1dQWVDV3+ilLWWeUtv39IlFY4bNMyyBwm7NrW2mDZIcQik1hvhrVQdNBXd
jGeabI+vy52hW1gjuB0dS0WhwNimf2rKkoOeRyOiwrjTKl5Q2wMOu8tu295YiR8nPyXdxi7+FBF2
QNTV1RRwTjeV7BmHNwRPYJfLNhFe3mmGvPu+6RsBtZXkfpngsJV8vQuu7NM2KhQ/nCnCKxD4vd73
ir1cHHvN+lJjpVHIcgFZp8At9eZOvjRcdruSZ8T1P3gIX5F1VnASQGuMRJl7BuTbjxyVE9/OqGbe
HjS5EVc8KI359l9weVynln9/uSQnK/kiSowU3dll25o9Ma+WEIp18ey0Gw5hdBW37zqXYt1wyquW
vUg3GUvImB8vD+eOUgnzCtMXqJubfoyEx4sCY0XM5mx6zLUEii3RaereiHRa08G6GZcmvJ74OnYy
Ctj1os2ikhFQRITaMKL7zp18P/v3OtkgGy3cxXd8vCv9n6s1Jd+V+GgqIPyjJ/UoRd9+yZpPJSMk
GU5yj07Yrk9yKHuEf6574mBA0Fp9DhwjmlEyIa/OvIinYFFKa67+PhGu/+DGAoJYrf8Zx4KpBBAB
PBjFJHppSjXd8lqaKZ7cDGZmgyYe4WveBiESKZNLE0nbtdQHZOJcZQXziu+5HqT4QJ6yof6e6n5N
zPuctegTfbTJDEVgoTOUTrP1v7NmavcKMIJL7RB5lBp36mMUDCPbaCGkL8YgoqFm+CYGzBG27wjb
hQOuceccqjxqup03abv5bdMgx4oT3JPSior4uaUWimvNSyncxoRwtmALKGBFM0k3zhE6R45UO+fw
aNAd+wQvM29wqihX/qzaPJfjVEuR9f5sK7UkgctZYMhhVsm4l+jYo0waNyNR6C7qXeFgxAFpsN8w
Q5XtRCTj3IDY4xCQuP1wZxytrq5nwvGjtLH7xb3+LzY/jQ9g1MAIYMgIRtzB3FRs17+Y0oXt2yzw
bKMWC9w/P/dTKkx4HEI4MIr3y7rkQRon5of9EIlJmz6QMDyzIc01yVWC9eyAzOybAVtZKzp+Yt/q
2AUr9jYg1TEZ0OpEpyr0RrTVbqy7NebD1UtpzBH/rLw2eHeMWC6KFrLkRpk3k/alFs5eOCvfs6PN
zflAjMAZ5tES6bGs4DjVykf3li20tCb9/LtBfllKUJpf2ZZDhBjj8rrdn6JAfQQeAzfMF9wxrG5U
quHuj6g6y3ciImQtCWW0jVn0HToAW4OQI2JbUbJcf7OriECfgbsdr2TK+RkDGN8FZjooeULNAHST
nTUQzIyC9o62AqDocYb10lt4RMPs/b3lGEVnN7ewu0oSix0YJyEpgJ1FIW5o4/Zm+rWXzEIkUDLo
siMKZdmAvMx3fpKNHp3epqFrFAm9ytxe4g6ZQXt9T4AA52BXfP3TxlX5zDLu4D37GOpcf/rzNNKb
LyxTPRPN6+GJiiaBgxsMniDmp13xXvb1JziAxcjBSE0Me0ARKbx33jNJxgvCF4ftY6OlmgzakvJw
Psj9FeKFW15vQphxxaMUEawSoi4vpZUxfnXLI9EnhDK29wXARVC4VdxL61J3wPSCuTWsnP3Jec55
ZhCpWMt9lB3zBfGHK4Xk4K6B0ZRAdXqMGWQgTjZDgW9S/z76TONBBOXBdGFeTUt4MJkpgT26f4gi
ZNhgxfDvbBi/egmngpm7z9NytiIKVXajE9vsv5oRwaYCBwNMyP2TjGqvmdp0f4iuCS8I1R11AgTd
dFMnWmfHpoHH1PcGfE8xi9sPE5BiJKCOqMuD+ZY/MuwCSogKroFi8hq6B2s8opEv3DvDJUKx41DB
ywU3XoBeN16C/0Lndg4tYWc4xeZmEfkNZUMHq6havrm+hSIK3eEqVOEDyW5oHYEwPSQOPtH6eS0o
DxGIqLmQ3c4uZW7E/41G9Y0sOHTYCf1b7X96M0iO1Wted/+6ID1IGCyYZfnFnhHPdr/P9fvgJVFw
lC41m2Rf4fUHHdkmYMbOPsbB0q2Y5HblO0C4heTmGbN0QK27CAiUlGQkYBZyXU1YCGzMs275o2Mn
VF416vVs3P9t288zD/S1B2DLbH+FxeTy7ZZ8wi1qTROeldH8tBln00UMJ8Z2Al44kBLwdkBTugT/
d9CcQ0KwpI/TwLrR6bx8048FQXkgM+R6OhAFYKsZ6FELQfqt4etpeNP8x8MIJPykeZIBRlsELv2V
l1ocA8Km78fSco+dgm10/u9bZsGfwjFd/jHsLXwBiET4NZj+qjZqcKJdimyAdCvbqvJNgepA8mx6
bZdihs9g8LgEbjT55P85QE98pBr8cNBT6fh9k4V9fiWiu3IjbY/GwbGvGKd4i7kpr+70oAWMHTkx
/gBAw1mI9r/LTTJrCqCUOWTMQJ1vdEM0w7QOId2jt8Sc1zTPbjcTNy68//0jnhDYfDQeT3tYGVhB
9XY4WAcn/Vk2MxkwYrMVh1KK93neFJivwZ3MwRqehxLkxwpXp7srCnnqeHcknkdQ9pOFUyHGYY1Q
lNdZVlHJibF5aU+QTNAUHVHYAD0yJJcvAYp3AVHKf1yO6HZDZeZIpMAz17iH9vGSy991Q9/uaPnJ
Eqh8d3qOP/n+6FzFr81RrTRw0NHkFnKyHvcsyMe9FDfoiK+WUadiQJb1xNb4w6JBJ1FymZBwvVC1
HG5EeXPXn5ILWqGKY7b4RrwaYumbKyCAEHhzu1OIN+dWuMjiraAlemSAlsijbwWrWaUlfCp8qXK0
uUF9GA0V5VCeu2PrpUhlsi/HcIshPOJreRJbBdS0kPexr4eLeY1OZ87Xslld3ZXIbRMUwEf/8v6l
+0lE1RYsKiau/zT2ctICHmlooattR/SJ6XJK+ImiFADYYKo0vGvMTo6oiTDaKCnJQ7YM70iWOTzF
oyR03z5Hv4kfnEZALV2Z4/Fl22X8jKOV4snK1p9+RYfkdvP4FfDGoNRohu30WMphb0iz9U2zp0HO
wos3zWKHv0Y2EtE452CS/Uo4lf8jUiMdILdrq+wEF2zNdCbGvQVG1M/Iv2temg4Oza0uw9jCIJmr
PeJxR/IvtDYTITtU6Ntsxem2KhG3c8FZK1YRe6W8Xf81NdK0iZnT1E+x4VI/diTBEHlCsDSYwUiU
cNLKKM5lhxySjuV5rFDydcOzJZ+gJB1YmzCwLdopSMriw1AMYINiJWdJxCq20A0anlLZShT2NPz8
LkAYIRbTa4hzvCeqdLzKrOb9F+8zM5mzrQe8kYqGb74FfdeYmQ78RSa4lT2Ialy5vj6zLmkKYuv2
vzxbRPaGxHSGhERqrgU8RW5hJ8+kPlKowhjt3XdcmM9TqT4krZ0SZoMyGHoI/CQexFBUOrJ4aFeK
mn2Hl8OjRX01bOyGe9kYpjYbFP+aqiTGa3J2ZIYrOncGFnNZkzf8ofXFLLWqSF5NrzBX5+gJh61U
tuKTzpteJC8S6ymh0sEQ8d6mEw03rOILYNZZFEzy/IEC4l6N6ybikqYz/bPvVxOY68IEHCvlnxGR
CuW/hDth7VVne481Sfrg2aJC2vGdipZ3ow7kRW9bZaFO/1soAb4Y8Gr3evyMtUlavqvo4fQHLPbd
BMmW+HOW4apDfjgvcqwStvua19TF8otOQ2olTVIrGyo4ryfFzZ95OZ5XQLVFv44AUMLa9pW37643
WYuum+UZogZUQ4bt17dZ2Hy8wofKaC7jl3PktaGWRUXAjn/1bs7VQ0sKd/icabnrt/d6LL5oJRvj
peXghRJRo2u+k/jYv86BgPkM9YQbmTRe7nk5qKKaT4C4Z2KgIZPJ0muD6LLZDKAa74zOlqTa+zfw
aAFyUghfTLwA3B9O09Vl/F8IoxOviK4/po4AfesIvuAdeQ5WwNFyB565fRTFYgBxYoeDKIpcAkpZ
T1TywAOJ9m9LnkLsyiBDAsGTm0MIKRvRLDPBk8QH2cjTgjlcabxr8Dw+N94lJ5EV8D7LJEiLnDkZ
xZQQqP3YHBAKQcCpsKvTgavwvT6RwKOe+eGBckIkd6FVPZKkzuxOjvvk3lOFsMzFaq7sSCa5aRQZ
WBRnJKgoDzBzNhzl97iPcmXwyyc0KF+D4beBQWw2b5G1AUILYcFaDxJmnV20AQ5X+o3dHoPAGHLc
EimzQ52S6JQ7dnPGdmaYTeWrYY5XcfxHjqf8sx1XOlC6FOx918/cPbQ/zkbFVbAZpy9wuqugr6wJ
2en2wyh60+z7x7KCbXFTLFgBkARGKGob5Iu3ds2dtFgniEh1CboDlizKD+FcEsenjuoLICWlGv43
PjJT9Rz1WqWaY0Yh4HlHwirasoWM6yXHkmrmvNphokRAXxhRT49PW3UWdQKwN6rwLWBv/D2PcJYW
MAv1UWDBIDVESbljnGA0QusX/DlHw19ythseDRrIoSMKsQ8SSVJ2XqXT/et7ukdOkW5b6vOeYFGg
2OOvQHfOdXhWDqaqO8Pf0coYj+85tieDVxc2wbplxXn9W8HidOpUMN3UAjeSvPYLIg2xHYp6vrG4
oS6okYrp36T/T7qFCzjqXmIcexiphn1i05pSQx+xZ0Lgp0L3VQmpPcgkHi8F5/TxbQTLZ/jbfP+n
irXEnCjKL0Gq71zJozHbXPzM9HGvQgKKs5rfgi4NUd/eqsnpAi6Hi4sjg+N7QwqvZ7EgyVOOpLFC
AEZGhd4LXwpf3ogoycd46kg996E6jwYQzy3K+CLnXyVdRCFXvg7C2GdD2p25FLL5Ndodwphu3EMp
RHgx4o2GjgXgCbBQDlTbBPtEQojsSiVIsqYwGwu8BcAG/2P439bvs4vNk3zbSKEiPUk10DLa6y8g
yTlCcfCFJEX/xvjDXbwX5WkQBIIK4L9uD/VG80LO9wBxExtI31BGg75gKthbl6vQH70tBvpgyVuC
RFehEpXoe7xzX8h7CRMIJvII5yIj5WlwiRTf0sp8XpvA5KVDFFNQKFXDku/RoR7YJylGpgeTGqJE
J/xlb/KL5wWubbKXf31Hpvxuy07JdzikVoHecZfM2gd69v3hmjIZGIilBKj32Tq71mA7DPifVkPx
SFc6YjaCKsofs8ayC3T83DrpFBzhNYFZVvKapQgah3eu3VpnqKyOUyNH/tjkYCJbCnz8YBmTiiZy
VQVi4U1siPu3IU13Hs1nFdeZePmgy3vzTLbk/qMgNUZUyAW6Dj4XEQGXDhJky4MgKnIgoAi4xIxT
O8AQvto5wA8ejY5Lb41JNsDtAJKNdE0RKBoNB6NEiT59HjsoQq8H8gHXXDHcdO90ObhkXwVojUpJ
IBjS6A+W5P/rdUhW3sRKctlORTphfSpCLeX+WrthkmBwrxCRBIsFrxdNO25j5HCMADkFXiVQIveV
2WvlqWjaCCSAH0Ek+He6NNPy/Lf/3LVIKd5EC3TfCwO/Uyi7jyzRjrZeQpY+Nx6gtUzMEIIllxwC
ar+HkZvQLu2UqC8XmkMFL/FdtaL4BipHCYCwe6OgQs97Iup9dGAllL3KUzfWSh4xEELNC4UW/lgP
LBw3gjTgusto67hVAT34C4C3EVW7DcEKHq/NxawDpcMqpzgQVF4S2uWG8OcuCsSNDlRYi01J8Adh
hbpSbCQAfjrffvmnEaPfSX3h37WUkLgzqDDjGg/wFdxNbsjbfEPk/mL3BUH97RFcYYW2bgefiLtA
2rM2CzgyEo25HO2vZlt5BhjRjjhDKnEFcFY0dSrwWUzeMSstjEDTxzF9Jd8pD9Zf26LyRTLtoIVj
9jktq21s2OV5+LgBjtqYpNk0bg2sE0WrC7tnOkt0i02jaYAXBNLDBBdUsEueOmA/mKtswDJhr3yc
b9RKDAXxnMqPQTMH+G98epLhtgnj7VmsrDrY4ovF6jtcIIS//CIRaCNB8XCjuzTO8cS2Vs9iMVvF
j/zbo4U5ZT8a0OrPZKAUQQvxjt85MFiwUmjotcgVS4zU4M/Uu58qSwIHuVBnzhSjvIs7CVc0MEeR
bGUtwpHlOMwmF0Mrdgc7EMjkPv42/K+dAIt5noFYX5oqoYy+Zaj2DuqR9JFP2sctefnfWxi9wDcT
eQvVzIvqZwt2Z6so2Fkxmx+PB5FAdpmZpMQ3rnoUDHSjsmO3AKIc2PAypQ5Ypji7/qFw0hF4Ee2X
Wo4Xl/5krKDfeEEtwadc71pLW9jBJAbeSwhrCI7GiB9XhKIzHcQCs2dUo8LHqBOhH4jv8LbmaTYV
BIZlrWDQr2FZ0vFcGzipu4WvHStV23sDa2OezJqioyxZaeQK5ciDzu6Bn3Alu5jdXjZ02tv41CzB
KO+YthmtDWb0Sh1Bj1bNs+iPQgeIddPJ3zR6EKQ3psH3QmIeCGahwnzOiliLtPcRRfpjnX9lN9z1
w7UjOL1ZBAeDG82MP/kP2IphDcOJSNTEC772WrYdpPf1eEuzijcG7f6HzwRggoPkJjAqtIV7Cb+y
bmrIjNYMe6PkSd0eddpl2Ta0NKAhPqQLioTU5FF/p1XM92QMUwvxoCMEK8FtrRCdNq3+pr1b/0eJ
T9yGUmMcDuKE6sil6Ct+5cDTGOcr/58sNJEdPsiWo44fZvHbIEzogQZRX4M1jdE7q13TiD2CqO2c
lRfGyhMYdKVycbFyKc4ZrcJZN1Ij/n3H2MytWNyL+A6xAnnwZCDLC75YKPYxivgwCgR4eZpP/y3U
/XBrxH+tSxd6tPjOMykzAmdobRIHAE1udz5l+53Mq8hazaSJ2+FYJYXmQMS1c/RSKl6+cRZsIN/h
d0vc3gLstjYnLxU66k2QDBAIDBBt/1ac1Ymm0w1U1Rk12IHUtJEvNhD0+OH+k3MVKA4oM/hIj66U
1auW2YIlKoxmHfYUsObr7vKNgRzu7+YXwQKGkdk0JBNBlv9yN0txZI1M6wzYwt4aAjGEDaLJudXH
+ADFumPWtRLFYFLd8Dlvh3tY9XESicX3H8bum0+n6dsKdGBm6shJSnK/a/xYtapDe2v83RYH6CL/
SQAQo3frNymdGNQRTJS34R9UsWYZIla5HNkf6Bq26o71Zh/cpYx4FL35iEjLmPquAySo0cLcmdDg
TMCYAtQ8gqXdTXqCBsonf8sXxd+0I29HeEps9KKqUpN1mXNeZitAyUhL3u8HrKB6LHl2P73q8DcD
bIcs3zHFJcZDnD+onyY6Hf5S64CTFlpdDMqStSY6j85IKwLHPJeeNIBkyrx4LQbmpaxJkaMHSBlb
swBIQS/dfbgyA0ZdLDHQKjTd9bouIKD/W2ZSko2zatOrjePhfgJUNcLyNt6cYcaafXVDEiI1iDCQ
k4bKYtAXrUDEt+vPuY2C+74Ul5BEVwDCgpd9uyze/uFkWh5EJI0f+U0nh9aPxjSEuf7kruAX8b+L
qju6TtrkhqNz+vuSUCoEjRdcoP5y/taawhyR1bLDYHSAzYQ1ZZj5YCO0yomChnBL2q054IbEmgOw
wJidfLJyD1pYpy5e4zci50AGh/kQXPVHQ0bCSCMt/0zhos/wkIEhr2ANl4kTd5FkoedjO/4j3fbh
jnGnUDsipTM6vXSr/JH//xacvf9tEUEnCctN72PZ26if+ZzRkUzjYGLwIE55geeg+PbN7AENqFzj
jp+aUzwV5ao47JId8dvgU0zQFa5h8ZVr+u5RbyV5TuQI2Ze5U9vK4KE9S05PFmUBvbOeB9Y94VYB
mrFPLwR0cxpDNC9s0bGuyp+nAmM5whGxsIXTMi8/znQg8EgO1HgCcG3NjKY++7FhfZzgT8tGKBz1
kJux1D/Nn+MgZFhGHxVk4XvAzuG0WW+KAGbzH7NPVcx7d16sgR6DmXDZFrawqlNuO/ry89ExeocA
O8XIdpW6kGHwCTeEsQILDTf4AzW81w8H6TJuYe97e//kG4g81lICFAh/iY7GoiNpCSY+zgLgq8IG
W5N987/PuGg62dOBYjj3i/3yCoZKyjHPyEipFpUF+jj1XBH4++OMEJva/6FVoJfGn92WQBo46Keo
fORe4yyhUN0A8EMyUQojlDj+R1X4SFUftPyZQ10WW4GybGlBWpjGjql8HNtEkb2Dtl3UBlkifldR
Mkm3I1jA6Oai0YeUXyMfIXMRNJyOJWNYZGy8vxFXUWEz5x4lgBmK48IvTmnfenMX59/YE9sVPKdH
zkNLy8/WSCRsQFU59K1TUCg6ZNxEkQcprIB9LKcCu4nujYWmaLActZtMXH7Bu7TAgUj6qs+FEtjy
JRnXgcHq0p31nVGuycsxgH7lShEGzbjMGcnaP18o+16ebUeQExkx2STeWCDGGsOy3pUvBciw/LXw
A3B0rGUW4bZk6+5a3ROWzzvWoC1iUIe9YyEzh2BR414qIG83TAxVdJ1fMCzxvMVZCIZLdytd6MIW
f7z2yFOpKfNGbyTWddl+/cTp/QT14bjGwTIg4TIOVCNA2/SoDKormZBpUcSHE1kmZYnH5HNOei9L
u7H5cJApQF6sz7eNqAWLoiqU3uPc8W0hssyQIJURifVJA7ngaXfB/83NqjFzCyVwDgfzBKLq/1nq
tnMmx8JmRJ/eJ2B3zUqnnSQuNJL1VwA2t0uVLIMd7nzK2z6xUDbqAT2OR9tyxZseaPCcyJN4Lugj
5hegewv5btEdx9xJddnfehLMUboe4CL+PcySjS7DFFMk9ex7RyaGMZvlTTQmmKzAiitbRtVlrMzq
021bRFVxovXzc7bBheT2YKbTcZF2o+51j5Pwm9sSq81h0paUFCixh9SFvy7Es9sY4EbA7gkLPTN1
N20/V4n8nM0Uc7qfatGAajJpaY6lYOExGrIgd1WxzpFnit1XnQPclFp4U/F1DuNDcyKRIJyAV7/i
QMHfeQLpTCW0XkAwwjruLHzVSv9poB3ya5gZ2vXmd7olyOYHByAPk7QaFiuNYNlx0TwiQzDA6sXr
6DCYVJDVRKgfJtIvxo0WG75yKWKbdKU9yHNT991tfIm/Xu5UWIFYbhWQfzGirRwnfTE8pfRdfCc6
S2sZFLfJUok1pVbNDvZUbvbkOTi1zs8mIc7LudNK1k1ZWpkMKHqI95TYUQG3w8YyWDK8n8Kr2EYB
oalNwiMYb+toIOj57bi5ZTu1FEX34sRzWEENRTmjjYXqJg+LojA8zioXB7tM+Oq/drDnLJgmWuRP
wyLDT7TRDprjPOFIADIO3I7IfLkfkKePq4L4WreNWvo4vKIQrU3gnj8brrEJCfswjTA3DJ8r7QTn
TpTiTzXO65S3Q6Mq5kOYHYYoowSCtca/BQnQoI9cRbOacApms6gCyEBvNia61vFoOnIOYWc9VFqu
3ELfWDUOyy2/cv6whaJYJ6r+pir1ki0TzhvvYk3UmKtFEdA9UfdsT7m70+2KYbMb1LVeOCxdarRZ
bOhcFLZKWL3ovb3re/eiQTKcSm/XuCVf2C+z7wsjxF7gduq3fbRGgg673rHqow3LRoD6IqbPWzaX
ZZrmlMkAd+84M3yD/8gVqkwAzriNtpZJmIwqNeeXp8WA93dcbbF6BnrRxzZSwLMQQmRdY7mYdL7L
/n6AHPdL5O1jjsjBud7AUsfE/ERmZPVUaajmXRPvPWLUzlPiIObG8jfDqRDNFfkrwivmSsNeY87J
oD8V61gojPfhl6hYmibtLWPIcVQDqMbF7eaTDdleD26dQ38WjgRD3vohVj7Y4he8gWQCYtF/BPPj
YL2FL500HC6la1JFKT3V/PCKV3Oj7fOiXRgLbXkPUzPhtOIYnYEoFivigTQpMIlUItKQMVmTXH47
jB3oM4VbEA4yNtyqSgqa/0X/E+v6FAB+t4LnbG+WkWbhfri9qhUQtKpUep30TQDOV9KSdPipNRmg
LFDZV440xnOYXqMje/yLKH2PtiV0yB3VQ8eBFhaXD5ze/rriaVbyAmgr9Vcmue7RaDBHDkwfFmfr
XzASkpMOx5IL71gidBWCNKQSw/YzYsylyqlIDw9pZx3yFyubyuv1KowjGJag0hULdGD5bo4DRHeM
WvpT0EUjTuEIm2n16TmRlj1/HwmYqL1D9yOyUC3eC7qnR/+QCsmFFHsl+GuS18vomU3xOUVQnekA
Dt+/92/W+T0dEACPV2F579L1jXmYxzeCOEP0fZpMim70vgMFTexmjEzyRHox3wwBg02pPXdKIkHe
2NxbryY2hiI0iWDu7O+nHZmYjpJHDeLMqnLFELO2cpnfHototawfhXTQfWKo+EDYXJZn+62F/cDF
DIQhLtg41zLfkYjMMZiysTmkkwpw1Mddbdkb3SuaGdiQZ6YkqIeXJBA1L+jdDC/Yb/N3zQ819MNN
b58M6t/VlRZj/NkbwBTWIybLE5aXsWkFfBGnDR4bCJYKfNvoC/Ul8kWvvghhq8woUhtJW3dO6GP5
IaF19eQ2M1w/KZsXahrzaRubnmCrY1+zhVWNBqp9YP/kQlSA+773yfSxtdpUSjTgGMRKZ1VKh/XH
P+qhC5dKEwjd5qAGTuqQUgCoJkbEU1wxqezR4yBoGGjNQ7W4x0hHEz2zd3usvG1f+3FbwlIXTsDe
Ps+urBkRlcZ5u7AkIx3kID3kvXScxMzeSzgppt+hxxAcq+b4npNlt7O286C65mBdBNQ/5tfOQx2K
TqdzE7r33mlBiHgltchADZ1ankZJNiLC5vqXphF6ufRzin5BfLfqX/xaQlZkXSwVbKsn1f2uwjF1
cqRILe7tbE/PrFA39aZiIq7XqrV8XgryZTTaAlgPcU/b4xED61J0fSgbpbHzX6QePdjjkw7VW4PU
jmwT6Nh4XVYUscLyyWn/lozU8SauCeXPlk+6EtBHKxMoBISOMXY9a4nmVlFz8ccC2hTVIsEGy5Lv
YMFplnQjAP6BYc6V8rHezrOqDIRhkVEkostUTs5+LvL7WW9aLdVfZy5+vjQuZ0py0h6GlOF6TixW
hew0xKc4ylHdV/4U8DfovYAgPolZfk6URwVxiPzcziS9DZ49+QqmVgxIbzlfy6fwpOp6nuokn4pg
IZnBjCm/R93v7dBIP8Nqyk80wLY5fyLbihAvbC0KY5ynzB+CO78B1IPLiVQTeREXkbYUuTrOFDYQ
UQ816Xekkmxg3AwMklVnL2SFbYVmZ9tPTCrogkIix2/NHKr0GC2FnZxS4vrj/w6CGYoT+x58hP8V
ppNU2O765hvCZtV0MKFQOJUKbzM1/2AOgU0wvfKFyviaybAiXHNtCydrBklKmwoeqWVsuI7ng/9F
TBByrjk3HeRRSXP5LPlWf0Fs7Fz0eiowgSL/hGQBMdkap1A0coc6YqTEFPSgq9CXosm1elopBr+V
QQw8FmtmTl8vx8J+tfVlYQHsBJMpdRF16iXWDzb9Zfpy3O/H7lkRS3HelshAfbzK76x6xISvzsnt
AG7ev68adVmcwTTkYjwgUZEzty3RrziG16uNWpRkTL8860i9XwMwXTte9FmnQPZPf62qsDIt+Yuk
Q82zb3Rqh32eVpD9ENO4t+yDn771iNdlK22Je5u3lvLDbCNbC3z8l+xjODYqdkYmmdxipi7E4irE
pgDxETAdFNYuIismiKl1mLYASI+PV4bueQR0YzBBjpZl7AREWsBtCFpzRrvgg99b5pGKDuKIeNfJ
1ndOmpHKbBGyXldxZtNRzTsvFYAKOdXRMN+gS1UB6yecrnd0orpvHA3mVxg8aLDOpsIeW86ssMto
ISTW8OUEhoVH0GcFWs/e10YQ5KUhTuPPPf0Q2gkYMdr9d9ROxA5bfaoELL+JJAruxRMHgPBWBWLu
o4k4ymFl7NzQW+fvNLDvMqpTLLQoi0CsCleA5XyS6m+8HK0l+VpkiHhxHnbn6GK9p/JKKFQv4qgR
hjS38YSnEwANs0RQTVncebOJw6gT/LXx7EZ0kLbhz4C7uSV5bTvtw8TPQubHBsQZR+6JYHoddHRH
aFKjXb3y4Bqb2yFG1+ExSMHaYVtr4Ogn1rast/y0orhtCoHEQPB+hsyFdLvt/SsyY1SkhwPWi8/Z
c+Wiph5xnsIbuNHfHj49hOCfsDXKGLXYVhwGJyjiRVQ1oDP7fvichWWvwWH6yM+JLDGLXG3L0vhj
0OBO2oah5MXqd02gFhAXcN5TjCsh//x3LJoPkwfrRwElHjEmVlsggFjKy5IHgVvI8qGRmVLs53wG
lNjQ0wcWaaHU/HfTFPtchfbhArt/stgsN4ld6dMvz8+JYGACAv51RH2ucDZNMRK93hCZTWnRA0Rv
zo9CHdrqVeKlRb5zGFbtmZYJeFLFfl9H2y6dWzkk3hdRb2P7C+h631CaL3SIjoC8CO9c0hUqEpab
gN6A8kj4q4aoyMuFGUxzeV3xxx9OTJv7ciOtIX0gZOw0BYMjo7LchR4BAtSEXEikTifcZr4wPbSK
YZuLaNjth0QafVP83NKZOghFfWcDU3d+SNQ3wSNuk7ubOJOD/byuIk2TcpRKUCZj6Xo9oQKfzkvI
XF4hJrt0g4uNQe+82LmLXnqORdoEsY6LIyErIOsrfs4aYJMXd2/Mb9QR9g6szvgpfiIuNesMCICu
YGT7pdZsSPo1a54k5mR1OVqOdfxwwAT4wkSTZURF46tVMk9h3YuSwJs+Me8cngOY8EVJrOSi9SJ4
OcJHrDp80qARHQqLJBsi1T6YMjDZeYhvSR8JQAnlKrS5Kf14Wi0dbdl1WyM0d5YxVQGvwdlzxvzm
iuDhPjhsNaa2lFxPjSDATMOyGIa8PuF7Tp70cDI+xjfEyenKqG7R/VLZQZ8VTyyacujUUth7UN2s
bJ+iY0TYx9Rup6bGsZWbIE7a0TkUXbgK7zjhm3RpjRz2LsM8/NaKQaXFvt2ITE8tc+OFsg2DSooY
oDpdAPGswrVqjYWF/X5hWv8jaKDcWGUXbe8wgvljcupqcHTk7q8EiWITTxLOPvfknR9qgRiV3TEW
p6eeKbri7kzjew0Kbj4iZrSsE0RqwfJ9ZrBXk9cxlggTLXWYZtgeTMR3MUjUZDGjN4E77J7y5ul9
2zDdtUSJuRfemU7THLfvnc938iITXhOL4HPHgGDhwRwt0Zy3RiVlnNdQosHQJg/BOREXxM770Th8
vyy+ksBvkVJtIkRihMexu09w6EGIjAugPuzjYOiQCLIjHZIOcplwQnoHEWC8HzPDbYw1JIbmzL7T
8MRxhy0TGqWVflvJafx0SzYNr1H8GiG1yBr7K0olAlgTBZjGQN85GUrv+ashVyRlgrE7e6XIFwzq
jH/YrQN05N3/OOeZmJklef2l4w7tbWQ5t0I+8kqxDjjh6X4nivn3pGvxffSIyyCb1YoqHfmRzo6H
1kBpYyxvCjjPWZekozLEsxnVkoqyIBo7BBjW5qv96bWjpnHrUMkCqLwymLpKapaL6ncXYj6L1+To
PoBVngX9DfwbEqjRsfkYIQkQHrsCUErPPqlkpMmO2bS4d/Q6QPGeI3e/AjkifGqZerS4UEl3q0kQ
87kYC/I8dwURBbke4sYtSUP3PpFap5XuV6+CZLvvNWRk8pOocJf0vTMMGow1BKaLESGkJbLAXcFW
eCir96gPi/cyg2jagjqGFOINx37dHRTA/jOlSwk6f+7CN7I5P+iC8mivE09+7EsTGCb3fMGHHgsj
ZvUEJoKnKlJrI6MBy8p5R/l2lllJ7Jc3s6TQJnKuAZrKqdoJPrM+Ik9+yvbS1WTFMmjqBpnOQgTm
mk/OLl0Bi/ljfIeRdu89f2pfT7oi/bmddCIyuGBOSS2NMFN+WeAdQk9nmrpIDRFxVAMAA6GBlxS/
a5JiNznUrp1ZsLZJpUpGkicI7n3CfvQcnkEzHb+vsP5nri7iAz2r0DVOa6aIWYjR5RCCS/v9qYAC
wXhuuvtj+heREChO9HK+Qiudogk9y6LoaH/IQqyyjKywf6LSxGbkzdlzrD+q/1SHWcG/KMA7N6tD
KFVNtNhlrmjAtfuOeY9/0zjBUdoI2szWgfAS/hn+RA3oBVmdSvjx8WfPkRe/jGhETw0vOKNh6bpa
3Vs3diRHfJdqDkrAtfiwqJluP5cXPA7EFnoy2sP08ytbV62XEboSjp+EFtbAmzYIg6okM4Y85Gii
lM2u8wxvOqA0CcdQAUZbe7OcD0BldKgFF2xBmzUiebq+PVsNyvMxm3Msq2dl3oueFfCqWLm6ukvg
5UrE8XGQG2I4X57KqFXZ/bI8gAqZgT2TLY3M1+CtfTQTYXNa7schb9LqRu7GC5ZF3cLApidKSrAj
iUYMhpQyJMVJwxiTRFCPZ5ZW92tOxXSlbnNlvTvYwi3Vbb5dzQzz9oLZQ1QX9ub7v4rxQBiil/io
LOjkSsBDI4XETbnofS2PNgxKcAn56u4CJYwWyTwv2UAlhJPMiXBGqA8SCn09PUuPGXX5IY/SRLQt
j3iaroLwEvJjnDWCb81fzCla2I2VxCdvVsPmUqt9puD0pDQbU7qa9PBFasPA8DKxMAqv3WqAmJvZ
kLcW/nc8EohpTPpBMxzl/4VwgWrLmjaOe72Jr2DGlQR10GrETDwvCvhqBsnyY0cCN7+t4rEspCVw
4Y0fWGaBN71c28UjbcNYB++2O3XhJKmIA1B84A/8aQ84+D2UhVGLkssAMTHYlQsUnuAianNsJUOx
YNOtJ2P3Ow7NKnQHL023ooZA+rZx/ycPvilRIy0kqWhLN1EGmMU/9Fy2+E7Bhr74fo6ueD+NC4ja
LSr48msymk7tMBoe2N0jvlBYZ2KTlbYZKwu7toY9tA7wRygxkAnFWPJOzV6HpmCcmNQg81WOsE/U
PbpC0XHNyVsfkt7+TLuPU8r5a6eL7Dqq5wIjCR3y1GrpuN1BLSmRlk/kZncZ1/BeOln2vO7MU331
U6Rz/nwKa7CBumNswlre0+Hzi4hL1tlWhSzVPVj8sD6pHj59Mh58MzM0pt0xjdC2/kZGVaHgH7zp
CT6oTziJO2NsYqIPqOkQu0x4fNowId2YaWrff/K2dJyqZmvPghAtyK885LM7/XGbxWEq5+68dGD0
h3I0gWZa5FWq9kZZT+6ysPKEdWMUXv5foJE2GJ568qp8hZv2yzD5zvAuiq7vB1QgTp/7Ig8dMg9M
tfpGxUFv5bAknU80KPZnaK8zTwxtfqF4/y10r/E1ZdXaxjMv+A94gc5giW93ajQ9IVzflgxnltuw
Pf+g1TrzvnZbHuEdca1PWCOuIUpeQ98bOnidEriDXu837AmjreL33g7PGfOqAoWSwJKqlG4mpBkh
KXLkXM7bbbTbZOc/IYm9ynviFvUn1EbsU0ieXkN13zFJg/2TINg8g8EwoUgSyTrfA1L5zJOTY0O0
ucSTFXWvIsyWh118woTVHWu+c0Npnynhcj1Y2wg5eesabI9TlWun1kcG5krH2g50Uw3IWxlQtNMX
va+9QDe3ZzlZXPMpKs+92PBORoDfQ5PBxgW5W3/cE5oLXD7aqJbyJrqv5EAEf4CiqIZnoUVlMLVS
XD10dzjR7uhlWbnyD4Q7RNzNq19Fi1YlW7y028bIFw1bizzxAnWW1jskc3VU2y5ocLdivU2/yDZN
3D/RNHjPXRV2Nc8/S3hFYTDooad1xtwpf9xuXAaO/tN85ptG4d/V2LE67e1wqM2YCCOSiWtO/ACX
gNePxz5RT+F6pIAgF3lfB56pUx+QbzwHVVwnsvcRBC/0k0mwu8QSn5qRlILoG4WZRMlfW+4ZjvKf
GKllEfbMIJkcx2pm/qiH/13H0r/E/kvYL3Tzk4gGT9ehjtKFliOhpBummgo6IxKVWLshPXff+yvb
oNuUDAHjWTH6fnYcWe+Y0kcd8g7M0fRFg91hzjn801mjqFxk99tg0OxQ8hWSNOoTBH4lDuHZLhNb
W7rnq30/b+vcxjR+diGyWeYcK9vzMKZ1/tD0ihirivC89F2V1vGgfa/CVlD7eyWYHolM1b2TOeha
WU8LPuvhKOwH0aWyi+M61UJtNb+w0Y4pO13QmIAEwkRvKpg45De8d8g9ly9vdbVMAMPRNrfp/28j
7yQnbuhBX+mvyZwSAXJaRfCnj6wNPz+qfQc4P9av4uYcMaUrTi1FwuA+M9+yfGCiovT7hPwayxab
24t94bzx2GaWiiy/ulH15ONcTYLqt6LY8EvWfV77KxCiZbUTnSCcwf7N+UyjR2EZ6kiY2O4RoSxp
b42OqkQu9816Dwg7eIxCdZlmqlGbwqWB+6Nan6UuUSLam4WSjt3miNzIr+i4aoHG2+4JQB1QAt6Q
fQI70EPj3oYYisTIaKKNMI15a5vitJ4RRN36DwlVyDAl9uo+HoDbYwhLse9vr450fNAklM5lKi1g
/4s3I1Qf9KxlyhIzAXk6t2w1teWa8t5xPg2dBaQSyQuMFIu7TyHmxQhxg27jccGPVXSQ/R18/5ZJ
bZ1dp9CWFBSXXShmixjxVSsi2IdgQ+I5rO9e0dMCTRCE2YBlc6q5JZ1f3U/C4KVG9fUTppaMFtqb
B22IHZm+tqcQNtYzddJhedRKfV6umab8NrLROlbY4P+ifhLpbT2RTzOGQA7UYqEaxTNg2bn8nyh3
VF4WrS1kfUqn864Yrqu0tzrIcjqOLV1uGmYh6Begg62CZQX9T8h7Y2D+SF09rslmTtDhL/eHL1Yt
Z5xHNVelH1tVcSjwkLRqg0/847x3f9qDutY5AtoUsNyYiKzjLHcxCvlyUsDwyc0fFcu8q4WZd3L9
Kw0YmjOlMmyhg/tOivl+ruUiKyOZqGShp1VRmzfqLSHB+bM8aUmmNtpSaD2em88MycGd9LWPmCUH
JfdQUoOdiriWTAuHAyi1zB/rTiK8voib6/S49bSHP6J1qGZv04XcvBI+QHTNrRqzbOfxuUQ517k9
P/MR9toexHmoXKwUtPKIloJj7gG5BdbM1GsuTVjtKmpdKIQynhJUIVyo+x19ryijWA+D+2jpDAuU
ecX40XBteXwlLUiunVqgQFmq8yrET4qhsd9t9KSASxoSR+PB4FssFLVfy5rMr30IqZVe0oFnoaeT
XbQw4hNoSwLWCt48V9fwX6Uq1qI78C1fTo7n6/kLnxDKOtJG8WeSZ8f8DMaMvIKsQ8l5VEwPzDIu
YGed6i6MfeCkOwcTlCFPSVpPQulGqIvAXYu8bIsKabXoZF2wRY8EW7Ncoe6YpLoIKFDpRSeGZYfI
1V0eE8SXVhS0yuyeXll1XBeXGHqMAf2ENfBfsJhm8wPijmcxPSkLTCW6QGChuaVyceOZW7vTYFGx
OuZjxTKB9ZFJ1S3tn87F79bkFHdcs1X5GgMt+se1bUIf8T6x+lbhbG8+86HDX3d4I3sxNHM1nSl/
jOqRcBbHF99lgf9pESMPn72Cf0Yx9mexCcvwrqvdOvsGmAHOJyguHblHxU8IMI9lPzsO5gh8cuLO
7OyLooNEgrZdvGA7RBOi6HYF7wHNZcKydWiNhmfR8Ow0XLDWhnFjG5Wa4ruaI7y5qGFa5WiA9Qus
E0y46eeNpw2e5K4Ni3BypXpsiLcrvDutLSTbOB9L200HxyXZyaDLTF28yXZuUMspUi1v1RuIgOWl
zYezmk19Dx7DO+ZcJcBT37COJQutXFqwtQ6LIr2qzpYnLA8G7ys08BhRGafTO+a7qjY1hkTzUNz9
d0lzkY3Ktzee1Bn0dBTXJHCAUlQfX4aZMghJbt38k6qOHZGRf/kzY/hAfmC1kvn1uT9eF3G765kE
PVuYYeqyxjT+Ml05gwKBcWoeQMtbvYtOj8P6bO2sXpHZ/eUyxxuP2AfBvt7nP4R94QijIVKOWJ4H
tzaMUH5wNN4RBNRhGvR2KSYnC6+J6zLiYwuvhWs+d9Gm6PTquLIy7I1SKfUqQkCTM0Z5V60iQTrO
XA+JlwIT07/BF9i4mxkJA1fbPsdUlUZMjFajOSWIB/b8mUGgLI2RYDY9/8Y9db2BevDhIbf81bO5
DYSne9mnEc38VVHHsU9A9UbMmIDbQo79sZnFE4Xvkqxp1D2Oxt/xpIA8XRZeMcrMO91zRLIa6FC+
1HaVkAD1x8r0figKnnqzo5ey2BcUSspsKrw4YqBC4WAQrMdGbxONFyKU+e8Sx1S0Ne02clB3lSx5
6F90zinTJPkiLjTl4uZMO0MichkpghaLlMLSOKpTHIChYZYJi44+skawsGqWvkbk3iDFDDIbwNsw
8zJeGi+SXhYc0wpk6YsXvbI1pMUcerQO4fSiGr4YAOYCfUEwUW9+TIKOvcnjVQR7KzwUaakz383n
rw9fx9xqYglZFvL8bFKL9Yr5u/nyk8cwKZsRFI/ddfGh3oYAziMvv9s+pwbrsFJSshmhwKT8p/0l
c4nhJdNVkmsfHOXE+HnU/ufpHdCq5Dh5xaIqGpoipccOU+Ogd9IaO69fec0qttiK1E9v+YPHsu5r
XG3bpqI5/Ea4eE/NHu8Tren/aBnC336+Sf7yDPE6o+wpmINUVkWwCmSScAoCJhufsOKpyGj/VNng
dKIGOTyCOP60oRjrqunR0eROfd/w6b+IVFmoli+R8/4/7/IlgYjVQz5ssGTEYJiUQv7mwEGigvzW
k39tXN/G4ztuEsMBDApwflAyMvdFb4fxtMebSa+/73c8b3v25nMBMrz27gCssgilwKWqbjxnhlJf
8zfD9FsyAloZXvi2un4abiy+S0WFw6MBjiwI4bqIAbDreus9hqE3YBCB4h1V6Id8zlRV9zjcjJl0
SXCnvHe1vdtYj1yR5EjaZx5xRu7E9TdprNq2Q1woVeJQFmVjZI09MsmS/seINA6UhH4BHmdo4iQJ
0fbm5YZYF3BfiPNdXbtwcKkHOqofk71ISp/Fx52PoU+c+9bTCODRmcho4CMcCU5mImnrbs1xzljl
4rJTHh/siYS5Nh3ZK24HITgLj7jrGQOwnbYp0JK4mIfoofbhNHHOjAAWbWPwGMIPaUFciMxEZehc
/TH7zKAVNfSqTsi+iVQCNi7MtS7IRz/G3ZCqkQMUQo4+rvxk175MpKurIWO4yfnY1+gR0DWH9sgw
ciklUSWyMt2cI6dIR9baQojhSGsZRPiMPKx15/HwzzuDu4417oTqFXzLvDVv8AnAkSVLplLTQ//i
3dqZnzHXIUoGexH204tU0C91sYYbDPK3m8v46tR4b69j8vuLw/Z4hmMZIbRV/u3Qunf6jybCNb97
kJwWCOM3ked+vqiItPkJb18bWb6xphWQsZ1EUs1YLR9PvzEhCuQLngNCgVaXdccV3bTwkV5eHqWR
rZVgZ1Dxk3QRLvXbiZPnONfG0aUDOvGdRajjKdHL/RukdvMA7UxNuIDTGsP4mrQE+jCB4QvQKn8s
JH2QWry+zRTEaDwfOdMUEtMuNjlAu3CBay7V+jYWJiDRKWJD1z3p+Righ7zzyYuJDvSaDZEnWuVZ
tw7XLwFXrfLo0/ck+hyZ7x0dX/G+xikC3saqppkR4IqPZFTuaX9SodlYe4IVKCTP0mxnVPeSfxGU
HF67AJZwGm6X4E5uj9s17dpx5VHJb4VGHX7r/7XeTfAEbN6W8MzFLbonJJYDXTO6EDCfy90Y3KZ7
1yiyhqt8AM+IRTnzTaSt/izWOR/4xufP6+bcC+fnOyoNKN/aYlPHuqX9FDYDtJ+iYFjD4aBcbCJ6
xS2xeZs7BDC8I0UalHFajpXRzrq5EZQgsMwSpEYnU/rZktiqOxyFL0nOwCeQRN90iMvq16tv9IBu
m+8WjYMaxjVWmq7kRPVgh9bhTcU8mZLebE1nMSHDuVbmlkNB/vUwtRqu1l0saisBrx+BT/0wGAfm
PTGtATJtXtDxaQMQfGxg9Zo1uquiGx+yCcevcfASGczwCNBCnRnZc61rbNUJD2T19Hfy7u0ULWkI
u3CV0gStvguKu7+PqGjSpYL5FXvJeDFgYyuYqIABoah5eHGmtaJpkRNyc0NVxN9mfxEm8Q13OS56
o+j6X0EDLWKcBjClYFQCevz2US0AQ0lXh9NTLllQvo729D8yyrSqQPt7ILYDCnRdTeZWP9oY6q1S
QXVhbouEyZYT0PIn0d36sHIFo+ZhbFvNhFKc20xg1HCpy7PP6CmQ0CiAXIPUCfS5urjVFkwHgpfm
+1pai1/7UHWdwS/eDTGWG8RmxA1ySr1xsnyiT3vSR346A50sIhUh8UOKa6JXB2XsxRdi//h2NPg9
qwrnoUBMz0sWIM7oS1M1Bd1+nuPC9saWpRokallxMVjdjWf16FnNHCLNTdnazvLMQmoocC22xg3v
kWOu9asHygQhzqYIu/QaE5/Ag5xJz6AiJlb24sXy1TdZn8AV/3rEINYOfEI25QoJN97aOs5q4Q3x
sEoF+bfQfc2v4hjizVu6zfYxD3zo4CQtjHArPYErtZHFTHDrwEzlNOE24Rd9QhPfsLXKLmnIvCFE
DMc2Y2NVpUefVhXGgjhBmigSabsgXZPPOmnqXVEAMo8AmUe8jt1CjN7pF9uD6+evU7EtJGad54K1
va/onfGnOxhvAO7mLXeyOKCPwYtc5wpNdvveeAjOMe5IDlV6BKl04EKV8sraKZHnzJaPkmJQLOy1
SprI8ZYK9GkLo/i1wxz+9ee6TZAx5XMZHKPSH9CdTBDGFVjv5YKlm3DzgpRWgAHuLkvKH8pmhcZl
3k0THTrh62eXdqBdxJR1GMeZhIdDxFa15/kN+hDreTrVSXzRf8KS5350xNj19g+z8dI6OmxHkM2o
Ds/E14iTk2CiuWI/r0ViaCA2N1YCg773XvklRvTOzZWn37AiMO7gHkXV15daGZlEFiMPx97Zbwt1
FOSj6eeqgM6X0WO2B8K6BqAWNzFyTboVLMz78Hp2bByiiFT7IUPbN+Yw+9SWf0Mqpm6BZJHF5S11
tBHmzwWDKLnVtnwTHoSRUxKbgPeKXLzobu8RgFYNFoXgeI6aqwA1dqjLyIw5Un9MyyURRNf0EUa0
hLmVqpaeFTjyocSarNpo1km6hwyCUTZ70u/Kq9xqe8zAAmwkQIN+4TWOK/w741g3y1AGmXtNVZ7o
8D730RI1QVkxRsjNBgGsQzHTzYXM33et3Tx+ANZgUSHptlm0ClBg+TnPQES2aDS6JSnw67SvRdjg
Jn+yFvAfrMhiOkOAty0+DgBvlYfJIDTC8oCuLc8Mm1wayHrw7MZx0QjaSLhP9li5NKAVNHNLad+z
njZjV2BYCj/0IEz5ZZNuG21A1xzfZ0maG16zFGC4HcPslIaCE/k9hJskbnTSezTtofF/InTnL8X4
AtUABGXCpsOBZBs0x7C0NM2tizkDe9lAzXnNlmySZXAPRXMwcrOlvpipvwHUcIN0j6iZDyZqhiTK
zoYgXPT8iYJr4HSyhuySDcBiSaUJJrQBXKRxvbqJry3YqwLu6CT4Ny96xj9BUe2tpqayVjDt0dyZ
O3gLCMcgzpEpiImoWJ6QWbkyv5Wod8zvwxkQstOvSBbJTebldz5P5Nq0aLcZSzPdlXnkL703k34N
ULMkhBnyzR7knIQpVc4fbGOAX+YSJ78fW6GE5vCfo15+IDRrmSwuCD3B2BZD6EfwhZYxgvZ6zv2Y
lZvK7yTSRwQDmZWA4OwXa6/52r6bx81Uc34dX66vznZ25PK/0qOiesC2j90DU7O/TrWmTLr1PxBZ
xeF1ckxWQ7i0ViM0Tg5XErP0EnZLd2hwSsycLTReckJrSalluQHeCCCT0mBpxepta1ZCNJ/XgyqL
eOGc33POXf/2pHT5xYY8ZkGJw8xM+dpDsauAs17gmugOTrDNpQvmF+wBMxglK7Vi/54k5YsPQJHL
E2V0oJGgSpYKg7tfX+iWGxH4lVsn3NCy3YfbHU0eAeZLh/aOSZoZdVk91jdGyQW84cxdGEzeghMd
XO8L46eIvTs0eRfT61j8hGMafQE899zau2ue2QFRMDEr/5lO0YHRKuhkTg7tYx5ftCCs6ztibBpd
eVoCxyV5rUE7Zdq3ZfGdFPmTl5sY2o+ceEoN5c423W0CLcjltPykhiYCI09ddYlemnJISMEsxzST
AL3+5WIpjKSZaJ2jXR/gJfqkkk0V+iUMITrxaf2cI4ZfyldVnf7B4gq1jS0G8qRphh8FVRbNkic0
skYK2ukVQjlz1UN1zv1hXuEVowgz53KGdoL8OFBNDwgSRsISlkr3l3H6iL9MXxBO6Wu+nEtF+/fU
29sIAQqBP3CavCBco/f/Mx5h2JKAUm7mLur9+PTfqyYW1LIBnubfWEcU4Xe2VO5/cj94aA38Wn97
veYeakOjZGD3ArwobPUXcQ3/zoc3VvAZGKtU9LGwhkEL2afJMViNVKfJ4Re9aNXA7AZ5P6tA5628
BA9020rJp90iRrjMzLJvTblgDn5MgLqcsEZzzScWjWDhhgs7B2GexSBHew1SU+17MCkYz5LS3NkG
OKWm0fzZ4n0WH2Rjo4RH9eizPG2T+JCUtqkS/eh+aOf5dlzk/14HGeYx6a6AKVjPjxHaEDmgVEbX
YG9X2sJI2S8VIt2EZZl8mUfdfMRJmeuPzI0QBNCbvC3hok/WS/cBijyrh1tZXMu6eOlTn+Lpphad
I39szwZbBK9WPdoJbkkEAvdOrTHHtyXznaNhyA1hzti0NuaPTYgxJ5Kxv0uFvQuZHKUx15DIZzNr
/lJmsyj2ML+HHtHjpm20CwMX8ENNm3nT7iR8DYVu0lHqhLiBsE7FSmsBcsI7u87pYNN+CHuEVAXW
3twvl4QGk6fjUM4G51j1vbQWnqp2tGAzqxtG/jS/Ms/APWcdteuKjezGniTjWa84lgzNmxjp78wi
ppJ5Ml2mw+f7Uuk2eKif28IURcf7voMJSu31nEwheisMYrpZMiYbCuDarrz5BNW0OnExS2T9cT5C
ERrOwjdqVaCS/MONAbs0Is0/071H9hN7yOcnLU3i6koTcmDfrpZuxVVOY+tqs4vmej2ayac4czbF
e/d6bFXpc1SlfwaCPLO98eieuZTegKaSIjgkcE6c29JAI4hAXHog6P+pud+4CE/7nchOZjJ56Ek6
+z7/kJoMtEu4QumlwiytrjAdL4+rf3yyRBm7cI6Q830CtUhehyGL7Wv03cXft77gRmq11fGM7bnZ
V8O8gW4XRr8HBgRLYtgDFXF10YI1tE7blGMJwT5mVCzmgPClOCmVHvTqH4MpWyb7efySgiXero0G
MYDfao7XcsqAsDfVFMnqLc2k4jrfZ0sbHetIiz9bsmabw7kWjLEHlImmi5c9JE5RMjJG3SWbuztw
6q0zDjw4UVzJHLWn9niWo5jp9gdtp6/IKmzxDFtjnoLuqvZ18USaS83voeVRFBJRQEAGmSqkuUXq
95JYqq2UhITZV02JUkQTy6IB/5+EPuiJz3EXWVjHgYvtX96XBaYC0CAv49h8PaOXjCG7vlN/m4l+
nd6Mwn/23tWuGy3dIg75riTZA4QFMj8mVilt45emMDTpzjmHzaUpemM/24rOP9VKIOtkFI8P4Xsx
e6eOC1Hwg1JgsYcS/8K1wVJLuxG0a9ggCUQ6XUlvPv2TFpw7UtoC8HyOa7wDdofKhrrzOP66AhLH
j+Yne+ryvK/hLLRU2EfHY4stq9aIGvTRij2hQitBKo5R6nsccvnWEv5pjjQFXKUD98VYH3IuxmXW
nN8NpVT5sjJcJwsHNr4KSv6muHdHVMeK7tNLx7+DFzsw+RSaDtifKC6qGY3BxblBff9YkkAjtivW
mlegTGYU/AgbiqBxiMhsNXtZ+WG3W16WFFCCDhr3+aPV/iahJKau5TDt5IIaaFcSYWkq0SrBr6+D
FRVzWFqODPf7B4byMclTq/aAU/nOWXYEM7MuuPCoiMb+7N6PpkpwMSnLkVr3//8tke30byDJY4J4
CjhwwQfpIL23nDvm6q2rNUaqG7U90GPLS7loZ3L6KQwvePh89QP5r7jdqXYxvO9AKpO+0Jmp3djK
cyWdvzreVoAu5h2uT42odmk7oVwDKPb8S6AVawI7uUT+4BPpg0FI2Iuk74HU4VQxHQYg+11GF6YX
sSt/ciXwsdD57iTsjoVsViHnviIQBiq2b3EDFLcXqADOftMPfG8nIGcssOX2MelBwWLoyTU8HpoI
lHA7K7xkNaLezoKbU7BPvSG8FZ5iMsubRAEDrYMvQPN3wsQuuEUaYYv5/wcxQw4oVRX4XTQWbpaF
wdVeQKzM6u05MdKgT95C9r105UyoaV1HlJuf5WZLhqT9kw09wjU6rppd/PxUKwyjqNS/1YpnHCnZ
0fbWDi8OOp9LfNR2Y7T1lz6MjArIyR2pngZfg+qUdBtZoLhxFXoGbn0lAHxdZLRjFN4PQG3YY/SE
UB/jUuhIp7jnLSwPEbeJdSX5bZQeHfySqBsSC/yDDEBxmHCEZDDm907ZDNHuoohWiAEI4O40b8jY
mmhuJ8QfBEgItSM6Z8p/2nCbrvibo+NI6CspPqqxmRC0dFwDOrZfHRb+5tzawJhTo6auUvprxfQu
//X/aASiRuF0L64iMdJuc11KHS9/lRrlMh9+EgaA5GsWVM7f+A6AtxxoRKLr97/AQyAYA2nW5Vgs
Dauzc7Z9pP7Z0lAgmIJ4Wzk4xGzUzESVSLubMrDvyb9YQ4r4eiTY57QFu9xZvwWd1oTdT4t8CHNX
2legjJhU3vswsQ7cu5hTx8iMO/8RH/081BUZeU4gmCLRVGGjudrb4G2M4CgseeLwaj76msjhLwvU
liMNlwwG48CEi/fV6+GEJgz1/w4zR/xhxiIr80K76fF/0DUh6IDz/9VzxRSk6nyCIeCeHDWCUvuw
dUDsW/jXB6Ny/306KgEIO48IIVkJ1uY0wdPKv6TRUbsFNeLfanI39P0/9dy86N5RqLjODOi1LDC8
zO5Vi+6YV9NscFvBZyWW2GQO2TpNXz39fkLbyzRJvMEraw/4sLCYK1NfeFr/MPzHAn+90GuyniHT
dbwbL3r2UKQLuBaZKqkjWldwhx+A/zLJ7f+kvjj70hEkEP9qrAllbl4uD4ykn1w9Aqc+NVUnEZT3
Un9J6yj9Rjg11v1EYfsEWfeitClhyIl9+qs47JvnTYM4wJ+KuZS9ygQ3+gBwFSSSb65RYu9icslf
K/0iiYYfYcdUgtglURDlJ+vMIBJWUxpLBaU+5uhPWeBRn/9HZYomN5HS9KL8lQIeGC9/RdOW41jr
dMwTXG/ajgpjUxk64FNLzhqTOeyGM07uAzpLVJ2bfxdRj3Daj3WTvpC7sMcaNeA+f5YTpziXTUc3
rxj6QDdq0gfJJpL6b3LoLWUOrglRcdVARoA6MwSwdu1twUpLBNiczs0CvBPnC7WuTUKHj49Zgyow
p6xbWVuibK4wPiR+LRl/8YdfasA9wYn2F61O4E03p9iXiVF/ZwEYtXOUs3zncJWmVipPQV8UW84n
FV8RhiHpN36cLGrHFhrnN1326JbDtrfW2Y1ANJss6txTHZ5EGba2nARPAd32VtLSFu6gpIo1P/8o
Vyjl/qSru/7yZR4JcOEjA72kKaZKUArCcBq9r52jso9hj3lCLeueFYeofhJP+F8JTGOMS2d13oyW
ElcKcQ60TSMsJzuhqSd8rtcXG8bGMCXpxJSh3ZPeqzaC63E9LvbZ5aORVQpKbL1fN3onI62CPrax
trPQN98i5OFomHnlUtGvIUhMlVUrJaR1QM99HvIPBVL0DIzsTF+adGxwO9B6OzA/mLpllewsKL1l
1uC3oJBFcwCDwUpkT/rJ3CkYXQm4TCVqIsizGPmCQNG7YDOmvV8y+WryRxPxxgJxOzGEw8X5mxDI
1fltpfDToiKg8ulwJqQpp5WSmnI46ZXG42JRNpSaJYbKbDJUXsmnCC5yeLwuLTeg9hOSyU7DVV9h
tC4O+LcmQ4tiCuMv1d0cH7Cj5e7W7S9voDK0VDE1QGWW0BzanKptC9o44RRBIUOvs9U/hjD4A1+g
KJSu4LknKyFweTiYX/7R6+guiAQqZXmbMb9BOFEHQ96I6JfA8sGYZn1bXi/eVm6mUIGGMW2klcpe
pN1Q9sOsMsJo3M/pHKW+JGBki2cBqcSXKkhE5H1QGww4G+oeqWuPKkisSLPRM0P4AyFa1DF5gd9S
fxq2cpHBOwh0lqKE47KUn3QJuP4GZW/JuGDF8p2Qu9LvyLkNBJGL/TlVRaPrpoJnpS6xdCb5XNoq
Bd04CCMvrLFvLQHO8IgQyBh+QWV8tCDXEUd9ln0w1jQBqQQpNz++fC9d0SDebCvmeW0RKFXCknJW
0+Q26VFsbMyHuWO4xpaVL1iDMvwBcY263lx/ObvHd3wA6jDqwhAih/YX/Mlv6YV4uT/whANbXXxl
dH3n4OJXtEwG6k7rKYjV+fG/HPzngI824aL2TJhR8HCIb/Ef5gJZIgBhIsNjH1a7TYR8o57TleP3
ySoW+ee7hu2PlhPf5dmWL1OFZue+DKDFCMjJF4HccYPKp7OhUrB3wQTaqbz2/Z0bKk8VS4c+1FYu
9ogoymYUcVw6kbKRsU+VpWLM2c5yalViR2P0K94hkDu+KJCe/72GwVjkQAyY5Kkrqob85rla3GFv
m9fzqI/HSAHDnR2ep/KRxAiDo8LM290AKgdnxC7D6K0T7vCSuRukjvT5v8uYnn5UGds6+i4ydyCB
mfy86kDdhgsabNhHytpOQxuVvBYtXnQXdhqsEgrcoIdpt1VqYTM3gvpV0ieb+nn2wIsAm0Kbim36
iu5FGqELf7X50Vn57ur5AeUR7MfWk9+mV58yC/794eWvhor0ZD9WpoEyCdpKs06dUxRjkQVfnLBi
RUjdPcTUZsEp4PgTEtOTVgjCM6svy/T0sgTuGVT+8dtGEO3QWZRlxOS6CLNQv21RcP6jEAp0q9y+
r6gpBdIpHHQGs1gzAiji6iOyvLM7MazuRovsZU3HwgkmrQWOQqeihVwwclMuSbtdxLN8+XWR+97Y
2PU7JAyUs63PybCq7ACDcfgKjsbl5muEX3aeUk7qpdk4QJDsjnIHxO8B+bcugKGS9e5XF/0Pkovv
l01AI2/ECQKfci3rpolk1URiSoeadRz1n9OVmUKY/zFmMa8iX9y5fIr4hTn/6WxQt87j2E5T52qn
wh4Lnunxcv890MYkU9cgDJkqyYtN7ET17otUf/aTseO5zKOUbN25+i0J2x5o2aLgsTY3un1bBC3S
4H/HSnK+Z33YMBlXF3E/AKE5lKMR1igpc8pZZESJRzESQW73qFc8+W3JLwhhsOW4UXBVhtvEc1RX
4biqftH++CfIxPFd2VvPVORa8EG7iw8qKjEFYYAnixSYkrvX6FXscvPl2LtiPzpihPfqxANo66I/
hzdwr3VTPkoyug3dZudnIAVU/xShZMlcleDXBVwfTdOGmbJUBenMm1Qa6/5I27c1qjAxweXt0G8X
vKFBJl+NPYSBtClDx1gofmCsaeOMBwNhUmVP6RLBOYm5ormRIIrm1bZbnTeLdBa9wAG7uxpfgZo5
UlHCi6xmnf5zPVm1yAQGIlZvJkxPkH9+WkJT/O/N8eVpQP2PWEaGe0AUe9MCPyxvMTc2yhc2LVUI
YGohF3vIfQS5E0Z2RYH3PYq/AaX08scEW1Y6pNqG/JpVmy/67g2klg1QleF1JZRkXedM0fSvaqb/
swxII3poGFyTU5UGHR+WkwYESi771kJzs/L5nDTiGIA/X/lf1xeeQi9EW7TyLI+MKKBwQ3Rtok/r
7bVfrr9ehYPpqfA0LFJmUGjFnbiMuwS7STLAdA6b5kQUG69a+bxzKC1WXvWC8P2aaEiyupjW/w0C
tQYZ3Si7fiCSN75oRjagdhqy3mGzmjZF2ODadUsTTlDBTiJmFIN8hySrN/2JHQLQni1qLF0ovbqH
Rc37tDweaNy+nx3G80Pk9fYOhqwpqKyXVW5eHFOjs7Cg3oO3s00ire/FpgxHjOriJrgzePiQh8lA
WXcEMakyp8X9TRl6FCI8asWZFFHPhKzB+rG1GPYujWjyRtLbYrXAVkIJwfdJCGn+90oSqHhkLXLZ
I6yRCZF4ZB1oiNX3OODG4DNaVSYifJRQYIgOWJzg1A/6IK/xJbH80/K2KVD2ZHz20pDYPz1VTQy/
0bVEZEyYPqVqCxICQdrCXIvnbdu8Vm3d9I7VUvU7ONJ3zdwvM7UW6n8O4aTZyn09GwefzdK6KUtM
wjDpxb7Ke+lSf5x2W0oka+F2J0sfASPBlHhhglcwywnWRea/u7kzKsKnvifJ6G5iqeqqjVJ3RJHx
KeBv+eJKJygl43wmh1llQhfu0tggueANFUlorahAmcQDNvntKXdmj+sW4epat61lbI+njqus5Cs6
YawBTQu4hpIiDYgEZOojYiaqLw+uNUmkRaXjS7QWmd4K5dfXMB9edPGUBgnLfiicKMKdJ6AlL5dC
wHMHe6M0/ia394V/2EcOHY6pFIUPd6rBBAFZTZzSlkx6TLTwZ8w87bUbNF5xuECighB1fqUNC6jQ
gIQEUO0t+MdGIdkEpsdFQvwmhjStsQyVyJxunU2RtU0/ca391yNLO1E1q7GQpqeDk4SQKTH6pIRk
4IB5b2wECEYVTVq0VFDPSvdX71Q650xZ9HjJJttGlDXv/kDHDEJiL4YsdIffVjqWId/nEF/QZ4MC
4qcL3J9cM3vc1Ad6pFr1xsljqo6P2QE23r+dAKDF0FUNzPn7tnNmNIsofbpdBHkLnXF7cG5odmFC
8lA6agVzLDNnXKnzntIXWFbX1BNMiWR0ut6/ZqqE+ox15nmzUjy7ByXSvM6tvx+rJKrvyt31adWD
/yPVlpSB+qvRcsCeBPI8nV1K/tZmoPPcn04PkB9BF9s+u2WcfG9ALVWIL1zs3zcOqDOmzeVL2O+l
3hjeRIRPrL531j4KaYfT6NjPgDrhEMQgzL3aiqo0VKAKA+KMvoKbeTY2cN/5AiPtiRsLDWacwhDk
Mcfmv1RVd6SeoEdW3P9JCCvusnvLB6RaLTKCTchEt1EqB+1VBzhyzUpwOSfUxxO3EhkfZxll2VtH
KCPoQ1Kp1inCeteUgvdBFaeHgtG7D2s9Ibs1tbs+dhmRz+tglckowVQd/QQrpOjtgj4FVqLerT6T
pvCfNzdmI5j9DFegOotSwbB/2Wrsb70MHrK1enTSxNLlQdyoi0ie72FXC62JmmTxizcdIjPQWcxt
bQVTZCaVHFif8FXzibfAWCpLChxrkf/0WCH9Ut7JmJJVy1EwWeM/3jjhp2XEIwJggYpESRCnb4zn
CJTU461S8x2FF8zyIoIpB5WD+OrW1R57Y+BPmLQQlQiHorLG7nkQrcj/Fmt//F1lzcn9yGb1N8al
oyQxuyc3tA3HiuSUZleW69blSYUeEDXBiB05JO+SXejrXnMpKkrOzTHu9vKl15nVyTajv2I9nhal
EdRoYBgwOUV5dyikGJTP5j0bgwahe56GqKY0HOiYfCl2RG/sLFgWKd9LYFkxtCAsvgmxjHhhr7AV
PQBb5Jyl+7TOQxWHQoc2iaYhom8+cBzHl+vJJF9jP4PbsJkWwB+8YnohKUjdZhfrRZfTxdYwbAk/
UxDlLs2ECmhIrcecyDH1aRjBAkYamk2Q8SuWyT/D2x0SQuSic/ND8o5FFcYxj8GBpQB5Anr/3O5A
P9V/NWoyoYWbL0blcgJxWdg4Pg4cdPLiNmjIk75Cw6lKpxNDkvE1K4kbu5I6PJPdDz+Q41rDIChP
FDR9sGuNurtbVx3EUY89vwwZK7D6DpF9JLNihk0nhd71ZpsbmmFd98WOewlJzbF3eLjdiA7E/DBo
VsPaAFIR84zOaE9Mop7E6koL4q4Wxmj4+LXA2xaGydjzODCYb/p7otauDqUpQv0tBRaVXReu6I9x
owLo4nPkr6P+oVNF72Q5c2GTWksipxjWMbmsGwzp124boghEKtI5ZopkQECAf8lAcpmqR0B8CN9T
5vhicEdJlrrvlG08+uLTMts5caDuj/a2ss42EoLnK4G3qZGhoESgg6FltljYBW4HLM+kXKiYB8Ij
OcKdrLGTmQ7jikOYATzSsVq3xw1e1t0Dc+XvIE6SSfud4edsL4KjhIhYkm01DzCs/38Hsdd5xxb1
TSrW4YPn4r5RK+nKPrVk5lbdknwR+R02zbttDvGOHBxBT9njuxySCx7UIciPUOFvXFNBi1uo7t3l
BAgWMP8EwIdf+lTJHCbMSSkB71UBQBo1Pym1PfnseBP0q8mxMNBMqO5R5HJXof+qoSe8JVDLU6qP
PjzK7CvevW8CsfWQ2M1tMgFpvBxr7xQWTDUcIFyG5xUfnJ7t1oQQJOsCNj1wCr761upP++6MAz2r
mLIppMwRoT+jGm27GRrb8QFQdua4SKCWva1zyhWQNIxLTlsvfvWDVbTxVZVidx0X9SxZp/kDiJct
5Yiy3pFfuKtXMd/Q4Ys5C144eYWyxs7qmknAwOHk0qOFIsSUV26OpPYal77iTX35AX477vWAfdC+
9p4l9U8PTtmnG2/QWBZkybVyamZb4mfhAX+Fsnxq+cxB+f/epGT0+UlzRuvXOWPFhz1ejlKWf84R
TyxiCnM0KrWzTFfj8ZDHTVTL/IsBB20Yedt5oiFhC+RvRZDzW1xizzOHFFJIdGDnewWAtaRr+yfj
+VCMhG8be45MSGLHMettVSWMqmok79kI77KfxbW0xhHFsWkWseO6fk8ew0/m0dRGTMfT6hb4+2/M
w9d3H9omiL356LYierMw7y2XAXcMQfaSAXzt1Pc4PORFIlpdXdIL8F3LtsEnlzorOGAM+NUNuVsC
/UcQP1IsJEOZ8V6vJAFI5Dsd4UUeXDju74d/+AlyeFlDIT15d/AEhXAdsrOIHXNVpvzEXmFmhpTu
mpHLG3kn/bwNWCP357sS7gxzoE+ARsfeRe4NSrkSN67ARAN0fRUMwh7nqcRrHjs19YPVcQqYLBu7
Y7XXQM5l/RwniB/KCwmM6VW7PF452I4LfH+ojhngggXDLyUpeav2Nily7wPGqsFH6UdkQW6TAwUG
c4W5htzImI4q2UDhUIspyQCju2d5Vg8mTvQak5oMMS1UefmmrN8Hmz+s+uW7nlOj1FSadIBwsXdb
BaUqWyqJXnDv4jPtVoNxguwhyyw2GYwyQxYKJZ1Z6jird1WUu5mgFz4UjlQzwFJXdQ4vyMa0f/GY
CLwZkVDhVkt0rp1bZaWqLwSYKyXMcnC0iskUivnQoBWSvQKduNVUxK6m+BIxe6fcjSreAWb9KJFc
z0eQXFIQW4PiilFgj8T+2Fn8Ni5eJQpqNRWoQ5/FJdnaM3YdlyQ70CcgrajbWZLGoKP0vHAwSVBR
E8C2UXCfv+6o/vs2qemGXJaB9GtK0sOXbAz1oxF4mYiFXasOVrraRbv6mV1GyDq4YBCYgU0LN0UJ
SY2O/5ZdVNFwkNKBjE8zpKD9SO+pGBVMlPi0ywVhjK5aacPX7W+9hw4GKBAXmqQxajzK6zTlE+EA
AogMA/IlRslS0Z2CPheXMy13ajodlzCIfhgZ1geTKFgzfUM0jjp1zCedg+Vrc4CzfJYoy8/B7mne
IxbwpW5WftGA3xLW/mGVAaa4KVroQilisKJPVOfzB9SrSLoI0xD18SNKLG9gRdh4rsQRr5ELUK1w
NKzqhh61GOYFmoY/cJo9qgKHVkqGc+W3cVx6wA3Ts0Ld5L9Whej7nUSRJunUENP610857XEnmYmY
SvrrZBAZLlxlf9pLCz9Ye7mQWdIDIJTAuKLAAz3oB7/8qO19ctQysYlwf2BAMUiVWPa1FJY5aX0o
lNvPD8i0YQa5/5Xw5i3dBkiru2FFIlv1ypDBoLmIToQvbNx1/V5k1iB+HKlYMg5rrHPrRj6GlLxW
cULK1CyZuhfKvt6Zs7IlZtSXZ8qk6UD9JCZ8//xLJ1HswCTomdSTdQ/ZUQCSTPhTsEy4BP+TNJ2T
8cMGtPCmD7ePRgHNqfNNUdkcm22wkvWwmLKfa88h+t3ez82nHfb+iY2628lZgZbQTBSy+0zZlVru
GGCt/FKELmpSdnu/igLj1+4kjF+7lIRYRu9W2uGdfqv7GO+VNpFVJ2HUwv71g1Fd5txzGHek2DwC
kErpXfHJKIB6OLhd71uQri/RnPRA/3FF5z21fihcxEqPrMiVIC4NGMa+byQETJaZhn45cCtorH+3
Oj8HEXmLCKGvo9Qw0V0AipQ1JMsypXeUS5T/sJigShWLrBPB55Z/EDnTaGNqWz+KaIIRHxTQatlj
GVVh8XFuShgsE1gdXH5Mqf0yLLOusLq/1kd+mggWFBxgTep/bYWiEhJJoyUWg037n9IsVa7LRudr
P9Tq1xL6I9ucR2KyTOQ14i5lpN+5oFWnKBSVN6izsGZQXBcOgiXE5796/KmxbrPE2Qwp+0GBs0J6
nYtXK0kpCB1f+kpmN5rMMe42oYyEwuIwdmRMLcvxV+dv0xsRllaDjW5fxTCWUYa+joeCTF8SUyG3
eks3In2VTNqTC3DSfLa7cU85Zpg2+MUTpAN2pNnVwk1SOEFmwb5dbfOjsyJHBhv4nY1ctYsmD+yu
XITntwCz8lBLldKy1ZyORK6jCC1CISiVjnh3sr4EYz2rpeSkCMEHEJ4EuOozUAQbbxXgd0zhiGOL
yVUmYHKJU5luYi526io87dHTeYpPk38pQ3YS2d9QYJc3k/87/qqM2e1I16QO9/XFn+TyUMgtN8pX
Ul9j631NmPhBltN+ov2Ev8FtzsbcShs51B0ull5HzLhoeBv7eaMr/JJoLbtQe6CAfcvotkGW0QK7
679L/UQp7/d5d7FlG8aJR0wEDYJzIIzqTReVWI+RUkrRq3tSHXC6+D2OnDekmcZGSqrjT9RV3R6O
0pS8+vL67un7Z3l/h0I+6Tt8da5boHtQfMXB6cA6GGmPdzhpp51reKCIfq8YtA0Fe5X+M9aTRJrL
6SBpgeYJSoGSgC2XX9/8+uvpWmSfIPt6ork8r6CPoVIs7bYY2OhyEXlxKcX7RF+sPZh/ui2DL9Ew
LnV1roHIuGcAUBvLaJA14zTM0qFQFrYuzh4u3GlFJue48q04kZgKlUJLHcD0pFyphDjstJVo/Jjy
mvSxzISGnu+hdBl2BHUoYub4r+4Sxqi8Sz9x2cG25gtFw28yWYge3fK6b9fqypEqvI+BCpDwWEmT
COrxXvt+2+W/z9ynyIJNyIJ84yhdHz4hiZQYyymBmObmB3p4vCsoDzcTKFs/+wc9qbjtVYluw+5I
xwVDuQq8MohE5C8Ypa+4qEFOr9QhgD5rs0UbSthRynj3IEc96RgwIdF/nWKH3yedpaccPSciwQmG
jUBaeXTdhQVH++IyObhsa5QjLOhiC3aS7DraCdp1ualOwT2h9+mnXbOcnHAYhP7K7qJD/i74VUoA
oUj6vQondmAxUO1bLXjNxMIcHAHvGHlJDnQSAzDe9KGyGAu5CVsJQvb0r7pq7omeNoLXGOxwJjep
LbulOxdnsDvP8Rqp7qh5iufTAce70edVIo0VV5KKHEIyqZqKMpIsOxM52x9KN/SS3OlzZwUW3uHf
2guar2aQb06imtaTs4xDkqRN2TnLSrD3RwZDtwflnwXCicHOgrAVunbR65B7uT875fc/HCwxuaXv
JddoZ5A88QuXEL47tW9wsUBQBFDhd8hwVol+8iJ/xOkz/GoucxbH8FxVLzmwAy5Qqhc6GomEty+g
jtS5G50/MlSNZG3dGmrNsPtNTkfZ8UE/9tbSHMmtRmYge5W9+XrvhoYXGgYwqPzT7RveZL5vmMuf
Qr3VbFcQoz13TQ67ovgHYTO699yY4GAVsDMnE4u+1eFexHT5UIVZYKlt9+EbHvw/MMCrpz6jztL7
oG13BfepevpGaUrE92xA7Pjw96sl8ORP1bLUfruwfLat09bbEaFS+Y927i+ZY8uf5wShxiy2SGT+
A8dvTycq4zmqQw9OU9qPxbmsh7gVS1iHf7uB19G3RD1dKWPvmvGZoBgZsZiiyXqaCNJmHjM8EMNF
hWoDBvhYuI5MROmQzUQ4M/Bl2FZwmrnIYmSn8JWmUJI9hMcb8VHbWU14mTL6dDbzUklpdIF43zbX
+eFsb4ndu5JO2DXZ/SbJXk0hNjw/6muUBH80cKNcLIdqwDjpRv1cdKQBhZvKA000wfg9gYNbJoLP
HGAnktGyzndkMtwShkc/qrfyNPJCVayzIY0uJ3jKY9aVjFnR27JCp3wiV0MdFj7g3BW+vKkb2wTf
/lA+aPl8VB7d1QQKDc4o6vswcKKxxtCABxzJ7J1JnywJpD4g3YMOIP614m2T7vow9bYW7DdsPlZ2
/STQtzpoMoyYxhUo7c8RjGr7xWPYq+mquIjjZcFUKRzyBdsYa33g9oReFehsmw+3k7xzi3dBF8AU
iLoB0bDW1r2o8Qxh3oaOOOsl+/BkGOW3ig5W1FHCn5CJ3wn/LnnsAvEUcM1wswvBnuAhubLS90K1
FRYvqxeTSzoHbzcCKjIsDyClPLwisB7pIaCq7AWqYEAnabVLd6CP2sh0qjlZqwTal5/YKC5Maf6x
odh00FJ1Fu2i0Y5EmttjTbgKwp5yifdtpAh+iR6QtgaAHXlNudUOt4Ln5tq3XL4C1eDgwvNakTfK
W2fhWTVRQhKywoY5SMXI5UZHaeQL45/Zv/JqRAhixHoOlIE5wIskAL6C16gQqa55lvBYJWZ8dCzU
YKjtPXy8wvFpsgG1JP4J25CX6sNUimumJNXFdzhXY3xZQaYHsg7Q+gEMdDCo7pFG90gBv7AMrEk0
y7CUOUM/m5NjjKyTVWlkc65rfgr4ETC+k3OQACuaAXzzGpjaO6fcoBjWZ0E0rihHP936apNDZMTs
OAgWlqhDpZSpOjn2Sifb+gZWBhUDYy6RiWikS9dhkjJZcrcEdrAyk+5JGxaqZV/YqiwrjKgs0GCx
YUPU6oVUTx7Al2+YSkiASJML3JQM5PegMp/7W3aTLPh6XUzmfJCjwp7Jpyqt9kyVRxCMqk9JzTkJ
rHoF95dYv/ijHUFzRkdoJr5JFJk5dIIXCOktii/d+H/y8FWVt9JSvuX6qbFiGuaO4FT4DmyFFuaY
aUuIXmHr8DHwWZj3HGt2JuB8JaVHZX4Tmxhf/tfbbbRoUdAm91ectQbdFcmPaDIqKKwVlkWCmJXJ
JpbkoztmkdcwdyEJl6F6Irw25s9EWTsSjPSIi5XwSRrltagIslKCns6lgstXe8805rSp8M9NnD1W
2K+6O3qKjDV7gGL7FDQ7TyXStYoKiiMRbvpvMd5FurWqZ+BJITCVUH+U9170Mx6UHfXaC8v75CsW
Ixe2wuOnWrgy4+01OTqPQbX2At2g+a38XJ2p4/VVPgxoG9Jta4L9NN/VMbLN3jb36N5KNN0KsXc0
opQWgR2KfTCWW0qNj+4nFR57Whh2WGOSnfboJzT7RLZ28CeLNX0WqrzYdkOqh0yclR3ABgjRFh5R
SJuNkwPDGzT2SeYsaNrPGwQvjSdCqkSIOmDVkgdQgJIZqqHmBxKExaL9vCtk5DEzkO1jKM0eDa2H
O5Wth2JFtM7hbwM1Mgdcj5I2m7/2gi0gDVOQUcKmAPujLvIi2YGvjJh3vpjApnVGRhCPJDmKLCrx
EchG0LFJGBRLU6jjSxJVgiIjyk9Rg5nH4UJuGoiPZUe9oZJ3p+pCh1Q2yGRgBZVWX35/2l5AW6P9
4lNkEiA1a6euHgcfHn6YqIXRX/RqOHIQGEPWubexMNdrs4A3kJEcG+I208gkWk/nmU/dgBvlWGzI
gtGG66B+bMIBxDrmBzciyYNX1TLwamgorTfTz21/Wpqw88isWf9DMsym33EBE8AEWGpaVA54XO/G
wys34bv5lmCALNNDSYJ4IvOEHNO05Dc6loC9OhKv9OcsFVXCn11GgcAvQx9GkBdtFUvfUHhU6M7F
GBtOT4B3DEDaImHdv66M2CkKEIRajJ+aG/R7NHA79LbsRZs+palV87nOJV54WU3LOeA61rLaYJcK
Ob/DycSwBxByQGRqshYjGrTQ8O0274qV6ngAK4Da5o5wrC7RNJ9u0/vjky0+r5VkDd19fAeVN26M
PkkolQhgOpHRcOuTI9OkukQDQ8KYZz8xPnyUEVtK4zpzjjIKZ02xTQVFoYcuXD22lgPLYd/ANmnH
TAf1mN/Q0zu3HLOz//El7Rs3vqtn+Ggfa4gO0/jfIcmlHjzk9J5C2kFKESWhEYYO9ZyFCpAeyv6T
M37QKyu2+uMpZN9wcLA+DVGQkqwvL41IMKgAipsq5JqS0uP09vkoL8uEG0a9Uek/5mcE8B05wYuJ
3w3kYZ/x1oNNd7TTix8d/sLQKJ7150By97YMMJGD9Yo79Ubn/doL+kx7JpGhDtDzFpunGxes8yCW
78kEqvPU+xR0A8lBOpc+t0yMIJPodUYZAc936BHDC9hOseftTSKq4xvAR8qRVYeB4W8pGir6cvQR
y7SJIsS3AEhD5IU5HmJx8FiKnxnaF5UK33Vn6h4JcuLpKeDUKnn5hxOAeGooMiK563/cqBL2WjnP
6+IiyRYFGlONWPvEWIbUnwL+pealfxPRhi69EfhSCzPFEURczb+4/M43FEbHicSSbTbafGo0gLwO
uMMvbV8oyfg7Nn+YN5JD3WVkeMMM3jK1y2i6ppztXwNt2RR8UcCaU08bU2F2KiHH7QuAy1FEMiX5
ZVWTsF+nDwRTGkGDOgfvRQwfKNBSMD2zY4eYG4+Az63ke6cLso4NAXXrzFdYJuxUA4I5qiLqcvxw
RyWx30nSLbEwlSI6OqKAjOBTqJ3dCqviV7TDmzgJmgnDf6K62e790HCffg1W5+6BjYemRUMvzY2n
T9aF1b3YgvpcjKc8rMzmEvrcHgoVQHz5l0GrwJ9D657orREHp64S14jse+A1YxjtypWazbQDDLf8
l76mKyZriqMzaFnIR2187fIFKEkAVHcpOUf8izbPIvILMWPQGuB36dnhABrqgPa+xjKX4LMag7Fk
qBL+CZbu/QxJOHCyiTSiXhdeelWNcw2PZbGK8kY8++8o/mL4d5GfKxq3BaGb9moa+VsrA6qg6cRP
J13HrZuRULAnVTJqeoMBQzP2xKK7tdD1WuplrPKmD8CP1n50HExkhumeyxK1NB54GlOt47huGvE9
j2ElgDlUwGUBKTk89zWO1GZ8r6KSD9QADBYfbA/TysPwnYq5LIOjIkHwDX9PdGlUd51wWFsPRN+X
g+8IA44NqDu9PUVYH93XVEbiJPmU0QtzEl4UClrGlLK/wyJ53AOmt0SiENeuitFQkFu+oJk1Ailz
mNcKsVaB8OuWteCUPSHkBfwdo4WhqJ1fUTnUkD9sTo/9RA/JIJlEI88t+zmdxXjcpuVz0nWCzPHW
wvusxdc+XkD2wRv3hV8K05t2rEMyRT2waBElRGmUMgabSl6B+JsAEFz35EMx7ylLi2i/3Dy76cpz
vbdpTiGdsBl3r1t2Osb6yhdZuJ3QzCIoR5OUTOkuCEE1AdnRLILummvigx/gXxHjOLpbME9hB6oQ
8S0yI1DR6jv/O2w9T+Dnwnnc4BVTbvOUdjhBpVZYI0+KvWT1JFUA1b6e+rY2ziWReSVMkr0L5pj6
ZwLjdHehLAWdSzo3rxaFCx6r63ADyOZWThK/u2i0NRmPJ2zkGWK/ucMq7f92YLR0WIHwJ6+C/Xa3
qCXMpB+nbR9w5VR5pfyAuayM3j5sYOKdFBNnZaej3nw3rGCd9GaGaU0j96K5ZPI5/ax5dzZHgLCG
CDXqnB7l+iFKQUCY5s3UMgxNUWlkvWOc3qtfuRcYmSw6KByGa+AtqTKav6jW+Z1zWoNQZLmJFYrR
qsUrJP4SqynjTEANd47zrxnvU9okUhHrG4sUQOoJwM9wv6E+C8HbzlOLVfV0Fyjmx0a721WXFowc
mBaSpn1jSr6IQsoO1h0NIrp4aoqIJcEiJdhSJaGHhzvE6oSsSErfiHSJUYV2GcRazfjznAmHc1Dr
5I/ApJBKXQFZZ79j44i0TmAU0O57m0G4VBy89+0fjI9V0+O1ETiZPxrX1/H9YGZDojimFJtGg944
jP8JP9yBsUprNGiqaSIkeMVLpvPSVGRrqv65OQrY8N6aFI+ChiOlf5KDCllzip6cX4ruhVz9bwVa
h/QgT68YmDU1a4UGzfx2upg15D2YbPYJqxm30nQn3q8Go6AmBqfXCvonyzu86BYGH6Yls8S/Mipk
/MkTTc2eC099l5rnpTNLlg1PjzwK4DnM3NCJ3EGjxBPLfDvuW5WeQwkuFMOkkqUGymC8IPCo/7jV
5tVoKQRTUTG3DMmS00iitUq9qvwI8mpIgOjAR2615rI/6PxgISWmnrcRaAy/tIZm9rpEUqyClVyM
TzimIDw//J1b6RVbaruMf0KbbMVAuRJTiarbf+jbubjoItT+NYeSQ3k1dss2Y1AQ2qcor4IVOcGh
vDXLwV9d39xPVWOQ6Icdaq3U5p2pibt8tK6u/Rp8t71WrYSCA2S117GtXZ5S4dqUDDtvyh5hf8SU
0zjxSZEdJLCRjILN15evC002stKJaEWB2HHKAfea1F0fWOFtYAuvpzaLtCNHuEtNCTb9YBgj9f6p
yddw66OKPOz365E5CrZGizOyqr+4CSA+bW9lM9cL3AOwv96Hfo9Sy2sYbW53orVD3bM/hfAm/3t7
wQ8pUzozm/Fq9M6ZWeRNh0n3ieIYQnoNVGJMBdD/QGTy4IpY3cE5gdH9t6Wjt73ccA4eSKswGqxW
9GgZ7Lv5PTSFGociGT0ws3geiQUnTe4YwkAEb0n0xoP677BOt/Vst/79QMsc0nEjf5ax/e7Or0i/
XIpJhSv+XquFRMKfYfXPA8KJh1hjipnm3FJe3IdeZcMvI6reT1WYmCtLuIg49n3/WLS5IQzuXgKs
2CfJOALEIRSTKfl1tpvPyAE046p2Ht05a59gO+3Ejn7rXNUOX02HgenMWXEfwBtz1ycIxok/u7vD
lfhI+u9bqcih1FNXd3PLLrz/wjIc0ljL730zkhHWYtPYZTEO5y4QrGKWvesz95kDvdqNMaIzIKNF
H2ADBS93UVAY8YQ/CBEqfEevYd7d8NpxQP092XFR6R05cLwKodsjdWwEZ4a81l7Z5AviLfLvN5Jl
FZZF8kgkYfdDKWIS+e2UmFZPYDYCBhyGYX6vnFRqpEqXhT4aE434Zb/ipmzhwI5sd1wVP7zjv0K5
+ywm7uRdWYirkyiz51nqCKkFwNctSxjk0BeLcUOjkCyDIgcETzGybc4LsYxR7fVUqalSjH//REpt
ARDvgZh6RkFBwJHIBYpaBbSsVs/+0l7pazYUEgkqS4IySQiFUTSPVnFiSAZFhcEh7CWifrZ5Bj1s
iF1aPPAmJT7XDRBhlkK1AKIPsFsT8hFoHagoQfNowvOpGmPLXrMPoSxa4B7WHZc/YPl08vmOp6vG
fMW3wufk9LImkAnxCnPCg6A6IdYnU6WvGmTh7EfDryoBaOzJUuj+4F4PpE/+PetmjWTvEOZhIZm+
DYOfpaGyPrdUSWhirD+r4vXtdmpZcQsiXD8N9YrUXROL2HgkgMpt7Vhjf5DxAF6m5nB3OzzEIiIs
JhFxpPTiwoZdcL6Sxk/6iVj5HxMGu/1B9jiJQ82zdJuoaQgCISQXXKdkrFS2qR7YecY/pwaV8vwz
jaa2MEYD8VvjAQBLwdU6zDNahekVV4zuRU2dzLEoLw9SWsYL0jTf70Wd1GHGZs2oMqXUcBe+VtwY
wlkqj2nq4Rpv9e6N3d6FIzvY6PoZC7f0nNpsID0XvFsEW1GZDbt6Q37ebjStTU+Sc4FBC9QbT00j
JNQYzj8jEvUgbyt4o+GMd/Tmf6YBZLeNxLfpUs5uwWXrnurc3ZFgimYmPZixW9YsqQqN/KjXSCgG
4wRzYype4im9loWHl7l6U5e5aMo2IlodwgYRVm5CtPnzEl2diZlOevb3smj3altGZJjn+haeDMsA
tnhNQxd/guZmEbvix89AerQIZnA/91kHs6MPea9SyS5zC1tdkaB2fWu4jo4z5RwLP/IC0HsNGXbB
8cK1O+DstD2mbRo7k1u28S2OEO7fr+DsupnImhfx8aqoqhfthQ0XZ6IRwVXXz3hOK7fZOWItcIbW
fSezzIhDETBHIO+gBeLZm6Suzvr5aXqb55jpIzgvPhZxfYIn9imevOt6CVbpXApGfvZsF4jhlOIH
tMNOXG1+PP2PhreKyWv5PtTGuLa/jpW4eeEDphZGQ2SXZNjriVFQK0uX0OKuuWsSoHywpe6UfsSY
p45DMVc/T/XL/+Q9tw4GwNKGjKkrGKzxTNFyRM7ykL2rVj/z7WAWBL3vfwuBJt3PttnnUa/zWmHR
jFlSwWPYl9xZDEbyfswhJwflLsrfbx6LjW/IWBAGJG1ZWms1TUOP1Q+rFKcVcMIlivAI+gLl1IHP
CM854Ho/B8nJez2NkJxPB06jCMhjE2qTRORjQPzu8D/QtfkAZUk/G87iwETTlbSmS+CicgfeGNfh
Z8GDXqyy0jmgg9doDEsm959mONavG1vZGD9/iRloeBrOEXyov8/v5wN1YM6Xlm5CmleJ+z+d4TuK
PJsLbkpTb0kAhySB65g5f2biuHkjySZHUcpT9GucpXQ7pZLg1MltpWmoTdCCtHaoelcvqhsSP2Yv
Hj7IroHHnmPGEBCiU2R0clhPmJ0eiP+vZYuOY+ayTKAMQRjVx/EeNCPsgZfpwZ6NB/MFCoPhoFYS
2gZzmru9YjOgHyYg+4pwjA4Rcp8o1tEakheTQ2vixc0cVfl1wD56XzM4nKZO0RbxtdEpfa2kO040
ZOWqPb1CrSFk+YvtbRRnKLQCaSimYxghrSV+K2E7QDKBRdZdmsZso/+O+NZ8wooTRznG6aI2rKSz
nqsjWTcp++d+xq1AOjhdPELLCw4Xo9T8Zk1JXIbX2wsMpU3e2Hyjqppu/EnAES/+q8RDcwoVK7rw
v6fVYY9sesQVcnCVB53YGc36QCdCp6AWCPESSH1Fnr3WHpU2Nai351frUe/NF/7fjpc6l/DLarDv
MUu+r4AWDniQDmOLbKdDbaV6z/87PFZxU5tVklHLBmVfLk04+mZoSBiu74xzXUTJg78Wv1QqCJC7
vfw9S0NG/ijznPJ0mu5TVHr7L2TIX6MImHb1HnwOodBIqs4OGjOXFGz8Elxz/ANFbmn9JxaOAYoi
yT/P74zEc0hGDeR+YYd4LGukVYlMb7YNJhr6bGMIXdexx82DQDftWS1pH0yx9sk7h2Mitjj117aC
Pc5KvDfcOXGNOcxX62BgwtXA64XPF2Amzr5kPjeGC0AUKvwvPUgmhTthkE2T/WJLv/WHDCBiqP5u
+yQJo680dPiUMn5bVbsTDea8nh9Dz3NMQK0cZaExnXcc6nDHHX2gYrWCK87ToP/r4Rpg7Kcdnh7a
+dhZ1XqzFHQwJAqvMBSoHX5LnZlqPLf15WViZ6io4qwdPunyvcGnAHLmX2U7jVMrDwRwB0rEvtT2
QEYhdlGt7i5ltskhkIRKlZ0h0BInsTVlbAevu/XNrEfDxW7ySUzYS6yjcC8YHKDzYhfaUsIk58Fu
Kv6sKBRxJs9k2+Hv6P/rFC1K7Yfl2tX2qOHC/SQp6+dfwLn+HswRvqJyuD11gYbD1Is5vLsodJYk
cldT9meZ1ZjnQKEu4sas9pDf1iF6OF+U1jgrdzqWRRqjvJtquzbOIEchzm9g05yNKdK8eqsqSjmv
qkuhmFRAx4rS/0vx6G4prsnv1HSzY6wiKnroE3tmqqFityiyrlHo74G4AfDxPE4jgr/3zqX6+zNF
ASFPE6gGaQTofmZFjXXMTFFcoTk/PQgtW6F2pKL1V31VDsrck2m82Ax5P7QIMhSk8z39d8DWg1yr
OD6s3hHENSuV+OeEYBOHKMgOI9Xp1ud4sM5iHaopmHFk45EhvBI54v5rzeSo0qk9Xh/G+4BCPfpC
WFHqZjOrG11cHOcqkwRamx86qG8JF/7nhMsTU+/249JEGHcDz4OngEVAzTa3l/cNDpbmLw7DzG9d
8ZytWeVyu3fPpiWvDYnvhdXqtzPdYkl0Wtq10tip0WgO0BFE5CS/vNpcO7/oJICDGsLT0nzaaLkW
HSRrOT9UdVPVVqQfG2mySnClgMmkv/jBjY3U34Esnj9RJd5aUVqwarLsQvE4mhYZA9PbWZjAqo8W
wUqHTSyHMrY7qkHB/Tncjhj0ejqNAF1EhBXdP3b38JgNTKpNX+rL2AkmANh7Av2gs6xw7w5rXYiJ
MaB2ZDWg+xiQvG/ENXju/Sa36z/x9ilEu9kzZ/gydPpc0T1+poUhRZqz5fQ0fcMzCttDWUeNX+Wz
/WZIMp68E2b9t7kwpdpFmYc0I3N+/rXLcB67c94NAYPjczJt1N/c4IIkYdTd4LETAE2QIlodchRJ
opuedKyEXSZeJA3l8HEFN1DwjLWI0gZ/Y+WwqyrzouwWEWzhF4u1M4XUxI9nHoYkDKq4zwluo00K
lKSGB4io5cZTeIrtOq3oNzgsU/qgTx2RQJeeW1vzx1sH8TUL64R3AnKLNubK53RLJML1tX4R1kBe
W4fjLe9I+sChJkzvw+njfqnzYD4gZsn1ne3D2MiS+5v/5/lTCExCriNwySJThlXzraAnTie1nZXE
BRKDZUj/aYT2BzLVvNjS2d807c9eWPwXsNLVC4LencdbCvupCMeNesysiHGkmCWwItQtCLU4w5Zq
8wmizdaWi/isShsVUShCAX1Z5CcxBA3af9h7c6uiNLsZ8pfEZbJsiusEg4EeFHHrozvKpv7t3sUu
qpAjvyzy8lnzyMWZqbn5+EQeOnoEhN8Bqtdia/E8Ywz6mQOIW61JkLJ8ZVKbqLL3p2K923S/RxA7
bIitICWEWVvHwxKS5wxMQZdoD2gDPJJt2p9gVWY5cr3L449xACgFyOfnIZkjm63RSOOKHtv77XF/
i1iECi9AcNxgA10p1AiXV4XMC3auqvgFuXofntZAcs+J42zGeju/w0Q4cRpCAyAFKgUG/NTKcWo+
WUflmq/IbLekVQmMED3HwCS2mWKJQ82i50Nw41vbywAt0IdMq0erRk41he+zdTEMAKIm/tpya/ia
7LlAkqFTlOh0k16F55FWZljjmqXgB/ae/AAF08VbT7N6+ge8NYZYGXphgz7kZGKGAGGUm8MHeaet
jeDtqpkCPJ9SdNRxZM1z9+6d2TamX5Go+8EHBfAOwgMqvrtROWrhcXm/scHI7oHBJRImUCWgJCDT
cV0zFWcuKfhNqj0sipAy7U+7ICABBoTD1iLtu0YzFU3ivUhFh+CPb8t3GqD7ZhYVvOoC8SGD4uzF
yG6GBhVA73Acb59qzJbtQarLQDyZPeFG/qaO0QehJK0Cnr0YGNxo62E/xwCfxi252e2uRPckTZci
dIDkCa3/t5/MNxryj/mPTZkg0JSyz1VHtVj9ikYGlOvfLVPwQOs6zdHcSkwjH9GpbgpF7jb+2Jo8
8GaRxk9yUBszqHhWfpW9UrVMSzXihs8vUMexhpsfexxdlhoFi9QZFhxX4+kaq9w8moqZcxEOnOCy
BbQIOeesHaeHyqRWr6RBSYEff3pBoUy3tt0MeoSeqbFEcIev9zoP0XoZM8XCRZ6HzEb3THMC1RtQ
jthXhL2Lll0PI9UKoXSfvZa68KvLeA9RipqCF+9jZH+DPd4HQ276TgVWMt9AIq7ECmX1YsEZ7y7Y
eb4Rg2igXHD+N5bDJgMGJg262fBsSrCExomL9I28zvM7CJEBhfbHLD/8dTDvXfJf6430GBu1ItLL
VMq9zxuCY48d3T+euGOCtQTVxK70fQBad0GbdXeAL/JhGQxzLCl1Z6XzJSrtoOhyz87Qlc8EPyEy
CgMMka4m97/POn7GrTnHKYcxzh6B3wcYqiMq3+LjR768Y7iksJcCWHL9waZ0Wvhgs1hTaBUDLv2A
HbVG26NQ99amgul42fp+T0v+hXTwbGs7wFr2RAcezMAwDWIrlkfegOlV/XAZvwo/9MBP4gXe9Wks
IBj2Ux4YRiSgPfYDpNsK6x0dEEo12O995i3bBgOM4yWCjy+vU2PO7RPhR0YZSwkbKCQfqdcg/qIx
MMqDEiJRv5COgRwM6C6PkAV/w8+O9lk1N1/yJIYIzkA1pOcpVp6SrE0kCT1rNLJS0ftUWc12Fvjl
Xv0aOLDf938PT6Pfg1M4ZCFt1Uvpehhu64Eo66+HWW0Lih2jqSbmV6nmE/Uyzvi2DQOKIjPOT5ci
6kRpI0hCnIEW54UhFL6czy+k7zAsMFnPhzLG1YjY3XeGMQOQdlQ9fJtjcvwXojaIfuLSyUhCTxON
XhXJzWBVQpYHlvRfNr1qV1Mq9268NG4y4/096VD3A+M9MKLkZwbI7gGw2kBYy0cq3F5ALPFDtS2B
yL7WIjVxpFMl8UeTct2icMq1z8hQ1UXo6cYPiW0aLXzilBUdawAHoAW5FTDbBVFdaZdSjH7VVLrh
NDbzGcIvOwk4FzWVVBxMSvmiuLpwWBdKNEms7oVY62FjXHeMFs8E3r5wUH2bPWokW3N9pgUm3tNO
azgXvTFoic3UUFVcAPBnToreL69z3+M9Q5jyT0k1Ov94gYhN9E0FPfmW/4traBWqhPThpnVYZvcD
q0TGv+Dxkqi4IsUCbpm9o+b4ifQL2c+w0MmKWLyd4f+7Nw0x9EDD8qHdkKDzJuVP18GAmfWIH+ot
ILy5xxPvHAU9nSwVqARo1JCDZhHRok29tVlE/VAPABXj7AcIP+vuwuEI4N++WV9Mp/E4KjXLky7n
Lm05KL3B4s04ENGlqwADYwQ934UBjOkZvzZIyO7Yv05V1sqxn4A02n32h1BiNzzJb3EOWcORTOAD
JaHaWcEw6+ZZveAHi9O/txmnXeNnfiza80ZBOxZk/Ictk0CDg/GQ+6grTqpq7K3VzALnL0BOhMyv
/SGq9x7o4OWBQnhYnQ/ldeVRBkYyeOSpvwTDZ7sUh1D5o8GoVIeLTMzTXqX4B+FygcgfG1pCSEv7
3QXh6CFCFpMTk7kLQaQRIUamCxHlrOTIoHOc5R0rfuO6DqQI4ITw5vquKmYgYV4l39l5/rw5rdIm
/ZG6P5tTTG28p5fkiQG5WKnq1jgUIQ7WtAaUJ7VPmegft1NKtNoT3zyLPNAyP5hzZ13LHOixYi+Z
H3rpUe9LgQPU8XpPAAcNtOL87fCKFmXSxNjGUOcktjIcrtbpm832HNAfqXoyMlKSweQtWQJ2bRYj
Un/TzAxdxcd8uOBeGF94HiCU+JOfHE53JZ5yzljHvizWot0gNuqcwvbi3STKrdn3lOSF4ZMG0w71
45oF8+L69vYUyaCwTKGFzoK0awtPbqMUypOByy0kj5jJos9ox7Wg5FM7ahfcS9PYH5wYR9l67ZJw
nPtjmwTiKQihmO58L679dxh4jNkTfasHfdTkNbqXJ2vcyWaAQguRN4Ye4bI+iXwix7I+72R7i4KV
mgm57LNwPQT3nd3tfkYMA6gmqrnAVV9308eW6so2GzKIJ16i5n5izjP6KNDgwbAS5yBcww3PWfQd
ZlyhEU71/o8azEsr6BhXF02p/wWY8z5VM95mVo56lYxoMnFOdCQW3BaopxXSQuzv90sJbjBlBMzV
K5F14MTplTJGscOWZX7BHUJKRdFQBeJ4ZBrmNopqG4xrqoVguNMgkurMn1gL5BAziu2g772wmCE9
Q4jIwBwqlWTCwRUpWL4u7zqZd9Sd2MAZubSK12TVd12J1ebnznOGUWjipTfj6kZF4ONk9R/WW4hR
ebJRgEeJ+fOmSLC17SUyGIw1fMPGy4MyPWcn74SSEDDpD/sBFL2NuOoQXm90Szd8I20DTyyxxCIT
k2ueslcZQANuH5YRATQlmZZxB7uRUqPULoasrJAEyvgDVhVSiBs8tBDaSXx9SUCVZiu5lL9IbhKm
pPeQP6V7+4ZgD81d8m8fYQsyd5n1eF5g4JqwEAV+JlD62gUwahM/QGXmPEA07X7J9h8wITOOVfA9
bQ9tdm02uGXDWrRVAQqUsJ8pDXu6j8Om0YHProXp8yc+jNoJ07Ez6krvLxsDUnYKNqqhNEgouxBt
lgBzTkTW+9OFETJA4QciGqPhiawe0+5Lg9sADdDcewbZ8U3X8X8Q+KSa1GtxbP1LWh1sYEtYOrcc
QpHZfAvvwZE02p+VP8i2hcKtFwl5PubC+jydjQOHTDVvj8HBZfeGteHAw0qVjoYDKEQ07eIxouJ+
R1bklx272fVU5vgbOtdCybH7BEcI/jun4TztQJRZn6G3pW0hOJMhW/mlDrvxAS9OLmdkcYZp0OvL
DeSQFGKxFlZ/ONVZunMGaPGPi9B19FyxFfiYDXJMtODWBySLT9i1E2kfKHkH7JnEVHhu5aXYl3Xw
18nkANgBfJIwnQSosHj2jhUldD2ugCsmSXjrNGwmH+eV7qyL8HCcDLFaY8w5TBI6i+buU4ZmGiF9
TkTXwDPJndOYALVoGyR30KklTRn5ui3mT9Fdp0+kMpLhmcywWwwEEzsFM8ovGUGBG3HzhVqHzp+E
tmfqZcIKUYV0DC0eYS4gXm2ELwJJ0p/vDbepg8xgtVc7NRiSwEBIG4ZvIT/Gn+KqUX3NUEWAX6h4
fGnz/9fsowMkoz3ijtAHEfCsWMMaYfsnIdsxcX8LImAJxKn4XGBgHkJK1lvcgc1JX+LgP9ZmusbO
QqfJee8b8UYqZVgYaU+AJ5sMCpvrfQ+LGzSrP+jIIJ1vpvhX5SryY6bAcZfEnomay89a0qGhjfZ5
ugmlWHqS/b8hBVbd/uHULGnwgjweCX3zPv7vY1Xaar+iXnijqx7vig3xGH2CJ5xC+AmiVX1NwOCZ
7Nd/g/5KMtP2Hiik0YVMyiVIrDdTQRc2XdjUv/NVmjILQ8+2Bthq1TMK1YJzqJd/k2B84I1g5e9R
VKguQkySRwmhEZC29SBK78og2OcgaPZ7pl6N3hTzetRsBIVx1I9M+WWi5+AmPAKZBfMJfHShBRv2
YIBFO0Du3p2pglnkPVDQGwrXjjqMeDwb3aJ1cDNFWWH7mM1xgy4zo5SfFySfJ+9/oWbVAftzq4lT
poQamIIjMHbBicoL7dl9jFsMxr8cyn2Wlf4caq1MFoFweEtw4k9Yer0pNDjG26mTmDDTsVnj/i1Z
VMSfqeycofYlzG77yEaDKtIFSEK7tLEf6UEYQ3Dz1RUIT5l2+ce74FV2dZg9jwP4OZ63xof5afVO
mS2MrINZUTsr17+wPtp4N19TMHxZbk7h/xWRWbv5D7Jm17MHcO8qAehmK9xPet6x/gyiW4R2orev
wl6DVa2iy3j3hvG9y6BcYr4nW7k1j2khk9+XiYYEENXpk98DL0Z189YrBeYY1gG1/QW0ZvSPmfdT
tfv+gtyCTR8WBX6Vy79dONdK6OJAfGl34M+XQ/o1EqSq5vWbjJSCZCgVi53ovlaRv2r9wRpWHsRn
oyqcjbHb0mg2Mv/XXOZSYs2m2sOSLCvvFcr9dTsgDTTqgyLp+BIhH48jxVkrK+YKobNN67f7qjj/
gW3m7mXSyGOSGztuLLLpdjuyvxn+CufVH2aAxH+5jUWrTUtyn//1e/eDZfOeh2OJeXSbcgMaFUFr
ft3bpQ4ndEEVDSnCR69dAQH3Kw+9p0tq92xeErNAHccCVwuuM6IGcPWmMoEEenIQVsuMwUwBiCda
sQPpmGaVmrQ6hCjeDm9Mp4MMhwCEU/rU2a44jjRoL9cBoU11bvWw6t/ov1ryzC7atZNQVw4ETzER
nxyC+mprzROzSZDkhmCg+dVF58Vw4azsXGG0tZVkeY+y7OprEJ+gwrTteL5BoRUqxmBG3lDk0bqd
D2UwKH3Hkh/YSZaCrOq+E/T4r17yYuTgpnKATg7sjB7LjdSLZNvxuIlalBidiBmg5XQ6rvlYBi8R
KeQdxlXt5isbTFpVc685P4f0UAn6on4ia00vhYoQKJTUTUvtjoagfctpOAKGkYDqYJPSPdE5Jglx
IDfC6Zc4l3xTdv+JxWOx/r81zOEJMRAgeD9MwXdObbfmVvggDTKAJJKisVh/x2oURRzIzkMjy2Eo
5/tyIoTJ1ZqRsrqS+eM8RYpPSEzbfX78pZssV7EOBG5TlwkFI8cG4090abyLFlv3DD7jhkYpQ6f1
diKebCKDAbxndDVyCBk+l9einOajgHMlut5f3DpqdWU5OlzMsOFM/g/6baGZIikQ4Xb64GoJwRk1
GnUUhmX2lu6uXcMbVuQFmdm6yecvCQLc08rw6fDioBEWxqTxn8UEMehejezSqIMiTedB4ZO+wKSR
pBvlwx8/tvmAFru9Li6wRIZHH+Ad7G4ETdYVkD8gey1IL7xBr+xh5Wxq/skNwRdIILIIk34Eu5yn
a0gRYpo9b0imAcXhi9zFIgpHNmkc3rxgAS0O5CNZ3yUN2UUIcskyy/u0V0KA7QKTIPKOJPOwIXBJ
SQ/mXNCAGD/hMf7MOl5FGBLzOpmKI+bLpUAczHg7xr4ojo0dRc3i/wWYIi12cP6/q0GcmMdI7lmw
kw55mAL3ysdlVLQcOgHR2/SwZDoz5EH3k+PDOy33cUwma3WJjQcU+H0QA4APeTS3FAfnDp1/tCY0
saazDOJ1KF48RdXEVcXNEJ5Aa8VFgC0aOq5owjX9tt2EptCkTYi77/5r5yOMnHW5teAkJXS1uHFG
ORxrbdA+EMIPiAkeZmKwpDjpHLhvxTEWmjYXZ3Jj0lX6CZMXOBAxfeY8i14bK4oS5BEQj+DPRQ61
4X+/oErFhZyysCtqWjR9xXtuN/QyYTKGJoUR2np/q71DZo4wX1IMwl/sI9hgBPjI6r/ys7RV/T+D
AZPRLe9ehEOqERS0JdKM8dOc6GwHv+LiJcv40LlNxJRxrqCx2WERQy+lNfIrgimmi5Xa4HAJfOwV
o1wHsrfR5g2WbaNPISAJ44s5v576FGNwabuIYMeSAff+dfyeLttlT5/80cSrdiOvaiZ3Laggrsdr
YOxVGgb3noGExcNsQmixsrkPFhdshFMe2wd3hawbEDNeKN1Y+fLBAGWvKk+o6K6wUhOCeCtovcO+
HnDE4neaROwHguB7mBx+2vRccIVRkZfyGNDEd4lz1nQrGScO0Lk3aTSQXeE4UUnGZP2hLkPYxEZI
xRJVm9+n61m88FJewbaCEnjvJmxyFv8YUI/h4nwFB73gVy9iB9ZA5sORS1URlxM/jLAoKFzC3klI
QZFdPSR8jGBc68keKClne4+mGM8+PP7kCT6Oj8TfjPSqiXMjZFNWeHYH+Pcwpkx14Zjx+v6+uKi8
U9lAcxV3XF1WCz8gzZNMJH/ipMqfU2bfqeLA/y4tEz992t3xjSBnleRA4VgHp+j0+6gb+wZ1C+tU
ibyEaNesqmnkKcX826WmX+lZ9G8usNuS/Owm620kzXH2fKOGCbsE4ZWwk3CluaHSZcJIGY2BMq+g
9+g3BNg7qF6O6hdd0Q3RJmQaekfWWbGx0/Rf6CFFzJ1ro9VxCgrsMkXLrZR36ZqxMAf/tpTllVNt
0Xi3EwS6WFY0vUxada4MNLYJBibKN1Fb9/K5FaSDm6T7jmw+ywkERKBgXgO2ryAMAeKGgC396CA9
OVGmt195LZ8EjtQLaXt7OG7/+xdOtS2MQwNxOHbA50Bdthtt8w4HhwutW0OaE/FckMHavP+WiinL
ypmmboEQbCbn7bUCsyfrla/zj1J52yVYk0/kecvk8F54MIdhUxgGiBRpEAWKbuP3578NyJZoqv/f
W8NR1EILFNl9cQQwyefo/jU/u9++W/Y3G23sEFurQdPY2dFJTsxhmIWAwgW+1SZg7jqiD+wB95V5
KijU5jUj/58QURh+bA0dGISm571uN+kY90Jbpw5Ol9le/8KDeGv2eh3bkzkAKoScHJnhqTur+osN
GBS7EdLT9ps2P7FL3nXtQhOsOQN+6KycEVI1ambrsNptGQbrAci0YzTlMNOJe1tDxzMUCk4ULINt
I0shpM2b44gKiEvS1yH22S7ClPBceZDCWoOgqOhYam6EPQ8FrCFCTADWBtEiX3PHw+zamIu3R2IJ
+j6WLlg6oUoSwDPTliOfMaTxydq0nt0iKpPS+skXnKGXNQBjJb8PTDojDeNOTx588IbY/UoFSIy1
0DQbxWMIOua8t61i5RLrWfeuX7AdpMywAcODoUCjF+um65Aez/hlBUmK5H4o0mLWdSXMYMWDKHBw
eTW0J3VtE26hbyPMnzBpnJolnUY6Ru/hYgH6kF8AlhcnjJYLsgMmZibYwyXCk/No4Sm4bJfFGDUW
M7fDSrUzvapD8kP6PPg3DzHZIkMfGas38PBD99WTFyr43gJ6O8/dIUFcO/sCkiUcaHStdny+6zlp
w3W7mlsknGzbdQrXdE0z+qSFdsX3c4WefuCb/0k5sUSr7lwoURq8tyAtBU+fCCCgPc6mYw0JVYCn
C+GIHGxKhuOnO7CL18XSFENhtl8tj75uhol8oUi2r25dOwAU7VFB2RxyU8wA4Wzct021USA/ZtPq
k2qkFPZXPJ+I+66eijirLZat8sGJt3ZS8HsjV4KENsN9elPSvzR+stIyfsr8ceDNKDFAhdSFrRRP
FYI6slypk7y8IH636GQDf44ee0/wb0hpqskL83kOh8P8sjgxWnlyxkqLDpaV0sSSRHxjLLsPq+T8
f0fyGyjQ1Ael8w/ALTi21d+GpEOdz5LA67Q+jxNmkGvBs+r03muxBI/1A+/rxlGuEe8AET255pXY
FqtiHG9DTr5LtjPEa5G5XbG18tRLiqW/B4x0HSEiVX2RrzU8FdJZMygreuPGH2t5VTSHA5v6l5Jz
zlHUdftW9F74FGy6VwjS3JabVBojEh1T/JslxaMo5RfpZZSSXMctmV4Fv6wvp2Bxdkj/XbEgio47
oNDsZEtmRQVaOkdYrQubo5C2V23vGJ1XEmXjmzWEjjkLvjcwV6ip0fjE50K32dWaSzO3uneHFqQV
aG8Rwkl+kxTTIqv7ADDFHcJpoofzWZW8YUHQj36y5cj9KUf+SR0Hf/zVKNjrrUQZy2zVQArdcoF4
rJhFgrllH/MWX2f30pjfjFys1Y/ScCYfXC/gdzGBB+2MpwojRxqzfwEVJmPFe3ej/sJyHwifXv5S
f4K0mqz40nVNmiGjYNMnr009L8xm2akEAbZqUejfMeem7uBeYzfRJYnnxxKl4vq4CmFGaOujM1cq
LeX1UDJhBljR/PXr2efelnbXX5lbHEvy63NNO1AX8smOjlWfXn7vSoYGBru+HtwR02KuK1Ns0lK/
pZc2qbhKRslyhI1eyoWdHPijZ2e8Th1y4xIodUQO5xp2zlLnBB19oys+ex+/4s/oPG1zqJKgJl2N
qX9adVWaMhPtu+y8NaevkiJeAUYS8RWk5yW+8VTyp3hDEvpHRc00B4aBu2ldzdGA+aclC/AfutgZ
sS9gd5k0GH8oH/M5Z3JCQdoqr7L1rcciLbgYRuvRRR8qTiISp7kRcSqk/VU0xBZ96VOtOPJJGmxp
yCoJDNF0D1tUQiE8fYLdaiPDW9K9xydf3Ld0hX9jXZ6FeP/kbHovE6kaplAcW4UKaBNrd7SEcDsR
9TMnV0PuLWIC/8pDxM1PTYGNeRU/SW/1AbuCMPwCexzEQmSdWrFaIDgouDqMXshMXaMdhSbyd8H5
+fG2hyJQvMkb24WHnttfgnKqKwnqVTj7xjCq3Y0HB76MxGmVsWT2iVrKEhCRT1XtRH9Cg1z+mnl+
PPrkeL7R45kd+fu5Wxx2cK5RDE2lhnSmZyv195Tno3rvWJGsEs0GHlPGk+ERMbpb8XYCXJclpNjz
/uW6HwsHp7r4nm0H8V2zG1zW2z/QmF+veNmexs80S+Dn8DpP+U1v1cMlepSZfpGEMSKBjOnczfjE
oYRH+jDyfKanSSypW+103cBNQv9mSRWFnixSTkOy19W+JodMGC9e3NU4p1yKnjAm3zF1H2/P9T/N
DlGpKnzP9cFmVgcCjr2b6RTa7Su9MQ6J7MukU/np/czp+qK7sczfN5SxpFIQPvMvjRZqCFo1B6Hi
xfemF800xaTevL/I/cSvLmf40+E4JOYQ9ccTkToCDYfAMgOniZ+qxFOHn6xZX9+n4gNdHay5lFRs
vq97XhccEIsBFROPg+RIiyATNeu7jo3xf8NOzXgXSg2GvjON8Ks4E3/j7YOLfRzsOf6EHv93T13A
gS8pamAp1/n6y1+cNcuPudd8DO1aNYPHRUjckyM/uaAYMYuXVOA0QrhxvooOsF4b5kPLLcktUtWu
vbSPQkeLqgtP/hfRODKingTq/lJgKTECIb0t184Mp1sEIexe789CJWNQ1exKcZufx9/4pqHpUnZ+
57uNnbfpdqMxgg4hJhpLYzD4mOTopQkIpGG9fqjlBj55d7/6nkS1dj37jugotPOZOicmby8dv6Dp
QzzQYd640cH4zrpaWbf3Mn9CV8M4vegvMWwr5BlDLvNeKL+Rgibu55GHU79XU48DD1YUz3TJrjsH
WLwyg8676wWdfWIaTO/6pV+55B9VJM2/uoYnyj1W4lFiQhWojV58z01kLWg7FyYkcbkKOfEGakwr
K6sX3e0XyGIC89lIMkhb5hXq8yhcc5bbJKhwEG2rpOpF3DNZD7tLJszu04P2QOx47Mf8rmyNluvq
ObW3ONO9MkuuFGXecClckzU+Qewodwzicd5MSg31XlzPlge+sHk3zEIKnhKrDnK8O9wUyCUPmgRG
+bXNzgXD6oAHFS8bwRBoLNvaVSwgJ8x4JU/XdR9aB5FV5ZdAUt0+tKiZJnl977R+zk93GgWh1MDQ
1k969VDHiYNdZ6yu4eJdLElanCUZsknrsL1xJ3vKL8XlSStW20pe1KJBMvo1ETtT1SN5LFZI4LHN
ztA7EkCyv123IGnfhOZELRBRdIToS12SvdL2uxlovzG6sd6upzGXIlxzzG+HjErjVPDj8gaELsLG
0O3vpY43ZYCGPOdwHyjsDlhMy8oGldHzo4TqEzktK+lzplu5xvpFIZlDnefnu2WlD86gvAsnS5jX
FgZDCHrnM2FT8g0MdX45DyKoqvPFtkHlhV1+gnDglxRHDbUdw7TyYZEM0zLrV6kLn9RnByo+BKmT
Q326BmL6cw2k2Y2ZJmENpuWR+5CIDe2wxvIQAYaVefaTQzC6OkOlBZuKzt0CAc0XK63EgAebCsiN
ni7IkZw7EQuTPYv0tcuU3g9LYerqXnavN4wjGRcl5xSFhhJZ82JKXyqr6ABI2E7Bki1IDHCOveV9
ZiEEjILv9cVsqQRnfar/bTStjXBog0kayCNcovqqEIYk4Ttq3YTc5hwVlpSguHkMNLYlaXTT5sUC
PsG07CrzV8V1VIKyv9iCxqsR79fUVkexxCO/VZTuZBDlPmhH4xSPyJazo3qHMu6iNF6cJIdz5G07
WhJtqtGsaJZuP36tfp7k6GlHlPS16hOHyA26GcUVgkY0KOUinMi2c/v43Ynfqb1OAPkhbp0TwaiT
EPt9tMpdc5MXOii+O8lwVSAiRv6bYr36AUB0mfKIjh7HWEHaUH0pKJerS0bbsOJm37pdfecFX9Ex
63IukiNQKjDgEmAIT6k/xl4/9M4qFO457ApSkUtg/x3n1bdliZMyjs9sHfXCMJTP1RF7bIQEl4R7
9TlksSwSLCItzG1Mzdn+5QFdxEQv5gshqtmA1iTX7bpMdkrk7gjJykLFq6ZtDJX4r6aAKsCqhSGl
V1OXQjXgUpR9Lv6MfQ/ef/s+24wiGPo1/OEncO3RzyF/np6zE73I76MZTdbA4c+cMBCf2IXWd6/L
D7QDto97xFKWgOMNhLT7LqdVQ/WdGU66OG0Dm7jhido0uELwXb/YprijuUG62oefZmsbJ0kdaiuZ
JAZjcQj2E3cmYgA8TUALDGg9tkptaHa3uniiSxFuKXs/ruwh88NU2FiNK78F9nnLgCc/992qs3cd
bQIikmXA6yrayo0Y+XPDMrbHcdKbU/odAH70E9+74g8tDcyMNpTMpf+vGcL+Kdxa2wmX16X6oh8f
k4Q/5/s29EdagVMEBKmOQTvb1PvbcD+IvJcl7TPqTK/basXVZzCKqidQiBs/+ylZQjcH2JB17paF
laJjpnaoQdzDbygf7mxZtn5+E6WAv+vZG1xBb85kJ7SMYW9cR+wWDNs4L5QfVC9fNV2bUrX+6Vrr
xNY1VLgI8yxnGJUL73IzSa45mGAp/PzG/dq3dS7/+aETNKQ4J2G6UaHl0A4Aq0T87vtNANWRF171
FeqhkAmTiAzgJYxUgPfPyReD/UMhjqebY7mYmuhXyjKC5sTeId1KHu32vIKxGMHelFQNW5iVszlj
lj7lMp+e4fkBQEl7utFPw2MaCFeASLE+M0J8+G0q4m1CBwzbxD8adhJz3+Fc/5N43Qx12f4cVjWb
oEOmgxPGRZnCuc0vE4wCXXeCW+IicPRo1Mgi5oZIAOm0rfUWI+dXFM5oqfH4uu2e3QHrMAf4pOJv
dSGZPuDxfh6MlvkbfmN9JX9tgXNJRhHyb5yeyIQGGA8n4xOfmmIs10RYhzKBYWqpeRyxIgATKxvF
xm1EgFHjG+RzXDnwtT1qk+oe515UODRBZgOYBqXdjv4vWh3kG4OYkmMaTPhGww+gYE6/CV/9L49t
JHU5QvJo4kK+DnVv/92MyZGDPIO0WXSUOMQ63KiI+dtAoBjvAOh19PwbxmJLuzTDfyNY52HqW8wT
rAGSF7xSP3gPptsYZahlWBs6TIUL+qVPlNtxW86EAzdCeb7HDBrOIzqN2bxzlnbaos07w2p6FTu2
1Qc2w2qX+EPxmxC6HIQyHrmcFBs5VMd1UpQHsDtShUOnLquNKm3Wxnq6nBE+NthJZL+qyTlUVeIM
KVTUVGrTiEkh0BLs9xO/OVlmTL4i+wpX/6OuY3WPB66xAXrsDktJqBiHJ3izRowXkktoOeqZOoEt
q5Rs9zOW5SXG6NAlidyV/nJHueN65i7ulAu8lewvQ5TZwA/4BN6dXjalIGH1jr1VOYg53BwzkFMa
lodnfk5Hc8jyVE7+1HigtyLKq697ZuzjbFYa+mkhWWyNLxvK00XferqXBrU91StjMh1Sdpb0m38n
WN+tkRznIJUz0XX/Agv3NwH5JWoyhdVFffqy25L/yfD3khVlSTkSWyx9mYCnectJveGAQhin93nA
OmeXwqagtuHFXI+SnDoElS2VioPKMyMDs6Es9QbHYe2dXixbldwqzKGvTaxGwA7px34aUZL2pNBy
LFl0sJT84BUphYkqvGFH+/d4pNrlaZ186cKJgxtY+z6fRbeu7PUcbWh7sbjjy8fPR5CvVFaoOz2G
wx0vuhE+1em6TAURYHXIEGsl7pwAGVO6IbWoxXWrNnUbjdjRWPXiUmIDEPYRZIRXawwE1ZpKTnf2
k3UusTXJpQ82rIgmtBTpGOunAS6HJlRrxijoIgHSkFfypaG0dDt1gumW6JTIGGV/vuL7bjt3OsGs
E2NFpmi1WxI1cek2ZhS/+8Xim0mwhzlcFMISkSyqofwb2BB/qKt3flWkyjTwgcmG53rN/sx4KOUv
hwi0mX3kMm37DnVqDN5g6j5t/CZtWtR6CbrodTbHi0E/mZiqyFIAR2hUEUKVjdpQyvR5g9/pTglO
PG1fPZDbXTF2E9KmZ/3mqYGuBDRJOnDlpvUz2jbIfl9TAzCm/BvVdNBBL/B6O2t8fU6J5r/gy7jR
0eIuaCT2H4E13ms7gbqHnVyp7lQyOXZabjt7vE5g4N/Gm89P0kgjGBCeQpRCINe+PLn6/ib4piT9
hiDHGDeVPtedOJpkBf2a0rXwqLY5R+hFn3BREMNJtY79T9BLCVecxjixbWIImeDipIW1+ymrlukn
ERPN+V061mZGY0v/D+q7FE+brOn8P3HcAib8R8k4i+VTauI4MDj9Ikm6R9ZysZK/+amoNkZWt+Vs
Xm1v4azXSZWff57WnBkcsym7vgC0g5oC92JspFeWAKaPGfOJ5Ka0G7XVjJCcZac6fhihqJ0d48/c
FfVlP/FIP/6VWdu6hKCxl1Ue96W1hT50KjnyCV/El6P55znhbwK7vArVbbJL6p32qK37GYIzRug5
nhsHfpT5faJJ+/4wyCeLqYZAX6i2PzORTrNdlx/IXiHSLWH/DMfm31gL5oJHlFkAHAfaVAqpNTeM
3dH+Ez9zSZlZpJ6AyszzJ/S7SruTgYntWqb2pjcqfKy/61p8pXdCyRWgZnQCmL480Xc10/EQnh94
KnXXdx1HOP0yphs1PEPEtRDj80Y9egsG34wgQjIMHgsLi9eY6tFOQQ97a2OtMc2G0mRqrofKy5Ph
HUr5uD7UPr55jCWTu3Ma3iBlHeU63sy55JcvFyTUNQzrId9CbMGfFLujVoVQFOVg6y70I4lBTbAm
9ZFR8dDIAz8R/dORXCTHk96WAEKlwKWbTsa18W2hTGIFPF2k3IIV082mQ2gidO4IhQquzDLLZAPj
+nmR7InvY84uZomjW/bSVQXN4HP3qAqiw1tfgGij1Ft1dOkG2ONQkj91b0Mg1mW4G6VLEVkhuhyP
aI5RWjhTFPPb3LnaPdd9ecM24H09J9JqhPhuGp1DycshyU2wxQ4FKG/bDul7A98PVNRFTEQZ6A/u
AAX3LlAoQS5ElaNAUoDYScDAQdwhTt/oofNJTKYejNiZC8MCJdpVqg+xmkYKHysvbaWUoXMwYFDK
/QPvAAAkc/QgBdXgF+kVJ0ygpU1R0uF/2ll5I9bM4h4SIlQrqZaEe2h+ygonXU8QU3izcGo6lrj+
+A85s4ctCpuBhw1yYfa5hRtRPzOea+AU2BloA61uAdcxQ0zv6p1VAPwlk3f5YaQXpLIEeb+LGYro
5WCIcgRJAPqVlaOq4okAp7D1hinx0djQHrQoxhGPsKAF/fIeCO2p7r91IDiCY9koR+NRY/C6ZhTG
68DZT6yyumOASEeyiQrgoPKBSsaXqbRGjyrRZ6cmIY+Pgb+25zhe21H1IZ/dMXgZYdi1Y1gvFb1c
3wRo5ZKEKpybWNyzVcn+lOgak1jRF7ITXo482MEqANHyRBqJiopN8kEWdtg4RlDNilYs2hkmKvM+
izEGnVi497R7MNuasWqSDAa0kIHOpi1lHFzA04tUqdICCZgyYj2cdgqDRxTlw9IommWpdPpabyp2
wsYxGoRCZKu69x3VDgSZYfuqXFJfpKXORlBIUgHaw5oo+KMD7Fhu/GX4ziNsuuhR3HYbUiL7EV/U
RBXBbgFygAqzb0iX8rX76QqSS/fDoqz/JnQTsBf8h/TuuOyQXH0i/3dWPTTwPLvs5YQ9XR/VMD3N
WzyQMbFj0FM+rdxyJFPe11Zpn0xeI1K8YsB1f5uaX8zl8ZQ5PAXxokBJCLek+8XpH/Mbthaa0rvw
tE3Jq1/cJDm2+TfTg5H5BxhUkKqL1Gc08mcb85NCQdYqT7V1vBSH0ZJ6ijMRgyW0AKHiabyNWqBL
EoZ1qol8xVlRyScoqoEpigu1tytjbpKg8zuGidsEjC2Cv7CXc450Mgo6+rMceZhra7MSnV16lRZ9
IeTaEKb60A/+I+WksUJrYAx8Q3uA2rXhZ1ByWyHLDdT2/B3+nnGWJQaaFEvrkRAlkL5DTx0o1xSp
oSoxzAvc1zFj/Nc5AOnEdjGsWgR7hW6VkgJTvoz+atPnR+itbWgN2tXPUxrL6BbrnC8QiGjdP0zb
4IbYEioeBokwCmchfh94hyQzhXtsJ+fgGwFfaf1FzX1QMP1FQClRyFEkLWbQxRa5htTNvNtmlZw/
or22JVHxSOZhlmKZWChmOZPme7QauiPqlL9byPfyfrjukjLHyqbuXCX3FborEUEhik50BTlhUkJv
bx04d/WCR4STrYAOB/f07gccTHH57ff/qu04eyadd8WPFTk+Qh7LNiR0V1vngd7ihytwbHjNOq0w
nbEbG494VQPPVtVA7FQCaTDOcuQTX0XzSleC8W79jxzmlsX0L5H1bgTQISJL2j+79DqFGp7EVIml
rHK0/l73YW2pR29PSM4FSYUOQKgmSkIj0PQrh+jrsfioxxHvhAe/z0mYOr2R5uBIAhsgA/bVedzc
BHWnokPLSrtS3IPTFrOwcUeeeS7HugVtHIsiaw/375EC/XP6IzdasPji01TH7KkbiIhBTy3RHbeI
o1VvnywU6mTfqDM6EYRbOELokX5cwYc+mUkzCxl8JlMBjOf3BjpCLoxpAmA/FYEbIC83BJMrH9hC
SB8OmGAVid0ba4Px+vjeDniAHpZmdPsplNiNOloHyzK08XbBRPPwpC5gTr2t5S5zNaHqqCsczd+J
nIv+B88efCVd4s0tbuT1cRJ4rAxw3XDrTREfeSCc0WXDmfZjXxdw5plyhdA0rGM33FUgVQascB+h
ZDm8FObJJ2ac/KbxkSYAxmj88XogJfmR55956ATykn4qA+ys6QYmbECfXTlGmxWDcNPjNzVLBz0H
BsKwICRuNo1BgjhR7kTjjdgtYOvuPrr7/BXhqpKFLSN9j+wwgF7srxGqt4fhenaRZjd11pRv/PFy
QKmhupp0ikFDNJt3Q6oFTQiJR9ZGrHXtKa1qHi3VD8v4MwhNIx8W51OFj9+7vyT3VSNMIGDOE3o+
molwZ1QKGJFNqBdepdXdaGdtPPk2YRSyvc/T9MWJ8dF0fGRyDFqoy1EylIjbtxKT7PWUZt2Q0E9A
hRiM9Y+KzQnAsTbAIl2NeDD5VLzilo2KimEf4iuY33eszW3Ilibm/EYPcZeRswzC49ok0tiAEeGU
vhy2GREXdti8rCsB8rsebeYgvKqe8MZVKH3YrTJm6b18KAY8kxXvSPkH/uotzEk69t+j6Cj0qOSZ
Qugiiksq/pdL4ISq+Sx+GSKnqszIiK3jxxkNLSmRDhyYz+sIsQjltFNE/VUI3uaXdy4qdAgqGT6y
kkp0hh6IVvA5HR/GCEINPdDuo0u0/uDHWz70KVR+kG3fVkq8pwz4Cpg/0gxm8HmSQsgZOg5YhgKL
ZvkgTbXGZfuqIeQYkS3qj2QMoqYJrLfIPKcuHHY+zUYMFTnwD7z7P7uBfMVItr18BYZtrpK4lC//
lg3N0NC1X7Lz1jM9pSFmI/vOjQlTSd1lCH9OJ7q5NAgvodMudHCD0ifIUeXjGr+43kcP9OSiwM9r
zWrDlhyrv6pPqXO2ORfUQXeYPzt/aLmXhdILm4nK/m7JTthRFfKRPCwMYuDufA5WDCnWdZSS0dW5
AQlmiaHU9muOmtfvuT4jw73iFIpibSwP7bnbgVbnHUx/qYLzIjUKGWWOqRmkjrXgg97gF0o07Rzf
xIAh+OlsPPJzIDZhtdUNxTc5YLMs+RrYFA4yISlaZRaYJJ2TT7Q0oRYtpVrX6LTfPbD7pEaT/q1t
e0IfgV5UlNg7EOxhrriS37UnPsgwJLIzuLjMqzXF80nXNdrLlx+QD8iVR7DV+SZ7cXq/c3EkT73u
A3bX/BFem1obgGg7DIFLf0Mslrv1ivbi25ak+sG/Qp7HTahD7QrrqT0pz2nJI1xpZ7AYqsaMqs2l
A5kZ125AWDsiU4cUXABlVzfnbWuxMjwqj67nHaaF7t2oD23M9VftXPv5dvgV0FPo5pQuNCiTFN+A
0Idw+JwlbaTNu5k8gBmUzhb6BAm+l15p31WaivhbQ0obPI5GUr/AC9ERfte9Y1suL43a0N4TI8kM
LrvZTllvShLHUNJoBTHIscOO4gbssw9Lh4vn9PeHUNeeWIqI24DPWznWkN8JPjl1JLE78TQ8dx3z
0jY5dYhO35ajhBICf8Hs96+vXZm3FuVXjGS2FW1kxTzaPRFfFPeaGtl4J52ZSSU5x/69I29FimZL
HN6LfJDvZKAGNun64oxgYIGCytM1EJkd//x2vnIbf1PHs+JLinqLdBkfe7w3+3trQ5S4FV9FNlk0
t+8hjsVcTe5nVKbnAoLVV6JZocHtbsldhQrzZ/AirBRRbWtCfUO7lc/IUBJ8eyCOadGNe4pr6Snu
6bNFYstpoC4H+QJlQpA+jn+HS/fE4/V1g7S09yqumGeqrqihuuJlpRM/bfKD9L10PNtOZvEHgD9A
/u3iirPz77rkmu8SdhsFEvnLPtHAGlEqWpwg1Go575vL4uYdadwEJPiW8yDcRXBrZybp9kfGOGnd
VndsRzcVvmOKhLBoZG8q4TK6t/iJwcy+cDSc0ODqLSokwQ/lYU90EW9O8bD4PK0lEbTLiUZbYVYe
o6NskrsGGNs2REythMUcOHP44CKuk3wWmHdzzM+loyl+7h3HsUOcAkp1DokPmEnxaQBQEyV0Qj2a
HPrS59wN+7XDRIh+dZOFWI1ZSNxmNwyULB+pT6C1nZlz8R+opQuj5gzZMZU5RJ/yUeMkYr/RZ4/c
9RwMiiYkdaWUtRpZLRIeQgFTTnYOLKTqkOYcfliwj3rO8N82cmHigPGLw4qm7QfPFci6NmNP/9lI
4nQl77WkWpIP3tmfDeZF27d9GSyozvj/Pnypl7zCd1+pKUpWrvtEwtSVV0kGkp9iTWCU1KnHygS9
6dShJbvHYVvwi9NZSXkZoA1Mj/9VUAapHzhsX/9o8YqbrdnS5FK6009oF0o2kcK75Q9UJi22tGlm
0G58vWk1T+mYqZLwRVODiCtXbw4gEOpjMYaQaPfjlbCEbyRSKPvv5qhww9W7LnVgCgvRKaY5qaEN
hP3i2eh++Ow81cp3QA+gPbsJwWoviC5NsxWnjTiNNwOm+QCpceZ0dRJnjHBVD0GLAxi4klcEmROS
Osu8QwTLAC7BT9U5pInQTxXfoMatiIZqJG/2uWihiR+U5HtuzkC0lxL4/gLTAggzdAF93uX86ixv
N7gOO5bPH4N00VTSF0qCvCTc5DHQ9EItZzUAFJn9iAiN+anL+6Ao1A/4IGKTg0kcCoHPCGnFJU+0
JxANIwGuMXbLnF/n/3GD+KZdZUnYMXFOiyq7ZC/KTnL7x9W9EMQRWIF/vluK2T3qFBRkyGsur8cM
2+uXYvqewqYLJC8gvj0S3WrGBSHJXvmqhuQma22RGwoSg8NZhB5vBuTmoK/GSocGS4vn/NhR2xck
wMFEXYM13+F6oCkGhrw2LlaGsCg5pC2ITf+z3+cFRVBahOIvbhofEKI3HzVjD+AE24OKmL437GUW
KdKOCUTtOuYRo5/kHI7Nus8hmmu5aXlII1x3HyJKRbPM70MyWNbqj3hknCePQk+vft/DtdZpI3/O
1qYsq/sdLoroI2BX6iGIUBOG6bN1sZZo8Ei0yhvFSLgY9BqKEKxjiI/CzBjiu4hJ1Yw9pTw//6oW
z0QN37l1WnzaFvzrBTMLzUxPlD4IvVViGo36bv8l6yAG7M8DfeCBKw8lAlDndVrXWiFLjIMGerbu
6rlfksQCKyrHlyWY2bGUv0SQR2OtSspntzLGIVkAybsHdD8peybhogLEH1TedoaJNlmMM1DpcOej
r5sRmXoKB/hs+Ow6dmxZ+MhFMIuoCy2sg9zex1/pvY83PhIcBOKCz5nH2nGb1PkduQBDaMThrvVc
LrgeLp1KlstiX2BtcyDSL32uIVgadRn2COBFD56cTDkWiGezIYqzTZhwJFzZxa0s6PQtGehbEPmj
W52aVQHRRv9bRjcBKoXPeF5LYFl79jqjXDO13yS0kREXETXNy42xRUczC87IbLLSsmrWHyLyhSLB
Z5kAav7HyN2VN8ojR+KNgaEpJu5kNZde2mpHjl0Dlz8XTt76xtUwZvoJfTnyYtRKYlNPqlpJJriy
9KUsM+LxfLzeqqiI+chNceF49mPDO4RfRSZimmavEBOzvqV+Oc+nehuT1ErCCeGAKSL3roVmLDVu
53gnxdil+r51oz958IMXzyrAleXkKulyuibupany70hNqJ4tagSG+pu23VZWQEy8mhmCcMcgK0jh
cnU+Rkx3MPmWcO/2p5Hx7FVQl+JK7wG7GtOW8fPlF/YtnVKEjOcAo6HwOmrQkBorkTamAMu8jMvk
pKAEwjluC61hrWnYRlP/ZgSNnl16SVf4mmKyXhOfjUyl+v7UncgQU/rpdJ0lRz1Xt5cnRt2OPEd/
xn7tWYIaJDvKPvXNUpSltg2XMvEHGLxod6dPj4J9FZ23ct1HaCYaURKr9sGB8aZk7KU9GVw1cc2w
Ck0KD+A8B/AcvdanCHWi0jmkzw62sJfl4pBwJhYi/FpbhxcdtN+2r8Bah5ObAc5AuC0zCjuwsjBj
xrpFTy3w4tykx6LhWAF/V+G3LZLQQXrYhgC8wX8r5VVlqmYnL+Co+PZQAJnz8T3I2oPvQ+HcEmxv
qDk4SF5PHZ3kB52HtxqWD/PwaZfFgxop+ZNBLHtpZBq/7/aA091TjWLevQYfPR+Bwx8LbCQDJSFi
utIWJnXUeo5SloNBMNSH8RIDO8IdkaFOAVEeT3AYi2KxP5v/hPW0dhCHr9is+t3OhqU8LfoPh1eP
tQGngAkUWDN4cGMOvmCjMESj0Fwd9QXDXDN5Gqasj3lD87cCN5n1g5DMSklFctqG2HEoFkoUhkKz
tA52Jg7yCRxRI1kGfRfTDod1moUTlasM6p5cHkQ35gh5CTG2jOOKwEAZAy2n9ZbcwYt3wEnZHpSY
rrsPemSDXGsNVyPRb0+dJBPKhlZrWI57k9SoreTvEPWKkIuziMn5rkArhfVs5/Sfp2v4Rrk6Rpno
m7ycP29tr/4ffQ+nL/fXccNDWGFsUxzNayluEnvm8S5w1gRm64oN+ObE6ZzL0R2fwspE8DRGk//T
y3WOmee3KwrJ5ZfqcjHA5vSlXIAnkHmtlWlxQSzRvSsBsdSYBFDeVPUL15+ErDRS4Fy6rSXcX+WY
Ng7vg7WK6CN64wIwtluDCRH7vtqlMUfZu0WE3jW/+DPHlaLD29KUS6BAnUx2qGi4vODtNv4IoOOD
3sQatY7v/MYuLANGjxe6ZvGw9q40F2u231i1j3pFByU7KOf+oTB4qMrA9LCM13PhqDHdbPoXdyGY
QY4l/JlS06Y/cBub8J8bFJXZ2pdJsGTQFRq4tiHkEzfD8m6nS2RwsPl+YACS/9fMt6qZmS3e/UIa
TDt6iGkoIKW9VPMrudz+1yXOYf3TtM3tLva86/zuFeKKxMS/HeyNaz2cenaBja5khs5ZHxUZok9o
YqyCEAJE0fPei2P/N1KHmavK58OvE6Oknq7pkZNAXnlHHJS+sBi938dCC/jZ5v/BzbFE0GZsYraB
RaD+hfj2eI0tB7oV5LVonFiAjZ6UfwycSwHKuM60CAa2ujFtQE/F7byHTs3vDwOTpGbbqRJzBRzJ
P40M1bd9Om8afZHkO3R+SxIqKnofm24D2iqK0rK1IbsXJn4R1PgCd3nQx+IByxtkN4mIkmv3t78z
h67rYmJlh7IOwWyBT4Vj0WJBN7a8Et5egGyHxjIdqANbiUVseBhMVb6xupWcbNNQRcVgNypKTEhw
pLsp26kslWl1XWBubkSW70pjvnIX9woSokW3Y/WzM7q1YEf8lWuO6BPUPmhmfCN5YYPdmT7n/oXk
B20HmZS2/oKR2JBBj6LZr9vn44W7Y/+1vYRq+PgvMV9mJ/cFiOgFfHlNt92adHG29+n9O0QG6rkn
uRo0DqO+EBgaGR3MI7JaRueRR31MzjhRu7+wqT1+ATABX0QRDJXtYtIKDpxMh2aQtWrgrnIJGSeN
dPc21FBIHLb6iG2VbzHQvHOep/JoJaRc/Vn1lBC9VibQN2qnLtHqHHvO66zjrlVX721bwg+W+bJb
aZzdLBwp2Ha33n8R4naX114iYAAkkOVNtEULdzIJewfTUAgIq0uUAcjIeMtqBHxQDzIvNDwz1uJy
hATnJkz9iAaz5KLY+s1DFzrYA9JuJt8rSpqZTtGab4YbU7pmP+RYYznPeXmcnH5NmW19ZA70kHxY
jo0cHflGQWvaH2SbXv3by1tPGA51xQn8YaJTTgUzJDZAjrmv5xmrSajLQGvY9do3mRgpAEGsbN0p
cpKJ3Tna4zV6VeEWAhiezDOh/qKsz13Lx0hgM60pFiT4AT6kf4keQr6ncmd2EjSpXq1GpROSzXfF
N37QQ0OXwx/p9IIAH4wuz14F+wRFBLX1pnrGXY7wqwxuaCUTowZWViCuUl8e0SknDvptJJhOUkBK
72K7MTrC/i9KNJHsZ1l7mMGHSerEU4EKEiYj6/+4ScHbNM2xSs/ow/OGcW6TlhVvb/SvA0ay2ppy
1dEPjkwNZtaYTG9AtThBzFaOxO48SdiVCikiDTCLGOF23nBL8SdxpJXJFR1PW5zTw0548Ol4pCRD
06NI/MoKvgld/IEbv8GglftM8FlK6AKhvy88wXpct26eX2BLkz4CUhxqHgiJ5biVP1RCUJCUp69h
KSkQKf9xhWnorMLcVBBfEQAM/EK/MwKCn78o1g82A6rAWoqz6WxxBBJ1/efozdNYYmgY+Ka6Pn5T
rPlDTaY9Ex7IBAfySPgmj9Uu3Cvk/letlNrfMN2Kx5WZLmUZrJ2Rt/hWmB3IeYS2KFviMDx4j64r
hyMSs+ND1F+UozTR8yIKuPGGAADzqkQXGXCzMXlOD/6lzV4fOZ+8CtrMj0SLCDNGRmF2HBBM0fWn
CzbeWeX/MjRlfrrIz1Q1NWaDnP2iKyCSjCIiy0TB/jvcuwRD7gHOTt4PsVdyJgayvYTEXbvTU8cq
tUe4tkJpd9o0iMJJVCyNRJ0qBdV9j0NDqvnh+Wk/3D+ZbTDydUNIis9aQmI0jD0FITRXEHsOolng
EhLv7gTI8c9HF+FFn4vBrDUvxVhppOK38feOYdEjK2Ld9uaT2dXlmb+YzpO4XwxJHDlbWDd2E/rv
rMY3T5l5siNTguYAdZDP96loRgnrCuej4Gh8XUQckwogD735EXCckD/0s+XU0pxHaAPfz4mqD5m9
WBla0gW/1syPJfCChMl8nYfP0iU19UWnEm7aXIiIMTXXHuEo+lPdf1DLw8CVMBKJp+UnXtuiGTiH
ky1vfeeg41JHg+EDin8yQ9s4kiDUR27tDzOJupfx8BQ+J83SnVMgq7eil2VeoopLd5XFg0wel6oV
cdC+UOfjumOZlwGd675q5NRydpFBxnnhw3fQPsR1ZVJ0UymlQY2hGM+2cH8py3sc/Ptmdi76SBNg
Hr6Q0dAtMhsR2/McAkIT8THjt9ZM2MJaupbVn+ISyr9YKbS1qsTlVh7s1hcba8REYUTRJ8MOVquw
zAe3bXk7CyCRVCCva7HklsY6GMVECWcmPdUkwNUQidJfHl9L1My7Myka/CUjozYEohDOd5QjTd+h
P4GyRnMDeKvS/Hpr2K6hXmBwI+mV3ck8uiaMnVibdMKJ99VTXrZ89h0eH4iIg5DNC81aj2J+cTrR
W3vRVuxq11eLNkssSe0WppYUhyi/h4VrQ53NHdqH8pdCEoscA5/U8SdyysZSfvrMEmr2e+isM/ND
8Zj0EvnIyJ0cHnYsdI+YRi4Hr+ZtAHF98isAbhHrUh672yrpaEwXUnKKGoXYktzV5NbB5RaTCwKa
Dc8paijQoi1o9T620H1PQugVMFJorkuGgT0v8jlePzW7B/zx/ivNrCYQG2Xo2O2wSfUAwf4OK+W2
RtHfd5kvo5YMcP5ogSp0t/FzmuS/C5XnbHUow7JYU3vfAnrIFSegYJBpjyzXBjGsca6hJJe6YNrD
km3YHovh8vhHCffQx681/4UF7F2HNbsShzVtP4UXJ6Xikyfi7Ad57giw7g0WTsgsjwsd+X3iNgEU
v+VzyYpaftYVymSNd9+co7HWalKDftbNaQHowjX06Ufkk0SI2Ifp4YvKpJN633pxGnyp8YBKusy5
7GFu6CqAXv63UOv5PzV2jKvXuxlZmuPhHjPUNwGxufuhleXnmhlzWmx1SCRbrB8wnCGh8mlSf+vq
2HfiPcdjmG5FxS3FRRIT2m9iB4HEmXP9vbenNzXK+IwUoo980hwbvAKoxBCx0qN/tkK3n8TkXYwl
U2swMI9K9RIv45U5/SXS2S2v1EDSaHsV5Ms+PvdyvkMlTDpNEQZlkaXa87tQQVVehEZahEHaeBrf
cB5LVWxHMbC5nbt7m7bUGZtOn4xTG2eGrMlcCf6BTbLNH5yLPPYNwcvu1w+vehWqDmtN4W6zy+Xp
szQ9pOAUbkxQr/TjMB1HEpUBPbXNDfUuWd3wpp4trKSnwj+V6BTuHQFxYtZMyGaGa9bBRrn4rV32
XsFqIaKkxpTlq93n2j6wSwXWb6CLriTwGCHePwSFwXxUZPfXz4c1on2ddMmlaz443KuZsHNs1nqG
JRKBf2HX6aNKWFa6dpbRSMPp1DAhsPq3btF3gINQHW+9+0NY7ZGruP8BRrwikR/To0VRLjdNi/j+
24A7IZxSzkN5myGdV1jofjOGzt4CMP2jS3QA3sT0Hg34OjRYmoEMQM3j/1UrXz0E4z97v21EGgy+
Yd+X231bTVFRO6zRYOl5Cr1/K8Ow3xiHfSyUyzeTXKkvaGpJ7pVa8p10i2LqJuWAW2z+a7nLIK9c
gtLK2LjrxI1TLr5AuMu7SVxLzfOggy0HnBqRQzQQpof0/U1A5VYUjfmXUubJt2SkFLDJp+FAl5kH
PCdSYB1bYfcrgL1OeqBHydw26P/xa8tqLNtG1g5xXCDxbjUTCE9x089r/R4svDTxEJBHV9STnune
AIWo/B+0CKuMzV5Z17tH8pOJxXBdGdMNIkHrxG94Qfado0QW6q6pPmBhCzgrBoV6DrEc1h0PaXL/
cEI/Viz5hxKstZYK0KExBWRuMGhvvZPlKO2pnCoqozPcikRxtIf1S+b0D3bDj++K99VuSfBqp3ov
6WAV1Gam1XAZgmD5knefYtyOkI1xmeEd93VDdjRiRjNNyPc9hQLzliBVj4+koG7xb6mrddmHnT6H
Zgb9ixW6vWRvplLwMhlDiE416BmEROoQVacNtLijUCDxG5D/Kpt/Eb8BvQ6ZwY+avIMs0wEomQr+
3NsWB9dwIj4GM5av7oPcsfyHS7UzxOgPZ4i+RWIuzS/ZlRVP1oPy+vM75cSthYnI7TzQs5EagwNs
wcXUWAwMXD9ufho2Sbq8UZYKEXA7LrLQrjbvXWmjftaGe7YQ4rtSopC9OXjGknbL5a4IuEZ2QaTQ
iRBm5v6xatWONBIBHXrGBJ+oPDbeVI1pttkgMnUSV4NLmRzVdUDDgpv/DNGTVBXzJwhC6cab8p0S
n0DMsyGKY+AquhgeL8XjeLkZAb0YnoXc/0uMIBbTnqek3RDMnxaPKdzm9CM+J63T33pE8NSuMamz
eq0gHROpjtxSgxRbpuzRFlAzA4WmNrmlgZk5AWAtEu6FW+o6hc/yMArOVScEE49nHg659JX3nKks
G7Dr35fopgjCZxdGAoBiavtOODStEk6B8tvtEYeOBdfjr32iWTUhMlbcknj4sQaj6e8JOzHFMs38
WN2GBrELhDqTPbRom0WjqTjkKgQLnPPqoEKhvy3Bid4hYik7TpNZJs3isfQzTHNPtfGpUgMUWjUc
Z/K1mhc/08KzACWG9nssW6Eb2wfVAezalHGqeJr/PRjoImHCCWJ1h7v90uSz9vzipGvGc3GAHRWa
7ee75wdiC2JxgdxQw+3HDi45H5kWsOAf5nTdBkiBXeaxxIcVJcsFmeTdP1OhgC2jp91JsHT/oZhZ
A0N/Hanl3XD/7SWCSN58Rz2xrmP7em+U1wZtA84hH1dTH3ctWiR3Hi5PKJCWjOjTh4Jh5pwmPwHT
NoMf7keOp/z1OfDD+V3iQYgP9vwEHzx9f+mCMcZKusBMtw0OM85GqktzDbHyTgNr3NhCBrOVDz3p
ml5pN/B4YaSIVyaZNGVrE82RyL9atiEEKBVs8NZNFA6dePIIypRAJ8/qzAW3Ji/anWV3VulzCpiC
GH+eSVvNG5y470CJXfPXsDUhaElGl+fm3zbqaLYUJofdlNusaXXHuBhskzZQ339bUnsuxCxyfWca
XvEwEISgg4f+K397mWHbUfCaYq9YCgr/K433CrDHsRqQeAPbFR7KMpOo3sVn6FftbOW6scCpLPSJ
UStDrDciZyEQS2cMgoRe5MsuqJ6+J/jmqDSPZqlCe8TMJjbEH39M8GDtS54kM0hUDU1tchEi9G3t
di3pzDO6fPBCuv37yK4uwgeHdDVg5WZ/y+se4sqmeAAOGWVtpkGUmKPJ2onFSLiNjzSuB5ABPIgU
hlegwxSmsFJI61ObgMMqCToWppFSuVQzTHi61fjserRd78j9kgzz4L6ubQ6x0qQiDja7mbNzL9EZ
R6/MzI+0yyQLK3Hjnn09WTIAhbqGXcRPOO2eD6559IEW5tTMT/3xHhwbOShy9bR3aOrWF5zqu8qe
Ap4V3dVTmrqex3OerSmNg7xy31c60mu4yjwuJ9Ebxft9hcQ6o/Wz5PpU8G6JhvqUjU4d3scdAzBm
RLsj6KcKhqS+fRaQMMuk2OuckkugKEVsjTKm9wQrCdYu1nnd3Vr7o7UvYrYBgTVDkPJ89VApBndt
IDbzhbN7Ownybuffr2NGOtL6ppGaGJDzO1rjpQogv9eSOev872394wpZ5VO3NB7dHYCyAlGMYdkk
QXQmXyCLf7ULnLzCucNYxBWI+df6aXsa5jbkUvX+gQgBic/Z1AoB5e//xJGzgvyla3thOSbVN0Ta
A4RKiAcLN9GUA5O8yBo8ICCSIhoRM7JDoUyWJpxzXChH/RSchE8QYKHgqvPjk2MlqwGNoNiXVE5d
OW/REoe6fn0qbobG4S/9Dh6FCKI2fDADHuth7gHJ+O45cUJ9ZF0enNkEO6XVRcpOj7EuZC1ZYzQW
lNuh110fHOgXoh0PXxuvCWPW9FGi6fxT2qUQCaEe/3QQcoGPF9wxgOfxewcrDtXHJXmvRL18W/MZ
bVTBANaW6diyEtRcsfXCVnQBToC0R7IL09B70MgDqLYiD95ae8LNADUDpbAsmCbrCfVwUCfmuTd9
IDHM2m3WtkwHjWWO39sAyJbopNd22BFZDelkEJCghgNPVV25Zrtl+Os3AhC8rc4Lr558Zvh8xC+G
tkjo7vRS4XV5Z2LzIasSSyjYW+DHVgZIsNWrZl1obiYA4fcMHUq3UFBeWPzdwFuof0T4eeR4D1YE
KAB3gz1nyOO6jWlgDq9oHLyR5lcfOFlhNTThwGiceBGv/uKRXJSGMkKBmm5oWrv4gvQSL/FurDKc
gQUa4fNUK8bCZyvDM2R+TC5tyz3rwSLkHVahRzvSfBTPwnRVmeyGdJn5d2gJi+MwDOISGwnZgsuS
UfSYvlsPoT3L0JPOIJwIiLZZzzutpsuLoXPwV6aJ98W18FWPAz8GBlXCVUce2J1ZaW0oHvWw4037
vSGTj35nUo9sb9qlv60o+chbi4Iu7nMgKSw7Qmk2SYnyN66WlqlyoPUWzulTEqcBRszxbtgPu9ov
FdwF1DoRwYpTUENqt58iwwRKahFqJudviWJqa77qgxlq0hOEr4AV9lpPuO9Xuaz5sGcZH9QXkQLV
iROl9xEg/sd2GBIokKOxxL7M4dyTtqpVHaN0srXBwFtHj3lsV+23BGv17TsbJu8tXBC4bH1OmBGj
BbBmzVxGFZvYzYF5PcGa7XbNmLHhxRLtZ+Oys+3Rm+ixZgsz7qql+uWLe3Span3MwmRQtb6oKvD2
qt8fGsPi8mZuTyVJ+s53hbbw/eGwdJfcq8mX94ihXcnMdq5GzXPIcewOgjadlaL7jKOzazO5KJwi
4x7Hjmqzmm6KDsaeAuiT/w8TDP5sPbWBDfQtv48pvzca0JJ4wYe8bUiA4lw7v3SKqQcONBNPNdVr
gv2iS7QeGfHrQuun94BinOJDruWm9OsLYLGhgoRW/WrpPK9R+nIpWZsdHofa1qk3cJCGbMEEhZss
2B3HBxdO4XlmobacyOyxpmC0JEdzb/xYibooP5fNZ0J20RUU34zetqLZTZCl8XL8cGweFfXJ46HH
9hAVhL0CxtkO0x0Cefb2wu+9HTXpm6yVXjdYmC4MW/gIV+a+U7dm6dOh+0GMt/xKYrjF3KLf2uO8
THwUgjQ2/Q3ATKYwmdsFBKVbB7AeNcTGDlm+Ryz+i11wQZFlIhR1sM5SYjU/4YAmSV44DI5xy/0m
LNUE7zSc7iAmRlR9FiFEPKXE/fbcXVAn2IVq7xo8o3VlRMhw3tOqV6qiqw4xiksV8w5bece2M3Qc
HgOYSi/cPRVB6K4qP9cX9ejVgyZTxlyXbz5v2Gys0jtPbYsqhF7rIymQZm6chS8dbEcuhms2gqCd
OAPr7SxmwNOLs236I4Qg2cYZ2aOH6cEwHGWEAmzrFLSodjW4f3RemBSgM7FDHfSiZLVBwEDT/Tes
8LYCOzLtOkkQ5R+I6mok89/fgCjup+X8mzMOlZQVgYR/6WQa92cZF+0BAg8rpfYk3DVoY4WRwWF2
YaTuNIs7+BcOra0Q0orPAaHJuvAeF8HT/N6EJzkTGARfQQ4NlbAM+Hl/TvzfKKn/sxOrSqBbfc2X
dHOr6W0CmR3KZf88udv5epzIvgtgM/Vu+dm5N+EO3+mUnudFp+TwnFaZuOjlPwDlhLdjLwIr64Jq
bc3HkTh4YO8gblymL/ZceaHw2zD6lv4g/G0CWKI1uQpCrpT0F3ezru6h9/OeXMxnXuQkUaGLq89x
bSTEXgsEQn0t4oTNaUT7oaBJpgDZ7rz9fXrbxLIygCJ/0RmHUavFIdZnit7UmY791uXQyvEHELz2
bkouARABaSedWONQOpSHJjI1Hh2BY9NMnUJtbBQEF4dBXhrWAN0VJflwVVg9IT+dCjiUzB9mITTb
dbvqgDubyPz5e+FYyeZ0XqjBFo4LOFwpMXWqB2bKZo3t1hrHHbcPKcYrW+brXtXtmiDzWDAuNEUk
vFMnWn5y35JvK+PW9XaRxm9rwSZS4Z6wxHsj4FFJNMn9tga0ChnSD52bS3i72i5AMEMhWmuQRy54
TfxKM5iXx5PFG5YPC7ymc+fSlRfbuydiDNx8VSMcnleaj+wiENiKANaFtfKf4Wf4SEvDMuzBSHtl
eMltPqOVj7QlJHSqpEjuRtLVZdsfbHCglJRQEK0kHj2mi6Uyw0dxStw/A3KsOIUjEpFWYpKG2o2/
i0Ns7e73CFonmJMHzJqqv1V+pXziG3q645UbaUqXjziQ2UEsVsS/Fwwk2nao8S2qkx29rmtM++Nv
ifK1VMRfUrjx3gSCx/Rdu0lOqTzAwC+MZvmE1t5sCOcsOQoKt8O/8CoD1qZ/JYgQs5V6icoi9BEx
QjjuUK2bYKMbyQueqo1fVCKGUvbHtTNfQSTfGuD3gK62XIUCHWk1Y0o/AahtRaofdgDRYftJ14UX
4OOY3IDbQEoxuiK1wgDBbLasjeot5B7h4ZD1riWIVmbTkvySs2ptPSBnsoKkUaVqVRbQJ0QehxxC
V7NJgMUtE5yHPDqBKOBDahMcxXsrXcWAiDcQAdUVO0BqRDyh0MO/zZl0D6t44uN21oNRJJQ1vwyQ
rvksfVOChlDjjW4tJ6Uaqqws1VGd1nYGrCkwZ6jtoZ+ng4DI6FWXNkj9CCrkKvqiqWoTsnvFfRny
5j3nGYyk7ChxcDj5CrNOANpvoQDJzAMRPrB9hrjAPDCeKjNkrSkiKEUT3ivFB6ljEFJRMbFpSwEP
eVT2/uqkQVse54pBUM0BlsgNUto53cxQp2M/I9dzWtn8hrER1mhEnC/wuKxz4duUyNwHQ0tmbxYY
2ipXSfcEARr2k5wwtQZLG+bS8O0bDoERihIxMlHPFfu9uPlU+Bz34nGOIrT2zB6sFnY6pkl8Njxl
dgdwk8laTYrFkPGBBOqGAjZSBcZJfCPPVscxRtaPz2VNsaTwNDmFwSQ4hwwvqU5mphwS5CkpbL1D
G8z9KIVMl6FxkT3TxDxRYSowxhLq4yl2SO+fnD0Qmf/lYJRFbsYhZAkloEMj0EL8MXUKHrIc2vlt
poGon0vbyEfBgTnYDMzAppsycUBvgE3xskNnc+kvE+i8VEEJgV1n/EK+Ohg/zwK1/3/BqEIbAEzb
HEXYbySOMGRqWQ7Nx72onOnHHggkWyEJ12OcVffJCbXCSyfgTw1FTGb6AFd8cmeHDp+gcTZt4k7o
nIz4LgSLtlE/l7PAa+fEs3r5g7iM9bgZJWbMgew7RyO00cdXeAWauftx2ftZOxpRgz87n2Pu40AR
YJedxcrX5BcnUsX2zDhN0SEeyumnedBqMfA4bjyZPFf6yAMmzIF12hLH3MZ9BbMPhNZj8H/HEyWk
gBBcv0Md7PYqAMGb/FpwW+jhdk1Wsv9b0YeeMpLU5nky7bWXxP5iadONzhjBrh5rbjuw/94Iz1Yn
/K3OATIn1a7O/AVavukfZA1y7NYO4wOVt3dhfokC8GCXoQunranQIxA4jE081cdYFbW5sb0J6JH6
u5TCfLlIfZhjonClCch5wSzunl4hkiT/Uv6Gxkp7v8QCVvY+F7noaDhe6zNbg46J6BIuFq1nxN9H
jjNEiK4jni47SF6u1mfZV/jia+x6s9ytpevh/VNh4CBDAY/ZLx799LDzy+zLw8p23QpvJw/tH3nm
SPI6ugwd+f2dAnZdnM3fJHXAEI0ItqVVUndIl7WYhEIjZCU2xWryQovPPJHc2ZpDdxvmMTQPwqjA
gaxD7cfVhhmyA6C217h2uHAOEfqOV2mu2cqU8k7YdzhwJ//Owq/Fny8cAHR/2Fr6YQzdIU19NqOr
pNOSXaGaUhwupMjpV3JqgcNSx3nZEpKRIYtryxCtydnLyCykyrtLO/QN5unN1WfBupC027Je8x79
+boUBEaB4zL+UywyRlFouIKlvRGHqEfUNsB5NFZtDAn/v6PTQBfGmt94CEweuyUtd90CvjYYh4y7
NtVM54TL0o5Owt79jm2OYk5QE5jFVcFQn0xlkviOqYhN+bTby4DOeDbqy2VplDxQZfA3EqGTeKGI
8HrQF3PPyThg6FmaiS6qhY7+1S4lOUgJg1PYXk6d916zmQ25bAFfUEZODQqipDjYFievyYL8Kj5W
xDwXKoE2n3z6vvfnjwFtksdLMWqlHBiBBgsIxCgVFQ9seh2Rd31VSA+FDj6lei+VxF+3ddL617L/
o6ehKiutNs0eXuWfkaNQKYRqbdRA3pn2srCs7vFz1FM4PDJ8IFhzc+54bZlVvr8s6gdoaSKvAkQ2
/7rTvnkrjHYt4H/oZRFrCFv5Zkwe26sAY2vsMzmOjA0ff1cbhw81zOkKcnzDskDLx14ikStED+kA
UVQj1zK5KgkQfuRLlisS3yHxqU6LX5fbNFgpwSnEG+brXgvUU4aPbVSkMcyRRMEnbIvUk1qV/jcK
W3WkrkBGNiTJpaTxWO3jAmRZYx2QNddkpI7YhgsyvTUzaXoGEOmiFL7NBvPP4LVzlRjfKJ61M/zw
Dh3xR1lwj+0Mi80m/fR7BzhNtRh42FYWuvinf5dSSpGeDCIgUTeNr3BohPWC/jwPWjwAhSU1MJSf
JPVAKRAtOZbUjTIxGpZLXTbWvnPgLs+ps1KvDKTpZ0erpG9cZYDEgnX3VQJGV3gzV06POF2bCF5z
+97oJZIS1s7tthS1fPC6snZvMKizTBYPKXbSV4j+D+oATK1L8C6vIVOD3mlbKlL8Zh9hsq6P0W2L
SC5KXKJ5/Yx5XioL8n5YWWs9kfC42hXui00b4U7YpgQ1c4SzgQl+to4fZuiNx7TGB3tbTAtn2FqA
PwFhffE1ns9h/r+xUsnuSl/QIjdiYb2OsJ7aZpE2TY8GdCDOD+lR+RBtcvZcBnv2UAW199+CEPF2
gUvxWdETfkzbrDgCe790H1vn4hFUeAUQZZHGzFniON9byVe2UnO7I3GecbYsYCzUCDkLNWkYIMQn
Ppd7aeq80oj2xOi8566o9BdO+8nLM5/DP5c3vhBW3CkrGL+CeORjlrCv8FqIt4Au1XEXKvtpoS5o
EQ4a6SLUUf9VfZRxMOawmoBgJHiOkfPsV1C+PLKdv5KxgQCO5BV/PHh369SoSCz/TcmEVtTBrZY6
cqc42YqhDfbJL0zEyTd2CAXuQyI0p0S4fPQQsZBsYe3uSkUXe/vqmStt2epTB2ISPZVELbxlVkHj
UGs48dMrzY5KL4oCTlHJFpxOCzKiUmpn7LJVJAOZh9PGcEF4xnGzsK6WTIrx0VFXhJKYKBbt/Hfq
Yhpl/Rrr6afKiaoU5uByufa4zjrJokG9O7ayXBuz7QsG5P2LhjJDo6tNLM8QLPxw5GT4CDzWjSih
gkGrLEHZZIv8Qu4RUqtlMKWHAmJjiCYpbqqOoE7WSKL3gZnrhH36gRbUzpcBrGiUOHh0Lihdo4H8
nIMVlSMGncEbb2O3WLUMbMWuNK2JmOLXb73hFH5U0m3bxnWm+ekh5UAH0voHb4CIwvrh50l5wTN8
TMEZRVQ8Ibqy+5fjBYvd1MWQcOW4y+kSmdTrv6RsGWLpa4psrxGIKYR46dJrcVwwd74tkVq88M4s
O6HwPAFE9JB8bZVpaumEa+MFApseMEWjxERI9TJ4NFzRH2iMbBa5X83XNVGSA1GPIcEi4iOIujCz
K71fy04w6ebg+sGkMaUdVdvMQcTqOyJ2EpCXTSMyxNV5Y4iQPbkRuJd7JOinHkkEpY03mjv4XuOw
EepOUiqbrmk2rsxz4bhcGAinJDJNf+xGnTC+nUtVzPy7cP2nrO6KBwtdJaOTwl5OhmwyiWEqnR0c
RwUofLB6blovmr/LzFoFBcaIhI8fvqlgoFWp0id3H9fzOvV6IwDJ35nTsqZXq0tYlg6CYkB7CHle
tRknWAWiklmfmYFOiOl2ZBYFTSfhGq/71RGbmIlnBnUNalQ6cP/hq8wGDtac35rD02j9tAPLOiHW
qXoxq7s0RHKq5Jul3xXwJHcJuuctnOHdNajMHj76bFXdk2lbHpWMToOGrmiuqddTgPI0FYqsbhko
AgEQ78RioRDNlZ1sXjT8xUZhyWCJ3fqemb9W5viNlQ9DanqbLrs1LjpWVqBdIrvXf7fqDfJRdzyf
bHAJIUlkKHsQixjUwqGEAj13Y678MPQeZ4Arigi8zlPMoWrstkY1N+4oZgehcrt+Yxshwp0TJJto
KLMZoO3MgZS7LvEy6w1HX+A94kTWZ1hX5Hlr8TefiIzqbT9qhUCNm1HTqPaopmuzgCuiKAFHvBW/
q7EOJPYhaWqVqITcuAllXYsPYLUTbc9jgS22n3fMOb4ZsdePx9H19bAOFGv9TiTPEksgszrK3JnQ
dsY43LDLP7gW9aMgY9qA0BsfledUP7R25aYuRiOO4JekS+EXyLmd1rHBln9qoWn6RVvu7Jw7xGD6
WugrPxiznuiEISgvTA0LegUgz6I4TNiN31HQKbnL0or1z87h09mmehvkwTfBI2fga2GeJ60blAtH
8CVjCwpz6NF1a7ZBefLdG/1BZiC9NA2ldrmr7NAozQ8cxJU9OzLSB7l8oyaRE4/KzLqI2bv5epEJ
JMAYdR/bPfa5sqFsbi70IGdhZ74lYEjEzDCh85lfm1t4VR962GQaJzGMO1feHajQh4YqodbKzxeg
roRJN9DtEYq4TEtfh9tkDZ5Vh/b00rirkqL1NhqCQCAxNI2k15nIS0RAZgLGNH04WIMVJcRnwZsC
PET6FsiWK8QXH0W7h/6fMcc0J9dVOXEKc8PuzYqQPuf9cJqekZffOXd/zyVTwZ+vZvvc9UM8r/HW
p4NnltROTiwf9uJyEdgZz706omRO4FEahqvevI51UQ8S/Nse9uoKvLXQnsV29NyPsTPPIO3wBQiJ
uMADfziald86QPaXCK8oty6Kef6Z5AaHvCYYkW6ZZ9XpevFX63Lkc+6vGCZ1l2HchHSVGdVCgAdk
ipOrKKH4WyvQqkFNytvBEkra6bHF495uN9R2Aev5N9zNdZw7wYOpw2Oz8AX47acetl1AUttcQ27+
g+Kb1k409JP7k6Cp9HK2NeH7e8vqDL79+unb4rHREPu3Hv+Voj8mr7cdKMrNVckhdxCc2XZee8Zm
+eKSl7CdBIfQMCKCZi9h8haX4q2WM0y7V+/mi+zmenOhUF43uZCEBK/uIbmdr4MQE4Wv5zTbKdtH
TEDx57IVnMWFBsR1K1SC1ErRhQfa7ZwDpMqBvXdAitALDvxfJxjvm8rScNuSZLaLv6qKf+y5tGM3
AT23OQjfx9BNlMj1SDCuZq2T65E6hp3v8KCnszvCeTbpEJyBX7tX2bLXcZeoil83h9rweHT7EbAL
x5iR/GHVqSio8YkR+NdMQ5zf+ey1vdHmxAYfjZ6yL3pL4loBY/E76oMMArW7Q/FpVW5Xm3WHm7Sj
5o2wBVWZNT+LY//wMxeUzZaGNh62AP1/T4QX4aJOpdRWqpp4DhJ4Fn9szaELOTmp4SaeV44/Su5L
3pNiN6qQQWsrZaV6njS2HeYMFKfV5ahK322CDeNhQYfdrkuC8P5neZRkQcRlVoxzAQ2YSE2nBUqz
ToJ6VDdtRqcEXGx0s8guNEzhOYKEbQ4EUCJ54LIdOFxgbItgELRWdWEYvGSuwgCr30k+4ih7F3o1
ex/KXURLfbVV4vqII1VdYhj7gh6uF3Hn3rP24S13uIsqG9n5PSKeLx/Vh4KKQ5W5qiJBsUcHDUAX
qAXcshyuKz41jCViBfT1r/S09RbgipaSHoRCIiXx2Eu2VLwD6+Yx9jT/yAJ5eqwyEAF5zWqw5BOS
1dphrGS/g81GB86AbhqM/eA5sgsrIr3pM8AzEiqnlJXnFAq3bs49mc769pY3ggwjoiUyUMIF2QUh
Ti95MaFRmnMZGOkDevuTVCWBrxSd9kKYWemYku0wwOR5Qdc250UNAacJh0CDY39YfcYdApsQX6eC
nOCXe2GgDPR8PWmgHHNhIJnX7Uzzgk8YgYmgJIJiugY2Xby5bkTnjrz+HSpT0cz1+9hr0ic9hAnX
CLLQnaRm5jzMtDmNXjHyJFE4ShqAID6wlqgTE/n9vIgKdl0mhqUFDm16knMPpVN9CLUDB7Hh9D72
1q5uw43l06Dsr66/q7tdGW70opQZQ2JTb/xTDmBz59meqZDlBrsZy/ZUZoehzaPNME0FNSlWUTcf
j7N1a8ZG2N44jo+U16pgp8N8oJbcKvNGVhEVSVSBRkK1brvKufOQBUvaUbd4dcMZGob4clW15g9I
jQYnYtWaj9QmBlLfeKso+Wt47hYJdHuE3ZyYJLk+bot0XCTHOkj8lb/gdLiZUGQZfe6EGRtrmK87
3fRNm+K04BtzB3xcxoct0uHG2R0phuwQoBqXS0DQhVZY7Y0zdkEICcGs68JO2zPuzKTdRWtigYy8
ol/IZWTFEt9hfQPVXXjtsWq1IadcGzeiFoT80/+8GtHSJJPoKVWU2lfmy2Rvz1o5ypwDOHjHCdst
SFclNl2ZACMUhjmHOp7GdSSYf50+dHfj/JbNsLYqkr65UJhMP41CEg5TyQAQ4X+k/1/gpRK9Iyo0
e1/SrNqJfpkOQrV9EX/M7ufUSlCgYS5v6jfC253FPBr+gjKryofKQSl1oi81mzKxn1re6RPmWi9o
HTJrR9PDmIxqwCknMoh67JhygxSZhq228KFpRVlUP1iaRDO5+GD6QMEINX9bAdVaf2yk5sWNOBq6
F6eotJqplz69NuSG101hRWhWwem2+/RdpCLUOxB4C+qp91SdIqRCap4XAPxnVFmA8RyCGdYZOYaB
oNZoTF+IGk3LDpXmf8uRVwNkPuGq2lK5NVF3fOfNf+WxXbmj1STV08KiI4h//AZy1O+55BliJSLV
iGE/AB99eNw+8g2QPIDkeXI2Jakq9K0iI2TE86RM4/2Wuq3MYo5wc7v2429O0PNODZKnsKkbEgnW
kSsn3wODbtIF/QZQ6swIDxtRMhYa+yXn+QitQ93uH9CU3/UVvL3olWwIG6FrA7jOrhZhwkc8sn4D
l38tNrJ3DjDoYa8rcYnqBS9y49z02S4OzErGugR8KgpWQvME/298CbjYaY97l19RWM/9r9Km5oHs
r5te8bVFWUYO2EW3Lmc21zjdhP3AplEt/Oy2gqc7D6eTMDR222BpTFLzAgqthz1gWWBhRojPc9js
ShQuPwzgGzJf0H/tOUg7lH3Nv52Q/qGaNfrqeGGMVWUP7sVV0Pj4qQfEhdDfpeUiUJEIhuUcedXS
g4ZuQo0wzuvOzOhsuJsmd1Hs3wUfEcl8m8Yyx9xwkdw6fUW+pjzF+LVDbQmGZr89qPCnuIDW0099
SBJuZqYpwIXEa93OJEsKLtRr1qG4mxg1FPmumtLbZwLK8QrdkgSLn2qrN2gwGfarOWjYrpxp94jL
2WCCKGaZCF9LEVG52xx6lscI48f4NAOLP9+ERK5JqRkfxjv6xYli1vICezfXtdRa67npf/Ijvk0j
n/WKUz1n+G0opvWicElj2SyBCZFi9UYJUdAYqsD/DlWFUxmLULVyHfBHInYFGna5N1VVojqNvwwR
3HQPVb4jbCAHeFfE1vJEmMX0ei+bLTxnOVLJpYYtBckBqQSNrAPVuu/loqVnXh+RkrOxxjNtgGiw
u+ZQ/E2N7V8f51TQJ9vw6C+aZm5ZQCThO9QlaVx/F/TDCEaXMQxURXsiVpBBQ1FWUUcgUdSIDPMX
yw7BY4fDTPV6mL8/lJC+5AhAXW9c+6UFPUbe0rXCQ3yiw739PQIT9g7Kpzugd8VLx1NURBIZRqAV
v8C+9GlSZpoz7W8j3ncL2C0WvmTJDj/EtovsgwuCBTcHP8JlnIeX8V9OPK28lvrHZxYs9UlM8Y31
+qMgmfjzWK64CjQOQQgR4ePsa5sk2LkXP0MUMQ6J/J+P/c5BsGHNVbcpWAe4yt6rzZH6NUDQZQZT
LckgDd8jUdmVL4JxD9vaiNOMEIHtx5EYY597rozZ9VvHfA7kwt4EqKwzUrrwCK+IKbao+c6eALoY
9HD3jT/mIF1y3OVheFX1ACe2JUI/iNyQSyi2lSLMdYHG9pwstQTXhsJ7H9i7DDzp0a8fY10CpkeB
ttNWKoieKgwzYFyrJB8og3vGLFJKFl3mhPnmAo9JCINjJJRJXfaCLr/+MeqI50KrUV2cpUHhUGax
UYL+mmroJmovamswGLfCI3xjHRgK40SOKPaYQBLJ2gY6ASBLHKdBtuhCdbn8hbrb3EV1sgshulWW
/9dD8PgoXYCOz8KPAPa7ord5718ugwzbM6DUWX2JjMrle5h40iXa9AjTnBLtoYeBmHlbHzR+YJ1i
nhk0jE4O3KlG7ZHmxntNUOmftfVrrsqWq0pDBOIRyrMVUsypjNAhqTzhgwIOMV42kAzZKXwCdaXA
fiMqXfN9X45hW+rj0D7UbWqJUyMDijjyFh2YpNBDOKef8JM1ejUUIBoMHPDlhTO1WkyGrpvJaDDT
vKpyaW8NYVqepD7vR3VojTFdVR8rGMhl4S/1XOD/SFqdRIPQr1FvjvbT66TN2YXKJbk8jsDFz8p9
oRBWLGaVBDSPjqbZFARK3rut4NYDCGOMoLf7MKRHY4gTqyuSChDKCzyUYMFInddqr7NVBEVhyzE/
AFy7bU+mEQEy8E0t5e+zje4HKj4FZSSKIB++84Tr+f8rI8lM1y4iJeSVLpDMXcM/ZyQBg/PmeGNp
dP/YlRva50squGVaNZr4S3bRBj3xDASfDW/uNZ8kkVeMDQs4DlAg98SgKv4kmyKzi4KoNW5Xf7z7
UMt8PZsfVaTAuc6PQK7M17Jf6KbFw3t9J3cKPY5VqT6m849DGs9qJ/dGrlRnxPkk6u01gBFyLGx+
b67oHYkAIgRKIRCrBeUpln5E3I6kfrOxN4q23geHx4ZTPLXyZ4UEA6tC9j6FBwf14l/Jo7TytP5r
B8h81z9r8oIjhV/ENrlr3uw+eWqGx1RV510/o7yS3Qm8O5auVi+LxxGiset6HP7maEjhmVyBzJa+
NmJ7VoT55ibLfz3wg13tBGWaSTNs+IUDMZkxTj8zJLB4YOZeyXud+XEALQbmQ0LkNVJ8uq4mhyLy
wNIAgDoeHk0E1DjIBXa5TvIDX/f1ZdtD+W+m5wSa6oYKURQRvU43oYr74flMnEbyBTT+bqIkXN7O
tVCWN6CvmZGzJB+TEyyib48Ah2j3NC/tOAVQO5yFxkVtJGWrnCbHH+/M+isZz6DmHa+nEkrzFNAt
obfaxHBETxgKXbMO1gXpYuTHYZThuUVwQvdBI/9e2Zokx//nHhfRblrpCHV8qkQsLrsGCvMbYBFT
mEGJFww9IPZMiF8MDOE4w0AzomI9EgnTKWrpzU3nSm4t/oNsPo0V/9da0buWmpOzOvxrxZPASBba
Y80o/tRa7XoHMm/9WW0USJstFK7hEdfMEHsi2AeOOgK92EyYWOWqV8maMsMVunZDxVVOdGDIvEzj
boS5hpabebmIs87fMswqETZbE5I+HorNgmmAdTefgnWLPTSYXysMvCMDUqMNOeVctVhS3/E/U6ba
2Um66rDxr7dZgYbpdAl1zR18qezphYcXe/i5pcmfJNBWXOXONX/84k/CANgSolEMZBcP/3Lm2x0B
kUjsDBbAl6vQj7WY5pyCPeMOJh49IN5yq+iIJhxye7XX14rwsbLQOgzcRpJjA8w3FbiePRDYMKdT
Gm1oh8RFRurpaSqsPD4WQ5r9Fu7KOyAehIqWp1OOxILsZddwTjMAxrQrFLSMLR3rgOq9Y7Fw80Dp
Xdv5Ue1VScmjMza6JOG3lfHVtG1nAWfAV7lpbfEkUXGPW606+RGHNz/PP4QVvX/56PX+kiP4sjcw
sJJ6LUOMlIW9xHXQqYVKmXrYlq7yHZoMV276xj7YPY2u/aUmq1piHf52e52PbqaEcESWh2YD2Qpe
Bn0wkolKxqEez2bZv7wbBPRslRh6XKdsiw1LGVerMByi6x3xKIRKIyOfBgvz8t7KtYrQT4LUFjOb
UyHEaitW/dB7NIwKtQP0BDyKHy0RU5fINN5GDkan0dOOvHLPVX4tNDoqtZ7MGwFbbMFUboaX8NZ6
8ZkUvRdUf/xtHASI950jBS5/YtLmuyvArNpCoIyeJ1ufRCoha9i/2loa/soCU0GSupLYE4MjnESI
cx5UdHA8oMS4NfWuSgr8KtR2UzF3XT5O858Ft0uZhKY4VDUXnTgl2K3OKSX6m+YIOKJ9sv1taPip
rlfF8AGSeGws6cy8caVw5cGUj1jYH2gSpKs4Lh/g+ofD4Abr8b4hY67Qfj6KsIeWG7W4Kiuuowqj
TOLnyEYa8z9Wzfs315C/zs2uKuCgNI2Fm2yex1CUl+niOwqUxch1C0X3wekh0jzyaMK5GEH+no8t
o3t7z7ExnDeYyry1OcJNoeUZxIv7wLVa7ToXW3kHBEDBFKyqKKKdz71DenT59Smeuc48rQ5sa/s6
ufx6yE9HJX8DCHEA/yFLbpQ8KaroxWiKy1+dVj8RmjD/+6YFUVVRObsUI9wpVOZIIaULjpXAtW/4
61/JPGtxvjZras67x6RmNgal+JVccHNmd0xuxfzhMW6mNqTK50rLGiZgmGLOuBPTvqDucboBrRjP
XrxzHq/qezBhHYAWWxLKmjgIGqETK+yHeoSE4Lwv6yVY61sa4KphGfa6Xt8D9Jp+gj3uLxUizbDQ
DVAwnMvymv40ISq39Gp8Fzbhq8FD3QUekG/sLlcnokzpFqmO3QqDRDYyXgXF+xUwrIPigrhuRsjG
qbq3sX1p4vquvlBej661TUzJDuKtyrFSsu8eE6jsZHKXmbC+R4hBLzR42XeqN1/8LREl5yWbVEX0
qF8dyKD0zheKdbJ/s00Y+JyBxf9KBYmosnS4EH82lRIgjbDeAdAUm3T5fhE6tJMlMHJuBLoSI7bc
/0wkAwHL2FRQHsBNt1kKgEVq4mFNyGkI9q187/LCCLUw97CbBldgkVE5WPAZkpAyXboUJ3T9VFkP
2sWD77ybhXkZgODlD2AiSv7TWB9TMjDPck/mt3GY/FMyJJbw5Odbtkph0Y/XMZIYeEsBldY4jnX/
6DwXsWvqv2UiXvlYt+/eFBwiOKaffI+WcTjmFEUM4wsSt7fLwQgoD5frwCvJ3//Rh+XypxkXmI88
MZySypnYvpc6md3rNVR/EJDJ5pQUzaIwemVKdU3O3h0kQqpPYSt8eTGSLWOKOBMEnpWcBRsjDm1T
NDRa5FLQ82KewbGVR+//QNsgK+3n1Aa9zhX+n6sYMOYAb4KDn7mTeAxcja9KPSC9kGk5ZCJIJjze
Z34v64h4B+FuPeO8RP4/Gt42gGI1LDyi8t8VRl6FKjRn7lI9i+Tf+A8LeXjJ6dQe2W+jHA68dm4N
HV5y1C7qyeWg2IOxFgApnlIRMGpmTiuhX2l7Nbjo84hgWzhajeHVJSPsEmVdnNA9a0lasMfgz4ck
ja2IAE1R8YW8mzrhnTouO/sRMzBm6cPE8LvLUs4UMyAuZPFq98RWltfHiHZEDSTQJTdMIM8QJffx
YOD29S2eekYtJNo9wmmB2CnCM0aoEVIqDRq0A/a369CHRlq7FI89PmvfICVLktY7OkOmSVLyvjQG
5eOxT+BfVYKuICex58nJQ3pEat5snS6ZEqihdfkKTA8NiSK9xlVmLUexQKZlNpssq0PifHaRfFLP
6dsTkRe2tERkbeRYa9EAR0fzBXvTKhWIrlJCbZ3a5kO2OdsaUGhgYDiY8mSwhXg0KWmw5sZQkezD
OHI0CMwCTSA59xmsPhqW2AU+odWfpW6M1jUbaU7KI21SXtSzimBxoU0v8v0HzGHUvqgh5wjy5vp8
7FFf5SN/jg6HwD/Ll3ExL39702KoVrsagNlGhKCwlkoCb7a5JLVqs8jZicAPM8ni/WYtmIKRaYDm
VCYi7dK+w0bOPn7trVS4bhiE3H0Es5ICauM/xwyDDoi37vZz6W+02NDnzm+7M+TNwOe3rLBbEKkx
gxxPyTqpzCSDVuYoQOrroBiejFccfQleuRVIqOm6EE83OxTgnoIf/5u3HUJzSwK7V1VX0LoWUF+N
/opBhLf0z8fXSa97ADuiJ3wl0AmYV/Gdarg1ggU/jjGqd0RNvuztsTlETqJJFK9egPCmBY9SQCk7
VQOA8LJv3w1O2/dPx1d42lzp6x5VCDEbY1fFsvlnxp2yE44IYrXqN3dPLYDHhJBXYgZS5oV+E/4X
W5wI5Wr6ClGLSjGJId+eDWQwjinzjqIB6tMuLiYA+zxp/Cz3m+36NKBCx/g+FOf+On2hfvhcUJm2
HLZ85+yF9cKqsMoTz+i850GQ7tFDGAIDUvZVptdNuX+gEoAQ20q1v6caG5qmBGMjEpI5re/SQDmz
zzQfX1dR1TrqEZOpfOaSGZyvCMOBkyvfG9VRQEjskBTYspZLpGYlLD1mT3dNHvyrssegBInxi2//
JbSQba+ipME/jz42yVQs6LGaCftGw657J2qPBZEct7i3je43RVzMClum8EDMe0TKYXC8LnRq8axX
7KEQMS4xywSzdwifnypzXMqoGSz8PC2u3o9Rj2xCHTfcN6xCIU+tEAwCk2J7qPRMS3gODFSJK5Y8
LmcQK5IxGiYM0D3Xpn1c923oqEhVZCd3r2aXu1yLHE2F9ENaIf4OUmxTBqtJQrvOB93bu1CIDHFI
UWGMpREWnubY92TmDPICA02x5oV6/E2SmnF+sKqNeqkS48YRatx4g3F+N/NIkIe4ZDCUISUT7ROJ
IYofA9EQrT6cEEt60yT/dd15HIkMO8QdYXc9BNZCW9gaoZYZkdTpC2S5DzF3Koy/FwV3pcx4lLOZ
zZBD0avClJ6b8uGw+OwNOktYBx/A2kAmvhwhphyLDYCb51dgUDGoioJ0tCzAPko6EamRc+U4Wq3W
2x/qg+acQahTSNmAj/lNrMyL+vAboJeFm16OkNYHnK9RuVeYO77SLw4XZSrbvMHK17Dnn7C07P38
DlEyWVBF162nGnWBleuom8G4W2b8ffnWIPYoI3SkzNfw5Bas9OIeSIw8F8eir9Fu3RWqz+/K9Lyg
P+A/XncM2W4G1aGtv7Ri7kQUCSA2i97OWMYnFLe+dQ1rZB62Wo+2clg6Npl2qv7qeSek7vQE2ivz
XPWKUSP8CCYFB/s2aTgMAQQlt/npKkgsxjh4ZKYKszPcYtyz1VALLZsenTiUHqtXxxnwXoM4deOo
2OV5tqK0zL/WIdn61WmPV9bVIz02CxGZIqcdapx4unb3SB/x30Z8NdsTWOSgLDE7rWZ2d2QR3BCj
NLwa/lA3fUnDDV0VWx3Xq2fiN5LD5hy1VQyIoDueaBYO27ROtWzdtwFmSDviFA6VU/uganSYeKZa
fScm+vM7cKaFTDQBPWajIrwcmOxQagCuXzQrMcv3URL6C+xnGzkTQf1qwHj00au2ltW/4mnD0OJa
SY9V4mQm+M954O1OCxptNgIQS0rU+c/Ascht5CkgwSpOG8b0T15eLg1s2qKgTbPbi1cJsfCOB+p/
6tdFYrqzJzkRYtx0IpZ6VrbYV5m/sOUVw6e9vBNaI1Vtbx3cDRQdxXyToPUvIgZfxpIw1+OHNIWl
1NcQ7dP+wYqfQ2TEgFWVWC5vsthrZZkL97J+tWFygYVZD31rGRqmYhKUzQREPEttrCxgkdEZDril
rUfu0x7HUERbiVwnbyQHWr/HWFdupwP7Z3T8z6yH5b2zGeJMmiC7kBSkVE/jVZ8T516O1l7z7XvA
TnkMkXpmslq4ioGp8goWQK3xlaC32jfSXYqWi33jvhr+4vVSJTEP0frL0rPIqa+9qqPuzMrJkczg
18IZ92F2s3tfQuW7jops9LViwHhEw2eyzxuUv0rGbVPNQ8bWGJGkAythdUcYgGgihcvDFl7UGoDC
mwXb5brkrSltfaXtwyZbjYtkOacGe73oFPigtA9bCP+WqdhudKOq6bdGVEN/EQ8s00gTc+DR+Pca
ZUgPFeaN/zQbKJNEaLW9gqj5WpOgqkG64L6NC7VSj9e96MPRPrSX+k13M7PPFbdtj41rZ1JicVGa
aEtWUMBra3ANDVnsZlfa3DTONwlosz590LZYeFqxygJlOr+mKAJFSDxaD5lRXHFgXC9XB+xpHo1t
PbvqfW94Vy+i+9H4pfO1EGA9XgwAofsjfiHW3Tcf2c440JnpsdellquJWeHoRCgCedydAgE7s/EX
yxUOLa7eucmLA0MwRSUWAqxxdYrzt/OjoFaX/3LKZAXM7iA9Yy30pelTJhLfPCGVBbYhj3dIxW19
xnkq1hBNobumV9HeuT3PXuyImvzTT+bzFNh9Ol1nzHijhPyMXh8VBfY78Bqy4dFgcUAvAdGuvFtf
sT2RjTkeMkCf+hy3ZMmbnKV10oAmPLnAfOpqhAlOyOLaT0SzWi9dJwr1Z7xP2pvk3LVPu9tAWNZV
HcQK9ipEun6R27rElHPSsTT+RxCZf4SVliaCeSCR+k9Gf5CMWO2XhnqwG9RBgQjuvq1tRkq2JwaW
73VQ7JL5S9izFjkZCT0v+7XBaYSq4B3alN+UpfplwRtAZKgNwhBth0RRJO8G9rtbO6XPtLf47h5c
kNm1D8ylTKBeqIMbwOx6L5wgVH3lS/qbb/ktWqkwlQqoviQdiEnGP87BvtI00/bxi9YMLr0Rnh0B
VPgjU54L1+h69XqR/GYMlXAV4PQSq+TwVklOyHronAUB0aJ9EKX8dWca07pZsa1Micx8Cjv02fOE
WEFXUDD7Ag7Lz256wDegnV47j3kibD8cmEvYF1eZnHDmUhu5+IxFPZrkdCsMuqfgHTMBYwcBn86I
aINmgIoziG/zO0BPy7jB6+z/8ShUvmJiFeY19XH+GFfkmPFBhjbWm0p1EfMDJ4l1C7Aq8KcJIQam
/Htm/se2R19MwrdB1DGj+1dNwD0B3RoEE/0fVjmUBeGBXTftvp34fwYxhJFSWW2GSA8bCoVLPpNb
82Z+tL0QjFMzbrZzVnjL+ocIRI54WoHBq6IS6l83sFtfWkWrares8DmNAryOVcXMOKhybJ5ILC1S
srs3g9fBIvdvbCJ3cy54S7tmyh5aRZPauegTUvhUyNF3wSm93CQfL6Kr3sLW7YcQ2kPQ7FqsOQNQ
nRAFFJrsiMwUcKLLEAtvDtv97JthcgjQPBFpvoutpotOctsnPHqw3Pmq7z8QfR/lPmB545yXANJz
bfqfclrE6qFEsLZsvf73AX85zqNbO4EAbpRDATMa4Zq18xT3nHZwLAdTO0oTCBKF0jg2VoMrRYSA
Rg1j3ATAJRBLNkwvnvOKP8X6trzU9haVCKevYk77WwHSen2ycMftZn1TvP1Ia2ln6C+XxOsqshfv
naytwETwlthYk5lwXOmSW5BWN5upr5/QAvtjsIn9ANiJZkJPycfu/BXCME9AIgop4HmeUxzkp2hA
Z+wjHCqDNDyI6ciIU1XHuUoBFWYZ6rKjT8I2FDG6wGyk4w7Q3gUkIdaZy48iVW9PjBv82MP3sW0U
M/GSUrg3kRoSHLTJ4CbD2c804NQZZzp+OGY8PFBrwIIJdQIlWWrUU2rz/6cdTyAyAmlGESyCtdSY
oYc6FPfGtU5IjX5GuDDgAIr10CXefQgDnnp866pz/fpITSrci5A3cjXLj+DCqz6eSds0IPxXL8/7
R+RQXHs7hMMedAwmK18jUSiBZqf+N9F5kFGqVFvlPrQGC0LYpm05zF2L4UAqZw0tkMrzlaATfnmm
G4vENkGUZvHdGhzn08ccMxkLNztqSQMFNt8tCUrEL90Si3svVZa15x6hKRzb6B4JAEjgGiD7JEZW
su87bpS97Yjbq+15PwyNi/Y/6DLdzUIE2WZS/0otr9iYbd2J8GdI17E3He8wScfc5uQKhEFftbNz
G0UhRkMdRulg8EUAQubjnniAeJ/skYc51oborUFhTx53g/K7RQARWXZGjMaX19j8N2npKllenWKy
+tnUMMk2/GavYiSODxOssutdKoYLq6E5Zkc6g4Zwh/YMOid6KR65BxmhJ1co6ib86AHZTtsMOd/0
VzD5NrOvckhi0XN+mMUNJNdpc+P4jcHInZ3uJZmWqxh9UTSnZ4wOWOO4DSPcARaQ0mf4hcVh74OT
tmjxFIVBN0WrbAyJRf6n2PxYC8QHYLig7j/JEM3fiuM9hgKTZGTiToklEZ5yplptYyqwyrFNFUZ1
KOAvjE5Vy09wvf0xEeHRHp2XukGlJZc0CVE/cqbKYkxWt8CsrMJnWUGUbX4boj3WdALSMxFd51Jk
eXgcWD1+/WGRPpAeqPKtjvqdPIrkc8gdw1qW3VzS+tOMdt8AYAhC1ra0adstPsIBjliZj0SD5wxk
hxs3tl9pO0DA7l04mIrpxdXwtlqukg1g66p03KZ48ztf+FKoiX7ouCtkSzLO4MhKhbiTI0qR7XWi
Z9icpmau7IsSwuOjhkpHcOld2Fsh7WAH2T5jJhXEAVpqFBDoNC6/EENEutR57QX+nKomDwNkDREn
aRCJYVG2qq+BoG4JROgr44kyQPEUmfy91LFp8Ef8FijjBkyd2/rnB3k5S3WxcLT7wcaHfYj7fjMd
5qOVy1BYAg/IAOuqP/n5EnsBDaKzqB5CDJHqzCjfwp3UveW7HA36YHm+QvWWOuFvbPf/4ofjgQpu
KUjjFGakTrgbQRrWCflSq66/el22LWU8zPLUIrJXElkl1tV0/MUmWsOMPpFACcMccPqXIroySkOV
cr7R8uP//INltP5wlUmi4ZFjKyVmgTYJEoMFR9tsUhvrxJAEcBcL/EVz13wQiPFBbg+EP367m6zw
OrKtmJKFaDkP2toxQxh8u0NQjHZwMTNZI43wEkDSyQFNEgvCNVQ6WKj9f7DCTNz3fikFkQocKvhK
xo2C8zpEXGI9lkPLeTRfhnzWJyy+WtABMVlRkj29939bho6YhRH4ke66qwU4e0pHY0HRlA+knl2D
gqWvwkAkuFhEC3jKT664w0mipoHWVAI79hpc7OGep3R2pBbZTktTRQIe47MuA9IhAYCwwywDTO5c
WFOkjBWF/X/AHOqGzYggrcjDVoH6cu5uaL+Np0YlVHcqTIQGCdFY0V2ULdel9lKIzVSymn6lzLBv
u2JtNjITjmfuKa6rz7MWgFXzRYOJ4Lxfk3sshrXq3/XcyEG0b8nkTAO6hEQfiRaWHXAFbUjWHlHp
f+5/ZDAZZ5jNHYZDR4+DneGjlvRX/fvF3Hc/snKqzqKtjRo1kj8N573E4EadxnwzPzMYQ8n1p4cD
g2ma644UrfxuysGJwaaLv/WqbZoKrsZ8Ea752yrjkFCVgdxrqQIuiRcT9OXf/zV6FrHOafGrSAhe
DoOOJwsYlKnrH6R8iTLNL8rshMGRHJ6BtSrkvQ1/+qX/J6guHERBnGpLvync4CRKKowkFHfBC2Qd
nQLiSAKzt7QjGhi3Ao6l7QSEGA4hBO23/WSvRBsk39c1dtNn3l14KKOYBuA2FEGhKkZrAxns7wXX
FhCru9ED1VIdKwMAeDImY8BoV+VfgRjaONCpaSXGw1NoYZmxnLxeMIw8EeucGaNmZV11hLWwNqkO
CtzLTeYqqHZphQGEY0GSKtdDVAIcOBFfELZwxd7/lQ4hkcDHlfDE/+/gkJGb/NH8jSOrBUY7btvp
edZylLsS8P1HO+kqghGHDd7hKCKWFbNvfcyQovXHyup1gyQL4VKZBZpzZFZUxN8gr1xxh5d4JVHg
X0hnkMfYa5NYEISpON5eLYh3iBQLPIeR5AMvD6ZhP/JE1ZUhpWG5EqMfZHHLPoOMwFtgxeoQWOkJ
I2JQ+6NYUxWS7dLxLvAZoSOyXsrtoAP0aKFa2mFrJ3IdWb2XOWlj0rs5ue+jIIeuAiEmZ9CG6Ags
wjN/JeHYeeul7R4OeT/AC/47t2ADMixk8xahTgi/vmN7H3caQV6obdQwGylfDwHdeh5OUK6pm4Zm
887WozMeJgjmzJeCyHZigYYPM8ITO5+pFMdPg/2yZEtg73KT4Vb2NuSBdF3NR/ayaG/Y5VhEu8aK
h20otZrlpPnhswkOaX4Kagt+yxDatICio+4x+n879AMgszxJX/5aYOSOHCe5aOfYjA+oxBFLKtm/
UxCZL75AZdwlLUOWo/Qd+8mx9BcsNd2Fn/IQHmlFN3ckx33k7gwaQd2UEqhUgz5EI7WZ75J7GaK5
JfwLBn+N4+K6Ten8tfKrFdgFbS563N78HTKbKuU77kQBIPWus64YcvgToTVqRhcN0trkLIFZm1D/
/YOK0xcDuNYRYzB2llTjFoNP+9ifYpUxqhsgRnU+kqWK5SbQlz/FacXM1vj7L0N6u1wi0D6c4kie
sCf7x4H2WQWrg8lMjakCN4hD3GE8oss1W+M5yEKp6VDqVF3Ab/aWk8Am2tHZr+WrVF50Iw8BThvu
yjX91Sjke6o5zzMuSzc39fjTvgD3whQSq0IAwYE/zEeT0mvE83JgpfNrCECZdcYlGOHwFyf6OmSC
gSRErT+20FDgAkyBq3HnVjiayMwGc3yZ+r532ZksGKgDbuwbHi4S4jPR/ksEV1rmsFxFWDvCUKHC
xa1GGlSwHswjG12gwRpYgypJL3DCZRuVT59mXc0t9pSWPV7xB7ljjjNP7Miw/a5BqLeRUZ/0PoAp
sNz/SBOiWQ0Sf3827jI/tUZ2y6ck2Q/OF8JDeaJgbtB/GHTC1loSZk0Jipkb4lbzOsp+/41zI044
fGnycj8Xj9QuEYXbR0euzqWapktPggqpxzti5KPz9J38W5gUJgVE0a7PMsi9iBaMh5+E/d9cQLdZ
ackDyW5voP2bM/0tVAZfre/zEyq1+gFSbnpiQJc3HXwK7w+2oeuHbd1orTUQex8UYWav64prIrW9
vHCNumZqQWl/flk4JIu6o0HSLgzyQsdJjBjtzaSGb5UcLu4azmm/Tt7K7itKXq/9f4iaAlUUDHt4
amHFDSk6EchrAVMh4tRH4JQCDW+xNdGbyU/uEeSx7M281SKPAJe6tLDn0M9yxaIbOfJ8i61+o+H1
Cv2WLw3NdpG1bC29Ir3SWNA+AuFyK8dR7CLSv/J4Vxt3+Do3YlwDhHvD0gDK21pI497jZkPdBvUh
i7Gq7eqbLX5ZNFEWKScuwBjxTmnhf9sj2xP3+GulupuCoI/N/SIEbMvaj/CpxdUVz+aG7yhVmnYh
Kc1F/nHqpRJajczr1MOeosepqpiwGapXlm7C3yCcwEmyJp5QWCfxS2ybZL49ZDstE+vqGd2RAE9N
45Lc5/zsn8CStNeqh69YbK/ZJDVir78JlOgqlmB7KFGZqyeC3O+8WawmD0wOQarVq9skuYl661oF
IOk7CDeAQstf+PfqqErbqaVDILb2lwAa+eiWBlTtGS/gW+ya8uR8lC+5ByndCsxxajnDQ8cWOQ26
9HY+rcZCy+Vbl7w02JpBR8dQIE4Ffu7pJ8bnjYQ2OBBnGB8xIXcl+yYgFAhgFT7hioUXlzbKZK6+
kUd9Bt2/0gjXclXrPAaeDKSLSwobo80nRl0wOiaOD1RKaljwRMQy6gurrd5MaY3+WOcvUDxyvy0R
+QXmIS7dhkAfLI/28XjDLnPcN7Wsqh8IxOBLpBtuNNpS4FsWIMN9Lcoo2CadMM9tStB5eZ9ySpr9
Vyl52y979hc09gwDPqzeGcu/+XuY15LM29RqEwPHhL5WtB2UHLGehTy0g45aM1+IaAf9FRrnjJ0N
4rHjD3pM9gPyW2IweZjYQzjwRpuCezJ5LUy5paoRSkDxlE2pRXvmTyO/BHEko3HGk2UF8kh6/Vvo
og3XkfPqM1dBs5RushCWnh0dgwsW9mpugBwlS1J1onX1vmdQqjXuamwA+jLfOcqT3wkJG2nL0NYV
JZQWb8vqS6YoNk3wF8JJ4MjfBXzAteHi51zrYXP5ThdZY8cYQRTJ/MYfGheVod73iJNtORCU8Wk/
xMJhRvnxP4XKkrvm392ab5Phe1tt2HnYsvsCaLeiQIJg8r6rdH5gGqMtN4Wj4727MqhTbHRsKjGo
ojzhX74vECI2SsJ7h82eAQOogR8PNEtSN8WSf0DPy/7dSj1WP7qXLepi4MacQx7sxcT+hRPBNn1X
Lkc+rJjyewgnl6RdcTfCEA9uSgz/Ti2Xm+izp/yKWjm/M+b/9NYVusXr3rBQPGbErwVRQ3W32MQ+
iTC/dYIse07Tvadl8ifHfzhCU7fn/OOqAMmz8RMWtYAbGZvcMqE3rvliMTc/L3sVx+gQZ0KUs5X+
pwlzk6sCTlD/pnDbscjps79I8KDG4morKMA7Tjz8OBXKPVakbPS2g+x99GF3heomd+n0NZ8xjCC4
ZS3+teRqG3N97U/PRU6Z37kPje7SyRzkvDLU13Y1vHbXoJQeHvBz8h1v4IQkvXj+KUYUqFt/bL3a
U0zJshfAfLzCHU4a59z3Rlefgb6VoNuge9BNSWrbO0HugxpuhVokeWqmw2gPPDnGxqnIwqvFXInI
fUl5cHTvFt1+onkd248Ci6ueIFbB+GmMZDQMuPbgTNPDqJguqZjA422MSe7OFm/1EuNWJZpkt23S
c4FEEXackQnz7Tc8Nh77C6vgUO/XlflcD4zabWUKTZDfER5lPDFjN4PeLKA2Lxqd6lw89Jjiy4Rt
aa+vq3H6w/c/SM525kewhxnJks7naYyP1TsJNL4ss8EOa/gSUDUil0USpk+ddNLk2TFQs+C/ziIZ
wPwG7iPcBfPaF5f3PDHSOpiJS1jXx3r45Q+KRB1cvlKu7u/5asYVLYUu+p5UblfaxA020qt+Xd9I
0kskIaSr7ow0e1EEkoOH9hzNK+x1aGeGZ2BtwR6CqXOxMRfBPp8xqcD1fXYmxTYEWHTcVIle4mmB
Ueu+N7MX7yqUXj0v3bEnYd+57pWDIFkWZcjIMo+CIcEoT2+/WKp5zf+haQeGsYxMt40rIEJwV9V/
Glx7bEXrcp1oxPK/H/pgaAGGcrD+nxzv/fltzu27mcm5C0W8HdH6iQpTYLnNwU7cJiLvpTFuW5eE
Pa2vGjyusLygnR5aB1Q9ppy8r4EYRurIiYMoOrXoC1XoRrHoIvMl4+9rc2GPDVPdI+dPRO2VyBs+
v8hDfPWZcr/PnqIj1ZNFG/+X26lQAAg+yRK7HFh6r1GIAZCTodSRiTCYUELCK/wWjZBRVHCBCUBG
3rb8zPtMsWD2QKeZb7wgIC2bRPhPE8egqL3AYO9MdlnTQ8a74SKSP3LM243cw5GpztdTuJNGn52f
nxem2cOyqdbTGmTwW2CLtiJYoclIRNcMCZDdoWMZqSpn551/kWB/8kVgPl/COTHE69Z8jbgrpH26
SLZB10huric0Den6SOMTFGSK4bCMZ6/XgzJ55SmASWBi+VgrewHX/sU86L8hBl7X66lskLIWhSp7
MCZYlqdXdu0grbrr0faHBAUMrnmJOupyYnNrjSnT/11AY+zo1ZGM25P9AItOli7EvZ9NnzOo/Mw6
wbRoiiBK5es7Hg9xI5nLIC2mxs7pU9cvevFpN0c6j5xUxCc315Yp156QJGediIIz43bDN+VivIhI
rGszs/Bq6x3CpWCu+j3VnRDDg86p/v5+eYelGas9XndO9WtQ+tairSsyANmg+zwsj6jCnIUzT1Ju
vj8JA1vdBnxz/TZhq1x/YE4+TyurQaU4Bm3cDT6Bo8YfuLm8q23oJQtnSpJ6xkAAxWK2KQara88g
t+CYSZ5AXtZ84/v5ieQ1E4rEbuarF6386JmzuKNin5Kl/qo9O3QeTVRZych7q3NFlxc6dE8I7Agk
7HqWgfbB+DYwuH4RbUqaKh+yANDozz5iSDS8B9ODN9zf3AsT0jXivzbc8AaHQc+dPOmXVlR27ftm
9yQHpu2DeylTBdBiM9VTCnZ5jLJod1LnYQQP0a6is1JiWkOdWa67O6cuWS+8g4wMAHuDsVJxuS5b
Z7Q1Fkoh323Bg0/BD9eQwNSTDFLXSZ9ovKjcrzg2wO0yAEm0bK/sSB4OVJTcPS7KHjssXnPq1Ubi
zj2RxYyMdyF7thYQMC+3aeT7nQuwP5xQxoo0ZtuPHC9IW7ISTfQ/ewIzYI5AgLc2rD9x1XFENwgq
apllkwyjEGEDFH2J96Y04FHuk1TtohTb3/kvsBeJ7s2i2kRTXXwBsKSAPcw55J40V1O4T27PnfmE
b7Y7kAfdNJ90j7s36IBJc7eZeA8KMJ228gF+/ZKKDAPBlb0k9wSfc06Lkx1NBBquOsCCklDR5CJm
GK8uzwvK7uveUzZrnMDAJGY8gAj9SKqNOcdxI/pEG7N6+4n+Aa5kf7D5rQUHdC4BOdMy+FpDoGQf
UzI/DzJqcNc42x9Dl7NzLeGCnnAgrkQrnpKIEPmkfnRP3GL3z1RrbkI4v8IrCh1Ni12Gnx7421qk
+pWayyWn9ILI/YSX7ITZcpR/SUnAUiif+D9v4eoB2F5O5W+DrR/qBigZ31vl+fzCOKvE/eqeiuVC
CrSGeLttb7RB1mXhSnGB5s8MpDHCKA4nV1u28fvY5dEE6kxXj9PAukV/E5dfvyiLKpwvbSp3AjmI
HhmJG2LV+CIfs/X56EeC2haI4vVqJjQI6jZ9061V0xFr5JJo1ZcJJ5cnv9O2+KgXziMHHl0FnZRw
RlG2DXkrvD3y48MwBuyD31QkMrpd34iyKq/sjrn0yERubTHNpO6K7Wgep7adjgC2tUtyB5CtPHvn
QTRqitO8foT7IzhY1qsrwGqr0lnISx2G8OT8LfFD+2hi/6Rb9IAEZoxAXn8t1A8g6l3vjK0wmweL
IJOvxu8DQj8IxC4cZ+cxAo4BdhmQgZ+jAt/IN+FyHbKBrIjjSkxWs6aTi9qXoowRBrK5bVboMdRF
VBj0mlDN9pVjj0k31DftXhdcRqE7D4fI3my2+mCDyVPexIpFaUFGwC+Wf2Ieh7GrqsdI3tthnOkT
SheWSTwKA33BM3ucAE0Md9UbDvtwse/xjFA59GzdxCo47QDUOyQXalNlwChGBt31Cg4eg9r7kZRx
FkHxVCwaDO79vma+84s562fv5HVyPT8e3tRZaSAWA06J5wXKKw6V7qCjaAYEP1GMc/lHn/6SZom2
jBQ6cNBY+IUmOA/bP/RluuRP9VZkhXybz5XJUS/SNtl7li77OZuVm+SyMu+H7QC5XLy+qTwagLki
eEMpjcuxHOwrpFswa2nuKR1g3VzWvWillX6aTRakNzXanUYCkCnL5MvkRuoUfHfgg9NAon+M8KL2
Hn52ICvFy4lkgKqsfBVK7Z7QSYm+sq0ZwinpN4I0bnfC1o2BYCGuXmoDr3zfiOdMDygOFPQTFUw2
lW7FEGiVcJg2OW3RDrxCEN3mETo6y+G/jIappxkTrkPMcF2aeImfYOv6C71ZFdiqrapQZaV0hwwW
wn25J2sD2O1EI8ingo6HDGE8WkUjvtEpfnwRWiwHcyCI7gMD3YKJtq4TuzOdZRKbP0XtNDGXyMcN
HsLScQ2PSdtfjMvJd1UKchv7G3FqaP9mDQjXfYVH6ZR7hevpBKF7xd8ZC8RC2CXCzUtn65crIDEA
aUIKS9wME07VHAyLsm4YoxsYuRr2tpvpcl+CNyNhz2i9dpDpRM176+bd/o0Io70IGcNUirPo1U6a
GN6+bj8Iu6MHjjh/iMxnBzR92HGPXHsmrhi/wSxr+uZ0Fxp4hInR93A+M7/8uN87MCxBErmT3Yn/
iNzMuDJGcRvE1d1mwW6XCEC20bmdaC00lKsu5cwliO9xw1ws02obkDrqGpsGoytchvjFYJKOLYKm
WOSydR9/89bCWnrZpLh+rz2JxFvuJbPdiMRRLrYjfsaAbX5P02+xNeDnsh0jlvaNzh3qJTZmP05Y
IJ7Mia1emRg7qioHZaSZqJa+em+EQINCaJO+mifvOUYuhS3u9BxmehMtCVezVCqKiIuFZb25QmzI
3yigz0bUHZeqADvEUqWxyRs3bwTMfiDwEgsJsBYYzmF2R1HzWTnVCn0vX+1ZehnZWdRQZwtViq+u
FLpuIkxEwM90JOYMeZvRuceTfsvDRsLmMCU5zCxUL4L24GpNLzO6P587uNIu0JONV/DVIscpKB/u
yWquQv3aK6kTkpQP4wI8ONjaSSGnbVfCPV239vZK+yiFBjMUXHBD6+NYCnP7LPBspGZCyJrav5Ci
+uVFqwpPE6QIRvqXVD6jryAYWoxZzQeu0aL+w9RovTXqM+nUV126JPFbLNpe9l3bvSRUpTmH9TsB
Q9li0cSboeQxtRnneD0zMZBAWM5hFBJU3Yr6trvzlFMkJptQuZMarBa7gMV4EpctWGiLiuVHSHBg
hEr7Se23h9g+W0jehiVjzv5JiUcuiTbE/c9tHOpHNKP8fac1nV6DyJh6yeBTkhcLf+JVmZJrb0Oq
IVHHX56ivlrrufx1APs/tJ/bjJOvTxkYVHYv2GgHixYetsviFzDrNPkU8rT5mbgppCtCgdry3HQk
gAumXPK7jbSe1T4FE1FXsFVusR/30ESe0ydvMDN5EYqzILl5fcYFqsFC8Tv1B+0/m/bXyPKlQWbS
VbMaxztMTVgWis+nZRDliRUbQb4TLpeYPYaRTE6oPHwP6+7/W4oAxivMq59/seztFUWaoxjzSjK7
zDiHOPjt8VTYzJOTtMxfK2j606n484qv+Mmoixxf+mkP/GLSCjSsxIbNHbH5VhOfQ+2d7CTr3ZRD
ojbOubzsOvWsklB0G1eCPcGHBNU2SrGhkfqmxg4+XM6t25bh5F213D2aaled+MhihYS4aEdT+75C
dkMEXfqLWBVmaagJ33JnpBLV+Kg/a47HUbNNTV999DnHwXa5OADHsfc8amVKIRi2t1MCmbXormMp
Fnu9hcHfGsxaa7fUwspMm3IpMKnzGEKEQ+Wao98Oxj+lyblYr9RaMzzW7nCGfPCq+UgZQ9yf1jwz
aJ6XF8SFDuhIw4NyAxzihuAgqHEeAW3uLcRzL0np+pWSMoUIAILCqBJJ27y9Ga7q883s5gxsEiqL
B9JB8ELTIskU5D7cqNeMKJBwKTCPRR7YhAri+e6zho/ljicxXa5uI5/OJ0K9y5ijYLMm2B+BnYFy
4JXSCpqN1uusw7UBK16p7FWN4mqvW8HXmaa27DJBaeIEZBcBB+zxOuckpwtObOFR0aZ4DrpUZP8v
2sS77X9pALL+z+qY52G0FJj1VFt5cH3HRgNh7ygl2vSMFg+ukqur++UNH6ViOqFWvrZJ4V3T2bIn
5TnBb51t2bFi1qedubMk3CT2vqM6uOVu4s7uJ5uVIQomlcl9eRY3aPLtE8Zh6kO33TGA3e5whrY8
43Ly+Wm6dTHiqqZdTmKwY0OqK3McJIrkWbkbsDrIyk0wy55AApEv9eSWqnHb8TftkZXxy/azB19r
BcRoFv/PAducBYJ0gt1/Y1J5Cuy3FPt/q4mpjve9LarH7bKomr+pKHaq7hGhGxPGI8ZPyabLbgvY
3+ZdpJmmVpz/N3RH02im/hMzBb3Zb/VnS1FvB3DzHSmZshywZ0SIbjWmwZjzkPB55Qb5WB8GjmRx
QwcCHPOB5KMNd+ggDjMm6OcZ2HGC7QfGMN6AwkJUGzvNINypJCKeoPM0U/Jbeu4enw67gGPsiPdP
GpanIGiYoSLSwSI/xEzo19fcQuo7t2xbqcMCQOIB/uCx5QI7Q8vVkUOUlgSOFCR5hcrz2Qbe57a/
D/jdJ5ZEOLZfZwVIAqYt2aPdpTm0j/rkvr7ePo9SRz4UP7FQEIjbzqHudNcKQrMhKrIhm9j1fEsR
hmdP4oZz1pS0iWA9Df6+qRGC8B5l/YUgbI9Tq9WRm3vuEJwOoNbADFe92EextGs8+Czh+SUrcJFy
vPK3JQa2EYWAb6HD7+1QeB7uPazJnB8y+fQEtSfn3rypZQbwz7Ev7XtNPaH73BrJ63LE7fl4bLXQ
EmnM9dM3x2JrbCiC0IRJ7ed8lILMpZQgIHCMZlJBOvTcc5gYX8G2gOzHjbYTws7279FRqIlYYkqq
dqkUMfu+1BiT+45/ub8Ec3k898aW/Kw8DCBBtn91SX12VBnGy/3D2uQFAKxEbeE/EUDi3XNL4iz0
hjActbHdhUbbTeVsCIQEQMlGYw9HGTbIwpMY34anT0JMTjPIc2Edvy9hDowEiQ1b8NyvFWg966kl
zQS+xTK1XPO4lD9cMBWtLIihQzKhV+z5Sqv/aYA9EGBtkuiYEx3PvpA/6DiWc7S5OzCjesF4OGVw
qsm4G282BWzlHPfKB7B7UAKSzQoD8D3Wz6o4ugFn4knCzXnt5vXxHoWpPI2FRUxsEwvxPQ7dP6uU
/HDUNbKAkgf5rYFFLi45/PC3G4nNg4x3qrOCWCAWLJsUaFKwORHvW8q76oYhiT5tMrUkm/p9bhAU
NJc93fVD/hMMG36YGYAkb+P0rXQ/YCErNWD9bE0DZihX6WCIODWIQnlsB1B+N4hadQmWsqY7xkUo
5QLiGIWLJle3OkH6KLt/Xm9vg2pUYgCXSVIJ5kBLmRgezhVOBinwldRU1ABlDMd9s97aKETDWVcz
5rtlSkiTlGHfM/01l9fQoaClDJ+SVNshvKMZaLVbNKwNZBVIcNu60zaW1xZzuREFbtpYqol5PXmo
Qelm3PGudEtaRxn+EL5zC/RIGbli3R0oJvL5H74sB38v1oagjJH41fS+grMOgasnMlmfYbV3ifBO
K+jBkroMeE37Z5w3NPbAvNBa27YMN/tmJsj3VPobO0pBxNHlc8duW9idyrH87t2e3mxNVhHsDu9j
oH9Igxg8PIWGsBvdIaZxSt08cgiH6iiPLLZHv3tZUrQQbAwZTeO7ue69jj6rpV7TQ0VF30zA+Nt9
ZVDxb+pgno3NNobeMRwtOS/RZzqcy8EuGrYgJYhcLZBbUfEJexVf8HjB0jD6pdWKVDxCD59ngkOu
vs0AYZw7TG+h3d6eflypHWYRUuvBHegvFtwjJlal62chdDz+gkudMKzm9L+32mKcwdDFUJUnopWV
Gavo+Rm6F84X8EW7ucu9Atb/kBnJLpZnJnBWhVw6b7T/aUdqX/yNBu4K2n+wxQswYhvadDoq3twx
p+AZBPVLvuJxBP0oE4Th2cFOoRniDKi5tbQdEVwRx0p3Ux47PxhGw9swtDZlDD9IQnJgjhb+l63j
28NmltKXgPvItpPZj3kLhFx89MyewiUgchLgu0rWsyUY6lbBQlADK7trf8x7CFlPy7clpThU2H16
QgRU6zcXKbxq+KVJ4alluNzIQCAQHxuJxq9igqyXDWNY04UTLHT2jnuYeS6Y3pKeOkU6Q5B0oSUn
S2r6dRgYHdEr9Y3ZF5jmviamz1KkWFiz+DAQ4i61QVnC3MDC8uy3N614Zqr7acASkZ4ZVGwWvJKg
kmSUZkk8v/8HdQc7pTHYfrbdbOL9EJGNnu5A76bhlMF1NIFNsCL/ddyNg0s610Q1IFnMlrkYg9cm
q79i+X/k0TfumPyRzMnJHEoEvnxsRE6E5PkXUwF/DKmNH9yhQ9rxtBYbRv+s5rj8Eijlb3Xxpfy0
umQGkBbbo7fQm9JRPV/Bod2AV2uOW7l8jDcytvPEXWF2tFLs8Bb4rF5vJueVT5mBGxe3EEMVdiXz
urbwSVKvrDoiSfBzOmLO51i/om84Ay4fNz1/z7WFJ+KjFFinHV9UgW9Gwbo6m9ZfaqKsT7nhDOUz
DBkn0hrlkI0Hjo642c1/KLkEnJTFSnzfvLLwAgSj+3UN87fkQkpPnVK/PT0NHX48bkgclmWziixZ
0QYEGljPqgflZImnhnqsL5atg7j1LqFSuqquJsLEqpO/d0SCW5zlsg5+oYFbknekNSVNSl5/C89V
ExUWpqhemh4HSzCHtyPwXn1Z1h6WRFCyJ/FkFr2MZhg5WtImc87BfvCE3ceXEdXjHV8cHMIABMex
1fbF4VyV5J6HVvU63hG+Plvl117zk8BK+iiCpVhgeVh3Z/J9U7tz7aje5J60o9O4Fn6yxyZ+OKMz
JcEsvJz2MUSOdBZ7/ksGjvdiVj/T/4Pw4zqWvpywDqstHyQkO2vJroVK6EYB6DF6SqEcjAO9t4CB
ABRfMfC6Bz1bKxckzVARLju+yXJgi31AUPqrVA3aRdcpH7d9EWtuSUQrnMd+KN2Xpx+9ArF+SKhP
grL4uzP7Pr7hXPATG7GVDOKtuuYl6uXxGMMDf0/fixZBKSzinJ3GNsvs98HfsZ3vLKysLKoCsNlG
xsL5UFtxuvgRaaD9F+UUKh6hIi/Eehs1ax8fXAd6VPnTTH4ACvomFzEo406unNup85jQVkMda+Ot
KREAhIW9hvlhp7Vwza7/3bt/e7fCAQpkROMVC1JMcJAGK8L0GUTLjl3LvHExMi2yg3lDMzAknGI8
BvSYy7+EHFPojGIEzgqVEXI+XZoiaAJoi9w5rpn+hkiI8IpuohIbCXaXqNuiQy9TE2YYMOngLfTY
jwvt+ogXYduvuXk+t9OVU3eos8JcyqXuaArHUjPoC6RsGNXRhVg/3zqTGECN5N9mfZtFY0ZpqeHZ
UrqR+cRz3ZDPUPt/y26PsDt4uRt4Sj0DSYuceHbSW0uvreE/X/6ckmvLTl1w5vEvo2Yn9WzAZ1D0
aUhxN8yZHZjGXQfyh8DnZTEFzjy1BxGgNXdJvTXIM8dUlp43LXFrGB4Qn4iv7fUFPmvyb8T+ZgR/
iip4uYB8XczTPh84K/hRfeLXn9g8jr46hV41hVJtbAZ8H/eGgApvmJmx9J54Exn7cOt64Y5tggHR
7i12t3/XABteNOuhNRiJMlQQM+Pq+4N6ssMDViUsXfjUum3rQ1f00Of+iQpis1KSLQCuVS6mWigS
YhI9UpjjPYfJxBLDlMspDChGMmam4tvQBy0pmt4jQ15oKapSyYxqLlXI9MGcX6HL9LeTvSWbumYm
gt2GbT/CkNvvto8J8Ge20zKJGX4M51X1E3DRsgHDrfcquKOTL2rp/rGY+xgTNrq6PRf+Vqx5NTSk
23er+cgoCGUlVmBG0n0pPFRnIywVJWYrtMyN4o/MFZ/jpPLWtE1lD1C+ianKzMUdp63P/JS0/RzJ
W/TAt0XN02bEEB0lIJWvXAj4LpfzfxyU3sISYF2YxSpt080oZfqwANbb/jVeCZevECKwwq7IGDbO
5AspqYvdnAjaK2HL3JwxcIGx+tGToSzkgrxkygdOOlzrWE/O471RbkmperH3rOVOv7YF8D7C1Gsq
rxEaZDiJvs+ffXt3r+819ITCApX1vhZ776Tvso7pSiP6K1qKBy/wJVOP927rSbIKKmJsnFsiLr8f
ijy+l2GScxRVLh/5zTiJi4dkQwyb4rAe6CNXbLeLpqy9Re2lZv8Fbnw1/Eh1pRvzARIhxmzcZRd9
sEilrUMsWpkzD8e7rQy6K9d91/Ja8mV/N1BIpCXnazPcvevJmKtxQwV91Ae2wobFXLOkE9KW8oUx
OZbU1H8L+rqWF7jQ+HC68RbtXrhKTn+3ImG+5l4fJokSYYls4DMuyfY30HiNjL7EflmCKTe8Sgfs
4LEkM+FZWYpVgOi0kXKv55HiIAWw7bydVD8ovHhgFBA96cXmnir1WWAVBPFskCR1azfC9kL2z5nq
tpBoW/AExPZWvlM/3lNUsbTwy0fyTYjwRy1ZDKrnT7WaJNnNpmxBMpmU9oiAzUw8ddhP8uX9njam
Fdy9LMmhghZv+hx3pi7wVNYZiNksJVaAkx31WhpX6zfhGBRYk/VLA7CII8+tHqJ+ZXGNTC46WUZd
LjXj7FJhWRbIZx8UuyjJ0us8PR02AStuktTDcr3GUdJ/E32xVuR/T9Ju0LLjUVmzNP2p916CijqF
9TRHAmqjyLlPtBZOMuahdEY0zt2n5+qApx33tu+nu4hP8Vfma+IZI+CquAXj7sPK27nrChMu+062
hUuDzbljarA8lGNR+7iImMA7esdSh/Hz7twC0q6TLyoqagqpeb4SOkrIDM7a1xVCetiN1p4F7cJX
z76m9BlGPz6B16CQxD553Kxb6cqsQV2MH/ca4INCYnInB4M2qwoCcAyFpG6mtLUMZXNDNle87y3B
FijDk0sv2W2tKmXFB7pc6b3dV+B7zI7Lm1jEWnK9cay7zDSsW4H4PrGKDzXV1rWJEoKoAUojEivG
3YqH85ZC0gqH423fwPHJtAvY7LCZrAGVs29tCk3x8ArpAktnMd+/lQGuFoaAKtpM5helRLntUpO8
ARoddekMV384a19UE4ZpSd6wfSwpPbq1WrfBSiGqyvxqS0ULKSuyATo1fDdmOrf7y1sv4GfRHj0B
Z6JO3TlmFoQiJPq2oDCSlGfJGyowVLHptcyxB++17XVU5Wz+SoQRSLwb3FoOcM/AwrkqvqNSclLo
JvrYKu48aJY9AghxhmkxzOqfHivomaaEjC1a15Qf5hFhXgUsv/jaAzqSiL48NlxTA6V/TyUOxvsO
gmvQGaAfUX+AWkgsuj3XBRZ8P5AD+EEnTHzVGTdN1eZwnWgqhonlMkutLZFV4zMTZwGxLNcCjgE1
W4rM5Os2ugwon2dM+GfZmOD3PyAIUVB/cXK8j/O8z/lK9+q6lsFjyWPtyE6fu6423A6bKk7LmQQT
ki+dB26sK8/qpFnv2D8Waw7BAf2bNNQjYzqT3G8w4PjvZTP7EaIbQpZ1U50s8GaZU68xI7YwC0Qi
qUn5QonV0gt0Osq3JPL2o98CtHRIiCA+Che3dchgbJj7TeMP6ZCAQgmjzwj5FYbdEZG9hepunTUQ
cx52G2NB9VsaJDcCtHy/th+YXp1IT3/R/yTtZMgdhYJzJMaJPSvr23d7INltVRi5YyAmB7pFXbq2
H87hKnKhhbZtuuVQSAojnlid36akVz5Wdorm9RUcohjLV/Q4OxJIVsq6DucuLQVR3A2FFK8UNZDc
nnDgvZ6TXwvQMWsxNljVmt1UOHqk8vMymsepiVNM1cQnz5bFSZmqDWt1MtSBd7sv6c6cc+e2B31H
+QHKZjWW7cXxzNLCVM2yFwfdZgyJ0YnKveBQUFMikpGOS2iCOw5X08Q69l7Rd3n3b1LCd4vSmAt5
OGAZRFSVfX90cLpiwq5sb3sal1zzIyOIZgk9O0RyISoz/KN54ynQwWtTV86RxetOj3x2d7eZBK09
hIi/OiN2nvCfsZHGXrLUSCbtHXOP3CVYOK8Z0OojTBjUkBqVmFu/lCa7vAhJ7HC5ZecZFNgKVeI4
tI9Vc5TgkA6hZW9K8UYc5E0kPKNgXBYT99BLkiiiow8Oe/HSjKOCLnnv0Ue102sckDdjnPgFhRJS
tU55VydjwCIDysRgNkgCUzG77JkuhWKmhNXUm7YSCxwuAfTJmg2Voq877QPsF1feo/4G4vKWd3/L
1DwZr7bQoth5yA966shZlTQ5aVmev/agtQLWN8Mn0EwHGqgrnQ1rFsV5jpnoLFEtMtiJp6gJu5DK
00keDP8s418eKboFGl7KZuDEofTNReZ6ww57yY+pnsENajBeVBgJzj0eX8B8mbA3O7aQOW3E6T1z
iorwb7ds7WBfmKYfirv5ODSYdlmyo2MAMUeQ3Gb8httSif8bTNZGfQR2dGxjsAMZvuvyfG+uZSN1
DyfnyCKSjsKsX11uQk8HGdb6LkVDOoySO5l84Ajv+wlfZRolTAZNP9kmD8Nj4GI0sc+HBV9k103g
giXFdABLVvhiecFO9kzq1o3utyh69fyStDt8eqC1CsdtbY2dPoFk4E7QAbPiH6SiI9dCSIfcCJFn
5QzO+/InT74zu78zGYKILHe1Lr5uhJWBrxAfb4/yFfww6R1rYWNTXeMcEM7LiiaFLq2OnD+Gtod4
I/M1mL5IX2W+8S3vL0Mp8xpHG54T+ZPWWf+vaFPl1XfYR+NDVHB3nmkUrBtMs7O1YmqP3KpoyfDp
ERShc4hZDEjSDY06Uo0taWkEaNRRMXHX66cOedSBpcVYIHryHzKQFVC6e7nOp6BwZdTGnL99/6Fh
5D/uOFYWQiouYOy9iCBbPMWoWGCFODHMW0kIUb1CPpKd1Czc6AoHI1h6HQ5LYAnnntu0PtLmjkdL
5WhFuBjcfGG/NQgYvko9jhHyk01WvruBWgZz0M03t/dLwtCMDAsklq/6N55PqX5P0T8jxQ4rQM2l
FQAQJ6Yyt3CaYn5hLtJvCZ59AfCDqk4AZmJLkhntNflZlpVKm7251vBk9uKc25uktX+oKU5PL2lD
gQR3SQcoDjsYcSpXhXGaJ+KbGriaqb8u3l8h7iezx/POhk+6HjfXPgOa7HNJ3LXbxkQHGr57aew7
sfXN1+88xz4ZtOyTkREQtn0cxamVPYbVWOVPWDH+kzaB/EbV9O8r1PhZVwhECZzpTHrRN5UDSr3Z
C5Yr20WXG+pGwaCNSVaDj+vaw2J93kSeRuA+d36EgDjBeZj4reoLXlNMmOhq4mWa4zoCSpTmtLx5
qGNhlsc1z0tWM9LKouqGrC9KvugmK7N6axyetYq1OH9lZYykwZOHPjS3iGX3900ZziUEHnyvxSli
i7eCoRdjNQRxScz0LUkGgbgDW4VhBQuMGXHmrfLUiYytN994JN7HFQvoV7HJdaWeHc7SSCHd52ge
ZT/4WkuS+4CBrYTRW7vYoPglp4rHpW1698d61osxvfcVMOefKgo4STdUgyFYU2CpjOVnjK/kkLWJ
5a8HYVfQNjYR2QfHPozAPKcci6XTGiPp/mPey6GO+NqtAq/OVaRP75bJH/e6qRcfH24Pf+ctdVVg
BvZSTi77L2hSq4WGU9q4/5WgmmljelpI6NmtFL2443Xf71+phT5qmV0jWgTEN+6NyNyIn8vjQ6pk
+lK6VSCUnjZChNsvH5zSboVypaqA1PCDZjZq4EXmqh6S0CW6WCJYEjQT5UOyqLdEOhQ8RTqBrxv/
sbLFvqUHCkj2pjReWMkThQkx4czgmeXGQUaFQqUVQPX7bvzmQagygnwhyibwWuCY+W+JqvB5vKug
P3jP14T6K7LipvD3K4XOg5+3xC3K4aBH6hggnEC9MUcwC8DsnLBiGnyFj1gsbC+He4N1CjFuFvdr
IveLxTFVaVgMc584U0y9e/cT4L9iIiGDK52/eQg7eBDqKACz9FFvJE4L7As4hGqvj1iXHjAsm6tJ
h1nymWM4M3Un8EYl+NGO3hStaPBI6AweUIyntqR0NkLlIJavTc3v/9/DwP3GWVrjjMcp2t3w6M39
lonm1OFEA6iXV5LCV0JLDBBHgsoLk5yChcXx0VwssUwlHXVfkp9O4IQqv1w1yvixVqsqytDf7Y2G
yCGfHfl0JZ/yjCbYcB42KCrsKIonWLrrVQx+uFAt+PNn86h45dlvRI+lJ3pEsRCq+vQglej9VgrS
00ONyfrE8zQnlULLLN6ZaUbk3uNLEMjFp+Jnv5TSGBfL7+6bptfD+2rCdA93+NeO9ZbQMp6eQqce
WhZNBcNla7/JSRf82cbhjy9sEH0f7dZZYgLKM2UjLj3TK7U2BhPXakXw4nVM19PULatuqBFW7wDq
ttouVdHAY+lfGotBnUAbE/9JtfelAUWzpgP5hICG4irsuKxJraIH/hBEq68mraCo7yN6wqj57q5+
3X3dLpwdvHlEwyBv4DUFd3Yg3GN/q06X6HP79LxXX/XkNAgqARUH+J2RiTFBJmtYMQPvvT/2MlzU
a82dHQn1xTXUmRyF8k/vwwyVXtNy1GQYsD9qLPE7z60TFmlSZDqshfdCYm4t5+Of9ADjf6gMnKvQ
oCnNNZ11kul5krmdcm1DDuf8kQVBRL/teUolR1gsnrHSyYu+baknL19C8cNBy4SwTHBJ3AF63TZz
9V1UAYh0VApM5Ni5Mr0WMnhbOOT+Sj+q62TtVKeRWwmIW/bsGzI76pqRdajFLmDlxkBJ35+5/aLU
XB/cZMKNbYAGnt7uqpXSawqx73j4a6lsm9UKQkOsTmVOkJNuHPcPQ0DZ4i7R/z9ZRtNGkybjlELg
UDuoxgVSeXXaDF9MwLScghYizQY+wWRWmvNkCFstIgAZ4Hr2r75OytKWnu0II2Qjz28CFtLSU1r/
4y6Y1jC2cb1BpsyqYR0BkL3FHZRSwNFy5px9lcJNUdqsvkPMsBNVCbXgcnjU1I8Y0JFh9nLNXdKA
NuQBy+385jJ5/3VH/Z+RTfvOUxoeBcLFeEr1GAo0rrvoSTtX+KenkkhHV9+cL6pIyfKZ1VBNoiOp
oWwpZ55uKGHiRJBoEl2m63SsIu3eyv2fM/HpZgXDUDLuRjjxxZkqKbjcXLg/iYvTSRdmxQgOE8Cx
7+xgpGoKg05+cx+cftCBYeJZKHA2M4dLIduq4yu4NLdabLPcFbNzNDtXT9YK0YF93yvOpSmN+pGI
S3uVXA/T2Br2jMuE2z0Ci4ppOVmbQEG0WCORlf0rfrLTuBfnBlU6NNrdhgn/FBAfniehQTF2YI7T
QWeHys86/32DyLjv6S+0JL/fKW9iv+kuSgwj9ivBXbkkxtkcilSS3a5ggFL1xrKHcfIlZXf1o1DR
TY1sCO00iJ/aI4sHQm/7pBLtVwSHkrldsH4rft3me2sT+73dleNVb/bDMw2VE/y7FwK/mODYcPCt
7IZo7OtP552h0XkaZ8VoOCG2aNBb27sdaQI7OinYs4pNzxSvLpx3rmzOAkkrdaNKOy1xWdoR1drd
YAIih+ACDLXqYqPwLTe2xjOMkzVF0lnvgskGAkzl/15FMczNYwzgGnYymA4X67SgPxG6ApeQGpTG
J/8dSaO0+d7PjYqnw4Jw7/wrqqTiGYhJNpGfRYDtOTWDcI8RiQTleoXcV3N1TWrJbyX1MUUe7tdg
vV0R5s6ngDx3Jq6BsoSHnv/M94MeE/im0gQYRkayq6T4a55jCNvehEMT6c5fwHqgNKbu7ZWqxDd8
brN65yFzAkUBh1Htd8XkRIWchSOkVLKy2izSUxTl6rkI/H0qp44m879J75o7M6VSXLVeVxWW97dr
UhWlcnMuaGbQoFX30KpoWEb2DEcYefDLyfIKVDLE/0gqUTnrfT674gryrpCUoAT8Mj0e/g9zyc7W
4RM+rYNsFr7R6+2cvd7RUVGNGTr/hy3Y//6kxUQXK/1I+O+5NMWRrfj0RuTaxh9qxNS/Q2fXEqfl
UCvQirSTXqjZCGjcndH6obsOj9c45cu/nC590ijIqU1SKMVBJLKgeaC7pHmNzSkky0fHs+SY6xoh
mI7pN5JH34RoD1Pqry79X/gPZrZCk5YJa1+7H1+B7iJoo2sRTA95Q7jEIxrC1yTig7cukSLP+O4h
5BruOda78qUwDq3WzXXJDDNnYwM7NjGpo3vzmuGIjkSZq60tC06MgcmXZESgS5gOCKsyNzJr6MgK
CRm9gceENZATidQk9z5w+4Z8EWlJO1TghMw2cU8R5zT6IHnvZWIDYBhwGVcZIduZLkZjntEzQ1vM
QgnxlXH6rPMW41Vdy1nra/l3EHjeh5GG7V3yBpIHgBNGuhDPntI60UzKHlWMC+3lFF0MgPEHUEVd
shH6wkg8Ebi6cqf1frtUZ/XJnWf/nwl/0e8GaKLsw8JOjHf0BnLrGFklBtWjw62b7U22PsmIi6Ln
cK5CEFYMTvVHe5xsrQOFZ8teYCMsNe0o1DE6PGD1DP5z4AjY2MfsxCs6pT/7bBKmFCj5AaG6ogDC
2/qBnmqCCVPfBnmTCtHY1CivmEs25gdgrajvIby/Afi0AQ47OhWrBW8nmOU6ZyzD6ujZ8z/rL9Uf
E62gJncbUgTlu+eZqQqc9xzPYHWeZAcIqkWGhHZQ74FQvV5soOh4kuh+d5CmzCxdjitG/rI39DiN
KAGIbLJU73VFhzBNiAekv2GuC9z5Uy3jEAiXfKsoXzWTaxxNXk4jllpcSE9Age4Bck+tiK1jEwuy
QRpcp+aCDUBK/ivX4VZSdopSJnfU8wabEPfOHGBgHaFqVa+6gb6OZ2p1zGkKtjHJi+2p9gAPhnWa
tcijcjlaA9CCCLSXDHtb/MAHRxNVtw/5DL8bDI/Afp1Qfy0rSjkxwocVWDIH0JbkYN5eBGNm4r4w
jn3Vnkjy9b21a3+O6Q+UdL4zr7ICKbgWF2v5x9F+/ZjFLERuhxdZR5TsqcHTumXl3lDD4t9e8gyc
P1NoYhqqVKU4FN+mZpN146+fybcmuTrpmILDmlD6776C6zAMHhnX3o6UBhdvbE6j4ri/jjPA8xSC
LBLfTR5czfoLX6QgPwEJ5Wn1kmTNe/PxoeoJpFQQ9k02FEqLv2GaksJ/yNpskBn8rd+6UShQvloZ
AsJjjoLjl4+/Dd3g+E9UXZC1kzvoAmPlTVnlbDjc9R41LcxGpnYVtSGJNMFwzzrcZwrwoElWpzWD
XoKGpeR+DyRjBVMrgTHIl9rlfOB7hxca1PjNSLcI+OSm1IpJlLm0K0FlSC1cG2m8ykUlwXtVU52D
HmqkcvCUfst/3K4lfi4xga5usmsehfjujY9AoKJWjEXaXDAcNnl4wOqJb97046sExjLfrxHLkRTc
FtvuIRzbs9KhmrV16kDk3YzS3TTXWRyP0amMdeecwXfFGM153EnBoGHBKupF/2cynwWq8Nx76XP6
jMG5/oTDJYTIsRANqapu5lZjsYJepHyBFPQ47+eT50pdc6vhmSq1LDDcEMBu8DJrMgJsMIeMknQC
QbhEoOe37+WzAwJLeoLWgC1XXQjVnxcAb68bl7tDB40NNmJ0qjJ8M6+RxoVYdaxwZNpNTqOnZcKG
sVguiohPkfirH0vFcGfmcrDg6WeczG8ULY+tQTYVgfnq1R63Raqr4ogeSidIYnrdHi1hz5tJXtox
tLaRLwynfKLLEEk2W7CWg+xMjdwzyFrrNDW2Dn2M+5+O2edsT6HravoRebIqU6T4DRWQtjpNoxPB
1HigN+AoCMjKZrKrPobo/kxq3aNblhMVi4jaOAjHzmcagFCOOYU/HlmZs3WT4PP59jp56oX8PlIy
Fji+tOmJYiJL8X7aq+NDf28ndlOOuBzQLR20SDiLh2Qi6AFW8ipUQv4KY8ziejPLAvuBPgx8LtK7
w9GXEZYPYSwvqHNCGeE1WX8b+sHIIC1hI7Lbxwj1tQAhbtvDczRy/hjW/agJMjz/i5r0VBDYQ3UN
GmKnX33/3Yuk6g7mm53sUZN2NnaYi21n3ZCPAjAEGH2bqxtgQigArdGZkzhytistebfQ8QDjGl2A
yU9/fq8X6/NhRXTmkP7pbIENECFW7SsGTVPXVPilFSeUHDpvH616IIpdA6pB9ArGt7Loum5Lq5qR
XEw6f7T+3Kiu5Oqdr54mEF5Aq4aYgtox+VLKuDqRkUI6UfYSeQZbDjC0KoOtZbrCxu3b9ufftnRz
irpZn3WBnBPigi9NlfemlZzPRH+A8dGd5aWTp+Qy7TgzgjHVKUNCckleenE2F2TaDB6fH6S++OcQ
zJUOBuA2CJC11rbg+BgpGmV2QlvbmKAlrGZinVBGxJ/vbWnaxkKG8IiNTkkThYgRIxwhABr7vxCe
uy0NHZ7w76Lv0fTrpdjXIuJRWxSVSiza70udBUQ9SGlXxOJWQahRqyKVHI+seV3PNrTULf1BimD9
t+iNGHFpdXhyAJXRO56Bxfk4HCogkTMbPW/eHcSkhD+dIoOLnUODUiCDcKo9AVW3zl+3OqoxTrlU
YixuRg8yBrjqfqUljO8orvzR4yTYsHlFqT3Dk3Ja0CzeQwM5/pjSh1GndWPxpC6lmgwGDvzmuEIV
19V/Nj2dhK9ls0zjU26jA/IbpE1rcxaBL+yc53e19ig7W6iid4GsHSV9bhfuZYe89ngwldjVJn1L
II5VdNvOSIPblzOk2JatMB99s5HKorJ4Qj8eOnIJKGf3uVwI5/SUCIJrDqZI9vqUuOJYHgGzE7Lk
bgXq+V4ZLNTr6arp9DhbexR9DRtGsnzGO+gP9K5cv7JRuDpRcafSbbn3zVhvw1LpE0A5XrwDZZaD
VrfzdFeHvUmJzd7PKYsFxywBW77ilcHMnxVDkLtmXe1Ntnvq6FB30HnN+8vU5x7ZRqB8ZFcLEXU9
8CXb1Tq9xu6YFzi5SXJTwIr+1z/xXoRN4SXZ2kYQqVk5phclXBJo7gkeON414gLJCza8HHfzLzBV
uAW2tC+X2+VZuQ0k4PnjLTrJld+dxUTFE7s0UmaR7wa12icCi5lhFtW7/C2Xpzol+IN0I4SMqqwz
mffzKu1CDaXRiV3N27Kbq6G8TvxkWuniQ47p3JXprnwvTFYNY/pP6KiOYo/HnCNSr5jsvK1MBhRo
E19gWobSTH0bKXAdR8dJVcgq0BCDwx57eSeGyAKzu7BK4podVBdPmuGYdAUv8SzEChdQhORQw9VF
Rpmpd8p0bp2UWYP67DQvlbl9jG8B+co3rexSRU9Hfa1IlCOF9qTy8+FEHbBfIwcWhxhdX/hI3mMs
kNh4nl1dPUgYGPX/14dmo6NvyUBGX8Wo2iV6/0EU3aecW+L/dFW9Q3h1OzTh6fB1e5ojdSU0q7bm
zdVk1BWLh0pDGbo7hHJbvlYmsVejNDdbYBJuS5l+uD4/uqQXWfMNqCUi+tZbEH/hX+y0WnnXcNtU
uXHMTZ85fxvmJFaWe9Q4Yr7ta36Nykh55ePq4lOqDKJn6TN1BZGFFJ5UWboLBV1p43EtFvunhA2u
O294+k4TJewz+f6v6/zYqhljFO8bZdKs1c/40SHVRFdYClpOEMy/rZFMBkgLjSpL8p53yk6KwtYi
Pc3AFhCm6kylrDips2heUbLELZo0BuSlRjmfKuC+hLeUg1NYUrvPTogbrc5yw8EB7qXw9cs136Cn
DjpMLEkGMhQmQD4p74TBByPJEsUZPUO/xSO+uoIaaCT1WGMelkmOzzxb8vXIJcEEPsbspm4cAwz6
PpOszSjITDCPjKGjjB5zEw5RgpIp0WOBu/H6pQpC5rEF8SVse2qLmKxOciMfmx4mDNbKGd1iQ1Xv
IPpXYPBedO6C0x5XCIQtBUB9XGUguooYC5ak26oVnBFmDtEmwc6F2mdm1I6BPNYlH3+KOVx/4LhH
OwYbvGTFLS7sXC7w6besKq559+XrAvIX2NXM9n+yU+U4u43sLIjFo8WdgGuSEv0MpUKcLNcxZBDM
A5yCgjZSly69eHj9FuTrrQXI5C6YlRkLnFMgHmOu0DOO9Qm1Y/rrr85b6Y7ePJW1aZvEzKNDLrPK
51pI3ChQB+mDvGUPcMk+PBHnYvTe+seaDRw5BHn3R79zCiGyNbdZI1l9A0rXdHXfMnb2hRTwZ7uN
Fcezfg8UBegNK7u/mg0STmlTpfLbgXRCIYZntuVaYBfuG5iwS5neiaIuz5UDszmRpAPSHnD1UR/H
QRLucRsOn4t2Em5BQ6FsIINpXdXIqm2XEn4vqmUuE3ps5HsWvCBvM7ZPXhvipDAIuOH7DdZ7IEuN
ZPpiJvLDtw3Hyzhgk4MScnIy5RHwkSBvolrHfp5i9jTWpkEbMsOxocs2UWiSP1xgQO5q4PicAxKs
wzvMG1TMT8iNStnQy1hob+GJiUflONJYlLqzGa4n/g+B2ysYrVmfrsHU6Dl67Hig1qhNOZomAFVg
IBJO1IHiI4K4+IoMPbEAAXqKH4oMYd7cYxRiX/f7FLPcSf3TwOpc/InXEt/qc17lbyzbJQF6yLs+
gEk1swAcYAHlQzuMQcsQwL77YOQOWekagWYH00uLau4UfENlSyHf/EIYLJLd+C8zLk1d8do3y3Ys
hLjv7GDqMTqZDFUqF22jtIRexp7DJHyT7Bm/lMvKOVIOquvj7CYARn2u6OaxuWy8RyM4AVDUCTqq
GoPXrTctEMUx1yVCo8j8CFLkNnPUpp7R0pd53RIf1Br+EydzwsNW0ahf/91pKYYT2AOyxpzkagOE
LWeB2ph7LXgMStumYUi6qxNcIemrhpX7gAIEWAeTmPxQO13uQitwLH4jN2NC8Zwf6EJt3sjJ7i1N
uoGbE/fgrJZRtIl/1t8Yba/Rc7IaGGVvxQG+dZd5nmevoIhfdRfIB2bJH+U4xhZF8sPFYQRG4TYp
qFK3QnfD2N9rBcaD2RuPYY5BtuQvk+VwiX5aVKXyafXyP4NLHJtqeOp7qCg1hwwhQdueKkoRRrYv
vS21HTZHnHN4R65y/IMQj5IcrC3LArNFYmjowN6Gfkh1Ou4GysBPF6/2Ojsy0sX5n5RCg+RqGJJW
xjZmTU/Z/+r+50TfjBFscLJ0UbCOSBrA1peb4riOAG1ReFeWsB4Vxs2l/KAjlOBFzRRd1Bv2xlsL
gLPAvLNoaT0IeKXcTppKob/YonVhA90M7JZTQQqqHGwJG5cMYuRpfLJUUz+26OtepQAkl5nS9YZe
Sb0cxfVwTc/goz0Trd1ylWUbFQRhTKXTtdfynEjMqrpmG7dApyHMv46fUffR7WOWJdCS9oD5MQ4x
9zW++4nLXkK29YEzIPTYCLPmdwqzmR/YRaS6Y1sLiPw3denknRydUX9fsIPP2CstNcaDBWOuAGYZ
jjWg8Xm4xjmRmRjh/na9evXjnBqATNginK412rubXQjn+C7OMN/MuQYNpan5uAdv6MYCELV//vbf
dZvRUZvkK3q7BeGUIdK298j4Qim/uWKxDseRY/LRoEKwMbROrn0Ab2QxUtKJKDngy8Lis1Whp2lI
AmDxk1nxrU7Lkqb1+54ZiG1nvmC0Eqk8pfE3A4pdCpSIA1EIWymC7G8pT/PW1Dj6fL4Z+usAOP5M
leRTcJsmGMn4JCnII2HATIuPwz/IXu2y6PiGmbstfY/y5m/QrWQSs2o+YyXRFqszwOEllrFpeSwp
SoXzbNcYwLWOEbAFi3pYtKt0aPeHY/2PwChUvFrt2jSFOYzECeJQQb7gLsSINc+U1Xng/66vD03d
jQ6vHl8YGMiQmAeOdlyXQsH0NCOuTogMFL7KIoVZ9m4+Mq1ups8hW0VvwKyRJ5yuu35cCK0phkA+
hhkOFvSBgxfOtsgeCdkZtgFOYwCrrEb6cHV6BgMauIv115Sjna+7+7mRes+TQ5qZi+262vyJQzQV
jKmfdKPgal41OF1pCp+AJ3BA/wBgt+lYnLs/L4LwOYt/IyPgEe2cOGJIZncBdswl85Srkf4K6wCB
5ofapMz4oywJDNgrd2RWEHwCRtOEmT5zuqv8c4BMbQtc5l55Z7RB6NTWIza7SGsXSTmPFsaihmlQ
9BVdvsVw8+JyC0Y7BEV+gn9Bj9WfEK2+JL9LEpkExWpX8rsejbbrt2mLpuC+sGTE41oBOCErLo9U
3yK3nzGYZjIIBvNuBy2KvSe3WtnYomRT/xB+L9tXvxOkpq06FziKgoV1e0hbRUsXHOO/265qrOs6
02x3crscLejyaTaJjWyFfXjC7XjKgicFvhW+3Zmf/MjCvRcf8p+Ficauh2h8adPrt2inH6GnwrDP
q7FWkW6t//HdeMJmkMFui3v9/SdY+uIPI9eB6tyoy3OFmZo67S3bjpEsp8Yd/w2TxaqsEPhdlgf5
LOn3G/M9a5yOJh1MeX7ec4uRD7aUcpFL38g9WCF/OvhJFt7NaUGLe0fo45B4bLyYFDcF3++4maGA
LQkN21ISvjcONjgEbZUrZ3kRwrCzyH17mCbFigM+k0TIYiJp+bExuLliCpONCBrkSfmWaKDoJw6V
opCtL8JfTI9YuacSlGXL2kC8eZlPyeGy+f/+UuFiETTl9eAhNTIyFzQLXgNZlun0eZ4X/kejfDiM
07P74PqSG4MWsKS5dfoV+sp9SrJ/846v13El4e1/JYFUoAvK+ovi+9Uf8TAldsQuvBypPwNu2Dcf
MAKfOpwQCl64PGNZvxf2Kc4njIwb6HdlWiQoPpHRgUc99QJWoxI+z51n814Y7OU6umGv8Dj0vUXX
MPX9JPFsybfgI6x5IHPcNWrhIjquCYpx1UgjkeFji88UnnLFcfM7QWhDBH+ISfXH3Us5PbO49XA3
OE3inx3FDZXXXrOv+65YtFcJunv+moCv2D4P0rd1JYawdJZlLpzsaOdnrJhbbaJPXuqjLS4oCpCr
ETAC3A+lBGu7bQhGHzz/S1AnY1B5Ycb0JeH9+GJofQIxJiWkCKvilyLBqVhAGbERTpYRkQm9q+a2
n7wLrL7quQjRRs/Fv0d7981Rcf5B3uVwBCwRXCTFy3W1ZltlrgIwPtpJN6CaoJh2ZbFncSRpePii
9NyZodjnWXj3tBEZoncoNAuu5zHQbqY5vkG525D2fBwcC00pQzpqcxIY376iT63vXucU6fr//fLz
Sis8YHxgEnwpZ0SJTX32BfWzj32XjxoDqJkkoiLdwrN1zEqYT9MbfK8Bgzfld7bPYDAm4/20pabG
o4/DfzlGnvHAhlY6jbHca8Dav3jeGC21+fVixFbSpzxbbk+vNEebpqXbVuvScNDtnDXc9WBSi6KY
jks4TvGtaodSYCUdVaXWGA8q6Ofgl5bzwIvdVXjYbl64x+/ifY4njg7ICUC9tjlarzskN7C++/xZ
7y00rBCVS+1Ds5/gRyXm4abt1ubabMWKHB6rfd7fqJISKE/igEtfQUd+vx4GkyXUzB5/3BU8aP1l
TXTaRww3wXWYwjgeILYmJp8XBYdR7lnbXTViK1ecVt9Ih3+n9NZFrxD3h15B0zNKm6t3T2ew9RsV
5NY+lEjW74KGME/7KdSLx4TMcWJTAN2ppJeTDV1j0vz9TTJG3SMEitCKUBf9XrFybmsyTQE+cF2X
jBFCtpQwBvW45hUEwt4NL3yqZ0I4FHinN92cnwU9YvQMixg9cHhsmykrPUIy5MWeu7A8qSVJi0Sq
eAtOx0UtzOwxxnS/ORdJYtUCg6/rMqcmFgiCsrdBBvbPz3gvldRwEbD47FeynRG+3fJ633UiUPqe
emg/ZlMH39j8QMbLvi54v3XTpKC1ciUWEfwqDgb5r/M3dbbyFb+0fsPnX2q7Inyu2KPuJBs9UsFa
HGPJoL5jhzzd+7BU/BpK+MKaVLCPVv1dhHHR3tKfMeYGdQqgjmAdq1dAXqPQ5I0VGwbOjnMCPwKd
0CcNk1YNg3e0ieB1cgTE4XhMOQzC/5VYnvsHPsPAEHZYrNiEYN5XuTEGk5jRe8n4uw5Byob4c+nK
zlMtfjRLAVlKVOLkKJoZw+KN+dBUmwtdIpLAPGW9S3hM+DzYO/Rt4Xiwc/Gd25jwK+k+cCADaVDx
EB5dqkncVu46Yrr8HhB0JAZBW/HFfHNgpCvbnp7S3hFx0G4CCxMYprJfY7AmhuthvyO+ABBTbT7W
NqvyP/kWqKHgn3+BqvJJCtNEVDgf2UxVMYOsxc1RSbrTXdz7ttXNryUXbxkNdJJiOMRavLduBBPo
gM/arDjHN8XHaHT+GGEWp8PkAqUwn9Db+SrXE7Pqp9ChsVodmf9ZVEqyovPtSCD/5BBq7xS9fExR
vUxyh8mNyVD+L+ew3ahXE+W5clQUAnipnH2e0psVUmN6Oq4/pmXDQU2ocGWBjFMX3H82bOWJwmLF
LqNduc8W7BQOzhyQRcs0cxPWb4GHDcl//T82Sw6aEoQiStOZCCUgEVut52PzbctATIV/g/YtchXD
To5nT41NImoXXsfGqrx/yp5kHDZ495TiXv7BUOSe1iAZSpgFodSFKxrKqEFLTQEf/z+h8TTsTuzS
rxssMrocxkZqIsyC/ydM+FeBe5oCkU+FzWzcZgzqFivhBcQXjAuRWHXOg+v/0ppguHQjY4W1g5pe
3Jxn9yzourpnxfHfoSspkYCmCOr4ZViuJ4qmu5oYS2wVx4RBiJDENhT5l6vaDC4119gICtjxs3ne
KeeiwDaPWNLQYJckMAXgaENEcBLKC8q7tRjXVTpN22jJaKLAXihiy9sHC/GF7uezJfdg8HHiULP9
umkZw5e4bHyohs6pUL0cjrhMlxZpMObJxNyV7kM3cf+VLYrN/UaEn7uXe+ZWA+d4f4ZabKOZLK3s
r8onypWcIWafJDRnzjRzXgZQiZsVfL542LADksc2eR3hV8JZs3P1NDa9vY/yjzeZgB78j1zcx0vU
ofGJWwQBUEqPwpyO675vnMrGn0B30NMuCxCvBFe7eL8sB4wFivzcDiMIEqMMyGUqT2MQmeVarKGI
B9hguvFUbRzj0Ahr4/IsgdVqt1vydk1lGk+x9WvvrJOWLnER67EO47lJzf6XtfbbUH/jsbN9dzgw
OeTu6dYet//EPjqqyHA2LBIii9zuCBGMO1Oih95jRu01a3K/pf3SnDbo4fEuLjnUugBAQTXhKvxo
xXu1P5mrCPqr7gNIWGjhnllMaTsPUEQ/hI5kdi8mQBWFMVl3J3kMKaQOahLUrMnS5A1d+YdnOUXw
Ek6Z0Zy//QcrycDWs9PkroA1d8Rt+JWcQyNyMz8uo6XJnH+dgyKs9wSLzfWFPCa8o+VkifoRc5B4
XpNUpZSbMv2CEx7b/07GBBOFXE9LF8no0ARy27VJvdfZ36S4pdlV4u/ub3Xjn7bfJ8pLobud+2t9
dwunWWIDpQm3RroHWgc4FJ0C309llQS6J1G46neSx1FSvmLkVhv3JlkArDAS2TGGeOFldUYRYBz3
oqNQIhINvS9UgkHk506g36V8tTR+usS1MkR7ZIg2TEqv61L2zCxz/8Ww9ZcU2AiKb9JlZ7Dtr4dD
gL0Q/b7K8iWirq96FoJFNkmqetEVjY8deHMKNazSacihuqWY2hDGejYoK95OpxNfdvPo6nqeyqMi
RRfk4KRpuRGCK6cmD7MqmhA8Xur7NJW9T0226w5cjfO9K6RX03HCbFs07W9zdfi5e7rioeZnDCAM
tw1iG7YrJbIczJTf1TW6S8BkO8HyC8muAC3ru93SbNJFH8rJWOi4PVWopQtZ7PQ+n/b7GI1TdAFN
oDWvzoEQSZ+T34Op3P/6DfFgdgJW/WSI+l4D0o/rBUdJT7UJHetlPrCF7XZAiv9oazXCDHaLD3t5
otj+KGHv05a27tp9/Ai4jeLx5R/+pJYfRYm62J0SfDBq5YQpI+huQUg5g8Qoj5UqWPCDinOuFRR2
L7TKyi8yadjgccM2b0320eeUhoQ2M54ak12gngL+kPibKDH88XaYxr1KDiTmcjWu2TKJB+/qhFYI
u6I9dGD/oIyC8CiXw9nsvkAruN0So+oWzmN3xsc8aLuADyAXupHWmjCMZoQX1tVfFnT+RrNbFTmE
JfhrZgYhnJezk0V1EvL/iUCSmC5jjTXy5auou5G3oPpnQQ13s9LuLQ9yklU/0IOrifY/R8Ms3ow4
y31h7kRqGsuaIpqiZWRTZwz8/Kz4ac1NccoRTkbtcHrL1178WjjII8J3N6d2lDR+aCq/lfIBoys4
yzf1I67fgvifFAORgWo+Ckih2SlmKewQdEC/knJIqqErjyf14Ka9xwFwv+t4/gDU91331jy+65U3
otrIW/K+Z8TYV7oE2iqVbFAcq7zlqbb0h4dMwThIuJu35QqqNgDZiy/n1PoBQ6GdAaGkJY1HRgPr
jP11LXQXlyN7Px5NbUBEk7KjAHQEIMU8xlCdXxqAxQI12Qefie+2XHhxi3FSGscWQJQWv3IdmoaT
B+GZnBQSnUel1lx8WjZDINwpx2fsHcIQKwdIeaQHNldXUZogLcaXMpZShKoHTvIlqgJztjFL9qQp
+ZdmuPeP2A7LpTWJRrIE4RLjtnCCER94+LKcXjdyZIscn3o3opIIyTEvBRqInEmf2eXdYxYQcszt
VjG4Jxo108/cOG4xrqRebQq5iB5KpdBq8dygmy4kNv1/VMSJJWL/lNVajwbSF0Ebt0OVquCcJKw6
+nhLpZ2WIUyzi1J14hzp0rKWUlcd9NhKcBo3HoulwHI9Cg+cY50rQ55MRhxKvtokJixg8/+cH5r0
63O4T3XCDVOFlehW8HvVunVcBaIWsLUEZH1AhupQDTCzd5uBIjN0hfLBybHX03g6jkNkYmpbUTgC
IZnGvpNlPDueOJVICvPn0eMot+irCpxEfGjyujY8Moqx+IfQH6uTjSJtUiwThsKeAIxj6LwGDobS
jqCElTgVlkfqttaz8w2lY3nO+f3bwzr8D9bC17bdp1rpqOekpN1T+3z/wnv+XD+Ipu1+312fmRyR
+n/sQ5qtwirVgSEFKKfkPoL1I/ZN9Yv83buLHzLaXBK1sCEwGj50yvUN+35kHYzNdpkSkus+Qo+O
ljsgcDKHA19WbnF8tXk80UTdzJCYNBgPbV2ow+y0a4bEBYGaGeaTPxSiU5Oz3PGHGnuAdGTUjpNW
L+dcdYziCjicdG9HN3o7zyOIbMzTyg2NsXNu2veq65Fut7Mo8LgD5NdjxyZ/G66fXcZRjapdpLaS
2p0BE5cXJtndBX9iytbicf9IOFlTesJ/9hUdJeuciKx3y4tIljUIIBaJTYwgxNshFRRw1IhpEZpG
yJt+dEG4CwbgtMvrC5lptQ6j5HQmKztrrzfCKNi5E/blWtHAiUL8T0U7IfdIyr6d9X8aJfXWvmNX
ncV5WjT1qksdaEZa729Eod5Wx274udcGguZlWbMEjeGl7ftuijsktKKTjLYjNFlke4pusZRhJL6r
xblSWoneDuX9rLq1FsINUAeirIBFqfxpfAp+fPQ6+Dtt56XDjGLDdpy4IFYMQuhUUJ6pJmryWcpi
NYLyW1wy+ikgUDvYfQQaxeTQzU7NOUxbUWDDk8/MNmfd/LVy+UFda6Y4qbPdu4/oTPI32/DmL6Kf
2E85yJpjcqme/NKZtFfyZGeyvS1WZgqhBihvzoOQa4yQDWMQ7ygvnFqCCICGRkRtgyXP2+A3wBTz
BIApmx8TKbhEGK7amreaADDE7XX6OIr8sjUMhsTwFNn1pSrEcNMV1CTPoSNFPtZkMXoY2R2zC/Qo
fvhthDgJsh9oXv0Go+TsCMmX0Q6ESJ6yr38+C5aXTlpgKGtIW60pAu6FTKlxkJviVURHdvV+noP9
TMShOc7jO1qgU5E73mjwxZLOhbU5o+YSzRyMFXpWwG1X9bObfHTF75zC770BPsMgHYCTriWh/qEC
oLeU82sOQh0ISw6bygyqDVtAI/w30NNzlnkFN1CB6XuIIUYbJ1XI/tCl2mg1v6qoppdFxZhH2f1d
s4QQihCUHhmGnWAmYnryifPqjgTt3jFwDZWnN7wFrb8PZB4ZIMKctTQWSIj8kmJ7bNF8q79bRuLX
+Wn51qrcKoNS6Na4cy97LC86vWZvN4jWpwzbLy/uGs/fgEMhsyoUe5cpmupQoMpdwQ7Va2+pjk8P
HHbKJ9aJGf91P1+3iXFxNG8ZRI32yjEaYI25EF2hOANTyA+u8hswQN4q99bSiM6mIpOS1MaYs+PJ
SxSEzy9+nEv55G5reabETguuj82UlhSxn7wpteDlqZKekrxyw3Xo/T1uQIAmAVdriPK8YnFzOv8I
IxkmCxyK2JMqXri14CXeeOQgquBv6BDeM3cISD7AKws8XbBOrbfLHt8MCHsihBG04f3I30+KmU32
3qIpjtsYbas2rQtnrs25zUE0rpPhjnvwW3BwBOEPXmc/jz/M7nE28gDXmXEEjGt7+gI9qHu2Kslo
BVf6jlqoVsBsXDAstnnb8nNnK+N/fPJb7wfS7CvDY88pq9tx9O7OcC3v5iY8WzjwPDUkGzsW9Ali
pOjZEWStESq7y5FELqLpcs60hMQdmV1JSrahef9p67XrIsMeef1H6Up4nyabhKlAM1gmcNdOdRjB
yF6avmy8Pj0OQj8bj7T3cb31MMw3UlCFJuk5fUgqV/NfzmeI31TGJ6qpUvVBzkyqqe1GuOUkB6Lx
p1130ZkcsqPTA3xel/tuujPo/Shv75TeHqWRwR1OQVpVjA7yF4mBN1dTxd/h7M1e9omGPStCdR94
9jmtp5f7j7jaf5zhOG7Y1r42mM1Hp4ZG468LKioBk06Gv309Xh0TGk+omy/WtlPPL3MTyZFdYHSA
JYmxMZaV7tDrX11IkcR1mWolC9x+z2CRp7ai2d0D0GkG/9hkjdZIyLjC3+QR2R80VDowrhDNn8Fo
UIb2n2ngUFX7xVMPEmaVbjSgDbYjuTOh9b5Qi9TC/pGYRn3qA9Pa5Rbf1R//ECU6KUu1oHNU/qYu
iRWUbiolF0wxaELhdFHbDjxzpk0NwIYrlbpcME/HX3tBY7jj6lDY6VCja6qoWqxWohoRG8st1IVv
rABG6nXd8nu7TjiQ0/7Zp6dHwkKU9B76YJ5HChNmpT3/G5IKGxgnqnztOz2YIYTHUYkSpwSwo1N0
268K0hTMZetsgRK17at6tOwDgeIaMSZdY29TEpKQtI6fg1emK9auxQIMM+JuOOpTO7v1bDkDXO/p
Ixn7lCw0Oq72YVQBM+0XAJ7kEImdbQ5Sk505+NRCArXy4DYdbLTe38JMkv9Rj++leSeM2BVPN2yH
4gMEtgk2/v6kKztctOazGGCmIZoLf7jP3cJJlrZaPapTvtZMCrtEi1gAnufqUbsdr5+9eGs4FZRO
HrvECk12apC3bKN/Y3X+ukusnrEchHQuEhO5O74V63I/oN28WqWLelxEfX64knp9AymYgoQ17mw7
MCYskVivK4qb2ATaww8NBwhQwLg45XpBZrnHebwxRXAMl6D4p79oklorWJXeAJ2NKZApvCcXXJAR
1D+1fmILAIAssKs1m8d/heMqg0jYOgxLiPv4tfuntxlEHE1YsWhl+79SVnpTfYKIK36cwFc7zpg4
Nxnuy7JJHYbdTXp9IJ8nNkOZUwgbfOXe9tH8vB4X02dOTDo+YvX7+6E+Gt+0lLeE8KIgr9Y3LN0x
QPlo20KKHQ4tWLVixavUJ1w0tE8afL1JOku0r0e5rbxxlGWd/uOTpMzkWsbZKLYGCA8OqkIpafWE
z0QTkeOL0JBC23KKIiHvnoIT3p1C6s/a/k4p8/k3SWue7BCubJ9D8j5uua5ftikBgJuzval4muH4
aOqg2sLV3Iub/lJX1p2fj15kudwz9+3WT2s9ywzry0Iern1FFwfNg4i8TCeLlDIXdCCP1FrC/Nux
Uxnz+QOUcP9q1Za3p5Lbl/OqiqQyDHq9gUmmCPoUF6hINbveHOXlCJB7ZZiqm6gpEVFAUMhyDbiA
sAPjNW9Kj8BoN5NKCxQ5mQz+mcrvbuB2kFl+o9AeAj6Ww3jkWmQUGwcGRK9s2hRfyp8RlntnGZHF
JL4Og6jodWke6H+go/sKHLNvYGOeUIbq3e9Z7ARF34dUMuMttWEDEisag8uPxepQgsuz0PDEvKlg
uiHTn+NMA1CY/AxD4D9gmfTriYid/ENTgIhUa3LKVCA6L1CxudPVJTfaInALTdaAE4a0VWnEimrN
t5G8Tal8hO/jYpzkS1RarIniUfn75688MCkEi5D4VV0GxKnF1KrOUG6IPRBXz7FeFjiXShw6maKR
Q3Vz0BpBu9JnpIeJ+hSlL7NqgHgqs6TFSa6Uu4RUfsZc3GtumW53ic7TpGob7d8elZYfZmWJfqca
6OI/jI1PQ+prJHgyofF2U41qKh007/qiYIj4I31shTRLtTOc1OhJNSRlMz7BbpCNE4C3y7voWuXo
kAammeCU083c4m/kNF4FjEO/0f4m2E/R75tceG5EoGFoR0cJGILIDd5FIz3FISyQHxAQM2zVbgKL
/HV9IqMMWF+0ApdFAtLioX5V6bWRjt3C6fVIx6ksiK9UGAvI0oK0MC3ec2bDNs1ZHHcN0OoqoAiL
esa7Zs2Z+5xUdMpjsWV7fYze5mQpyu5TDXjMsXsmxBS0wDHZRwxwM4rSh5Y34bIncsArx+K7jc4m
/XHZnoJ9fRyFCLcYOXk0MQX9fEEF5VRj5obcKSf6eKpj4Uly8GAvQN9N1q7ORgF+Ai/FSPZMZkS2
ZgwQD2dN+SJ/6Kfj9/agtBw3GVYpG1Bx2ABaQwmo7PJncaJmbT3Bb5DXjYUWfJaXP5DhTdVs30Qt
c7wvAyxtdDAD/2cEcsq8pnLJEKg1uh98R3Rdpb7P1yXWv15Dn6AE3kIfOQVQxqtA1NL96TJilH/H
L6dbuUZa/gCTvFrh66IWMhMWy/9dLSoNi69VUK59NBCrgeNUj2aC6oX646jMVHIKaS1sM2eqIpdN
UcT+R1zFZC1mvt9p+TX5sbOCyDcvH3/u+zcMsP/D4rwoON2L62NcfFb8d7cp9kMBYHEA4g4NYQ3/
FkbA5JKI0xLBe5pXi2GI7zFUMpK0dOrD/09ZwHAPstTePpWYeGv2wM85KHVX8+E44OGA0De0RC2C
1Zylxc4Oe9ufX4AIkfCIdC6D3kRwl/lePcZlGUQ3cGJI74VQGVYHBL+3ft8/d0+t2dPDz+sY9flh
Pab6cJtsi4fmng6KHAhceObbWo9ts0cmsHZNYNO/qedCmuEYOqsyAxI48CxDGdp69af7U7QaoSU0
psrQjFuQxiTBLytq1GIdJl9S6ynDWU2o/R37I9fuC1RCeIErXa14nrnpzelbxDuRnAymywmUCAN6
kG5lLRVkFx7QXjDZ4Bxo44l2j0U5Qyi2g8aFLX1HGzFMARXSQVtgoNsU9XIoNE+reTr9RWJNS61G
iqqv+qO28mCgdNkpy0w0P3AIRzYJPQyyNmS+Iho3xUx/UgUFBTdggy/vu0NqL3METz49Wa5W4xll
017VMAxFUDN3MoD56Llg/jen4ohlqDmO6D83wYoUfTPnHEhZMJOIl77ybFPS3OzcoS3NTbD23AD+
osryXVa3l1e9udeAasqBY5aPyYFsu3fOzgDmyQA0jPEvU+WsbnPKGEzdusZJlzyaNuih2wcRLrhg
eoScfI7NDGMs8pCP+czmf0cjvRmXmBcdbjyqMx8SfMMdvCo+5lIOfLjLRjNxipiirjKePzlhYh+9
j6Fh5x86F7AEDwAcJGrvFxRK1IpW/uL9zCcC0Fwkfmi2AJ5Nh+yqgQRk6587JrWKKooNjERjgi2K
f+rMMdaVfHqG8XOSzwBR8xUySAmzUdvTPLHMYjDDjhZWSzoMxFKvZsLT3xMW4g/22Ju22z2yjAb+
CIPl3u1CcsSiEXoIp8Yfg2HFngKfDlub4Lkg3tyD/twfINcSL2rU6yZ13TxN3aL4vbtHzngdL/38
RNhY3z6ZHk/GwWy1Tds55DHa9eb9oI8gpdX2fXPG0h/0ZUhf7k9TJLmviBP/XEZB1HfNz84JehRY
xI7PxNSmarfL41jhQzJnV9HBHZrWfFQlqxPQWtMNjky9Oq0lbtUGBX1o2aOH/hDULGZS6SNVzN5L
QW5dqr3Iv1kvu0jVwePPGJprEmE8kIks51CKVox8uaflbJ84QztXNXS24pQBC4zQGHUntDMv+1TT
7q12MRnQrf1cJAh7q6C+nCCRrYeUBfZnunWJLZ8kr/f8Wq8qYaosRjbzcsM4pZ/TVar4k5twZe+5
Nxu91G+ABuOVsMHThJf0PUnJAcm+mAC9diyhStRSk47wDt04jbYUKGO2GS0inlWLCr4dKb5RUBub
h0jx6JAR6cDBG5PNdyJjN+H9A/Ha1JqnHu+9f9mAtpdJTkaKF2bx+sinAkYE79EQurJ5QMntAiGv
czvgFFtD70R1PsTTI+K7se3FlSuw4XHGgUNhfeVvcJEOS3UEkTP9I8GXLu5rFhl1tM/KBvNbf0MG
5TBYQ54tPcOIc8mpFqgCwfKeoIo3SYWveHoqr4dVpp7NiGR85FmN7MCHPL4tD4tbsP9DxK0aDs46
IJgAZnSAcZj+U986/1R7QkMif7vT21M6UcVrY1PjMNLmbe61UyrUsKXd937K4RkgTza9r/q/qfMr
dZixWn+SOY0+g1aARVSVCPBMk6PguUWVx1wjxMvlOZdYGRBiGiNEl/l/bWc5hkPsvOHR8IH5xIWN
K2vpgpddhL3CIxKg1agESu7CsrBslzkqWrboYRtZ+dtUZIOTAL6bfg/vwZq4y7mde41LlUC+8DTg
eflY7qDvDr1o118hB34V0HOJM7QPhI3mwy+vCMmLHNbdB5UBtoStw/WN3OEwwR02eMQWZFnMk6x/
1aawBBAkAHfu4LzPNaSANgknl9b8jUXh1iZ1cmEvkFcYEgrk+a2H9iM/2Jjq5dSeuUCcm19VFMoC
rQiC8HQE6w02o/RLomhm1/xFSqRcDB/y0FnTTnID/qY9z4Yizt9jd2/zO4hh1GEkl9MCc1TxHdmH
pkz4oj1peGnUcUPouN1tbx5yulLgGiikD+F+wKqTKCiaHgWtWZ8Jp8dKVzZJ0o8Qaga5hM0BAdj/
cSQvhH5h6LDyhgzskjibSjGyte4G8mGlcl5pTlN46/B4ZDACY0o3loHm1oCczMalO4fAVRsrYDf1
q5B+FUNqkqeBuGoOUPPwR/cSTt1hH8mD60/GA0BksBIj1pDUtlQ/Zg5YASp4xLVGqqNEVqqR5P45
OKkmaTIjSUjFOEjKdAdV9pbqrZH+O+gcfo8+2L6LC/2MfnaEEJUq1rsFIRW87FAIkRI2oI3fQ1MS
4ADthY7Gb0ko9ImbXcHErry1UFJm0vvpZotkzFg2dARDnuOZLlvPVFxBrwFDyCZMeI4MC4FF6EVh
/v77Gn1Ix4+3DW0MNHHhX6+Rky0kOmPAFyzZC9LanTxGFGE9CFlpgKDXIQ9YZ7PnBNqgOdAGnbCo
QCtY6wgZKkbSIrTHLQ+DG8h/JJRWFWa9AmLwLXyeq6IZExkK9NQNSA7Y3y+pRKs0T7RmRvn+DQhS
LOwRmd48i8+43VN1HNlPOltbKOH5geTXuTL5ePNGAGnguWzEz0qo8vFHEDHtgQb+ADz4IYttPlPu
BMC06aum9XCPSuzbbzlr7UoDU0g9/p9rG6tJb7gCziAxGWo9pURjfXhANxZhhjYd+zrLh0fPSq5w
hYNxbgDRf4bL/ZKLS3V0kRZKMhGNDHXDYKYHf0k+a/AW+OJ2O7mgdQ6pWZZbMByurFXcg39O0qym
JFQse3fYLmU1CyF+Q7xEnpfnjS24llRB9ZvbL0DrwUrEE4ZrgRw5QABEXF/Zy5M9EBGmIVKdXuFe
SYvEp6Af0IU3JkTVRGX2uX4PLC7yNfHvvPqK/rzGuMtKxSW5lts4s26+ucvt5yU+GopSlzZsV43b
aJfBwV2TIGEq4wk/aPEugjX/F+6SQFw67k9D0p9pLaVolJdLWU8UP4UC70B/oGLExZGvf0cKL+U+
CG1zT7aQmWexlegJ8bqjSOmlYzRzr70s4pDu6v1xaert8ZTvtMXGzt8EU/7EPR8YwtIqPvm/Cz5h
YLmAZQXTe201t7Wd4PGAReXDgUoU+TsHmhjplmTqSs90hRskt7nGWAbaG7838Ar7TtzaCUHZcPuG
K2GWO0kWXkpaJmfhklylNwQT3hyEdi89qmfMdfTSd+1W1/Tg/bVuT47vL52IsjSGmMiAAG02uPdV
Q2nR+28X1Y1pRWvAxQ2pV2adCR0qRgmxZzPWLEZeL0mcJcQSz/Kol/0ycNUssyTY8XxZmfi1cNhX
u+3gdlV8HT6NqHQm79iCky0Thl3Znipd4arDSHzXrtjL6eRVnMysOyUcXt3KgizjuA3Gb1xNsmsg
h2VpwSB+nl3cDQDz04psuhR027b01NfqD0/HKG8TgbAnzg38tFdaFUiGTfHZb3eOP1bK0CXPrBdm
Q21lXTLSPFcomhcm4B183TZBuSeh3R6k6C2To9XxBPZY4acIk2El2cpXG7994V6DIjT4gxLUwCpP
ZrilLcfyzu1KH6wdj6n5WkSSXsmK6+wX3ex2GuGMI3bSrvUCMryOQodpKyAPljpyqTM5I8wezc4p
dipvsqDpfoA8Om1z1T8/6YmoAFUonC1iS1G0RxJUKB49i5Q3vYXkwaYkND7Pgg2CP2bBx/4ZPpKu
TC6jwuQLwGnpqjooHXk6nJGlasrwyRPDvFnzxPipaDgAtzRyWvySziTxu/9D3X8fP9NA2GoTZzXc
e/XYZiwk3cJN8toQwuBjdXmBKMk9qdlbTc6K0YxdAoyJVI1y2eH1OyAJd5ifmNFyN8Ky8x95J49J
kihSR/2l79y4g4X6/jSvV/8Ho3n0xKzok0tUQxxhtptX9pyg0a3uVwetgF0KEwoQLEaOom4XggDk
ihX3kN85L/pyU027OS4TZbFpUiKjQZS/nAiaPlU9cmp/g2ny8mjbbkPppmLzLXlXedxNQ82Va917
LiZF90VpS5bpx89Gyls6kTkT9IBb19MSOVcFEpNNJ1xYwGPeUyv3RvA5KbBniRresA5YXLwj2kp4
KJz+5WCjnHqptzFVOLyXA/JrIrpn2lw8BRs7h8vV5m3pYksDcu/5CBeCGl0xr0zPoF9CzWNtpTWZ
QZSMxcwH1luklG6SgmgZhb3T7ZqQp8MBJpf7H/7hFopFPif6sWy9YWg65nmsDmtIOwvR8kd4oFrx
TC4sRWfKkKG8aeaU9qRCouUdDIFjTyBw/KPERvxFvKYtvVGWPgbXSRoCKMwFUUbRejHzDqODjPCP
qU9dQfO8E04PgOkEtXu9hrvGAHVaaUAWJDYRtEdGek7UZINgpKwM2AIQxBBBeGSWqpOjkB4Kbvup
9+heccDeWfbOa6obstlE5xWbSL7r9qjlg3xYbLi61zhfchzXp1ecD15Wayb4UCwcn+HK4lw6gDJO
8BkMX2spSWoFPvqzXZ4YwRJ08YA4ETHm+OFnpm7eDzlKNE7fz7AhONoAIGCtrp9N1u4rLfcA6HFd
yI5thQ6yEqsuZTes9Pq/mtS98PQfQU7ApFGrMQ/PyAYz5AyuFnTDIo26LETXMzZrX6WzaLMfGiyo
OFw0GM/G0ZcZOWq47YeLySKle74CL5fr0upSr0PqCp+1WL48gzEJF9jm9ARbQ6Yv9M+BWqKSoTN3
KQvZsw+BBOn3o9xeIu01yvqOw1xglzQgldIHGvrzqhRgbkCbd/dayD7qhqgqRg0E/Ty8mCFAbp7/
d9+d4DyNJwswGvGCzN3HlT93Rfj0sWtlvo0e7QimHcjIw2fnVCamCXAD4fVq8vJiWzOM4ICLn4M0
H60oc8hfAiix2W8qXgYu9rIcBbeuv4fik6D7KaJuaKuVYx3W7Mu4sbhB6TnXM1vMAnGj5HP86Hym
p9zZMUpX55gGBSedtU3OoyxcsEamXsQuymXv+3E9m/FCcHNpwNDwmQzVNELOztcjNv2jCCueKlFY
8qBK+E+W7Mjs/kBRLylcGxJz5J7xJze2n3Cr34cEtVdJjvJUmbqYAbTwOqBR6abTaervKZttz6d/
OqNJsman/TXi/5e61GihY9qkiqWDlEc/jgXiQ21usvW2t/DQ60ag6GV/FdMnOfI7nkeUDqJHVSts
VkHEkUL2VhspbnKPW1JwGAGaVQJZQSX9cNNKMzdNziCxRv6cb7jXTGMx6miAEp73wwrMbWOTAiU+
k0jQzLcTc7sS+TKVRyaOeVHWlewltosu3OpdvclONCQlqqLMQmMZYAtFYZ4H07oQJ+AuFIGc3nJK
GzMcPV5W1EBSBT3UoQjTyTMvBl5Vq6X8J+Uqb8PjTJwKDqSUKicRf6tS5mIPbPVPW+EpSURr6PYd
iW6ZVXcU0Cv/HEVrtqie1vzqbKiCMW4OAeHMdjS8F04TPVzjb+j2T8Fg3ffMMJwAj3N1yEEuQDxg
XE9icRn8+fAc6l/9lPPmNDv8dgMC7bfoK9zzDNtUWvSUwxvNVRXEOI5KGReebjDXdVvp+/So+VA+
8dKiXmsIN2HHrhFeiEk2jAuFM5hV47NplxqwZcUYQ6x9mMEgtImbkgkLfa2Lof0wX3MnuJMCVPWo
dRK3HnrjbEetei0npBOk8S+Y6GHekwsNFghPtaPX4JoRA3I/f5o6nEJCZ4KKe4TrRzM3Xbk6XR9F
CNQ7Jm3jolmI6UNNX17icqhp4r6/YCxyFdTzL0YtIQ3cC6LK3t9PZCwsbLQE6miw/t7anHeeroRn
I0710y9ZOrvMX1ERVlvUtXjuTRgdrFah5hxOolPc9Q9HRqcp8tKuUuNsqhnV/0BNvdBI+SmtdI/M
fothLCcNk20ly4IS97H/lUvCswki5bDMVN25yFQ+C4bbsVFaG9sYUwfXehwN5/XlVSI7eXmqsesw
JHOt2wDvYOuWN09Wuxz4uW+kA5nXTnrlnLzMQrEQ4DW2aZH68ifav5bV/Aw17hwQbA0cmM+Wb6FL
Fw11kR+lDrw8gPXPY2n8YIzQFEAxkqscysr54imiQggvmGrv3c0p2PJZrNAyvJkS9+E12kbRf8Wu
rmOwBLVLoe3aa8x3ErIs+xLrf7ySdNxC57nXzZUlOzurikFTrFUfXIC+dv5lfNPYMu4LUKN4Uj1X
8g5kNls+NtQLZN2ykHF9ohb3Wp5piw+rC1Ltxegt4jK4D4fevHQiLPHkuT+O0J7stD6K/Z19hD54
InEXQ2uazDuSc5/DW8mSklN82Ems8DAzHPeNzDkffT6RqS0h84njN50VtmSrgu6bWwZexZOsl8wF
8cAY8A++UqC6aPjym6BfBQKBVDGSrry3VLAv6zf3yqf/Epcb32P1tOvdfFVAkd9PnUHHDygffUV5
MgVe7tsolx3fudP+ut6yziuoULvLB7zES+I8a7kOL7iqxb1ZYbLPJZ5Gqxg+FBZDLxywouZOwVo4
deC15GaZ0c8l2kziKddBCH4pCqUoQ/PD9DDY2IprRnQ+XbfQHRZ86Ujh7DYvm+Dbcqq6+LF8ewqF
slnHZt9w7BvALo8CYTFCztJNBqxns0sWbzSVRDOXK2Vnj2CgftI+7LMZWCr11dQ/KUM9Pd7zxcjg
c9wQVWQFSFu16f+bVkJwcvCIcNmSzVGsMYJ/XAqnMvfmJGkK9+nbLQwJO9NBwYcaMcUSyHAkjIFS
LYYEPVGZUtcM4G8wqXaC9JfVbjOCDjlFG0hgNtrPHGeOh/ZUYW1b5CT6N8N8PDETo8vSCTpYhgri
AB6xr25IppMhcdKKpyCfJmkBVNAPeFkx0vQ7HVBIwFlT3uDYqWNUQyIKNvxt3TEjHDHrEMnYhcpQ
zgVkRC5kPlejBhhv4fEfhCNr5hVI6mDVg6K/hanbbp4rUAA6mGyD4UV4gVzwGpUpeBiAzPc6rKja
LXGtk6FAWJvPaLXq2okaLNXwOEbtROmkDR2P5/WnGtahSRSuFMDoYwd3OFS8assOUiuOsBK+tF/2
7hn5wQaBuho9jRmsGqWi3pMuJPPWafp8GzxGq1LTXw6z3lgqfSsdWlUYzEyYqSF8+oBU/UrmkrZy
K80CnHTQVgb5WhIP8PVLeBcQqdpELoIbRsxUbQrRbyBv9fjM5WbewR4804X8c1xXchThK7pIvkQ/
wtGufMrjamj7CWqYSMYgedx6DlH91ZQjYdTHy7MSWs57KktNWQyhr17k0Et8gcO5WGn9VMaHBvK4
oSpmsMh3h8ktuOEhu4IPh74nJgY0FohpEaEODnTdeFiCFriOVQYWeHNLCnHQ47L1e9+9IfohBrZn
T5qv5IV2Eday5Of56O+hMMFeTbcBUOLBRUGb346CtRAKKUYokycLnBClDxX1u1Q9o/12Wyu0+Gnr
lhzV8MqopKYzFVkS5GfbaRf9ytOb/EMo9X4+ZBZcicQRwOIa84WlWjiOO5OH8hlTRdRs1NzPSl/w
sXeTB30K8xTJk7GYoIDUSM8aG3fY+ZyQvkJIUpMtIWvyYKMJ8TlP97lA6eDGKr0swiDtYBtKVUrR
neMzLTI2r5L/x4T487cxAdyJ8c7SbsmPho7a5oamsNlP9yN2b+NK7g45JM58PtQrpq81DQeZsGgN
35NCb/QpoLMVolYiYbFhyeQ9b/nhSMv8tORaV2kPp4WXF+iQCiRFXA0SgLJBWzXCD6aSEp/QOFpj
IoA3RhIUr2ojcIz8IQ4Xs3iFCUf0rgy4k3TvRUgknWKAsrkWfJkmgEbhD6DkGo87dfXMho17LR4t
UHEUuLY+xXaYPuDULFIf+eMEdFyWH87aTTx0Y5Vpjfy9WTsrIAQH0Z96dDqCsScFFwDBy1Wqb9zE
NPuAgeBIvaNUzAe5gryH9O7/OspLeFLA/f6PFCMtZ0jnYdeFHMVoktJU9eMKy0AxFJ1mLge/mgKD
eDdO2y370JIbEUdrSDh6uBpWewCJVNZYt6m4uubDBOvn3AX/qOmCW3/Ohs116dTRZDTwOH5q4bg/
ooQibYG2AZutOS6KWCPQUI+U+PoXqpDaFBCp7aOi/zfItA9q47nW/eQqmymY4UBseyWkr9qtKLQZ
ZduE5qtyyT5hr3/slWt+CYa8xnze+y/InCWkMMeBe2I7f+Y9+VCzmh8bUQXe2AXAZjMgUWpwjSAJ
Ul+EpWdk+VlHFHsOIEouHqhBc8R3m9YD2VE5/qxoSTjy5k5jmPUYOcQa48mMEtsdKLpNIl3fCo+X
ppuCfSvRoK9xTuCYKafEqofNlxHgB4vFdt5AnvPzl2dHVXpw/03NW0c/nhqaY87GN74ZK2g5+Es6
my1ICv05unwP3ybQYMqdAXaPHU17zzLAIbz8vZpYVRqQAKQ0nIT6QDH+NLPP+GY/QFRjaJiveivs
z8Nui7PO7A4ZbMR0QEMf+WvpLXhFetRET7me19q7ooyHsg6W8TRsKLcRtfsG2w/4AaS8Rg61A04n
t2gOSQlrBa4ieMD46ASsCbwU8uZM4qi4TYUXdp6KuBl1KPzsIpnrbNrcqHCVawyli7s7gIEbG9ck
ivrlENz3iylfdrE3zt4OLjFka9V2MWSYI9/mJPfIguqnv56Y1UjSk9qNADZKn4094WDZCFk7aafM
fVIzfCbkxkbirGmZYOlDfL3fPHUyVQjYtmNAuJJU08a/AfadD4hWXyhGdEvmc42sPywMt6tgl/jB
NocQHnDwH8jKl7Qj6HuyA97/IhhGEugjIMX/gE8dXFPR0XTq9hSFwpSQiDv8G7T0KgF21wtFrLhD
BXDJf1gd3lOsqlvV3q8k0nyLfNjO1rtXpVPYxLVTH1uilRrxFJACUAowhPlIMc/uUQaqBZU9vema
rc5BdvPSZ5qymmMxnw0ZBhcJgMWol6ga1x9em6OX8wdDUyyNCJnhQGehD3J4TP1CkkRlaXHjg2tx
+2v6OagHPPcyVZ9XFTIkYsGB0na2taL6O2BFDPBYxc8M4PBzE09Rtq7XWsHqU0NHEfi/Tk+FlZRQ
bKLxloDs/SWisD+5jBtYq6qaUtCGwaUdLdfkU/p9cm0bj79WX6p3K3VfjNE9+aQ+05YVWHqk6GMB
5lIqoX7B5kI57ucSBKomzzULkD5y2dk4fqcDKEmpWPFYewxePnrto12DswWK+Er5c8S58Vo3WD01
QvROIRIwSYPdZU/QXMHf94oOXYRs5IOoLPAjcAPrvjw3vVnK75Un1K8X1DBVdqtSzx7wEwpT25Vy
4zhdcqBpncXgNbg6Pjk96yFZET/mfGOXcSdlZqy/2hPnuZT3/KbvBYEj1yw2OSprR2wUP0qbQEj2
8A3dKm8J2jshssHIPpIAIfIuRiirftpPulNVqVfyiOnCfratvYnJ+LB8sMM8Bt8Ydyp2mUA6qeJJ
1+AZnuQT8x7MC4ZsTcXZp08BHWywalygwh+f9AElTJIrMgqgdmnYVR8fD50r4GyNtSgRD5JZjSCb
cQbPz2akzccamQUQvpH1oNn4fkDBwm3jDhxXIHlMnNN5OhMxidz4bw1Q3M4NMMpplrj0WE/jpVD1
mISWQY3KwX2lZw1G8n7dVAbhK02JZDYX+tV5BSdVwJf6rrM1bUNK5d3hPa9ABRQBlfKIvp/73dnR
+A3EaGDsI9aEiz0jLv5whSZsfF9XZc3PLuAc39ClS8QRNdceSNdg5qTL/2lPpQLy5GQ10audGBEN
35pHdfBzKTrMOb5ESDPui9LXe2rqPWaNGoU99wDS70tuWekfVas2yTyfVj3jH7k9SurzX56/wwG5
ybUMlpWV1r9uZIi1Kf8MOz6njWyCwSFh0TY3NEiHriG2rytzV0Rr6S0Zils6MJ/8NQIQv9Pkxq4J
Z2paIu49aGlJXL5oYeKtDloecCcRERXFqTAjJgQe0lIuLaYwbUB1C9cGf/r573r/lUwoTnZu2Zfy
7y4MxbTNarllj650gUemVxMqwQB8SU4sGG3Z9O2LL94LyCadJtU1KWU/DzowXyDlDw4ieTaF5t6M
aNjuqMM+N7XK2r0SCKv4Y4D3X0+KltMqTR1JfH+CxFdQ5LKS56CzZ2KipUu9FWAtfAACGUd8W5i2
sj6e9Txy1Qv5yWk87CKJ03JZZOLzH4VwbAq9hC15Ml6d7AmNhpu8/MtEAqxS5gKpfsIReVW1q5y+
F5sMlyZIAxp2SFh6aRryHyvThnTSA1pKLGFubGVB08ycKW5ArcVc/b1qHZfRu9Fj0Rzq/usZP2a5
A1wDwB6ezsY8dbSKjapFEScAjQ9fCy/6Yhji+esaPTlPU96EMEiGjCryBXq0+r75oyyQKekF4qwy
n97ytWwuznlhm3BI/r9sJ5Zue9UH0wyhAudFDaKihowMNp7/7mDyGbd9NsHYoAsgIQBX1pHYAOph
a/drL6INSwei0vRWSOt97v03IEVBzf9044Ba+8qkQ8PlLzY5plxwBrQ9SGNXBSxoS7PxDMbZLaXy
H8gKY04ic5cicssuaNXSy5EYjjVA7J+cWG7d5GVyLDgHlklro8jBwK6LU/7fYFNQ/7p21GT352Sv
3H23IkXIL0OtQVBMzbc12Q5syy2HWRtTWH/dw00oH2xnOTsEsz37da5XBppbPzRFNSxUbMPKLFhI
tkAGcjXHGFTPwms4dKvdQ2aWiXI3qg9rNEHQSYC6vv/OAeZNI4JYGsgvH/fXEK760mozKfF+pIBH
hrpVgl6+mytg1HPNKV1bzpV7j7AP4Dxe8zjeHMvvwotZKFKiFVP5KLOQVagWYaB30V36AUVTrg5U
xE0eLw4UohsuVPiRpz/rWErIj8obI05MdBHkC6VQVJYcxx40jiC9sr4PJXQG89VHkZvcakgPMzDh
z1dWO4iw+gR9uIb4VjjNPuiRQRH0A+HFvr7ds2ZzRa5E8nrjE48oywplw7UGgmDJfcYfP+FHONFI
VFuphvwvc8zevJ9OFkwovK+9yBbDLyBkuuxWur58VE9fqvcuKXPCKRKifSlJpBCkuw6at9qugaNp
lta+7GIS7t7G2rRKoTX0xCDOnrEkTgoCEaTwkHuYZU3SwHsCd615EbdZ4VV+gDPwe2MvAQuYJ7mC
PgZG5FoetZ7eaonZqha3dmzvrrv7DBP+RPUp/w+4g6Mjyp3fgjwkIsnTe9eyQB5Z1F7np4p2UnJ/
w+xJaDQ/CRSsFN+cPyDqQW1EH7rYuU+fqXXGShfYnGrBrA5TVkFKVRoDu3Cb/WEzWoZQ5kuc8WpK
YMWHAI3Y3ci5atvovdi64HAXJn86AQIcQ+lAzNz4gw42c6zFIwHPtZgD+lyT41E5yponQSNGne31
dCmQYGnjWG8e1js9dzBAAa8jN5S5f3FXxH0rysfFTYuzUx40a6k+b1hPaSXRmx4hX1hetzFRNdNH
jpW5pTMd8vg8+2Yr7N3VEKoYOq/WoN8sP5sD1krcfDNCt2en7A81pXCSWwnnBXkP2b4ze/jYj4m0
uJRySGfwcbZxKBLFzIcvybvv1zeNssyvJgmriZ+Ou6Ac7YLDat7B0+8nOsg7gfnj5+/fyNzcZsWN
hrvig7g1fovfhS0DTr4Flc4I11UYVYevQgWE7v/dk2rluWU6ltkneLrnFiC9nYtrQxmYY6s9gs4f
Q4tBe+iRuxwp4y4UpEy8ZC8jLX5fEVGYiymcHUvXjJzKx0MlRrxczFnSrOVbBAlpXalCfxKjYlJu
k1iu2yp7BBk3LgohmiCkTObEDDmg+3oV1CeN4voRGETr4ue9jBDqtwPbL6YzfYMR1loJC6C1kcXh
fheOmADXbnVHChcUz/yHbl6FSKXblsGM1ri4prctgAJJe7095J5c7n7ymO5dJCAwzysnM+DoxB03
6OUwOLhJz0J+ylFSBpY+aWNhjDhi0N5cqd+mG30TT0AwCJqRxlRIgo6/44iIxc8y6msEK0WGjEl3
BpMFPHpfSLJNB08twBTl5qlj255EvEtXVFrNVs8mEYZuf7ZCt4ysniJrmtDhffuEomvtcvKHm6Ip
uMu5/StjDkO6xqluFslHhhEjR/O8AZA+EbgdfyNr2DlAmPaSo6wwiuEP4VF3CGLWVmvgtEtrBp2q
YiFxnMedPIaWy0z3YyBOFrjRf5xgpay5rWKCT6nnKWnqDjdajIJ7RoMRU0DepdMbbzIKxHXWva1i
I0C5k3q3+4flR+Bj/nZdTnXrCoBSyFFNILwgmNSD4ZbTS/HFy8GweeAMq+sJT+mfiR/D/VKuvaZg
nchP64sYd4iKKVaWBadbnuct9DXP7TIQZZ+Ym76GvYE9G8h7deun6A5kM3TWFVxLzR5yz6PVv8vz
9BKIFlS3a2zVmTCm34c+G0+J7Z/bjOCMAHMm/a+EiKbEVwx5qmBQqsS/fGYczwi6w/fFREwpQ9g2
sJ2iZj9lbITa3C0QvfRRHo4qEWNpZGevaF+sYxixnwNGxeDYGcimorYEednB550UX5YrQwrTBBkp
Rd29LK0noDL5ZUxcFWn/MQewpKp/fBvwbPwUCR3Qnmvm70DrKj2RrwxWuH+YKMrR8PtfTG1T/HMB
JxvMdMkGzOwQ6c7CK7wvyTsB9sPY8RJcAHpn4Rs04A2oglRpiGmvs5GvkekWVs68XElT8xsSD/Dg
Ry4uv6FAtUNO2XAST5O4dqXiKnVWThZKBTRpqQYDk0jB69NQXRAAAKUrhxN2zTJiXr5VECIMm8L6
VAYGHl+9lqlg6CxNIMXRswArUyLeJcV3N5osUGwRYxKyb4nvbz6kbGTbKmVC50wMS5ALV8zEwVkI
zES9jeiKYSgelQBCCRuuWQn+g1TjeJsVS8VjzBj3LmmH6P9DYKgcP190kT94rR6bR698YjX4AHB4
vLAnGxCeftqteB+t9JuSjxbXAJ2+Gb+l9+Bm/D5NiGUtk2Q/eSsYFkcGP/vltixsATL2rfCGquSa
CJX6S2iK03xEULgelYV8kNdsdfVZIMsH9KLquwwZxjH4fTDIAZME4i6tZwGTkL+9v2l4q7zlUyBA
Qj1GjfiQFL+6lutrne4ml8BaswGkmWSKMXNSn7q1hq5jwaysZQECD1DjzvJxXVuYTOQcfgJx0KrH
HkBRzlGp6D1+i1fEWkdWpC7Iafwctmeh3xiRKAB9EUX0F7N6sHaW1W28iHGoDODYl+jdfUzssgx2
CDEaghyU3BKscn9IBRyGKjIMYDApQpPKgwaZJsEfsoLeqH0pHvCIGBt6HU0Yr2p4n9XXY9N8WaPH
3XdjpqR/FlK9z+aUPINJyC/NekivGY16vaHUPiIJjZXPA47G4vc7Ch5odNvsQNIoKN/t1dMILOjw
4ABEB5rUQ/Y3FojbWxL525mpJMcO/ecOirKtKhZESEOnQviexXQdv1runDSKwoOAPUtp/rfMJE2G
lcS1TmAg6snSMkuDxQUbD3iRl6lb7mC7lsagohuR0YfNypf0rK7OQ8gJOuKcPiNkjXrfqNcjD2Sq
mIfhRlCQCC0oNLUN16eaaEquzYrxTTtc7qz7mIOgQ6wrgqXIHIDUWy08uPeXpCznfU/oOkiwXcEn
sOrcGht+jKAd+IPgV4AJ391FTxtXB22RFyP4L9Qjp/CbNhAcLqNuL6fqaf+HB0QCsTnCzCfP8JuT
l/yWl4WiBI8IXSsw0g8JicdEXhSDZC+MnzwjO+/Vwk7v44Jbg/yp9Ylf7YKbFHy2r9jiN1w6z3t0
fYvXfkJ/kx7aUQYEjfci8imnt4vvWpBQZEA8tdQgPXRbL7YLpMNLFKhQmOzNIMr8RaThl0O4uwiK
xmDH5PKyhwEYQKOGDMxY2xI/wN8ChvCBir9oBZ346PoGErth+/u4GUXndgE7bvNqWOct/Q1VjBXx
BjCSB1CQ7n9cgVbCt6OM71enEVNC2APnq0DcTnCwQBXH/SrGAVqJB7H/WWSLJd1dd5vrwXLsTADt
ULe+w8Ey8MH/wPL5a7+qqTZ6R1BwYExkFx2VnwjwvhdqSsAnVkGShmdhqFlh74ykzmCq/c2pbLmw
wALI40w8nN8RPBD7V6LeaQcT14iyXHFjpkRihohiJWh99oDzQN4EftlIX8jnRG8x4PU0vQ6P/o/2
fv0M4q8Y7bUqrsrwg9LPW5+ZAkTg3jSIfQKpJlD92Wdh1tP3HxyzRNbI2VwCejVltFf4s/pNtGBO
Gn8TxCmFmpGs3yluUi0xlYoSTm95xGRe4YRz9EHY0kt13m3glD8WEr2PwIUpEpJb0z5ZD8VCF/xb
x8yeQrgHdPbJ+umAjHYth8KWIACQAPMzSUYdFGQnCR5i9lZQIYjWQMxl2u4criAtT3da2gi92hTp
fwwogkn2U9FXWZ///BdlfPSD105/ph5FYn/Xd3R5mfey28wZekUH2gCuUpfCbWWlMAXeDPmJP9mU
rqopWikrMgvrEQ9+FpyokQ4wZ6Oh95Cm/1SWqULxzfhKPZ0gnmyUnxls1qImzR2f18Q7hjNnUqj9
3CIIw66SRSZ+JQPzN91ZvplDVm8AoouePM80+6rii7UiQFAsrd6GO0sO6uPe08GzAOJB2NCXfdpw
h/9oB3CUE+jTPJhKERx13bIhtF0ha4Uy8VB1uySl4JYhYSc/QSsu/MlzVOgvkj/TKn7RHGZ871u0
wd84K97eSILvIIriYiSgkTG5wEyBMlIAmwekNDhF+/tfwNxIM9Xc3gHDdFkqC9Tuu6PRKHdFqJ5E
iLZw9/tS6iAvGWnp2Q/mlJAs6ftOQbjeOhul8169+Us8M+XN//2ArblDqhMN/B9gl8xzlehSuNwi
BdPKAbhOpl1ysU4uZnYDEfc7VRv91KTlwVak4CRDJtRSABlARU8iAY6BryP1TsNSauAirzYWg3B5
HVRWO9B89nmg5RiIICYCTLrW2+JKZhc2rE/W59stwNsZ3/TQThjOobV+hWXC0dKDLgFzI7XWqtDj
xlCKhttuB1LQLKP3roH7GUvsxdRLGJLYA7v9YbhbU6JccUBB+zdnIzUUpMlBsOC2a10jyUBJnJt+
NiwtfoTsjpHLio2xfoqMFaL3Pbyx1Y3VfSKLlgc5XWb9U2Uat1Cu26EQIiactle7dC/BiV8MhAHW
WXNJOWUWJnpAqYwBvG+1hVfMd10olI3wTwlERnno9bpPEs3L7wD8/Xp1OiEJCV2tZQbXe34DFA0n
bbloIrVBrH16/vdaCwYyvSqGW3Qr1eJiPdHzd7SooI+Pt9NPEcUoC8nkeRZChtxN4IEDIzD0Sw5G
pFzCFa9DCIUZhhGkMB4IWXztW6APcmMe5pg7l74Pk9jSU3iiMORaWk50NV+2pMeownU8o20qKaiU
FK1fujOsys8j4OL6+KZNPYS0whXSVvC8bu/M20x6KtftKzZM8UjQ5KP+C+0/ayEVMM5WuZPYlovU
rWMTqNt9MJxhManH8bRzHnzCGIt5l0e/TWhJ9mDmkxp97eMskiNrggKr8IRbI6OQQ/A3ALEPRuyf
XacB6zK11b6l7O/WH5MKRy1cjK3AQlz6dPmSocK1JLiR513hTwQ6nwv2CjcJYm35WTiNGPQzb4bI
2tjyDZcSmiPMVJn6eLq3OOUstjRCiHcVNEOZA1zf3KAuqc20tj+ivbnA6UoYRIERTik7BYdFXAfd
XDM0RSuiYmdFx7wmdcCrmyhu1fsG3ODqxyLLCknJ8WH/vLx48VcGLq/9JVQTQPxkhvNJ/qte5c9K
5LscHbFAP4Yf2LBXHqJey3Yfm1Bs2CEjXV2sK3l695GbaMvnO8G5poMT33ASw+ZrwxmTZNhWjYhk
kcz4q+hCu/YvtUP2vNCv87vrEtZ9rstLVygJOsnh6MfFsR84wp72EVBxOfJfjwjdYYY+71KwO8GD
+ST0kPw5VxY+lrQxXgYcJg7NKGoxJiw2Xjqlc41CsCOyiq3rx9i0cHoxZFai0YZ3g7vdHZ78qDnO
hz5dFB+1NT0YxY7YbUVP6LLpLMMrauTust+XKJRB6wChZZ6NcvbkfFzqftZ7SPp6VDFgeBQS7b/M
yusIFT/XLr3JYpOZQrh18bb/AIa91pfGV1UQNattBSORidX1PoXLbkcNGkvHHtWJIicqONscqmBW
+kTdy6LrAo+iPFi0UUOFuY3vEZLBeP0OMSDe+oam7Q6ZGLyulhhr7Ty8bTELpNTPCrN8bUzOkslU
r1Vkt+zANvRYcZY+vxvtMe4jgBNockBuMbrkOo5TRREDiaV8/AbcxIc3Q/kdH/VmBS9TtMR4ou2B
mWAN250qFPm8+xFcenB2buwELZpFDPWtOwXqWoKmwVFVbVSO4T5BABOhUWlx/7JdFUOKHrZwS1bb
lERSg3rncsIAUwl6/BFkBvaVe3fvT7yLyAQliXUVffRInwITJxfX7I6DeRbUE+Y2Ae8i/aWTjJrv
XjBQIWML04JkA37jRaG1R/kbYH8qqJ4Jona314211a2dKnc0IDJ6dLZvOl16yF65BLtAk5amHzgO
xYJLxwKXqUHpLTlw3JHSNYbBMrOediKEEkDgWGOtc8KLCHLxjKpp2H8dadfufLAXL1fVU7aQeph9
XWMBKf4yBUPjJ6qan/l0vNlrP7O/iXe1ZDJjsnaKotUTFzk8sdZVf+adyUxAnoUiyeGsLYFd9bcp
rnfScQ7vwrC66wbj/nArfLjtY5q0yOzZCYO4kMkLE/IV7eqxCyMZes7VEij/rA1DsCu4yjL/3O+S
7gvL/L7Z6bl4WnIUMgAgl6sQkSlLinA6AA01y02Jw7AdUuPLpjN+LP/3BQuKYTVfEkbxFFv2YQAe
LteIsQyZx0z/gT8azQ//5bOFcWMFDajvB+UORejEc1IVUxOmV2+a3OsDoKI0PdWuq3R3dL18tK0i
JOrEy7wr5kTRGhSI1sJDvssBnAjD5ZIEIAjuFXiGg5M51av29yRAeq+u0ZgLPw799xRneKvRgdu6
FgzrBXQyqCX9CyexpBrp+f/q9FfB1GxkvVWg7wn4nNv+H3Q0t96UeXSK4Xx7jzbp/SYeVPa3zWGE
Y1QDFTnuNNKxEwt3cEzP5TV5n7k9yz8fut6hg2M1ySRouIKRaDNpz4mjcF+w1+IcXVjwe4w/8qVx
NGdA2mTPKQPuG/869KaJsG1PZCFDZdkfSuRSk2toecyc0lWI3nwExU3o/k3wmkF4Z1dMLaLlwUqe
/xxNKXRzols/sVGKoTDs8HfnlzB57in4h3afXzlI8l5kexNX4/A6mCt6VcJGC/9H04vTONwbMXNV
L4cqEAiTwok3QdHhTYr1FikETzE2hkjYJBzR/cvkXCklom0EN0udrIhy7bJETTKxOyVP5xl3f8oH
61nE5abFPqBqeqI37I2AgdmEZkScIdc+nGTlF3wZ1E7kMVrRyVfo1kk2wDCuYEGcVjs3H7t+oFvQ
fs8NLiCL6F4WfGxzaYsz8d7IDF3YU0UU/RR4J1vQm5Wd875+T798e8DFNpIhuEZxu1NGG1dHEA45
HesPfgGu9RYXkhFcVz9HYg78sXnBOgwRc6Lp2yu8rNoOcxOl0E+LmKbtjQvtsjghYniuesA0o5J5
IXexogAKvQZOAB0Sn6Vj58udMPfzEg+EBCBExtdQPfa/gf4dSxAzdGL8UmSpSJmhSaVepHWgTM2X
/Dvkx+2s4HR4aWPjWBrAFdCJr1W3fvIM/1PHk5wRwMU8D5efPcE7A2k8inynvzcghNQECr/tP6qh
MFVAGxvcjd5tlXz79pGQhxCl171wU9nm4YZMINA28dsfclIDKak9T/Mv0aQRjBQX5f6rC5pmI8Y0
yDqyIwuJuCPXgmR7s9kL53Kuu0PDuk5fQeMBwZj+HRg5ledpRfYLxlP58SeFf8zMwEW7JSf+WWX6
jYM3BYJLHrdAJHY3Ne8e1ncDBYR0O+vMOy2Q2iEjMJeEkLnGCw3Yv3CPIHHI5J591MJ3GATxCEjv
y604K+4UiG/xnZ9gAPK9fBcWL5FkL72wxKpF9nG/UsZUbEN6eY4Z8PO+Bflwl/UIu2wnV8QRKMLM
KOC6ox74XDt6fXLQxU3EaaMxV+zXAAGiogMZTJeCjlcY79RZezd5fJl2SKTVnuWcLxp4BJq+hxuE
M805yZAIcpqLOv0VdnjjkHKcxEraZAAqC+yuey2mZcM8PV1uxlavgdPyeHzr+bEjIfHfrsxJ6cIt
ohf9EpBEWv1yupuJCq9zU/+VL0zNpDYg4BzptFMDsXeKdPa86FOz8yMtMXJoNBUH5onVRU0hk6oS
uM41B07sjwS253ouAscAdJHZ45DGP2YpxAQuLpYgivQiluBns1aFdOB0yBzWD6ZcUHBjWn+uJtN9
kw3Ntzxn7um/R9o8nJa93f6P2V/d113tHv2rdqxGfTU6wqkUKki0fSYvS9Eat5Jcx/0Q450jKvnv
wElyuMcY1l2HLUEnF+dQMNZwT9BJZfVyZZKGgFPS6jvfVMhVvRRcfelJo8M4oOR4Y+5rghEiHmDl
PmscjGpAzp8lZ9thTya6z/DiT/l4Xc8Q2U+arnQQsik8D+5nwfiy2367a0Pd6KbQn0IZPwsxY9fr
z1l+G3QdyWNfYp5wVE/+3uCY/60GS82cUCvSov66mKBw5SyeqxlsjfZz2kqqm3zVA6J2Ozhbwc3f
6YsMsADcVVhIMGwEUoL0ETsJBcIu0zBJ3aOpUTTjOoiDacRBqSd/N72fc/PspK/YzkW9XX7N457I
ABfkCaM+sy82WuHu8kAfMtaCwra90r4b6SwTFVnoWxgAF8G0A/orkgtP4eounmqL4464/su9myZg
GC29icT9X4mG7ZDSik0LTboVs1TQ8aZcWdpXVQwcJQQrw4JYQrpAx8Xmc0oqhOHHMEBPnKP9bJIX
xT8gyxGxVlc9whH8kapyJra0JDFotob86+1f35pHIRuYET6o/zwES+k8wOBypZscWi8Fpf/b5ViH
n5ZiBNolOE/8It7DoIojclc1sqqzfem9NYZ9R0qSTX50Znu+vGUgN90pRLPhbLT8Y4RT0I1qS2FO
8GTLDI0eky5RcfgB5J7DPR1+6VF1UYbMagtYyPHVH/QwLH/Ch73Fl3TYbfSUWXveMwwjGX30T+eq
8htKMvQb1PWkGvoVcrLmwlCtQvFwJkKZZq/YdneloxorpZ9NmBjBNjJ36ubokLHlOWdRWPsnU40H
tJFrqA3exEWYDUKOfbxPCZAQR+5NLoHWW3DfgdbUrPgi6HbsMqY1okClAkejVG9LRaM6j63b5OiR
PwZBopslC11DLnbGgcuRsJ3pZQ4sSiTI4LeSbCooTUT8Dvl31TIFPpsLEgnXzXfc3Xy7g771yy59
EystSp04R1S0pFAapGZpYPN5oQ2I+wGeilEdCHQNavRlsKxqhwLSpr1daRu0wzR2NZM1W+7UpFrd
m4zE2zypDMTc6Vonjn/T8rpfCbMPMOMlPKOkHxEouc3vuR1vRq84oCdYpRwCCwXsk3KROfr0oMOO
PpH8zqKBWft5zupLQgWgWx8w5+jbnDEhRu2Vw4IHw5QldPEHHru6N7c5Mpv6IHlXO6qkmXUXRqeo
U+iNJ8yp2GhxN5HrkMShcvIyae2Uu/dtrVbRLTksssAQFtpijUFzqFyyVuAKkHEhnR2RVRFx8m/m
BNwPUN5NCNG8pMTx/K9gh+SldFwxZuVQREn+6I5bCijdJmu4+rcOpKqXMN/ARTzYkdgOAiOk4SEK
LmgR+0UXRODs/ZTxcvCFq3wmH1/zYI+RuPbqpHAZrXelUe3hyHP7eCTU3xwGFLsslIfoSZ5WN7lJ
ZZYj5NfHYkXkc0edP+KQ2HWHaJFlx3lTkaT96Bhkz/SlmnMmowbocJXiHmaPdNADRsjJyEm9m85g
cxgKvUgZw3XHfaecqH58Gne084RnH5vNJ3kVPRFhBZnMdEx6tOH9w6ZNqCpO0LjAR9G5HI0Y39GH
17RqDF7meWmcn+xQ+lHpX3TisGZqH50Kq9E2TjtF1SGNSqEe4g4l/MXqrVlOyIoOBqCvqrVltAeO
aoJww0c0dk+kdFAGWyV85if7zQsA33MNvja2kZOSkYzDLtGGobU01VJcXhiXhOsxn18Wzokuze6t
Na4QDMcvaiBWMJMoEwskVouV/u24Om0DEaTv+Et0pZgA/RwVb07CRaKL6vSKqYCBwZQO4nIFsRwz
h946X38hFqjcROpW/NtojIOWtOO8YcNW3ar9AVDZ1PQdJvFe53XwHVY7NaepL9Ev+4lewjIcuJjp
CRSbxAWN8xbHVnJgsXwVdfuLQjmTTzXekVZelZngBvVdecX+PbR23Okm/nBFKV7dzhIKDf1MduHY
9ZcG0HuYH0eqJmyX8hqLeicTMXLXyGf9VpnVQvpZ1qPdPeAGx9fL1PZGhDL0P0sAcNEP+PzA6SYL
21bFm2VrMekLtepT3CGfPI9InNsl1TGytZi4f0j4DYyDK+stcHlQVQqAh0AOvXy2/NRyEdJKwGEz
2S+57Bxv4Izqqgm1O1sE79xbhX9Y949EM5XKC1HR0ohADEaYodjsm4QQdCqUEEuTz5cdhhxaZb7b
Gsg32fHnLwuFbfVDSyfyA8pcQdyPiyr/velCr+15zXOV6MnZSJcaXTLjPxhOO6PdNQhY05HwXJDH
lKn+215634YrkN5IOz5SmNA/19Q9oKVWy0Pdb/mKKKMjUTxvv4lkeVMJ9KkaJ07UPWbsyZPUpCoV
9ftubmFfWXBmn65TuuARNvj9bAsoOrpqhZubd5z/tdA8usPhFua76yfx93v7ZgVRH0/DcOsH4pI0
520yhLnAWQ1tZIlgf55zwG7ecD2G8M9Bqbrw2VcLWKCkUtpCbpJuQ/ut4lOrfFH/jnPb6ZO1cV/w
7Q+JGmJchRVD3riVwjaNdK/k/FKJXuS6hAY5TJt7wr/P/LgD7vo6hsTV26QLJzZjsHOnFBcG0BBV
tUihxsDXMDRuJpNRPLFpVw9C2HWDiEIIrV1U92N75RmDun1PpZkOzuAiHN+Ck2lpbgPNpJsMk8bA
RaCqurXI8sX9yn5SrBXTju1Ao5NSQGlKsCNNbz2PeLH/qOns7A6CPcYFT21E5B6EKDPmU2yJ8WTg
qa8/Q2TdFpfA5kBHVXouwuhmiutynD7c1JvQpD8jBfUHa9O/DxgGPxHffuQa+2oZCZ79MadXT5o5
2ucSdnLJrtJghkGlrPGciKC6hfwKuzMTCl9m/XeZEtBGs2gLZuOpOY3fvehI1ZReWNpghxC+oggm
EGAM7Fx3cAKKlbB0AiQzXawPSTey/bpTO/UPhvQ4u+9556DnqpBQdBmIxv4fKkYacwKbgXrVy2OO
pljRljWMyWsnTghNc6eY2HaSApbMA6VHy279RPXrSZ3mllKqRkZd2aiZhb3FM8oFWxTtXfF1lRnd
9TgyYj4OxkCNsTrlFvhwCQ75AgMqcNRXhJj7Izfu+mP+xPvrOQ0oEv7QVTDU58eVvN5/32uMMVYv
YmlVS8yOVB1CPY1N3541UeQAUj5t0Pq3B2CEAW1T5+gEflY+sY7jGPooobpS6GWO4Bp7DUUFLlIC
+NiohZfs8XH42HIwhck3UEvUXjDPVJLsfGmy0KT6i96elv9syW9Km65vz53hz4B+Kh6shLGkiYzj
uhtZtXVvksOoXqpwPtGWzMLtLrEiDgLJxu5Cx81mGb+lAIApwWprz4SX592158iToMmxbFo10cl9
YkKhBYwe4iwSbggPbs9iQXgn2Ioa67AIg36eG1SkatgwKYlSNWIzwUk4qMyVAx5CLUNi3Hf5MDkA
edNaaVYqbR8i3uEdBU0fhL4FKdrj5EjFxfvxMi/XhXGX5h3mt7CxCL4uYhydZP7v829Q+bXkXiuA
n3iWVZq7l2MQkMDHKednsA7vs7Wd0/k0bXy3u5ZPPG8jpcm1lMySFUCslpl3S7mAxiUchix1aIw3
g0CnHnwXxPyHaLQPgl1suH5EqdhsvxQGpCUOxY1hKckV9sOnJ310Vnj+njHUzXqkxoVRsr7etBCR
5Y2dr3HCe/hJX0cww0Dk+RKy2jbChdAOs1u+3arn6LvHHYX6OkmHLYZpUnmGxttSEq39VtChzfLK
lxo/gwLcHpAOaSz/PSMeTwGPf6uquFhWoJY+/Pnyq7EsuKsOPMB80akq8jsyb0t31OvdYiAtP6RW
1WdU6O9J9dmFwT/cyFXIdtzW8/mKuwRc2H9C8A1hDDVs/0uIbgvcv0O0E3AjKaNAV4iOutJ0I888
3KIq+gbgSmPlG9y0B16k/nrWsGUNXkU0Q/XwjrN2ht/swYkZv3iqTqLf2XrpbAsA6bjscd9F7up5
gYjieDlhJ9bGUnMqJnBwyKclTYd3ZUM0yB7xG3cPcRfSdtvcjU70TQHHDLH8bf76rfnhRUOUvC+G
IUu5Uo9prVIhqBiceKam2FAfH+FDv+YaRDS+P9XwrKfXiBIitgIsjbtHyl5TGvrQhu3MbZ30sHi1
+4ehgj1Qj/ftJc4zoLsvGUV12tFWe+oODeqZi3+Hrc61HPIPLCV1YERfUDL17K710HOPG3G7xeWL
efW+c1PbdXD6tCSVXb9HAkvnSxdUNsoYYQpUijNvAyCq7qf/Nm6Cn0uLQyAewC/xUthEzbCmyNUF
yW7yiG8ogx/0l3jQRcPeqlgnKUrMdgM95y8SdoU6Vn7Q6ysRmdY+pAxPQVVOn5MRkyMqmBQUhsLT
PE1PNxrB9jbCMi3aQQxvm3eroY1FMeMwpsFfCliN7VmTRyFz+ykp/6G6jJEjLboM+csuPsu5dSm/
OsIuSQIm8pVEVMpOKxZPmIkEsNSP0+YBHdggO4Z1+Q8q63d6fgDBL+PR7phoJ8h+VbFVz0vZX79p
6XMffHNF6AAxap7gnl8o2SbTRSKARa5bgxb5BzYDVBRJByDZuMup+mxL323Ww+2pt2YUvUYqWxZg
szCf5tnaG5Z/+Z8+GnLH+UnqmH+nje+xOizxLx9bVdDvORzaelV4Yb7iK2bVJg0pYH9ljq8+zVvl
4poq2aTs7xJC9B2n2syDF5RDd3Crr2RuX2g9A2GGn5RxuTyzChCV7dBjJSQKTL48P1hV2d5bl/Nw
HhWyBBD+X3idcaG1L5rBL9UqqZ9e027tyd+nofrUT8/UNt4vmOkeeBdgxync/NjmCYS+YuDK3yK+
BzRRUvHQgd+q25tkCvh/RG5UcehQHXNbKwxFWPzcrmg318bgNoV+3PDh3oAO56NAB1G8bfeN3xVI
Nb3udsSw+k0w1Pt76mYc2pB9SusoI9uIbL9QPcOaOQ4blgLbIT6THEqHSmRy66HEJTCxDN+e6Sq4
9PZM03kwNY1i94ciCsikH0vvWf603eZPKgMevHxMWn4cGwV0oeXOkXImoy7to/yuaPgczZ6D2mfH
7c1USn6SchwLyyN73cpFcbp5Y4pFGxPM2xVaW4blLC1nTXPASdPqWEcHrFjnNsx8ikOkgUGAM5Vg
knKqIwQwK0G4nGMt05HJhbU3iRADYPl/9wbTwxxz0prcudvvicrYBcT7+1EmiQ4IMoLmi+2ObfXc
6zY3dMt203nAGr7AjYO6u79j3hHityNJ5diIPut5zSTzTegoiCMEj8GDxEsq1WA61Q2IAHP+gZEj
dPzk04T2dDb13BOLoKq6wfw6QbC7Rn13snbBfP1KQAafJcDhM8XvAQAlEhXfDwHybolov5p/Pk7c
ykAYztFAsT6kwIMgu+lx/OR39yTgip+NVFVDtR+qM0tYfNyx5y0qxWfBufgmaAhpA5EdGHp+CUu8
2dP17mgqKDEG0x15ijO8T9hhFBbPDWgWrscmri90du35uwsAltZ2xR1VtMKCC+QEC/5Q0rurrtaM
Jr+M9h4mycsHlKL1zSazvHEADsMdLMctonm9Iodimw0lYkf0nR2cpq+/emHfUfdQ/sBgj7Ac/VtH
3q3/+fSSu6usdnShRgiHsaTqTxjl6smilS2AWzZg2KapRbaYsPA8g642t5Vknd5IGzIE/EWdFDco
0NdNUKQUZ+QjYn9fQpoN7NYxRK7AABx8wKcbYPmhyvpD8qXOF1oD+f9/acFwKbvV41yuje4ax6WI
VCBemmbA8Ovs5U0HCYfF0E5S4NrGsX0+rQQbiQZbdIc2ul7gJVlcJDBwV1ktNW4Pk8lsKi9AR9f0
hI/r+LtMBSqL6pNtlrNBdV+ZS4IHv7aStwB5YUcY3cOk5k7HXTREEF/b6vgGSEx1yFNmzFEzg1+1
0+x/Xxv02Cve/itSq09hXNqTfXsP1hXT21ziBT0r/FR8jdA7WKuNLO+VaCwBJLUEqA86ukvLKzng
Ta3P9KuNJ/cMhorW82a1hhy4+tsh4uIMtq6oEj0flbJ+9ySVmxx1xZ6eNkozLC6+zxuBJBBVWFD3
vMdzKNpej568+6SOkMgyKMvgpzOKbZsG52/AKBvhdVDjfbL4QUfCv976uNx5Ht/VmXjhav2tYxf3
76jmylPZ2QFsu2k4nc9z5k7oWDnp35PXMHBIkcXkc/HmrSY5A/LsQwPeg1deLRqpoiQw2sCC+IDp
SuhC5zZPvx275MUC6Ajc+dXhHLtFUS3INFkueD7BNObd1xH220l6CYIzuL4rrQ+dtnpsiBC/TD6y
p4GGo8vpCZ7b0scHrqianMg2Xr7NLO8+SWcF8onXpypjZXHsp47vqdGFQucpMDDszpIXtvfYaf8R
VQuujHT4Ioii+CunXtcwT0AYNQyVvqHpSq2SbUdDuRfP+IQw3dvGPNEsDHycfe+msYD+UiUjj3D3
xymuXLE/RNHj2IyNgGY8NygfSXm1lCdQ0ulYheqQQzRSap/2kC39G0IvUHWAT7dFF9oKOfe5M0hQ
BKW7oVuFTBSxXWb3luT/+6j2Tv7HWjDGhgGs2pmuXobQQIg+NqKmhk6LDPtVopCrjYshHyNIIJB9
gkdMJc7Tw4j+3KO8GDxZpjZQjPMT4FeLAlyAF+m3PGP+aUTwEWRXFMsGG+9aFyiBaSxGGDQEx/ud
IehzQB6pUO8Hh5zNr2BGIX7QijTFrMBZVxe0qKGJHF8qAa4QmnnA8KM2E/df6xN/zw/YlKF7KIM6
vz5+4LfpteiTdXbqZpmufVwzvqoKBnBXP2gbqqHsFkI/x6/pgZD1ivag9CNRAMczp8k0PN1oil3m
X49uyCfYtVRTmXujAMUzKkmZ8jnTbp+ns9zEvH+v/me1KQNpI8Q8iA62dGKM3R/7gku6iIXLg0FF
Blo79yryL6Ux64x9yVgR9axu2qPPPQCvRK0FGXIzEm9XHDAksKAsPdUEZBipEc+UwWRuQMg+VDAt
BC7r0glgMSX7i0Ci0W3iU76Mk/JS4NGaUO2mBI1I92MYH6YPwk0IiXN98Mzp6sGKIQ8hpRGQKL0j
SzAnR0qp9FVnroFg686wLRdT1XyYO9d5Q6rrZ58nvZiRz+b7juC5xLulLIHZWShzC+h1o7RfQ+yQ
Ajr4hupHOMtEUmRNgwAbHnM2BBXuzIbGPrGwdbFKBi0US3JQTKT5JyTFZwbkt/oF4n7m+FpYMb7l
MSSuCqU3OC35/gLASW/9IOla/OCZnNuInXf86ulUJddo8ThKZMMflHWCOkA8dqlAeirHRd6O51qc
kKLNCmpbCdL4A2lUUsNHFOQQ4ctlKZ832AjymB6VSjJ07xCY5++Z7gm5g10xlJAIdvjh1d0LX886
Z2V6unS9PqPICEiF32gNdI3F38iybmQI/t4xMdf9O/0hZ/yRE9AqWggSvJ78jsVI9dFoBNLzODRt
AU1aY9aWRfycckB5JQnM6U8JKerz1AJ51r3TzdaVU4aF1oL7Cr+bAQwwWBDS5ohSj2HGKZfLDCJl
EaOBV6HFp068S1yViy0WrM0rPnpBC+NXgWj0/miqlZz4h7pPORK99LjCYLKrzbkxwZ9ct4ceAI1y
mgQOfBOK6KjvqFLllLCMV2uu74H7zgWn6JqO4RAWNo9FSL1tczjK2AYHfyP9ZDu0/HSzRODQcYi0
7eFL38G7nGEPlpLlR7fLam8NDAmDPUifBKSMKgsOpfp7b+rzr020qKTShPhYtGhSTWBhRZhgZrG/
x3TWon3FNlRXTZu2aRDsUL/jN1VnuP+OdmxNeOQNqOhqJB+I17/9vDjOa6Qw11n1T8NwaaiM+e5P
1yekDq053eZ74TM1UK6O7Meu2R9dZwk3RV267NqIUQKz7kMYbFrcPgkxKC/q2sZoo9WAkMusRYnR
MSZhPpOMvNbhIvrO8XP4Oa1a966Vaa7H9m4vJa2Dihmbriql4zeMlr8ZOCxBz4TuOLtsF/37wd6n
9AXNc6OlB3ni3kTl4bzPfXOf6mp3kmDziqYU+x4xzjNiuqsPuwwQD7SqqfgutDZEZG7vGZup/hf4
GLid762WQd0zeLHfIwqyBdHjhinw/p4EliyRtuu5VswNj/CEkngI/p6d+GIGX8gkeG6IYqaDtE40
2JfIlptkfpOoPnhtbv9COQe79VeljKepX8bcW1xw2xbJ9TBJMuo8vNPuzl2SH4PhzlAtYWr/CbuC
uHSOuEkM86lgiZkQeMngCh6I8BX1/nQJYsYvKMlD869HPjasjOoprSDU75WdBMUtubz5q1IJH5JA
VA6HKr0LsOjF9rSqYajHSPEx3tbvkQ8uo3Ry7/8tQSDMX9qdzQBrQUfwuFqc6y+bQtaSctwajRNN
xATdHfaGZrL0IeEV2LdPJ+afElQxayuBacDeveN0zn+96Q1uSuvZJrHvOBzSikCX7Ed4JPC+NavV
PIbgxrteI+zXhPBErBEz47i9IwWfZvxnBHrd8ix/xfodtASGeo5EB302qAcsOuFziQwUir6wO85y
2H7VZ+GMLBu99X798FCLb3RCozDKV73ssbnqCcxSyGcLlRXI4IraqELoEIi+nc3UcCfKgRyoXqx0
LBHEfnS2bPWJPYLdJNfzFh7h4nttr8xyxs+rHbyf4bLbCJvJkK92rZvL7C5y5QoUFkIua2w+uUhM
rm8QDqGh5ADdaYoPBLS/NZrlC0MGOb/tQrmHt8ndceHxw1AVCU2Rsh0yhrXpdSKCuCwm7leMW5PO
uDOcDlHmv2/Ts6HPDuQgkCsCti4sjUWjSIrDlow/Id2ZYaCeQDiikzYf9f/I7OFRvlYKo4aBUeKq
0+9yf4hN9Y/yBqWagyG07KKWDvCE9qkw1TQenaFx+QblusL6tI6HitkpBfXvzL234SJd4nMF9ids
yOaWCJ+yjKmLuaHX8JSx7wnOnZis6ghRDtu2tENUWXnlZ3VxunfnK2FyaYk3ChAMkrX3b2cc5uRB
FK1HHLzd3rjtjiZrdn8W+hnBHmqxZVkgYL3CoSS94j2R6Ba27sOfRFnmhoMCplOInn79BlldDeUE
naTKvwdak30z/pkpeWR0eUoUKFT0ZdG6WUbgx9g6yYCiI3k//r7Wx3751+JUQm6HbkZJwjccLjpg
LWt4nNGu3jMnRO5MK2D44x6+Jx43wVcMh1kBZk9LDAxFFIBW7gUOd/++2lDjSNwbfThMngfk7CoS
Ui5AHWPV/GO652vYqN5perAo1pOuPaz8cgD9QgcfGK5GuGogvID7Lnu2IWJBQkIsBHDAwVjL0X0g
bz8H55XQpOA9llIk+nncY01MDtrCk+G4bDOrRxaj0eNEGVBvPN4WDYoJRa6umP/vkcaK3fcZ0Ii5
v75u2edSExqZwgofMiH3zutJNAfrXqLWSv58Z3xNKtChyfx5MtwLIsbqMb2E/TAPob5+NwryYKgI
yJH1cyA5ds/vYlK9IN7g8MuPwsoPNmrXWWSA2kBce5PcKKwA76z4FpvcsRFW8MYPRUxD6n94tXWV
vJSlcf1jzN+NoTg+HquRwex90NXEuxVg4UpdbSMY7aTsUpkGNgK8fGcN6FzkF5CbkMqaTho84cxf
0pkR0e53LD4+U8ypgeniLzgAxKLgSpKLucQe76ElRoxmVHZaGP1yzMBABH3mrLYJ5lHFhCFd+chF
8qHgSoCOTcRuNCzFvJUNWXGg8CP8MRwRTLWGqu3WoVBc77inIjJS6ZlyWPxDWz4vMIC8NcPqwPGS
WqW0Ji8/87/mlFVeI/IcDU6N57fr1fSPH00a1Q/hbv95TMgJpGpCxcXgGzFTJ8cU+TFBYys2KUSa
5QBiv7FQTq/yZ2oqUrlojPnMpwlNVnf0OR9gifUtPxMma0CWnYAjrWqx1PYxqB3B+EtWJXcFDdDI
v6Lx1TDzLWDeZvRhE8cYU5tP3x1ZszAYr5wf+H0gjT55jxJpXZJ7Q26yBo7hol8ZjZoB2VMK33Ig
sC2y55Cc2UVqx+zSibq6NNUxiBziYE16pbelHGPIV35PwO5XvS6Udd/tw4QWKhWVIv+QCQFnMubX
E/lvxBqUan3/HEy8lywBAhTWZWq789Z5UFpQUg2KpiTBgLDPLUfErefe/CFUt9bZ+/u9mup2HDP5
pl1UL5C8IuDWcCicA43aLTo5stufiWRgW0zkf8Ee4thp9uk1jjRghW+n3Ayqo3m+ME7WoJGvH4ld
AhUXTe8X/Ihz7p/ti3Ypn6JMFl/FspLPfHh5Ud51toUanOEcu6wAHrdf9ypFfCZQp3+bZjIcTUKt
btr4luzCd246gBLkPLQn1yhGdKyVhGxjtw6Qh+OKq8UN+5jMFUubthxDqsJ1L9PpVo/MytCp1xqq
x2hEooBEol7NpNvk0UJq5Na1Zcb5hDGnSmcoTybG8KYPY84f2jTHtDu2fGOfarxHm6RKmtogajRs
24ghcecBRNs9Gu8aHiv6BTG6vVSFU2Ur3p2Fs7aFMuEm+HX1rKdKqK3JWwPo255wL/u2aOjCyDTS
Ht3KE4UiJWFJZKndGO8HTD5wRCrYOV/1rcv5qEAUgR36+gt+3l7xMZZE0JHeTxsS1PLNcr3vhuWH
E4PdEQMyBkbT9Dz3wkQwGKFOaBVk7Q13DOrzD3Kj5CCHCX5L/A46PM1KwwACJeP+bCoVruwGKzXK
/utIQ3HR3/jRxjzQnImbnvwnX6uEAwhD5/wFo4VJA4xaUSS5reeCUn61rvjR+HXMsWdgTbhMVsBH
0Zz7T85jmGwW8zuxB/W6cmeUemHfx9hd63CyOeaVgvKKMJ20vPm1ExdFuXKMAWSx/d7gY0NyP/4d
6k8wTCfhlTTm+GcULZXzVRviB5MJMxnp/yn8GTURRgoBcR5bhHxSZu7V4HuBjgv85tLDGiKF/qEm
mO48hZmlovht2ChFmb6Dbh2iCFi6dg1QtIIX+jAdquQDOE81J6zxUMr5JyqEoLt0q0tkAojsL+/M
bIH4HkZZ+pNaezhnt4Bl81MGZIoWad35vpZIRrA8PUYNKKMc+zwAA5yFAhNOXmnCoi3mBw6eXZTi
WnLadxJT3ORP5GEOzMw2Xe/hADdw1aslnqYCqnaegJhk0gVL7FOYxJbu8tHE+/fG4YOyhrOtKkrP
E+w5xk7UdGNhgKbzh3o+QI0pkCfFIb/1hzhlz5Rt4FYPtdlNrin3pX2vWpyTwCZXNU33e/gFMmBt
PGkLStSq6fksUotLl7EZXhoZnypIB4lGWJ1uZ8FXyEUjx4F/fqkZ1rX/cmjapnzcWifO6oKFmAdK
7jANQnukWDd8jPgr5g5uHFj7tBhXhkZg8MbhxT/1dKo8dNtGUP/yxEkebof//d6dPmiiQztz2VTn
9YEcPNsj+iRBq3FpY4mI/Lznxj4bcvybLJ8miXcm5VcPEcP/EZFmRwKRKRDGgA6PPn50DIeOPchk
YGe3R9JUlP0/+MQzkl1dGCIA94aMznI0mGMrfsmP9M9wxA++ddmUarIG2Z/dzmRU82ekBDu5C0Pb
OzhHfDqgwXLVke3dDx7GUojIwYIbLGyLTyiTimnnjb5twYLefH6iTWxuy4VP6nMMU7OOXIziyP+z
a/B5KkJ5XA1kmkCjOytPMaJUT6hgKKaqjIeRo3OpnCSwKOWmkqDk78iR+UmytcksisJ5fDqP7EQe
gxwMkIiQ1FZZOppeEE7RMtKeTEtciTn0tGFEho34pYt3BzSWjxbOcqZeArJYoKWqNFdjG6hMiNxJ
0MFmGZ4HR86baSJFu4mH/jng19VpJAyvC6F8h34VIRthVxKjHRoVa/EfQp6KYy6tbFV/bz9aK6XH
15RaMvoPo2EMBo5E/06Uoen26ZboiGuXAf947ezcO7H6aJ5mRTfuigHnpnTmfSLEwSevWeDYYzLY
RX6BDKrBcWJALeOqu6gObK3+ASDVm+Duj33eJvINbpGTDq6R7g3Kcs1FPWnWkld1yaGPUpsFcUB7
+2Y3dXhLLAQeX7II8Cyo9pWF17Qsr141vxCJN8wK+a0HWASRE2WyhjgtsJ3/EmRiX9OPZRx2VVL8
O7p/06IWvwdW4xb0N9oMbr+5UdV4INTmPC41nb3AUbY8nLGblynnLO7cEXJL9wlv9m6FytOfwsyo
DXsqYfcNH/+b+8U1aTJHiOKgB5JRJNBDPh3oHeHMPbNZcO5kqKJaDlIdwCgtgqzyzbXdiWltGFic
YJbmYzFWmWJLqHPTeVtxCzuA8R5YrTMtKkTDCFO5mPBpYdSEAf95vWF1D6Mcz5bQqycUpky1L2nb
AyGEv4Szsu7tDR/I2gyODAiHJWsInZEmFrLuGriliR1/Rgl7T/slixDWB2t5fTJ+RnQNQs6Sd8u7
OSmu7sUk5U9l4o/g6qTmuzdUJnon7U7Mbp+kQ2f9bj73vZpIUiyM33fuQP5AtmwauvL8cTk7BQHv
rixiaVkC38Inr/PK8c8Peu7kdvOLIHupz7smZBH2nMaSBcUYNWNsPd5wnMFi7qxfE+bQ52S21cb+
Bisr63iAIYP35/u6R+Mt3/2t62VTFg8mpI2EMFIXGuxldAa7hRkm0U5W0ORqoEGeKL3VtnVuxrcg
eKncMmKlJYO3UpMXUnmHwJ28DmT67gOg59X/WJb2nquqb8oV23tBWngyIgtBBb1y7jB1+gPBsuyR
+d3Uu9iXgeGsUj0O6m2gNnvrbQ0g9gHWfy6CMZf1+s4xE1BA4gNtsZuNHQQ4ORn9/F8tko8UzLWY
UjFdKuDCEMNdOtQZ1RmSPUjLhASagIOZsU2kERkAEXFVpHZfzFRjEqL0t/KDj8yh/bg5YCnucahT
WW4vWAKuZ2L7m1mtenvrSHtdCtds1GYy5jtdx8WzqWFudhvexAOjpgb8S8nl+zmPH0dbIlqJewkc
ueK6ghM52hjhaKoqW0eqJXzPTHGtScaiss2CJ6PymARVnJPSQ25PGMFqr2fVE7M9koqMcSXfVC+K
k06rRi85R10dsOO8E2ijULUQo5i7gbBpb8MO11ZaR4bIyIJhFr73uS1k9N9ecvlrnOF1E+dPIins
ovgW053gz40suMrcDbmr7/yZwBtvsJ9QqgKteCPrhAv+GT4ZUjP2i4B8WVx2gi4D42ihP5wxSN75
XODw9J6yswNV/9WM4DEaUmWCvd7S75BnE7S7RNuY6Gxx2h3gzM2WA4ukHAgr9XZ5qZQnGcvzg7km
64kl82uO+vF+Pr+qNtlDnp6hnn/GANzetYRdxz4onjHVM2zAuRtCJLmV7xVLUZ7G5SwKl/bDC0mu
E5P2jUSvrppvCAmUHT8aw8OKjzDmVlfFlQIbcIeECTI04m8NfhvxCqSB9IcclexaKqRxt7mbJ5Pn
m0RA5eVX1lSy7dBEfDm5McWEAaI1c3Nu6gLD9xyl6Y71so5HD8jorn92qkVylCGeWYVimEi2U+kB
eRrQtDOW0iK9twdmQi3vq8SqSN7q+jorbYv0vittmbFbGaQHL3wp+uXduTi01rUALWGsBJz3IOB2
iTfJmioUxEvYweyfcqNIxSmwIR0iBN02c8x5Jt78h8UFftJ9PKcpggp5KdlVgKwzWaGWqgeoHffG
TvVm1TK5ySuKvQn7npDjzpVxPf08I24Cd2lbvdMWt+ctVbmKhOsTD/bo3ealiVyIe78KPousI7al
+XVkHIKX1zYpiloWgsjeazxgtYVnLeemL+ZhlCysQNEaAr27KOPkbVAJ31xd96Dqowrq7/CU4KRV
XyJHi3MIYdAV/R15J8JD38JPXK7ueUnBh/3tRW1UZbj+ysiTR1e+/pgEKPiVS37PFK1cDQYZOA6m
wLQ5TFYJOpRvxXQ6M1Ae4tzzIUQH6J8+6jxhocbeVjZZxLN55+PflYPV4og0XcKrPxrB/ej8lJxT
Qq5bwkWjXfrxbNxW/nnNcnU4lwla35lRxAuzTFrFzqmA0qCcwUML4gyYiexgQ9S+CB7w/b2MTrws
Qo+X6BZrlJi7+ZYtwnCUe7d/KeVMCY8UFe6zv9CDsIbcMWvehbJmJz/3jsu1bh6qmaNMW41hIiCn
hcmv8cCsikOj6HiCNKn4nrzB7dWfw0VIHPDoGGxFrEriIDelwhnbVwaDaSlR55KGX39jZrzvLFUa
oe1gPuAFdvdQ6iPXFI20gJlVjXHqNw80y/1FseOjYfCNFHqjybQwzzIgIh/N+azj+Sm5RmJkBt4u
OZB/68TnBSGKqGoPhNznZ2By7b5LlLOJLhdYSr1MDu2VT8wKzZVvKmFfFEWN1EVA6v+JxvZREUoB
LRQJ6IahgFVHyfkzXxnKv66UB4oYLHuQIu91TEcwW7GmsT0+/6p24wmJnDJ+0eoQI8xUkV3poGxc
RNiWjB+4j8BjNAJC6Z9WmLBt2AVeKWdmlwtkw8VuZz9hXP9jSp0583ZZzw3IV+bD/iln2cK/dD+P
oyGVNNC8GQRVbhEgqKkkRG3z8kAbBBaftWb0A0fMwLasqVY6ucxAVimCv5t5GPpVONudPSFBymzn
mHXTcJbQ55d+PA4uJl1Sw5usbpK1yJN0x9fkY4Ms0DdcDk50NZB3I4y+BvQxXZADyFM5JbxzPvxW
qcN2qat1wJlj6Z4FvrU+GDgq8P/Y9d1odM0/M6iTFHhi5NUf/9gO1MhT4P0scrNINEnYcUk24Kys
UKkYiUVPue9JstiV3LN3YNqOwHFawdGXGyptVCOsDUR/4SU9grBrlI4KDDKaR2G31XTUWuz1amsG
4RzrZF3/omZx8OYavmhzG/Ep0p67f5YcW5l3z9q/99NxaQhJu3wnWRacmeXwbypLsKsQ6spjGBnp
P0oSToyIHyp+KFBryxen1ABcY7/1d7WkC4Jamc9I1dLZGyfsVS04p9mCw8tFq8t93BocVUEcDHOZ
dJpOeufDoizGG+O5MBxIValzgkj0DfTiRPpatQNaoH3LXjQ5rhNTSFZRLhC6vn4pqPQ0LJSGXRCj
8faSX8mA2PepPNJRI2XWprR7IG10BGa1jAzioIwOrB+BnRUIzS+7HHJnXTCJ2+ME/0z1dp4fFeEK
23UP73vCt2GLgrTmqPFVQgApFNChNQjp2pxpvGMgBL29h0Ci/8hGe25p413LVQ+qKv/ew15xrsuz
ENHoXjC3yrN6wDz2bLMiK6tX+V1Oa02Qu11Vsr49yGhr/XVnkLnqjrVLAM5TdDQTMLyr9VbFPE81
gvD01d5JnobcJNZkvoa9+IRymWi8HNy4YFLTEVpAUR3LqzHtv2HhzBBmDD5r5X6BUkUUvkeBOQFQ
U1cxmQl3eljOMZw2o+l3IB/8FKVZPpPlwg2VyUxqWyS6lj15QyQVBAX61WkMB/ZTpl+wRBMaD65n
ZGcx02p3s1bapkgDVNx2Ik/oDDBtMoJy1fhubVGJFheeYJ3ZH2XKxtl+mGgmDbsFnVBsaO+Q6LAu
a2JV+5t+Vh5Y/WtAjppLJjm6tD/9N6wALOBEU9HXvmfvk9vyIFksyYTNqRKwgmZvQA26vhW7bsPn
DMXnevAQNm++SYsgBFIUVwFBdrezMEDa56nY7kl6OphusekaUPmPOcyA5Lrxw8dksSzNgkdyNRnD
E+jZD4EazbwG891EXW8GozkDyMbHo4zQhfgGOICQioJao6X40htpw4PabnfuxjbBQ3cVBs5NkoGy
ZOy1gL/dE0QWnaelZecwRwr/opBs3wiSoJfjwQoKUCL50WLl5sC0BWDIPXG4OI7mRHpUNUbrM1av
TFPsT4fNAyOGUKZmOjWAUh4ruZ0pqR6G8rcmOMh+TlaxkHMY73+LBolMq8PVZZj1UVJZeG9nVWnh
pMz2FSHiyDMo8DdJ7KOcQeJE3HZj3btnF8M3wAEf6C33v3BO4X+yNiqZgo4tj/L1ee6vJ2yf99GK
L1wurscpUWhsFP4eJ5OO6TFT8WBKLjgSLqwiofceTo+yJX2czbPGfv0D7QJp3JmU0+ymCwqA0Te7
Ybbx1jSqvuIHMY/tpyF8BlFOvfm2Wiyf1PajZr2zd3QwjfbCPofqBsy3Wadb2TyBSrCoD8ulsq6I
qp06skIZCjC4ulHU1hHf26ovGaxzrETrQbYu7QTS5HDKWFhHCvYxCLcfeDPABAhz1y7L31U2JKz9
UiCrRU9Ma1y7Re+MNOZGHBbfGgfNoV7XOozceeDVBrV/bsf1C6JNBaVHNVrz21XUm1/8QlrZAQGP
QsHwT3Td3wO13e2srbb7k0V2eg9+0CF9a9Zwl36yTwd4f/wVvWC7JkwJHLCg0eeAOJWRPZMxwNt9
IETTsg57fn/3Nt9N3SfUAJ2SQaT8PIQzSVe1t3Crl/ZxQia2ABWMrxoc7Xd20K4vzg5FZ7O7Re53
OSHpG+AOPRhLrMSUBkgBuW6zTTJMLlKgxh8q7z3C/UO62jvQpW0ACry7VzXSdxYXWn2qUfxpI4xw
YuhPB8RlZIR1o2Q1BkYdKjGQdIgnoTE6UNHrFwTYMFfUxtvHxS+Tn213L8SmXpauuN5ZgPxZNAmG
EE/ScLaFK1HraMcYyj1sDLZjba/4c9VXKnegRF7oaOP5wc+XJ9qT2tleBt/TtAhx181v1XGS8kW1
7C0bvol951PYBgEyZwnsWPLDHEZE8n64MkYLFHnMPV8hA6hQeywKxS+4L3qyaELPvDnButXz5vth
ltJ2NyBAxg/IIitSdG493Mzkusaf3j3YTKc1VI4Gi+9GqEi8FQBuiq69qzfb0HJPBT6BkySbpgSv
WZCYNa/MGT9lwmFEsIPUro5x1b91B9I+b1s92mSlHXI/q8tNoywm2wNHHgeHvVupRM43KOT+Vy16
7UXoRNK5xdZaLscDv4QZdWFxTy2Kp6+aNXtUMS9xpEd29JtV6RosYDXrYS5zpYh2pY/ngmQE/E/9
Z/0bkFstWr8q+52KN3WJDhtPa97yzpWIcdnNFnEFx2g9jebhz+mutThlJXut8fsaajUP/RI3Alls
mzvCek9/8AmN4/xSe2Za/ehMBq/phl9Cc0a/ObRKTo5DeMrftQRvbXWspfFz7g1uL1YchbHbgvad
U0pYeJbat+wK7/sJl7yUSfwHbUZ++gHpbgYOTdcQsQI0R2lKBTpYg3PFb3V3blz5zTve7TfrcZCL
7Boo/FLfQD/zlqYBEy/TtE7d4LvUsqO1gHTCalwWUwRJrvwH7LGoHWKa3uOUXgymNwYa45gRv24a
9GtxGVgqIN+3FVmf2UBihu0Hi+9+QI+FjRdL86aRt/pLPMGZVw7qByi0fcEpncFd7iLOINw2k6wb
ZCmHcsQAfUVT17jPq15iowhMxwe7TH9XQsB5cTY4bj2R3OhFLeMQDjs9qUZjcY1sJERHtBQPN0Jp
KkMRXnFANPt+ZRTRvadVReeKdUbWIUuDaP/Zaor34udk+2FQUZ63LhosrlYiodb2nK/vRoM/P9+r
OB2AGQC+xBCHRbnORkwOqIcQahqIYqzDJfhlqlhNKnxK6X6o1qvp4SO7Men8Lm7qaZDJacXwbKLw
7PF84ckq22gx8LvFnI3o/R30HNI43asByhnQBM+in5E0l/OEwxXSkd0uUtLNfDKGOFqDUAU65ywy
bEhcTvrEs4Mlxml4HIpL8LH/FQ6sy6SvfiZuhg0Gx3kE5iXE3jGbx5qlyu4Dljrq1ZfwTehMHqX6
DmrHVR1vSYoPXYw/daN/te5JksiI59B75ANqkC6Ar6cVkefTAgWG8foq7CC2loJpA981B0VMbELu
zunCCkgO7kQu4VCM17DQTMLRXudXyYFWLEfg1Zck8nJQFLrTAUlSi3rJDbluOTfa5Y3mTllxD1s9
W0FaiYx5Y77x2ldFpuqTQXtKMXCsCTXMLScOSyojTep0BXGQLcUU0KCxYKAd0LAZcyH7OaF0jDPW
ZbqI9plIMESBtpGxnbFNWurRFbzDun6a5Ck75Sp/djD8NJmIqZq+prI/OZ2+OBmTu/sOqeiecrDa
arzl56u9Ero4irWzKX5fTg88Uap+OXd2LP3pXsO0ArB4SXAl55288C16LhDgv0kqHUGAMrQegK8B
CVqOk5B69lSIPsQ7Ialk4IsXla9mHZGhUInwy/JMyeeWloJNgr3F7aadmp7KhYZ40KBCmfG22noV
dZYDz79DTNoZpYkahQuKjJa0r22v7EPmNGz0izB+Mvqyl6UjP4UkbT2dc0RmH5aUUeeCMbBQoJ/J
DXr5+dOTnHabliO32pcYVnCpPMGFp60hDTSyOmzc4Nf/7ftma6eYJ5NEKhtM95VKAHDl7i7Da+YU
yvTjxfFSlnBMKYT+9Cf3q0UlYVb+2fE794yjJ2XU5D2Rw8U0d5WErqyfk/PunmUXu/2L+Nwm6t/i
tte/ZALkHI+j36zUPejstUkkn4ha+GRTWJPgBHeL8Vgr1xWJLUjH/b74P7Jfu5DPRXVGIXmkrekv
CQEDL0TDrw7rULB4B7DwDmqfKxu1LTWaFxO+2OwO8QfRCR0YEElReVP3v32jMHHtpTq94eB3Gyze
nbHEigBELTnblQMJc4eNsPR/V7LcdrlAIYUflJd5kVBpYlKpKLgKmwkMpSmlm4U7ehqzDMr4ePyv
jHg5DZNNn+mE9fyVNN5OdiTsSgHrWNKZKk5jKd28Ziy5hXbpsF8O3sZJb5OaeqcDODPdsqZ7rS9G
CSD+CDwnXqlMTanPZw6LH7ag9c4rvaDt2rZ6RSaKbt/cSM7VUc38GjE6klPjpyh01OrVKaPAg4QP
sCHHsUehKqnqdcbW+/fJ4TBHe3Ecwxp2WB3xFFCzz24YFJKWREpXkBxsC9RoaTCLfY3/S8Ok7e8U
J+FIIy7SpmRxchAjfmPfa2Vg4VvP/Hp/iZcI4txtKMcVgL/U1qf6M/7xQKRYnjuIo5hMRaYbZP3t
E/ym9XkPUjEoi9j34f612sE9+cFwc8QhfiGqIGKE5nPQkH6k5TGgeSUBINPVUVS+AQs+BmjasOWu
Mvja0cshb8FzXT2Q67sKhY1ZjVE/P7bQof1acmhOnblePqdT+WFI/NmjuQ/kCqdrnhUC0VmwkyD+
iwbjVinsymtXa+UR4PlP9p/I9JP2u8LRBmxqHp3MfqjHGcq5G29s4qFMa9iOB+YWwtTWJaWrrfGS
3o+1UXJSqR/8AyNobhIuzESECRsk4MR28v0qx6WwVZcCu9/X/cp2XodlF4w6MrVxV6JqgZ8bG43p
ORmQDrC16QxpXRSBQhyET5KwL5bc9AQc94735KkN+zV22CAPZBrjmKbtB5WEd+s2yp3LCrZQdC2y
dvWcBKiiJht8bqy36h9PGRkuhQSg6KsCo8N9pYJCYUGlsoOXtEzApA1F52JmL5RPNURZLQ4eNEBU
yI/Om0/HGuh60/qxfHRQv+aY7puBOrHTwMYkw7VApEIuZYu4mQQdmuAI4szukBhcnJSMoGbngy8j
lT1Su5lnbGb62shFXGjR4OgNMcNwkeNNvcdhFZh5YfdqElfi9lJshFcWZr/bJW3rP+tRQgCccUD9
X3dNoCiY51UNnA2Migv5xUHPa1OiuEq0izhqa1cJ8r0q3z7+zxU+2sK31yBfSNCfa9ZPoar9lxAh
lur/rpvuu6/T8tf4xhLYYICtPPqPU2b80mUXr6jKoF8/2yfmpKyhHk0eK6VTSp7jj2kXFooc02EH
/GQg5Roo5FS2NAg7MAzPFNPVafQ/wZeowe0A3y4eX4Y7siga8N5YHrvwvAFyEeZeRqELb96n01vh
trZoat79CIpMZdLn5rVfg4SFGcZzRZNSyZl/C2fJdZGJhsOUTC+FdyiE/OtC2qBveztwa/zePGSJ
uA66PlqzNRBAqssEMYUFZ2WZ/AujzXAe25jhfJ2K0UfQOszMWXuk6NEWmMNJRixjMM5wOub2T/An
rTxaridnQDqlE2O++kl5aRG2x0JuhzxPuTjT0Pj+a6evTkzh9OaU6SRkImSfCb8sFsmPyqRzEEq/
KgWddpsZeSyAMX97cnNWV9ZuDyScOUQzNIYgWiUSVynZYr5kDtG/xuEU9BIdSQL3+lhb8viq9KhL
RxxER4VVNczjUmnAMy6a3fxQ5CD/y6/upiDjhxnJAnXQoSgR3gk8FQX5hl1f9M9IKFEPe1HytDpU
9/7w/VnWkXsHkEz+8NCdwcb3oc8wMpa8yIcDU89hrl6hK+mec494K5c3EFU+L2rDwd+pmZZKRjHs
opEz+5R/5fHVvZNVRXCOOc1GsqBFQKiz80oN9403w49dxwAojlnVMcyvR7RtK8OFQrbcpHILSt5D
VLf68qQSp6DCfwYKCQ85D09A0OxpGpTggvh0UfyiSnq7jfeTEL8Mcch4iFmF7sgopdazJzU97miu
AJzxveywp3sTD+VYOQsW1yFfrgS2tf0kgwX6lwailn5MGgTNBzqDg7hERhDCXk74owf/kbHqzG/N
BhmcyuD2IaXXqaIfymukXdLv4mnNf/dNuPnLw7uBMnl29kFT/+GgCCjq5Oh5sIZASKJr3qQVp1Kc
kv/DCLzUQTKFJFN12AoHKn6ppM3YFZyPxpWsKFxWuz/Yo4NoDs1gMbPzc3xGcDYZYcLkZpoD28vI
Jmp/coml5rUGSUNFo0qyDerJM60hHr4vrpkJ2HXR8w2LiSybV0xb4xI4mEErwlBvQ/ZJIH93UQek
c0Zb6MKJWndNgdrwfzEl68VnmOcI09q/hz7QgS58x82t9UsnxL3PAz/fD76MXftCrM+UGeIeNkSE
TxGKx07sTy5+u1zUBCnmkhnuPEK1DwUEWZxjnlu+EmIzJtX/YwhsNodHEoY36T6alweGI6gqWhOB
6fMog9dQ7ps7+HMXg0LehyCsKxT/umltDrJLZ0ZVuyTymrOD49Z0LrBX9lChCWLGTd/mHVytuIQP
R2WoyaeP/RnETbn5jnUwl8T4nN6ndy3SMbeQSOMpbaKEInQystPCybKoJjN4hbO74ttA5nUHXT4V
3JG7EMOfnFGepFiwldMeYsiewpxZAKvwisV6pwJeW+yHyWV+sifYmoUHx8dVi5E5emwh+zt0NDtC
HrK8qVC3RJAcUwtPVI7B5lI4pfktopvDJxfqkSWbsr/F0/motNa2hVSDVmQJZr1lJ7KmzDb28O5q
Q7xBqTibgWiaciAcgrD4e9Q4Mw1jWSQ2WZbb0mSexnKrG4X54bCR8UUK83XF19l6zmI/WpZ4gJ7R
R47AnOK4VzRlf97sQoM18c8MKSIlSRfrjHXO1x5Ob1a7MWw1SPhWARTbJc1MZgi7inpor/BSSh3M
xtd+jk0YlQ08EQYJ/70K12VMrBW3XszGRml1yI+EQ9gDbjsQV+TOSURsKrVQ3pFQZzWdVcXxxcbS
MXPV/s7J8zKeVTDUQka6I31lyuilNGnjaQwm4O9PILZ8R/yzBGRUCxUlgZx9DSD7OfkaEWS6QHvE
/Wsh9Dc1jZz7Rjzm+UzSEOOfYgeXc9QcJb4XaUgCHu0DxwUUss5iiuTdJZrNp5HPUxYnGiOinRUx
YgiVO5MRGo8ubKsa0+n4RKV2yf+cviBe/EEG9Nrci3tOEyGegB8Yw/YKcLAafC2pCTwpkghlhKl8
ea9mImadRVO9nlSoosFr/+uE+wqqUkj1rji5tNXddacrG5Ro8JKt+jcEtaAZdmNe+C0oC3qUC70g
dBd34PFx4zWsm/4ajot16jbs0aJYKexxv98ilTnxq7v1qabm1TKgpQRxPRCxaQ3y0cPXkvmlrcdr
n4NVM3hF5crYKdguMIDArnh/bje2yL6egMIgVTl6tI5n/jecTWuvu2ZWYWW5uirlI9axDWtW7ZIk
6l/O8u1witr5L+CUB56hKkWTTFBdoDZUp2A+wq9JPOEarWtQSTf+Bg4NkxTvZ1R8Xlra8memi+1t
Rf6rAPoKflX2SNAh2KmRrV9ucLAxCSFEWUfIIMBLS7SYXtEM0np0cm49yteQGSsXkiYSmYVd0R6O
icF7fzhgidbz84p8Kfia4Y4P8V3hTODlExbC99wcDnsWYFOTTF4fsWzv8x32IkRoOn9WfhuZ4pED
Xu86ivglrLSSCAenKf677/tVBWgyE0HrUNpmT57QxBTbitzgc8jeQ7JM59Sjwn/o9YVJ/6DkVhRZ
kajZTCRZSdigt2ToXwk9yAFlPwohg/zKKpjzyw03P+hwtuReLvchD1mihq02E0eUncAwuQVhURag
ShJ/OSXdk1KyvfwKqt/inl+CBdn+aB1qJpeOohhDQTubpQy71LJEAJ6HNipfrgMMWEVslBSD7ew8
G+vzTxZPneoL+V65TkNsgEPRsIrnK2561AvUozyoGCdgMX/CQF5uZsfn+Yk+R5AvM+JjEgLPyKhl
NUBFO1j3hmz3mZ02wH56yjVnOjOVzAC8JhEDf4haJ2t7TM2/5a8MGsnocmxbSlrXEKPwyAibHX/c
zUFcUg9DiUzH2+rXPbCi5aJlfu2/ccWI0qL5kl2CEvWQca0dUYYdFvScUXzuu4o67o6IGJvMh/x+
Y4DH6kR2dWtOIZtktzGNlOJscQ6zbSavhQpae9ma98P5zLrE6LVtUqYRf6rJXTEXlP7dwx/eMMjF
G6msRdXgGp2CUG57UL/9+m1G008shoxB7reCqwJijL2DXU2kL6Ni9+rVUx0iPy2yc76cq6ZYWpzY
CvwqH7ns1u/U6ZHx2Fk/iwXBI/nR53YT4S08I9eK8r4wzfh1OqaJhGLAP8JaI2eVJRpK5LUTL2ab
q3eT6eCh2Xrf2zGjdXpKpIBPByqhK7rxXu/+8Ee3F9pQvzaNmJ1DL/hLhBrZ1u3W7tIpbyK7HVeM
K5ZiTY4KbFnXhS43KzTw9gFHseRCdAjm+QNp5s9ccy6JDRAIY1F8l+FHlryX6BIAzuYtl/+k8ZN4
dqxSkIT2NDydwAW60H2hM5PF9fFL1GhfV9NKYfplI9LW+WjGkjleEnLBOpbPIlwT8kqCK8Mcav51
pWZqPfT26W0/oxzn+ovNuTPO9VCs77Q9ss12yx8TKKIU+9EIjOfBttFlvG8i2oQ3iUgQGy/IZGz3
iLTm9nM7MCzQP4cHnneyNInPWVdETckKHwRvbjS/QaNYJRrhmw4xZnWMLlBVXP7KX/htss1yPs3c
FkV1RmvKaWVFLNy3PeIuYmAtKOvUVogHtYio2t9zxeI/cJ1F9jJzwdZOlnLBK5HnTvlU1CnyItNB
OUcNl4ODHqilpMYbaurCPnOjppGv8tiakxSQyMefp6Dn4dWBrr4wjrI0eFWaBCh//b6KYdC51xs+
inRI1CRFz6izwRPuOw+vOc6lEVC7AHF7hmrJHrAtmWdwm5HLV3tw08qzBwfjgyGjGr273rY61R4S
raP3JlVxIew8nDJVZXJFuWufPl9X24UlwaLjO7BkDQguKBcmcxEPwyOE2JXwXNSLDz9JM9Bs685t
UCcPZbWM/gEa5SiRMwFUr1HUsavA85RsFiiHtkeupOoPDkFPkuVlyC19ZayrJdGAQMU8WUMhyfiX
Pqup+yy6aNK7xBP5H7rjCuzUwHC+4znhJ6+ZF+VOIqVWNqhv2g4hCDaOOfDAdaURaa9PGkbVBm6T
vaNWo17CMpBDOsB4hhO0eu4kfYREIzWiSOy8E7lelzmn6jbG7ICkxnqWIG9wo80ZkUXGEVmo9524
QpCOukuVybR0SWItyRri9HUJeZsMHnc2TRtXeDAzorr33Gw6+TyuYZweRJp0wVevM9fttNAJ/nGj
aJ/z42PEAmhQV/qe2fssF6wyW/s20H5Z/liocPcfk1Pe988zrCOa5a73Bri9tyqs+elc1QH2HwvG
oiJ0u9qWdA5ED6Di+UVhjEoa3a6xJD9QoGvGkBVz9q5mOmqdhh3S2PldGuWzKE86CG/tqg3aISyQ
cUffqeUf+qPe3zWMv/w7xOwagVoHNv1bLUwVXvhSWza48u6zJXM5E4yH7RKtNhcIP5XVioutAh2/
tGQEPIF9kGJFO+qme0mqYyy7v4Ufbfc1yakM3hQT807ihqar/ayuWNNP8QCdzyhmS7iEvkx2wNZJ
+qVUpWIY5XxVRa+yn8YfXv60h2Ezc3OdcBTY3wGeQWBYNl0rwcQfKEziI0Sap+bjS859pLQcn2AZ
GNvTSlOCkUHoQr6QJhWEx1Bxn2XTST4cVp7WAAKp0atEt83n0KWF3Cn8bs515KbK7CkmENnG0kmm
szPlofuYknjo2FBg43NkBLw3+VeLWR3O5egw5IuPzqcOkuwfNwph9Q6SgYHExf45ikH2OIrCAyVt
6oQ1WNVB1hdkL7/zaBzZvvOn2mJkE1iBhBktybcOEGtpAZhi3G98WvfXnFVBBg8eIn1Uf0Ti7o9b
zORT0HUKfh+Djzf+1QPS6ZrUvGJaCTHi+R9ruWLf0NOuwvgGY/2W1/Mw3UE278vUScoIMlavCNBy
jBUBs5YaeBuOWCNTnnkG7BVTA1jzxrbJGySHe8jN/R3AADW0gn+wOdjLKYOmoLtPbPxfFqHYLi3I
v7AaNxvIFILKs43uLJ98TZ1wWYj+B5+CsHkgrzV8ghT0mTT2Sdw/42nzmF5CuFxJbqvuRMNf7VRJ
L7aAgg3aVOcCQ0+GVrcSf5ZjTJSdxkcu1Y8hHdqKkdFK1buxa4cmHg5kGgX7OfYsrIdQ12WAfMJX
jSthNczvkUM0guqvaMwiadw08Vt54jkL1xcHHIPLyQyCB3ZOz5wSimoyHxwBlKMZJpL7VxgTtFXA
GC7tb6nnITurknS9JfwoFMEE1b9d1tp+EIJ1/s+tICPRic9I6j/AwWzkUwlpkiMKniROtkTTjCG0
gOSmJng9jIF0iI7AGvsnfjjc+PrxW8pLSil27mi07a+CVCqxILg5CnvlnQ+30+35YSWJB3vQWiQ3
xrjVuPsQVvIMUlOHSstvxclIJQr1VqFqabqmBOy/807FWCgduTO9If1N9wx3U4SViFxxFMn63nfM
lmBCOlzrLK7MGAulBr/Vin30VtEwVQB4c1os4EI2h+v8GHSh254DBGunQXR40abVOi+IBMpWHLYl
jbQFMGAXe1AHuROxCgXMkdtG2lgbpxs5CzVWQNAwYPaZhyS/KpwF6gNnpXiEvZMv8CfcT/dDONCg
nZ0dLdtsRUAX4U1MlhSfv0J19A54CcKow5w+S5NiBLSsYVpNPgWtPeLw9afV7yBjEyRW56WrcmAA
Z1oo9EgiLd5ehVdvO/43nYlq6zsQBo1HS9wIxhENLL1gctNfcZWn3GPDTqHqD8yG/kmQe2RC0f/0
uv2Ok/DZgOfoCQHjLKRz3W9osWW/EaP57HsY6sH9DavtUEPiBv/P2e6nQdWgkmCV5vv9HqIAFM4Q
6F6F1L400benczLeIWYmz9uTAjKbUJ9zBtTYWBMKkXOSzKfyn6kTcMh17HNXZ9kyv7DrZaFOQxuk
gIZ11rBiE2i0gtNxeA9nMTN/3wCy2S2Sv6pqiRx+h0q7OwS5SpM71EuszwgyzQlGfN9ijiOeWdUZ
hDEz23hbPzU86mEKbVRTq19ZPJKJdMSIG65qiQrxi7TinnuA4F2j9YYywNn/L4UdqszMpPWKu/pg
QXUJ1mcoZz1rPlcILX16HK1QiwpjrB9/lf+c6bvtWf4icJJGZDBwMO4Byo3EOiO9Nsfh/Nh/49re
BZUpyhUB6lfoivP1yFG1zjNkmPBfYcqhSsG2bsbzJH1FQeK0GjdAS10knv9+SDzU0qLegnlpKWkZ
QX0yCc5E3pUw5b5jdfrwgEkVYHGVcq+p+baGtYrNUEjeyqciB7NKiQQPTeAX/zPW9rW6EqC7iRe0
TCgf8vO4L8Yaf/kkrA8zAVvOfm12+Pu0240Wo1oouzv1sf3P0wFt1yqztbfM6DI56WsrCCazYYD8
yuZaPdvCOTNhdT5/ty3wK65413rajhc8HRxdv8Pnx3qV2mwTgVcNhtXEcU978K1zgDAhwlKVFGDF
NWh1FeMTyfmEGoRFuuqqX+Nx7kG+96EaQfgOSCVO1z8tAb2txahHgTz062SCapc/T5dcZOjCeRyB
eOWO45wGJ3bSBsXHhUtGCK5oXvHtlhWT24gwjQ7MSxc2GwS6IQbWH1Wahrv6tu7GY5S39xfMqtXl
p3imXdHXwu/LJ7gQdZ3+9lJmR+H8HWHcoBcUqAs1Sbjx3lvdArlFnXBYFMc3CL7Guz8rSTN1W6Q6
0LLyEc6zjCWRQIySP55EvqdR2zd/7JMHnuiWUn2fZI4QH+AnASbkNjsp+GGl7QFXpwP3phkI0CnT
fVYz73aw+hIcBi70d9MeDGPRA6GTmX1YmlnJ9K8KDKwezqGUkEyf/oVxX8AmsaD2q2Ou9ZpDDww5
rMFIWj5EmIvmTFEEqsnoljoter0oN5Oc8LFDQzdEQuhpgYlzZ/VA+wSZ7zyvVTCPml77khUVOrVW
vX81ZRAjFEu1CTt29ztW8KfrPFlGMhXgVrs/RjwUPMLTSNV9PrZy6PssEi5vnvqiyCyPwflsI+iX
1CzGfY74Td5if7J9QqH5kUnvRc29SPEoIUKfpL0J7ypdGjfvyV9fujNnWDviLTGsfTT4m7ys070f
OrxLAbqo3rcwmgRj7CEuRMMZll2WZuT7Uq35VIV4YCZEu7HHT3OQTrPW45NEZm4MkCqXINvH0lFy
H/A7uL1YvFelzlEDI1E2XtFRUdEbRfczuJ7czPdDT00oGzefDuhWAYokQm+r/ApkyV2lrhlFWGMp
Lgt7Gndxv9BGRhFcF2PkcbqlREESamTTfhTw6hNbIsmKyncoWvLYHBSmN8NVfl2iN6HSqPUNSWNv
7V16Xoi6qFP2fYRmTrYk44yu1QAR2ERh2DepkIq2Zg16gMq6OQkCXcG9B54qm09jEhuiVzikMKML
hTgkhu4RiOz2TGyYPQg9lU9E8PWuzbadoex49DCH+LthyH7ZukIwBNYXPsSDYO1XjnsTExCb52sN
D5EqMEvSvyKVjTnqjf8/7JpmbQqGIyad9PjQa+U9tx5i15VZpLH+Q71nUJRWKtIS1MZWf9ZaStV7
jQ95lPBOrqWSFT6PbzyQHPUlhQ/TEkyBNjbWXIB2pt9auqDx5KPjZg1uTjN5sX9lkQiTE87/Aair
fby4k8dwV0AqmvEZ3LzkVij6MHDKm8KIV3zARCr59DfArLFnI7xmr4rUVFAlsA+Gth2U2yMmf/cT
hT3CavxZmhdMfMG+Ym4R59rEpXo1maj+CQtbPzwhhX01xCv/ccOgnKQNh5V04CjoMHOkK9Ztw4C0
QJRnc8VjPEAM0B0jP+PjaIm6RQ9EAWQs5kYVUQYzgjylDkQ/CgKx66efecvrATWrKfe8iJr0z9hP
9bDo9BDryZTvY0XZ0Og5i7cDY8MeUgALgXIH5V81S/Ur4AqGwQLSz0Ohie7DoJl/6BBbz+JlZs9u
PMWjEwIbyEsXnWqLghwBApyotwmSpxF22YqM+zSTnhEuSXExPPbXmcaTADnE1EXeiM3dcceQnHZF
Lb/HotmBeJ+47H0R2KVpp+gWtVHkN9GS0W/OEXYJhexSST/LoqqgXnuQ/eODDTCoYaxdZJ+PSkN4
qTu5iEsfg/EOzmM9UwjUA+C57nxXxjMGsZTKSMM9XYh2rLX86QmPmFBFk4BEMPnFN/MfQAKUAwWh
WrskFQP3+5bQd4SEjC+79LwL67Wy2wq40oW31H53FJo+RD8DZnlD9ZB3nzCvLH4ety3vXCWpM4iC
I9LtDACAK16eg5TQ/zTc8PooaPFpNBWefYRfIZpp/P0IXPYgKIQMq7GNi6+3dG3+MT7M0ddv/EqC
zTG9sm/aHlE6F3L0vTWNLFnnTX6Enu4SWjm88aHakIBtAC+/SFJ0aq0ZbGz9bzxLmYHkvjnF294x
NcwYlo4NixvbY6kiyvqsGO3wskU/SAZot9vl/OKARn+Op/VBR/YdhwvwS87o3EIAILcMYm8h/VPd
mmMN0rVoSpcn3XimslTPcMPybnZqEmsHs1KvBCDoaKmz3E9t2lgY/rrozO73FK3t0z9//dTjvsys
gbYI+2uEZDOTLsc/11gRqP+VJ5lFeEj/Zc+HY7Zx7G81EvpFB+0tJEI7IJG0wwnR6t4mrCJhnmMM
RbMNbTq63s+jq4jum84DOoZWhswMrIns1Rj1xVVv01j6VNcoZhQKDwj7YRPKSfP3prhwKuUGNtRB
JLRpAk9l/bhYo8Dft8/43iXpBqqDmPXVE0SapFolFXlxSJg+bJ86GaUC2jhezI/z7tlbQ4T6dVIv
0CgvLNGEQSQpb2a8QLjb013G2xEPCG7PxdQCnRuWkHNK7m8IeGgjriYqOAWqcWFKRwjmh020EYnh
piuosylQGalXR+vO62xP2ABa61JnVXwuv11EFe/UUfs3Kleh4//9s7Yx7D+WnW0iTbGUAU07v6ly
vW0+JqbC5k5emnBseS942eoGuQiA5JdZBTZ2PsQzwvJOOFQRTVED+ZysuZd4O+ZacOmCMGHePYkP
wLmba3Fs6WMmBfHSEBnU2yGnjKtDbXLomxXy8mJdvcepeEdtbiIorWrsmdgjsTjWRQc0g3S+pCnx
dcdretmLDwHdN3j/NitBE0vfVxS3liWhNxbkEqDE2tDO0xCxo+19iFLWHUrpjTov9X7xGraTyFGf
hpx+7BzpEU4448LfwGm05qpPUqzCsI8LcODZZt76leoxurPnOi07/6pfpYy4iveBpekpJ2S7WUeD
RK7mRC9+4pegdnOT6i1kJ+vjcCK8vWn0seNSLGuPhuER92uyytmUPzQ+qZ++sdZSDqxK4btOg8vd
Y9/zbkfTO23keW6lxU9Q5BB15qFCyjs9/sZNC1bClG1uE3mcqfsgmx1WuJWOvrGX8uT1UaXMrWDh
kX6T0t+Od40MNyYQ46R0xkeyn1UDrgmzScpb3TicqStp01NBl0WKhenRlo9uBsc5hxKplJ0n/e5D
CAIaaTU0F0CWhaSp8mOShEbsTSCAhbmyMOpJharC/4Wd3qo6EAxmcdLr+gToEv1l8wp21RNrtntb
vIfSqkGp1NF12VYzuyo0xV/FckmUW0UmlIUxRCaKVxK+SXlW7nsmRGMzxIhJc94TICczhjTZBMz7
7awVWtJDqJEPXsn82K2qr6Cz7sou7YAvC4ivBpnillMVZQeuszWRJUZjLtixX2O6bDj//LoNvhYp
O9M7pxF6ZIB6kkccG2pI0/ScAVkOmcTKy1uyHImnwWqN/5HrdeUjDdnbKfTyvWh2jFvG/WcX77HI
Wk5VBmEDTRK2WGuTAJ9z1VVXl366NvoDh5CLArK1l03MPZwWW52FA3vyQe0N6rurGnN+RP2gMIeF
2P8USOk1hiBLOOde3pdq5IFMd2PaUwt32dF/1+J7/i+5Du1SMPTIJ7zgNyN2FnfLsfMx6VXdOuBI
W706unQXZha3cFambYfc4yOH6rAEFOKC49LVsWwn7bTnavtvjU1A95irRYTMXAbdf/Sm/MUOI3gX
35qfu1kKDtXelyG1t/Ne5IEvJ9Uf24+OHIl4xBZZWROqBJlY15KIMWpFbCLuYL1G3ybbEVf34xDo
nKG+9b4KZ77Jz2PmWaj6eskIGvIk7MXl9muTqgRWsqmm/8d7IaYmMCudkKkxyQvGDmho3agdsFjp
gD2EhWFz9UGZaGg+AE+udWOB+aAcCd0Oi1kD/yDyIu+Swj5XP5VYvFvmYUfwmDI8mjzp4YY4Avq5
bHUPFTklPxT6n9EhSJTt39fy/b5WgErtDUzDszZDPsUEUEf2yKp6Ox6OuTupPFpWAD+YDoGbnPvf
Bm2kfWO3Klqt0MsJIK0nxktxejZJpaiMBGJvtexRsm/KI7vbhfC6Ex2/y/SNGRM/dAnLA08P7JKe
e0WD5wGrxIYWot399ZMltWwPIEi5LrMrVkYrBiD2Xr64kqs8BySYYEUeOsz7u9T08CRUHj2ZDgHc
hM6XVYw85g1GtyNdOn3Up14SxfK0QVY8AZw+WlgxAaP9/ar752rH0jI0wwG/KrSyVhC3zLm8UnNa
oO9ujcHLV75WLrjaMbekY5hFCsw1rY0anG3EqbGZKCTnsOlbEbukgH1CEGstt7cKDrAbvaMfw3sZ
6y97/fht2E7IIJW7Syt9HHThq1YWzTvyuqDQetGMKUZat7cYZM3nOoRcmpU6c3MUx96Rq7xYdB1U
mrDBy3DanN/w+ars35Y6e41HbSe3nRT1KTMKbEbzZHB8HX/BhpehWIgGJyAU4ftkVDLWvmK6WUDJ
chfCgSwliF16811+MXNOm1XD1laMPwCQLyPVDRRgNy4zuEUb24zVZakFFZXFALBA4gAYb7RPG83H
YNp4ND1RgzoaL/rbpe2AndSRxYAv/y6bgu6uLOkb1w/qrmPV6AVD0ilCv0yAHrK4V2lDFOuCsE+c
i1rVG+1O/bouNpzs50bzPpoJgfgfRv1+RY2TphTSYsq2odZJ7t7NUjzh9peXJjhWIAPW+WlcWa6e
aOHPueD/p1npezsF1W5aW8O3Yp0W/9jitzEnP29GunUDOxW76qHeT7EkgoiNSHgGmjJE1jghvwGv
L3DmS1eiABndi3UOIFjJwtcHpdhLDYGkiosDNzY5cPBhX8nmUhnU9DjSH5CPeI67NORq4aqAqEyg
QpeD+U3vughKf6Kv4HhaVsdqYXz0vVf2JBfdEW9YERyPBI6BxJ5BybDxSd6eRLHsdukBDOfV4qO1
I74c3t6TZh6WuibfgH5hJlxF3Zka8nAu/gesvfmYJ+ocGcxMmWnTm9ARJUVNrIgDqw+WyAL3Rlwg
Z6VpcolwcYY7lhyxbnhVCtPmVrpw9OH04XDIjXWB0FUAX5zhA0ofsAmO4aXXFWR/4qtpggR8Ir7N
og39tmZkniW3WC1tyhR7Zbc0kq3ikTnuT9jNc61CQv6MBO2/HIlWBX12hYGkZOHcnA9ZBGXtyaNb
Ex1IUNyzkDYSvdSTQvH3jZ+UM35NRQnCaABEmNaUlRG2b+8TZE7QD6wQ15KDXL383xd7d0gDLcp6
JzsURs1PDjVzo+1QPOnzIFkAyE4ET397Q1ktNsp5m/WvnTUUrNmuH1wh98rIg6RglbntZDYMR2h0
tA4pEfFwcGEimhaLlfcvDDlnFRuAkrfnasX0AwmEowco+bF364OcIPoxSi8hrbKGdaOsKCTBKZ9y
tdM8mI7nZk5L73/eC80iepkvCKcctHf2mfufO2RK3WkoGqSiE9HX4r+t71ZlRNQvepgJ3floCUJY
YJy+eDntyTPg9zOHThtv2dt2zipm/FUNmzM8/Km88KZh/6/47li6HolSUr1jOU18qlg4a5AzfOuW
h5J+FMFbBfVSY44QQkZF7aTHWXrOeylZ7rudNlhZTv3h1x/u01T48FAA+PU/8/LHl/YVYMnImfl5
v38JTiXD7x09Ax1rlFc9Fx90cxgslC1cBBp8qh4ARVP9ecrfpYzER6FCTh4wG5bh3nWA6yZuf8/K
Btww6354j4VTduosegtpVG4rAFwqcGP631ODymFT6TurRwp1kAurjfJLf81FWLOtWc9H74hlmLZi
cSjC1a/+p+mIiXW6YB0JBlJDWMubNy0ongZzhxg6i/8XxhQgYGB0pbXkiFQ2Rzo9QLPWXH+0DVF0
5mXhXvW+QQI7CdZWOa+rkc23hsABGKKBzbXi4l3irLZ3kFK2OBWSUeth/d0FUra7xADUMCNvIcCR
At0YVf3vEjqyDc0iDbRIWdOZwrcWwPDqkPfvPIU0yutukhPKzWuYCfcBBf+B+mKl14x+Cgg5PJSS
sonWErlEIVbtfIiUYNQ35PfqVIyE930Z+zLAOJDVU4KohQ2dvufp2NFRYvIH2+1ux3rtoNFEzmKb
6YGCtSBapn5SsBYjGU3aWjjnQVzxL6jnydbbnSwQLKVplstJ8LydgHKJe0CrzLh+ZPFi6cAAeMgp
VwMG0OJUShN3JxknT82CW4SwCb8+KirLDuxdC3QbXwd4zmlZaC9MbSRfDTfd0+h6b3Z0FNYVng4O
wfk82THmroxI1olOwazUaaHZi1AKYe7uqmPCgpO91mmlaJPFbPVnpU9yZKsqo2UsZKpNZK8lwckR
3t06OhFsDTDlTCgGf0CG3JI2GZlEw1x97CxAMDQcTaRT9zaym/lpiiwqt0LGPvT/k9dT2OqYsmFt
Mpym+vGhGLouveFzS1XFgXkWHU6MuIyM157piYa1K+6Mc5YVxkKSG/Xa/HXtyMDTxqvuADE/BOqG
zo87wzWXkxEFJWbF9ulVmpR/N/65CMe60CenYnapAMI3VdaZ1c8c0YuFypBFLLhCEHNbvMJvDByC
P3TWKPemrgUYVp5yzvah84kR4p12td3QP/uPwUHmW6VmBu/SjRoojJO2R7GMp1upk3kSIM1DNpn/
FVXlxeUzSnhfvCr9TqhDthpa3fA2CztTHdJiyG3zuTRSTblsJVTpVcj2d+b2CpXh1xD7Q0tSmlPh
kg3/+tLSl5mzmiPpNRGMpllpudQIVjO97gFBYbHeJ1e7+6wugrlfSR7x34yFvNXOtpMydDAqX14m
Zm2yIcdXJly0OuYXs92Huq4lsLbIL91s+ji7QMBR9CI/9Q0qW6nLLahrF30pwOF90rMFNGsMSpQw
4D+q70f+6p+g5jBfutSaexGRUuriPY8kc+axtqK71qss2gTQlb15rb3ZswVOz8ndClDqY0/OsWkF
LKSXF84vvMQ5PoWregPFbFlEAvwyYmnl5gO+vvrRqGI0XLcIw5cwEwAgp9VkjSKaOP7YflrBH9jL
E79EF83Oe1vBJlvOrb3+XNOvGbBWlA3FJGcpTGbHjyLUFRhO7Ast4D/WcyQE79hh4rREmzjxVA8K
JxB0zUAKTXD3bK+FAvxYlkYF+WOm4qPpksP5ze9gnZvV9GSHSwtWIqPSQNLwnEpW3FgzuIhlKyft
HVeaArmieIR7ySdPUzF0AXyr1SKCnEBnjnugjeKX13HhHG3zQXFTwkvRoMWvRQWHILFaut9YpxEu
7CyXDd0Gr3YJbvjwOzKTvWNB7Zr/Rf22S994duPLbFzQZMwz+36wx2e2gL1jxZbv4gu+tDfOmCvD
102dVdkWUBYaolzHMtE85ojZy/FZje3PJjQ0eJ6x1VXmrXf3yHoTZ8gIFy0KVB7V2POw8WmUhQAv
h1UzU6Gw4D1AAHuBJsHOmKY+4uopB93iPREiZ2qYz3pbG0Q5oxONA1YzI/Y+KNpMJqumtU6U47Q1
SyzGSj3lEW+RVdU4B7djFW3XdjdgH3XaqDDpWZDn4LwKJMJHc6BT35QoPTg9ce4Par83wuRLeNMi
Hh152NfD0Paxj2NKV9ERX2xr/UkX+I5PeHPc16uvEw479yVN2xeLm9T1WG4zzCuarFyg1KNtjvZE
htYtUZU0xQoVtkdTPdCEWbAlWV3qvkEQ9kXs0obvu4kTRiSCxeSisd0gCut0L3xD2xQ0svG2rfDf
rabQc/KJZm/kDPq4CemqdTC/+mH+1KMYxVadWN7GOc+CLDJJc0KpaXwxyErmjZnvztbX/swc8IIa
LiL/EENGe+5ZZKDQA44wxEmbdZ3xfFfv9clLf/Gz14VfrddBsgL6P83mMR5ULT0JFy0H7TUvpmIk
jFAlik1rm/D2bslFYzINQTMlmsUmyCsv5rGhreO0TGZKCD0sUYE1Uom8VUpUK5YCQUaeZ/64V336
4Eh0pPVLDrTsZer4PmFUFvmszPWT64RN2eYyUXf4Sa2X3bQGzlLzHMBtTmk2t0BCnHzRb3C2dxD5
9Rk0S6fjWQWnciNomv/Ci1E83nUVnuUtlPYjYYRpaRzhcTCN+vxy2eDcFICudrrH6N+qrX+WkgnQ
jpmb9kEn0nmUG6Cw190JKe6pYP2A8TjjFgGFWuRurLo7obhfMOs0ZXKt3q/euZYQdtRq2JqvF3xs
d2KSJKCo4UtjLZTL9vV9TQkcNJh9NIeLDL7Wa7TnCghZiJ0OldQmqzoZ7mWFiGVNlPm/2U1Z1iCD
V+oOR0N7sEVOutdEY7s5qTEfRXypcBa970g3vtWyMc8aB0pcBQH68beuGN78pEYnLXvs2ERf/rWV
0Ig5AZ2lOYw3XPOClzvjdgMovkG6oA0TgTwKHLfS3QcN8uwVrcRYCvgva0qQwDzbAlShpWYg7xM9
ux6wO0oKp0IlCyVBge+8zowGtSZDVnl4dJZqEHi1j8LAliYsNjmIFJfd/cCcUIA9wEZG/ObwQvTt
ltBZtxi2xpGif6TWQ2yS07a5KIrVcN8yg2EJqzu1DCQL5UpVCO5EtYHgxrB6Z1teHt0Fg62+olv5
A7fkN0qrHL9xEpRrWITam7nQUHsCulikk8wt4n1EUFfaWpaFov6tAUso8bjxLXyrSvJOom8sUD9D
0lbpuEqkTfERkEIXRUUYCO9Qoz/nNha3trLdckPzt11m4J+60O7lydce7ZAHS+uAZyl3pyO6MK/j
+fpUtFucTdnYsD/lhX3J6jLxpZcnmY7KgeQW9JpLPveGb+JKfFmkFjA/J4JhGu9UnEyL4eOA4W28
UbLaC/YWeiPCQzZoFZawAf9yOFQCScrsQjqd50tqpt1x9telZEZs/yjiwQc2gr0HW84LlS+l/kQ+
EgVQscZmtrQ95uVwxRlILvUB12fyweNd3BFd7cUcXggXiwC9IZYcFxtcpc/DBw7u5KSn4ZZBNN/I
LgGnNOV/CeawtCO/ovkIimfY/7+81knJyWxxAR5I5VhMBJViPZuzLS3nU2bt6lhaCT+56tHd6JQz
IDx7fnTBLuoQTJCBgiZMhcXhV40mFbUirhO3O3B+kMqLztNcfNpuG7NV4bRnoN8kZ4qnFF0WJKs5
G2iDeKO8O4QxBMZWcxgHq7Il8ABCGkPPc1LdT15lFDClXoDsoP/OhBQg6qMO+9q3dKv7+wSjq1rg
tIINIMl7kz17dg1yGox1/hhoTTKeKjh1orfIntLrW+hxAYcryC8p/EJ6sZDEkowl3a+43NqpK0nE
9stOP4y25NNntv9gfpa15QrV6XPCUKZcD725SncHpCf3O6DvnN0AnRoVkUbt2/3fuyg1F8cIaUqS
Nd0I11Gh2U4bwDL/nDS5686jYlmtoK5cffm7OGw49xTMSOqGtApVqayXJGqOHn9pjfCYmQ7EO7KD
FhhCxgrdYuorAhEYUU2IObIf62uCm+WZLNe/8dt4sQCVK/r2J55oTqhpRCcWRKhiBD/EV21k77yK
kiX/v5+jhgQAk2qgxain3vMflWJAosYMwO3loHpg++HLZjEcwCgAhusv5ivWTKv+ZVSx0O0iN30A
cMWzvnAeYoPxIxKJeI4ggQS35KThh7fZNbto9wK2ZoQo6bS83GE/jwDQWYnyexAJ6mj9KaWH4Sdi
SKDdBNMEelXv40wqEja1tSsuIyuRz5h7hUjDQ+Opz5dDHMmL1Vj4tAe1nD9mjZGSvT0/RX3izLPj
RNJWGnU8JJ03qtgvakMfo7HyS+lYTEEF6mcc/CkZJmmV1WjtRIhk3PCNgV2Nwc/DilteVoEaI7FF
rVbfjTJeOFlVJmmPnfS8g+ak4iexe8oP3g0N8Ij+p+FDxc9XP6fep0jCUWoOfYtEcMkMOQK4cr8e
1SA6qb8DZbaI36vBV0n00pUa0ITCsAkkqIz6mdcAKmZcg+35sqH7naC+eBv9CKNnjG3FJ7yCe+MI
U+MNSGeFU7M5SSyFZT7QWhT2wxZshywU0ZQX5KXIAmxVUbnpWNQzcSr1AhFn4no+Qau/iKGGbi/a
6cNjWuXgqfEyccKsckKqDaz1Ja5cFroi82KeCcgeHjE/PaYkQCKhn9/2OFVrlhND1IKD5td9kBj/
4XYNpZla1fLI594eiXfHTQZGZsBOk/e46rPr5uJZoxjnKYgZYTT8gbVpui98SWL7jP2yEtSBQk9d
nx1IsbXD/lXlOGVBir/LvjM8r6JF1r8+mqlCWG+Tcff2Hh6yDRhfRbF4Dl6H/rR2UdWZNZsrqaIt
AzLAKzkUqPyfaouT7xbyZRgoWrSIEkRj84+R6xGZRLTXa2jBimMAHtOfXw03TZ16H7GYUmBr7Rv/
9hc4t2qX8kW24cy7DilAifZrewzCozo9oEH+zps/J0RSlkuraRHRPBIDiHgB8mhmbcT4M8ZnIQuf
9xf5OfaHG2TxrqF0+WIhiQIkYlNxpQSEYqw7exNGwdmakRBA5c/7r4SNm4qPB6upnOynjraPOxRG
VOS26E1YdbFZSquUstPg376t6lnYOyQ66+Ys0CC0AhIclbAyd6BK8QaWvUr4DJaScvPEHvDXHgky
6EZvjuoPa4uzKgRpLER4TY18ROUYCLnXkM7NlXP7nc91L14DP2nXT02urhZJyvlIRZhapBwD+A5T
/nM5UmgG1Ov+t716Dc6ppcyGxPUHb4fVdhbypNTYDybq99SHrDXOfEyej4O3lCYKLekpbaRTqsw5
u73BB8qk0PHi6vnc/1ypvzCFZwAlxJWilJtKSTEX1Deqkuvfu43V9bBw+MfWNm5HB3fm9c0jEwhF
n9qoGjM3cSBjplnbS6yYa+C6RvWt+/KMMmcZjlQfqmSH/paIFzm9W7tf/WO8kJbOzr4wZRt5FzoI
G+LIKY8GX3oU5GyjB7sjg0xYrR6KxDR7uucsn50mgRz2N0mZXanSTUvWh1uev29VK18JmsKNLH7D
KXZKBbllmOrCW9Pr2IVp7VxsPS6F19h4vSThaINE59gaRIQahFPcpYmvJaYyJAbZZi/I2Ggnr/W6
yNm1ozoLrZ1TESOMldg+kzmhM38AoR1+BgK4cHNXnGnnMnZy68qPQW2B/ZPUFh1GOXmpdnDh++Rz
qx7A7hYdCc5mYqXWmhaajzYSUfPDTG972K5ygNtW5unyevD4ZeH81+AthWrTZag/koz0TGjCXtes
qam1QfHZxO/oLkL3LDFuAuYbzdzU1b2BHke7nkCwa0V+tU0QQH7z75hTmrlhRcvnOYr4zmEfJWN2
Elttkt4gdSgG0HS8qgrf6Jh5ju5o08dCyXSdo+9Kl+sJtEzIivQtQyOXTRLd3PueAMM/oQtbV0jE
eAA8DVgWbhkeMaMWxlEe0T96iYi4vc19omim9cRn2qv2nxXkcYdmWRzAWWHvFGV+SsWm8ndv2weh
7iI1dE9P3KqzhX5dNXJ4+dI5KKFs1VbmE5ttbFUbJ06BYKOYHPhngGaHKhx0lE1uU/OSIm5Pwpqz
cjvALl9ELWhc+qK1v+NkrLGykZ75eTA8ZhJoqRl2IrY1b0PO/odGH2kD8leI5UwypeTO+oNaiYb5
jpiJsiJcIPpFP5j+GJrIGAmESXsfxtiVghMLxApIrFjp9jd4TuT4LqyTSRG1TUNxrwzGNecZyP6g
BMnQ6HSq3Vu8ymqFa0IMzG8bVkxqMgCJcXmfhNb1+ZYzVp/mVoPNdqPnCm3re4cOJDMWx6ZVliYC
L5EATYsPzPnmrz0bKc3mGf11qbAdHgPgIot/56PmnXagNoHGaF/FGiFyUZOIcMmextfiyJTtWZHI
vqjhLUs5HqejWLjdBQO5h/+XuJyhR9XSy3THKShMe9LH/5wHPCXWXygaoX2wz4d6BR78+zaTGo4N
r9JJ5Q08u9MKYNHYJXd03HOtHmSY6G4vpdk3+EqUSLi2TFmL9sTZsN2o7Ow4KDx20rMtq3Sd7vXV
3gA5D8/eYRCa9xmiiC8DRGS/vceo4Kmvpil43mZpVL96Z/C/LKAIg2aX4MUfSKfcvJtNabCMqTeQ
G3TNhbDvGmsyrJ74PyCausIQmyGx9aP+4jqjW4rw1BUTcauaOk7dqVe1Q0NhpeQjd+evSXa49xUa
ltmMDh+JliVlBaFMvY48a+wX3cyGd3Tqh3UYsWKE+MzMgCo14DXfFPorXF6OKQZVJLVAUQYuUy7H
F9NxGRgmywtnLo9wiyCU8GqHhwc8RFhPMba6sXW0olGjsXbsCtBKQ5XfmHcidN7zxiWbZYiBLYUr
RrwonpY0OkVlBieSQGEHrzTubwcTDdQCBBhcwvzDdwy1bMTF9chVk9ghPh4S1aXKdEv64qMzPxKI
mhaAxrODcoyHT1R+Lqiy1QUNFhZn8okWa6rxsiyJMg5VOLr+vbCKWzflP+3rKD28kseAOkwzKs1w
rBUfrZHUuzuEYbZJHphEem/gwE0WG8LNu9QEfatIt8YhSz5/2/UlTohdTVFHGgLwPzf1yjJWI7nb
Pq8E/sQahxn/3Tgw425p+JGwHr8t1jeVCUgA9Ro9dWd/wsvXh2hUTLn42/n/im50i5Bvi2h2mlCf
Kd5VVCAxUCFZWaqb6p7KAzRphouF/gNBNN97QXQv38j/LXr8wa9th+1EeoXnybgEJFU87wSAxJxq
fVtYEmB7bnj/H2HSB1qyvDtD/qQcj1rWwJxe3hPiBcdy8rBHeXsmV6CpNgPN6nmDeMOI4T/9KOK/
fs+ppBGgcMMyV84sUC9fuw6doDg4AWwH2yOLd0jlB2KuI666nVyqQBnL0a3ZoBma6L+qiUzDWGwN
/gjraQd1Yqk7fT3REcol7kLsSLEA2f209NIEyYi/h8VrnyRL0Hfq28eTedxr06wGKsW5ondwIGJ7
hxegN90tn1es2gwk4KL7kksQCZZZDt/NSt0E7mPExvtXhJEumoMa9Z0pOtJPruGtSaF/1cTHK1+m
Pcq8k/aL3SHFV5KaJcJTOheuKFlHRpKXmQ7rn50keb16lh4rIGrlLPAkP3ICMNogBYAnJ4eNs4l3
ob9V2MhghJhyVytfSITkU1pJ9Ja3gKZosBBC1JjLZ20meAkN6GXkuJU4SC7fd35+rGOyC7LVhYOO
KFhAatT1Hr2uroLsbNUgdCULQ2U9lMP1t0ZK5Rafv2K9ix8VRuYGnrme6cJaoORpyC3qmEnc+Z91
R+cG6YZB8TPyaOgKS5+yhvA+QHgKxhqIbKxytoLTrle8zGYSaa2ufMsYaDVseWlU9z0Vyv8mMIOd
nMerjy8dFFOTw5qzpecECKZPjktO1zTOU1GFyU0kdL+t9RK7LfW3p00F7nYvIdwvDELACQDSC3U1
7wkNDfMzjvY+OXpplNp5gzHACNPV9uyZUgelDCxsi0D1P+7+yz4KZ9lURmo9Hj7XTeiBrtO8Q9FI
TR0pwEujS+dz60wln7JaKOV3CKnVnx6k1Ohl5eJVA4VJsB10vbTA0eWr+2A/P/+NnzErt/ckwXSy
POJooU/8wWXFzNxvefv6QVnwxscHXKZ16j7DSiP3+rqCs5DGKhCq90uU/WBfaBe6DURf35iBmSD9
mbwSgyy7ugKpt7n+9QPHlvPux/WW0gUh6BqsiBPc0ipRl0iDoMmoQD34OZ1x61jjhUq/Kt2n8fqe
q8tvfJQdCdyfPKfOp9OJQo8jm2mDfkUAWJJLhoaTAj5YqQuHV+JkKgEczuq34NXyout4WcXj7kxs
QiHQfvGULyqmvKTl5FlI+dj9fzD3clAmajB9n2+jo9HmOv+jh5XR+a9KQeNKHm2eBmCS2m2ibiLL
i3S2/zSbB6zgcIAjm0cG1YGKRh3wOyUXRuL2Yax8UmmvuPmpHoaVX5lYIsPNWTBXynA+9Q8poNYS
ofX6B9CAJgbo9svrkjAH+T1wqXgkbjOWqR4/Kz5YQ3mf4cYn0k7qKLN5TNIekk2avnGGZ1Qm7HuN
wDBvPMHXfhoYs9uY7UXNJaFnxp3a2cfYloMrvUffL0oKLwqOB8RE3hMFn9n0nu/wz57UHyE8rinO
Q9Z6rB69kUwwoqJ1X738zQhjlXYfx8P2NELibgTZ0UdmWIA0C4u6nzTjUOxmJ+ktaCNYqiB1aaRi
3nPOR4pjggxP9ABAujVPgbFxOyB0C97OJfQS4hKpBidpidcmZ1Q3o4HAcxHXK9FXfoXQDnSIoJ9f
Ngb/ULWT032/btmyZp75HIwfzatp/qbh/1kXP2jBclns/UMTa7HKW2noTybEML14we4obqZBlRuf
jfHQkRz3Xio8l6GQeWVGd9ssDYOzrc9wPKTtsCoIW0/kRA6puY8nyO4lyPwnqlH4i29m+S7CBavy
p+eqXNMbHdREq2p8QUkTpvU5pceJ6GBXg9HoOxElTnPAfcOZiDQJvoVNNatLYEmDf66R/VAbJsO7
xZSB6aja9q04kdqv39tzH729mpo9PI1WrSrGOP/8qSUE/Vjfk2wwUlLRHu9H1M6JLKuT6Si9HnD9
ptuWK6HzGGdi5hfLTak87iZ1z9hBb+BZOCVhtn7/VNVCOw+ZGpZ8XQoKAveKhyMn9sX5+hVoS29a
+9+L+8PGAwa0yOWBMfAacvynJEt6+5Vfcw+c/ySforPDqyy+3i8ly79Huuk0pAVNIDgB3RwUeOpa
evrniLh1QY3pR0eTRlxiePVBppNYRHDTvo8xyxcy5W4VomNdooFCrXAJcVeWFD+FLgvOwxIM+PDT
nHVAyvOam6Y6NcdARyiH8Fms8n6O428fKEDeFQYBwet0ss2wqscgEtMqfD+G1B4TQSyZf/vvXGDp
OriyTCDTMzmz4a3XyPNyKD1xDJZ4pscNYfv5khf18DeCl420xFGlxsIYWRpT9WS8rBcBwu64JUfg
oSO37nB7qixPK0v9cjKAefK+Dn9wxR3ACjbUMFP8KPR1xd+N9mt6tVmmqE6KnArARixymg1kQD2+
v0xSdLpnfSTu8dxIm+7Qea6+vwBZ0WNWxOhP6EJKptuECaZcHJeM1CZz6IpLQTZqzNn+EVxAe5eP
iakVgwk0uH2HZdn77/v06rZpJ4NJgx/ehxjmSmsd3FzzHIjegVSqRt2/3JdznazA2qy3MNWrIXdv
pUaBEbltrKWzAIGPqGuq8Db6R1rmoiqbseVre3sdCSU24oA7i7Pr2dfb6tCpsQOSnVahXBlw45Ck
gooGiKpn4qcrvKav+XSDJY5CPgOTJATNkpb6uzvfxhOlQxB2GfoU8T3VzyVriucCqVydE/FpicdD
2YSe3+tXJSSmqVXMfzKTTGLiYWzvEI0kOZT0K546QBMiEMKzSsXsDh3BcHIBMwXpSWKDxcYpwpCo
hJM7/sN8sQfj8uhib+TUVt9/EF5HmSFAtTwv4AdcOU4Yvme0SSQUM78dCOwcooPtvGy3Gq88g/tM
19wBB7d1Em3aIkAYimOAH8Gl3/Py3b128s+BShyYYq/KMF+FOfLnB0bsULMi9Hy1Y9rljN07Mpf5
zFMAxrfI+vuVzJw/fcl38+NW54RvZM2rC3/m7t0Nyn1rwkZ52/zYd7ZMeDHfqKNnQmaYhxLlGL8C
x24e4eyV3aCX2g9J3kBwRdSvtmS3dLm5qd16gF6AfQJTzJhzfwzPF2ZdEK1/AgBGhYjrm51y5Gjh
n0ySQzMZ6/PRlUPlcTYj67XOf8bK5Q0q6i8stKfIE2IInbrton5Opp3yUSx3vVUYGm4/L56iypDx
gzUeOCRD+avli+s6FS79F0qK3AIsBhQ6a4BtdXso9+ShJUvPunc+8GKRNfkPjzYYEdEt7iHNj1g0
+jxwHgrSRZJpGEc0hgd9WhWyaST+0QNRCsNdpqZul+Baucy5oPEH4EF8WyzakBUyyYQjPRcNffk+
FhNhL0K/BKkpNWPBl/6A3w91ndPTh9jER43Xq2pquEbgxczB5eDYa+q3aa86n53AiGLZM+HU89Cf
QZH/ExDmCfRSrA/41L6kWkUl+OjC/52LhnVmHLMckI70EGL5F1ilcRGDlfyOiEQ5rh5gLuCngpcs
S0dcaCjIf293DfgWeuVAhG1D5Z/YTd9Vlv32Mb5Y9XQozf+DhT9ehZfhpYTPpQ223U22cC0OmdkF
0cJvxdwuBDZoZnLdweSuG2F0cNXpPmHjQ+WbVTVWa58GSNKB4wovOvDyHP00kNW1E0FqhwznXJHO
UO/K5/APCI4glnrkwdDC+0elxsR+IZNavgJbm8xeBmRW2UqWiJxjC+7S0TyYXA8NYqLI79NMWlm4
WVv+cCKaVQ0YojJn8iy0FxEtqzw7YNMhAjW4Gswa7TbMmlJPlIF32g/YyQOjkChAJ2YW1xBzJ2e6
SDXAhG7yMRhGJYnrmgtx0fPQJpOyYXlZgukW5ZYuOG9CemBndDhOevGPFcL7y2L4e6hwrvId1BFn
EJSeMJBr9HQHKV7hu0a2zfhRfdK2KvyQzAlWwh2YlBlh+5psp5De00Fo02hMCfcQif+l21umscjI
lSvS1XH8wh8YFcLaVzEV9bJkKgVwPjCoZVQKuDN+Vf2mPKIMr+NlbMR14BS++4aNPO+7fZVOB5xs
EY0QoZd1EaXcj/CuOO54B+i8Mqn9ysasN/VQoPixePd7cJ2X0qHbE/KYox03TbEpMi0Furgol85B
RGLFAQJFnDKmv2RMuvbXUK4mctwpJJF9NajS6hSggnp7AJUdVuJC+/T8IeVmwupSCzm7Erjelh+l
laYN2BrW4uOXQwAlB6Q3ZewSkpPvwQcbSvGdZYk98vFnZZ6xAEQJ8F025LaAjA82f1A1PxyBFEH9
qonFQyzO0TXoiuKDiVb3OoQ39JCjomK31d35q0d6gYceONU04Jp/2xlSnDKFu7azpixm/EsaG3YB
IlwtXBOVn2FY1Va+XicPapOIV3DD3ouSlfKUPSiw/of1BDocbFTf8+VNHxU3PPOo6r4GT0h7YtiO
HksWbZqnhtxPTZUP7K41DzQSA3IABBIp/9si3/2DQ1GQF2ViJBZbAEoZwpxUwIGMkYAXTb6pkdi9
kT7oqeIuo9m3pX3W8fLkFLYLNWDgTRCh7kdJHGdt9SsRumrXFQQcvhssMJTNeYYQQ56qkCIN+ss4
wJ2OtlvGOInMWwZwMKHpqtc4yt3svyNvAYWV1EnIeqPd2AuNiX5RoB80X/hDhIXKskrvRoGYcra6
zHY+Da+Xn9FKtxPyYMlaMY+c3eQBZVX+4mvJkiBUg0RKvlGCkXBWC9vcy4HW1cq8vebcm5WXJ4O9
vqkpo92SRraTzWsqpGVwmST0JmnqUasb7a/EfWDRpcC3wnKLhXxwywq3Hbv26xBQefLteCjhXaq6
yElUByvGPT4Ybqm70poDFcGfyvc/fvejxP20+0qDnVnY1ruqpAMOfsim5BLl2ewOazToKCcKX5lm
fkbd7M9TNvumv5s2LC0dKEnjtm6ZDjHCVMn9W7+gnuYuHeFOGtOXosEusOHOil8TdclKq/q/OB9I
OMesVFWgKI0GZnlCUrM9UhYfGHtpxJqxHwih4kOa1f8P+D2xCFPWBtsnacsSOVsqkETJnM6j7RIM
vIAe6ddBYZe1ZKJ17R8NK27R2TL3EYHLbQ0YkIPk6EfeYNiyvckwCFBwB/pNuiOpUfFA/B3iJNLV
9ZItpaK+Wjjv06k5e/M2L6HZq7f+uqXcApblkD9QvqwvCaV74m3EKtL2jfZEaG23DIofgGwxCVE+
ZlNpGvR0xPGWUkuevMXPN5+1Te9PAHbQRxIB6M4N6mxxPRra0PwpdCV9L0TXKmAnFwKfjZfhsBeD
IZMchlYrJB9Vck8bybAfLQBbpsb7Xw85ZCeLa9kjgjD982rcL4MkJOJ3LpKjBu/feTX3NfbVdAGd
LNL+7m7GV6FoQ45FFrK2ooKzBOivmoeLGPR9Iye1/7ouMSjwL+cxr3TkthXP3Je1i77EhgWjOfkM
gZP3uzh7pIeMRFlDkL8Ln5lp1lcEUe9H7VCtGixANc4+Fun3GJmcDMIYoVJkuhqOsqwby2mF3gok
Ay8Vxrt5CM2S3WXJLxf/6U+pgTDXR60jIvDn+S3xdzcuYe/KSsqMODmQ22ievDHCLhDk90ftUfN6
EZ3MeryQCuHk2NoCJYQ8W1cBNbev85HzVUlCKrIhF6gqSsgiEHfp3aQ7EJzEVC1a45l+hab2bJqj
bM0mCQ0qZJUyD2MMinQZMFd6GmuvWoKeVHKdGp19LdmPCA2rIKUPJtqWn+Hhmn/Imv1BBjPQExpq
93W5RZJ0GqV14EsAg19Nd5vadokgw7rfQ/6moGzBDbzHbpqEujvcoF/d7tXx/RRywEQpNvUAacX+
E826j5NYFuFhYQPy6K5/1ItAiE8qVc3jzzqsiSCU78uZst80/ndYwfmftxdVvuRZTCodKbVO9uok
NhJ9hxSIOMOvZJLDBfdpzfoMbcSyh1TD9+TUYtDETG4zTZzZCEtMRz5XlSK0boOMwQhxmXNCwC6m
TlsKgZeqSmZ9bj1r3OAOR3M576MEO7matzMNFrgnXhvSzv13+/fA8/77+0Ql8c1oBfndARfK02vW
d/uJ5Si8JZYJcJmy6h9OjKLtYcuqKaC587bs8q5AZFjtjMI+wotac2xX4muGlC+Uh/5GwF5+X1Zq
BdzvvvklsLeuf/1whupgcLvvLqN2a+UZ21p5ktj6ZXrVBL5q3Gs96/LFiI5SOwGQXVf9uUcwl4rg
DzvltGiek9ed7BKQtpOODlvJPrZkvBKh4dltmjkvoapqPZviumo8fhK5EgDTd97QpdHuC7UFxANG
0idxrbqTSS0Bo/0i2HlPPpbF/ChzMVc9VXlzS/K4C4P9CO5yDVSikSemsM5COjwSbvnQN234tDyH
5fdecc3ixCU/2aHRU//avz9KPdEmOgdkSKb8BgZTM6CdedXx4DtvJMTiQFDRrlBsQRRZBO3Gii6H
bc9KvcRLHRe08MgSoDB0w6g0sqUujNvFi9ZIN3Oiu3qmUjFsSMZx/dw0R//ED5cljQP+gQKsSGwM
ZWNH4VdBBze2BL4iqtxfEN7Gzy+uYKVVi6qPWFEkRIXDYDgo/xuzc9HNwzCSD5LG/sNzS0Aujhii
csP3wmXrF3yK/Oajw2X1mdhi5pGlQTVu+faM47r2kkEmm/AEEKWVqn3dLVaa1e+2SwGv//uHa5/f
e9uJE13YYo8WjKaWQshKwsOoDIb2AnVJV4bOjetSjEzJKzBPKm1Ol9H+koC99A4/+w6ecfGp0qif
lOKaqkdM46mFZ35Snxyki1SkCf9z/+rmnFKy/PYzs2kZ/f6GTWS4T6c4t1RBta+AYaBKnJ224wl+
ofppUg4G0mxaUS46bUt7mhlmGBf/o2q4mwfIsB0B7MYcIMgfIG93G5IYYgvVqCFvYF5jb2/IUkNU
22tEkR4ceK7Crx88XFKpPHDSXZmppVi+rbqO6ru+3eMFRSSFaFvCG1MRiYmoWX8B/FHtKqklhOWc
B1NqYGeMUvNlbxBsirtJNuHhEHljO7CE+ZTD/Q8+JyT+FHu0D+OoEEW+zYqDV1q93m3vFS03WDlB
h4yYsc/XxjCA3wEMw0X6/r1f5S5x3FCvsqUQWXdXqrMVaJUau+g+2O6WF1iUPvZVyDSNmCRdRgQj
8HExTv5QZ0JRXMTKoBFPwQV3AnPPmdg7+mc52onzdWbdaPGdICojz6x1h2rq0a++8jrsjcJV0Leq
Gzfj/+PMDpt8W1i4ibsekzb+mQQtIEoau6T7t3KBoI/abxCPd9cjNBj/yeFB03E2O9/1LKllg1a0
gzqe5lJtwwJR+a2PGh1HP+o3WnlQTjaHNfKm3IYTfqsEdxkSodom06lfpAPa7ZKs5owPhXwySd3x
m+7NGT1pPd4s0cxlVmq8XCXbTZes0ASX1EdLkn8myFMic32lxbXT+39SfXI2ndaO+f1znvRE/oUr
jqWoz1z34JJXmoYD8QbMdiyiJrQ1nt2h+to9TJpnhgnKJ1AosP1ZBOF/2nderJydpxMKUr/yB4Zt
SiptKYOM3Bxk1gSuMuZpNtQHueFusgQVHSF/t0h6SLD/7GwumXOLvyrIaOnw6G3aCbpaSkGhBYV6
Ui7II5wyGV/eps1hQCaxJ71nrnG9eh+rXbWX5bvOe2tuTeFnTtziuPR+NZrWgxn3HS7wSzeIJM84
TsipwtMuA283ooRh1fYJBP7s2SnKrG6dr0mCBX6fafEG1T1VPpq3GZhNXwd0VkMLry6wUGTx0QCj
1P0BhDAEBGr8nkCt+Ved3iqxINQOIeCTsoLn7s2MyQJwSTbSfYKxE9+/tZf6eF47p4dIWTRki6g4
GPyYEfVDanVw1+g5sIGFWvdS5Zfx1bAVfDGe88P2PYKkAgtgYD8XpyT3O4UAG/DasYQcuUz/LPIt
e53qWQmacuXVb47aGaDLgzfhR/f5npB0svKurnMkw8ROrkjXolzj+6JC/EpNXkIpmjahtjPwBTml
1wdm0YM5uQckaOLN8h48Aja8imCRrBkKrJVv1urjBSnZUkmTfdyn1Rbu6iVWzDJk1Jxfu1dSt4GG
ieP+1Tdrpvnpk+MnhK75yIUjk/H5LliZs/W0LX+biEaMrK5LU++WCo58aCjngfYaP0DIJhdwsOgg
Cp2TAKizIUxxTSr+OV33gp5R/rc/wENKRQqpo64BfPsiL5fSZkKqBXllY6H8y5N6IppM2fe0LXOO
HJvkUkrlDTPe9NB37qujBSc+eVegbVLm03n9PKe0OrIamfndFWXQbGOaDdWPVvVYBFqdHtNNRuER
Q4PzfHHkEw2tsa59+8PNcGHR3p1UPhwhyxZq4OuK4DaCG+ITy20IH+GbR9ubYxJFIlZNYYQqB8Yt
oUQVUE1voNCg/lWahAVuVenkwBdoG0zMrS3G5uCXKYB96tuSt0BRLiCR0Qa+z5W81ee5MuPnG/9l
pD3rNKyOEh4YqL5mVfLFShFPQ+bfexil22WXR+qOXN8wCSCyL2wJhjUS+yyekWSAGey8NcYBzA/P
r+qP0Fm3nIL22LUJb96dxBjEwkg5gAOSBAof5Z6z5k7xqT6ym5bRc6k9tbcREnRCJTLAKHTNcKAv
StozmYWO/cyueQKqHEdEqO1Y+dVTjXK9c1vfFI0milrNY02UFe0lYYJl9HhzN81ilo/IscGK+psI
AR4rrgQq3Jp61Z9vJW5FBSX70vPKlKnGpqOJeEABDzsPLiZSnoCu/nF/Kj6C8CBs24r20yNSFMQM
B+c9OVHe2wA0SO5yVsNLQgh3DZ777pxVdzn5GWvDtaPZzIB2rJhPYS+cyXavg5woyD9LyaKXbTRO
Vh2KOGlMR2c4HdkWovg5cSAA51aOI0GH3ifkeoakGLeNRILVennkxuvC92rpzAauLj8tp4trckYM
ak6bV63z6wdMOjRRCQ8u+Jj6T9fqOyWpoXi0gXEKMI9n5ptv9+BU/TcixtGj2b0ZNnu6V80wBJZB
vKRdAuGObsVsv+baBL9dQ+NTZ1R7ZhjUvBa2CrgSsh16u1hR5UyU/jIqyb8uKO1gD3tUpHVz2Ivp
ZOpc+UJdQuxBHmZZWApnH+Ur5nygk5LpjXgJxyXBWz05h6mzuAMo8KgYXZiWZvnGnv6vk79GB8UH
35vFxN3jiRR4GW7BFHPNV3V4e9YB4CNqtwgH0wcD4dt55acnUf0QA+RIkjPRAoGfyss/RSS8HeFh
g4OGf1CJbKc5GnA+GQF+h+IPlqk1EX4+nNrGg/pO9wk+mb/JZSKVcah+vMC9Gi4kI8VYX3Y/P2LN
XCxoUae0hxv6nQ8xY6yqU56lk40ABjBYN3RwOAX7o/tbPHfPQXBmJk5q3oow+IZhjd+mb7F8ooB0
HM+2OViibgfCzbkV1x0PpJHi+wLieJcjbhnrc8X9iHRbu1/OUJExFoxmeEoINuikKhlqW+2sMvmv
poBzVSyGXgkimuA48ySmF2EEVsA/PLtVewIRl3Xh04pADIbHBkrHw03pJpy5ctKXgT1JGlAhOFpL
dXixZ8a0RUZ4qyFRz1IUv6SoGOvVFW4quwz/p9zuVa4dqscfhheaNr+oLz8NjNQR9JvpjdJld/AW
GZXwU6mvPxEn/8P7myCLG6YtOLv7+p258wRIclMryWo53DC8jWOHIwyc5Gu7MTMMhtKBSWExHtIq
nXsRI6DqpWoPSH9BupUS5YGvhx2SpeEHPjdJSqiVy4gEeLH6aChLMYsrx6E3w+0n459PJ9Dt6KvL
taT4KjKeCWweu9FOb6JTUflx0bZkEcOespASt0uS1yYpjDlLtEx5Qbp2E1fLAvAzrK3d0A6HGl9S
IAFJrIrgNHN+KOqZBIQSaCXoyyGVDFouuFsAwAqkQKCc2x7/01dbonjdjg8INp80mCev0jUUz5ra
Kf/jhwzkMDTFGhKAJPk1NPDEdKpcVXQaoghgGFRWw73A5MnmBk4/ZL8iv1LhQpBAQfwzidZ0yODL
r4YSExcUw/0wcKPaCJela4DG55U1HRVa7stjNhbAMZAdcjmmi2CI6r1XqkmCb4muar1+2xLhRph3
aH3d74adRJEBHiqi/dKxeUTm97cWhAv1rqT9Vb0r3cRakDiFm0IMV5Svv5Uvt3g+oj5LPlvu+zPZ
HwQmH8uaJSMXKNw49ksh/h4Z51klMbsCUrtVhvkBYZlPesMHHr6ytgaju8LMguJYdCZ+8q+utFUG
1Yt7GNbJzPd2MMi7DEwejrYXcomZFDcP/cL7ckreBmpOT8nYTE+ER0K1FZnMNrhnTWJBd6FcpyS5
58ZpDsuQS9XwEXQ+PuRHvwUAWA/ZM22IN3D88vhuDOui7hQEcxY2rSJosWM3eTtHESUYZ5lWs5d/
fhjUQegiKi14eZqz6dgjS2FQBWn1xL1sRvdRikxQj8lq2DGwgFtIvxAwNYCnJx9Ovvbw3iWqJ8CU
Z/OGYSGV5ze0+2AbQSIXMJoMngbz/a3/cqZ+R0sIz5BljO2srUE3cnqIk3BXD2tHBy/29Omtz7jf
sapggW0xpVPj+8mmbQGSnxE230YdEFCvvbO/F3LGDIIj2x5aKkQqRbHQJvxfbKDJ81bwJ5SQlyDv
j6goB5GMFIw0+LIy0tpIyVVla8CFnYiLWSZnTz5aID50oejXBH0hK88yc7zZW2dOV/LXB8fro4PN
l59IoeaT6/dofJkArHplSTUakwPV5m86ZI9kXBl2nmXOFHw22mP/LQPe1q47IV5tNSTx2X0Wh/Mm
31Pdr/a2ktxmD3D0dkIB7pIeosMqQ6TvqgGte62jnubvJatLv7MuvEfrX8Dk7/APUT/+QbXb/6G0
6SaCf5g+pS6Le7iQk7eBNx6Nqu6eXFtLrC3pD+vOcl6meeC55kunnr/FiC0JHZXtYH6kA19kYK4z
AkhgIu/8DzMLHSrpxzAABTTdO0QWerIoZtgop98TTwwGQQA4yP9OOmU9jLDz3XAOFF5cxdmJ0/ID
cs3rmcUFE+zGV+viuS+SDhYotKqupVlleKqi+mhQyFd65kvgqChbRttHJt8hTae9C4TKn/hkwtrp
JVIv11zEeIJSntaMb3klqPZdNWqRXEIB6Fiw7a6OdDugOP/Bzfw2p+D4eKPh8XhzJI2VEDOdw7EI
fMpJEIlqJAPaWUhiTQm4tBQqI2CblI8wZ4uqfoTTcjZ20kgBI7r+RGY9lz3UGqXchDUtv93dALCh
l0O4ejQgUkhQHZ0ZkyoOQgbYwWYalR7ZvdJ2SWX+4SeR1kPFOmkuV23pBvn5YSehbdndRNXxG0Iy
DHJorOm045d9QoYBJ5bki21fjrAZGcEIFCAbP0Nfa9KKJ24NDxZdlKgNPOu4DJZhi5xtz4+K30KP
h09xQjRtnwUgwGk6U71hRZed3b0NawXH4DUVtg20BKEDn5JXhAQAWyIYCLhWbcd7yvHIt0r8al0F
1ui41HjsiiPdUHNBH1H6tcRim+X+b+R2oQB1HxG+UQBSko0nklVb4k2FkNogtWYMwlPu9CGsLy0+
l6vhQ1I8Oal+htIt2kgPeNoPhzKRwkFdBTliMaiFjfDRQdDejOgVDEuXVwP53b5qiY1moK9z76KV
1e0+vslqNlSaOn7vgqdLwSBxZrp0L5CZkFWsXROuOIxK6CDKDwrV+F1osfbgyFBNbQPoNRPCkpQU
h2AEr1A8Ud9WzhnRoJeYvAOthum9+8va5S0p1n7nqyD5ME6/sf5Crao8q9MMIFz5OYC66CgT55x3
Z3LBcG1AQGK5xSA2kUzRlHtPo8rZCStl1orEFw3KudifVlJzWM3f
`protect end_protected
