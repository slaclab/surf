------------------------------------------------------------------------------
-- This file is part of 'SLAC JESD204b Core'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'SLAC JESD204b Core', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

use work.StdRtlPkg.all;
use work.AxiLitePkg.all;
use work.Jesd204bPkg.all;

--------------------------------------------------------------------------------
entity DescrambleTb is

end entity;
--------------------------------------------------------------------------------

architecture Bhv of DescrambleTb is
   -----------------------------
   -- Port Signals 
   -----------------------------
   constant CLK_PERIOD_C : time := 10 ns;
   constant TPD_C        : time := 1 ns;

   -- Clocking
   signal clk_i : sl := '0';
   signal rst_i : sl := '0';

   -----------------------------
   -- Port Signals 
   -----------------------------
   signal subClass_i   : sl := '1';
   signal sysRef_i     : sl := '0';
   signal clearErr_i   : sl := '0';
   signal enable_i     : sl := '1';
   signal replEnable_i : sl := '1';
   signal scrEnable_i  : sl := '1';
   signal r_jesdGtRx   : jesdGtRxLaneType;
   signal lmfc_i       : sl := '0';
   signal nSyncAny_i   : sl := '1';
   signal nSyncAnyD1_i : sl := '0';
   signal nSync_o      : sl;
   signal dataValid_o  : sl;
   signal sampleData_o : slv((GT_WORD_SIZE_C*8)-1 downto 0);
   signal status_o     : slv((RX_STAT_WIDTH_C)-1 downto 0);

   signal s_sysrefRe : sl;
   signal s_lmfc     : sl;

   type dataArrayType is array (0 to 412) of slv(31 downto 0);
   type charArrayType is array (0 to 412) of slv(3 downto 0);

   signal dataArray : dataArrayType := (
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"10111100101111001011110010111100",
      b"00011100101111001011110010111100",
      b"00000100000000110000001000000001",
      b"00001000000001110000011000000101",
      b"00001100000010110000101000001001",
      b"00010000000011110000111000001101",
      b"00010100000100110001001000010001",
      b"00011000000101110001011000010101",
      b"00011100000110110001101000011001",
      b"00100000000111110001111000011101",
      b"00100100001000110010001000100001",
      b"00101000001001110010011000100101",
      b"00101100001010110010101000101001",
      b"00110000001011110010111000101101",
      b"00110100001100110011001000110001",
      b"00111000001101110011011000110101",
      b"00111100001110110011101000111001",
      b"00011100011111000011111000111101",
      b"00000000000000000000000010011100",
      b"00000000000111110000000110000000",
      b"00000000001000000010111100001111",
      b"01010000010000010000000000000000",
      b"01010100010100110101001001010001",
      b"01011000010101110101011001010101",
      b"01011100010110110101101001011001",
      b"01100000010111110101111001011101",
      b"01100100011000110110001001100001",
      b"01101000011001110110011001100101",
      b"01101100011010110110101001101001",
      b"01110000011011110110111001101101",
      b"01110100011100110111001001110001",
      b"01111000011101110111011001110101",
      b"01111100011110110111101001111001",
      b"00011100011111000111111001111101",
      b"10000100100000111000001010000001",
      b"10001000100001111000011010000101",
      b"10001100100010111000101010001001",
      b"10010000100011111000111010001101",
      b"10010100100100111001001010010001",
      b"10011000100101111001011010010101",
      b"10011100100110111001101010011001",
      b"10100000100111111001111010011101",
      b"10100100101000111010001010100001",
      b"10101000101001111010011010100101",
      b"10101100101010111010101010101001",
      b"10110000101011111010111010101101",
      b"10110100101100111011001010110001",
      b"10111000101101111011011010110101",
      b"10111100101110111011101010111001",
      b"00011100011111001011111010111101",
      b"11000100110000111100001011000001",
      b"11001000110001111100011011000101",
      b"11001100110010111100101011001001",
      b"11010000110011111100111011001101",
      b"11010100110100111101001011010001",
      b"11011000110101111101011011010101",
      b"11011100110110111101101011011001",
      b"11100000110111111101111011011101",
      b"11100100111000111110001011100001",
      b"11101000111001111110011011100101",
      b"11101100111010111110101011101001",
      b"11110000111011111110111011101101",
      b"11110100111100111111001011110001",
      b"11111000111101111111011011110101",
      b"11111100111110111111101011111001",
      b"01101100011111001111111011111101",
      b"01101101110001110000000100101110",
      b"01110001000010010000010010001111",
      b"11001010010101100100111100010100",
      b"10011001111100001101011111011010",
      b"11101011000101110011111100001000",
      b"00000111111101110001001001011001",
      b"01110011000111000111101100001011",
      b"11100100010101010100001001101011",
      b"11000001110010010011001111010110",
      b"00000000011011111110110010011111",
      b"00011001001111010110100001111101",
      b"11100011110100000011110010100011",
      b"10101100100001110010000111001001",
      b"01101100101010111000000100111101",
      b"01100001111111110000001111011101",
      b"10001001110101110010111100100010",
      b"10100100100100100101110111000010",
      b"11001001001101111011000001110001",
      b"10100011110000001101110010101101",
      b"10101010100111111010000010110011",
      b"00010000011101001001010001100001",
      b"01011110010010110000100100010010",
      b"10001100011011101010111010011010",
      b"11101011110100000100000001010110",
      b"00001101110000000001000111010101",
      b"11110010100101110100010010110010",
      b"11110010101011110100010001000000",
      b"11111001110011010100011111010000",
      b"01100000011000110111110010011001",
      b"10011000010010000010100001101100",
      b"11110100011111010011101010011111",
      b"10001101111000000101000100100010",
      b"11111101001000010100011001111000",
      b"00110110011101100110010111100101",
      b"10100110010101101101110100010001",
      b"11101001111011101011111111011101",
      b"00101101000011010001111001111000",
      b"01111010011010111000011100011111",
      b"01010000011111000111010001100100",
      b"01011100101001001000100100111110",
      b"10100010010001101010001111101100",
      b"10111110100010101010011010110010",
      b"00000111000111111110110100001110",
      b"01110100010101110111101001101001",
      b"10000001111110100101001111011000",
      b"00001000100111000110111100110000",
      b"10111000011011010101100001100001",
      b"01111010101011011111100001001000",
      b"01011000101011010111011111000001",
      b"11110001111101011011101111011111",
      b"11001010010001000100111100010111",
      b"10011111110111011101011010101001",
      b"10011110011110000010100111100110",
      b"10000100100011000010110100111000",
      b"01001111001000110111000100000100",
      b"11011111000000011100100111110011",
      b"10010000100011011010101100110010",
      b"01011111001001010000100100000001",
      b"10011111001100111010100111111110",
      b"10011000010100000010100010010000",
      b"11110001110111100011101111010100",
      b"11000101111111100100110111011000",
      b"01011001111000001111011100100111",
      b"11101100010000001011111001101101",
      b"01100111111001110000001010100101",
      b"11110100010010010011101001101000",
      b"10000100011001110101001010011000",
      b"01001000011001110111000001100000",
      b"10111001001011111101100001111000",
      b"01100100101101111111110111000000",
      b"11000101001000100011001010000110",
      b"01010110011000011111010111100111",
      b"00100000010100011001110001101000",
      b"10010000100101101010101111001010",
      b"01011010100100110000100001001011",
      b"11010010100101111011010001000011",
      b"01110011111001011000010001011101",
      b"11100100010000110100001001101110",
      b"11000110101111010011001010111010",
      b"01101110101101001111111010111110",
      b"01001101000101000000111010001010",
      b"11111100011000011100011001100011",
      b"00101001000110110110000001110010",
      b"00101100010011111001111001101010",
      b"01100101000010101000001010001011",
      b"11011010011101110011011100011010",
      b"11010110011100011011010100011110",
      b"00100111000111111001110100001000",
      b"11110101000010011011101001110110",
      b"10011011001101110101011100000001",
      b"11001001001010110011000010000010",
      b"10100100101001011101110111000010",
      b"11000011001111101011001111111100",
      b"00101010100101011110000010110110",
      b"00010011110001101001010001010111",
      b"01101010100100000000000010110101",
      b"00010011110010000001010001010011",
      b"01101001001001110000000010000000",
      b"00100110011111000001110111100111",
      b"11100101111011011011110100100000",
      b"11011111111101100011011001011110",
      b"10010011000110011010101100000000",
      b"01100101001011110000001001110100",
      b"11010100101111110011010111000110",
      b"00000110100001001001001010110001",
      b"01100111001100010111110100000000",
      b"11111010101000100011100010111000",
      b"01011011001010000111011111111000",
      b"11001101111011001011000111011110",
      b"11111110101010001100011001000001",
      b"00001001110011010110111111010100",
      b"10100001001111000101110010000110",
      b"10000000010101011010110010010100",
      b"00010001110100010110101111010100",
      b"01000100101110100000110111000101",
      b"01000110101011111111001010111001",
      b"01101000100111001111111111001100",
      b"00111000010000000001100001101111",
      b"01110110100111011111101010110111",
      b"10100000010011000101110001101010",
      b"10010101000011001010101010001100",
      b"00011011000010100001011100001110",
      b"11000010011101100011001100010011",
      b"00110110010000101110010100010000",
      b"10101110101001111101111010111010",
      b"01001011001011111000111111111010",
      b"10001100101111111101000111000100",
      b"11100111110011110100001010101010",
      b"11111010101100110011100010111010",
      b"01011100011011110111011010011110",
      b"10101010101011101010000001001001",
      b"00011001110000011001011111010101",
      b"11100011110001110011110010101100",
      b"10101010101110000010000010111001",
      b"00011110100111011001011010110001",
      b"10000000010101100010110001100000",
      b"00010001111010000110101111011010",
      b"01001110101110000000111001000110",
      b"11001111111010101100111010100001",
      b"11010110100110111100101001001001",
      b"00100001001001101001110001111111",
      b"10000111000100011010110111110000",
      b"01110110100110010111101001000001",
      b"10100000010001010101110001101010",
      b"10010110100011011010101010110100",
      b"00100111001110110001110100000111",
      b"11111001001001001011100010000111",
      b"01100111000011010111110111110000",
      b"11110011000110100011101100001011",
      b"11100110101011100100001001000000",
      b"11101001110001010011111111010110",
      b"00100010100011000001110010110001",
      b"10110111001000011010010100000010",
      b"10111110010100001101100111101110",
      b"00001000100100101110111111001011",
      b"10111011111011000101100001011100",
      b"01000111111001011111001001011100",
      b"01110100010011101111101001101100",
      b"10000101001100010101001010000001",
      b"01010000011001110111010010011100",
      b"01011000011011001000100001100101",
      b"11111011110101011011100001000110",
      b"01001100100000010111000111001110",
      b"11101101111110001100000100100000",
      b"01111000101000100000011100111000",
      b"01110010011111100111101111100010",
      b"11110101110100000100010100101001",
      b"10010101111111000101010111011000",
      b"00011000100111010001011100110111",
      b"11111000010101110011100001101010",
      b"01110000101010010111101111000100",
      b"11010000101100110100101111000100",
      b"01010101001011011000101010000110",
      b"00010100101101101001010111000000",
      b"00000100011100000001001010011111",
      b"01001110010101010111000100010000",
      b"11001001110010001100111111010010",
      b"10100000011011111101110010010111",
      b"10011010101110101010100001000110",
      b"11011110101010100011011010111111",
      b"10001001111000001010111111011101",
      b"10101100010010100101111001101100",
      b"01100100010000111000001010010010",
      b"11000110101010000011001010111101",
      b"01101000101110001111111111000001",
      b"00110111110101100001101010101110",
      b"10111101111110001101100111011111",
      b"00111000101100101110011100111100",
      b"01110100011111111111101010011000",
      b"10001100100000100101000100110001",
      b"11101101110011010100000100101011",
      b"01110000011010010000010010011100",
      b"11011011110000100100100001011010",
      b"11001010101100111011000010111010",
      b"10011101001001101101011010000001",
      b"10110100100101100010010111001000",
      b"10001011111000101101000001011000",
      b"10000111110101000101001001010001",
      b"01111101110110000111100111010110",
      b"00110111001000110110010111111001",
      b"10111110011010101101100111100000",
      b"00000011110010111110110001010011",
      b"00101001000101010110000010001011",
      b"00101111110101111001111001010000",
      b"01011100101111111000100111000111",
      b"10100111110000001010001010101110",
      b"11111011110100001011100010101011",
      b"01001111001001010111000111111001",
      b"11011111000011101100100111110000",
      b"10010010010011111010101100010010",
      b"01111101001111100000011010000100",
      b"00110011110100100110010010100010",
      b"11101111000100101100000111110100",
      b"01010111110100100000101001010110",
      b"00111101111110001001100111011100",
      b"00111000100110101110011100111101",
      b"01111000010101001111100001101011",
      b"01110001110101000111101111010100",
      b"11000101110010010100110111010000",
      b"01010000011010001111010010011110",
      b"01011010100110001000100001001000",
      b"11010001000001011011010001110011",
      b"01001000100111101000111100110000",
      b"10111000011100101101100001100000",
      b"01111111001000011111100100000101",
      b"00011111000110010110100111111111",
      b"10010101001010010010101001111010",
      b"00010100101101110001010111000101",
      b"00000100011101110001001010011010",
      b"01001110010100010111000100010111",
      b"11001000101011111100111111000000",
      b"10110000101001001101101111000110",
      b"11010010011110011100101111100101",
      b"01110100101011011000010100111111",
      b"10000000100111010101001111011011",
      b"00011000011011010110100001100010",
      b"11111011110110110011100001011110",
      b"01001111000001010111000111110110",
      b"11010001110100011100101100101111",
      b"01000100101101111000110111000101",
      b"01000101001110101111001010000011",
      b"01010010101100101111010010111001",
      b"01111101001101111000011010000011",
      b"00110000011011010110010010011111",
      b"11011011110111101100100001010111",
      b"11001111000110101011000111110110",
      b"11010101000101111100101001110010",
      b"00011111110001101001011001010111",
      b"10011010100100000010100010110001",
      b"11010010101001100011010001000000",
      b"01111011001011001000011111111111",
      b"01001100100111110111000111001001",
      b"11101001000011001100000001110100",
      b"00101010011011100001111100011110",
      b"00010010101000001001010001000110",
      b"01111011000111010000011111110010",
      b"01000100011011010111001001100110",
      b"01001011111001011111000001011101",
      b"10000101001011001101001001111010",
      b"01010100101010100111010111000001",
      b"00000000100100001001001111001010",
      b"00011010100110000110100001001001",
      b"11010000010001100011010001100101",
      b"01010110100101011000101010110000",
      b"00100010100111111001110001001001",
      b"10110000011111111010010001100110",
      b"11011101110000001100100100101100",
      b"10110011110001011010010010101001",
      b"11101010101111101100000010110000",
      b"00011111110011010001011010101111",
      b"10011001000111000010100010001110",
      b"11101101001110010011111001111000",
      b"01110001000110110000010010001100",
      b"11001101000111010100111001110100",
      b"11111101001001011100011001111001",
      b"00110111000101100110010111110101",
      b"10110110100001011101101001001100",
      b"10100100100001011101110100110000",
      b"11001101111110011011000100101110",
      b"11111000100111101100011100110111",
      b"01111000010001000111100001101101",
      b"01110110100010000111101010111000",
      b"10100101111010000101110100100001",
      b"11011111111100011011011001010010",
      b"10010000101100011010101100111000",
      b"01010110100010010000101010111000",
      b"00100110010011001001110100010101",
      b"11101101001110111011111010000111",
      b"01110010101010000000010010111111",
      b"11111001110000100100011111011010",
      b"01100011110111000111110010101000",
      b"10101111001011110010000111111100",
      b"01011101110010111000100111010010",
      b"10110001000100101010010010001011",
      b"11001110101010111100111001000010",
      b"11001000100110101100111111001001",
      b"10111001000100001101100001110101",
      b"01101111111111101111111001011110",
      b"01010000100101000000101100110100",
      b"01011011110011011000100001010101");


   signal charArray : charArrayType := (
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"1111",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"1100",
      b"0001",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"1100",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"1100",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0100",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0001",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0100",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0001",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000",
      b"0000");

begin  -- architecture Bhv

   -- Generate clocks and resets
   DDR_ClkRst_Inst : entity work.ClkRst
      generic map (
         CLK_PERIOD_G      => CLK_PERIOD_C,
         RST_START_DELAY_G => 1 ns,     -- Wait this long into simulation before asserting reset
         RST_HOLD_TIME_G   => 1000 ns)  -- Hold reset for this long)
      port map (
         clkP => clk_i,
         clkN => open,
         rst  => rst_i,
         rstL => open);

   -----------------------------
   -- component instantiation 
   -----------------------------
   JesdRxLane_INST : entity work.JesdRxLane
      generic map (
         TPD_G => TPD_C)
      port map (
         devClk_i     => clk_i,
         devRst_i     => rst_i,
         subClass_i   => subClass_i,
         sysRef_i     => s_sysrefRe,
         clearErr_i   => clearErr_i,
         enable_i     => enable_i,
         replEnable_i => replEnable_i,
         scrEnable_i  => scrEnable_i,
         status_o     => status_o,
         r_jesdGtRx   => r_jesdGtRx,
         lmfc_i       => s_lmfc,
         nSyncAny_i   => nSyncAny_i,
         nSyncAnyD1_i => nSyncAnyD1_i,
         nSync_o      => nSync_o,
         dataValid_o  => dataValid_o,
         sampleData_o => sampleData_o);


   -- LMFC period generator aligned to SYSREF input
   LmfcGen_INST : entity work.LmfcGen
      generic map (
         TPD_G => TPD_C)
      port map (
         clk        => clk_i,
         rst        => rst_i,
         nSync_i    => '1',
         sysref_i   => sysRef_i,
         sysrefRe_o => s_sysrefRe,
         lmfc_o     => s_lmfc
         );

   StimuliProcess : process

      variable v_data : slv(31 downto 0);
      variable v_char : slv(3 downto 0);

   begin

      r_jesdGtRx.data    <= x"bcbcbcbc";
      r_jesdGtRx.dataK   <= (others => '1');
      r_jesdGtRx.dispErr <= (others => '0');
      r_jesdGtRx.decErr  <= (others => '0');
      r_jesdGtRx.rstDone <= '1';

      wait until rst_i = '0';
      wait for CLK_PERIOD_C*200;

      -- Apply sysref
      sysRef_i <= '1';
      wait for CLK_PERIOD_C*50;
      sysRef_i <= '0';

      -- Run data
      for i in 0 to 412 loop
         r_jesdGtRx.data  <= dataArray(i);
         r_jesdGtRx.dataK <= charArray(i);
         wait for CLK_PERIOD_C*1;
      end loop;

   end process StimuliProcess;

end architecture Bhv;
