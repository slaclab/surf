-------------------------------------------------------------------------------
-- Title      : Heartbeat
-------------------------------------------------------------------------------
-- File       : Heartbeat.vhd
-- Author     : Benjamin Reese  <bareese@slac.stanford.edu>
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 2013-04-30
-- Last update: 2014-10-27
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: Heartbeat LED output
-------------------------------------------------------------------------------
-- Copyright (c) 2013 SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

use work.StdRtlPkg.all;

entity Heartbeat is
   generic (
      TPD_G        : time   := 1 ns;
      USE_DSP48_G  : string := "no";
      PERIOD_IN_G  : real   := 6.4E-9;   --units of seconds
      PERIOD_OUT_G : real   := 1.0E-0);  --units of seconds
   port (
      clk : in  sl;
      rst : in  sl := '0';
      o   : out sl);
end entity Heartbeat;

architecture rtl of Heartbeat is
   
   constant CNT_MAX_C  : natural := getTimeRatio(PERIOD_OUT_G, (2.0 * PERIOD_IN_G));
   constant CNT_SIZE_C : natural := bitSize(CNT_MAX_C);

   type RegType is record
      cnt : slv(CNT_SIZE_C-1 downto 0);
      o   : sl;
   end record RegType;

   constant REG_INIT_C : RegType := (
      cnt => (others => '0'),
      o   => '0');

   signal r   : RegType := REG_INIT_C;
   signal rin : RegType;

   -- Attribute for XST
   attribute use_dsp48      : string;
   attribute use_dsp48 of r : signal is USE_DSP48_G;
   
begin

   -- USE_DSP48_G check
   assert ((USE_DSP48_G = "yes") or (USE_DSP48_G = "no") or (USE_DSP48_G = "auto") or (USE_DSP48_G = "automax"))
      report "USE_DSP48_G must be either yes, no, auto, or automax"
      severity failure;


   comb : process (r) is
      variable v : RegType;
   begin
      v := r;

      v.cnt := r.cnt + 1;
      if (r.cnt = CNT_MAX_C) then
         v.cnt := (others => '0');
         if (r.o = '1') then
            v.o := '0';
         else
            v.o := '1';
         end if;
      end if;

      if (rst = '1') then
         v := REG_INIT_C;
      end if;

      rin <= v;
      o   <= r.o;
      
   end process comb;

   seq : process (clk) is
   begin
      if (rising_edge(clk)) then
         r <= rin after TPD_G;
      end if;
   end process seq;

end architecture rtl;
