-------------------------------------------------------------------------------
-- Title      : AXI Stream DMA Write
-- Project    : General Purpose Core
-------------------------------------------------------------------------------
-- File       : AxiStreamDmaWrite.vhd
-- Author     : Ryan Herbst, rherbst@slac.stanford.edu
-- Created    : 2014-04-25
-- Last update: 2014-05-05
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description:
-- Block to transfer a single AXI Stream frame into memory using an AXI
-- interface.
-------------------------------------------------------------------------------
-- Copyright (c) 2014 by Ryan Herbst. All rights reserved.
-------------------------------------------------------------------------------
-- Modification history:
-- 04/25/2014: created.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

use work.StdRtlPkg.all;
use work.AxiStreamPkg.all;
use work.AxiPkg.all;
use work.AxiDmaPkg.all;

entity AxiStreamDmaWrite is
   generic (
      TPD_G            : time                := 1 ns;
      AXI_READY_EN_G   : boolean             := false;
      AXIS_CONFIG_G    : AxiStreamConfigType := AXI_STREAM_CONFIG_INIT_C;
      AXI_CONFIG_G     : AxiConfigType       := AXI_CONFIG_INIT_C;
      AXI_BURST_G      : slv(1 downto 0)     := "01";
      AXI_CACHE_G      : slv(3 downto 0)     := "1111";
      AXI_ALIGN_G      : boolean             := true
   );
   port (

      -- Clock/Reset
      axiClk          : in  sl;
      axiRst          : in  sl;

      -- DMA Control Interface
      dmaReq          : in  AxiWriteDmaReqType;
      dmaAck          : out AxiWriteDmaAckType;

      -- Streaming Interface 
      axisMaster      : in  AxiStreamMasterType;
      axisSlave       : out AxiStreamSlaveType;

      -- AXI Interface
      axiWriteMaster  : out AxiWriteMasterType;
      axiWriteSlave   : in  AxiWriteSlaveType;
      axiWriteCtrl    : in  AxiCtrlType
   );
end AxiStreamDmaWrite;

architecture structure of AxiStreamDmaWrite is

   constant DATA_BYTES_C : integer := ite(AXIS_CONFIG_G.TDATA_BYTES_C < AXI_CONFIG_G.DATA_BYTES_C,
                                          AXIS_CONFIG_G.TDATA_BYTES_C,
                                          AXI_CONFIG_G.DATA_BYTES_C);

   type StateType is (S_IDLE_C, S_FIRST_C, S_NEXT_C, S_DATA_C, S_LAST_C, S_DUMP_C, S_WAIT_C, S_DONE_C);

   type RegType is record
      state    : StateType;
      dmaReq   : AxiWriteDmaReqType;
      dmaAck   : AxiWriteDmaAckType;
      shift    : slv(3  downto 0);
      shiftEn  : sl;
      last     : sl;
      reqCount : slv(31 downto 0);
      ackCount : slv(31 downto 0);
      wMaster  : AxiWriteMasterType;
      slave    : AxiStreamSlaveType;
   end record RegType;

   constant REG_INIT_C : RegType := (
      state    => S_IDLE_C,
      dmaReq   => AXI_WRITE_DMA_REQ_INIT_C,
      dmaAck   => AXI_WRITE_DMA_ACK_INIT_C,
      shift    => (others=>'0'),
      shiftEn  => '0',
      last     => '0',
      reqCount => (others=>'0'),
      ackCount => (others=>'0'),
      wMaster  => AXI_WRITE_MASTER_INIT_C,
      slave    => AXI_STREAM_SLAVE_INIT_C
      );

   signal r             : RegType := REG_INIT_C;
   signal rin           : RegType;
   signal selReady      : sl;
   signal selPause      : sl;
   signal intAxisMaster : AxiStreamMasterType;
   signal intAxisSlave  : AxiStreamSlaveType;

begin

   -- Stream Shifter
   U_AxiStreamShift : entity work.AxiStreamShift
      generic map (
         TPD_G         => TPD_G,
         AXIS_CONFIG_G => AXIS_CONFIG_G
      ) port map (
         axisClk     => axiClk,
         axisRst     => axiRst,
         axiStart    => r.shiftEn,
         axiShiftDir => '0',
         axiShiftCnt => r.shift,
         sAxisMaster => axisMaster,
         sAxisSlave  => axisSlave,
         mAxisMaster => intAxisMaster,
         mAxisSlave  => intAxisSlave
      );

   -- Determine handshaking mode
   selReady <= axiWriteSlave.wready when AXI_READY_EN_G else '1';
   selPause <= '0'                  when AXI_READY_EN_G else axiWriteCtrl.pause;

   comb : process (axiRst, r, intAxisMaster, axiWriteSlave, dmaReq, selReady, selPause ) is
      variable v     : RegType;
      variable bytes : slv(3 downto 0);
   begin
      v := r;

      -- Init
      v.slave.tReady    := '0';
      v.wMaster.awvalid := '0';
      v.wMaster.bready  := '1';
      v.shiftEn         := '0';

      -- Count number of bytes in return data
      bytes := onesCount(intAxisMaster.tKeep);

      -- Count acks
      if axiWriteSlave.bvalid = '1' then
         v.ackCount := r.ackCount + 1;

         if axiWriteSlave.bresp /= "00" then
            v.dmaAck.writeError := '1';
         end if;
      end if;

      -- State machine
      case r.state is

         -- IDLE
         when S_IDLE_C =>
            v.wMaster  := AXI_WRITE_MASTER_INIT_C;
            v.slave    := AXI_STREAM_SLAVE_INIT_C;
            v.reqCount := (others=>'0');
            v.ackCount := (others=>'0');
            v.shift    := (others=>'0');
            v.last     := '0';

            v.dmaAck                     := AXI_WRITE_DMA_ACK_INIT_C;
            v.dmaReq                     := dmaReq;
            v.dmaReq.address(2 downto 0) := "000";

            if AXI_ALIGN_G then
               v.shift := '0' & dmaReq.address(2 downto 0);
            end if;

            -- Start 
            if dmaReq.request = '1' then
               v.shiftEn := '1';
               v.state   := S_FIRST_C;
            end if;

         -- First
         when S_FIRST_C =>

            -- Determine transfer size to align all transfers to 128 byte boundaries
            -- This initial alignment will ensure that we never cross a 4k boundary
            v.wMaster.awaddr := r.dmaReq.address;
            v.wMaster.awlen  := x"F" - r.dmaReq.address(6 downto 3);

            -- There is enough room in the FIFO for a burst and address is ready
            if selPause = '0' and axiWriteSlave.awready = '1' then
               v.wMaster.awvalid := '1';
               v.reqCount        := r.reqCount + 1;
               v.state           := S_DATA_C;
            end if;

         -- Next Write
         when S_NEXT_C =>
            v.wMaster.awaddr := r.dmaReq.address;
            v.wMaster.awlen  := x"F";

            -- There is enough room in the FIFO for a burst and address is ready
            if selPause = '0' and axiWriteSlave.awready = '1' then
               v.wMaster.awvalid := '1';
               v.reqCount        := r.reqCount + 1;
               v.state           := S_DATA_C;
            end if;
             
         -- Move Data
         when S_DATA_C =>

            -- Assert ready when incoming is ready and we are not done
            v.slave.tReady := selReady and (not r.last);

            -- Advance pipeline when incoming data is valid and outbound is ready
            -- or we have not yet asserted valid
            if intAxisMaster.tValid = '1' and (selReady = '1' or r.wMaster.wvalid = '0') then
               v.wMaster.wdata((DATA_BYTES_C*8)-1 downto 0) := intAxisMaster.tData((DATA_BYTES_C*8)-1 downto 0);
               v.wMaster.wvalid := intAxisMaster.tValid;

               -- Address and size increment
               v.dmaReq.address := r.dmaReq.address + 8;
               v.dmaAck.size    := r.dmaAck.size + bytes;

               -- First in packet
               if r.dmaAck.size = 0 then
                  v.dmaAck.dest := intAxisMaster.tDest;
                  v.dmaAck.id   := intAxisMaster.tId;
                  v.dmaAck.firstUser(AXIS_CONFIG_G.TUSER_BITS_C-1 downto 0) := 
                     axiStreamGetUserField(AXIS_CONFIG_G,intAxisMaster,conv_integer(r.shift));
               end if;

               -- Last in packet
               if intAxisMaster.tLast = '1' then
                  v.dmaAck.lastUser(AXIS_CONFIG_G.TUSER_BITS_C-1 downto 0) := axiStreamGetUserField(AXIS_CONFIG_G,intAxisMaster);
                  v.last := '1';
               end if;

               -- Last in transfer
               if r.wMaster.awlen = 0 then
                  v.wMaster.wlast := '1';
                  v.state         := S_LAST_C;
               else
                  v.wMaster.wlast := '0';
                  v.wMaster.awlen := r.wMaster.awlen - 1;
               end if;

               -- Write strobe
               v.wMaster.wstrb(DATA_BYTES_C-1 downto 0) := intAxisMaster.tKeep(DATA_BYTES_C-1 downto 0);

               -- Detect overflow
               if r.dmaAck.overflow = '1' or bytes > r.dmaReq.maxSize then
                  v.dmaAck.overflow := '1';
                  v.wMaster.wstrb   := (others=>'0');
               else
                  v.dmaReq.maxSize := r.dmaReq.maxSize - bytes;
               end if;

               -- Done
               if r.last = '1' then
                  v.wMaster.wstrb := (others=>'0');
               end if;
            end if;

         -- Last Trasfer Of A Burst Data
         when S_LAST_C =>
            if selReady = '1' then
               if r.last = '1' then
                  v.state := S_WAIT_C;
               elsif r.dmaAck.overflow = '1' or r.dmaAck.writeError = '1' then
                  v.state := S_DUMP_C;
               else
                  v.state := S_NEXT_C;
               end if;
               v.wMaster.wvalid := '0';
            end if;

         -- Dump remaining data
         when S_DUMP_C =>
            v.slave.tReady := '1';

            if intAxisMaster.tLast = '1' then
               v.state := S_WAIT_C;
            end if;

         -- Wait for acks
         when S_WAIT_C =>
            if r.ackCount >= r.reqCount then
               v.state       := S_DONE_C;
               v.dmaAck.done := '1';
            end if;

         -- Done
         when S_DONE_C =>
            if dmaReq.request = '0' then
               v.dmaAck.done := '0';
               v.state       := S_IDLE_C;
            end if;

         when others =>
            v.state := S_IDLE_C;
      end case;

      if (axiRst = '1') then
         v := REG_INIT_C;
      end if;

      -- Constants
      v.wMaster.awsize  := conv_std_logic_vector(AXI_CONFIG_G.DATA_BYTES_C-1,3);
      v.wMaster.awburst := AXI_BURST_G;
      v.wMaster.awcache := AXI_CACHE_G;
      v.wMaster.awlock  := "00";   -- Unused
      v.wMaster.awprot  := "000";  -- Unused
      v.wMaster.awid    := (others=>'0');
      v.wMaster.wid     := (others=>'0');

      rin <= v;

      dmaAck         <= r.dmaAck;
      intAxisSlave   <= v.slave;
      axiWriteMaster <= r.wMaster;

   end process comb;

   seq : process (axiClk) is
   begin
      if (rising_edge(axiClk)) then
         r <= rin after TPD_G;
      end if;
   end process seq;

end structure;
